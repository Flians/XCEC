//
// Conformal-LEC Version 20.10-d207 (02-Sep-2020)
//
module top(RIdec64b8_720,RIbc62af0_23,RIbc62a78_22,RIbc62a00_21,RIbc62988_20,RIbc62910_19,RIbc62898_18,RIbc62820_17,RIbc627a8_16,
        RIbc62730_15,RIbc626b8_14,RIbc62640_13,RIdec37b8_688,RIfc8daa0_6634,RIdec0ab8_656,RIfc56348_6003,RIdebddb8_624,RIdebb0b8_592,RIdeb83b8_560,
        RIfc98798_6757,RIdeb29b8_496,RIfcbd098_7173,RIdeafcb8_464,RIfc8dc08_6635,RIdeacb80_432,RIdea6280_400,RIde9f980_368,RIfcd6868_7463,RIfc8ded8_6637,
        RIfc7dd80_6454,RIfc56618_6005,RIde92e10_306,RIde8f300_288,RIde8b160_268,RIde86fc0_248,RIde82ad8_227,RIfc8e040_6638,RIfcd96d0_7496,RIfca1e10_6864,
        RIfcbd200_7174,RIe16c5c0_2610,RIe16a298_2585,RIe168ab0_2568,RIe1664b8_2541,RIe1637b8_2509,RIee37f00_5095,RIe160ab8_2477,RIfc8ea18_6645,RIe15ddb8_2445,
        RIe1583b8_2381,RIe1556b8_2349,RIfe9f828_8159,RIe1529b8_2317,RIfe9f990_8160,RIe14fcb8_2285,RIfcbd368_7175,RIe14cfb8_2253,RIe14a2b8_2221,RIe1475b8_2189,
        RIfc8ee50_6648,RIfc45278_5809,RIfc98360_6754,RIfca2248_6867,RIe141d20_2126,RIe13f9f8_2101,RIdf3d900_2077,RIdf3b470_2051,RIfcd6ca0_7466,RIee2ff08_5004,
        RIfc8ece8_6647,RIee2dd48_4980,RIdf36718_1996,RIdf34120_1969,RIdf31f60_1945,RIfe9f6c0_8158,RIfcb4560_7074,RIfc45db8_5817,RIfc8e1a8_6639,RIfc7d678_6449,
        RIdf2aee0_1865,RIdf28ff0_1843,RIdf26e30_1819,RIdf25378_1800,RIfcb43f8_7073,RIfc8e748_6643,RIdf23488_1778,RIfcc2c00_7238,RIdf21e08_1762,RIdf20788_1746,
        RIdf1b760_1689,RIdf1a248_1674,RIdf18088_1650,RIdf15388_1618,RIdf12688_1586,RIdf0f988_1554,RIdf0cc88_1522,RIdf09f88_1490,RIdf07288_1458,RIdf04588_1426,
        RIdefeb88_1362,RIdefbe88_1330,RIdef9188_1298,RIdef6488_1266,RIdef3788_1234,RIdef0a88_1202,RIdeedd88_1170,RIdeeb088_1138,RIfc8efb8_6649,RIfc44e40_5806,
        RIfc57860_6018,RIfca23b0_6868,RIfe9faf8_8161,RIdee3900_1053,RIdee1740_1029,RIdedf6e8_1006,RIfcbd4d0_7176,RIee22678_4850,RIfc98090_6752,RIee21598_4838,
        RIfe9fc60_8162,RIded80c8_922,RIfe9fdc8_8163,RIded3be0_873,RIded18b8_848,RIdecebb8_816,RIdecbeb8_784,RIdec91b8_752,RIdeb56b8_528,RIde99080_336,
        RIe16f2c0_2642,RIe15b0b8_2413,RIe1448b8_2157,RIdf392b0_2027,RIdf2d910_1895,RIdf1e190_1719,RIdf01888_1394,RIdee8388_1106,RIdedd0f0_979,RIde7efc8_209,
        RIe19e750_3180,RIbc625c8_12,RIbc62550_11,RIbc624d8_10,RIbc62460_9,RIbc623e8_8,RIbc62370_7,RIbc622f8_6,RIbc62280_5,RIbc62208_4,
        RIbc62190_3,RIbc62118_2,RIe19ba50_3148,RIfc479d8_5837,RIe198d50_3116,RIfe9f558_8157,RIe196050_3084,RIe193350_3052,RIe190650_3020,RIe18ac50_2956,
        RIe187f50_2924,RIfc47870_5836,RIe185250_2892,RIf142ef8_5221,RIe182550_2860,RIe17f850_2828,RIe17cb50_2796,RIfcb5208_7083,RIfcbc6c0_7166,RIe177588_2735,
        RIe176610_2724,RIf13fdc0_5186,RIfe9f3f0_8156,RIfce40f8_7617,RIfc47708_5835,RIfc47438_5833,RIfca15a0_6858,RIfc99170_6764,RIe1745b8_2701,RIfc8cc90_6624,
        RIfc556a0_5994,RIfc7ee60_6466,RIfce8e50_7672,RIfe9f288_8155,RIe224aa8_4707,RIfc55808_5995,RIe221da8_4675,RIfcb50a0_7082,RIe21f0a8_4643,RIe2196a8_4579,
        RIe2169a8_4547,RIfcbc828_7167,RIe213ca8_4515,RIfc47000_5830,RIe210fa8_4483,RIfcbc990_7168,RIe20e2a8_4451,RIe20b5a8_4419,RIe2088a8_4387,RIfc46bc8_5827,
        RIfcd6598_7461,RIe2032e0_4326,RIe2016c0_4306,RIfc98ea0_6762,RIfc7eb90_6464,RIfce0318_7573,RIfcbcaf8_7169,RIfc8cf60_6626,RIfcb4dd0_7080,RIe1fd340_4258,
        RIe1fc260_4246,RIf15cf38_5517,RIfe9f120_8154,RIfc7ea28_6463,RIfc8d0c8_6627,RIfcbcc60_7170,RIfc98bd0_6760,RIfce2d48_7603,RIe1fb018_4233,RIfc55f10_6000,
        RIfc7e8c0_6462,RIfc8d230_6628,RIe1f6590_4180,RIfce58e0_7634,RIfc468f8_5825,RIfcc2ed0_7240,RIe1f4100_4154,RIfceedf0_7740,RIfc8d398_6629,RIfc8d500_6630,
        RIe1eef70_4096,RIe1ec810_4068,RIe1e9b10_4036,RIe1e6e10_4004,RIe1e4110_3972,RIe1e1410_3940,RIe1de710_3908,RIe1dba10_3876,RIe1d8d10_3844,RIe1d3310_3780,
        RIe1d0610_3748,RIe1cd910_3716,RIe1cac10_3684,RIe1c7f10_3652,RIe1c5210_3620,RIe1c2510_3588,RIe1bf810_3556,RIf14d0b0_5336,RIfe9efb8_8153,RIe1ba248_3495,
        RIe1b8088_3471,RIfec4dd0_8360,RIfec50a0_8362,RIe1b5ec8_3447,RIe1b46e0_3430,RIfcb4998_7077,RIfcb4c68_7079,RIfec5370_8364,RIfe9ee50_8152,RIfcbcdc8_7171,
        RIfc46358_5821,RIfec5208_8363,RIfec4f38_8361,RIe1a9b50_3308,RIe1a6e50_3276,RIe1a4150_3244,RIe1a1450_3212,RIe18d950_2988,RIe179e50_2764,RIe2277a8_4739,
        RIe21c3a8_4611,RIe205ba8_4355,RIe1ffc08_4287,RIe1f8fc0_4210,RIe1f1b08_4127,RIe1d6010_3812,RIe1bcb10_3524,RIe1af988_3375,RIe171fc0_2674,RIdec6080_717,
        RIdec3380_685,RIee204b8_4826,RIdec0680_653,RIfcd70d8_7469,RIdebd980_621,RIdebac80_589,RIdeb7f80_557,RIfcbe448_7187,RIdeb2580_493,RIfcb3480_7062,
        RIdeaf880_461,RIfc43928_5791,RIdeac1a8_429,RIdea58a8_397,RIde9efa8_365,RIfcd88c0_7486,RIee1c408_4780,RIfcc77f0_7292,RIfea04d0_8168,RIde92438_303,
        RIde8ec70_286,RIde8aad0_266,RIde86930_246,RIfca31c0_6878,RIfc59a20_6042,RIfcd1de0_7410,RIfc91448_6675,RIfc97280_6742,RIe16c188_2607,RIfc97118_6741,
        RIe168948_2567,RIe166080_2538,RIe163380_2506,RIee37ac8_5092,RIe160680_2474,RIfcd1c78_7409,RIe15d980_2442,RIe157f80_2378,RIe155280_2346,RIfc3f530_5746,
        RIe152580_2314,RIee35368_5064,RIe14f880_2282,RIfc7a3d8_6413,RIe14cb80_2250,RIe149e80_2218,RIe147180_2186,RIfc42b18_5781,RIfc7a270_6412,RIfc5a560_6050,
        RIfc96b78_6737,RIfea6fb0_8216,RIe13f5c0_2098,RIdf3d4c8_2074,RIdf3b038_2048,RIfce5bb0_7636,RIee2fc38_5002,RIfc91cb8_6681,RIee2d910_4977,RIdf362e0_1993,
        RIdf33e50_1967,RIdf31c90_1943,RIdf2fda0_1921,RIfc43658_5789,RIfc59e58_6045,RIfc96fb0_6740,RIfc7ac48_6419,RIfea0368_8167,RIdf28bb8_1840,RIdf26cc8_1818,
        RIdf25210_1799,RIfc91718_6677,RIfcb3318_7061,RIfc919e8_6679,RIfc91880_6678,RIfc430b8_5785,RIdf20350_1743,RIfc7a978_6417,RIdf19e10_1671,RIdf17c50_1647,
        RIdf14f50_1615,RIdf12250_1583,RIdf0f550_1551,RIdf0c850_1519,RIdf09b50_1487,RIdf06e50_1455,RIdf04150_1423,RIdefe750_1359,RIdefba50_1327,RIdef8d50_1295,
        RIdef6050_1263,RIdef3350_1231,RIdef0650_1199,RIdeed950_1167,RIdeeac50_1135,RIfcd1b10_7408,RIfc968a8_6735,RIfc91f88_6683,RIfcdfc10_7568,RIfea99e0_8246,
        RIdee3630_1051,RIdee1308_1026,RIdedf2b0_1003,RIfcc7d90_7296,RIfcd85f0_7484,RIfce3888_7611,RIfc5a830_6052,RIdeda3f0_947,RIfea9878_8245,RIded5f08_898,
        RIded37a8_870,RIded1480_845,RIdece780_813,RIdecba80_781,RIdec8d80_749,RIdeb5280_525,RIde986a8_333,RIe16ee88_2639,RIe15ac80_2410,RIe144480_2154,
        RIdf38e78_2024,RIdf2d4d8_1892,RIdf1dd58_1716,RIdf01450_1391,RIdee7f50_1103,RIdedccb8_976,RIde7e5f0_206,RIe19e318_3177,RIe19b618_3145,RIfc8f3f0_6652,
        RIe198918_3113,RIf144b18_5241,RIe195c18_3081,RIe192f18_3049,RIe190218_3017,RIe18a818_2953,RIe187b18_2921,RIf143d08_5231,RIe184e18_2889,RIfcb3cf0_7068,
        RIe182118_2857,RIe17f418_2825,RIe17c718_2793,RIfc448a0_5802,RIf141170_5200,RIfc7c9d0_6440,RIfea0098_8165,RIfc57e00_6022,RIf13f550_5180,RIfcd6e08_7467,
        RIee3d900_5159,RIfc8f6c0_6654,RIfce0048_7571,RIfca27e8_6871,RIe1742e8_2699,RIfc7c700_6438,RIfc8f990_6656,RIfce9828_7679,RIfc583a0_6026,RIf16cdc0_5698,
        RIe224670_4704,RIf16c118_5689,RIe221970_4672,RIfc58508_6027,RIe21ec70_4640,RIe219270_4576,RIe216570_4544,RIfc3ff08_5753,RIe213870_4512,RIf1696e8_5659,
        RIe210b70_4480,RIfc58940_6030,RIe20de70_4448,RIe20b170_4416,RIe208470_4384,RIfc8fc60_6658,RIfc97820_6746,RIe202ea8_4323,RIe201288_4303,RIfcc27c8_7235,
        RIfcdfee0_7570,RIfc44198_5797,RIfc58670_6028,RIf1608e0_5558,RIf15e9f0_5536,RIfe9ff30_8164,RIe1fc0f8_4245,RIfc7be90_6432,RIf15bb88_5503,RIfcd8cf8_7489,
        RIfcd8e60_7490,RIfca2d88_6875,RIfcbdea8_7183,RIfcb3a20_7066,RIe1fabe0_4230,RIfc90098_6661,RIfc90200_6662,RIfcd20b0_7412,RIe1f6158_4177,RIfc904d0_6664,
        RIfca2ef0_6876,RIfc97550_6744,RIe1f3e30_4152,RIfc59048_6035,RIfc907a0_6666,RIfc90638_6665,RIe1eeb38_4093,RIe1ec3d8_4065,RIe1e96d8_4033,RIe1e69d8_4001,
        RIe1e3cd8_3969,RIe1e0fd8_3937,RIe1de2d8_3905,RIe1db5d8_3873,RIe1d88d8_3841,RIe1d2ed8_3777,RIe1d01d8_3745,RIe1cd4d8_3713,RIe1ca7d8_3681,RIe1c7ad8_3649,
        RIe1c4dd8_3617,RIe1c20d8_3585,RIe1bf3d8_3553,RIfcc73b8_7289,RIfce3cc0_7614,RIe1b9e10_3492,RIe1b7c50_3468,RIfcd6f70_7468,RIf149e10_5300,RIe1b5a90_3444,
        RIfea0200_8166,RIfc90bd8_6669,RIfcdfd78_7569,RIe1b2ef8_3413,RIe1b15a8_3395,RIfc973e8_6743,RIfcc7520_7290,RIe1acdf0_3344,RIe1ab608_3327,RIe1a9718_3305,
        RIe1a6a18_3273,RIe1a3d18_3241,RIe1a1018_3209,RIe18d518_2985,RIe179a18_2761,RIe227370_4736,RIe21bf70_4608,RIe205770_4352,RIe1ff7d0_4284,RIe1f8b88_4207,
        RIe1f16d0_4124,RIe1d5bd8_3809,RIe1bc6d8_3521,RIe1af550_3372,RIe171b88_2671,RIdec5108_706,RIdec2408_674,RIfc93608_6699,RIdebf708_642,RIfc934a0_6698,
        RIdebca08_610,RIdeb9d08_578,RIdeb7008_546,RIfcdf7d8_7565,RIdeb1608_482,RIfc78218_6389,RIdeae908_450,RIfcc8498_7301,RIdea9d90_418,RIdea3490_386,
        RIde9cb90_354,RIee1cc78_4786,RIee1bb98_4774,RIee1b328_4768,RIee1aab8_4762,RIde909f8_295,RIde8d578_279,RIfea8ea0_8238,RIde85238_239,RIde813e0_220,
        RIfc938d8_6701,RIfce5e80_7638,RIfcbfd98_7205,RIfce8ce8_7671,RIe16b4e0_2598,RIfea8d38_8237,RIfea9f80_8250,RIe165108_2527,RIe162408_2495,RIfc779a8_6383,
        RIe15f708_2463,RIfe9dc08_8139,RIe15ca08_2431,RIe157008_2367,RIe154308_2335,RIfea7550_8220,RIe151608_2303,RIfcd6160_7458,RIe14e908_2271,RIfcd1408_7403,
        RIe14bc08_2239,RIe148f08_2207,RIe146208_2175,RIfceb718_7701,RIfcb19c8_7043,RIfc93e78_6705,RIfce7938_7657,RIe140da8_2115,RIdf3ecb0_2091,RIdf3c988_2066,
        RIfe9daa0_8138,RIfce8478_7665,RIfcdbf98_7525,RIfc776d8_6381,RIfc93fe0_6706,RIdf354d0_1983,RIdf33040_1957,RIdf30fe8_1934,RIdf2ee28_1910,RIee2ba20_4955,
        RIfc93ba8_6703,RIfc77de0_6386,RIee27ad8_4910,RIfe9d668_8135,RIfea8bd0_8236,RIdf26458_1812,RIfe9d7d0_8136,RIfcb1c98_7045,RIee26cc8_4900,RIdf22ab0_1771,
        RIfcc0068_7207,RIdf21598_1756,RIdf1f6a8_1734,RIdf1aef0_1683,RIfe9d938_8137,RIdf16cd8_1636,RIdf13fd8_1604,RIdf112d8_1572,RIdf0e5d8_1540,RIdf0b8d8_1508,
        RIdf08bd8_1476,RIdf05ed8_1444,RIdf031d8_1412,RIdefd7d8_1348,RIdefaad8_1316,RIdef7dd8_1284,RIdef50d8_1252,RIdef23d8_1220,RIdeef6d8_1188,RIdeec9d8_1156,
        RIdee9cd8_1124,RIfc942b0_6708,RIfcde6f8_7553,RIfcd1138_7401,RIfcde860_7554,RIdee4878_1064,RIdee2af0_1043,RIdee0a98_1020,RIdede8d8_996,RIfc5c9f0_6076,
        RIee22240_4847,RIfcc8768_7303,RIee21160_4835,RIded95e0_937,RIded7150_911,RIded5260_889,RIfea76b8_8221,RIded0508_834,RIdecd808_802,RIdecab08_770,
        RIdec7e08_738,RIdeb4308_514,RIde96290_322,RIe16df10_2628,RIe159d08_2399,RIe143508_2143,RIdf37f00_2013,RIdf2c560_1881,RIdf1cde0_1705,RIdf004d8_1380,
        RIdee6fd8_1092,RIdedbd40_965,RIde7c1d8_195,RIe19d3a0_3166,RIe19a6a0_3134,RIfcb2c10_7056,RIe1979a0_3102,RIfc923c0_6686,RIe194ca0_3070,RIe191fa0_3038,
        RIe18f2a0_3006,RIe1898a0_2942,RIe186ba0_2910,RIfc422a8_5775,RIe183ea0_2878,RIfcbecb8_7193,RIe1811a0_2846,RIe17e4a0_2814,RIe17b7a0_2782,RIf142250_5212,
        RIf140bd0_5196,RIfec43f8_8353,RIe175968_2715,RIfc79b68_6407,RIf13efb0_5176,RIfc92528_6687,RIfcb2aa8_7055,RIfcd8320_7482,RIfcea200_7686,RIfc79898_6405,
        RIe1734d8_2689,RIfcd7948_7475,RIfcd7678_7473,RIf16e170_5712,RIfc927f8_6689,RIfc92960_6690,RIe2236f8_4693,RIfc795c8_6403,RIe2209f8_4661,RIf16ad68_5675,
        RIe21dcf8_4629,RIe2182f8_4565,RIe2155f8_4533,RIfe9d398_8133,RIe2128f8_4501,RIfcdb9f8_7521,RIe20fbf8_4469,RIfc41d08_5771,RIe20cef8_4437,RIe20a1f8_4405,
        RIe2074f8_4373,RIfcd7510_7472,RIf166010_5620,RIfe9d230_8132,RIe2008b0_4296,RIf165098_5609,RIfc41ba0_5770,RIfc41a38_5769,RIfc92c30_6692,RIfc418d0_5768,
        RIfc79190_6400,RIe1fcad0_4252,RIfec4560_8354,RIfc79028_6399,RIfcbf258_7197,RIfcc1df0_7228,RIfcd81b8_7481,RIfc92d98_6693,RIfc5b4d8_6061,RIfcd77e0_7474,
        RIe1fa0a0_4222,RIf156188_5439,RIfe9d500_8134,RIf1546d0_5420,RIe1f5348_4167,RIfec4830_8356,RIfec46c8_8355,RIf1508f0_5376,RIe1f3020_4142,RIfce3180_7606,
        RIfce8fb8_7673,RIfcbf690_7200,RIe1edd28_4083,RIe1eb460_4054,RIe1e8760_4022,RIe1e5a60_3990,RIe1e2d60_3958,RIe1e0060_3926,RIe1dd360_3894,RIe1da660_3862,
        RIe1d7960_3830,RIe1d1f60_3766,RIe1cf260_3734,RIe1cc560_3702,RIe1c9860_3670,RIe1c6b60_3638,RIe1c3e60_3606,RIe1c1160_3574,RIe1be460_3542,RIfe9d0c8_8131,
        RIfe9cc90_8128,RIe1b9168_3483,RIe1b7110_3460,RIf14a3b0_5304,RIfe9cb28_8127,RIfe9cf60_8130,RIfe9c9c0_8126,RIfce2208_7595,RIfce9558_7677,RIfe9c858_8125,
        RIfe9cdf8_8129,RIf147110_5268,RIf146468_5259,RIe1ac2b0_3336,RIe1aaac8_3319,RIe1a87a0_3294,RIe1a5aa0_3262,RIe1a2da0_3230,RIe1a00a0_3198,RIe18c5a0_2974,
        RIe178aa0_2750,RIe2263f8_4725,RIe21aff8_4597,RIe2047f8_4341,RIe1fe858_4273,RIe1f7c10_4196,RIe1f0758_4113,RIe1d4c60_3798,RIe1bb760_3510,RIe1ae5d8_3361,
        RIe170c10_2660,RIdec4190_695,RIdec1490_663,RIfceaa70_7692,RIdebe790_631,RIfc954f8_6721,RIdebba90_599,RIdeb8d90_567,RIdeb6090_535,RIfcebb50_7704,
        RIdeb0690_471,RIee1e190_4801,RIdead990_439,RIfcdf0d0_7560,RIdea7978_407,RIdea1078_375,RIde9a778_343,RIee1c840_4783,RIfc957c8_6723,RIfcc8e70_7308,
        RIfc5e610_6096,RIfe9e8b0_8148,RIde8c1c8_273,RIde88028_253,RIde83b40_232,RIfcb0bb8_7033,RIfca4b10_6896,RIfc75d88_6363,RIfca4c78_6897,RIfc95390_6720,
        RIe16a9a0_2590,RIfcc8fd8_7309,RIe166e90_2548,RIe164190_2516,RIe161490_2484,RIfe9e748_8147,RIe15e790_2452,RIfc74f78_6353,RIe15ba90_2420,RIe156090_2356,
        RIe153390_2324,RIfc3ecc0_5740,RIe150690_2292,RIfce8b80_7670,RIe14d990_2260,RIfca6730_6916,RIe14ac90_2228,RIe147f90_2196,RIe145290_2164,RIfcee2b0_7732,
        RIfc5f2b8_6105,RIfc753b0_6356,RIfc74b40_6350,RIe140268_2107,RIdf3e170_2083,RIdf3be48_2058,RIdf39c88_2034,RIfcc1c88_7227,RIfcc1850_7224,RIfc965d8_6733,
        RIfc96038_6729,RIdf34828_1974,RIdf327d0_1951,RIdf301d8_1924,RIdf2e2e8_1902,RIfc5e778_6097,RIfcd0328_7391,RIfc757e8_6359,RIfcee6e8_7735,RIdf296f8_1848,
        RIdf273d0_1823,RIdf257b0_1803,RIdf23b90_1783,RIfc95d68_6727,RIfceda40_7726,RIfe9eb80_8150,RIfc75518_6357,RIfcd01c0_7390,RIdf1eb68_1726,RIfe9ece8_8151,
        RIfe9ea18_8149,RIdf15d60_1625,RIdf13060_1593,RIdf10360_1561,RIdf0d660_1529,RIdf0a960_1497,RIdf07c60_1465,RIdf04f60_1433,RIdf02260_1401,RIdefc860_1337,
        RIdef9b60_1305,RIdef6e60_1273,RIdef4160_1241,RIdef1460_1209,RIdeee760_1177,RIdeeba60_1145,RIdee8d60_1113,RIfc961a0_6730,RIfc96308_6731,RIfc5ee80_6102,
        RIfce6150_7640,RIdee42d8_1060,RIdee1e48_1034,RIdee00c0_1013,RIdeddac8_986,RIfc96470_6732,RIfc75248_6355,RIfc74ca8_6351,RIfcb0618_7029,RIded8938_928,
        RIded6610_903,RIded4450_879,RIded2290_855,RIdecf590_823,RIdecc890_791,RIdec9b90_759,RIdec6e90_727,RIdeb3390_503,RIde93e78_311,RIe16cf98_2617,
        RIe158d90_2388,RIe142590_2132,RIdf36f88_2002,RIdf2b5e8_1870,RIdf1be68_1694,RIdeff560_1369,RIdee6060_1081,RIdedadc8_954,RIde79dc0_184,RIe19c428_3155,
        RIe199728_3123,RIfe9e310_8144,RIe196a28_3091,RIfcc04a0_7210,RIe193d28_3059,RIe191028_3027,RIe18e328_2995,RIe188928_2931,RIe185c28_2899,RIfce1830_7588,
        RIe182f28_2867,RIfe9e478_8145,RIe180228_2835,RIe17d528_2803,RIe17a828_2771,RIf141878_5205,RIfcb12c0_7038,RIfc94418_6709,RIe174f90_2708,RIfc77408_6379,
        RIf13ea10_5172,RIfcdc100_7526,RIfc94580_6710,RIfc946e8_6711,RIfced338_7721,RIfce5fe8_7639,RIe172998_2681,RIfcdc268_7527,RIfcddff0_7548,RIfcc0608_7211,
        RIfce7230_7652,RIfc40340_5756,RIe222780_4682,RIfcdd618_7541,RIe21fa80_4650,RIfcd0b98_7397,RIe21cd80_4618,RIe217380_4554,RIe214680_4522,RIfec4998_8357,
        RIe211980_4490,RIf168608_5647,RIe20ec80_4458,RIfcc0770_7212,RIe20bf80_4426,RIe209280_4394,RIe206580_4362,RIfce2370_7596,RIfcee580_7734,RIfec4c68_8359,
        RIfec4b00_8358,RIfc949b8_6713,RIfcebcb8_7705,RIf162938_5581,RIf1612b8_5565,RIfccd088_7355,RIfcc08d8_7213,RIfe9e040_8142,RIfe9e1a8_8143,RIfcead40_7694,
        RIf15ad78_5493,RIfc94c88_6715,RIfccc3e0_7346,RIfc765f8_6369,RIfc94df0_6716,RIfcc0a40_7214,RIe1f9998_4217,RIfcc8d08_7307,RIfce8748_7667,RIfceb2e0_7698,
        RIe1f4970_4160,RIf152510_5396,RIf1512c8_5383,RIfcb0ff0_7036,RIe1f24e0_4134,RIfc761c0_6366,RIfc950c0_6718,RIfcc0e78_7217,RIe1ed1e8_4075,RIe1ea4e8_4043,
        RIe1e77e8_4011,RIe1e4ae8_3979,RIe1e1de8_3947,RIe1df0e8_3915,RIe1dc3e8_3883,RIe1d96e8_3851,RIe1d69e8_3819,RIe1d0fe8_3755,RIe1ce2e8_3723,RIe1cb5e8_3691,
        RIe1c88e8_3659,RIe1c5be8_3627,RIe1c2ee8_3595,RIe1c01e8_3563,RIe1bd4e8_3531,RIf14bfd0_5324,RIf14ac20_5310,RIfe9ded8_8141,RIe1b65d0_3452,RIfcecd98_7717,
        RIfc76490_6368,RIe1b4c80_3434,RIe1b38d0_3420,RIfcc0fe0_7218,RIfceaea8_7695,RIe1b1f80_3402,RIe1b0360_3382,RIfcd0760_7394,RIf145ec8_5255,RIfe9e5e0_8146,
        RIfe9dd70_8140,RIe1a7828_3283,RIe1a4b28_3251,RIe1a1e28_3219,RIe19f128_3187,RIe18b628_2963,RIe177b28_2739,RIe225480_4714,RIe21a080_4586,RIe203880_4330,
        RIe1fd8e0_4262,RIe1f6c98_4185,RIe1ef7e0_4102,RIe1d3ce8_3787,RIe1ba7e8_3499,RIe1ad660_3350,RIe16fc98_2649,RIdec6788_722,RIdec3a88_690,RIee20788_4828,
        RIdec0d88_658,RIee1f810_4817,RIdebe088_626,RIdebb388_594,RIdeb8688_562,RIfc9b1c8_6787,RIdeb2c88_498,RIfce1f38_7593,RIdeaff88_466,RIfc892e8_6583,
        RIdead210_434,RIdea6910_402,RIdea0010_370,RIee1d650_4793,RIee1c570_4781,RIee1b5f8_4770,RIee1aef0_4765,RIfe99888_8091,RIfe99450_8088,RIfe99720_8090,
        RIfe995b8_8089,RIde83168_229,RIfcc43e8_7255,RIfcd5a58_7453,RIfc89450_6584,RIfcc5798_7269,RIe16c890_2612,RIe16a568_2587,RIe168d80_2570,RIe166788_2543,
        RIe163a88_2511,RIfc83618_6517,RIe160d88_2479,RIee36718_5078,RIe15e088_2447,RIe158688_2383,RIe155988_2351,RIfc3f800_5748,RIe152c88_2319,RIfc895b8_6585,
        RIe14ff88_2287,RIfc51cf8_5953,RIe14d288_2255,RIe14a588_2223,RIe147888_2191,RIee34990_5057,RIee338b0_5045,RIfc831e0_6514,RIfcd3b68_7431,RIe141ff0_2128,
        RIe13fcc8_2103,RIdf3dbd0_2079,RIdf3b740_2053,RIfcb6f90_7104,RIee301d8_5006,RIfcba938_7145,RIee2e018_4982,RIdf369e8_1998,RIdf343f0_1971,RIdf32230_1947,
        RIfe99e28_8095,RIfc83078_6513,RIfcb6e28_7103,RIfc9ad90_6784,RIfcbad70_7148,RIdf2b1b0_1867,RIdf292c0_1845,RIfe99b58_8093,RIfe999f0_8092,RIfc9ac28_6783,
        RIfc4a9a8_5871,RIdf23758_1780,RIfc82da8_6511,RIdf220d8_1764,RIdf20a58_1748,RIdf1ba30_1691,RIfe99cc0_8094,RIdf18358_1652,RIdf15658_1620,RIdf12958_1588,
        RIdf0fc58_1556,RIdf0cf58_1524,RIdf0a258_1492,RIdf07558_1460,RIdf04858_1428,RIdefee58_1364,RIdefc158_1332,RIdef9458_1300,RIdef6758_1268,RIdef3a58_1236,
        RIdef0d58_1204,RIdeee058_1172,RIdeeb358_1140,RIee25918_4886,RIee24b08_4876,RIfc52568_5959,RIfc826a0_6506,RIdee5958_1076,RIdee3bd0_1055,RIfe99f90_8096,
        RIdedf9b8_1008,RIfce4800_7622,RIfc89b58_6589,RIfc9f3e0_6834,RIfc82538_6505,RIdeda828_950,RIded8398_924,RIfeabe70_8272,RIded3eb0_875,RIded1b88_850,
        RIdecee88_818,RIdecc188_786,RIdec9488_754,RIdeb5988_530,RIde99710_338,RIe16f590_2644,RIe15b388_2415,RIe144b88_2159,RIdf39580_2029,RIdf2dbe0_1897,
        RIdf1e460_1721,RIdf01b58_1396,RIdee8658_1108,RIdedd3c0_981,RIde7f658_211,RIe19ea20_3182,RIe19bd20_3150,RIf145928_5251,RIe199020_3118,RIfe98910_8080,
        RIe196320_3086,RIe193620_3054,RIe190920_3022,RIe18af20_2958,RIe188220_2926,RIf143e70_5232,RIe185520_2894,RIfc95c00_6726,RIe182820_2862,RIe17fb20_2830,
        RIe17ce20_2798,RIf142520_5214,RIf141440_5202,RIe1776f0_2736,RIfeab8d0_8268,RIfcc5bd0_7272,RIfc62dc8_6147,RIee3e710_5169,RIfc9cb18_6805,RIee3c820_5147,
        RIee3b470_5133,RIee3a390_5121,RIe174888_2703,RIf170498_5737,RIfc68660_6210,RIf16e878_5717,RIfc6ea38_6281,RIfe98d48_8083,RIe224d78_4709,RIf16c280_5690,
        RIe222078_4677,RIf16b308_5679,RIe21f378_4645,RIe219978_4581,RIe216c78_4549,RIf16a390_5668,RIe213f78_4517,RIf169b20_5662,RIe211278_4485,RIf1681d0_5644,
        RIe20e578_4453,RIe20b878_4421,RIe208b78_4389,RIfcd4ae0_7442,RIfc61478_6129,RIfeab060_8262,RIe201990_4308,RIfc70ec8_6307,RIfc70928_6303,RIfcec528_7711,
        RIfcbe880_7190,RIf160d18_5561,RIf15ee28_5539,RIfe98be0_8082,RIfe98eb0_8084,RIf15d0a0_5518,RIf15bcf0_5504,RIfcd4540_7438,RIf159e00_5482,RIf1592c0_5474,
        RIf158078_5461,RIfca3a30_6884,RIfea7988_8223,RIf156728_5443,RIf155be8_5435,RIf154b08_5423,RIfe98a78_8081,RIf1538c0_5410,RIf1520d8_5393,RIf150e90_5380,
        RIe1f43d0_4156,RIf14fdb0_5368,RIfcd2380_7414,RIf14e2f8_5349,RIe1ef240_4098,RIe1ecae0_4070,RIe1e9de0_4038,RIe1e70e0_4006,RIe1e43e0_3974,RIe1e16e0_3942,
        RIe1de9e0_3910,RIe1dbce0_3878,RIe1d8fe0_3846,RIe1d35e0_3782,RIe1d08e0_3750,RIe1cdbe0_3718,RIe1caee0_3686,RIe1c81e0_3654,RIe1c54e0_3622,RIe1c27e0_3590,
        RIe1bfae0_3558,RIfc44b70_5804,RIf14bd00_5322,RIfe992e8_8087,RIfe987a8_8079,RIf14a950_5308,RIf149f78_5301,RIfe99180_8086,RIfe98640_8078,RIf149438_5293,
        RIfcec7f8_7713,RIfe984d8_8077,RIe1b1b48_3399,RIfc4b650_5880,RIfcda918_7509,RIfe98370_8076,RIfe99018_8085,RIe1a9e20_3310,RIe1a7120_3278,RIe1a4420_3246,
        RIe1a1720_3214,RIe18dc20_2990,RIe17a120_2766,RIe227a78_4741,RIe21c678_4613,RIe205e78_4357,RIe1ffed8_4289,RIe1f9290_4212,RIe1f1dd8_4129,RIe1d62e0_3814,
        RIe1bcde0_3526,RIe1afc58_3377,RIe172290_2676,RIdec6620_721,RIdec3920_689,RIfc49328_5855,RIdec0c20_657,RIfc80eb8_6489,RIdebdf20_625,RIdebb220_593,
        RIdeb8520_561,RIfc80648_6483,RIdeb2b20_497,RIfc8b340_6606,RIdeafe20_465,RIfc491c0_5854,RIdeacec8_433,RIdea65c8_401,RIde9fcc8_369,RIfcd9c70_7500,
        RIfe98208_8075,RIfce4698_7621,RIfe980a0_8074,RIde93158_307,RIde8f648_289,RIde8b4a8_269,RIde87308_249,RIde82e20_228,RIfcbba18_7157,RIfc48d88_5851,
        RIfc99f80_6774,RIfc8b4a8_6607,RIe16c728_2611,RIe16a400_2586,RIe168c18_2569,RIe166620_2542,RIe163920_2510,RIee38068_5096,RIe160c20_2478,RIfc48248_5843,
        RIe15df20_2446,RIe158520_2382,RIe155820_2350,RIfcbbe50_7160,RIe152b20_2318,RIfc47e10_5840,RIe14fe20_2286,RIfca0e98_6853,RIe14d120_2254,RIe14a420_2222,
        RIe147720_2190,RIfc8be80_6614,RIfc7fb08_6475,RIfc480e0_5842,RIfc99878_6769,RIe141e88_2127,RIe13fb60_2102,RIdf3da68_2078,RIdf3b5d8_2052,RIfe97f38_8073,
        RIee30070_5005,RIee2eb58_4990,RIee2deb0_4981,RIdf36880_1997,RIdf34288_1970,RIdf320c8_1946,RIfe97dd0_8072,RIfcc3740_7246,RIfc48ab8_5849,RIfce05e8_7575,
        RIfc80210_6480,RIdf2b048_1866,RIdf29158_1844,RIdf26f98_1820,RIdf254e0_1801,RIfc8bbb0_6612,RIfc48950_5848,RIdf235f0_1779,RIfc8bd18_6613,RIdf21f70_1763,
        RIdf208f0_1747,RIdf1b8c8_1690,RIdf1a3b0_1675,RIdf181f0_1651,RIdf154f0_1619,RIdf127f0_1587,RIdf0faf0_1555,RIdf0cdf0_1523,RIdf0a0f0_1491,RIdf073f0_1459,
        RIdf046f0_1427,RIdefecf0_1363,RIdefbff0_1331,RIdef92f0_1299,RIdef65f0_1267,RIdef38f0_1235,RIdef0bf0_1203,RIdeedef0_1171,RIdeeb1f0_1139,RIfcbc120_7162,
        RIfcd9838_7497,RIfc99710_6768,RIfca1168_6855,RIdee57f0_1075,RIdee3a68_1054,RIdee18a8_1030,RIdedf850_1007,RIfc549f8_5985,RIfcb5370_7084,RIfce43c8_7619,
        RIfce0480_7574,RIdeda6c0_949,RIded8230_923,RIded6070_899,RIded3d48_874,RIded1a20_849,RIdeced20_817,RIdecc020_785,RIdec9320_753,RIdeb5820_529,
        RIde993c8_337,RIe16f428_2643,RIe15b220_2414,RIe144a20_2158,RIdf39418_2028,RIdf2da78_1896,RIdf1e2f8_1720,RIdf019f0_1395,RIdee84f0_1107,RIdedd258_980,
        RIde7f310_210,RIe19e8b8_3181,RIe19bbb8_3149,RIfe976c8_8067,RIe198eb8_3117,RIf144c80_5242,RIe1961b8_3085,RIe1934b8_3053,RIe1907b8_3021,RIe18adb8_2957,
        RIe1880b8_2925,RIfe97560_8066,RIe1853b8_2893,RIfcc3fb0_7252,RIe1826b8_2861,RIe17f9b8_2829,RIe17ccb8_2797,RIfcd3730_7428,RIf1412d8_5201,RIfcc4118_7253,
        RIfe97830_8068,RIfc4a6d8_5869,RIf13f6b8_5181,RIfc9f980_6838,RIfc9fae8_6839,RIfcc3e48_7251,RIfc89e28_6591,RIfc89cc0_6590,RIe174720_2702,RIfc4a408_5867,
        RIfce27a8_7599,RIfc530a8_5967,RIfcd5d28_7455,RIf16cf28_5699,RIe224c10_4708,RIfc53210_5968,RIe221f10_4676,RIf16b1a0_5678,RIe21f210_4644,RIe219810_4580,
        RIe216b10_4548,RIfc401d8_5755,RIe213e10_4516,RIf1699b8_5661,RIe211110_4484,RIfc81cc8_6499,RIe20e410_4452,RIe20b710_4420,RIe208a10_4388,RIfc8a0f8_6593,
        RIfcb6720_7098,RIe203448_4327,RIe201828_4307,RIfc53378_5969,RIfc8a3c8_6595,RIfcb65b8_7097,RIfc49fd0_5864,RIf160bb0_5560,RIf15ecc0_5538,RIe1fd4a8_4259,
        RIfe97b00_8070,RIfc8a530_6596,RIfe97c68_8071,RIfc8a800_6598,RIfc8a698_6597,RIfc9a7f0_6780,RIfc81890_6496,RIfcd5e90_7456,RIe1fb180_4234,RIfc49e68_5863,
        RIfc81728_6495,RIfcbb1a8_7151,RIe1f66f8_4181,RIfcd3460_7426,RIfcb62e8_7095,RIfc9a520_6778,RIe1f4268_4155,RIfc49d00_5862,RIfcd9dd8_7501,RIfcbb310_7152,
        RIe1ef0d8_4097,RIe1ec978_4069,RIe1e9c78_4037,RIe1e6f78_4005,RIe1e4278_3973,RIe1e1578_3941,RIe1de878_3909,RIe1dbb78_3877,RIe1d8e78_3845,RIe1d3478_3781,
        RIe1d0778_3749,RIe1cda78_3717,RIe1cad78_3685,RIe1c8078_3653,RIe1c5378_3621,RIe1c2678_3589,RIe1bf978_3557,RIfc49a30_5860,RIfcb6018_7093,RIe1ba3b0_3496,
        RIe1b81f0_3472,RIfce0a20_7578,RIfcbb5e0_7154,RIe1b6030_3448,RIfe97998_8069,RIfce5610_7632,RIfcc3a10_7248,RIe1b3330_3416,RIe1b19e0_3398,RIfc495f8_5857,
        RIfc81188_6491,RIe1ad228_3347,RIe1aba40_3330,RIe1a9cb8_3309,RIe1a6fb8_3277,RIe1a42b8_3245,RIe1a15b8_3213,RIe18dab8_2989,RIe179fb8_2765,RIe227910_4740,
        RIe21c510_4612,RIe205d10_4356,RIe1ffd70_4288,RIe1f9128_4211,RIe1f1c70_4128,RIe1d6178_3813,RIe1bcc78_3525,RIe1afaf0_3376,RIe172128_2675,RIdec6a58_724,
        RIdec3d58_692,RIfc723e0_6322,RIdec1058_660,RIfc59fc0_6046,RIdebe358_628,RIdebb658_596,RIdeb8958_564,RIfcb96f0_7132,RIdeb2f58_500,RIfce1c68_7591,
        RIdeb0258_468,RIfc9b498_6789,RIdead558_436,RIdea6fa0_404,RIdea06a0_372,RIfc81458_6493,RIfc83780_6518,RIfc4e620_5914,RIfcd3e38_7433,RIde937e8_309,
        RIde8f990_290,RIde8bb38_271,RIde87650_250,RIde834b0_230,RIfc42c80_5782,RIfc65960_6178,RIfc6c710_6256,RIee392b0_5109,RIe16cb60_2614,RIe16a6d0_2588,
        RIe169050_2572,RIe166a58_2545,RIe163d58_2513,RIfec3cf0_8348,RIe161058_2481,RIfcd54b8_7449,RIe15e358_2449,RIe158958_2385,RIe155c58_2353,RIfe9ba48_8115,
        RIe152f58_2321,RIfec4128_8351,RIe150258_2289,RIfcb9b28_7135,RIe14d558_2257,RIe14a858_2225,RIe147b58_2193,RIfcdb2f0_7516,RIfc553d0_5992,RIfc9a0e8_6775,
        RIfcbd908_7179,RIe1422c0_2130,RIe13ff98_2105,RIdf3dea0_2081,RIdf3ba10_2055,RIfc87128_6559,RIee304a8_5008,RIfcc51f8_7265,RIee2e2e8_4984,RIdf36cb8_2000,
        RIfec3fc0_8350,RIdf32500_1949,RIfec3e58_8349,RIee2c830_4965,RIee2ad78_4946,RIee296f8_4930,RIee284b0_4917,RIfe9b8e0_8114,RIfe9b610_8112,RIfe9b778_8113,
        RIfe9b4a8_8111,RIfcb7c38_7113,RIfc86b88_6555,RIdf238c0_1781,RIfc75ab8_6361,RIdf22240_1765,RIfeaa3b8_8253,RIdf1bb98_1692,RIdf1a680_1677,RIdf18628_1654,
        RIdf15928_1622,RIdf12c28_1590,RIdf0ff28_1558,RIdf0d228_1526,RIdf0a528_1494,RIdf07828_1462,RIdf04b28_1430,RIdeff128_1366,RIdefc428_1334,RIdef9728_1302,
        RIdef6a28_1270,RIdef3d28_1238,RIdef1028_1206,RIdeee328_1174,RIdeeb628_1142,RIee25a80_4887,RIee24c70_4877,RIfcddd20_7546,RIfccc110_7344,RIdee5c28_1078,
        RIdee3ea0_1057,RIdee1b78_1032,RIdedfc88_1010,RIfc6a6b8_6233,RIee227e0_4851,RIfc88be0_6578,RIee21868_4840,RIdedaaf8_952,RIded8668_926,RIded6340_901,
        RIded4180_877,RIded1e58_852,RIdecf158_820,RIdecc458_788,RIdec9758_756,RIdeb5c58_532,RIde99da0_340,RIe16f860_2646,RIe15b658_2417,RIe144e58_2161,
        RIdf39850_2031,RIdf2deb0_1899,RIdf1e730_1723,RIdf01e28_1398,RIdee8928_1110,RIdedd690_983,RIde7fce8_213,RIe19ecf0_3184,RIe19bff0_3152,RIf145a90_5252,
        RIe1992f0_3120,RIf144de8_5243,RIe1965f0_3088,RIe1938f0_3056,RIe190bf0_3024,RIe18b1f0_2960,RIe1884f0_2928,RIfc72980_6326,RIe1857f0_2896,RIf143060_5222,
        RIe182af0_2864,RIe17fdf0_2832,RIe17d0f0_2800,RIf142688_5215,RIf141710_5204,RIe177858_2737,RIe176778_2725,RIfcea638_7689,RIfca54e8_6903,RIee3e878_5170,
        RIee3dbd0_5161,RIee3c988_5148,RIee3b5d8_5134,RIee3a4f8_5122,RIe174b58_2705,RIf170600_5738,RIfc76fd0_6376,RIf16e9e0_5718,RIfced608_7723,RIf16d090_5700,
        RIe225048_4711,RIf16c550_5692,RIe222348_4679,RIf16b470_5680,RIe21f648_4647,RIe219c48_4583,RIe216f48_4551,RIf16a4f8_5669,RIe214248_4519,RIf169df0_5664,
        RIe211548_4487,RIf1684a0_5646,RIe20e848_4455,RIe20bb48_4423,RIe208e48_4391,RIf1673c0_5634,RIf166448_5623,RIfe9c6f0_8124,RIfe9c150_8120,RIf1654d0_5612,
        RIfcc4550_7256,RIf1635e0_5590,RIf162500_5578,RIf160fe8_5563,RIf15f0f8_5541,RIfe9bfe8_8119,RIfe9c588_8123,RIf15d208_5519,RIf15bfc0_5506,RIfc4d540_5902,
        RIfc9c848_6803,RIfec4290_8352,RIfe9c2b8_8121,RIfcc01d0_7208,RIe1fb2e8_4235,RIfe9c420_8122,RIfca3e68_6887,RIf154c70_5424,RIe1f69c8_4183,RIf153a28_5411,
        RIf152240_5394,RIf150ff8_5381,RIe1f46a0_4158,RIfca6028_6911,RIfc43bf8_5793,RIf14e460_5350,RIe1ef3a8_4099,RIe1ecdb0_4072,RIe1ea0b0_4040,RIe1e73b0_4008,
        RIe1e46b0_3976,RIe1e19b0_3944,RIe1decb0_3912,RIe1dbfb0_3880,RIe1d92b0_3848,RIe1d38b0_3784,RIe1d0bb0_3752,RIe1cdeb0_3720,RIe1cb1b0_3688,RIe1c84b0_3656,
        RIe1c57b0_3624,RIe1c2ab0_3592,RIe1bfdb0_3560,RIfc4d6a8_5903,RIf14be68_5323,RIe1ba680_3498,RIfe9be80_8118,RIfc86e58_6557,RIfcd46a8_7439,RIe1b6300_3450,
        RIfe9bd18_8117,RIf1495a0_5294,RIf1481f0_5280,RIe1b3600_3418,RIe1b1e18_3401,RIfc69470_6220,RIfcbfac8_7203,RIfe9bbb0_8116,RIe1abd10_3332,RIe1aa0f0_3312,
        RIe1a73f0_3280,RIe1a46f0_3248,RIe1a19f0_3216,RIe18def0_2992,RIe17a3f0_2768,RIe227d48_4743,RIe21c948_4615,RIe206148_4359,RIe2001a8_4291,RIe1f9560_4214,
        RIe1f20a8_4131,RIe1d65b0_3816,RIe1bd0b0_3528,RIe1aff28_3379,RIe172560_2678,RIdec68f0_723,RIdec3bf0_691,RIee208f0_4829,RIdec0ef0_659,RIfc7ce08_6443,
        RIdebe1f0_627,RIdebb4f0_595,RIdeb87f0_563,RIfc9b8d0_6792,RIdeb2df0_499,RIfcc6710_7280,RIdeb00f0_467,RIfc5ff60_6114,RIdead3f0_435,RIdea6c58_403,
        RIdea0358_371,RIfce5070_7628,RIee1c6d8_4782,RIfce70c8_7651,RIee1b058_4766,RIde934a0_308,RIfe9b1d8_8109,RIde8b7f0_270,RIfe9b340_8110,RIfc6b798_6245,
        RIfcb2238_7049,RIfcd3a00_7430,RIfcdb020_7514,RIfc511b8_5945,RIe16c9f8_2613,RIfcb27d8_7053,RIe168ee8_2571,RIe1668f0_2544,RIe163bf0_2512,RIee381d0_5097,
        RIe160ef0_2480,RIfcdfaa8_7567,RIe15e1f0_2448,RIe1587f0_2384,RIe155af0_2352,RIfc3f968_5749,RIe152df0_2320,RIfcd5080_7446,RIe1500f0_2288,RIfc84b30_6532,
        RIe14d3f0_2256,RIe14a6f0_2224,RIe1479f0_2192,RIfcea098_7685,RIfc92f00_6694,RIfc54890_5984,RIfcdcc40_7534,RIe142158_2129,RIe13fe30_2104,RIdf3dd38_2080,
        RIdf3b8a8_2054,RIfc57590_6016,RIee30340_5007,RIfcd0490_7392,RIee2e180_4983,RIdf36b50_1999,RIdf34558_1972,RIdf32398_1948,RIfe9b070_8108,RIfcb1860_7042,
        RIfca1b40_6862,RIfc5c018_6069,RIfe9ada0_8106,RIdf2b318_1868,RIdf29428_1846,RIdf27100_1821,RIfe9af08_8107,RIfc5e1d8_6093,RIfcdcda8_7535,RIfcac400_6982,
        RIfc691a0_6218,RIfcaad80_6966,RIdf20bc0_1749,RIfc61b80_6134,RIdf1a518_1676,RIdf184c0_1653,RIdf157c0_1621,RIdf12ac0_1589,RIdf0fdc0_1557,RIdf0d0c0_1525,
        RIdf0a3c0_1493,RIdf076c0_1461,RIdf049c0_1429,RIdefefc0_1365,RIdefc2c0_1333,RIdef95c0_1301,RIdef68c0_1269,RIdef3bc0_1237,RIdef0ec0_1205,RIdeee1c0_1173,
        RIdeeb4c0_1141,RIfc69b78_6225,RIfc6b900_6246,RIfc4d270_5900,RIfced770_7724,RIdee5ac0_1077,RIdee3d38_1056,RIdee1a10_1031,RIdedfb20_1009,RIfc7ff40_6478,
        RIfca4408_6891,RIfcb5640_7086,RIee21700_4839,RIdeda990_951,RIded8500_925,RIded61d8_900,RIded4018_876,RIded1cf0_851,RIdeceff0_819,RIdecc2f0_787,
        RIdec95f0_755,RIdeb5af0_531,RIde99a58_339,RIe16f6f8_2645,RIe15b4f0_2416,RIe144cf0_2160,RIdf396e8_2030,RIdf2dd48_1898,RIdf1e5c8_1722,RIdf01cc0_1397,
        RIdee87c0_1109,RIdedd528_982,RIde7f9a0_212,RIe19eb88_3183,RIe19be88_3151,RIfe9a698_8101,RIe199188_3119,RIfe9a530_8100,RIe196488_3087,RIe193788_3055,
        RIe190a88_3023,RIe18b088_2959,RIe188388_2927,RIfe9a800_8102,RIe185688_2895,RIfc8d938_6633,RIe182988_2863,RIe17fc88_2831,RIe17cf88_2799,RIfe9a3c8_8099,
        RIf1415a8_5203,RIfe9a260_8098,RIfe9a0f8_8097,RIfcb9150_7128,RIf13f820_5182,RIfc9fc50_6840,RIfce5340_7630,RIfc5cb58_6077,RIfc576f8_6017,RIfc780b0_6388,
        RIe1749f0_2704,RIfc7adb0_6420,RIfc7c2c8_6435,RIfcb2d78_7057,RIfc7e758_6461,RIfe9aad0_8104,RIe224ee0_4710,RIf16c3e8_5691,RIe2221e0_4678,RIfcd3898_7429,
        RIe21f4e0_4646,RIe219ae0_4582,RIe216de0_4550,RIfc880a0_6570,RIe2140e0_4518,RIf169c88_5663,RIe2113e0_4486,RIf168338_5645,RIe20e6e0_4454,RIe20b9e0_4422,
        RIe208ce0_4390,RIfce4c38_7625,RIfc9c6e0_6802,RIe2035b0_4328,RIe201af8_4309,RIfc500d8_5933,RIfc85c10_6544,RIfce81a8_7663,RIfce9c60_7682,RIf160e80_5562,
        RIf15ef90_5540,RIfe9a968_8103,RIfe9ac38_8105,RIfca8d28_6943,RIf15be58_5505,RIfcedba8_7727,RIfc6a988_6235,RIfc71cd8_6317,RIfccb198_7333,RIfcaa3a8_6959,
        RIfec3b88_8347,RIfc4c730_5892,RIfc6d688_6267,RIfca8e90_6944,RIe1f6860_4182,RIfc64e20_6170,RIfcaee30_7012,RIfccee10_7376,RIe1f4538_4157,RIfc63ea8_6159,
        RIfcaecc8_7011,RIfcae458_7005,RIfeab1c8_8263,RIe1ecc48_4071,RIe1e9f48_4039,RIe1e7248_4007,RIe1e4548_3975,RIe1e1848_3943,RIe1deb48_3911,RIe1dbe48_3879,
        RIe1d9148_3847,RIe1d3748_3783,RIe1d0a48_3751,RIe1cdd48_3719,RIe1cb048_3687,RIe1c8348_3655,RIe1c5648_3623,RIe1c2948_3591,RIe1bfc48_3559,RIfcc70e8_7287,
        RIfca7ae0_6930,RIe1ba518_3497,RIe1b8358_3473,RIfc598b8_6041,RIfcc2228_7231,RIe1b6198_3449,RIe1b4848_3431,RIfc82f10_6512,RIfc55970_5996,RIe1b3498_3417,
        RIe1b1cb0_3400,RIfcb7698_7109,RIfc4b4e8_5879,RIe1ad390_3348,RIe1abba8_3331,RIe1a9f88_3311,RIe1a7288_3279,RIe1a4588_3247,RIe1a1888_3215,RIe18dd88_2991,
        RIe17a288_2767,RIe227be0_4742,RIe21c7e0_4614,RIe205fe0_4358,RIe200040_4290,RIe1f93f8_4213,RIe1f1f40_4130,RIe1d6448_3815,RIe1bcf48_3527,RIe1afdc0_3378,
        RIe1723f8_2677,RIdec6d28_726,RIdec4028_694,RIee20bc0_4831,RIdec1328_662,RIfcbaed8_7149,RIdebe628_630,RIdebb928_598,RIdeb8c28_566,RIfc412b8_5767,
        RIdeb3228_502,RIfc9ea08_6827,RIdeb0528_470,RIee1e028_4800,RIdead828_438,RIdea7630_406,RIdea0d30_374,RIfcbac08_7147,RIfc55538_5993,RIfcba668_7143,
        RIfc4af48_5875,RIfe912f0_7996,RIfe91458_7997,RIde8be80_272,RIde87ce0_252,RIfc85238_6537,RIfc88640_6574,RIfcda210_7504,RIfcd5788_7451,RIee39418_5110,
        RIe16ce30_2616,RIfc884d8_6573,RIe169320_2574,RIe166d28_2547,RIe164028_2515,RIfe90918_7989,RIe161328_2483,RIee36880_5079,RIe15e628_2451,RIe158c28_2387,
        RIe155f28_2355,RIfe91188_7995,RIe153228_2323,RIfe91020_7994,RIe150528_2291,RIfcda378_7505,RIe14d828_2259,RIe14ab28_2227,RIe147e28_2195,RIfe90eb8_7993,
        RIfe90d50_7992,RIfcb99c0_7134,RIfc9c2a8_6799,RIfe90be8_7991,RIfe90a80_7990,RIdf3e008_2082,RIdf3bce0_2057,RIfcec690_7712,RIee30778_5010,RIfc87dd0_6568,
        RIee2e5b8_4986,RIdf36e20_2001,RIdf346c0_1973,RIdf32668_1950,RIdf30070_1923,RIee2c998_4966,RIee2aee0_4947,RIee299c8_4932,RIee28618_4918,RIfe90378_7985,
        RIfe907b0_7988,RIfe904e0_7986,RIfe90648_7987,RIfc9d928_6815,RIfc86048_6547,RIfcb92b8_7129,RIfc4ee90_5920,RIfc86a20_6554,RIdf20e90_1751,RIfcb8fe8_7127,
        RIdf1a950_1679,RIdf188f8_1656,RIdf15bf8_1624,RIdf12ef8_1592,RIdf101f8_1560,RIdf0d4f8_1528,RIdf0a7f8_1496,RIdf07af8_1464,RIdf04df8_1432,RIdeff3f8_1368,
        RIdefc6f8_1336,RIdef99f8_1304,RIdef6cf8_1272,RIdef3ff8_1240,RIdef12f8_1208,RIdeee5f8_1176,RIdeeb8f8_1144,RIfc857d8_6541,RIee24dd8_4878,RIfc4ff70_5932,
        RIfc50240_5934,RIdee5ef8_1080,RIdee4170_1059,RIfe915c0_7998,RIdedff58_1012,RIfcd4810_7440,RIee22948_4852,RIfce1560_7586,RIee219d0_4841,RIdedac60_953,
        RIfe91728_7999,RIded64a8_902,RIfe91890_8000,RIded2128_854,RIdecf428_822,RIdecc728_790,RIdec9a28_758,RIdeb5f28_534,RIde9a430_342,RIe16fb30_2648,
        RIe15b928_2419,RIe145128_2163,RIdf39b20_2033,RIdf2e180_1901,RIdf1ea00_1725,RIdf020f8_1400,RIdee8bf8_1112,RIdedd960_985,RIde80378_215,RIe19efc0_3186,
        RIe19c2c0_3154,RIf145d60_5254,RIe1995c0_3122,RIfc637a0_6154,RIe1968c0_3090,RIe193bc0_3058,RIe190ec0_3026,RIe18b4c0_2962,RIe1887c0_2930,RIfc62af8_6145,
        RIe185ac0_2898,RIfe8fc70_7980,RIe182dc0_2866,RIe1800c0_2834,RIe17d3c0_2802,RIfe90210_7984,RIfe8ff40_7982,RIfc72f20_6330,RIe176a48_2727,RIfcaf6a0_7018,
        RIfc61040_6126,RIf13e8a8_5171,RIfe900a8_7983,RIee3caf0_5149,RIee3b740_5135,RIee3a660_5123,RIe174e28_2707,RIf170768_5739,RIfc5fdf8_6113,RIf16eb48_5719,
        RIfcaaab0_6964,RIf16d1f8_5701,RIe225318_4713,RIf16c6b8_5693,RIe222618_4681,RIf16b5d8_5681,RIe21f918_4649,RIe219f18_4585,RIe217218_4553,RIfca62f8_6913,
        RIe214518_4521,RIfcc9578_7313,RIe211818_4489,RIfca5a88_6907,RIe20eb18_4457,RIe20be18_4425,RIe209118_4393,RIf167690_5636,RIf166718_5625,RIfe8f9a0_7978,
        RIfe8f838_7977,RIf165638_5613,RIf164990_5604,RIf1638b0_5592,RIf1627d0_5580,RIf161150_5564,RIf15f260_5542,RIe1fd778_4261,RIe1fc530_4248,RIf15d4d8_5521,
        RIf15c290_5508,RIfca20e0_6866,RIf159f68_5483,RIf159428_5475,RIf1581e0_5462,RIfc5ebb0_6100,RIfe8fdd8_7981,RIfc69e48_6227,RIfc5e8e0_6098,RIf154f40_5426,
        RIe1f6b30_4184,RIf153b90_5412,RIf1523a8_5395,RIfce88b0_7668,RIfe8fb08_7979,RIfcebe20_7706,RIfcb1158_7037,RIf14e730_5352,RIe1ef678_4101,RIe1ed080_4074,
        RIe1ea380_4042,RIe1e7680_4010,RIe1e4980_3978,RIe1e1c80_3946,RIe1def80_3914,RIe1dc280_3882,RIe1d9580_3850,RIe1d3b80_3786,RIe1d0e80_3754,RIe1ce180_3722,
        RIe1cb480_3690,RIe1c8780_3658,RIe1c5a80_3626,RIe1c2d80_3594,RIe1c0080_3562,RIfcc8ba0_7306,RIfc5d698_6085,RIfec35e8_8343,RIfeabd08_8271,RIfc5cf90_6080,
        RIfc5ce28_6079,RIfec31b0_8340,RIe1b4b18_3433,RIf149708_5295,RIf148358_5281,RIe1b3768_3419,RIfec3480_8342,RIfc483b0_5844,RIfc80be8_6487,RIe1ad4f8_3349,
        RIfec3318_8341,RIe1aa3c0_3314,RIe1a76c0_3282,RIe1a49c0_3250,RIe1a1cc0_3218,RIe18e1c0_2994,RIe17a6c0_2770,RIe228018_4745,RIe21cc18_4617,RIe206418_4361,
        RIe200478_4293,RIe1f9830_4216,RIe1f2378_4133,RIe1d6880_3818,RIe1bd380_3530,RIe1b01f8_3381,RIe172830_2680,RIdec6bc0_725,RIdec3ec0_693,RIee20a58_4830,
        RIdec11c0_661,RIee1f978_4818,RIdebe4c0_629,RIdebb7c0_597,RIdeb8ac0_565,RIee1efa0_4811,RIdeb30c0_501,RIfcb04b0_7028,RIdeb03c0_469,RIfc5e4a8_6095,
        RIdead6c0_437,RIdea72e8_405,RIdea09e8_373,RIfcb2508_7051,RIfcd16d8_7405,RIfc5d800_6086,RIfc63d40_6158,RIde93b30_310,RIfea7820_8222,RIfea73e8_8219,
        RIde87998_251,RIde837f8_231,RIfc7bd28_6431,RIfcc7ef8_7297,RIfc7a108_6411,RIfc7a6a8_6415,RIe16ccc8_2615,RIe16a838_2589,RIe1691b8_2573,RIe166bc0_2546,
        RIe163ec0_2514,RIee38338_5098,RIe1611c0_2482,RIfc54b60_5986,RIe15e4c0_2450,RIe158ac0_2386,RIe155dc0_2354,RIee35a70_5069,RIe1530c0_2322,RIee357a0_5067,
        RIe1503c0_2290,RIfc9fdb8_6841,RIe14d6c0_2258,RIe14a9c0_2226,RIe147cc0_2194,RIee34af8_5058,RIee33a18_5046,RIee327d0_5033,RIfcbcf30_7172,RIe142428_2131,
        RIe140100_2106,RIfea7280_8218,RIdf3bb78_2056,RIfc731f0_6332,RIee30610_5009,RIfcbe010_7184,RIee2e450_4985,RIfec2ee0_8338,RIfec3048_8339,RIfec2c10_8336,
        RIfec2d78_8337,RIfcb46c8_7075,RIfcb4830_7076,RIee29860_4931,RIfcb88e0_7122,RIdf2b480_1869,RIdf29590_1847,RIdf27268_1822,RIdf25648_1802,RIfcc9de8_7319,
        RIfc53648_5971,RIdf23a28_1782,RIfc823d0_6504,RIdf223a8_1766,RIdf20d28_1750,RIdf1bd00_1693,RIdf1a7e8_1678,RIdf18790_1655,RIdf15a90_1623,RIdf12d90_1591,
        RIdf10090_1559,RIdf0d390_1527,RIdf0a690_1495,RIdf07990_1463,RIdf04c90_1431,RIdeff290_1367,RIdefc590_1335,RIdef9890_1303,RIdef6b90_1271,RIdef3e90_1239,
        RIdef1190_1207,RIdeee490_1175,RIdeeb790_1143,RIee25be8_4888,RIfc6af28_6239,RIee23fc8_4868,RIfccf680_7382,RIdee5d90_1079,RIdee4008_1058,RIdee1ce0_1033,
        RIdedfdf0_1011,RIfc6b090_6240,RIfc534e0_5970,RIfca5920_6906,RIfc66770_6188,RIfe8f6d0_7976,RIded87d0_927,RIfe8f568_7975,RIded42e8_878,RIded1fc0_853,
        RIdecf2c0_821,RIdecc5c0_789,RIdec98c0_757,RIdeb5dc0_533,RIde9a0e8_341,RIe16f9c8_2647,RIe15b7c0_2418,RIe144fc0_2162,RIdf399b8_2032,RIdf2e018_1900,
        RIdf1e898_1724,RIdf01f90_1399,RIdee8a90_1111,RIdedd7f8_984,RIde80030_214,RIe19ee58_3185,RIe19c158_3153,RIf145bf8_5253,RIe199458_3121,RIfe8f298_7973,
        RIe196758_3089,RIe193a58_3057,RIe190d58_3025,RIe18b358_2961,RIe188658_2929,RIfe8f130_7972,RIe185958_2897,RIfc9f278_6833,RIe182c58_2865,RIe17ff58_2833,
        RIe17d258_2801,RIf1427f0_5216,RIfe8efc8_7971,RIe1779c0_2738,RIe1768e0_2726,RIfc81e30_6500,RIfc9ff20_6842,RIfca0088_6843,RIfc81b60_6498,RIfce5778_7633,
        RIfce08b8_7577,RIfc815c0_6494,RIe174cc0_2706,RIfca04c0_6846,RIfc53eb8_5977,RIfcc65a8_7279,RIfc80d50_6488,RIfc804e0_6482,RIe2251b0_4712,RIfc80378_6481,
        RIe2224b0_4680,RIfcb5910_7088,RIe21f7b0_4648,RIe219db0_4584,RIe2170b0_4552,RIfca01f0_6844,RIe2143b0_4520,RIfc82c40_6510,RIe2116b0_4488,RIfc7f6d0_6472,
        RIe20e9b0_4456,RIe20bcb0_4424,RIe208fb0_4392,RIf167528_5635,RIf1665b0_5624,RIe203718_4329,RIe201c60_4310,RIfc9da90_6816,RIfcc5360_7266,RIf163748_5591,
        RIf162668_5579,RIfc7e320_6458,RIfc87998_6565,RIe1fd610_4260,RIe1fc3c8_4247,RIf15d370_5520,RIf15c128_5507,RIfcc5d38_7273,RIfce7d70_7660,RIfc4bd58_5885,
        RIfc55c40_5998,RIfca2ab8_6873,RIe1fb450_4236,RIf156890_5444,RIfcd5ff8_7457,RIf154dd8_5425,RIfec2aa8_8335,RIfcb4b00_7078,RIfcd9400_7494,RIf151160_5382,
        RIe1f4808_4159,RIfc44738_5801,RIfc90908_6667,RIf14e5c8_5351,RIe1ef510_4100,RIe1ecf18_4073,RIe1ea218_4041,RIe1e7518_4009,RIe1e4818_3977,RIe1e1b18_3945,
        RIe1dee18_3913,RIe1dc118_3881,RIe1d9418_3849,RIe1d3a18_3785,RIe1d0d18_3753,RIe1ce018_3721,RIe1cb318_3689,RIe1c8618_3657,RIe1c5918_3625,RIe1c2c18_3593,
        RIe1bff18_3561,RIf14d218_5337,RIfe8ee60_7970,RIfea8090_8228,RIe1b84c0_3474,RIf14aab8_5309,RIfc6c170_6252,RIe1b6468_3451,RIe1b49b0_3432,RIfcafad8_7021,
        RIfcaa948_6963,RIfe8ecf8_7969,RIfe8f400_7974,RIfc67f58_6205,RIfca8ff8_6945,RIfe8eb90_7968,RIe1abe78_3333,RIe1aa258_3313,RIe1a7558_3281,RIe1a4858_3249,
        RIe1a1b58_3217,RIe18e058_2993,RIe17a558_2769,RIe227eb0_4744,RIe21cab0_4616,RIe2062b0_4360,RIe200310_4292,RIe1f96c8_4215,RIe1f2210_4132,RIe1d6718_3817,
        RIe1bd218_3529,RIe1b0090_3380,RIe1726c8_2679,RIdec4460_697,RIdec1760_665,RIee1fae0_4819,RIdebea60_633,RIee1f108_4812,RIdebbd60_601,RIdeb9060_569,
        RIdeb6360_537,RIee1eb68_4808,RIdeb0960_473,RIee1e460_4803,RIdeadc60_441,RIee1d7b8_4794,RIdea8008_409,RIdea1708_377,RIde9ae08_345,RIfe957d8_8045,
        RIfe95508_8043,RIfe95670_8044,RIee1a7e8_4760,RIfe95aa8_8047,RIfe95238_8041,RIfe95940_8046,RIfe953a0_8042,RIee1a0e0_4755,RIee19ca8_4752,RIee19870_4749,
        RIee19438_4746,RIee38ba8_5104,RIfe95c10_8048,RIee384a0_5099,RIfea9440_8242,RIe164460_2518,RIe161760_2486,RIfe942c0_8030,RIe15ea60_2454,RIfe94158_8029,
        RIe15bd60_2422,RIe156360_2358,RIe153660_2326,RIfe94428_8031,RIe150960_2294,RIfe94590_8032,RIe14dc60_2262,RIfc5c2e8_6071,RIe14af60_2230,RIe148260_2198,
        RIe145560_2166,RIee33ce8_5048,RIee32aa0_5035,RIee31858_5022,RIfc5d530_6084,RIe140538_2109,RIdf3e2d8_2084,RIdf3c118_2060,RIdf39df0_2035,RIfcdd780_7542,
        RIee2ee28_4992,RIfcc88d0_7304,RIee2cc68_4968,RIdf34990_1975,RIdf32aa0_1953,RIdf304a8_1926,RIdf2e5b8_1904,RIee2b1b0_4949,RIfe946f8_8033,RIfcb2940_7054,
        RIee273d0_4905,RIfe949c8_8035,RIdf27538_1824,RIfe94b30_8036,RIfe94860_8034,RIee26f98_4902,RIee269f8_4898,RIee26728_4896,RIee26458_4894,RIee26188_4892,
        RIfe94c98_8037,RIee25d50_4889,RIfea9170_8240,RIdf16030_1627,RIdf13330_1595,RIdf10630_1563,RIdf0d930_1531,RIdf0ac30_1499,RIdf07f30_1467,RIdf05230_1435,
        RIdf02530_1403,RIdefcb30_1339,RIdef9e30_1307,RIdef7130_1275,RIdef4430_1243,RIdef1730_1211,RIdeeea30_1179,RIdeebd30_1147,RIdee9030_1115,RIee250a8_4880,
        RIee24298_4870,RIee23758_4862,RIee22d80_4855,RIfe950d0_8040,RIfe94f68_8039,RIfe94e00_8038,RIdeddd98_988,RIee22ab0_4853,RIee21e08_4844,RIfca46d8_6893,
        RIfc5dad0_6088,RIfeaa250_8252,RIfe96048_8051,RIfe95d78_8049,RIfe95ee0_8050,RIdecf860_825,RIdeccb60_793,RIdec9e60_761,RIdec7160_729,RIdeb3660_505,
        RIde94508_313,RIe16d268_2619,RIe159060_2390,RIe142860_2134,RIdf37258_2004,RIdf2b8b8_1872,RIdf1c138_1696,RIdeff830_1371,RIdee6330_1083,RIdedb098_956,
        RIde7a450_186,RIe19c6f8_3157,RIe1999f8_3125,RIf1450b8_5245,RIe196cf8_3093,RIf143fd8_5233,RIe193ff8_3061,RIe1912f8_3029,RIe18e5f8_2997,RIe188bf8_2933,
        RIe185ef8_2901,RIfe973f8_8065,RIe1831f8_2869,RIf142958_5217,RIe1804f8_2837,RIe17d7f8_2805,RIe17aaf8_2773,RIf141b48_5207,RIfc542f0_5980,RIfc800a8_6479,
        RIe175260_2710,RIfca0bc8_6851,RIfc48680_5846,RIee3dea0_5163,RIfcc6878_7281,RIee3ba10_5137,RIee3a930_5125,RIfe97290_8064,RIe172b00_2682,RIf16f958_5729,
        RIf16ee18_5721,RIf16da68_5707,RIf16d360_5702,RIfe96e58_8061,RIe222a50_4684,RIfe96cf0_8060,RIe21fd50_4652,RIf16a660_5670,RIe21d050_4620,RIe217650_4556,
        RIe214950_4524,RIf169f58_5665,RIe211c50_4492,RIf168770_5648,RIe20ef50_4460,RIf1677f8_5637,RIe20c250_4428,RIe209550_4396,RIe206850_4364,RIf166880_5626,
        RIf1657a0_5614,RIe201dc8_4311,RIe2005e0_4294,RIfe96b88_8059,RIf163b80_5594,RIf162c08_5583,RIf161420_5566,RIf15f530_5544,RIf15d7a8_5523,RIfe968b8_8057,
        RIfe96a20_8058,RIfcb3fc0_7070,RIfc7cf70_6444,RIfc579c8_6019,RIf159590_5476,RIf1584b0_5464,RIf157268_5451,RIf1569f8_5445,RIfe965e8_8055,RIf155d50_5436,
        RIf155210_5428,RIf153e60_5414,RIfe96750_8056,RIf1527e0_5398,RIf151430_5384,RIfcd2650_7416,RIe1f2648_4135,RIf14f108_5359,RIfc7f298_6469,RIf14d4e8_5339,
        RIe1ed350_4076,RIe1ea7b8_4045,RIe1e7ab8_4013,RIe1e4db8_3981,RIe1e20b8_3949,RIe1df3b8_3917,RIe1dc6b8_3885,RIe1d99b8_3853,RIe1d6cb8_3821,RIe1d12b8_3757,
        RIe1ce5b8_3725,RIe1cb8b8_3693,RIe1c8bb8_3661,RIe1c5eb8_3629,RIe1c31b8_3597,RIe1c04b8_3565,RIe1bd7b8_3533,RIf14c138_5325,RIf14ad88_5311,RIe1b8790_3476,
        RIfe96480_8054,RIf14a0e0_5302,RIf149870_5296,RIfe97128_8063,RIfe96318_8053,RIf148628_5283,RIfc58d78_6033,RIe1b20e8_3403,RIe1b04c8_3383,RIf146cd8_5265,
        RIfc591b0_6036,RIfe961b0_8052,RIfe96fc0_8062,RIe1a7af8_3285,RIe1a4df8_3253,RIe1a20f8_3221,RIe19f3f8_3189,RIe18b8f8_2965,RIe177df8_2741,RIe225750_4716,
        RIe21a350_4588,RIe203b50_4332,RIe1fdbb0_4264,RIe1f6f68_4187,RIe1efab0_4104,RIe1d3fb8_3789,RIe1baab8_3501,RIe1ad930_3352,RIe16ff68_2651,RIdec42f8_696,
        RIdec15f8_664,RIfcc6cb0_7284,RIdebe8f8_632,RIfe93780_8022,RIdebbbf8_600,RIdeb8ef8_568,RIdeb61f8_536,RIee1ea00_4807,RIdeb07f8_472,RIee1e2f8_4802,
        RIdeadaf8_440,RIfc5d3c8_6083,RIdea7cc0_408,RIdea13c0_376,RIde9aac0_344,RIfc58238_6025,RIfcc3b78_7249,RIfc7d0d8_6445,RIfc59750_6040,RIfe93a50_8024,
        RIfe938e8_8023,RIde88370_254,RIde83e88_233,RIfc5f420_6106,RIfc976b8_6745,RIfc90a70_6668,RIfc60500_6118,RIee38a40_5103,RIe16ab08_2591,RIe169488_2575,
        RIe166ff8_2549,RIe1642f8_2517,RIe1615f8_2485,RIee369e8_5080,RIe15e8f8_2453,RIee35bd8_5070,RIe15bbf8_2421,RIe1561f8_2357,RIe1534f8_2325,RIfc3ee28_5741,
        RIe1507f8_2293,RIfce6c90_7648,RIe14daf8_2261,RIfcca7c0_7326,RIe14adf8_2229,RIe1480f8_2197,RIe1453f8_2165,RIee33b80_5047,RIee32938_5034,RIee316f0_5021,
        RIee30bb0_5013,RIe1403d0_2108,RIfe93618_8021,RIdf3bfb0_2059,RIfe934b0_8020,RIfcd0d00_7398,RIee2ecc0_4991,RIee2e720_4987,RIee2cb00_4967,RIfe93bb8_8025,
        RIdf32938_1952,RIdf30340_1925,RIdf2e450_1903,RIee2b048_4948,RIee29b30_4933,RIfc67148_6195,RIfc6fb18_6293,RIdf29860_1849,RIfe931e0_8018,RIfe93348_8019,
        RIfe93078_8017,RIfc672b0_6196,RIfca8788_6939,RIdf22510_1767,RIfcea7a0_7690,RIdf20ff8_1752,RIdf1ecd0_1727,RIdf1aab8_1680,RIfea7c58_8225,RIdf15ec8_1626,
        RIdf131c8_1594,RIdf104c8_1562,RIdf0d7c8_1530,RIdf0aac8_1498,RIdf07dc8_1466,RIdf050c8_1434,RIdf023c8_1402,RIdefc9c8_1338,RIdef9cc8_1306,RIdef6fc8_1274,
        RIdef42c8_1242,RIdef15c8_1210,RIdeee8c8_1178,RIdeebbc8_1146,RIdee8ec8_1114,RIee24f40_4879,RIee24130_4869,RIee235f0_4861,RIee22c18_4854,RIfe93d20_8026,
        RIdee1fb0_1035,RIdee0228_1014,RIdeddc30_987,RIfc684f8_6209,RIee21ca0_4843,RIfc68390_6208,RIee20d28_4832,RIded8aa0_929,RIfe93ff0_8028,RIded45b8_880,
        RIfe93e88_8027,RIdecf6f8_824,RIdecc9f8_792,RIdec9cf8_760,RIdec6ff8_728,RIdeb34f8_504,RIde941c0_312,RIe16d100_2618,RIe158ef8_2389,RIe1426f8_2133,
        RIdf370f0_2003,RIdf2b750_1871,RIdf1bfd0_1695,RIdeff6c8_1370,RIdee61c8_1082,RIdedaf30_955,RIde7a108_185,RIe19c590_3156,RIe199890_3124,RIf144f50_5244,
        RIe196b90_3092,RIfc76058_6365,RIe193e90_3060,RIe191190_3028,RIe18e490_2996,RIe188a90_2932,RIe185d90_2900,RIfccd8f8_7361,RIe183090_2868,RIfc76e68_6375,
        RIe180390_2836,RIe17d690_2804,RIe17a990_2772,RIf1419e0_5206,RIf140630_5192,RIe176bb0_2728,RIe1750f8_2709,RIfcd1840_7406,RIfc5f6f0_6108,RIee3dd38_5162,
        RIee3cc58_5150,RIee3b8a8_5136,RIee3a7c8_5124,RIee39580_5111,RIfea9008_8239,RIf16f7f0_5728,RIf16ecb0_5720,RIf16d900_5706,RIfc78ec0_6398,RIfcc8060_7298,
        RIe2228e8_4683,RIfc5a3f8_6049,RIe21fbe8_4651,RIfc74000_6342,RIe21cee8_4619,RIe2174e8_4555,RIe2147e8_4523,RIfca2c20_6874,RIe211ae8_4491,RIfca2950_6872,
        RIe20ede8_4459,RIfcc24f8_7233,RIe20c0e8_4427,RIe2093e8_4395,RIe2066e8_4363,RIfc45110_5808,RIfcc6f80_7286,RIfe92f10_8016,RIfe92970_8012,RIf164af8_5605,
        RIf163a18_5593,RIf162aa0_5582,RIfe92ad8_8013,RIf15f3c8_5543,RIf15d640_5522,RIfe92808_8011,RIfe92c40_8014,RIfe926a0_8010,RIfe92da8_8015,RIfe92538_8009,
        RIfcb5a78_7089,RIf158348_5463,RIf157100_5450,RIfc53be8_5975,RIfec38b8_8345,RIfcc5ea0_7274,RIf1550a8_5427,RIf153cf8_5413,RIfec3a20_8346,RIf152678_5397,
        RIfec3750_8344,RIf14ff18_5369,RIfe923d0_8008,RIf14efa0_5358,RIf14e898_5353,RIf14d380_5338,RIfe92268_8007,RIe1ea650_4044,RIe1e7950_4012,RIe1e4c50_3980,
        RIe1e1f50_3948,RIe1df250_3916,RIe1dc550_3884,RIe1d9850_3852,RIe1d6b50_3820,RIe1d1150_3756,RIe1ce450_3724,RIe1cb750_3692,RIe1c8a50_3660,RIe1c5d50_3628,
        RIe1c3050_3596,RIe1c0350_3564,RIe1bd650_3532,RIfcda4e0_7506,RIfc9d220_6810,RIe1b8628_3475,RIe1b6738_3453,RIfc4f2c8_5923,RIfce16c8_7587,RIfe91cc8_8003,
        RIfe91e30_8004,RIf1484c0_5282,RIf147548_5271,RIfe91f98_8005,RIfe91b60_8002,RIf146b70_5264,RIfc9f548_6835,RIfe92100_8006,RIfe919f8_8001,RIe1a7990_3284,
        RIe1a4c90_3252,RIe1a1f90_3220,RIe19f290_3188,RIe18b790_2964,RIe177c90_2740,RIe2255e8_4715,RIe21a1e8_4587,RIe2039e8_4331,RIe1fda48_4263,RIe1f6e00_4186,
        RIe1ef948_4103,RIe1d3e50_3788,RIe1ba950_3500,RIe1ad7c8_3351,RIe16fe00_2650,RIdec4730_699,RIdec1a30_667,RIfce3f90_7616,RIdebed30_635,RIfcc3308_7243,
        RIdebc030_603,RIdeb9330_571,RIdeb6630_539,RIfc8c588_6619,RIdeb0c30_475,RIfc5a998_6053,RIdeadf30_443,RIfc99b48_6771,RIdea8698_411,RIdea1d98_379,
        RIde9b498_347,RIfc78bf0_6396,RIfcbc558_7165,RIfca12d0_6856,RIfca3fd0_6888,RIfec2670_8332,RIfec2508_8331,RIde88a00_256,RIde84518_235,RIfcc35d8_7245,
        RIfcb57a8_7087,RIfc5a290_6048,RIfca3058_6877,RIee38e78_5106,RIfec27d8_8333,RIfca3328_6879,RIe1672c8_2551,RIe164730_2520,RIe161a30_2488,RIee36cb8_5082,
        RIe15ed30_2456,RIfcc7250_7288,RIe15c030_2424,RIe156630_2360,RIe153930_2328,RIfcc7688_7291,RIe150c30_2296,RIfc8af08_6603,RIe14df30_2264,RIfc9a250_6776,
        RIe14b230_2232,RIe148530_2200,RIe145830_2168,RIfc9aac0_6782,RIfc56bb8_6009,RIfca1ca8_6863,RIfcec960_7714,RIe1406a0_2110,RIdf3e440_2085,RIdf3c280_2061,
        RIdf39f58_2036,RIfc9a958_6781,RIee2f0f8_4994,RIfcdb458_7517,RIee2cf38_4970,RIdf34c60_1977,RIfec2940_8334,RIdf30778_1928,RIdf2e888_1906,RIee2b480_4951,
        RIfec23a0_8330,RIee288e8_4920,RIfec2238_8329,RIdf29b30_1851,RIdf27808_1826,RIdf25a80_1805,RIdf23e60_1785,RIfc55100_5990,RIfcd9f40_7502,RIfc54f98_5989,
        RIfc54cc8_5987,RIfc4b218_5877,RIdf1efa0_1729,RIfcc69e0_7282,RIdf18bc8_1658,RIdf16300_1629,RIdf13600_1597,RIdf10900_1565,RIdf0dc00_1533,RIdf0af00_1501,
        RIdf08200_1469,RIdf05500_1437,RIdf02800_1405,RIdefce00_1341,RIdefa100_1309,RIdef7400_1277,RIdef4700_1245,RIdef1a00_1213,RIdeeed00_1181,RIdeec000_1149,
        RIdee9300_1117,RIfce4ad0_7624,RIfc9e8a0_6826,RIfcc46b8_7257,RIfcd4108_7435,RIdee4440_1061,RIdee2280_1037,RIdee0390_1015,RIdede068_990,RIfcda0a8_7503,
        RIfce54a8_7631,RIfca0790_6848,RIfc50ee8_5943,RIded8d70_931,RIded68e0_905,RIded4888_882,RIded2560_857,RIdecfb30_827,RIdecce30_795,RIdeca130_763,
        RIdec7430_731,RIdeb3930_507,RIde94b98_315,RIe16d538_2621,RIe159330_2392,RIe142b30_2136,RIdf37528_2006,RIdf2bb88_1874,RIdf1c408_1698,RIdeffb00_1373,
        RIdee6600_1085,RIdedb368_958,RIde7aae0_188,RIe19c9c8_3159,RIe199cc8_3127,RIfe8ea28_7967,RIe196fc8_3095,RIfec20d0_8328,RIe1942c8_3063,RIe1915c8_3031,
        RIe18e8c8_2999,RIe188ec8_2935,RIe1861c8_2903,RIfc68228_6207,RIe1834c8_2871,RIfccb5d0_7336,RIe1807c8_2839,RIe17dac8_2807,RIe17adc8_2775,RIf141e18_5209,
        RIf140900_5194,RIf140090_5188,RIe1753c8_2711,RIf13f988_5183,RIf13ece0_5174,RIee3e170_5165,RIee3cf28_5152,RIee3bce0_5139,RIee3ac00_5127,RIee39850_5113,
        RIe172dd0_2684,RIf16fc28_5731,RIf16f0e8_5723,RIf16dd38_5709,RIfce9120_7674,RIfc404a8_5757,RIe222d20_4686,RIf16b8a8_5683,RIe220020_4654,RIf16a930_5672,
        RIe21d320_4622,RIe217920_4558,RIe214c20_4526,RIfc5b910_6064,RIe211f20_4494,RIfe8e8c0_7966,RIe20f220_4462,RIfe8e758_7965,RIe20c520_4430,RIe209820_4398,
        RIe206b20_4366,RIf166b50_5628,RIf165a70_5616,RIfe8dd80_7958,RIfe8dab0_7956,RIf164c60_5606,RIf163e50_5596,RIf162ed8_5585,RIf1616f0_5568,RIf15f800_5546,
        RIf15da78_5525,RIfe8d948_7955,RIfe8dc18_7957,RIf15c560_5510,RIf15b048_5495,RIfc62828_6143,RIf159860_5478,RIf158780_5466,RIf157538_5453,RIfca6e38_6921,
        RIe1f9b00_4218,RIfc61e50_6136,RIfc61748_6131,RIf154130_5416,RIe1f4ad8_4161,RIf152ab0_5400,RIf151700_5386,RIf1501e8_5371,RIe1f27b0_4136,RIfc60ed8_6125,
        RIfc7b620_6426,RIf14d7b8_5341,RIe1ed4b8_4077,RIe1eaa88_4047,RIe1e7d88_4015,RIe1e5088_3983,RIe1e2388_3951,RIe1df688_3919,RIe1dc988_3887,RIe1d9c88_3855,
        RIe1d6f88_3823,RIe1d1588_3759,RIe1ce888_3727,RIe1cbb88_3695,RIe1c8e88_3663,RIe1c6188_3631,RIe1c3488_3599,RIe1c0788_3567,RIe1bda88_3535,RIfca4de0_6898,
        RIfc5ea48_6099,RIe1b8a60_3478,RIe1b6a08_3455,RIfcbd638_7177,RIfc44fa8_5807,RIfe8e5f0_7964,RIfe8e1b8_7961,RIf1488f8_5285,RIf147818_5273,RIfe8e050_7960,
        RIfe8e488_7963,RIf146e40_5266,RIf146030_5256,RIfe8dee8_7959,RIfe8e320_7962,RIe1a7dc8_3287,RIe1a50c8_3255,RIe1a23c8_3223,RIe19f6c8_3191,RIe18bbc8_2967,
        RIe1780c8_2743,RIe225a20_4718,RIe21a620_4590,RIe203e20_4334,RIe1fde80_4266,RIe1f7238_4189,RIe1efd80_4106,RIe1d4288_3791,RIe1bad88_3503,RIe1adc00_3354,
        RIe170238_2653,RIdec45c8_698,RIdec18c8_666,RIfce85e0_7666,RIdebebc8_634,RIfcb8bb0_7124,RIdebbec8_602,RIdeb91c8_570,RIdeb64c8_538,RIfc85d78_6545,
        RIdeb0ac8_474,RIfc85aa8_6543,RIdeaddc8_442,RIfc4d3d8_5901,RIdea8350_410,RIdea1a50_378,RIde9b150_346,RIfc85ee0_6546,RIfc9c9b0_6804,RIfce13f8_7585,
        RIfcb8778_7121,RIfe8d510_7952,RIfe8d3a8_7951,RIde886b8_255,RIde841d0_234,RIde806c0_216,RIfcb8070_7116,RIfce1128_7583,RIfc9c140_6798,RIee38d10_5105,
        RIe16ac70_2592,RIfc850d0_6536,RIe167160_2550,RIe1645c8_2519,RIe1618c8_2487,RIee36b50_5081,RIe15ebc8_2455,RIee35d40_5071,RIe15bec8_2423,RIe1564c8_2359,
        RIe1537c8_2327,RIfc3ef90_5742,RIe150ac8_2295,RIfe8d7e0_7954,RIe14ddc8_2263,RIfce0fc0_7582,RIe14b0c8_2231,RIe1483c8_2199,RIe1456c8_2167,RIee33e50_5049,
        RIee32c08_5036,RIee319c0_5023,RIee30d18_5014,RIfe8cf70_7948,RIfe8ce08_7947,RIfe8d240_7950,RIfe8d0d8_7949,RIfce9dc8_7683,RIee2ef90_4993,RIfce51d8_7629,
        RIee2cdd0_4969,RIdf34af8_1976,RIfe8d678_7953,RIdf30610_1927,RIdf2e720_1905,RIee2b318_4950,RIee29c98_4934,RIee28780_4919,RIee27538_4906,RIdf299c8_1850,
        RIdf276a0_1825,RIdf25918_1804,RIdf23cf8_1784,RIfc83ff0_6524,RIfcb73c8_7107,RIfc51320_5946,RIfcdaa80_7510,RIfc83d20_6522,RIdf1ee38_1728,RIfc51b90_5952,
        RIdf18a60_1657,RIdf16198_1628,RIdf13498_1596,RIdf10798_1564,RIdf0da98_1532,RIdf0ad98_1500,RIdf08098_1468,RIdf05398_1436,RIdf02698_1404,RIdefcc98_1340,
        RIdef9f98_1308,RIdef7298_1276,RIdef4598_1244,RIdef1898_1212,RIdeeeb98_1180,RIdeebe98_1148,RIdee9198_1116,RIee25210_4881,RIee24400_4871,RIee238c0_4863,
        RIee22ee8_4856,RIfe8cca0_7946,RIdee2118_1036,RIfe8cb38_7945,RIdeddf00_989,RIfcc5a68_7271,RIee21f70_4845,RIfcb6cc0_7102,RIee20e90_4833,RIded8c08_930,
        RIded6778_904,RIded4720_881,RIded23f8_856,RIdecf9c8_826,RIdecccc8_794,RIdec9fc8_762,RIdec72c8_730,RIdeb37c8_506,RIde94850_314,RIe16d3d0_2620,
        RIe1591c8_2391,RIe1429c8_2135,RIdf373c0_2005,RIdf2ba20_1873,RIdf1c2a0_1697,RIdeff998_1372,RIdee6498_1084,RIdedb200_957,RIde7a798_187,RIe19c860_3158,
        RIe199b60_3126,RIf145220_5246,RIe196e60_3094,RIf144140_5234,RIe194160_3062,RIe191460_3030,RIe18e760_2998,RIe188d60_2934,RIe186060_2902,RIf1431c8_5223,
        RIe183360_2870,RIf142ac0_5218,RIe180660_2838,RIe17d960_2806,RIe17ac60_2774,RIf141cb0_5208,RIf140798_5193,RIf13ff28_5187,RIfe8be90_7936,RIfceb880_7702,
        RIf13eb78_5173,RIee3e008_5164,RIee3cdc0_5151,RIee3bb78_5138,RIee3aa98_5126,RIee396e8_5112,RIe172c68_2683,RIf16fac0_5730,RIf16ef80_5722,RIf16dbd0_5708,
        RIfcc4af0_7260,RIf16c820_5694,RIe222bb8_4685,RIf16b740_5682,RIe21feb8_4653,RIf16a7c8_5671,RIe21d1b8_4621,RIe2177b8_4557,RIe214ab8_4525,RIfe8c430_7940,
        RIe211db8_4493,RIf1688d8_5649,RIe20f0b8_4461,RIf167960_5638,RIe20c3b8_4429,RIe2096b8_4397,RIe2069b8_4365,RIf1669e8_5627,RIf165908_5615,RIfe8c9d0_7944,
        RIfe8c700_7942,RIfc9c578_6801,RIf163ce8_5595,RIf162d70_5584,RIf161588_5567,RIf15f698_5545,RIf15d910_5524,RIfe8c598_7941,RIfe8c868_7943,RIf15c3f8_5509,
        RIf15aee0_5494,RIf15a0d0_5484,RIf1596f8_5477,RIf158618_5465,RIf1573d0_5452,RIf156b60_5446,RIfec1f68_8327,RIf155eb8_5437,RIf155378_5429,RIf153fc8_5415,
        RIfe8bff8_7937,RIf152948_5399,RIf151598_5385,RIf150080_5370,RIfe8c2c8_7939,RIf14f270_5360,RIfc503a8_5935,RIf14d650_5340,RIfe8c160_7938,RIe1ea920_4046,
        RIe1e7c20_4014,RIe1e4f20_3982,RIe1e2220_3950,RIe1df520_3918,RIe1dc820_3886,RIe1d9b20_3854,RIe1d6e20_3822,RIe1d1420_3758,RIe1ce720_3726,RIe1cba20_3694,
        RIe1c8d20_3662,RIe1c6020_3630,RIe1c3320_3598,RIe1c0620_3566,RIe1bd920_3534,RIf14c2a0_5326,RIf14aef0_5312,RIe1b88f8_3477,RIe1b68a0_3454,RIfcd4db0_7444,
        RIfc4ebc0_5918,RIfec1e00_8326,RIfe8bd28_7935,RIf148790_5284,RIf1476b0_5272,RIfe8ba58_7933,RIfec1b30_8324,RIfc4e788_5915,RIfcb8e80_7126,RIfe8bbc0_7934,
        RIfec1c98_8325,RIe1a7c60_3286,RIe1a4f60_3254,RIe1a2260_3222,RIe19f560_3190,RIe18ba60_2966,RIe177f60_2742,RIe2258b8_4717,RIe21a4b8_4589,RIe203cb8_4333,
        RIe1fdd18_4265,RIe1f70d0_4188,RIe1efc18_4105,RIe1d4120_3790,RIe1bac20_3502,RIe1ada98_3353,RIe1700d0_2652,RIdec4a00_701,RIdec1d00_669,RIfcad7b0_6996,
        RIdebf000_637,RIfc64cb8_6169,RIdebc300_605,RIdeb9600_573,RIdeb6900_541,RIfc6f9b0_6292,RIdeb0f00_477,RIfc657f8_6177,RIdeae200_445,RIfce69c0_7646,
        RIdea8d28_413,RIdea2428_381,RIde9bb28_349,RIfc6fc80_6294,RIee1b760_4771,RIfca8080_6934,RIfe8b8f0_7932,RIde90020_292,RIde8c510_274,RIde89090_258,
        RIde84ba8_237,RIfc65ac8_6179,RIfcad210_6992,RIfcce168_7367,RIfcce2d0_7368,RIfc51488_5947,RIe16af40_2594,RIfc65c30_6180,RIe167598_2553,RIe164a00_2522,
        RIe161d00_2490,RIfc66e78_6193,RIe15f000_2458,RIfc6e498_6277,RIe15c300_2426,RIe156900_2362,RIe153c00_2330,RIfc6e330_6276,RIe150f00_2298,RIfccda60_7362,
        RIe14e200_2266,RIfc6e1c8_6275,RIe14b500_2234,RIe148800_2202,RIe145b00_2170,RIee33fb8_5050,RIee32d70_5037,RIee31c90_5025,RIee30fe8_5016,RIfea8630_8232,
        RIdf3e5a8_2086,RIdf3c550_2063,RIfea8798_8233,RIfc6e060_6274,RIfcac6d0_6984,RIfc56078_6001,RIfc6e600_6278,RIdf34dc8_1978,RIdf32d70_1955,RIfea84c8_8231,
        RIdf2eb58_1908,RIee2b750_4953,RIfc6ee70_6284,RIfc6efd8_6285,RIee27808_4908,RIfe8b788_7931,RIdf27ad8_1828,RIdf25d50_1807,RIdf24130_1787,RIfc66608_6187,
        RIfccde98_7365,RIfc66a40_6190,RIfc668d8_6189,RIfcacf40_6990,RIfeaaef8_8261,RIfc6e8d0_6280,RIdf18d30_1659,RIdf165d0_1631,RIdf138d0_1599,RIdf10bd0_1567,
        RIdf0ded0_1535,RIdf0b1d0_1503,RIdf084d0_1471,RIdf057d0_1439,RIdf02ad0_1407,RIdefd0d0_1343,RIdefa3d0_1311,RIdef76d0_1279,RIdef49d0_1247,RIdef1cd0_1215,
        RIdeeefd0_1183,RIdeec2d0_1151,RIdee95d0_1119,RIfc6dc28_6271,RIfc67c88_6203,RIfccb300_7334,RIfccd4c0_7358,RIfea81f8_8229,RIfea8360_8230,RIdee04f8_1016,
        RIdede338_992,RIfc6def8_6273,RIfcac130_6980,RIfc67b20_6202,RIfc67df0_6204,RIded9040_933,RIded6a48_906,RIded4b58_884,RIded26c8_858,RIdecfe00_829,
        RIdecd100_797,RIdeca400_765,RIdec7700_733,RIdeb3c00_509,RIde95228_317,RIe16d808_2623,RIe159600_2394,RIe142e00_2138,RIdf377f8_2008,RIdf2be58_1876,
        RIdf1c6d8_1700,RIdeffdd0_1375,RIdee68d0_1087,RIdedb638_960,RIde7b170_190,RIe19cc98_3161,RIe199f98_3129,RIfc73088_6331,RIe197298_3097,RIf1442a8_5235,
        RIe194598_3065,RIe191898_3033,RIe18eb98_3001,RIe189198_2937,RIe186498_2905,RIfc72278_6321,RIe183798_2873,RIfc61ce8_6135,RIe180a98_2841,RIe17dd98_2809,
        RIe17b098_2777,RIfcaf268_7015,RIfca6a00_6918,RIfcc9b18_7317,RIe175530_2712,RIfc72818_6325,RIfc726b0_6324,RIfccf7e8_7383,RIfc72548_6323,RIee3be48_5140,
        RIee3ad68_5128,RIfc71fa8_6319,RIe1730a0_2686,RIfcaef98_7013,RIfccf518_7381,RIfc71e40_6318,RIfc62120_6138,RIfe8b350_7928,RIe222ff0_4688,RIfcc9f50_7320,
        RIe2202f0_4656,RIfc4a570_5868,RIe21d5f0_4624,RIe217bf0_4560,RIe214ef0_4528,RIfccf3b0_7380,RIe2121f0_4496,RIf168ba8_5651,RIe20f4f0_4464,RIfc71300_6310,
        RIe20c7f0_4432,RIe209af0_4400,RIe206df0_4368,RIfc718a0_6314,RIfc71a08_6315,RIe202098_4313,RIfe8b1e8_7927,RIfc715d0_6312,RIfce6588_7643,RIfc62c60_6146,
        RIf161858_5569,RIf15fad0_5548,RIf15dbe0_5526,RIe1fc698_4249,RIfe8b4b8_7929,RIfcae5c0_7006,RIfc63098_6149,RIfc63200_6150,RIfc71198_6309,RIf158a50_5468,
        RIf1576a0_5454,RIfcdc808_7531,RIfe8b620_7930,RIfc634d0_6152,RIfcceb40_7374,RIf154400_5418,RIe1f4da8_4163,RIf152c18_5401,RIf151868_5387,RIfc4d108_5899,
        RIe1f2a80_4138,RIfc70a90_6304,RIfc63bd8_6157,RIfca7810_6928,RIe1ed788_4079,RIe1ead58_4049,RIe1e8058_4017,RIe1e5358_3985,RIe1e2658_3953,RIe1df958_3921,
        RIe1dcc58_3889,RIe1d9f58_3857,RIe1d7258_3825,RIe1d1858_3761,RIe1ceb58_3729,RIe1cbe58_3697,RIe1c9158_3665,RIe1c6458_3633,RIe1c3758_3601,RIe1c0a58_3569,
        RIe1bdd58_3537,RIf14c408_5327,RIf14b1c0_5314,RIe1b8d30_3480,RIe1b6cd8_3457,RIfc707c0_6302,RIfca7c48_6931,RIe1b4de8_3435,RIe1b3a38_3421,RIfc70220_6298,
        RIfcce870_7372,RIe1b23b8_3405,RIe1b0630_3384,RIfc645b0_6164,RIfc700b8_6297,RIfeaac28_8259,RIe1aa690_3316,RIe1a8098_3289,RIe1a5398_3257,RIe1a2698_3225,
        RIe19f998_3193,RIe18be98_2969,RIe178398_2745,RIe225cf0_4720,RIe21a8f0_4592,RIe2040f0_4336,RIe1fe150_4268,RIe1f7508_4191,RIe1f0050_4108,RIe1d4558_3793,
        RIe1bb058_3505,RIe1aded0_3356,RIe170508_2655,RIdec4898_700,RIdec1b98_668,RIfc661d0_6184,RIdebee98_636,RIfce6b28_7647,RIdebc198_604,RIdeb9498_572,
        RIdeb6798_540,RIfc40d18_5763,RIdeb0d98_476,RIfcad648_6995,RIdeae098_444,RIfcaa510_6960,RIdea89e0_412,RIdea20e0_380,RIde9b7e0_348,RIfcab320_6970,
        RIfca8350_6936,RIfc6f6e0_6290,RIfcaa240_6958,RIde8fcd8_291,RIfe8aae0_7922,RIde88d48_257,RIde84860_236,RIde80a08_217,RIfc64718_6165,RIfcae020_7002,
        RIfcadeb8_7001,RIee38fe0_5107,RIe16add8_2593,RIe1695f0_2576,RIe167430_2552,RIe164898_2521,RIe161b98_2489,RIfe8a3d8_7917,RIe15ee98_2457,RIfe8a270_7916,
        RIe15c198_2425,RIe156798_2361,RIe153a98_2329,RIfc3f0f8_5743,RIe150d98_2297,RIfcab050_6968,RIe14e098_2265,RIfcca658_7325,RIe14b398_2233,RIe148698_2201,
        RIe145998_2169,RIfe8a810_7920,RIfe8a6a8_7919,RIee31b28_5024,RIee30e80_5015,RIe140808_2111,RIfe8a540_7918,RIdf3c3e8_2062,RIdf3a0c0_2037,RIfc6b1f8_6241,
        RIee2f260_4995,RIfc70d60_6306,RIee2d0a0_4971,RIfe8a978_7921,RIdf32c08_1954,RIdf308e0_1929,RIdf2e9f0_1907,RIee2b5e8_4952,RIee29e00_4935,RIee28a50_4921,
        RIee276a0_4907,RIdf29c98_1852,RIdf27970_1827,RIdf25be8_1806,RIdf23fc8_1786,RIfc6aaf0_6236,RIfc6ac58_6237,RIdf22678_1768,RIfcdd4b0_7540,RIdf21160_1753,
        RIdf1f108_1730,RIdf1ac20_1681,RIfeaa7f0_8256,RIdf16468_1630,RIdf13768_1598,RIdf10a68_1566,RIdf0dd68_1534,RIdf0b068_1502,RIdf08368_1470,RIdf05668_1438,
        RIdf02968_1406,RIdefcf68_1342,RIdefa268_1310,RIdef7568_1278,RIdef4868_1246,RIdef1b68_1214,RIdeeee68_1182,RIdeec168_1150,RIdee9468_1118,RIee25378_4882,
        RIee24568_4872,RIee23a28_4864,RIee23050_4857,RIfe8adb0_7924,RIdee23e8_1038,RIfe8ac48_7923,RIdede1d0_991,RIfca5650_6904,RIee220d8_4846,RIfceeb20_7738,
        RIee20ff8_4834,RIded8ed8_932,RIfe8af18_7925,RIded49f0_883,RIfe8b080_7926,RIdecfc98_828,RIdeccf98_796,RIdeca298_764,RIdec7598_732,RIdeb3a98_508,
        RIde94ee0_316,RIe16d6a0_2622,RIe159498_2393,RIe142c98_2137,RIdf37690_2007,RIdf2bcf0_1875,RIdf1c570_1699,RIdeffc68_1374,RIdee6768_1086,RIdedb4d0_959,
        RIde7ae28_189,RIe19cb30_3160,RIe199e30_3128,RIf145388_5247,RIe197130_3096,RIfe8a108_7915,RIe194430_3064,RIe191730_3032,RIe18ea30_3000,RIe189030_2936,
        RIe186330_2904,RIfc6c878_6257,RIe183630_2872,RIfcabcf8_6977,RIe180930_2840,RIe17dc30_2808,RIe17af30_2776,RIfcccc50_7352,RIfcccdb8_7353,RIe176d18_2729,
        RIfea7af0_8224,RIfe89fa0_7914,RIfe89e38_7913,RIfcdd078_7537,RIfccb738_7337,RIfca9868_6951,RIfcabb90_6976,RIfca99d0_6952,RIe172f38_2685,RIf16fd90_5732,
        RIf16f250_5724,RIfc6c440_6254,RIfcaba28_6975,RIfc40610_5758,RIe222e88_4687,RIfc5d260_6082,RIe220188_4655,RIfcab758_6973,RIe21d488_4623,RIe217a88_4559,
        RIe214d88_4527,RIfe892f8_7905,RIe212088_4495,RIf168a40_5650,RIe20f388_4463,RIf167ac8_5639,RIe20c688_4431,RIe209988_4399,RIe206c88_4367,RIfc6c2d8_6253,
        RIfceec88_7739,RIe201f30_4312,RIe200748_4295,RIf164dc8_5607,RIf163fb8_5597,RIf163040_5586,RIfe895c8_7907,RIf15f968_5547,RIfe89898_7909,RIfe89460_7906,
        RIe1fb5b8_4237,RIf15c6c8_5511,RIfe89730_7908,RIf15a238_5485,RIf1599c8_5479,RIf1588e8_5467,RIfe89cd0_7912,RIfc5ba78_6065,RIe1f9c68_4219,RIfc5bd48_6067,
        RIf1554e0_5430,RIf154298_5417,RIe1f4c40_4162,RIfe89b68_7911,RIfe89a00_7910,RIf150350_5372,RIe1f2918_4137,RIf14f3d8_5361,RIfccc818_7349,RIf14d920_5342,
        RIe1ed620_4078,RIe1eabf0_4048,RIe1e7ef0_4016,RIe1e51f0_3984,RIe1e24f0_3952,RIe1df7f0_3920,RIe1dcaf0_3888,RIe1d9df0_3856,RIe1d70f0_3824,RIe1d16f0_3760,
        RIe1ce9f0_3728,RIe1cbcf0_3696,RIe1c8ff0_3664,RIe1c62f0_3632,RIe1c35f0_3600,RIe1c08f0_3568,RIe1bdbf0_3536,RIfc680c0_6206,RIf14b058_5313,RIe1b8bc8_3479,
        RIe1b6b70_3456,RIfcac298_6981,RIf1499d8_5297,RIfe89190_7904,RIfec19c8_8323,RIf148a60_5286,RIfccdd30_7364,RIe1b2250_3404,RIfec1860_8322,RIfc6e768_6279,
        RIfc54728_5983,RIe1abfe0_3334,RIe1aa528_3315,RIe1a7f30_3288,RIe1a5230_3256,RIe1a2530_3224,RIe19f830_3192,RIe18bd30_2968,RIe178230_2744,RIe225b88_4719,
        RIe21a788_4591,RIe203f88_4335,RIe1fdfe8_4267,RIe1f73a0_4190,RIe1efee8_4107,RIe1d43f0_3792,RIe1baef0_3504,RIe1add68_3355,RIe1703a0_2654,RIdec4cd0_703,
        RIdec1fd0_671,RIfc7b4b8_6425,RIdebf2d0_639,RIfc7b1e8_6423,RIdebc5d0_607,RIdeb98d0_575,RIdeb6bd0_543,RIfe83358_7837,RIdeb11d0_479,RIee1e5c8_4804,
        RIdeae4d0_447,RIfc437c0_5790,RIdea93b8_415,RIdea2ab8_383,RIde9c1b8_351,RIfc90ea8_6671,RIfc7af18_6421,RIfe83088_7835,RIee1a950_4761,RIde906b0_294,
        RIde8cba0_276,RIfe82f20_7834,RIfe82db8_7833,RIee1a248_4756,RIfe831f0_7836,RIfcc2390_7232,RIee195a0_4747,RIfcbe718_7189,RIfea9e18_8249,RIfc43220_5786,
        RIe167868_2555,RIe164cd0_2524,RIe161fd0_2492,RIee36f88_5084,RIe15f2d0_2460,RIee35ea8_5072,RIe15c5d0_2428,RIe156bd0_2364,RIe153ed0_2332,RIfe83628_7839,
        RIe1511d0_2300,RIfebfda8_8303,RIe14e4d0_2268,RIfebfc40_8302,RIe14b7d0_2236,RIe148ad0_2204,RIe145dd0_2172,RIee34120_5051,RIee32ed8_5038,RIee31df8_5026,
        RIfcc1f58_7229,RIe140ad8_2113,RIdf3e878_2088,RIfe834c0_7838,RIdf3a390_2039,RIfc5a6c8_6051,RIfc91e20_6682,RIee2e888_4988,RIfc96a10_6736,RIdf35098_1980,
        RIfeab600_8266,RIdf30bb0_1931,RIfeab768_8267,RIfcbe9e8_7191,RIfc79fa0_6410,RIfc96740_6734,RIfc92258_6685,RIfea7118_8217,RIfea95a8_8243,RIdf26020_1809,
        RIdf24400_1789,RIfc79a00_6406,RIfc5add0_6056,RIfce5d18_7637,RIfc92690_6688,RIfce3018_7605,RIdf1f270_1731,RIfc79730_6404,RIdf19000_1661,RIdf168a0_1633,
        RIdf13ba0_1601,RIdf10ea0_1569,RIdf0e1a0_1537,RIdf0b4a0_1505,RIdf087a0_1473,RIdf05aa0_1441,RIdf02da0_1409,RIdefd3a0_1345,RIdefa6a0_1313,RIdef79a0_1281,
        RIdef4ca0_1249,RIdef1fa0_1217,RIdeef2a0_1185,RIdeec5a0_1153,RIdee98a0_1121,RIfc5b7a8_6063,RIfc5b640_6062,RIfc931d0_6696,RIfcecac8_7715,RIdee4710_1063,
        RIdee26b8_1040,RIdee07c8_1018,RIdede4a0_993,RIfcbf0f0_7196,RIfcbf528_7199,RIfc792f8_6401,RIfc93068_6695,RIded91a8_934,RIded6d18_908,RIded4e28_886,
        RIded2998_860,RIded00d0_831,RIdecd3d0_799,RIdeca6d0_767,RIdec79d0_735,RIdeb3ed0_511,RIde958b8_319,RIe16dad8_2625,RIe1598d0_2396,RIe1430d0_2140,
        RIdf37ac8_2010,RIdf2c128_1878,RIdf1c9a8_1702,RIdf000a0_1377,RIdee6ba0_1089,RIdedb908_962,RIde7b800_192,RIe19cf68_3163,RIe19a268_3131,RIfc8d7d0_6632,
        RIe197568_3099,RIfc561e0_6002,RIe194868_3067,RIe191b68_3035,RIe18ee68_3003,RIe189468_2939,RIe186768_2907,RIf143330_5224,RIe183a68_2875,RIfc7d948_6451,
        RIe180d68_2843,RIe17e068_2811,RIe17b368_2779,RIfc564b0_6004,RIfcd6700_7462,RIfc461f0_5820,RIe175698_2713,RIfc46088_5819,RIfc45f20_5818,RIfc7dc18_6453,
        RIfcd69d0_7464,RIfc98630_6756,RIfcc2a98_7237,RIfc7d510_6448,RIe173208_2687,RIfc8e478_6641,RIfc45ae8_5815,RIfc8e8b0_6644,RIfc45980_5814,RIfe82ae8_7831,
        RIe2232c0_4690,RIf16ba10_5684,RIe2205c0_4658,RIfcd24e8_7415,RIe21d8c0_4626,RIe217ec0_4562,RIe2151c0_4530,RIfebf268_8295,RIe2124c0_4498,RIf168d10_5652,
        RIe20f7c0_4466,RIfc7d240_6446,RIe20cac0_4434,RIe209dc0_4402,RIe2070c0_4370,RIf166e20_5630,RIfebf6a0_8298,RIfebf808_8299,RIfebf538_8297,RIfc8eb80_6646,
        RIf164120_5598,RIfc453e0_5810,RIf161b28_5571,RIf15fc38_5549,RIf15dd48_5527,RIe1fc968_4251,RIe1fb888_4239,RIfebf3d0_8296,RIf15b318_5497,RIfca2518_6869,
        RIfc8f120_6650,RIfebfad8_8301,RIfebf970_8300,RIfc7cca0_6442,RIe1f9dd0_4220,RIfe82c50_7832,RIf155648_5431,RIfc8f288_6651,RIe1f4f10_4164,RIf152d80_5402,
        RIfc8f828_6655,RIfcb3b88_7067,RIe1f2d50_4140,RIfc445d0_5800,RIfc8faf8_6657,RIf14da88_5343,RIe1eda58_4081,RIe1eb028_4051,RIe1e8328_4019,RIe1e5628_3987,
        RIe1e2928_3955,RIe1dfc28_3923,RIe1dcf28_3891,RIe1da228_3859,RIe1d7528_3827,RIe1d1b28_3763,RIe1cee28_3731,RIe1cc128_3699,RIe1c9428_3667,RIe1c6728_3635,
        RIe1c3a28_3603,RIe1c0d28_3571,RIe1be028_3539,RIfc7bff8_6433,RIfc44030_5796,RIe1b9000_3482,RIe1b6fa8_3459,RIfcbdd40_7182,RIfc8ff30_6660,RIe1b50b8_3437,
        RIe1b3d08_3423,RIfcbe178_7185,RIfc43d60_5794,RIe1b2520_3406,RIe1b0798_3385,RIfcdb5c0_7518,RIfc7ba58_6429,RIe1ac148_3335,RIe1aa960_3318,RIe1a8368_3291,
        RIe1a5668_3259,RIe1a2968_3227,RIe19fc68_3195,RIe18c168_2971,RIe178668_2747,RIe225fc0_4722,RIe21abc0_4594,RIe2043c0_4338,RIe1fe420_4270,RIe1f77d8_4193,
        RIe1f0320_4110,RIe1d4828_3795,RIe1bb328_3507,RIe1ae1a0_3358,RIe1707d8_2657,RIdec4b68_702,RIdec1e68_670,RIfc5df08_6091,RIdebf168_638,RIfce6df8_7649,
        RIdebc468_606,RIdeb9768_574,RIdeb6a68_542,RIfc75ef0_6364,RIdeb1068_478,RIfcc12b0_7220,RIdeae368_446,RIfc5e340_6094,RIdea9070_414,RIdea2770_382,
        RIde9be70_350,RIfced4a0_7722,RIfcc1418_7221,RIfc95930_6724,RIfcec0f0_7708,RIde90368_293,RIde8c858_275,RIde893d8_259,RIde84ef0_238,RIde80d50_218,
        RIfc95a98_6725,RIfced068_7719,RIfced1d0_7720,RIfcedfe0_7730,RIe16b0a8_2595,RIe169758_2577,RIe167700_2554,RIe164b68_2523,RIe161e68_2491,RIee36e20_5083,
        RIe15f168_2459,RIfc426e0_5778,RIe15c468_2427,RIe156a68_2363,RIe153d68_2331,RIfe82818_7829,RIe151068_2299,RIee34c60_5059,RIe14e368_2267,RIfc5f9c0_6110,
        RIe14b668_2235,RIe148968_2203,RIe145c68_2171,RIfccfef0_7388,RIfca57b8_6905,RIfc600c8_6115,RIfcafda8_7023,RIe140970_2112,RIdf3e710_2087,RIdf3c6b8_2064,
        RIdf3a228_2038,RIfc5fc90_6112,RIee2f3c8_4996,RIfc742d0_6344,RIee2d208_4972,RIdf34f30_1979,RIfebf100_8294,RIdf30a48_1930,RIdf2ecc0_1909,RIfcb08e8_7031,
        RIfcee418_7733,RIfc95ed0_6728,RIfcdef68_7559,RIdf29e00_1853,RIdf27c40_1829,RIdf25eb8_1808,RIdf24298_1788,RIfc5ed18_6101,RIfcee850_7736,RIdf227e0_1769,
        RIfc5efe8_6103,RIdf212c8_1754,RIfeaa520_8254,RIdf1ad88_1682,RIdf18e98_1660,RIdf16738_1632,RIdf13a38_1600,RIdf10d38_1568,RIdf0e038_1536,RIdf0b338_1504,
        RIdf08638_1472,RIdf05938_1440,RIdf02c38_1408,RIdefd238_1344,RIdefa538_1312,RIdef7838_1280,RIdef4b38_1248,RIdef1e38_1216,RIdeef138_1184,RIdeec438_1152,
        RIdee9738_1120,RIfcc96e0_7314,RIfccfd88_7387,RIfc60aa0_6122,RIfca5ec0_6910,RIdee45a8_1062,RIdee2550_1039,RIdee0660_1017,RIfe826b0_7828,RIfcdeb30_7556,
        RIfc73bc8_6339,RIfca5bf0_6908,RIfc73a60_6338,RIfe82980_7830,RIded6bb0_907,RIded4cc0_885,RIded2830_859,RIdecff68_830,RIdecd268_798,RIdeca568_766,
        RIdec7868_734,RIdeb3d68_510,RIde95570_318,RIe16d970_2624,RIe159768_2395,RIe142f68_2139,RIdf37960_2009,RIdf2bfc0_1877,RIdf1c840_1701,RIdefff38_1376,
        RIdee6a38_1088,RIdedb7a0_961,RIde7b4b8_191,RIe19ce00_3162,RIe19a100_3130,RIfce96c0_7678,RIe197400_3098,RIf144410_5236,RIe194700_3066,RIe191a00_3034,
        RIe18ed00_3002,RIe189300_2938,RIe186600_2906,RIfebee30_8292,RIe183900_2874,RIfcdbcc8_7523,RIe180c00_2842,RIe17df00_2810,RIe17b200_2778,RIf141f80_5210,
        RIfce7398_7653,RIfcb1e00_7046,RIfe82548_7827,RIfca42a0_6890,RIfcbff00_7206,RIfcaaee8_6967,RIee3d090_5153,RIfc5c180_6070,RIfce35b8_7609,RIee399b8_5114,
        RIfea8a68_8235,RIf16fef8_5733,RIfebecc8_8291,RIfc5c450_6072,RIfce9288_7675,RIfc40778_5759,RIe223158_4689,RIfce77d0_7656,RIe220458_4657,RIfce24d8_7597,
        RIe21d758_4625,RIe217d58_4561,RIe215058_4529,RIfce8a18_7669,RIe212358_4497,RIfce1998_7589,RIe20f658_4465,RIfc77840_6382,RIe20c958_4433,RIe209c58_4401,
        RIe206f58_4369,RIf166cb8_5629,RIf165bd8_5617,RIfe81fa8_7823,RIfe81e40_7822,RIfc5c888_6075,RIfceb178_7697,RIf1631a8_5587,RIf1619c0_5570,RIfccf248_7379,
        RIfc77570_6380,RIe1fc800_4250,RIe1fb720_4238,RIf15c830_5512,RIf15b1b0_5496,RIfcd0fd0_7400,RIfccc6b0_7348,RIf158bb8_5469,RIf157808_5455,RIfc5d0f8_6081,
        RIfebef98_8293,RIfcc8a38_7305,RIfcd7ab0_7476,RIfcb1428_7039,RIfeaa0e8_8251,RIfccc548_7347,RIfce3450_7608,RIf1504b8_5373,RIe1f2be8_4139,RIf14f540_5362,
        RIfc772a0_6378,RIfcec258_7709,RIe1ed8f0_4080,RIe1eaec0_4050,RIe1e81c0_4018,RIe1e54c0_3986,RIe1e27c0_3954,RIe1dfac0_3922,RIe1dcdc0_3890,RIe1da0c0_3858,
        RIe1d73c0_3826,RIe1d19c0_3762,RIe1cecc0_3730,RIe1cbfc0_3698,RIe1c92c0_3666,RIe1c65c0_3634,RIe1c38c0_3602,RIe1c0bc0_3570,RIe1bdec0_3538,RIf14c570_5328,
        RIf14b328_5315,RIe1b8e98_3481,RIe1b6e40_3458,RIfc76760_6370,RIfc94b20_6714,RIe1b4f50_3436,RIe1b3ba0_3422,RIfcec3c0_7710,RIfceb010_7696,RIfe823e0_7826,
        RIfe82110_7824,RIfcdd8e8_7543,RIfcc0ba8_7215,RIfe82278_7825,RIe1aa7f8_3317,RIe1a8200_3290,RIe1a5500_3258,RIe1a2800_3226,RIe19fb00_3194,RIe18c000_2970,
        RIe178500_2746,RIe225e58_4721,RIe21aa58_4593,RIe204258_4337,RIe1fe2b8_4269,RIe1f7670_4192,RIe1f01b8_4109,RIe1d46c0_3794,RIe1bb1c0_3506,RIe1ae038_3357,
        RIe170670_2656,RIdec4fa0_705,RIdec22a0_673,RIee1fdb0_4821,RIdebf5a0_641,RIee1f270_4813,RIdebc8a0_609,RIdeb9ba0_577,RIdeb6ea0_545,RIee1ecd0_4809,
        RIdeb14a0_481,RIee1e730_4805,RIdeae7a0_449,RIee1d920_4795,RIdea9a48_417,RIdea3148_385,RIde9c848_353,RIee1cb10_4785,RIee1ba30_4773,RIee1b1c0_4767,
        RIfec04b0_8308,RIfe850e0_7858,RIde8d230_278,RIfea9cb0_8248,RIfe84f78_7857,RIee1a3b0_4757,RIfe853b0_7860,RIee199d8_4750,RIfe85248_7859,RIee39148_5108,
        RIe16b378_2597,RIee38608_5100,RIe167b38_2557,RIe164fa0_2526,RIe1622a0_2494,RIfe85950_7864,RIe15f5a0_2462,RIee36010_5073,RIe15c8a0_2430,RIe156ea0_2366,
        RIe1541a0_2334,RIfe85c20_7866,RIe1514a0_2302,RIee34dc8_5060,RIe14e7a0_2270,RIfc861b0_6548,RIe14baa0_2238,RIe148da0_2206,RIe1460a0_2174,RIee343f0_5053,
        RIfe85518_7861,RIfe857e8_7863,RIfe85680_7862,RIe140c40_2114,RIdf3eb48_2090,RIdf3c820_2065,RIdf3a660_2041,RIfc9d4f0_6812,RIee2f698_4998,RIfc52298_5957,
        RIee2d4d8_4974,RIdf35368_1982,RIdf32ed8_1956,RIdf30e80_1933,RIfe85ab8_7865,RIee2b8b8_4954,RIee29f68_4936,RIee28bb8_4922,RIee27970_4909,RIdf2a0d0_1855,
        RIfe84e10_7856,RIdf262f0_1811,RIfe84ca8_7855,RIee27100_4903,RIee26b60_4899,RIfcd32f8_7425,RIee265c0_4895,RIfc9e300_6822,RIdf1f540_1733,RIee25eb8_4890,
        RIfe84b40_7854,RIdf16b70_1635,RIdf13e70_1603,RIdf11170_1571,RIdf0e470_1539,RIdf0b770_1507,RIdf08a70_1475,RIdf05d70_1443,RIdf03070_1411,RIdefd670_1347,
        RIdefa970_1315,RIdef7c70_1283,RIdef4f70_1251,RIdef2270_1219,RIdeef570_1187,RIdeec870_1155,RIdee9b70_1123,RIfec0348_8307,RIfcb54d8_7085,RIee23cf8_4866,
        RIfc54e30_5988,RIfec0078_8305,RIdee2988_1042,RIfec01e0_8306,RIdede770_995,RIfcd7ee8_7479,RIfcd43d8_7437,RIfc88eb0_6580,RIfc9e5d0_6824,RIded9478_936,
        RIded6fe8_910,RIded50f8_888,RIfeab330_8264,RIded03a0_833,RIdecd6a0_801,RIdeca9a0_769,RIdec7ca0_737,RIdeb41a0_513,RIde95f48_321,RIe16dda8_2627,
        RIe159ba0_2398,RIe1433a0_2142,RIdf37d98_2012,RIdf2c3f8_1880,RIdf1cc78_1704,RIdf00370_1379,RIdee6e70_1091,RIdedbbd8_964,RIde7be90_194,RIe19d238_3165,
        RIe19a538_3133,RIf145658_5249,RIe197838_3101,RIf1446e0_5238,RIe194b38_3069,RIe191e38_3037,RIe18f138_3005,RIe189738_2941,RIe186a38_2909,RIf143600_5226,
        RIe183d38_2877,RIf142c28_5219,RIe181038_2845,RIe17e338_2813,RIe17b638_2781,RIf1420e8_5211,RIf140a68_5195,RIf1401f8_5189,RIfebff10_8304,RIf13faf0_5184,
        RIf13ee48_5175,RIee3e2d8_5166,RIee3d1f8_5154,RIee3c118_5142,RIee3b038_5130,RIee39c88_5116,RIfe838f8_7841,RIf1701c8_5735,RIfc5ab00_6054,RIf16e008_5711,
        RIfcb0e88_7035,RIf16caf0_5696,RIe223590_4692,RIf16bce0_5686,RIe220890_4660,RIf16ac00_5674,RIe21db90_4628,RIe218190_4564,RIe215490_4532,RIf16a228_5667,
        RIe212790_4500,RIf168fe0_5654,RIe20fa90_4468,RIf167d98_5641,RIe20cd90_4436,RIe20a090_4404,RIe207390_4372,RIf1670f0_5632,RIf165ea8_5619,RIe202200_4314,
        RIfe83e98_7845,RIf164f30_5608,RIf1643f0_5600,RIfce8310_7664,RIf161df8_5573,RIf15ff08_5551,RIf15e018_5529,RIfe83d30_7844,RIfe84000_7846,RIf15cb00_5514,
        RIf15b5e8_5499,RIf15a508_5487,RIfc887a8_6575,RIf158d20_5470,RIf157970_5456,RIf156cc8_5447,RIfe84438_7849,RIf156020_5438,RIfc51fc8_5955,RIf154568_5419,
        RIe1f51e0_4166,RIf153050_5404,RIf1519d0_5388,RIf150788_5375,RIfe842d0_7848,RIf14f810_5364,RIf14eb68_5355,RIf14dd58_5345,RIfe84168_7847,RIe1eb2f8_4053,
        RIe1e85f8_4021,RIe1e58f8_3989,RIe1e2bf8_3957,RIe1dfef8_3925,RIe1dd1f8_3893,RIe1da4f8_3861,RIe1d77f8_3829,RIe1d1df8_3765,RIe1cf0f8_3733,RIe1cc3f8_3701,
        RIe1c96f8_3669,RIe1c69f8_3637,RIe1c3cf8_3605,RIe1c0ff8_3573,RIe1be2f8_3541,RIf14c840_5330,RIf14b5f8_5317,RIfe83a60_7842,RIfe849d8_7853,RIfc74168_6343,
        RIf149b40_5298,RIfe83bc8_7843,RIfe84708_7851,RIf148d30_5288,RIf147ae8_5275,RIfe84870_7852,RIe1b0900_3386,RIf146fa8_5267,RIf146300_5258,RIfe845a0_7850,
        RIfe83790_7840,RIe1a8638_3293,RIe1a5938_3261,RIe1a2c38_3229,RIe19ff38_3197,RIe18c438_2973,RIe178938_2749,RIe226290_4724,RIe21ae90_4596,RIe204690_4340,
        RIe1fe6f0_4272,RIe1f7aa8_4195,RIe1f05f0_4112,RIe1d4af8_3797,RIe1bb5f8_3509,RIe1ae470_3360,RIe170aa8_2659,RIdec4e38_704,RIdec2138_672,RIee1fc48_4820,
        RIdebf438_640,RIfc49490_5856,RIdebc738_608,RIdeb9a38_576,RIdeb6d38_544,RIfc48ef0_5852,RIdeb1338_480,RIfcd9b08_7499,RIdeae638_448,RIfc8b610_6608,
        RIdea9700_416,RIdea2e00_384,RIde9c500_352,RIee1c9a8_4784,RIee1b8c8_4772,RIfc80918_6485,RIfcdad50_7512,RIfe86e68_7879,RIde8cee8_277,RIfe86d00_7878,
        RIfec0d20_8314,RIde81098_219,RIfc8b8e0_6610,RIfcd2d58_7421,RIfce4530_7620,RIfc8ba48_6611,RIe16b210_2596,RIe1698c0_2578,RIe1679d0_2556,RIe164e38_2525,
        RIe162138_2493,RIee370f0_5085,RIe15f438_2461,RIfc999e0_6770,RIe15c738_2429,RIe156d38_2365,RIe154038_2333,RIfc3f260_5744,RIe151338_2301,RIfc48518_5845,
        RIe14e638_2269,RIfc99e18_6773,RIe14b938_2237,RIe148c38_2205,RIe145f38_2173,RIee34288_5052,RIee33040_5039,RIee31f60_5027,RIfcd99a0_7498,RIfe86b98_7877,
        RIdf3e9e0_2089,RIfe86a30_7876,RIdf3a4f8_2040,RIfcc3470_7244,RIee2f530_4997,RIfc7fdd8_6477,RIee2d370_4973,RIdf35200_1981,RIfec0ff0_8316,RIdf30d18_1932,
        RIfec0e88_8315,RIfcd2a88_7419,RIfc8c858_6621,RIfc47ca8_5839,RIfcd6430_7460,RIdf29f68_1854,RIdf27da8_1830,RIdf26188_1810,RIdf24568_1790,RIfc8cb28_6623,
        RIfcdb188_7515,RIdf22948_1770,RIfc475a0_5834,RIdf21430_1755,RIdf1f3d8_1732,RIfec0bb8_8313,RIfe868c8_7875,RIdf16a08_1634,RIdf13d08_1602,RIdf11008_1570,
        RIdf0e308_1538,RIdf0b608_1506,RIdf08908_1474,RIdf05c08_1442,RIdf02f08_1410,RIdefd508_1346,RIdefa808_1314,RIdef7b08_1282,RIdef4e08_1250,RIdef2108_1218,
        RIdeef408_1186,RIdeec708_1154,RIdee9a08_1122,RIee254e0_4883,RIee246d0_4873,RIee23b90_4865,RIee231b8_4858,RIfe86fd0_7880,RIdee2820_1041,RIdee0930_1019,
        RIdede608_994,RIfc55da8_5999,RIfc98a68_6759,RIfcc3038_7241,RIfc464c0_5822,RIded9310_935,RIded6e80_909,RIded4f90_887,RIded2b00_861,RIded0238_832,
        RIdecd538_800,RIdeca838_768,RIdec7b38_736,RIdeb4038_512,RIde95c00_320,RIe16dc40_2626,RIe159a38_2397,RIe143238_2141,RIdf37c30_2011,RIdf2c290_1879,
        RIdf1cb10_1703,RIdf00208_1378,RIdee6d08_1090,RIdedba70_963,RIde7bb48_193,RIe19d0d0_3164,RIe19a3d0_3132,RIf1454f0_5248,RIe1976d0_3100,RIf144578_5237,
        RIe1949d0_3068,RIe191cd0_3036,RIe18efd0_3004,RIe1895d0_2940,RIe1868d0_2908,RIf143498_5225,RIe183bd0_2876,RIfc51758_5949,RIe180ed0_2844,RIe17e1d0_2812,
        RIe17b4d0_2780,RIfc9b060_6786,RIfc9ee40_6830,RIe176e80_2730,RIe175800_2714,RIfcb70f8_7105,RIfce0cf0_7580,RIfcc4280_7254,RIfcba7d0_7144,RIee3bfb0_5141,
        RIee3aed0_5129,RIee39b20_5115,RIe173370_2688,RIf170060_5734,RIf16f3b8_5725,RIf16dea0_5710,RIf16d4c8_5703,RIf16c988_5695,RIe223428_4691,RIf16bb78_5685,
        RIe220728_4659,RIf16aa98_5673,RIe21da28_4627,RIe218028_4563,RIe215328_4531,RIf16a0c0_5666,RIe212628_4499,RIf168e78_5653,RIe20f928_4467,RIf167c30_5640,
        RIe20cc28_4435,RIe209f28_4403,RIe207228_4371,RIf166f88_5631,RIf165d40_5618,RIfec0618_8309,RIfe86760_7874,RIfc52b08_5963,RIf164288_5599,RIf163310_5588,
        RIf161c90_5572,RIf15fda0_5550,RIf15deb0_5528,RIfe865f8_7873,RIfe85d88_7867,RIf15c998_5513,RIf15b480_5498,RIf15a3a0_5486,RIf159b30_5480,RIfc83348_6515,
        RIfc4ade0_5874,RIfc89720_6586,RIe1f9f38_4221,RIfc4ac78_5873,RIfc9f110_6832,RIfc4ab10_5872,RIe1f5078_4165,RIf152ee8_5403,RIfc899f0_6588,RIf150620_5374,
        RIe1f2eb8_4141,RIf14f6a8_5363,RIf14ea00_5354,RIf14dbf0_5344,RIe1edbc0_4082,RIe1eb190_4052,RIe1e8490_4020,RIe1e5790_3988,RIe1e2a90_3956,RIe1dfd90_3924,
        RIe1dd090_3892,RIe1da390_3860,RIe1d7690_3828,RIe1d1c90_3764,RIe1cef90_3732,RIe1cc290_3700,RIe1c9590_3668,RIe1c6890_3636,RIe1c3b90_3604,RIe1c0e90_3572,
        RIe1be190_3540,RIf14c6d8_5329,RIf14b490_5316,RIfe85ef0_7868,RIfe86490_7872,RIf14a248_5303,RIfc819f8_6497,RIfec0a50_8312,RIfe861c0_7870,RIf148bc8_5287,
        RIf147980_5274,RIfe86328_7871,RIfec0780_8310,RIfcbb478_7153,RIf146198_5257,RIfe86058_7869,RIfec08e8_8311,RIe1a84d0_3292,RIe1a57d0_3260,RIe1a2ad0_3228,
        RIe19fdd0_3196,RIe18c2d0_2972,RIe1787d0_2748,RIe226128_4723,RIe21ad28_4595,RIe204528_4339,RIe1fe588_4271,RIe1f7940_4194,RIe1f0488_4111,RIe1d4990_3796,
        RIe1bb490_3508,RIe1ae308_3359,RIe170940_2658,RIdec53d8_708,RIdec26d8_676,RIee20080_4823,RIdebf9d8_644,RIee1f3d8_4814,RIdebccd8_612,RIdeb9fd8_580,
        RIdeb72d8_548,RIee1ee38_4810,RIdeb18d8_484,RIee1e898_4806,RIdeaebd8_452,RIee1da88_4796,RIdeaa420_420,RIdea3b20_388,RIde9d220_356,RIee1cde0_4787,
        RIee1bd00_4775,RIee1b490_4769,RIfcd8a28_7487,RIde91088_297,RIde8d8c0_280,RIfe7dac0_7774,RIfe7d958_7773,RIee1a518_4758,RIee19e10_4753,RIee19b40_4751,
        RIfc768c8_6371,RIfcd05f8_7393,RIfe7dd90_7776,RIee38770_5101,RIfe7dc28_7775,RIe1653d8_2529,RIe1626d8_2497,RIee373c0_5087,RIe15f9d8_2465,RIee362e0_5075,
        RIe15ccd8_2433,RIe1572d8_2369,RIe1545d8_2337,RIfe7def8_7777,RIe1518d8_2305,RIfebdeb8_8281,RIe14ebd8_2273,RIfc649e8_6167,RIe14bed8_2241,RIe1491d8_2209,
        RIe1464d8_2177,RIfe7d7f0_7772,RIfe7d688_7771,RIee32230_5029,RIfceb9e8_7703,RIfebdd50_8280,RIfe7d520_7770,RIfebdbe8_8279,RIfe7d3b8_7769,RIfc734c0_6334,
        RIee2f968_5000,RIfccfab8_7385,RIee2d7a8_4976,RIdf357a0_1985,RIdf33310_1959,RIdf312b8_1936,RIdf2f0f8_1912,RIee2bcf0_4957,RIee2a238_4938,RIee28e88_4924,
        RIee27c40_4911,RIfe7ce18_7765,RIfe7ccb0_7764,RIfe7cf80_7766,RIfe7cb48_7763,RIee27268_4904,RIee26e30_4901,RIee26890_4897,RIfcaa0d8_6957,RIee262f0_4893,
        RIfe7d250_7768,RIee26020_4891,RIfe7d0e8_7767,RIdf16fa8_1638,RIdf142a8_1606,RIdf115a8_1574,RIdf0e8a8_1542,RIdf0bba8_1510,RIdf08ea8_1478,RIdf061a8_1446,
        RIdf034a8_1414,RIdefdaa8_1350,RIdefada8_1318,RIdef80a8_1286,RIdef53a8_1254,RIdef26a8_1222,RIdeef9a8_1190,RIdeecca8_1158,RIdee9fa8_1126,RIee25648_4884,
        RIee249a0_4875,RIfebe020_8282,RIee23488_4860,RIfebe2f0_8284,RIfebe188_8283,RIfe7e1c8_7779,RIfe7e060_7778,RIfcbf7f8_7201,RIfc7aae0_6418,RIfc787b8_6393,
        RIfc618b0_6132,RIded98b0_939,RIded72b8_912,RIded5530_891,RIded2dd0_863,RIded07d8_836,RIdecdad8_804,RIdecadd8_772,RIdec80d8_740,RIdeb45d8_516,
        RIde96920_324,RIe16e1e0_2630,RIe159fd8_2401,RIe1437d8_2145,RIdf381d0_2015,RIdf2c830_1883,RIdf1d0b0_1707,RIdf007a8_1382,RIdee72a8_1094,RIdedc010_967,
        RIde7c868_197,RIe19d670_3168,RIe19a970_3136,RIfe7b630_7748,RIe197c70_3104,RIfe7b4c8_7747,RIe194f70_3072,RIe192270_3040,RIe18f570_3008,RIe189b70_2944,
        RIe186e70_2912,RIfe7b360_7746,RIe184170_2880,RIfe7b1f8_7745,RIe181470_2848,RIe17e770_2816,RIe17ba70_2784,RIf1423b8_5213,RIf140ea0_5198,RIf140360_5190,
        RIfe7b798_7749,RIf13fc58_5185,RIf13f280_5178,RIfc79460_6402,RIee3d4c8_5156,RIfe7b090_7744,RIfe7af28_7743,RIee39df0_5117,RIe1737a8_2691,RIfe7adc0_7742,
        RIfe7ac58_7741,RIf16e440_5714,RIfcb20d0_7048,RIfe7bd38_7753,RIe2239c8_4695,RIf16be48_5687,RIe220cc8_4663,RIf16aed0_5676,RIe21dfc8_4631,RIe2185c8_4567,
        RIe2158c8_4535,RIfebd7b0_8276,RIe212bc8_4503,RIfebd648_8275,RIe20fec8_4471,RIfe7b900_7750,RIe20d1c8_4439,RIe20a4c8_4407,RIe2077c8_4375,RIf167258_5633,
        RIf166178_5621,RIe2024d0_4316,RIfe7bbd0_7752,RIf165368_5611,RIf1646c0_5602,RIfcd0a30_7396,RIf1620c8_5575,RIf1601d8_5553,RIf15e2e8_5531,RIfe7ba68_7751,
        RIfe7bea0_7754,RIf15cdd0_5516,RIf15b8b8_5501,RIf15a7d8_5489,RIfca4840_6894,RIf158ff0_5472,RIf157c40_5458,RIf156f98_5449,RIfe7c170_7756,RIf156458_5441,
        RIf155918_5433,RIf1549a0_5422,RIe1f54b0_4168,RIfe7c008_7755,RIf151b38_5389,RIf150bc0_5378,RIe1f32f0_4144,RIf14fae0_5366,RIf14ee38_5357,RIf14e028_5347,
        RIe1edff8_4085,RIe1eb730_4056,RIe1e8a30_4024,RIe1e5d30_3992,RIe1e3030_3960,RIe1e0330_3928,RIe1dd630_3896,RIe1da930_3864,RIe1d7c30_3832,RIe1d2230_3768,
        RIe1cf530_3736,RIe1cc830_3704,RIe1c9b30_3672,RIe1c6e30_3640,RIe1c4130_3608,RIe1c1430_3576,RIe1be730_3544,RIf14cb10_5332,RIf14b8c8_5319,RIfebda80_8278,
        RIfe7c878_7761,RIf14a680_5306,RIfe7c2d8_7757,RIfe7c9e0_7762,RIfe7c440_7758,RIf149000_5290,RIf147db8_5277,RIe1b2688_3407,RIfebd918_8277,RIfe7c5a8_7759,
        RIf146738_5261,RIfe7c710_7760,RIe1aad98_3321,RIe1a8a70_3296,RIe1a5d70_3264,RIe1a3070_3232,RIe1a0370_3200,RIe18c870_2976,RIe178d70_2752,RIe2266c8_4727,
        RIe21b2c8_4599,RIe204ac8_4343,RIe1feb28_4275,RIe1f7ee0_4198,RIe1f0a28_4115,RIe1d4f30_3800,RIe1bba30_3512,RIe1ae8a8_3363,RIe170ee0_2662,RIdec5270_707,
        RIdec2570_675,RIee1ff18_4822,RIdebf870_643,RIfe7f848_7795,RIdebcb70_611,RIdeb9e70_579,RIdeb7170_547,RIfe7fc80_7798,RIdeb1770_483,RIfca5d58_6909,
        RIdeaea70_451,RIfcaf808_7019,RIdeaa0d8_419,RIdea37d8_387,RIde9ced8_355,RIfcdc3d0_7528,RIfcce438_7369,RIfcb0a50_7032,RIfc75680_6358,RIde90d40_296,
        RIfe7f9b0_7796,RIde89720_260,RIde85580_240,RIde81728_221,RIfc52f40_5966,RIfc82100_6502,RIfca7108_6923,RIfe7fb18_7797,RIe16b648_2599,RIe169a28_2579,
        RIe167ca0_2558,RIe165270_2528,RIe162570_2496,RIee37258_5086,RIe15f870_2464,RIee36178_5074,RIe15cb70_2432,RIe157170_2368,RIe154470_2336,RIfc86fc0_6558,
        RIe151770_2304,RIfc4eff8_5921,RIe14ea70_2272,RIfce1290_7584,RIe14bd70_2240,RIe149070_2208,RIe146370_2176,RIee34558_5054,RIee331a8_5040,RIee320c8_5028,
        RIee31150_5017,RIfe800b8_7801,RIfe7ff50_7800,RIdf3caf0_2067,RIfe7fde8_7799,RIfcc8330_7300,RIee2f800_4999,RIfca0d30_6852,RIee2d640_4975,RIdf35638_1984,
        RIdf331a8_1958,RIdf31150_1935,RIdf2ef90_1911,RIee2bb88_4956,RIee2a0d0_4937,RIee28d20_4923,RIfe7f578_7793,RIdf2a238_1856,RIdf27f10_1831,RIfe7f6e0_7794,
        RIdf246d0_1791,RIfcce9d8_7373,RIfc63638_6153,RIdf22c18_1772,RIfc62990_6144,RIdf21700_1757,RIdf1f810_1735,RIfeaa958_8257,RIdf19168_1662,RIdf16e40_1637,
        RIdf14140_1605,RIdf11440_1573,RIdf0e740_1541,RIdf0ba40_1509,RIdf08d40_1477,RIdf06040_1445,RIdf03340_1413,RIdefd940_1349,RIdefac40_1317,RIdef7f40_1285,
        RIdef5240_1253,RIdef2540_1221,RIdeef840_1189,RIdeecb40_1157,RIdee9e40_1125,RIfcb7800_7110,RIee24838_4874,RIfc4cb68_5895,RIee23320_4859,RIfe80388_7803,
        RIdee2c58_1044,RIfe80220_7802,RIdedea40_997,RIfc98900_6758,RIee223a8_4848,RIfcc8600_7302,RIee212c8_4836,RIded9748_938,RIfe804f0_7804,RIded53c8_890,
        RIded2c68_862,RIded0670_835,RIdecd970_803,RIdecac70_771,RIdec7f70_739,RIdeb4470_515,RIde965d8_323,RIe16e078_2629,RIe159e70_2400,RIe143670_2144,
        RIdf38068_2014,RIdf2c6c8_1882,RIdf1cf48_1706,RIdf00640_1381,RIdee7140_1093,RIdedbea8_966,RIde7c520_196,RIe19d508_3167,RIe19a808_3135,RIfe7ee70_7788,
        RIe197b08_3103,RIfe7efd8_7789,RIe194e08_3071,RIe192108_3039,RIe18f408_3007,RIe189a08_2943,RIe186d08_2911,RIf143768_5227,RIe184008_2879,RIfc4bbf0_5884,
        RIe181308_2847,RIe17e608_2815,RIe17b908_2783,RIfe7f410_7792,RIf140d38_5197,RIe176fe8_2731,RIe175ad0_2716,RIfe7f2a8_7791,RIf13f118_5177,RIee3e440_5167,
        RIee3d360_5155,RIee3c280_5143,RIee3b1a0_5131,RIfe7f140_7790,RIe173640_2690,RIf170330_5736,RIf16f520_5726,RIf16e2d8_5713,RIf16d630_5704,RIfe7ea38_7785,
        RIe223860_4694,RIfc9c410_6800,RIe220b60_4662,RIfcb8340_7118,RIe21de60_4630,RIe218460_4566,RIe215760_4534,RIfc9cc80_6806,RIe212a60_4502,RIfc4ddb0_5908,
        RIe20fd60_4470,RIfc873f8_6561,RIe20d060_4438,RIe20a360_4406,RIe207660_4374,RIfc86750_6552,RIfc4e4b8_5913,RIe202368_4315,RIe200a18_4297,RIf165200_5610,
        RIf164558_5601,RIf163478_5589,RIf161f60_5574,RIf160070_5552,RIf15e180_5530,RIe1fcc38_4253,RIe1fb9f0_4240,RIf15cc68_5515,RIf15b750_5500,RIf15a670_5488,
        RIf159c98_5481,RIf158e88_5471,RIf157ad8_5457,RIf156e30_5448,RIfe7e768_7783,RIf1562f0_5440,RIf1557b0_5432,RIf154838_5421,RIfe7e8d0_7784,RIf1531b8_5405,
        RIfc52400_5958,RIf150a58_5377,RIe1f3188_4143,RIf14f978_5365,RIf14ecd0_5356,RIf14dec0_5346,RIe1ede90_4084,RIe1eb5c8_4055,RIe1e88c8_4023,RIe1e5bc8_3991,
        RIe1e2ec8_3959,RIe1e01c8_3927,RIe1dd4c8_3895,RIe1da7c8_3863,RIe1d7ac8_3831,RIe1d20c8_3767,RIe1cf3c8_3735,RIe1cc6c8_3703,RIe1c99c8_3671,RIe1c6cc8_3639,
        RIe1c3fc8_3607,RIe1c12c8_3575,RIe1be5c8_3543,RIf14c9a8_5331,RIf14b760_5318,RIfe7ed08_7787,RIfe7e600_7782,RIf14a518_5305,RIfca1f78_6865,RIfe7eba0_7786,
        RIfe7e498_7781,RIf148e98_5289,RIf147c50_5276,RIfe7e330_7780,RIe1b0a68_3387,RIf147278_5269,RIf1465d0_5260,RIe1ac418_3337,RIe1aac30_3320,RIe1a8908_3295,
        RIe1a5c08_3263,RIe1a2f08_3231,RIe1a0208_3199,RIe18c708_2975,RIe178c08_2751,RIe226560_4726,RIe21b160_4598,RIe204960_4342,RIe1fe9c0_4274,RIe1f7d78_4197,
        RIe1f08c0_4114,RIe1d4dc8_3799,RIe1bb8c8_3511,RIe1ae740_3362,RIe170d78_2661,RIdec56a8_710,RIdec29a8_678,RIfc54020_5978,RIdebfca8_646,RIee1f540_4815,
        RIdebcfa8_614,RIdeba2a8_582,RIdeb75a8_550,RIfc4fe08_5931,RIdeb1ba8_486,RIfc6b630_6244,RIdeaeea8_454,RIfc6a118_6229,RIdeaaab0_422,RIdea41b0_390,
        RIde9d8b0_358,RIfc69ce0_6226,RIee1be68_4776,RIfc653c0_6174,RIee1ac20_4763,RIde91718_299,RIde8df50_282,RIde89db0_262,RIde85c10_242,RIde81db8_223,
        RIfca76a8_6927,RIfcca4f0_7324,RIfc4ce38_5897,RIfc6b360_6242,RIe16b918_2601,RIe169cf8_2581,RIe167f70_2560,RIe1656a8_2531,RIe1629a8_2499,RIee37690_5089,
        RIe15fca8_2467,RIfce93f0_7676,RIe15cfa8_2435,RIe1575a8_2371,RIe1548a8_2339,RIee35908_5068,RIe151ba8_2307,RIee34f30_5061,RIe14eea8_2275,RIfce32e8_7607,
        RIe14c1a8_2243,RIe1494a8_2211,RIe1467a8_2179,RIfcde2c0_7550,RIfc687c8_6211,RIfca9160_6946,RIfcb1590_7040,RIe141078_2117,RIdf3ef80_2093,RIdf3cdc0_2069,
        RIfebeb60_8290,RIfc64448_6163,RIee2fad0_5001,RIfca7978_6929,RIfc676e8_6199,RIdf35a70_1987,RIdf335e0_1961,RIdf31420_1937,RIdf2f3c8_1914,RIfccef78_7377,
        RIfca6fa0_6922,RIfc62558_6141,RIfc61fb8_6137,RIfe81b70_7820,RIdf281e0_1833,RIfe81cd8_7821,RIdf249a0_1793,RIfc44300_5798,RIfcafc40_7022,RIdf22ee8_1774,
        RIfcaac18_6965,RIdf219d0_1759,RIdf1fae0_1737,RIdf1b1c0_1685,RIdf19438_1664,RIdf17278_1640,RIdf14578_1608,RIdf11878_1576,RIdf0eb78_1544,RIdf0be78_1512,
        RIdf09178_1480,RIdf06478_1448,RIdf03778_1416,RIdefdd78_1352,RIdefb078_1320,RIdef8378_1288,RIdef5678_1256,RIdef2978_1224,RIdeefc78_1192,RIdeecf78_1160,
        RIdeea278_1128,RIfc611a8_6127,RIfc61a18_6133,RIfca65c8_6915,RIfca6b68_6919,RIdee4b48_1066,RIdee2dc0_1045,RIdee0c00_1021,RIdedeba8_998,RIfc626c0_6142,
        RIfc738f8_6337,RIfcb31b0_7060,RIee21430_4837,RIded9a18_940,RIded7588_914,RIded5698_892,RIded30a0_865,RIded0aa8_838,RIdecdda8_806,RIdecb0a8_774,
        RIdec83a8_742,RIdeb48a8_518,RIde96fb0_326,RIe16e4b0_2632,RIe15a2a8_2403,RIe143aa8_2147,RIdf384a0_2017,RIdf2cb00_1885,RIdf1d380_1709,RIdf00a78_1384,
        RIdee7578_1096,RIdedc2e0_969,RIde7cef8_199,RIe19d940_3170,RIe19ac40_3138,RIfc64880_6166,RIe197f40_3106,RIf144848_5239,RIe195240_3074,RIe192540_3042,
        RIe18f840_3010,RIe189e40_2946,RIe187140_2914,RIf143a38_5229,RIe184440_2882,RIfc6f140_6286,RIe181740_2850,RIe17ea40_2818,RIe17bd40_2786,RIfc64f88_6171,
        RIf141008_5199,RIe177150_2732,RIfe81738_7817,RIfccabf8_7329,RIf13f3e8_5179,RIfca81e8_6935,RIee3d630_5157,RIfc66068_6183,RIfc6ed08_6283,RIfcdde88_7547,
        RIe173a78_2693,RIfc66338_6185,RIfc6eba0_6282,RIfc664a0_6186,RIfcacdd8_6989,RIfe81468_7815,RIe223c98_4697,RIfc66d10_6192,RIe220f98_4665,RIf16b038_5677,
        RIe21e298_4633,RIe218898_4569,RIe215b98_4537,RIfc3fc38_5751,RIe212e98_4505,RIfc67850_6200,RIe210198_4473,RIf167f00_5642,RIe20d498_4441,RIe20a798_4409,
        RIe207a98_4377,RIfcacb08_6987,RIfcac9a0_6986,RIfea8900_8234,RIfe818a0_7818,RIfca8a58_6941,RIfccad60_7330,RIfcac838_6985,RIfc67418_6197,RIf160340_5554,
        RIf15e450_5532,RIfe81a08_7819,RIfe81300_7814,RIfc6dac0_6270,RIf15ba20_5502,RIfc6d958_6269,RIfc6d7f0_6268,RIfc587d8_6029,RIfc6cf80_6262,RIfc6d3b8_6265,
        RIfe815d0_7816,RIfc6d520_6266,RIfcabe60_6978,RIfc6d0e8_6263,RIe1f5780_4170,RIfc6c5a8_6255,RIfc68d68_6215,RIfc68c00_6214,RIe1f3458_4145,RIfc68a98_6213,
        RIfccb8a0_7338,RIfca9b38_6953,RIe1ee160_4086,RIe1eba00_4058,RIe1e8d00_4026,RIe1e6000_3994,RIe1e3300_3962,RIe1e0600_3930,RIe1dd900_3898,RIe1dac00_3866,
        RIe1d7f00_3834,RIe1d2500_3770,RIe1cf800_3738,RIe1ccb00_3706,RIe1c9e00_3674,RIe1c7100_3642,RIe1c4400_3610,RIe1c1700_3578,RIe1bea00_3546,RIfc6bbd0_6248,
        RIfcdd348_7539,RIe1b9438_3485,RIe1b73e0_3462,RIfcab5f0_6972,RIfccbb70_7340,RIe1b5220_3438,RIe1b3e70_3424,RIfc6c9e0_6258,RIfcab488_6971,RIfea7dc0_8226,
        RIe1b0bd0_3388,RIfc6ce18_6261,RIfcabfc8_6979,RIe1ac580_3338,RIe1aaf00_3322,RIe1a8d40_3298,RIe1a6040_3266,RIe1a3340_3234,RIe1a0640_3202,RIe18cb40_2978,
        RIe179040_2754,RIe226998_4729,RIe21b598_4601,RIe204d98_4345,RIe1fedf8_4277,RIe1f81b0_4200,RIe1f0cf8_4117,RIe1d5200_3802,RIe1bbd00_3514,RIe1aeb78_3365,
        RIe1711b0_2664,RIdec5540_709,RIdec2840_677,RIfcc4dc0_7262,RIdebfb40_645,RIfc9d7c0_6814,RIdebce40_613,RIdeba140_581,RIdeb7440_549,RIfc4d978_5905,
        RIdeb1a40_485,RIfc9dbf8_6817,RIdeaed40_453,RIfcb8610_7120,RIdeaa768_421,RIdea3e68_389,RIde9d568_357,RIfc50678_5937,RIfc507e0_5938,RIfc9dec8_6819,
        RIfc853a0_6538,RIde913d0_298,RIde8dc08_281,RIde89a68_261,RIde858c8_241,RIde81a70_222,RIfc84860_6530,RIfc50948_5939,RIfc84c98_6533,RIfcb7da0_7114,
        RIe16b7b0_2600,RIe169b90_2580,RIe167e08_2559,RIe165540_2530,RIe162840_2498,RIee37528_5088,RIe15fb40_2466,RIfcb5be0_7090,RIe15ce40_2434,RIe157440_2370,
        RIe154740_2338,RIfcd35c8_7427,RIe151a40_2306,RIfc53a80_5974,RIe14ed40_2274,RIfcc6170_7276,RIe14c040_2242,RIe149340_2210,RIe146640_2178,RIfc7f130_6468,
        RIee33310_5041,RIfcb4f38_7081,RIfc47f78_5841,RIe140f10_2116,RIdf3ee18_2092,RIdf3cc58_2068,RIdf3a7c8_2042,RIfc7fc70_6476,RIfcd27b8_7417,RIfca1000_6854,
        RIfcc6b48_7283,RIdf35908_1986,RIdf33478_1960,RIfebe9f8_8289,RIdf2f260_1913,RIfcb7968_7111,RIee2a3a0_4939,RIfc51050_5944,RIfcd3fa0_7434,RIdf2a3a0_1857,
        RIdf28078_1832,RIfe81198_7813,RIdf24838_1792,RIfc84428_6527,RIfce7ed8_7661,RIdf22d80_1773,RIfc515f0_5948,RIdf21868_1758,RIdf1f978_1736,RIdf1b058_1684,
        RIdf192d0_1663,RIdf17110_1639,RIdf14410_1607,RIdf11710_1575,RIdf0ea10_1543,RIdf0bd10_1511,RIdf09010_1479,RIdf06310_1447,RIdf03610_1415,RIdefdc10_1351,
        RIdefaf10_1319,RIdef8210_1287,RIdef5510_1255,RIdef2810_1223,RIdeefb10_1191,RIdeece10_1159,RIdeea110_1127,RIfc7e1b8_6457,RIfca19d8_6861,RIfc7dab0_6452,
        RIfc7e488_6459,RIdee49e0_1065,RIfe80d60_7810,RIfeabba0_8270,RIfe80bf8_7809,RIfcb3750_7064,RIfce9f30_7684,RIfc7e5f0_6460,RIfc56a50_6008,RIfe81030_7812,
        RIded7420_913,RIfe80ec8_7811,RIded2f38_864,RIded0940_837,RIdecdc40_805,RIdecaf40_773,RIdec8240_741,RIdeb4740_517,RIde96c68_325,RIe16e348_2631,
        RIe15a140_2402,RIe143940_2146,RIdf38338_2016,RIdf2c998_1884,RIdf1d218_1708,RIdf00910_1383,RIdee7410_1095,RIdedc178_968,RIde7cbb0_198,RIe19d7d8_3169,
        RIe19aad8_3137,RIfcc2d68_7239,RIe197dd8_3105,RIfc5c5b8_6073,RIe1950d8_3073,RIe1923d8_3041,RIe18f6d8_3009,RIe189cd8_2945,RIe186fd8_2913,RIf1438d0_5228,
        RIe1842d8_2881,RIfc5b370_6060,RIe1815d8_2849,RIe17e8d8_2817,RIe17bbd8_2785,RIfcbb748_7155,RIfc59480_6038,RIfcbbce8_7159,RIe175c38_2717,RIfcdb890_7520,
        RIfc59b88_6043,RIfc8ada0_6602,RIfcb5eb0_7092,RIfc57c98_6021,RIfc57158_6013,RIfc58aa8_6031,RIe173910_2692,RIfcc62d8_7277,RIfc8a968_6599,RIfc57428_6015,
        RIfc56d20_6010,RIfc408e0_5760,RIe223b30_4696,RIfc82970_6508,RIe220e30_4664,RIfcecc30_7716,RIe21e130_4632,RIe218730_4568,RIe215a30_4536,RIfc3fad0_5750,
        RIe212d30_4504,RIf169148_5655,RIe210030_4472,RIfc545c0_5982,RIe20d330_4440,RIe20a630_4408,RIe207930_4376,RIfc88d48_6579,RIfc4bec0_5886,RIe202638_4317,
        RIe200b80_4298,RIfc88910_6576,RIfc4c190_5888,RIfc4c2f8_5889,RIfcba398_7141,RIfcd4270_7436,RIfcba0c8_7139,RIe1fcda0_4254,RIe1fbb58_4241,RIfc53d50_5976,
        RIfc9b768_6791,RIfc537b0_5972,RIfc4c5c8_5891,RIfc9e468_6823,RIf157da8_5459,RIfcb9f60_7138,RIe1fa208_4223,RIfc849c8_6531,RIfc529a0_5962,RIfc9f6b0_6836,
        RIe1f5618_4169,RIf153320_5406,RIfcc4988_7259,RIf150d28_5379,RIfebe458_8285,RIfc87f38_6569,RIfcb7f08_7115,RIf14e190_5348,RIfe80658_7805,RIe1eb898_4057,
        RIe1e8b98_4025,RIe1e5e98_3993,RIe1e3198_3961,RIe1e0498_3929,RIe1dd798_3897,RIe1daa98_3865,RIe1d7d98_3833,RIe1d2398_3769,RIe1cf698_3737,RIe1cc998_3705,
        RIe1c9c98_3673,RIe1c6f98_3641,RIe1c4298_3609,RIe1c1598_3577,RIe1be898_3545,RIf14cc78_5333,RIf14ba30_5320,RIe1b92d0_3484,RIe1b7278_3461,RIf14a7e8_5307,
        RIf149ca8_5299,RIfebe5c0_8286,RIfe807c0_7806,RIfc50510_5936,RIfce4f08_7627,RIfe80a90_7808,RIfebe890_8288,RIfc9cde8_6807,RIfc87560_6562,RIfe80928_7807,
        RIfebe728_8287,RIe1a8bd8_3297,RIe1a5ed8_3265,RIe1a31d8_3233,RIe1a04d8_3201,RIe18c9d8_2977,RIe178ed8_2753,RIe226830_4728,RIe21b430_4600,RIe204c30_4344,
        RIe1fec90_4276,RIe1f8048_4199,RIe1f0b90_4116,RIe1d5098_3801,RIe1bbb98_3513,RIe1aea10_3364,RIe171048_2663,RIdec5978_712,RIdec2c78_680,RIfc8aad0_6600,
        RIdebff78_648,RIfc8ac38_6601,RIdebd278_616,RIdeba578_584,RIdeb7878_552,RIfc40e80_5764,RIdeb1e78_488,RIfcdaeb8_7513,RIdeaf178_456,RIee1dbf0_4797,
        RIdeab140_424,RIdea4840_392,RIde9df40_360,RIfc8b070_6604,RIfcc38a8_7247,RIfc807b0_6484,RIfcbb8b0_7156,RIde91a60_300,RIde8e298_283,RIde8a440_264,
        RIde862a0_244,RIde82100_224,RIfcbbb80_7158,RIfc8c150_6616,RIfcbbfb8_7161,RIfc54458_5981,RIe16bbe8_2603,RIfc8c2b8_6617,RIe168240_2562,RIe165978_2533,
        RIe162c78_2501,RIee37960_5091,RIe15ff78_2469,RIfcd6b38_7465,RIe15d278_2437,RIe157878_2373,RIe154b78_2341,RIfc8e5e0_6642,RIe151e78_2309,RIfcb4290_7072,
        RIe14f178_2277,RIfc56ff0_6012,RIe14c478_2245,RIe149778_2213,RIe146a78_2181,RIee346c0_5055,RIee335e0_5043,RIee32398_5030,RIee31420_5019,RIe141348_2119,
        RIe13f020_2094,RIfec16f8_8321,RIdf3a930_2043,RIfce3e28_7615,RIfc56780_6006,RIfcb4128_7071,RIfce2eb0_7604,RIdf35d40_1989,RIfe88218_7893,RIdf316f0_1939,
        RIdf2f698_1916,RIfc7f9a0_6474,RIfce4260_7618,RIfcd62c8_7459,RIfce9990_7680,RIdf2a670_1859,RIdf284b0_1835,RIdf26728_1814,RIdf24c70_1795,RIfc7ecf8_6465,
        RIfcc31a0_7242,RIfc99008_6763,RIfc46e98_5829,RIfce2a78_7601,RIdf1fdb0_1739,RIfcc6e18_7285,RIdf19708_1666,RIdf17548_1642,RIdf14848_1610,RIdf11b48_1578,
        RIdf0ee48_1546,RIdf0c148_1514,RIdf09448_1482,RIdf06748_1450,RIdf03a48_1418,RIdefe048_1354,RIdefb348_1322,RIdef8648_1290,RIdef5948_1258,RIdef2c48_1226,
        RIdeeff48_1194,RIdeed248_1162,RIdeea548_1130,RIfcd9130_7492,RIfc7cb38_6441,RIfc97af0_6748,RIfcb3e58_7069,RIdee4e18_1068,RIdee3090_1047,RIdee0ed0_1023,
        RIfe88380_7894,RIfc97dc0_6750,RIfcc2930_7236,RIfcd9298_7493,RIfc7c868_6439,RIded9ce8_942,RIded76f0_915,RIded5968_894,RIded3370_867,RIded0d78_840,
        RIdece078_808,RIdecb378_776,RIdec8678_744,RIdeb4b78_520,RIde97640_328,RIe16e780_2634,RIe15a578_2405,RIe143d78_2149,RIdf38770_2019,RIdf2cdd0_1887,
        RIdf1d650_1711,RIdf00d48_1386,RIdee7848_1098,RIdedc5b0_971,RIde7d588_201,RIe19dc10_3172,RIe19af10_3140,RIfec1590_8320,RIe198210_3108,RIfec1428_8319,
        RIe195510_3076,RIe192810_3044,RIe18fb10_3012,RIe18a110_2948,RIe187410_2916,RIfec12c0_8318,RIe184710_2884,RIfc88370_6572,RIe181a10_2852,RIe17ed10_2820,
        RIe17c010_2788,RIfc6ccb0_6260,RIfc5f858_6109,RIfca88f0_6940,RIe175f08_2719,RIfc81020_6490,RIfcc6008_7275,RIfc4ea58_5917,RIfc42140_5774,RIfca3b98_6885,
        RIfc5ac68_6055,RIfc984c8_6755,RIe173d48_2695,RIfc9b330_6788,RIf16f688_5727,RIfc42410_5776,RIfc5f588_6107,RIfe880b0_7892,RIe223f68_4699,RIf16bfb0_5688,
        RIe221268_4667,RIfc86cf0_6556,RIe21e568_4635,RIe218b68_4571,RIe215e68_4539,RIfe87de0_7890,RIe213168_4507,RIf1692b0_5656,RIe210468_4475,RIfcdf670_7564,
        RIe20d768_4443,RIe20aa68_4411,RIe207d68_4379,RIfca6460_6914,RIf1662e0_5622,RIe202908_4319,RIfe87b10_7888,RIfc58c10_6032,RIfc50ab0_5940,RIfccd790_7360,
        RIfccd1f0_7356,RIf160610_5556,RIf15e720_5534,RIfe87c78_7889,RIfe87f48_7891,RIfce7668_7655,RIfc86480_6550,RIfcd2218_7413,RIfcb01e0_7026,RIfc47b40_5838,
        RIfc84158_6525,RIfc4b920_5882,RIe1fa4d8_4225,RIfc4ba88_5883,RIfcb7530_7108,RIfcd58f0_7452,RIe1f5a50_4172,RIf153488_5407,RIf151ca0_5390,RIfc51e60_5954,
        RIe1f3728_4147,RIfc9aef8_6785,RIfcbaaa0_7146,RIfc52130_5956,RIe1ee430_4088,RIe1ebcd0_4060,RIe1e8fd0_4028,RIe1e62d0_3996,RIe1e35d0_3964,RIe1e08d0_3932,
        RIe1ddbd0_3900,RIe1daed0_3868,RIe1d81d0_3836,RIe1d27d0_3772,RIe1cfad0_3740,RIe1ccdd0_3708,RIe1ca0d0_3676,RIe1c73d0_3644,RIe1c46d0_3612,RIe1c19d0_3580,
        RIe1becd0_3548,RIfce0b88_7579,RIfc82808_6507,RIe1b9708_3487,RIe1b76b0_3464,RIfcd5bc0_7454,RIfcb69f0_7100,RIe1b54f0_3440,RIe1b4140_3426,RIfc89f90_6592,
        RIfce9af8_7681,RIe1b2958_3409,RIe1b0ea0_3390,RIfc4a138_5865,RIfc8a260_6594,RIe1ac850_3340,RIe1ab1d0_3324,RIe1a9010_3300,RIe1a6310_3268,RIe1a3610_3236,
        RIe1a0910_3204,RIe18ce10_2980,RIe179310_2756,RIe226c68_4731,RIe21b868_4603,RIe205068_4347,RIe1ff0c8_4279,RIe1f8480_4202,RIe1f0fc8_4119,RIe1d54d0_3804,
        RIe1bbfd0_3516,RIe1aee48_3367,RIe171480_2666,RIdec5810_711,RIdec2b10_679,RIfce6f60_7650,RIdebfe10_647,RIfc95228_6719,RIdebd110_615,RIdeba410_583,
        RIdeb7710_551,RIfe879a8_7887,RIdeb1d10_487,RIfcc16e8_7223,RIdeaf010_455,RIfca4f48_6899,RIdeaadf8_423,RIdea44f8_391,RIde9dbf8_359,RIee1cf48_4788,
        RIee1bfd0_4777,RIfc95660_6722,RIfcee148_7731,RIfe87840_7886,RIfe876d8_7885,RIde8a0f8_263,RIde85f58_243,RIfcb0780_7030,RIfcee9b8_7737,RIfc5f150_6104,
        RIfcdee00_7558,RIfcd8050_7480,RIe16ba80_2602,RIfca5380_6902,RIe1680d8_2561,RIe165810_2532,RIe162b10_2500,RIee377f8_5090,RIe15fe10_2468,RIee36448_5076,
        RIe15d110_2436,RIe157710_2372,RIe154a10_2340,RIfc3f3c8_5745,RIe151d10_2308,RIfcde9c8_7555,RIe14f010_2276,RIfc4a2a0_5866,RIe14c310_2244,RIe149610_2212,
        RIe146910_2180,RIfc62288_6139,RIee33478_5042,RIfc71b70_6316,RIee312b8_5018,RIe1411e0_2118,RIfe87570_7884,RIdf3cf28_2070,RIfe87408_7883,RIfcc99b0_7316,
        RIfccf0e0_7378,RIfcaeb60_7010,RIfcca220_7322,RIdf35bd8_1988,RIdf33748_1962,RIdf31588_1938,RIdf2f530_1915,RIee2be58_4958,RIee2a508_4940,RIee28ff0_4925,
        RIee27da8_4912,RIdf2a508_1858,RIdf28348_1834,RIdf265c0_1813,RIdf24b08_1794,RIfc74708_6347,RIfc42578_5777,RIfc43388_5787,RIfc745a0_6346,RIfcb0078_7025,
        RIdf1fc48_1738,RIfcaff10_7024,RIdf195a0_1665,RIdf173e0_1641,RIdf146e0_1609,RIdf119e0_1577,RIdf0ece0_1545,RIdf0bfe0_1513,RIdf092e0_1481,RIdf065e0_1449,
        RIdf038e0_1417,RIdefdee0_1353,RIdefb1e0_1321,RIdef84e0_1289,RIdef57e0_1257,RIdef2ae0_1225,RIdeefde0_1193,RIdeed0e0_1161,RIdeea3e0_1129,RIee257b0_4885,
        RIfca73d8_6925,RIee23e60_4867,RIfce66f0_7644,RIdee4cb0_1067,RIdee2f28_1046,RIdee0d68_1022,RIdeded10_999,RIfcca388_7323,RIfce6858_7645,RIfcceca8_7375,
        RIfcdc970_7532,RIded9b80_941,RIfeaaac0_8258,RIded5800_893,RIded3208_866,RIded0c10_839,RIdecdf10_807,RIdecb210_775,RIdec8510_743,RIdeb4a10_519,
        RIde972f8_327,RIe16e618_2633,RIe15a410_2404,RIe143c10_2148,RIdf38608_2018,RIdf2cc68_1886,RIdf1d4e8_1710,RIdf00be0_1385,RIdee76e0_1097,RIdedc448_970,
        RIde7d240_200,RIe19daa8_3171,RIe19ada8_3139,RIf1457c0_5250,RIe1980a8_3107,RIf1449b0_5240,RIe1953a8_3075,RIe1926a8_3043,RIe18f9a8_3011,RIe189fa8_2947,
        RIe1872a8_2915,RIf143ba0_5230,RIe1845a8_2883,RIfc912e0_6674,RIe1818a8_2851,RIe17eba8_2819,RIe17bea8_2787,RIfc915b0_6676,RIfcbe5b0_7188,RIfce3b58_7613,
        RIe175da0_2718,RIfceb448_7699,RIfcc7958_7293,RIfc42de8_5783,RIfc96e48_6739,RIfc7a810_6416,RIfc96ce0_6738,RIfcc7ac0_7294,RIe173be0_2694,RIfce39f0_7612,
        RIfc7a540_6414,RIfc91b50_6680,RIfc429b0_5780,RIfea9710_8244,RIe223e00_4698,RIfcd8488_7483,RIe221100_4666,RIfc920f0_6684,RIe21e400_4634,RIe218a00_4570,
        RIe215d00_4538,RIfc79e38_6409,RIe213000_4506,RIfcbee20_7194,RIe210300_4474,RIf168068_5643,RIe20d600_4442,RIe20a900_4410,RIe207c00_4378,RIfc5af38_6057,
        RIfcd73a8_7471,RIe2027a0_4318,RIe200ce8_4299,RIfcb2670_7052,RIfcdf940_7566,RIfc5b208_6059,RIfcbf3c0_7198,RIf1604a8_5555,RIf15e5b8_5533,RIfe872a0_7882,
        RIfe87138_7881,RIfc78920_6394,RIfec1158_8317,RIfc93338_6697,RIfcea368_7687,RIfcb23a0_7050,RIfc5bbe0_6066,RIfcede78_7729,RIe1fa370_4224,RIfcd4c48_7443,
        RIfce1dd0_7592,RIfcbf960_7202,RIe1f58e8_4171,RIfcbfc30_7204,RIfc78380_6390,RIfc93770_6700,RIe1f35c0_4146,RIfcb1f68_7047,RIfce1b00_7590,RIfc93a40_6702,
        RIe1ee2c8_4087,RIe1ebb68_4059,RIe1e8e68_4027,RIe1e6168_3995,RIe1e3468_3963,RIe1e0768_3931,RIe1dda68_3899,RIe1dad68_3867,RIe1d8068_3835,RIe1d2668_3771,
        RIe1cf968_3739,RIe1ccc68_3707,RIe1c9f68_3675,RIe1c7268_3643,RIe1c4568_3611,RIe1c1868_3579,RIe1beb68_3547,RIfcdec98_7557,RIfc94148_6707,RIe1b95a0_3486,
        RIe1b7548_3463,RIfcd12a0_7402,RIfceabd8_7693,RIe1b5388_3439,RIe1b3fd8_3425,RIfc94850_6712,RIfcd7c18_7477,RIe1b27f0_3408,RIe1b0d38_3389,RIfc76a30_6372,
        RIfce2640_7598,RIe1ac6e8_3339,RIe1ab068_3323,RIe1a8ea8_3299,RIe1a61a8_3267,RIe1a34a8_3235,RIe1a07a8_3203,RIe18cca8_2979,RIe1791a8_2755,RIe226b00_4730,
        RIe21b700_4602,RIe204f00_4346,RIe1fef60_4278,RIe1f8318_4201,RIe1f0e60_4118,RIe1d5368_3803,RIe1bbe68_3515,RIe1aece0_3366,RIe171318_2665,RIdec5c48_714,
        RIdec2f48_682,RIfc7c160_6434,RIdec0248_650,RIfcb38b8_7065,RIdebd548_618,RIdeba848_586,RIdeb7b48_554,RIfce7c08_7659,RIdeb2148_490,RIfce7aa0_7658,
        RIdeaf448_458,RIfca38c8_6883,RIdeab7d0_426,RIdea4ed0_394,RIde9e5d0_362,RIfc41e70_5772,RIfc5b0a0_6058,RIfcdbb60_7522,RIfc78650_6392,RIfea92d8_8241,
        RIde8e5e0_284,RIfea0d40_8174,RIfea0bd8_8173,RIfcdf508_7563,RIfcb1b30_7044,RIfc5ccc0_6078,RIfcb16f8_7041,RIfc77b10_6384,RIe16beb8_2605,RIe169e60_2582,
        RIe168510_2564,RIe165c48_2535,RIe162f48_2503,RIfc4f9d0_5928,RIe160248_2471,RIfc4e8f0_5916,RIe15d548_2439,RIe157b48_2375,RIe154e48_2343,RIfc4e1e8_5911,
        RIe152148_2311,RIfc868b8_6553,RIe14f448_2279,RIfc865e8_6551,RIe14c748_2247,RIe149a48_2215,RIe146d48_2183,RIfc9eb70_6828,RIfc9ecd8_6829,RIfcc5630_7268,
        RIfc83bb8_6521,RIe141618_2121,RIfea0ea8_8175,RIdf3d1f8_2072,RIdf3ac00_2045,RIee308e0_5011,RIfcd3cd0_7432,RIfc84e00_6534,RIfc834b0_6516,RIdf36010_1991,
        RIdf33a18_1964,RIdf31858_1940,RIdf2f968_1918,RIee2c128_4960,RIee2a7d8_4942,RIee292c0_4927,RIee28078_4914,RIdf2a940_1861,RIdf28780_1837,RIfea0a70_8172,
        RIfea0908_8171,RIfcd4f18_7445,RIfca0628_6847,RIdf23050_1775,RIfcd3190_7424,RIdf21b38_1760,RIdf20080_1741,RIdf1b328_1686,RIdf199d8_1668,RIdf17818_1644,
        RIdf14b18_1612,RIdf11e18_1580,RIdf0f118_1548,RIdf0c418_1516,RIdf09718_1484,RIdf06a18_1452,RIdf03d18_1420,RIdefe318_1356,RIdefb618_1324,RIdef8918_1292,
        RIdef5c18_1260,RIdef2f18_1228,RIdef0218_1196,RIdeed518_1164,RIdeea818_1132,RIfcdf3a0_7562,RIfca5218_6901,RIfcdc538_7529,RIfcdc6a0_7530,RIdee50e8_1070,
        RIdee3360_1049,RIfea07a0_8170,RIdedefe0_1001,RIfcb0d20_7034,RIfcd4978_7441,RIfca49a8_6895,RIfca1708_6859,RIded9fb8_944,RIded79c0_917,RIded5ad0_895,
        RIfeab498_8265,RIded1048_842,RIdece348_810,RIdecb648_778,RIdec8948_746,RIdeb4e48_522,RIde97cd0_330,RIe16ea50_2636,RIe15a848_2407,RIe144048_2151,
        RIdf38a40_2021,RIdf2d0a0_1889,RIdf1d920_1713,RIdf01018_1388,RIdee7b18_1100,RIdedc880_973,RIde7dc18_203,RIe19dee0_3174,RIe19b1e0_3142,RIfc67580_6198,
        RIe1984e0_3110,RIfccb030_7332,RIe1957e0_3078,RIe192ae0_3046,RIe18fde0_3014,RIe18a3e0_2950,RIe1876e0_2918,RIfc6a550_6232,RIe1849e0_2886,RIfcaa7e0_6962,
        RIe181ce0_2854,RIe17efe0_2822,RIe17c2e0_2790,RIfc65d98_6181,RIfc65690_6176,RIe1772b8_2733,RIfea0638_8169,RIfcca928_7327,RIfc607d0_6120,RIfc65258_6173,
        RIee3d798_5158,RIee3c3e8_5144,RIfca9430_6948,RIee39f58_5118,RIe174018_2697,RIfcecf00_7718,RIfc650f0_6172,RIf16e5a8_5715,RIfc43a90_5792,RIfc65528_6175,
        RIe224238_4701,RIfca9f70_6956,RIe221538_4669,RIfc6b4c8_6243,RIe21e838_4637,RIe218e38_4573,RIe216138_4541,RIfc3fda0_5752,RIe213438_4509,RIfc61310_6128,
        RIe210738_4477,RIfc60c08_6123,RIe20da38_4445,RIe20ad38_4413,RIe208038_4381,RIfc66ba8_6191,RIfccbcd8_7341,RIe202bd8_4321,RIe200fb8_4301,RIfcadbe8_6999,
        RIfccbe40_7342,RIfca7540_6926,RIfc6a3e8_6231,RIfca6898_6917,RIfc73358_6333,RIe1fd070_4256,RIe1fbe28_4243,RIfcc2660_7234,RIfc44468_5799,RIf15a940_5490,
        RIfca7270_6924,RIfc5e070_6092,RIfc5dda0_6090,RIfc7e050_6456,RIe1fa7a8_4227,RIfc5d968_6087,RIfcd9568_7495,RIfc8d668_6631,RIe1f5d20_4174,RIfca4138_6889,
        RIfc8cdf8_6625,RIfcc7c28_7295,RIe1f39f8_4149,RIfc99440_6766,RIfcbc3f0_7164,RIfc5a128_6047,RIe1ee700_4090,RIe1ebfa0_4062,RIe1e92a0_4030,RIe1e65a0_3998,
        RIe1e38a0_3966,RIe1e0ba0_3934,RIe1ddea0_3902,RIe1db1a0_3870,RIe1d84a0_3838,RIe1d2aa0_3774,RIe1cfda0_3742,RIe1cd0a0_3710,RIe1ca3a0_3678,RIe1c76a0_3646,
        RIe1c49a0_3614,RIe1c1ca0_3582,RIe1befa0_3550,RIf14cde0_5334,RIf14bb98_5321,RIe1b99d8_3489,RIe1b7980_3466,RIfc4c460_5890,RIfc9e738_6825,RIe1b5658_3441,
        RIfec54d8_8365,RIf149168_5291,RIf147f20_5278,RIe1b2ac0_3410,RIe1b1170_3392,RIf1473e0_5270,RIf1468a0_5262,RIe1acb20_3342,RIe1ab338_3325,RIe1a92e0_3302,
        RIe1a65e0_3270,RIe1a38e0_3238,RIe1a0be0_3206,RIe18d0e0_2982,RIe1795e0_2758,RIe226f38_4733,RIe21bb38_4605,RIe205338_4349,RIe1ff398_4281,RIe1f8750_4204,
        RIe1f1298_4121,RIe1d57a0_3806,RIe1bc2a0_3518,RIe1af118_3369,RIe171750_2668,RIdec5ae0_713,RIdec2de0_681,RIfc82268_6503,RIdec00e0_649,RIfcb8d18_7125,
        RIdebd3e0_617,RIdeba6e0_585,RIdeb79e0_553,RIfcb9858_7133,RIdeb1fe0_489,RIfc9efa8_6831,RIdeaf2e0_457,RIfce0750_7576,RIdeab488_425,RIdea4b88_393,
        RIde9e288_361,RIee1d0b0_4789,RIee1c138_4778,RIfcd0e68_7399,RIfc76d00_6374,RIfe89028_7903,RIfe88d58_7901,RIfe88ec0_7902,RIfe88bf0_7900,RIfcda7b0_7508,
        RIfc4d810_5904,RIfc52dd8_5965,RIfcde590_7552,RIfc4f868_5927,RIe16bd50_2604,RIfc68930_6212,RIe1683a8_2563,RIe165ae0_2534,RIe162de0_2502,RIfe88a88_7899,
        RIe1600e0_2470,RIfcc9140_7310,RIe15d3e0_2438,RIe1579e0_2374,RIe154ce0_2342,RIfc698a8_6223,RIe151fe0_2310,RIee35098_5062,RIe14f2e0_2278,RIfcc0338_7209,
        RIe14c5e0_2246,RIe1498e0_2214,RIe146be0_2182,RIfc88208_6571,RIfc85670_6540,RIfc81f98_6501,RIfcc4f28_7263,RIe1414b0_2120,RIe13f188_2095,RIdf3d090_2071,
        RIdf3aa98_2044,RIfcd2920_7418,RIfc7d7e0_6450,RIfc49760_5858,RIfce5a48_7635,RIdf35ea8_1990,RIdf338b0_1963,RIfe88920_7898,RIdf2f800_1917,RIee2bfc0_4959,
        RIee2a670_4941,RIee29158_4926,RIee27f10_4913,RIdf2a7d8_1860,RIdf28618_1836,RIdf26890_1815,RIdf24dd8_1796,RIfcad918_6997,RIfc69fb0_6228,RIfc63368_6151,
        RIfc623f0_6140,RIfc60938_6121,RIdf1ff18_1740,RIfcba500_7142,RIdf19870_1667,RIdf176b0_1643,RIdf149b0_1611,RIdf11cb0_1579,RIdf0efb0_1547,RIdf0c2b0_1515,
        RIdf095b0_1483,RIdf068b0_1451,RIdf03bb0_1419,RIdefe1b0_1355,RIdefb4b0_1323,RIdef87b0_1291,RIdef5ab0_1259,RIdef2db0_1227,RIdef00b0_1195,RIdeed3b0_1163,
        RIdeea6b0_1131,RIfcc9848_7315,RIfc69a10_6224,RIfcacc70_6988,RIfccbfa8_7343,RIdee4f80_1069,RIdee31f8_1048,RIdee1038_1024,RIdedee78_1000,RIfc84590_6528,
        RIfc9bba0_6794,RIee21b38_4842,RIfc47168_5831,RIded9e50_943,RIded7858_916,RIfe887b8_7897,RIded34d8_868,RIded0ee0_841,RIdece1e0_809,RIdecb4e0_777,
        RIdec87e0_745,RIdeb4ce0_521,RIde97988_329,RIe16e8e8_2635,RIe15a6e0_2406,RIe143ee0_2150,RIdf388d8_2020,RIdf2cf38_1888,RIdf1d7b8_1712,RIdf00eb0_1387,
        RIdee79b0_1099,RIdedc718_972,RIde7d8d0_202,RIe19dd78_3173,RIe19b078_3141,RIfca1438_6857,RIe198378_3109,RIfca35f8_6881,RIe195678_3077,RIe192978_3045,
        RIe18fc78_3013,RIe18a278_2949,RIe187578_2917,RIfcba230_7140,RIe184878_2885,RIf142d90_5220,RIe181b78_2853,RIe17ee78_2821,RIe17c178_2789,RIfc9be70_6796,
        RIfc9bd08_6795,RIfc4ccd0_5896,RIe176070_2720,RIfc87c68_6567,RIfc87b00_6566,RIfcc4c58_7261,RIfc4fca0_5930,RIfc4f598_5925,RIfc876c8_6563,RIfc4dae0_5906,
        RIe173eb0_2696,RIfcb9420_7130,RIfc4e080_5910,RIfc4e350_5912,RIfc9d388_6811,RIfc40a48_5761,RIe2240d0_4700,RIfc85508_6539,RIe2213d0_4668,RIfc9ba38_6793,
        RIe21e6d0_4636,RIe218cd0_4572,RIe215fd0_4540,RIfc52c70_5964,RIe2132d0_4508,RIfca3760_6882,RIe2105d0_4476,RIfc97988_6747,RIe20d8d0_4444,RIe20abd0_4412,
        RIe207ed0_4380,RIfceb5b0_7700,RIfcddbb8_7545,RIe202a70_4320,RIe200e50_4300,RIfc73d30_6340,RIfcaf100_7014,RIfc71468_6311,RIfcdcad8_7533,RIfcdda50_7544,
        RIfca8620_6938,RIe1fcf08_4255,RIe1fbcc0_4242,RIfc6c008_6251,RIfcdd1e0_7538,RIfca9700_6950,RIfca92c8_6947,RIfcce5a0_7370,RIfc6ba68_6247,RIfc6f410_6288,
        RIe1fa640_4226,RIfcce000_7366,RIfc53918_5973,RIfcce708_7371,RIe1f5bb8_4173,RIf1535f0_5408,RIf151e08_5391,RIfc72db8_6329,RIe1f3890_4148,RIf14fc48_5367,
        RIfc72c50_6328,RIfc73e98_6341,RIe1ee598_4089,RIe1ebe38_4061,RIe1e9138_4029,RIe1e6438_3997,RIe1e3738_3965,RIe1e0a38_3933,RIe1ddd38_3901,RIe1db038_3869,
        RIe1d8338_3837,RIe1d2938_3773,RIe1cfc38_3741,RIe1ccf38_3709,RIe1ca238_3677,RIe1c7538_3645,RIe1c4838_3613,RIe1c1b38_3581,RIe1bee38_3549,RIfcb8a48_7123,
        RIfcb84a8_7119,RIe1b9870_3488,RIe1b7818_3465,RIfc85940_6542,RIfc9e198_6821,RIfeac140_8274,RIe1b42a8_3427,RIfc518c0_5950,RIfc838e8_6519,RIfe884e8_7895,
        RIe1b1008_3391,RIfcc5900_7270,RIfc82ad8_6509,RIe1ac9b8_3341,RIfe88650_7896,RIe1a9178_3301,RIe1a6478_3269,RIe1a3778_3237,RIe1a0a78_3205,RIe18cf78_2981,
        RIe179478_2757,RIe226dd0_4732,RIe21b9d0_4604,RIe2051d0_4348,RIe1ff230_4280,RIe1f85e8_4203,RIe1f1130_4120,RIe1d5638_3805,RIe1bc138_3517,RIe1aefb0_3368,
        RIe1715e8_2667,RIdec5f18_716,RIdec3218_684,RIee20350_4825,RIdec0518_652,RIee1f6a8_4816,RIdebd818_620,RIdebab18_588,RIdeb7e18_556,RIfce4da0_7626,
        RIdeb2418_492,RIfcea908_7691,RIdeaf718_460,RIfce20a0_7594,RIdeabe60_428,RIdea5560_396,RIde9ec60_364,RIfce6420_7642,RIee1c2a0_4779,RIfc75950_6360,
        RIee1ad88_4764,RIde920f0_302,RIfea4148_8211,RIfeaa688_8255,RIfea3fe0_8210,RIde82790_226,RIfc6f848_6291,RIfc5dc38_6089,RIfc76b98_6373,RIfcae2f0_7004,
        RIe16c020_2606,RIe16a130_2584,RIe1687e0_2566,RIe165f18_2537,RIe163218_2505,RIfcadd50_7000,RIe160518_2473,RIfc55268_5991,RIe15d818_2441,RIe157e18_2377,
        RIe155118_2345,RIfc45548_5811,RIe152418_2313,RIfc498c8_5859,RIe14f718_2281,RIfcbda70_7180,RIe14ca18_2249,RIe149d18_2217,RIe147018_2185,RIee34828_5056,
        RIee33748_5044,RIee32668_5032,RIee31588_5020,RIe1418e8_2123,RIe13f458_2097,RIdf3d360_2073,RIdf3aed0_2047,RIfc526d0_5960,RIfc42848_5779,RIfcae9f8_7009,
        RIfcb7260_7106,RIfea42b0_8212,RIdf33ce8_1966,RIdf31b28_1942,RIdf2fc38_1920,RIee2c3f8_4962,RIfc4cfa0_5898,RIfc572c0_6014,RIfc4f430_5924,RIfea3e78_8209,
        RIdf28a50_1839,RIdf26b60_1817,RIdf250a8_1798,RIfc9b600_6790,RIfcb9df8_7137,RIdf23320_1777,RIfc86318_6549,RIfeabfd8_8273,RIdf201e8_1742,RIdf1b5f8_1688,
        RIdf19ca8_1670,RIdf17ae8_1646,RIdf14de8_1614,RIdf120e8_1582,RIdf0f3e8_1550,RIdf0c6e8_1518,RIdf099e8_1486,RIdf06ce8_1454,RIdf03fe8_1422,RIdefe5e8_1358,
        RIdefb8e8_1326,RIdef8be8_1294,RIdef5ee8_1262,RIdef31e8_1230,RIdef04e8_1198,RIdeed7e8_1166,RIdeeaae8_1134,RIfc89018_6581,RIfcc54c8_7267,RIfc89180_6582,
        RIfc4b380_5878,RIdee53b8_1072,RIdee34c8_1050,RIfea3d10_8208,RIdedf148_1002,RIfcae188_7003,RIfc4b0b0_5876,RIfc74870_6348,RIfce4968_7623,RIdeda288_946,
        RIded7c90_919,RIded5da0_897,RIded3640_869,RIded1318_844,RIdece618_812,RIdecb918_780,RIdec8c18_748,RIdeb5118_524,RIde98360_332,RIe16ed20_2638,
        RIe15ab18_2409,RIe144318_2153,RIdf38d10_2023,RIdf2d370_1891,RIdf1dbf0_1715,RIdf012e8_1390,RIdee7de8_1102,RIdedcb50_975,RIde7e2a8_205,RIe19e1b0_3176,
        RIe19b4b0_3144,RIfc9cf50_6808,RIe1987b0_3112,RIfc87290_6560,RIe195ab0_3080,RIe192db0_3048,RIe1900b0_3016,RIe18a6b0_2952,RIe1879b0_2920,RIfc842c0_6526,
        RIe184cb0_2888,RIfc83a50_6520,RIe181fb0_2856,RIe17f2b0_2824,RIe17c5b0_2792,RIfc9d0b8_6809,RIfc9e030_6820,RIe177420_2734,RIe176340_2722,RIfc4f700_5926,
        RIfcc4820_7258,RIfc4fb38_5929,RIfce8040_7662,RIee3c6b8_5146,RIee3b308_5132,RIfc812f0_6492,RIe174180_2698,RIfcd3028_7423,RIfc7f400_6470,RIfc46a60_5826,
        RIfc472d0_5832,RIf16cc58_5697,RIe224508_4703,RIfc7d3a8_6447,RIe221808_4671,RIfc97c58_6749,RIe21eb08_4639,RIe219108_4575,RIe216408_4543,RIfcdbe30_7524,
        RIe213708_4511,RIf169580_5658,RIe210a08_4479,RIfca4570_6892,RIe20dd08_4447,RIe20b008_4415,RIe208308_4383,RIfc7b080_6422,RIfc59cf0_6044,RIfea9b48_8247,
        RIfea4418_8213,RIfc79cd0_6408,RIfcd19a8_7407,RIfcc81c8_7299,RIf162230_5576,RIf160778_5557,RIf15e888_5535,RIfea4580_8214,RIfea46e8_8215,RIfc77f48_6387,
        RIfc41fd8_5773,RIf15aaa8_5491,RIfc7c430_6436,RIf159158_5473,RIf157f10_5460,RIfcae890_7008,RIe1faa78_4229,RIfc4a840_5870,RIfc4ed28_5919,RIfce0e58_7581,
        RIe1f5ff0_4176,RIf153758_5409,RIf151f70_5392,RIfccb468_7335,RIe1f3cc8_4151,RIfc68ed0_6216,RIfc6d250_6264,RIfca9ca0_6954,RIe1ee9d0_4092,RIe1ec270_4064,
        RIe1e9570_4032,RIe1e6870_4000,RIe1e3b70_3968,RIe1e0e70_3936,RIe1de170_3904,RIe1db470_3872,RIe1d8770_3840,RIe1d2d70_3776,RIe1d0070_3744,RIe1cd370_3712,
        RIe1ca670_3680,RIe1c7970_3648,RIe1c4c70_3616,RIe1c1f70_3584,RIe1bf270_3552,RIfc784e8_6391,RIfcbef88_7195,RIe1b9ca8_3491,RIe1b7ae8_3467,RIfcc20c0_7230,
        RIfca6190_6912,RIe1b5928_3443,RIe1b4410_3428,RIfcb81d8_7117,RIfcc5090_7264,RIe1b2d90_3412,RIe1b1440_3394,RIfcd5350_7448,RIfcb9588_7131,RIe1acc88_3343,
        RIe1ab4a0_3326,RIe1a95b0_3304,RIe1a68b0_3272,RIe1a3bb0_3240,RIe1a0eb0_3208,RIe18d3b0_2984,RIe1798b0_2760,RIe227208_4735,RIe21be08_4607,RIe205608_4351,
        RIe1ff668_4283,RIe1f8a20_4206,RIe1f1568_4123,RIe1d5a70_3808,RIe1bc570_3520,RIe1af3e8_3371,RIe171a20_2670,RIdec5db0_715,RIdec30b0_683,RIee201e8_4824,
        RIdec03b0_651,RIfcaf538_7017,RIdebd6b0_619,RIdeba9b0_587,RIdeb7cb0_555,RIfc40fe8_5765,RIdeb22b0_491,RIfcd08c8_7395,RIdeaf5b0_459,RIee1dd58_4798,
        RIdeabb18_427,RIdea5218_395,RIde9e918_363,RIee1d218_4790,RIfcedd10_7728,RIfce62b8_7641,RIfcc92a8_7311,RIde91da8_301,RIde8e928_285,RIde8a788_265,
        RIde865e8_245,RIde82448_225,RIfea1448_8179,RIfc750e0_6354,RIfcc19b8_7225,RIfced8d8_7725,RIfec5eb0_8372,RIe169fc8_2583,RIe168678_2565,RIe165db0_2536,
        RIe1630b0_2504,RIfccfc20_7386,RIe1603b0_2472,RIee365b0_5077,RIe15d6b0_2440,RIe157cb0_2376,RIe154fb0_2344,RIfea1718_8181,RIe1522b0_2312,RIee35200_5063,
        RIe14f5b0_2280,RIfcb0348_7027,RIe14c8b0_2248,RIe149bb0_2216,RIe146eb0_2184,RIfc73790_6336,RIfcdf238_7561,RIee32500_5031,RIfc94f58_6717,RIe141780_2122,
        RIe13f2f0_2096,RIfec5be0_8370,RIdf3ad68_2046,RIfea15b0_8180,RIfc5fb28_6111,RIfcae728_7007,RIfc74438_6345,RIdf36178_1992,RIdf33b80_1965,RIdf319c0_1941,
        RIdf2fad0_1919,RIee2c290_4961,RIee2a940_4943,RIfc70658_6301,RIfc704f0_6300,RIdf2aaa8_1862,RIdf288e8_1838,RIdf269f8_1816,RIdf24f40_1797,RIfc64b50_6168,
        RIfccaa90_7328,RIdf231b8_1776,RIfcad4e0_6994,RIdf21ca0_1761,RIfeaad90_8260,RIdf1b490_1687,RIdf19b40_1669,RIdf17980_1645,RIdf14c80_1613,RIdf11f80_1581,
        RIdf0f280_1549,RIdf0c580_1517,RIdf09880_1485,RIdf06b80_1453,RIdf03e80_1421,RIdefe480_1357,RIdefb780_1325,RIdef8a80_1293,RIdef5d80_1261,RIdef3080_1229,
        RIdef0380_1197,RIdeed680_1165,RIdeea980_1133,RIfc595e8_6039,RIfcac568_6983,RIfcccf20_7354,RIfccd358_7357,RIdee5250_1071,RIfea7f28_8227,RIdee11a0_1025,
        RIfea12e0_8178,RIfc679b8_6201,RIee22510_4849,RIfc6dd90_6272,RIfc6cb48_6259,RIdeda120_945,RIded7b28_918,RIded5c38_896,RIfec5d48_8371,RIded11b0_843,
        RIdece4b0_811,RIdecb7b0_779,RIdec8ab0_747,RIdeb4fb0_523,RIde98018_331,RIe16ebb8_2637,RIe15a9b0_2408,RIe1441b0_2152,RIdf38ba8_2022,RIdf2d208_1890,
        RIdf1da88_1714,RIdf01180_1389,RIdee7c80_1101,RIdedc9e8_974,RIde7df60_204,RIe19e048_3175,RIe19b348_3143,RIfcc3ce0_7250,RIe198648_3111,RIfc7efc8_6467,
        RIe195948_3079,RIe192c48_3047,RIe18ff48_3015,RIe18a548_2951,RIe187848_2919,RIfc46790_5824,RIe184b48_2887,RIfc98d38_6761,RIe181e48_2855,RIe17f148_2823,
        RIe17c448_2791,RIfcb5d48_7091,RIfc995a8_6767,RIfc9a3b8_6777,RIe1761d8_2721,RIfc54188_5979,RIfcd2bf0_7420,RIfc8b778_6609,RIfc7dee8_6455,RIee3c550_5145,
        RIfc8c420_6618,RIee3a0c0_5119,RIfeaba38_8269,RIfc46628_5823,RIfcbc288_7163,RIf16e710_5716,RIfc8fdc8_6659,RIfc48c20_5850,RIe2243a0_4702,RIfca0358_6845,
        RIe2216a0_4670,RIfc9a688_6779,RIe21e9a0_4638,RIe218fa0_4574,RIe2162a0_4542,RIfc456b0_5812,RIe2135a0_4510,RIf169418_5657,RIe2108a0_4478,RIfc8bfe8_6615,
        RIe20dba0_4446,RIe20aea0_4414,RIe2081a0_4382,RIfc8c9c0_6622,RIfc7f568_6471,RIe202d40_4322,RIe201120_4302,RIfce2910_7600,RIfc487e8_5847,RIfc46d30_5828,
        RIfc992d8_6765,RIfca2680_6870,RIfc44a08_5803,RIe1fd1d8_4257,RIe1fbf90_4244,RIfc580d0_6024,RIfcbdbd8_7181,RIfc8dd70_6636,RIfce01b0_7572,RIfc7bbc0_6430,
        RIfc90368_6663,RIfc7b8f0_6428,RIe1fa910_4228,RIfcd8b90_7488,RIfc43ec8_5795,RIfc7b788_6427,RIe1f5e88_4175,RIfc7b350_6424,RIfc90d40_6670,RIfca3490_6880,
        RIe1f3b60_4150,RIfc91010_6672,RIfcdb728_7519,RIfcd8758_7485,RIe1ee868_4091,RIe1ec108_4063,RIe1e9408_4031,RIe1e6708_3999,RIe1e3a08_3967,RIe1e0d08_3935,
        RIe1de008_3903,RIe1db308_3871,RIe1d8608_3839,RIe1d2c08_3775,RIe1cff08_3743,RIe1cd208_3711,RIe1ca508_3679,RIe1c7808_3647,RIe1c4b08_3615,RIe1c1e08_3583,
        RIe1bf108_3551,RIf14cf48_5335,RIfc78d58_6397,RIe1b9b40_3490,RIfec5910_8368,RIfc78a88_6395,RIfcd51e8_7447,RIe1b57c0_3442,RIfea1010_8176,RIf1492d0_5292,
        RIfec5a78_8369,RIe1b2c28_3411,RIe1b12d8_3393,RIfec5640_8366,RIf146a08_5263,RIfec57a8_8367,RIfea1178_8177,RIe1a9448_3303,RIe1a6748_3271,RIe1a3a48_3239,
        RIe1a0d48_3207,RIe18d248_2983,RIe179748_2759,RIe2270a0_4734,RIe21bca0_4606,RIe2054a0_4350,RIe1ff500_4282,RIe1f88b8_4205,RIe1f1400_4122,RIe1d5908_3807,
        RIe1bc408_3519,RIe1af280_3370,RIe1718b8_2669,RIdec6350_719,RIdec3650_687,RIfcaf3d0_7016,RIdec0950_655,RIfc6a280_6230,RIdebdc50_623,RIdebaf50_591,
        RIdeb8250_559,RIfc42f50_5784,RIdeb2850_495,RIfc981f8_6753,RIdeafb50_463,RIfc8c6f0_6620,RIdeac838_431,RIdea5f38_399,RIde9f638_367,RIee1d4e8_4792,
        RIfcda648_7507,RIfcc6440_7278,RIfcd5620_7450,RIde92ac8_305,RIfea34a0_8202,RIfea31d0_8200,RIfea3338_8201,RIfcb6b58_7101,RIfcb6888_7099,RIfc9dd60_6818,
        RIee19708_4748,RIfc50c18_5941,RIe16c458_2609,RIfc80a80_6486,RIfec62e8_8375,RIe166350_2540,RIe163650_2508,RIee37d98_5094,RIe160950_2476,RIfcaa678_6961,
        RIe15dc50_2444,RIe158250_2380,RIe155550_2348,RIfea3ba8_8207,RIe152850_2316,RIee35638_5066,RIe14fb50_2284,RIfc62f30_6148,RIe14ce50_2252,RIe14a150_2220,
        RIe147450_2188,RIfc97f28_6751,RIfc89888_6587,RIfc8f558_6653,RIfc52838_5961,RIe141bb8_2125,RIe13f890_2100,RIdf3d798_2076,RIdf3b308_2050,RIee30a48_5012,
        RIfc568e8_6007,RIee2e9f0_4989,RIee2dbe0_4979,RIdf365b0_1995,RIfea38d8_8205,RIfea3a40_8206,RIdf2ff08_1922,RIee2c6c8_4964,RIee2ac10_4945,RIee29590_4929,
        RIee28348_4916,RIdf2ad78_1864,RIdf28e88_1842,RIfea3608_8203,RIfea3770_8204,RIfcc0d10_7216,RIfc75c20_6362,RIfca50b0_6900,RIfc74e10_6352,RIfcc9410_7312,
        RIdf20620_1745,RIfc73628_6335,RIdf1a0e0_1673,RIdf17f20_1649,RIdf15220_1617,RIdf12520_1585,RIdf0f820_1553,RIdf0cb20_1521,RIdf09e20_1489,RIdf07120_1457,
        RIdf04420_1425,RIdefea20_1361,RIdefbd20_1329,RIdef9020_1297,RIdef6320_1265,RIdef3620_1233,RIdef0920_1201,RIdeedc20_1169,RIdeeaf20_1137,RIfcab8c0_6974,
        RIfc7c598_6437,RIfc5beb0_6068,RIfc58ee0_6034,RIdee5688_1074,RIdee3798_1052,RIdee15d8_1028,RIdedf580_1005,RIfcb3048_7059,RIfc72ae8_6327,RIfca3d00_6886,
        RIfcb6450_7096,RIdeda558_948,RIded7f60_921,RIfea3068_8199,RIded3a78_872,RIded1750_847,RIdecea50_815,RIdecbd50_783,RIdec9050_751,RIdeb5550_527,
        RIde98d38_335,RIe16f158_2641,RIe15af50_2412,RIe144750_2156,RIdf39148_2026,RIdf2d7a8_1894,RIdf1e028_1718,RIdf01720_1393,RIdee8220_1105,RIdedcf88_978,
        RIde7ec80_208,RIe19e5e8_3179,RIe19b8e8_3147,RIfca84b8_6937,RIe198be8_3115,RIfc846f8_6529,RIe195ee8_3083,RIe1931e8_3051,RIe1904e8_3019,RIe18aae8_2955,
        RIe187de8_2923,RIfce2be0_7602,RIe1850e8_2891,RIfc8e310_6640,RIe1823e8_2859,RIe17f6e8_2827,RIe17c9e8_2795,RIfcd1570_7404,RIfccc278_7345,RIf1404c8_5191,
        RIfea2d98_8197,RIfcc1b20_7226,RIfc60398_6117,RIee3e5a8_5168,RIee3da68_5160,RIfc642e0_6162,RIfca7f18_6933,RIee3a228_5120,RIfec6180_8374,RIfca9598_6949,
        RIfc5c720_6074,RIfc6bea0_6250,RIfccaec8_7331,RIfc44cd8_5805,RIe224940_4706,RIfcb6180_7094,RIe221c40_4674,RIfc55ad8_5997,RIe21ef40_4642,RIe219540_4578,
        RIe216840_4546,RIfc4dc48_5907,RIe213b40_4514,RIfcdcf10_7536,RIe210e40_4482,RIfcab1b8_6969,RIe20e140_4450,RIe20b440_4418,RIe208740_4386,RIfce3720_7610,
        RIfc64178_6161,RIe203178_4325,RIe201558_4305,RIfcd2ec0_7422,RIf164828_5603,RIfc7f838_6473,RIf162398_5577,RIfcc9c80_7318,RIfca8bc0_6942,RIfea2ac8_8195,
        RIfea2c30_8196,RIfc59318_6037,RIfc4f160_5922,RIf15ac10_5492,RIfcebf88_7707,RIfcbb040_7150,RIfca1870_6860,RIfc93d10_6704,RIe1faeb0_4232,RIf1565c0_5442,
        RIf155a80_5434,RIfc45c50_5816,RIe1f6428_4179,RIfccdbc8_7363,RIfcccae8_7351,RIfca6cd0_6920,RIfec6018_8373,RIfc64010_6160,RIfc434f0_5788,RIfc4c028_5887,
        RIe1eee08_4095,RIe1ec6a8_4067,RIe1e99a8_4035,RIe1e6ca8_4003,RIe1e3fa8_3971,RIe1e12a8_3939,RIe1de5a8_3907,RIe1db8a8_3875,RIe1d8ba8_3843,RIe1d31a8_3779,
        RIe1d04a8_3747,RIe1cd7a8_3715,RIe1caaa8_3683,RIe1c7da8_3651,RIe1c50a8_3619,RIe1c23a8_3587,RIe1bf6a8_3555,RIfc63908_6155,RIfc6bd38_6249,RIe1ba0e0_3494,
        RIe1b7f20_3470,RIfc66fe0_6194,RIfc92ac8_6691,RIe1b5d60_3446,RIfea2f00_8198,RIfc9bfd8_6797,RIfc50d80_5942,RIe1b31c8_3415,RIe1b1878_3397,RIfc4df18_5909,
        RIfc9d658_6813,RIe1ad0c0_3346,RIe1ab8d8_3329,RIe1a99e8_3307,RIe1a6ce8_3275,RIe1a3fe8_3243,RIe1a12e8_3211,RIe18d7e8_2987,RIe179ce8_2763,RIe227640_4738,
        RIe21c240_4610,RIe205a40_4354,RIe1ffaa0_4286,RIe1f8e58_4209,RIe1f19a0_4126,RIe1d5ea8_3811,RIe1bc9a8_3523,RIe1af820_3374,RIe171e58_2673,RIdec61e8_718,
        RIdec34e8_686,RIee20620_4827,RIdec07e8_654,RIfc4b7b8_5881,RIdebdae8_622,RIdebade8_590,RIdeb80e8_558,RIfc41150_5766,RIdeb26e8_494,RIfc87830_6564,
        RIdeaf9e8_462,RIee1dec0_4799,RIdeac4f0_430,RIdea5bf0_398,RIde9f2f0_366,RIee1d380_4791,RIfc77c78_6385,RIfc84f68_6535,RIfc6ff50_6296,RIde92780_304,
        RIde8efb8_287,RIde8ae18_267,RIde86c78_247,RIee1a680_4759,RIee19f78_4754,RIfcd7240_7470,RIfcbeb50_7192,RIfc76328_6367,RIe16c2f0_2608,RIee388d8_5102,
        RIfea20f0_8188,RIe1661e8_2539,RIe1634e8_2507,RIee37c30_5093,RIe1607e8_2475,RIfce7500_7654,RIe15dae8_2443,RIe1580e8_2379,RIe1553e8_2347,RIfc3f698_5747,
        RIe1526e8_2315,RIee354d0_5065,RIe14f9e8_2283,RIfc83e88_6523,RIe14cce8_2251,RIe149fe8_2219,RIe1472e8_2187,RIfcea4d0_7688,RIfcb7ad0_7112,RIfc695d8_6221,
        RIfc51a28_5951,RIe141a50_2124,RIe13f728_2099,RIdf3d630_2075,RIdf3b1a0_2049,RIfca9e08_6955,RIee2fda0_5003,RIfc88a78_6577,RIee2da78_4978,RIdf36448_1994,
        RIdf33fb8_1968,RIdf31df8_1944,RIfea2258_8189,RIee2c560_4963,RIee2aaa8_4944,RIee29428_4928,RIee281e0_4915,RIdf2ac10_1863,RIdf28d20_1841,RIfea27f8_8193,
        RIfea2960_8194,RIfcdabe8_7511,RIfca08f8_6849,RIfc8b1d8_6605,RIfc49058_5853,RIfca0a60_6850,RIdf204b8_1744,RIfc99cb0_6772,RIdf19f78_1672,RIdf17db8_1648,
        RIdf150b8_1616,RIdf123b8_1584,RIdf0f6b8_1552,RIdf0c9b8_1520,RIdf09cb8_1488,RIdf06fb8_1456,RIdf042b8_1424,RIdefe8b8_1360,RIdefbbb8_1328,RIdef8eb8_1296,
        RIdef61b8_1264,RIdef34b8_1232,RIdef07b8_1200,RIdeedab8_1168,RIdeeadb8_1136,RIfcd1f48_7411,RIfc57f68_6023,RIfcbe2e0_7186,RIfcd8fc8_7491,RIdee5520_1073,
        RIfea2690_8192,RIdee1470_1027,RIdedf418_1004,RIfc57b30_6020,RIfcb35e8_7063,RIfcbd7a0_7178,RIfc91178_6673,RIfea2528_8191,RIded7df8_920,RIfea23c0_8190,
        RIded3910_871,RIded15e8_846,RIdece8e8_814,RIdecbbe8_782,RIdec8ee8_750,RIdeb53e8_526,RIde989f0_334,RIe16eff0_2640,RIe15ade8_2411,RIe1445e8_2155,
        RIdf38fe0_2025,RIdf2d640_1893,RIdf1dec0_1717,RIdf015b8_1392,RIdee80b8_1104,RIdedce20_977,RIde7e938_207,RIe19e480_3178,RIe19b780_3146,RIfccc980_7350,
        RIe198a80_3114,RIfcc1148_7219,RIe195d80_3082,RIe193080_3050,RIe190380_3018,RIe18a980_2954,RIe187c80_2922,RIfcb2ee0_7058,RIe184f80_2890,RIfc615e0_6130,
        RIe182280_2858,RIe17f580_2826,RIe17c880_2794,RIfc69038_6217,RIfc4c898_5893,RIfc6f2a8_6287,RIe1764a8_2723,RIfcad0a8_6991,RIfc6adc0_6238,RIfc70388_6299,
        RIfea1b50_8184,RIfea1f88_8187,RIfc56e88_6011,RIfea1cb8_8185,RIe174450_2700,RIfc60d70_6124,RIfc6a820_6234,RIfea1e20_8186,RIf16d798_5705,RIfc40bb0_5762,
        RIe2247d8_4705,RIfc77138_6377,RIe221ad8_4673,RIfcd7d80_7478,RIe21edd8_4641,RIe2193d8_4577,RIe2166d8_4545,RIfc40070_5754,RIe2139d8_4513,RIf169850_5660,
        RIe210cd8_4481,RIfcc1580_7222,RIe20dfd8_4449,RIe20b2d8_4417,RIe2085d8_4385,RIfcd0058_7389,RIfc749d8_6349,RIe203010_4324,RIe2013f0_4304,RIfc60230_6116,
        RIfc60668_6119,RIfcaf970_7020,RIfc45818_5813,RIf160a48_5559,RIf15eb58_5537,RIfea1880_8182,RIfea19e8_8183,RIfc72110_6320,RIfc49b98_5861,RIfcca0b8_7321,
        RIfc71738_6313,RIfc4ca00_5894,RIfc71030_6308,RIfcde428_7551,RIe1fad48_4231,RIfc70bf8_6305,RIfc63a70_6156,RIfca7db0_6932,RIe1f62c0_4178,RIfcada80_6998,
        RIfc6fde8_6295,RIfc6f578_6289,RIe1f3f98_4153,RIfcde158_7549,RIfcad378_6993,RIfc65f00_6182,RIe1eeca0_4094,RIe1ec540_4066,RIe1e9840_4034,RIe1e6b40_4002,
        RIe1e3e40_3970,RIe1e1140_3938,RIe1de440_3906,RIe1db740_3874,RIe1d8a40_3842,RIe1d3040_3778,RIe1d0340_3746,RIe1cd640_3714,RIe1ca940_3682,RIe1c7c40_3650,
        RIe1c4f40_3618,RIe1c2240_3586,RIe1bf540_3554,RIfc69308_6219,RIfccba08_7339,RIe1b9f78_3493,RIe1b7db8_3469,RIfccd628_7359,RIfc69740_6222,RIe1b5bf8_3445,
        RIe1b4578_3429,RIfccf950_7384,RIf148088_5279,RIe1b3060_3414,RIe1b1710_3396,RIfc9f818_6837,RIfcb9c90_7136,RIe1acf58_3345,RIe1ab770_3328,RIe1a9880_3306,
        RIe1a6b80_3274,RIe1a3e80_3242,RIe1a1180_3210,RIe18d680_2986,RIe179b80_2762,RIe2274d8_4737,RIe21c0d8_4609,RIe2058d8_4353,RIe1ff938_4285,RIe1f8cf0_4208,
        RIe1f1838_4125,RIe1d5d40_3810,RIe1bc840_3522,RIe1af6b8_3373,RIe171cf0_2672,R_58_102f1b78,R_59_be1fc68,R_5a_10279198,R_5b_102299e8,R_5c_101d0448,
        R_5d_f7f82f0,R_5e_be21600,R_5f_f7fa5b8,R_60_1027d530,R_61_10205ae8,R_62_10283510,R_63_f82b578,R_64_ace4e68,R_65_f8204e0,R_66_1027a0b0,
        R_67_1022dc30,R_68_102478a8,R_69_10286f78,R_6a_f7edd80,R_6b_101c3628,R_6c_f7fbe00,R_6d_f7ce9f8,R_6e_f7c8830,R_6f_101ffc68,R_70_f7d4000,
        R_71_acee958,R_72_94046c0,R_73_101ee420,R_74_102eb268,R_75_b320c50,R_76_ad80a90,R_77_1027fd48,R_78_f7ce4b8,R_79_ad77048,R_7a_102a6ae0,
        R_7b_f7e4c78,R_7c_e2a6ce0,R_7d_101e86e0,R_7e_e2a9cc8,R_7f_10292be0,R_80_b33cde8,R_81_101e2908,R_82_102e9780,R_83_f8157a0,R_84_f819358,
        R_85_ace8b70,R_86_be142b0,R_87_f81b770,R_88_b330278,R_89_f7fe9f8,R_8a_101cf488,R_8b_f8225c0,R_8c_101d4738,R_8d_101c4000,R_8e_101fe960,
        R_8f_102a0330,R_90_f7f4bd0,R_91_1023e5a8,R_92_10248da8,R_93_be2c938,R_94_f7f5458,R_95_f7c6808,R_96_be316a8,R_97_e2a0328,R_98_be2d850,
        R_99_10217db0,R_9a_f7ec340,R_9b_be23ec0,R_9c_101d4540,R_9d_f800828,R_9e_102970c8,R_9f_10221de0,R_a0_ad8d568,R_a1_be4eb58,R_a2_f7c5500,
        R_a3_ad88f30,R_a4_f82f088,R_a5_f7dcbc8,R_a6_10292940,R_a7_be138d8,R_a8_acee418,R_a9_ad84450,R_aa_be10838,R_ab_be31fd8,R_ac_acdaef0,
        R_ad_acea908,R_ae_101f8830,R_af_f7dec98,R_b0_101e2c50,R_b1_f801b30,R_b2_be16e00,R_b3_102e3cf0,R_b4_10291788);
input RIdec64b8_720,RIbc62af0_23,RIbc62a78_22,RIbc62a00_21,RIbc62988_20,RIbc62910_19,RIbc62898_18,RIbc62820_17,RIbc627a8_16,
        RIbc62730_15,RIbc626b8_14,RIbc62640_13,RIdec37b8_688,RIfc8daa0_6634,RIdec0ab8_656,RIfc56348_6003,RIdebddb8_624,RIdebb0b8_592,RIdeb83b8_560,
        RIfc98798_6757,RIdeb29b8_496,RIfcbd098_7173,RIdeafcb8_464,RIfc8dc08_6635,RIdeacb80_432,RIdea6280_400,RIde9f980_368,RIfcd6868_7463,RIfc8ded8_6637,
        RIfc7dd80_6454,RIfc56618_6005,RIde92e10_306,RIde8f300_288,RIde8b160_268,RIde86fc0_248,RIde82ad8_227,RIfc8e040_6638,RIfcd96d0_7496,RIfca1e10_6864,
        RIfcbd200_7174,RIe16c5c0_2610,RIe16a298_2585,RIe168ab0_2568,RIe1664b8_2541,RIe1637b8_2509,RIee37f00_5095,RIe160ab8_2477,RIfc8ea18_6645,RIe15ddb8_2445,
        RIe1583b8_2381,RIe1556b8_2349,RIfe9f828_8159,RIe1529b8_2317,RIfe9f990_8160,RIe14fcb8_2285,RIfcbd368_7175,RIe14cfb8_2253,RIe14a2b8_2221,RIe1475b8_2189,
        RIfc8ee50_6648,RIfc45278_5809,RIfc98360_6754,RIfca2248_6867,RIe141d20_2126,RIe13f9f8_2101,RIdf3d900_2077,RIdf3b470_2051,RIfcd6ca0_7466,RIee2ff08_5004,
        RIfc8ece8_6647,RIee2dd48_4980,RIdf36718_1996,RIdf34120_1969,RIdf31f60_1945,RIfe9f6c0_8158,RIfcb4560_7074,RIfc45db8_5817,RIfc8e1a8_6639,RIfc7d678_6449,
        RIdf2aee0_1865,RIdf28ff0_1843,RIdf26e30_1819,RIdf25378_1800,RIfcb43f8_7073,RIfc8e748_6643,RIdf23488_1778,RIfcc2c00_7238,RIdf21e08_1762,RIdf20788_1746,
        RIdf1b760_1689,RIdf1a248_1674,RIdf18088_1650,RIdf15388_1618,RIdf12688_1586,RIdf0f988_1554,RIdf0cc88_1522,RIdf09f88_1490,RIdf07288_1458,RIdf04588_1426,
        RIdefeb88_1362,RIdefbe88_1330,RIdef9188_1298,RIdef6488_1266,RIdef3788_1234,RIdef0a88_1202,RIdeedd88_1170,RIdeeb088_1138,RIfc8efb8_6649,RIfc44e40_5806,
        RIfc57860_6018,RIfca23b0_6868,RIfe9faf8_8161,RIdee3900_1053,RIdee1740_1029,RIdedf6e8_1006,RIfcbd4d0_7176,RIee22678_4850,RIfc98090_6752,RIee21598_4838,
        RIfe9fc60_8162,RIded80c8_922,RIfe9fdc8_8163,RIded3be0_873,RIded18b8_848,RIdecebb8_816,RIdecbeb8_784,RIdec91b8_752,RIdeb56b8_528,RIde99080_336,
        RIe16f2c0_2642,RIe15b0b8_2413,RIe1448b8_2157,RIdf392b0_2027,RIdf2d910_1895,RIdf1e190_1719,RIdf01888_1394,RIdee8388_1106,RIdedd0f0_979,RIde7efc8_209,
        RIe19e750_3180,RIbc625c8_12,RIbc62550_11,RIbc624d8_10,RIbc62460_9,RIbc623e8_8,RIbc62370_7,RIbc622f8_6,RIbc62280_5,RIbc62208_4,
        RIbc62190_3,RIbc62118_2,RIe19ba50_3148,RIfc479d8_5837,RIe198d50_3116,RIfe9f558_8157,RIe196050_3084,RIe193350_3052,RIe190650_3020,RIe18ac50_2956,
        RIe187f50_2924,RIfc47870_5836,RIe185250_2892,RIf142ef8_5221,RIe182550_2860,RIe17f850_2828,RIe17cb50_2796,RIfcb5208_7083,RIfcbc6c0_7166,RIe177588_2735,
        RIe176610_2724,RIf13fdc0_5186,RIfe9f3f0_8156,RIfce40f8_7617,RIfc47708_5835,RIfc47438_5833,RIfca15a0_6858,RIfc99170_6764,RIe1745b8_2701,RIfc8cc90_6624,
        RIfc556a0_5994,RIfc7ee60_6466,RIfce8e50_7672,RIfe9f288_8155,RIe224aa8_4707,RIfc55808_5995,RIe221da8_4675,RIfcb50a0_7082,RIe21f0a8_4643,RIe2196a8_4579,
        RIe2169a8_4547,RIfcbc828_7167,RIe213ca8_4515,RIfc47000_5830,RIe210fa8_4483,RIfcbc990_7168,RIe20e2a8_4451,RIe20b5a8_4419,RIe2088a8_4387,RIfc46bc8_5827,
        RIfcd6598_7461,RIe2032e0_4326,RIe2016c0_4306,RIfc98ea0_6762,RIfc7eb90_6464,RIfce0318_7573,RIfcbcaf8_7169,RIfc8cf60_6626,RIfcb4dd0_7080,RIe1fd340_4258,
        RIe1fc260_4246,RIf15cf38_5517,RIfe9f120_8154,RIfc7ea28_6463,RIfc8d0c8_6627,RIfcbcc60_7170,RIfc98bd0_6760,RIfce2d48_7603,RIe1fb018_4233,RIfc55f10_6000,
        RIfc7e8c0_6462,RIfc8d230_6628,RIe1f6590_4180,RIfce58e0_7634,RIfc468f8_5825,RIfcc2ed0_7240,RIe1f4100_4154,RIfceedf0_7740,RIfc8d398_6629,RIfc8d500_6630,
        RIe1eef70_4096,RIe1ec810_4068,RIe1e9b10_4036,RIe1e6e10_4004,RIe1e4110_3972,RIe1e1410_3940,RIe1de710_3908,RIe1dba10_3876,RIe1d8d10_3844,RIe1d3310_3780,
        RIe1d0610_3748,RIe1cd910_3716,RIe1cac10_3684,RIe1c7f10_3652,RIe1c5210_3620,RIe1c2510_3588,RIe1bf810_3556,RIf14d0b0_5336,RIfe9efb8_8153,RIe1ba248_3495,
        RIe1b8088_3471,RIfec4dd0_8360,RIfec50a0_8362,RIe1b5ec8_3447,RIe1b46e0_3430,RIfcb4998_7077,RIfcb4c68_7079,RIfec5370_8364,RIfe9ee50_8152,RIfcbcdc8_7171,
        RIfc46358_5821,RIfec5208_8363,RIfec4f38_8361,RIe1a9b50_3308,RIe1a6e50_3276,RIe1a4150_3244,RIe1a1450_3212,RIe18d950_2988,RIe179e50_2764,RIe2277a8_4739,
        RIe21c3a8_4611,RIe205ba8_4355,RIe1ffc08_4287,RIe1f8fc0_4210,RIe1f1b08_4127,RIe1d6010_3812,RIe1bcb10_3524,RIe1af988_3375,RIe171fc0_2674,RIdec6080_717,
        RIdec3380_685,RIee204b8_4826,RIdec0680_653,RIfcd70d8_7469,RIdebd980_621,RIdebac80_589,RIdeb7f80_557,RIfcbe448_7187,RIdeb2580_493,RIfcb3480_7062,
        RIdeaf880_461,RIfc43928_5791,RIdeac1a8_429,RIdea58a8_397,RIde9efa8_365,RIfcd88c0_7486,RIee1c408_4780,RIfcc77f0_7292,RIfea04d0_8168,RIde92438_303,
        RIde8ec70_286,RIde8aad0_266,RIde86930_246,RIfca31c0_6878,RIfc59a20_6042,RIfcd1de0_7410,RIfc91448_6675,RIfc97280_6742,RIe16c188_2607,RIfc97118_6741,
        RIe168948_2567,RIe166080_2538,RIe163380_2506,RIee37ac8_5092,RIe160680_2474,RIfcd1c78_7409,RIe15d980_2442,RIe157f80_2378,RIe155280_2346,RIfc3f530_5746,
        RIe152580_2314,RIee35368_5064,RIe14f880_2282,RIfc7a3d8_6413,RIe14cb80_2250,RIe149e80_2218,RIe147180_2186,RIfc42b18_5781,RIfc7a270_6412,RIfc5a560_6050,
        RIfc96b78_6737,RIfea6fb0_8216,RIe13f5c0_2098,RIdf3d4c8_2074,RIdf3b038_2048,RIfce5bb0_7636,RIee2fc38_5002,RIfc91cb8_6681,RIee2d910_4977,RIdf362e0_1993,
        RIdf33e50_1967,RIdf31c90_1943,RIdf2fda0_1921,RIfc43658_5789,RIfc59e58_6045,RIfc96fb0_6740,RIfc7ac48_6419,RIfea0368_8167,RIdf28bb8_1840,RIdf26cc8_1818,
        RIdf25210_1799,RIfc91718_6677,RIfcb3318_7061,RIfc919e8_6679,RIfc91880_6678,RIfc430b8_5785,RIdf20350_1743,RIfc7a978_6417,RIdf19e10_1671,RIdf17c50_1647,
        RIdf14f50_1615,RIdf12250_1583,RIdf0f550_1551,RIdf0c850_1519,RIdf09b50_1487,RIdf06e50_1455,RIdf04150_1423,RIdefe750_1359,RIdefba50_1327,RIdef8d50_1295,
        RIdef6050_1263,RIdef3350_1231,RIdef0650_1199,RIdeed950_1167,RIdeeac50_1135,RIfcd1b10_7408,RIfc968a8_6735,RIfc91f88_6683,RIfcdfc10_7568,RIfea99e0_8246,
        RIdee3630_1051,RIdee1308_1026,RIdedf2b0_1003,RIfcc7d90_7296,RIfcd85f0_7484,RIfce3888_7611,RIfc5a830_6052,RIdeda3f0_947,RIfea9878_8245,RIded5f08_898,
        RIded37a8_870,RIded1480_845,RIdece780_813,RIdecba80_781,RIdec8d80_749,RIdeb5280_525,RIde986a8_333,RIe16ee88_2639,RIe15ac80_2410,RIe144480_2154,
        RIdf38e78_2024,RIdf2d4d8_1892,RIdf1dd58_1716,RIdf01450_1391,RIdee7f50_1103,RIdedccb8_976,RIde7e5f0_206,RIe19e318_3177,RIe19b618_3145,RIfc8f3f0_6652,
        RIe198918_3113,RIf144b18_5241,RIe195c18_3081,RIe192f18_3049,RIe190218_3017,RIe18a818_2953,RIe187b18_2921,RIf143d08_5231,RIe184e18_2889,RIfcb3cf0_7068,
        RIe182118_2857,RIe17f418_2825,RIe17c718_2793,RIfc448a0_5802,RIf141170_5200,RIfc7c9d0_6440,RIfea0098_8165,RIfc57e00_6022,RIf13f550_5180,RIfcd6e08_7467,
        RIee3d900_5159,RIfc8f6c0_6654,RIfce0048_7571,RIfca27e8_6871,RIe1742e8_2699,RIfc7c700_6438,RIfc8f990_6656,RIfce9828_7679,RIfc583a0_6026,RIf16cdc0_5698,
        RIe224670_4704,RIf16c118_5689,RIe221970_4672,RIfc58508_6027,RIe21ec70_4640,RIe219270_4576,RIe216570_4544,RIfc3ff08_5753,RIe213870_4512,RIf1696e8_5659,
        RIe210b70_4480,RIfc58940_6030,RIe20de70_4448,RIe20b170_4416,RIe208470_4384,RIfc8fc60_6658,RIfc97820_6746,RIe202ea8_4323,RIe201288_4303,RIfcc27c8_7235,
        RIfcdfee0_7570,RIfc44198_5797,RIfc58670_6028,RIf1608e0_5558,RIf15e9f0_5536,RIfe9ff30_8164,RIe1fc0f8_4245,RIfc7be90_6432,RIf15bb88_5503,RIfcd8cf8_7489,
        RIfcd8e60_7490,RIfca2d88_6875,RIfcbdea8_7183,RIfcb3a20_7066,RIe1fabe0_4230,RIfc90098_6661,RIfc90200_6662,RIfcd20b0_7412,RIe1f6158_4177,RIfc904d0_6664,
        RIfca2ef0_6876,RIfc97550_6744,RIe1f3e30_4152,RIfc59048_6035,RIfc907a0_6666,RIfc90638_6665,RIe1eeb38_4093,RIe1ec3d8_4065,RIe1e96d8_4033,RIe1e69d8_4001,
        RIe1e3cd8_3969,RIe1e0fd8_3937,RIe1de2d8_3905,RIe1db5d8_3873,RIe1d88d8_3841,RIe1d2ed8_3777,RIe1d01d8_3745,RIe1cd4d8_3713,RIe1ca7d8_3681,RIe1c7ad8_3649,
        RIe1c4dd8_3617,RIe1c20d8_3585,RIe1bf3d8_3553,RIfcc73b8_7289,RIfce3cc0_7614,RIe1b9e10_3492,RIe1b7c50_3468,RIfcd6f70_7468,RIf149e10_5300,RIe1b5a90_3444,
        RIfea0200_8166,RIfc90bd8_6669,RIfcdfd78_7569,RIe1b2ef8_3413,RIe1b15a8_3395,RIfc973e8_6743,RIfcc7520_7290,RIe1acdf0_3344,RIe1ab608_3327,RIe1a9718_3305,
        RIe1a6a18_3273,RIe1a3d18_3241,RIe1a1018_3209,RIe18d518_2985,RIe179a18_2761,RIe227370_4736,RIe21bf70_4608,RIe205770_4352,RIe1ff7d0_4284,RIe1f8b88_4207,
        RIe1f16d0_4124,RIe1d5bd8_3809,RIe1bc6d8_3521,RIe1af550_3372,RIe171b88_2671,RIdec5108_706,RIdec2408_674,RIfc93608_6699,RIdebf708_642,RIfc934a0_6698,
        RIdebca08_610,RIdeb9d08_578,RIdeb7008_546,RIfcdf7d8_7565,RIdeb1608_482,RIfc78218_6389,RIdeae908_450,RIfcc8498_7301,RIdea9d90_418,RIdea3490_386,
        RIde9cb90_354,RIee1cc78_4786,RIee1bb98_4774,RIee1b328_4768,RIee1aab8_4762,RIde909f8_295,RIde8d578_279,RIfea8ea0_8238,RIde85238_239,RIde813e0_220,
        RIfc938d8_6701,RIfce5e80_7638,RIfcbfd98_7205,RIfce8ce8_7671,RIe16b4e0_2598,RIfea8d38_8237,RIfea9f80_8250,RIe165108_2527,RIe162408_2495,RIfc779a8_6383,
        RIe15f708_2463,RIfe9dc08_8139,RIe15ca08_2431,RIe157008_2367,RIe154308_2335,RIfea7550_8220,RIe151608_2303,RIfcd6160_7458,RIe14e908_2271,RIfcd1408_7403,
        RIe14bc08_2239,RIe148f08_2207,RIe146208_2175,RIfceb718_7701,RIfcb19c8_7043,RIfc93e78_6705,RIfce7938_7657,RIe140da8_2115,RIdf3ecb0_2091,RIdf3c988_2066,
        RIfe9daa0_8138,RIfce8478_7665,RIfcdbf98_7525,RIfc776d8_6381,RIfc93fe0_6706,RIdf354d0_1983,RIdf33040_1957,RIdf30fe8_1934,RIdf2ee28_1910,RIee2ba20_4955,
        RIfc93ba8_6703,RIfc77de0_6386,RIee27ad8_4910,RIfe9d668_8135,RIfea8bd0_8236,RIdf26458_1812,RIfe9d7d0_8136,RIfcb1c98_7045,RIee26cc8_4900,RIdf22ab0_1771,
        RIfcc0068_7207,RIdf21598_1756,RIdf1f6a8_1734,RIdf1aef0_1683,RIfe9d938_8137,RIdf16cd8_1636,RIdf13fd8_1604,RIdf112d8_1572,RIdf0e5d8_1540,RIdf0b8d8_1508,
        RIdf08bd8_1476,RIdf05ed8_1444,RIdf031d8_1412,RIdefd7d8_1348,RIdefaad8_1316,RIdef7dd8_1284,RIdef50d8_1252,RIdef23d8_1220,RIdeef6d8_1188,RIdeec9d8_1156,
        RIdee9cd8_1124,RIfc942b0_6708,RIfcde6f8_7553,RIfcd1138_7401,RIfcde860_7554,RIdee4878_1064,RIdee2af0_1043,RIdee0a98_1020,RIdede8d8_996,RIfc5c9f0_6076,
        RIee22240_4847,RIfcc8768_7303,RIee21160_4835,RIded95e0_937,RIded7150_911,RIded5260_889,RIfea76b8_8221,RIded0508_834,RIdecd808_802,RIdecab08_770,
        RIdec7e08_738,RIdeb4308_514,RIde96290_322,RIe16df10_2628,RIe159d08_2399,RIe143508_2143,RIdf37f00_2013,RIdf2c560_1881,RIdf1cde0_1705,RIdf004d8_1380,
        RIdee6fd8_1092,RIdedbd40_965,RIde7c1d8_195,RIe19d3a0_3166,RIe19a6a0_3134,RIfcb2c10_7056,RIe1979a0_3102,RIfc923c0_6686,RIe194ca0_3070,RIe191fa0_3038,
        RIe18f2a0_3006,RIe1898a0_2942,RIe186ba0_2910,RIfc422a8_5775,RIe183ea0_2878,RIfcbecb8_7193,RIe1811a0_2846,RIe17e4a0_2814,RIe17b7a0_2782,RIf142250_5212,
        RIf140bd0_5196,RIfec43f8_8353,RIe175968_2715,RIfc79b68_6407,RIf13efb0_5176,RIfc92528_6687,RIfcb2aa8_7055,RIfcd8320_7482,RIfcea200_7686,RIfc79898_6405,
        RIe1734d8_2689,RIfcd7948_7475,RIfcd7678_7473,RIf16e170_5712,RIfc927f8_6689,RIfc92960_6690,RIe2236f8_4693,RIfc795c8_6403,RIe2209f8_4661,RIf16ad68_5675,
        RIe21dcf8_4629,RIe2182f8_4565,RIe2155f8_4533,RIfe9d398_8133,RIe2128f8_4501,RIfcdb9f8_7521,RIe20fbf8_4469,RIfc41d08_5771,RIe20cef8_4437,RIe20a1f8_4405,
        RIe2074f8_4373,RIfcd7510_7472,RIf166010_5620,RIfe9d230_8132,RIe2008b0_4296,RIf165098_5609,RIfc41ba0_5770,RIfc41a38_5769,RIfc92c30_6692,RIfc418d0_5768,
        RIfc79190_6400,RIe1fcad0_4252,RIfec4560_8354,RIfc79028_6399,RIfcbf258_7197,RIfcc1df0_7228,RIfcd81b8_7481,RIfc92d98_6693,RIfc5b4d8_6061,RIfcd77e0_7474,
        RIe1fa0a0_4222,RIf156188_5439,RIfe9d500_8134,RIf1546d0_5420,RIe1f5348_4167,RIfec4830_8356,RIfec46c8_8355,RIf1508f0_5376,RIe1f3020_4142,RIfce3180_7606,
        RIfce8fb8_7673,RIfcbf690_7200,RIe1edd28_4083,RIe1eb460_4054,RIe1e8760_4022,RIe1e5a60_3990,RIe1e2d60_3958,RIe1e0060_3926,RIe1dd360_3894,RIe1da660_3862,
        RIe1d7960_3830,RIe1d1f60_3766,RIe1cf260_3734,RIe1cc560_3702,RIe1c9860_3670,RIe1c6b60_3638,RIe1c3e60_3606,RIe1c1160_3574,RIe1be460_3542,RIfe9d0c8_8131,
        RIfe9cc90_8128,RIe1b9168_3483,RIe1b7110_3460,RIf14a3b0_5304,RIfe9cb28_8127,RIfe9cf60_8130,RIfe9c9c0_8126,RIfce2208_7595,RIfce9558_7677,RIfe9c858_8125,
        RIfe9cdf8_8129,RIf147110_5268,RIf146468_5259,RIe1ac2b0_3336,RIe1aaac8_3319,RIe1a87a0_3294,RIe1a5aa0_3262,RIe1a2da0_3230,RIe1a00a0_3198,RIe18c5a0_2974,
        RIe178aa0_2750,RIe2263f8_4725,RIe21aff8_4597,RIe2047f8_4341,RIe1fe858_4273,RIe1f7c10_4196,RIe1f0758_4113,RIe1d4c60_3798,RIe1bb760_3510,RIe1ae5d8_3361,
        RIe170c10_2660,RIdec4190_695,RIdec1490_663,RIfceaa70_7692,RIdebe790_631,RIfc954f8_6721,RIdebba90_599,RIdeb8d90_567,RIdeb6090_535,RIfcebb50_7704,
        RIdeb0690_471,RIee1e190_4801,RIdead990_439,RIfcdf0d0_7560,RIdea7978_407,RIdea1078_375,RIde9a778_343,RIee1c840_4783,RIfc957c8_6723,RIfcc8e70_7308,
        RIfc5e610_6096,RIfe9e8b0_8148,RIde8c1c8_273,RIde88028_253,RIde83b40_232,RIfcb0bb8_7033,RIfca4b10_6896,RIfc75d88_6363,RIfca4c78_6897,RIfc95390_6720,
        RIe16a9a0_2590,RIfcc8fd8_7309,RIe166e90_2548,RIe164190_2516,RIe161490_2484,RIfe9e748_8147,RIe15e790_2452,RIfc74f78_6353,RIe15ba90_2420,RIe156090_2356,
        RIe153390_2324,RIfc3ecc0_5740,RIe150690_2292,RIfce8b80_7670,RIe14d990_2260,RIfca6730_6916,RIe14ac90_2228,RIe147f90_2196,RIe145290_2164,RIfcee2b0_7732,
        RIfc5f2b8_6105,RIfc753b0_6356,RIfc74b40_6350,RIe140268_2107,RIdf3e170_2083,RIdf3be48_2058,RIdf39c88_2034,RIfcc1c88_7227,RIfcc1850_7224,RIfc965d8_6733,
        RIfc96038_6729,RIdf34828_1974,RIdf327d0_1951,RIdf301d8_1924,RIdf2e2e8_1902,RIfc5e778_6097,RIfcd0328_7391,RIfc757e8_6359,RIfcee6e8_7735,RIdf296f8_1848,
        RIdf273d0_1823,RIdf257b0_1803,RIdf23b90_1783,RIfc95d68_6727,RIfceda40_7726,RIfe9eb80_8150,RIfc75518_6357,RIfcd01c0_7390,RIdf1eb68_1726,RIfe9ece8_8151,
        RIfe9ea18_8149,RIdf15d60_1625,RIdf13060_1593,RIdf10360_1561,RIdf0d660_1529,RIdf0a960_1497,RIdf07c60_1465,RIdf04f60_1433,RIdf02260_1401,RIdefc860_1337,
        RIdef9b60_1305,RIdef6e60_1273,RIdef4160_1241,RIdef1460_1209,RIdeee760_1177,RIdeeba60_1145,RIdee8d60_1113,RIfc961a0_6730,RIfc96308_6731,RIfc5ee80_6102,
        RIfce6150_7640,RIdee42d8_1060,RIdee1e48_1034,RIdee00c0_1013,RIdeddac8_986,RIfc96470_6732,RIfc75248_6355,RIfc74ca8_6351,RIfcb0618_7029,RIded8938_928,
        RIded6610_903,RIded4450_879,RIded2290_855,RIdecf590_823,RIdecc890_791,RIdec9b90_759,RIdec6e90_727,RIdeb3390_503,RIde93e78_311,RIe16cf98_2617,
        RIe158d90_2388,RIe142590_2132,RIdf36f88_2002,RIdf2b5e8_1870,RIdf1be68_1694,RIdeff560_1369,RIdee6060_1081,RIdedadc8_954,RIde79dc0_184,RIe19c428_3155,
        RIe199728_3123,RIfe9e310_8144,RIe196a28_3091,RIfcc04a0_7210,RIe193d28_3059,RIe191028_3027,RIe18e328_2995,RIe188928_2931,RIe185c28_2899,RIfce1830_7588,
        RIe182f28_2867,RIfe9e478_8145,RIe180228_2835,RIe17d528_2803,RIe17a828_2771,RIf141878_5205,RIfcb12c0_7038,RIfc94418_6709,RIe174f90_2708,RIfc77408_6379,
        RIf13ea10_5172,RIfcdc100_7526,RIfc94580_6710,RIfc946e8_6711,RIfced338_7721,RIfce5fe8_7639,RIe172998_2681,RIfcdc268_7527,RIfcddff0_7548,RIfcc0608_7211,
        RIfce7230_7652,RIfc40340_5756,RIe222780_4682,RIfcdd618_7541,RIe21fa80_4650,RIfcd0b98_7397,RIe21cd80_4618,RIe217380_4554,RIe214680_4522,RIfec4998_8357,
        RIe211980_4490,RIf168608_5647,RIe20ec80_4458,RIfcc0770_7212,RIe20bf80_4426,RIe209280_4394,RIe206580_4362,RIfce2370_7596,RIfcee580_7734,RIfec4c68_8359,
        RIfec4b00_8358,RIfc949b8_6713,RIfcebcb8_7705,RIf162938_5581,RIf1612b8_5565,RIfccd088_7355,RIfcc08d8_7213,RIfe9e040_8142,RIfe9e1a8_8143,RIfcead40_7694,
        RIf15ad78_5493,RIfc94c88_6715,RIfccc3e0_7346,RIfc765f8_6369,RIfc94df0_6716,RIfcc0a40_7214,RIe1f9998_4217,RIfcc8d08_7307,RIfce8748_7667,RIfceb2e0_7698,
        RIe1f4970_4160,RIf152510_5396,RIf1512c8_5383,RIfcb0ff0_7036,RIe1f24e0_4134,RIfc761c0_6366,RIfc950c0_6718,RIfcc0e78_7217,RIe1ed1e8_4075,RIe1ea4e8_4043,
        RIe1e77e8_4011,RIe1e4ae8_3979,RIe1e1de8_3947,RIe1df0e8_3915,RIe1dc3e8_3883,RIe1d96e8_3851,RIe1d69e8_3819,RIe1d0fe8_3755,RIe1ce2e8_3723,RIe1cb5e8_3691,
        RIe1c88e8_3659,RIe1c5be8_3627,RIe1c2ee8_3595,RIe1c01e8_3563,RIe1bd4e8_3531,RIf14bfd0_5324,RIf14ac20_5310,RIfe9ded8_8141,RIe1b65d0_3452,RIfcecd98_7717,
        RIfc76490_6368,RIe1b4c80_3434,RIe1b38d0_3420,RIfcc0fe0_7218,RIfceaea8_7695,RIe1b1f80_3402,RIe1b0360_3382,RIfcd0760_7394,RIf145ec8_5255,RIfe9e5e0_8146,
        RIfe9dd70_8140,RIe1a7828_3283,RIe1a4b28_3251,RIe1a1e28_3219,RIe19f128_3187,RIe18b628_2963,RIe177b28_2739,RIe225480_4714,RIe21a080_4586,RIe203880_4330,
        RIe1fd8e0_4262,RIe1f6c98_4185,RIe1ef7e0_4102,RIe1d3ce8_3787,RIe1ba7e8_3499,RIe1ad660_3350,RIe16fc98_2649,RIdec6788_722,RIdec3a88_690,RIee20788_4828,
        RIdec0d88_658,RIee1f810_4817,RIdebe088_626,RIdebb388_594,RIdeb8688_562,RIfc9b1c8_6787,RIdeb2c88_498,RIfce1f38_7593,RIdeaff88_466,RIfc892e8_6583,
        RIdead210_434,RIdea6910_402,RIdea0010_370,RIee1d650_4793,RIee1c570_4781,RIee1b5f8_4770,RIee1aef0_4765,RIfe99888_8091,RIfe99450_8088,RIfe99720_8090,
        RIfe995b8_8089,RIde83168_229,RIfcc43e8_7255,RIfcd5a58_7453,RIfc89450_6584,RIfcc5798_7269,RIe16c890_2612,RIe16a568_2587,RIe168d80_2570,RIe166788_2543,
        RIe163a88_2511,RIfc83618_6517,RIe160d88_2479,RIee36718_5078,RIe15e088_2447,RIe158688_2383,RIe155988_2351,RIfc3f800_5748,RIe152c88_2319,RIfc895b8_6585,
        RIe14ff88_2287,RIfc51cf8_5953,RIe14d288_2255,RIe14a588_2223,RIe147888_2191,RIee34990_5057,RIee338b0_5045,RIfc831e0_6514,RIfcd3b68_7431,RIe141ff0_2128,
        RIe13fcc8_2103,RIdf3dbd0_2079,RIdf3b740_2053,RIfcb6f90_7104,RIee301d8_5006,RIfcba938_7145,RIee2e018_4982,RIdf369e8_1998,RIdf343f0_1971,RIdf32230_1947,
        RIfe99e28_8095,RIfc83078_6513,RIfcb6e28_7103,RIfc9ad90_6784,RIfcbad70_7148,RIdf2b1b0_1867,RIdf292c0_1845,RIfe99b58_8093,RIfe999f0_8092,RIfc9ac28_6783,
        RIfc4a9a8_5871,RIdf23758_1780,RIfc82da8_6511,RIdf220d8_1764,RIdf20a58_1748,RIdf1ba30_1691,RIfe99cc0_8094,RIdf18358_1652,RIdf15658_1620,RIdf12958_1588,
        RIdf0fc58_1556,RIdf0cf58_1524,RIdf0a258_1492,RIdf07558_1460,RIdf04858_1428,RIdefee58_1364,RIdefc158_1332,RIdef9458_1300,RIdef6758_1268,RIdef3a58_1236,
        RIdef0d58_1204,RIdeee058_1172,RIdeeb358_1140,RIee25918_4886,RIee24b08_4876,RIfc52568_5959,RIfc826a0_6506,RIdee5958_1076,RIdee3bd0_1055,RIfe99f90_8096,
        RIdedf9b8_1008,RIfce4800_7622,RIfc89b58_6589,RIfc9f3e0_6834,RIfc82538_6505,RIdeda828_950,RIded8398_924,RIfeabe70_8272,RIded3eb0_875,RIded1b88_850,
        RIdecee88_818,RIdecc188_786,RIdec9488_754,RIdeb5988_530,RIde99710_338,RIe16f590_2644,RIe15b388_2415,RIe144b88_2159,RIdf39580_2029,RIdf2dbe0_1897,
        RIdf1e460_1721,RIdf01b58_1396,RIdee8658_1108,RIdedd3c0_981,RIde7f658_211,RIe19ea20_3182,RIe19bd20_3150,RIf145928_5251,RIe199020_3118,RIfe98910_8080,
        RIe196320_3086,RIe193620_3054,RIe190920_3022,RIe18af20_2958,RIe188220_2926,RIf143e70_5232,RIe185520_2894,RIfc95c00_6726,RIe182820_2862,RIe17fb20_2830,
        RIe17ce20_2798,RIf142520_5214,RIf141440_5202,RIe1776f0_2736,RIfeab8d0_8268,RIfcc5bd0_7272,RIfc62dc8_6147,RIee3e710_5169,RIfc9cb18_6805,RIee3c820_5147,
        RIee3b470_5133,RIee3a390_5121,RIe174888_2703,RIf170498_5737,RIfc68660_6210,RIf16e878_5717,RIfc6ea38_6281,RIfe98d48_8083,RIe224d78_4709,RIf16c280_5690,
        RIe222078_4677,RIf16b308_5679,RIe21f378_4645,RIe219978_4581,RIe216c78_4549,RIf16a390_5668,RIe213f78_4517,RIf169b20_5662,RIe211278_4485,RIf1681d0_5644,
        RIe20e578_4453,RIe20b878_4421,RIe208b78_4389,RIfcd4ae0_7442,RIfc61478_6129,RIfeab060_8262,RIe201990_4308,RIfc70ec8_6307,RIfc70928_6303,RIfcec528_7711,
        RIfcbe880_7190,RIf160d18_5561,RIf15ee28_5539,RIfe98be0_8082,RIfe98eb0_8084,RIf15d0a0_5518,RIf15bcf0_5504,RIfcd4540_7438,RIf159e00_5482,RIf1592c0_5474,
        RIf158078_5461,RIfca3a30_6884,RIfea7988_8223,RIf156728_5443,RIf155be8_5435,RIf154b08_5423,RIfe98a78_8081,RIf1538c0_5410,RIf1520d8_5393,RIf150e90_5380,
        RIe1f43d0_4156,RIf14fdb0_5368,RIfcd2380_7414,RIf14e2f8_5349,RIe1ef240_4098,RIe1ecae0_4070,RIe1e9de0_4038,RIe1e70e0_4006,RIe1e43e0_3974,RIe1e16e0_3942,
        RIe1de9e0_3910,RIe1dbce0_3878,RIe1d8fe0_3846,RIe1d35e0_3782,RIe1d08e0_3750,RIe1cdbe0_3718,RIe1caee0_3686,RIe1c81e0_3654,RIe1c54e0_3622,RIe1c27e0_3590,
        RIe1bfae0_3558,RIfc44b70_5804,RIf14bd00_5322,RIfe992e8_8087,RIfe987a8_8079,RIf14a950_5308,RIf149f78_5301,RIfe99180_8086,RIfe98640_8078,RIf149438_5293,
        RIfcec7f8_7713,RIfe984d8_8077,RIe1b1b48_3399,RIfc4b650_5880,RIfcda918_7509,RIfe98370_8076,RIfe99018_8085,RIe1a9e20_3310,RIe1a7120_3278,RIe1a4420_3246,
        RIe1a1720_3214,RIe18dc20_2990,RIe17a120_2766,RIe227a78_4741,RIe21c678_4613,RIe205e78_4357,RIe1ffed8_4289,RIe1f9290_4212,RIe1f1dd8_4129,RIe1d62e0_3814,
        RIe1bcde0_3526,RIe1afc58_3377,RIe172290_2676,RIdec6620_721,RIdec3920_689,RIfc49328_5855,RIdec0c20_657,RIfc80eb8_6489,RIdebdf20_625,RIdebb220_593,
        RIdeb8520_561,RIfc80648_6483,RIdeb2b20_497,RIfc8b340_6606,RIdeafe20_465,RIfc491c0_5854,RIdeacec8_433,RIdea65c8_401,RIde9fcc8_369,RIfcd9c70_7500,
        RIfe98208_8075,RIfce4698_7621,RIfe980a0_8074,RIde93158_307,RIde8f648_289,RIde8b4a8_269,RIde87308_249,RIde82e20_228,RIfcbba18_7157,RIfc48d88_5851,
        RIfc99f80_6774,RIfc8b4a8_6607,RIe16c728_2611,RIe16a400_2586,RIe168c18_2569,RIe166620_2542,RIe163920_2510,RIee38068_5096,RIe160c20_2478,RIfc48248_5843,
        RIe15df20_2446,RIe158520_2382,RIe155820_2350,RIfcbbe50_7160,RIe152b20_2318,RIfc47e10_5840,RIe14fe20_2286,RIfca0e98_6853,RIe14d120_2254,RIe14a420_2222,
        RIe147720_2190,RIfc8be80_6614,RIfc7fb08_6475,RIfc480e0_5842,RIfc99878_6769,RIe141e88_2127,RIe13fb60_2102,RIdf3da68_2078,RIdf3b5d8_2052,RIfe97f38_8073,
        RIee30070_5005,RIee2eb58_4990,RIee2deb0_4981,RIdf36880_1997,RIdf34288_1970,RIdf320c8_1946,RIfe97dd0_8072,RIfcc3740_7246,RIfc48ab8_5849,RIfce05e8_7575,
        RIfc80210_6480,RIdf2b048_1866,RIdf29158_1844,RIdf26f98_1820,RIdf254e0_1801,RIfc8bbb0_6612,RIfc48950_5848,RIdf235f0_1779,RIfc8bd18_6613,RIdf21f70_1763,
        RIdf208f0_1747,RIdf1b8c8_1690,RIdf1a3b0_1675,RIdf181f0_1651,RIdf154f0_1619,RIdf127f0_1587,RIdf0faf0_1555,RIdf0cdf0_1523,RIdf0a0f0_1491,RIdf073f0_1459,
        RIdf046f0_1427,RIdefecf0_1363,RIdefbff0_1331,RIdef92f0_1299,RIdef65f0_1267,RIdef38f0_1235,RIdef0bf0_1203,RIdeedef0_1171,RIdeeb1f0_1139,RIfcbc120_7162,
        RIfcd9838_7497,RIfc99710_6768,RIfca1168_6855,RIdee57f0_1075,RIdee3a68_1054,RIdee18a8_1030,RIdedf850_1007,RIfc549f8_5985,RIfcb5370_7084,RIfce43c8_7619,
        RIfce0480_7574,RIdeda6c0_949,RIded8230_923,RIded6070_899,RIded3d48_874,RIded1a20_849,RIdeced20_817,RIdecc020_785,RIdec9320_753,RIdeb5820_529,
        RIde993c8_337,RIe16f428_2643,RIe15b220_2414,RIe144a20_2158,RIdf39418_2028,RIdf2da78_1896,RIdf1e2f8_1720,RIdf019f0_1395,RIdee84f0_1107,RIdedd258_980,
        RIde7f310_210,RIe19e8b8_3181,RIe19bbb8_3149,RIfe976c8_8067,RIe198eb8_3117,RIf144c80_5242,RIe1961b8_3085,RIe1934b8_3053,RIe1907b8_3021,RIe18adb8_2957,
        RIe1880b8_2925,RIfe97560_8066,RIe1853b8_2893,RIfcc3fb0_7252,RIe1826b8_2861,RIe17f9b8_2829,RIe17ccb8_2797,RIfcd3730_7428,RIf1412d8_5201,RIfcc4118_7253,
        RIfe97830_8068,RIfc4a6d8_5869,RIf13f6b8_5181,RIfc9f980_6838,RIfc9fae8_6839,RIfcc3e48_7251,RIfc89e28_6591,RIfc89cc0_6590,RIe174720_2702,RIfc4a408_5867,
        RIfce27a8_7599,RIfc530a8_5967,RIfcd5d28_7455,RIf16cf28_5699,RIe224c10_4708,RIfc53210_5968,RIe221f10_4676,RIf16b1a0_5678,RIe21f210_4644,RIe219810_4580,
        RIe216b10_4548,RIfc401d8_5755,RIe213e10_4516,RIf1699b8_5661,RIe211110_4484,RIfc81cc8_6499,RIe20e410_4452,RIe20b710_4420,RIe208a10_4388,RIfc8a0f8_6593,
        RIfcb6720_7098,RIe203448_4327,RIe201828_4307,RIfc53378_5969,RIfc8a3c8_6595,RIfcb65b8_7097,RIfc49fd0_5864,RIf160bb0_5560,RIf15ecc0_5538,RIe1fd4a8_4259,
        RIfe97b00_8070,RIfc8a530_6596,RIfe97c68_8071,RIfc8a800_6598,RIfc8a698_6597,RIfc9a7f0_6780,RIfc81890_6496,RIfcd5e90_7456,RIe1fb180_4234,RIfc49e68_5863,
        RIfc81728_6495,RIfcbb1a8_7151,RIe1f66f8_4181,RIfcd3460_7426,RIfcb62e8_7095,RIfc9a520_6778,RIe1f4268_4155,RIfc49d00_5862,RIfcd9dd8_7501,RIfcbb310_7152,
        RIe1ef0d8_4097,RIe1ec978_4069,RIe1e9c78_4037,RIe1e6f78_4005,RIe1e4278_3973,RIe1e1578_3941,RIe1de878_3909,RIe1dbb78_3877,RIe1d8e78_3845,RIe1d3478_3781,
        RIe1d0778_3749,RIe1cda78_3717,RIe1cad78_3685,RIe1c8078_3653,RIe1c5378_3621,RIe1c2678_3589,RIe1bf978_3557,RIfc49a30_5860,RIfcb6018_7093,RIe1ba3b0_3496,
        RIe1b81f0_3472,RIfce0a20_7578,RIfcbb5e0_7154,RIe1b6030_3448,RIfe97998_8069,RIfce5610_7632,RIfcc3a10_7248,RIe1b3330_3416,RIe1b19e0_3398,RIfc495f8_5857,
        RIfc81188_6491,RIe1ad228_3347,RIe1aba40_3330,RIe1a9cb8_3309,RIe1a6fb8_3277,RIe1a42b8_3245,RIe1a15b8_3213,RIe18dab8_2989,RIe179fb8_2765,RIe227910_4740,
        RIe21c510_4612,RIe205d10_4356,RIe1ffd70_4288,RIe1f9128_4211,RIe1f1c70_4128,RIe1d6178_3813,RIe1bcc78_3525,RIe1afaf0_3376,RIe172128_2675,RIdec6a58_724,
        RIdec3d58_692,RIfc723e0_6322,RIdec1058_660,RIfc59fc0_6046,RIdebe358_628,RIdebb658_596,RIdeb8958_564,RIfcb96f0_7132,RIdeb2f58_500,RIfce1c68_7591,
        RIdeb0258_468,RIfc9b498_6789,RIdead558_436,RIdea6fa0_404,RIdea06a0_372,RIfc81458_6493,RIfc83780_6518,RIfc4e620_5914,RIfcd3e38_7433,RIde937e8_309,
        RIde8f990_290,RIde8bb38_271,RIde87650_250,RIde834b0_230,RIfc42c80_5782,RIfc65960_6178,RIfc6c710_6256,RIee392b0_5109,RIe16cb60_2614,RIe16a6d0_2588,
        RIe169050_2572,RIe166a58_2545,RIe163d58_2513,RIfec3cf0_8348,RIe161058_2481,RIfcd54b8_7449,RIe15e358_2449,RIe158958_2385,RIe155c58_2353,RIfe9ba48_8115,
        RIe152f58_2321,RIfec4128_8351,RIe150258_2289,RIfcb9b28_7135,RIe14d558_2257,RIe14a858_2225,RIe147b58_2193,RIfcdb2f0_7516,RIfc553d0_5992,RIfc9a0e8_6775,
        RIfcbd908_7179,RIe1422c0_2130,RIe13ff98_2105,RIdf3dea0_2081,RIdf3ba10_2055,RIfc87128_6559,RIee304a8_5008,RIfcc51f8_7265,RIee2e2e8_4984,RIdf36cb8_2000,
        RIfec3fc0_8350,RIdf32500_1949,RIfec3e58_8349,RIee2c830_4965,RIee2ad78_4946,RIee296f8_4930,RIee284b0_4917,RIfe9b8e0_8114,RIfe9b610_8112,RIfe9b778_8113,
        RIfe9b4a8_8111,RIfcb7c38_7113,RIfc86b88_6555,RIdf238c0_1781,RIfc75ab8_6361,RIdf22240_1765,RIfeaa3b8_8253,RIdf1bb98_1692,RIdf1a680_1677,RIdf18628_1654,
        RIdf15928_1622,RIdf12c28_1590,RIdf0ff28_1558,RIdf0d228_1526,RIdf0a528_1494,RIdf07828_1462,RIdf04b28_1430,RIdeff128_1366,RIdefc428_1334,RIdef9728_1302,
        RIdef6a28_1270,RIdef3d28_1238,RIdef1028_1206,RIdeee328_1174,RIdeeb628_1142,RIee25a80_4887,RIee24c70_4877,RIfcddd20_7546,RIfccc110_7344,RIdee5c28_1078,
        RIdee3ea0_1057,RIdee1b78_1032,RIdedfc88_1010,RIfc6a6b8_6233,RIee227e0_4851,RIfc88be0_6578,RIee21868_4840,RIdedaaf8_952,RIded8668_926,RIded6340_901,
        RIded4180_877,RIded1e58_852,RIdecf158_820,RIdecc458_788,RIdec9758_756,RIdeb5c58_532,RIde99da0_340,RIe16f860_2646,RIe15b658_2417,RIe144e58_2161,
        RIdf39850_2031,RIdf2deb0_1899,RIdf1e730_1723,RIdf01e28_1398,RIdee8928_1110,RIdedd690_983,RIde7fce8_213,RIe19ecf0_3184,RIe19bff0_3152,RIf145a90_5252,
        RIe1992f0_3120,RIf144de8_5243,RIe1965f0_3088,RIe1938f0_3056,RIe190bf0_3024,RIe18b1f0_2960,RIe1884f0_2928,RIfc72980_6326,RIe1857f0_2896,RIf143060_5222,
        RIe182af0_2864,RIe17fdf0_2832,RIe17d0f0_2800,RIf142688_5215,RIf141710_5204,RIe177858_2737,RIe176778_2725,RIfcea638_7689,RIfca54e8_6903,RIee3e878_5170,
        RIee3dbd0_5161,RIee3c988_5148,RIee3b5d8_5134,RIee3a4f8_5122,RIe174b58_2705,RIf170600_5738,RIfc76fd0_6376,RIf16e9e0_5718,RIfced608_7723,RIf16d090_5700,
        RIe225048_4711,RIf16c550_5692,RIe222348_4679,RIf16b470_5680,RIe21f648_4647,RIe219c48_4583,RIe216f48_4551,RIf16a4f8_5669,RIe214248_4519,RIf169df0_5664,
        RIe211548_4487,RIf1684a0_5646,RIe20e848_4455,RIe20bb48_4423,RIe208e48_4391,RIf1673c0_5634,RIf166448_5623,RIfe9c6f0_8124,RIfe9c150_8120,RIf1654d0_5612,
        RIfcc4550_7256,RIf1635e0_5590,RIf162500_5578,RIf160fe8_5563,RIf15f0f8_5541,RIfe9bfe8_8119,RIfe9c588_8123,RIf15d208_5519,RIf15bfc0_5506,RIfc4d540_5902,
        RIfc9c848_6803,RIfec4290_8352,RIfe9c2b8_8121,RIfcc01d0_7208,RIe1fb2e8_4235,RIfe9c420_8122,RIfca3e68_6887,RIf154c70_5424,RIe1f69c8_4183,RIf153a28_5411,
        RIf152240_5394,RIf150ff8_5381,RIe1f46a0_4158,RIfca6028_6911,RIfc43bf8_5793,RIf14e460_5350,RIe1ef3a8_4099,RIe1ecdb0_4072,RIe1ea0b0_4040,RIe1e73b0_4008,
        RIe1e46b0_3976,RIe1e19b0_3944,RIe1decb0_3912,RIe1dbfb0_3880,RIe1d92b0_3848,RIe1d38b0_3784,RIe1d0bb0_3752,RIe1cdeb0_3720,RIe1cb1b0_3688,RIe1c84b0_3656,
        RIe1c57b0_3624,RIe1c2ab0_3592,RIe1bfdb0_3560,RIfc4d6a8_5903,RIf14be68_5323,RIe1ba680_3498,RIfe9be80_8118,RIfc86e58_6557,RIfcd46a8_7439,RIe1b6300_3450,
        RIfe9bd18_8117,RIf1495a0_5294,RIf1481f0_5280,RIe1b3600_3418,RIe1b1e18_3401,RIfc69470_6220,RIfcbfac8_7203,RIfe9bbb0_8116,RIe1abd10_3332,RIe1aa0f0_3312,
        RIe1a73f0_3280,RIe1a46f0_3248,RIe1a19f0_3216,RIe18def0_2992,RIe17a3f0_2768,RIe227d48_4743,RIe21c948_4615,RIe206148_4359,RIe2001a8_4291,RIe1f9560_4214,
        RIe1f20a8_4131,RIe1d65b0_3816,RIe1bd0b0_3528,RIe1aff28_3379,RIe172560_2678,RIdec68f0_723,RIdec3bf0_691,RIee208f0_4829,RIdec0ef0_659,RIfc7ce08_6443,
        RIdebe1f0_627,RIdebb4f0_595,RIdeb87f0_563,RIfc9b8d0_6792,RIdeb2df0_499,RIfcc6710_7280,RIdeb00f0_467,RIfc5ff60_6114,RIdead3f0_435,RIdea6c58_403,
        RIdea0358_371,RIfce5070_7628,RIee1c6d8_4782,RIfce70c8_7651,RIee1b058_4766,RIde934a0_308,RIfe9b1d8_8109,RIde8b7f0_270,RIfe9b340_8110,RIfc6b798_6245,
        RIfcb2238_7049,RIfcd3a00_7430,RIfcdb020_7514,RIfc511b8_5945,RIe16c9f8_2613,RIfcb27d8_7053,RIe168ee8_2571,RIe1668f0_2544,RIe163bf0_2512,RIee381d0_5097,
        RIe160ef0_2480,RIfcdfaa8_7567,RIe15e1f0_2448,RIe1587f0_2384,RIe155af0_2352,RIfc3f968_5749,RIe152df0_2320,RIfcd5080_7446,RIe1500f0_2288,RIfc84b30_6532,
        RIe14d3f0_2256,RIe14a6f0_2224,RIe1479f0_2192,RIfcea098_7685,RIfc92f00_6694,RIfc54890_5984,RIfcdcc40_7534,RIe142158_2129,RIe13fe30_2104,RIdf3dd38_2080,
        RIdf3b8a8_2054,RIfc57590_6016,RIee30340_5007,RIfcd0490_7392,RIee2e180_4983,RIdf36b50_1999,RIdf34558_1972,RIdf32398_1948,RIfe9b070_8108,RIfcb1860_7042,
        RIfca1b40_6862,RIfc5c018_6069,RIfe9ada0_8106,RIdf2b318_1868,RIdf29428_1846,RIdf27100_1821,RIfe9af08_8107,RIfc5e1d8_6093,RIfcdcda8_7535,RIfcac400_6982,
        RIfc691a0_6218,RIfcaad80_6966,RIdf20bc0_1749,RIfc61b80_6134,RIdf1a518_1676,RIdf184c0_1653,RIdf157c0_1621,RIdf12ac0_1589,RIdf0fdc0_1557,RIdf0d0c0_1525,
        RIdf0a3c0_1493,RIdf076c0_1461,RIdf049c0_1429,RIdefefc0_1365,RIdefc2c0_1333,RIdef95c0_1301,RIdef68c0_1269,RIdef3bc0_1237,RIdef0ec0_1205,RIdeee1c0_1173,
        RIdeeb4c0_1141,RIfc69b78_6225,RIfc6b900_6246,RIfc4d270_5900,RIfced770_7724,RIdee5ac0_1077,RIdee3d38_1056,RIdee1a10_1031,RIdedfb20_1009,RIfc7ff40_6478,
        RIfca4408_6891,RIfcb5640_7086,RIee21700_4839,RIdeda990_951,RIded8500_925,RIded61d8_900,RIded4018_876,RIded1cf0_851,RIdeceff0_819,RIdecc2f0_787,
        RIdec95f0_755,RIdeb5af0_531,RIde99a58_339,RIe16f6f8_2645,RIe15b4f0_2416,RIe144cf0_2160,RIdf396e8_2030,RIdf2dd48_1898,RIdf1e5c8_1722,RIdf01cc0_1397,
        RIdee87c0_1109,RIdedd528_982,RIde7f9a0_212,RIe19eb88_3183,RIe19be88_3151,RIfe9a698_8101,RIe199188_3119,RIfe9a530_8100,RIe196488_3087,RIe193788_3055,
        RIe190a88_3023,RIe18b088_2959,RIe188388_2927,RIfe9a800_8102,RIe185688_2895,RIfc8d938_6633,RIe182988_2863,RIe17fc88_2831,RIe17cf88_2799,RIfe9a3c8_8099,
        RIf1415a8_5203,RIfe9a260_8098,RIfe9a0f8_8097,RIfcb9150_7128,RIf13f820_5182,RIfc9fc50_6840,RIfce5340_7630,RIfc5cb58_6077,RIfc576f8_6017,RIfc780b0_6388,
        RIe1749f0_2704,RIfc7adb0_6420,RIfc7c2c8_6435,RIfcb2d78_7057,RIfc7e758_6461,RIfe9aad0_8104,RIe224ee0_4710,RIf16c3e8_5691,RIe2221e0_4678,RIfcd3898_7429,
        RIe21f4e0_4646,RIe219ae0_4582,RIe216de0_4550,RIfc880a0_6570,RIe2140e0_4518,RIf169c88_5663,RIe2113e0_4486,RIf168338_5645,RIe20e6e0_4454,RIe20b9e0_4422,
        RIe208ce0_4390,RIfce4c38_7625,RIfc9c6e0_6802,RIe2035b0_4328,RIe201af8_4309,RIfc500d8_5933,RIfc85c10_6544,RIfce81a8_7663,RIfce9c60_7682,RIf160e80_5562,
        RIf15ef90_5540,RIfe9a968_8103,RIfe9ac38_8105,RIfca8d28_6943,RIf15be58_5505,RIfcedba8_7727,RIfc6a988_6235,RIfc71cd8_6317,RIfccb198_7333,RIfcaa3a8_6959,
        RIfec3b88_8347,RIfc4c730_5892,RIfc6d688_6267,RIfca8e90_6944,RIe1f6860_4182,RIfc64e20_6170,RIfcaee30_7012,RIfccee10_7376,RIe1f4538_4157,RIfc63ea8_6159,
        RIfcaecc8_7011,RIfcae458_7005,RIfeab1c8_8263,RIe1ecc48_4071,RIe1e9f48_4039,RIe1e7248_4007,RIe1e4548_3975,RIe1e1848_3943,RIe1deb48_3911,RIe1dbe48_3879,
        RIe1d9148_3847,RIe1d3748_3783,RIe1d0a48_3751,RIe1cdd48_3719,RIe1cb048_3687,RIe1c8348_3655,RIe1c5648_3623,RIe1c2948_3591,RIe1bfc48_3559,RIfcc70e8_7287,
        RIfca7ae0_6930,RIe1ba518_3497,RIe1b8358_3473,RIfc598b8_6041,RIfcc2228_7231,RIe1b6198_3449,RIe1b4848_3431,RIfc82f10_6512,RIfc55970_5996,RIe1b3498_3417,
        RIe1b1cb0_3400,RIfcb7698_7109,RIfc4b4e8_5879,RIe1ad390_3348,RIe1abba8_3331,RIe1a9f88_3311,RIe1a7288_3279,RIe1a4588_3247,RIe1a1888_3215,RIe18dd88_2991,
        RIe17a288_2767,RIe227be0_4742,RIe21c7e0_4614,RIe205fe0_4358,RIe200040_4290,RIe1f93f8_4213,RIe1f1f40_4130,RIe1d6448_3815,RIe1bcf48_3527,RIe1afdc0_3378,
        RIe1723f8_2677,RIdec6d28_726,RIdec4028_694,RIee20bc0_4831,RIdec1328_662,RIfcbaed8_7149,RIdebe628_630,RIdebb928_598,RIdeb8c28_566,RIfc412b8_5767,
        RIdeb3228_502,RIfc9ea08_6827,RIdeb0528_470,RIee1e028_4800,RIdead828_438,RIdea7630_406,RIdea0d30_374,RIfcbac08_7147,RIfc55538_5993,RIfcba668_7143,
        RIfc4af48_5875,RIfe912f0_7996,RIfe91458_7997,RIde8be80_272,RIde87ce0_252,RIfc85238_6537,RIfc88640_6574,RIfcda210_7504,RIfcd5788_7451,RIee39418_5110,
        RIe16ce30_2616,RIfc884d8_6573,RIe169320_2574,RIe166d28_2547,RIe164028_2515,RIfe90918_7989,RIe161328_2483,RIee36880_5079,RIe15e628_2451,RIe158c28_2387,
        RIe155f28_2355,RIfe91188_7995,RIe153228_2323,RIfe91020_7994,RIe150528_2291,RIfcda378_7505,RIe14d828_2259,RIe14ab28_2227,RIe147e28_2195,RIfe90eb8_7993,
        RIfe90d50_7992,RIfcb99c0_7134,RIfc9c2a8_6799,RIfe90be8_7991,RIfe90a80_7990,RIdf3e008_2082,RIdf3bce0_2057,RIfcec690_7712,RIee30778_5010,RIfc87dd0_6568,
        RIee2e5b8_4986,RIdf36e20_2001,RIdf346c0_1973,RIdf32668_1950,RIdf30070_1923,RIee2c998_4966,RIee2aee0_4947,RIee299c8_4932,RIee28618_4918,RIfe90378_7985,
        RIfe907b0_7988,RIfe904e0_7986,RIfe90648_7987,RIfc9d928_6815,RIfc86048_6547,RIfcb92b8_7129,RIfc4ee90_5920,RIfc86a20_6554,RIdf20e90_1751,RIfcb8fe8_7127,
        RIdf1a950_1679,RIdf188f8_1656,RIdf15bf8_1624,RIdf12ef8_1592,RIdf101f8_1560,RIdf0d4f8_1528,RIdf0a7f8_1496,RIdf07af8_1464,RIdf04df8_1432,RIdeff3f8_1368,
        RIdefc6f8_1336,RIdef99f8_1304,RIdef6cf8_1272,RIdef3ff8_1240,RIdef12f8_1208,RIdeee5f8_1176,RIdeeb8f8_1144,RIfc857d8_6541,RIee24dd8_4878,RIfc4ff70_5932,
        RIfc50240_5934,RIdee5ef8_1080,RIdee4170_1059,RIfe915c0_7998,RIdedff58_1012,RIfcd4810_7440,RIee22948_4852,RIfce1560_7586,RIee219d0_4841,RIdedac60_953,
        RIfe91728_7999,RIded64a8_902,RIfe91890_8000,RIded2128_854,RIdecf428_822,RIdecc728_790,RIdec9a28_758,RIdeb5f28_534,RIde9a430_342,RIe16fb30_2648,
        RIe15b928_2419,RIe145128_2163,RIdf39b20_2033,RIdf2e180_1901,RIdf1ea00_1725,RIdf020f8_1400,RIdee8bf8_1112,RIdedd960_985,RIde80378_215,RIe19efc0_3186,
        RIe19c2c0_3154,RIf145d60_5254,RIe1995c0_3122,RIfc637a0_6154,RIe1968c0_3090,RIe193bc0_3058,RIe190ec0_3026,RIe18b4c0_2962,RIe1887c0_2930,RIfc62af8_6145,
        RIe185ac0_2898,RIfe8fc70_7980,RIe182dc0_2866,RIe1800c0_2834,RIe17d3c0_2802,RIfe90210_7984,RIfe8ff40_7982,RIfc72f20_6330,RIe176a48_2727,RIfcaf6a0_7018,
        RIfc61040_6126,RIf13e8a8_5171,RIfe900a8_7983,RIee3caf0_5149,RIee3b740_5135,RIee3a660_5123,RIe174e28_2707,RIf170768_5739,RIfc5fdf8_6113,RIf16eb48_5719,
        RIfcaaab0_6964,RIf16d1f8_5701,RIe225318_4713,RIf16c6b8_5693,RIe222618_4681,RIf16b5d8_5681,RIe21f918_4649,RIe219f18_4585,RIe217218_4553,RIfca62f8_6913,
        RIe214518_4521,RIfcc9578_7313,RIe211818_4489,RIfca5a88_6907,RIe20eb18_4457,RIe20be18_4425,RIe209118_4393,RIf167690_5636,RIf166718_5625,RIfe8f9a0_7978,
        RIfe8f838_7977,RIf165638_5613,RIf164990_5604,RIf1638b0_5592,RIf1627d0_5580,RIf161150_5564,RIf15f260_5542,RIe1fd778_4261,RIe1fc530_4248,RIf15d4d8_5521,
        RIf15c290_5508,RIfca20e0_6866,RIf159f68_5483,RIf159428_5475,RIf1581e0_5462,RIfc5ebb0_6100,RIfe8fdd8_7981,RIfc69e48_6227,RIfc5e8e0_6098,RIf154f40_5426,
        RIe1f6b30_4184,RIf153b90_5412,RIf1523a8_5395,RIfce88b0_7668,RIfe8fb08_7979,RIfcebe20_7706,RIfcb1158_7037,RIf14e730_5352,RIe1ef678_4101,RIe1ed080_4074,
        RIe1ea380_4042,RIe1e7680_4010,RIe1e4980_3978,RIe1e1c80_3946,RIe1def80_3914,RIe1dc280_3882,RIe1d9580_3850,RIe1d3b80_3786,RIe1d0e80_3754,RIe1ce180_3722,
        RIe1cb480_3690,RIe1c8780_3658,RIe1c5a80_3626,RIe1c2d80_3594,RIe1c0080_3562,RIfcc8ba0_7306,RIfc5d698_6085,RIfec35e8_8343,RIfeabd08_8271,RIfc5cf90_6080,
        RIfc5ce28_6079,RIfec31b0_8340,RIe1b4b18_3433,RIf149708_5295,RIf148358_5281,RIe1b3768_3419,RIfec3480_8342,RIfc483b0_5844,RIfc80be8_6487,RIe1ad4f8_3349,
        RIfec3318_8341,RIe1aa3c0_3314,RIe1a76c0_3282,RIe1a49c0_3250,RIe1a1cc0_3218,RIe18e1c0_2994,RIe17a6c0_2770,RIe228018_4745,RIe21cc18_4617,RIe206418_4361,
        RIe200478_4293,RIe1f9830_4216,RIe1f2378_4133,RIe1d6880_3818,RIe1bd380_3530,RIe1b01f8_3381,RIe172830_2680,RIdec6bc0_725,RIdec3ec0_693,RIee20a58_4830,
        RIdec11c0_661,RIee1f978_4818,RIdebe4c0_629,RIdebb7c0_597,RIdeb8ac0_565,RIee1efa0_4811,RIdeb30c0_501,RIfcb04b0_7028,RIdeb03c0_469,RIfc5e4a8_6095,
        RIdead6c0_437,RIdea72e8_405,RIdea09e8_373,RIfcb2508_7051,RIfcd16d8_7405,RIfc5d800_6086,RIfc63d40_6158,RIde93b30_310,RIfea7820_8222,RIfea73e8_8219,
        RIde87998_251,RIde837f8_231,RIfc7bd28_6431,RIfcc7ef8_7297,RIfc7a108_6411,RIfc7a6a8_6415,RIe16ccc8_2615,RIe16a838_2589,RIe1691b8_2573,RIe166bc0_2546,
        RIe163ec0_2514,RIee38338_5098,RIe1611c0_2482,RIfc54b60_5986,RIe15e4c0_2450,RIe158ac0_2386,RIe155dc0_2354,RIee35a70_5069,RIe1530c0_2322,RIee357a0_5067,
        RIe1503c0_2290,RIfc9fdb8_6841,RIe14d6c0_2258,RIe14a9c0_2226,RIe147cc0_2194,RIee34af8_5058,RIee33a18_5046,RIee327d0_5033,RIfcbcf30_7172,RIe142428_2131,
        RIe140100_2106,RIfea7280_8218,RIdf3bb78_2056,RIfc731f0_6332,RIee30610_5009,RIfcbe010_7184,RIee2e450_4985,RIfec2ee0_8338,RIfec3048_8339,RIfec2c10_8336,
        RIfec2d78_8337,RIfcb46c8_7075,RIfcb4830_7076,RIee29860_4931,RIfcb88e0_7122,RIdf2b480_1869,RIdf29590_1847,RIdf27268_1822,RIdf25648_1802,RIfcc9de8_7319,
        RIfc53648_5971,RIdf23a28_1782,RIfc823d0_6504,RIdf223a8_1766,RIdf20d28_1750,RIdf1bd00_1693,RIdf1a7e8_1678,RIdf18790_1655,RIdf15a90_1623,RIdf12d90_1591,
        RIdf10090_1559,RIdf0d390_1527,RIdf0a690_1495,RIdf07990_1463,RIdf04c90_1431,RIdeff290_1367,RIdefc590_1335,RIdef9890_1303,RIdef6b90_1271,RIdef3e90_1239,
        RIdef1190_1207,RIdeee490_1175,RIdeeb790_1143,RIee25be8_4888,RIfc6af28_6239,RIee23fc8_4868,RIfccf680_7382,RIdee5d90_1079,RIdee4008_1058,RIdee1ce0_1033,
        RIdedfdf0_1011,RIfc6b090_6240,RIfc534e0_5970,RIfca5920_6906,RIfc66770_6188,RIfe8f6d0_7976,RIded87d0_927,RIfe8f568_7975,RIded42e8_878,RIded1fc0_853,
        RIdecf2c0_821,RIdecc5c0_789,RIdec98c0_757,RIdeb5dc0_533,RIde9a0e8_341,RIe16f9c8_2647,RIe15b7c0_2418,RIe144fc0_2162,RIdf399b8_2032,RIdf2e018_1900,
        RIdf1e898_1724,RIdf01f90_1399,RIdee8a90_1111,RIdedd7f8_984,RIde80030_214,RIe19ee58_3185,RIe19c158_3153,RIf145bf8_5253,RIe199458_3121,RIfe8f298_7973,
        RIe196758_3089,RIe193a58_3057,RIe190d58_3025,RIe18b358_2961,RIe188658_2929,RIfe8f130_7972,RIe185958_2897,RIfc9f278_6833,RIe182c58_2865,RIe17ff58_2833,
        RIe17d258_2801,RIf1427f0_5216,RIfe8efc8_7971,RIe1779c0_2738,RIe1768e0_2726,RIfc81e30_6500,RIfc9ff20_6842,RIfca0088_6843,RIfc81b60_6498,RIfce5778_7633,
        RIfce08b8_7577,RIfc815c0_6494,RIe174cc0_2706,RIfca04c0_6846,RIfc53eb8_5977,RIfcc65a8_7279,RIfc80d50_6488,RIfc804e0_6482,RIe2251b0_4712,RIfc80378_6481,
        RIe2224b0_4680,RIfcb5910_7088,RIe21f7b0_4648,RIe219db0_4584,RIe2170b0_4552,RIfca01f0_6844,RIe2143b0_4520,RIfc82c40_6510,RIe2116b0_4488,RIfc7f6d0_6472,
        RIe20e9b0_4456,RIe20bcb0_4424,RIe208fb0_4392,RIf167528_5635,RIf1665b0_5624,RIe203718_4329,RIe201c60_4310,RIfc9da90_6816,RIfcc5360_7266,RIf163748_5591,
        RIf162668_5579,RIfc7e320_6458,RIfc87998_6565,RIe1fd610_4260,RIe1fc3c8_4247,RIf15d370_5520,RIf15c128_5507,RIfcc5d38_7273,RIfce7d70_7660,RIfc4bd58_5885,
        RIfc55c40_5998,RIfca2ab8_6873,RIe1fb450_4236,RIf156890_5444,RIfcd5ff8_7457,RIf154dd8_5425,RIfec2aa8_8335,RIfcb4b00_7078,RIfcd9400_7494,RIf151160_5382,
        RIe1f4808_4159,RIfc44738_5801,RIfc90908_6667,RIf14e5c8_5351,RIe1ef510_4100,RIe1ecf18_4073,RIe1ea218_4041,RIe1e7518_4009,RIe1e4818_3977,RIe1e1b18_3945,
        RIe1dee18_3913,RIe1dc118_3881,RIe1d9418_3849,RIe1d3a18_3785,RIe1d0d18_3753,RIe1ce018_3721,RIe1cb318_3689,RIe1c8618_3657,RIe1c5918_3625,RIe1c2c18_3593,
        RIe1bff18_3561,RIf14d218_5337,RIfe8ee60_7970,RIfea8090_8228,RIe1b84c0_3474,RIf14aab8_5309,RIfc6c170_6252,RIe1b6468_3451,RIe1b49b0_3432,RIfcafad8_7021,
        RIfcaa948_6963,RIfe8ecf8_7969,RIfe8f400_7974,RIfc67f58_6205,RIfca8ff8_6945,RIfe8eb90_7968,RIe1abe78_3333,RIe1aa258_3313,RIe1a7558_3281,RIe1a4858_3249,
        RIe1a1b58_3217,RIe18e058_2993,RIe17a558_2769,RIe227eb0_4744,RIe21cab0_4616,RIe2062b0_4360,RIe200310_4292,RIe1f96c8_4215,RIe1f2210_4132,RIe1d6718_3817,
        RIe1bd218_3529,RIe1b0090_3380,RIe1726c8_2679,RIdec4460_697,RIdec1760_665,RIee1fae0_4819,RIdebea60_633,RIee1f108_4812,RIdebbd60_601,RIdeb9060_569,
        RIdeb6360_537,RIee1eb68_4808,RIdeb0960_473,RIee1e460_4803,RIdeadc60_441,RIee1d7b8_4794,RIdea8008_409,RIdea1708_377,RIde9ae08_345,RIfe957d8_8045,
        RIfe95508_8043,RIfe95670_8044,RIee1a7e8_4760,RIfe95aa8_8047,RIfe95238_8041,RIfe95940_8046,RIfe953a0_8042,RIee1a0e0_4755,RIee19ca8_4752,RIee19870_4749,
        RIee19438_4746,RIee38ba8_5104,RIfe95c10_8048,RIee384a0_5099,RIfea9440_8242,RIe164460_2518,RIe161760_2486,RIfe942c0_8030,RIe15ea60_2454,RIfe94158_8029,
        RIe15bd60_2422,RIe156360_2358,RIe153660_2326,RIfe94428_8031,RIe150960_2294,RIfe94590_8032,RIe14dc60_2262,RIfc5c2e8_6071,RIe14af60_2230,RIe148260_2198,
        RIe145560_2166,RIee33ce8_5048,RIee32aa0_5035,RIee31858_5022,RIfc5d530_6084,RIe140538_2109,RIdf3e2d8_2084,RIdf3c118_2060,RIdf39df0_2035,RIfcdd780_7542,
        RIee2ee28_4992,RIfcc88d0_7304,RIee2cc68_4968,RIdf34990_1975,RIdf32aa0_1953,RIdf304a8_1926,RIdf2e5b8_1904,RIee2b1b0_4949,RIfe946f8_8033,RIfcb2940_7054,
        RIee273d0_4905,RIfe949c8_8035,RIdf27538_1824,RIfe94b30_8036,RIfe94860_8034,RIee26f98_4902,RIee269f8_4898,RIee26728_4896,RIee26458_4894,RIee26188_4892,
        RIfe94c98_8037,RIee25d50_4889,RIfea9170_8240,RIdf16030_1627,RIdf13330_1595,RIdf10630_1563,RIdf0d930_1531,RIdf0ac30_1499,RIdf07f30_1467,RIdf05230_1435,
        RIdf02530_1403,RIdefcb30_1339,RIdef9e30_1307,RIdef7130_1275,RIdef4430_1243,RIdef1730_1211,RIdeeea30_1179,RIdeebd30_1147,RIdee9030_1115,RIee250a8_4880,
        RIee24298_4870,RIee23758_4862,RIee22d80_4855,RIfe950d0_8040,RIfe94f68_8039,RIfe94e00_8038,RIdeddd98_988,RIee22ab0_4853,RIee21e08_4844,RIfca46d8_6893,
        RIfc5dad0_6088,RIfeaa250_8252,RIfe96048_8051,RIfe95d78_8049,RIfe95ee0_8050,RIdecf860_825,RIdeccb60_793,RIdec9e60_761,RIdec7160_729,RIdeb3660_505,
        RIde94508_313,RIe16d268_2619,RIe159060_2390,RIe142860_2134,RIdf37258_2004,RIdf2b8b8_1872,RIdf1c138_1696,RIdeff830_1371,RIdee6330_1083,RIdedb098_956,
        RIde7a450_186,RIe19c6f8_3157,RIe1999f8_3125,RIf1450b8_5245,RIe196cf8_3093,RIf143fd8_5233,RIe193ff8_3061,RIe1912f8_3029,RIe18e5f8_2997,RIe188bf8_2933,
        RIe185ef8_2901,RIfe973f8_8065,RIe1831f8_2869,RIf142958_5217,RIe1804f8_2837,RIe17d7f8_2805,RIe17aaf8_2773,RIf141b48_5207,RIfc542f0_5980,RIfc800a8_6479,
        RIe175260_2710,RIfca0bc8_6851,RIfc48680_5846,RIee3dea0_5163,RIfcc6878_7281,RIee3ba10_5137,RIee3a930_5125,RIfe97290_8064,RIe172b00_2682,RIf16f958_5729,
        RIf16ee18_5721,RIf16da68_5707,RIf16d360_5702,RIfe96e58_8061,RIe222a50_4684,RIfe96cf0_8060,RIe21fd50_4652,RIf16a660_5670,RIe21d050_4620,RIe217650_4556,
        RIe214950_4524,RIf169f58_5665,RIe211c50_4492,RIf168770_5648,RIe20ef50_4460,RIf1677f8_5637,RIe20c250_4428,RIe209550_4396,RIe206850_4364,RIf166880_5626,
        RIf1657a0_5614,RIe201dc8_4311,RIe2005e0_4294,RIfe96b88_8059,RIf163b80_5594,RIf162c08_5583,RIf161420_5566,RIf15f530_5544,RIf15d7a8_5523,RIfe968b8_8057,
        RIfe96a20_8058,RIfcb3fc0_7070,RIfc7cf70_6444,RIfc579c8_6019,RIf159590_5476,RIf1584b0_5464,RIf157268_5451,RIf1569f8_5445,RIfe965e8_8055,RIf155d50_5436,
        RIf155210_5428,RIf153e60_5414,RIfe96750_8056,RIf1527e0_5398,RIf151430_5384,RIfcd2650_7416,RIe1f2648_4135,RIf14f108_5359,RIfc7f298_6469,RIf14d4e8_5339,
        RIe1ed350_4076,RIe1ea7b8_4045,RIe1e7ab8_4013,RIe1e4db8_3981,RIe1e20b8_3949,RIe1df3b8_3917,RIe1dc6b8_3885,RIe1d99b8_3853,RIe1d6cb8_3821,RIe1d12b8_3757,
        RIe1ce5b8_3725,RIe1cb8b8_3693,RIe1c8bb8_3661,RIe1c5eb8_3629,RIe1c31b8_3597,RIe1c04b8_3565,RIe1bd7b8_3533,RIf14c138_5325,RIf14ad88_5311,RIe1b8790_3476,
        RIfe96480_8054,RIf14a0e0_5302,RIf149870_5296,RIfe97128_8063,RIfe96318_8053,RIf148628_5283,RIfc58d78_6033,RIe1b20e8_3403,RIe1b04c8_3383,RIf146cd8_5265,
        RIfc591b0_6036,RIfe961b0_8052,RIfe96fc0_8062,RIe1a7af8_3285,RIe1a4df8_3253,RIe1a20f8_3221,RIe19f3f8_3189,RIe18b8f8_2965,RIe177df8_2741,RIe225750_4716,
        RIe21a350_4588,RIe203b50_4332,RIe1fdbb0_4264,RIe1f6f68_4187,RIe1efab0_4104,RIe1d3fb8_3789,RIe1baab8_3501,RIe1ad930_3352,RIe16ff68_2651,RIdec42f8_696,
        RIdec15f8_664,RIfcc6cb0_7284,RIdebe8f8_632,RIfe93780_8022,RIdebbbf8_600,RIdeb8ef8_568,RIdeb61f8_536,RIee1ea00_4807,RIdeb07f8_472,RIee1e2f8_4802,
        RIdeadaf8_440,RIfc5d3c8_6083,RIdea7cc0_408,RIdea13c0_376,RIde9aac0_344,RIfc58238_6025,RIfcc3b78_7249,RIfc7d0d8_6445,RIfc59750_6040,RIfe93a50_8024,
        RIfe938e8_8023,RIde88370_254,RIde83e88_233,RIfc5f420_6106,RIfc976b8_6745,RIfc90a70_6668,RIfc60500_6118,RIee38a40_5103,RIe16ab08_2591,RIe169488_2575,
        RIe166ff8_2549,RIe1642f8_2517,RIe1615f8_2485,RIee369e8_5080,RIe15e8f8_2453,RIee35bd8_5070,RIe15bbf8_2421,RIe1561f8_2357,RIe1534f8_2325,RIfc3ee28_5741,
        RIe1507f8_2293,RIfce6c90_7648,RIe14daf8_2261,RIfcca7c0_7326,RIe14adf8_2229,RIe1480f8_2197,RIe1453f8_2165,RIee33b80_5047,RIee32938_5034,RIee316f0_5021,
        RIee30bb0_5013,RIe1403d0_2108,RIfe93618_8021,RIdf3bfb0_2059,RIfe934b0_8020,RIfcd0d00_7398,RIee2ecc0_4991,RIee2e720_4987,RIee2cb00_4967,RIfe93bb8_8025,
        RIdf32938_1952,RIdf30340_1925,RIdf2e450_1903,RIee2b048_4948,RIee29b30_4933,RIfc67148_6195,RIfc6fb18_6293,RIdf29860_1849,RIfe931e0_8018,RIfe93348_8019,
        RIfe93078_8017,RIfc672b0_6196,RIfca8788_6939,RIdf22510_1767,RIfcea7a0_7690,RIdf20ff8_1752,RIdf1ecd0_1727,RIdf1aab8_1680,RIfea7c58_8225,RIdf15ec8_1626,
        RIdf131c8_1594,RIdf104c8_1562,RIdf0d7c8_1530,RIdf0aac8_1498,RIdf07dc8_1466,RIdf050c8_1434,RIdf023c8_1402,RIdefc9c8_1338,RIdef9cc8_1306,RIdef6fc8_1274,
        RIdef42c8_1242,RIdef15c8_1210,RIdeee8c8_1178,RIdeebbc8_1146,RIdee8ec8_1114,RIee24f40_4879,RIee24130_4869,RIee235f0_4861,RIee22c18_4854,RIfe93d20_8026,
        RIdee1fb0_1035,RIdee0228_1014,RIdeddc30_987,RIfc684f8_6209,RIee21ca0_4843,RIfc68390_6208,RIee20d28_4832,RIded8aa0_929,RIfe93ff0_8028,RIded45b8_880,
        RIfe93e88_8027,RIdecf6f8_824,RIdecc9f8_792,RIdec9cf8_760,RIdec6ff8_728,RIdeb34f8_504,RIde941c0_312,RIe16d100_2618,RIe158ef8_2389,RIe1426f8_2133,
        RIdf370f0_2003,RIdf2b750_1871,RIdf1bfd0_1695,RIdeff6c8_1370,RIdee61c8_1082,RIdedaf30_955,RIde7a108_185,RIe19c590_3156,RIe199890_3124,RIf144f50_5244,
        RIe196b90_3092,RIfc76058_6365,RIe193e90_3060,RIe191190_3028,RIe18e490_2996,RIe188a90_2932,RIe185d90_2900,RIfccd8f8_7361,RIe183090_2868,RIfc76e68_6375,
        RIe180390_2836,RIe17d690_2804,RIe17a990_2772,RIf1419e0_5206,RIf140630_5192,RIe176bb0_2728,RIe1750f8_2709,RIfcd1840_7406,RIfc5f6f0_6108,RIee3dd38_5162,
        RIee3cc58_5150,RIee3b8a8_5136,RIee3a7c8_5124,RIee39580_5111,RIfea9008_8239,RIf16f7f0_5728,RIf16ecb0_5720,RIf16d900_5706,RIfc78ec0_6398,RIfcc8060_7298,
        RIe2228e8_4683,RIfc5a3f8_6049,RIe21fbe8_4651,RIfc74000_6342,RIe21cee8_4619,RIe2174e8_4555,RIe2147e8_4523,RIfca2c20_6874,RIe211ae8_4491,RIfca2950_6872,
        RIe20ede8_4459,RIfcc24f8_7233,RIe20c0e8_4427,RIe2093e8_4395,RIe2066e8_4363,RIfc45110_5808,RIfcc6f80_7286,RIfe92f10_8016,RIfe92970_8012,RIf164af8_5605,
        RIf163a18_5593,RIf162aa0_5582,RIfe92ad8_8013,RIf15f3c8_5543,RIf15d640_5522,RIfe92808_8011,RIfe92c40_8014,RIfe926a0_8010,RIfe92da8_8015,RIfe92538_8009,
        RIfcb5a78_7089,RIf158348_5463,RIf157100_5450,RIfc53be8_5975,RIfec38b8_8345,RIfcc5ea0_7274,RIf1550a8_5427,RIf153cf8_5413,RIfec3a20_8346,RIf152678_5397,
        RIfec3750_8344,RIf14ff18_5369,RIfe923d0_8008,RIf14efa0_5358,RIf14e898_5353,RIf14d380_5338,RIfe92268_8007,RIe1ea650_4044,RIe1e7950_4012,RIe1e4c50_3980,
        RIe1e1f50_3948,RIe1df250_3916,RIe1dc550_3884,RIe1d9850_3852,RIe1d6b50_3820,RIe1d1150_3756,RIe1ce450_3724,RIe1cb750_3692,RIe1c8a50_3660,RIe1c5d50_3628,
        RIe1c3050_3596,RIe1c0350_3564,RIe1bd650_3532,RIfcda4e0_7506,RIfc9d220_6810,RIe1b8628_3475,RIe1b6738_3453,RIfc4f2c8_5923,RIfce16c8_7587,RIfe91cc8_8003,
        RIfe91e30_8004,RIf1484c0_5282,RIf147548_5271,RIfe91f98_8005,RIfe91b60_8002,RIf146b70_5264,RIfc9f548_6835,RIfe92100_8006,RIfe919f8_8001,RIe1a7990_3284,
        RIe1a4c90_3252,RIe1a1f90_3220,RIe19f290_3188,RIe18b790_2964,RIe177c90_2740,RIe2255e8_4715,RIe21a1e8_4587,RIe2039e8_4331,RIe1fda48_4263,RIe1f6e00_4186,
        RIe1ef948_4103,RIe1d3e50_3788,RIe1ba950_3500,RIe1ad7c8_3351,RIe16fe00_2650,RIdec4730_699,RIdec1a30_667,RIfce3f90_7616,RIdebed30_635,RIfcc3308_7243,
        RIdebc030_603,RIdeb9330_571,RIdeb6630_539,RIfc8c588_6619,RIdeb0c30_475,RIfc5a998_6053,RIdeadf30_443,RIfc99b48_6771,RIdea8698_411,RIdea1d98_379,
        RIde9b498_347,RIfc78bf0_6396,RIfcbc558_7165,RIfca12d0_6856,RIfca3fd0_6888,RIfec2670_8332,RIfec2508_8331,RIde88a00_256,RIde84518_235,RIfcc35d8_7245,
        RIfcb57a8_7087,RIfc5a290_6048,RIfca3058_6877,RIee38e78_5106,RIfec27d8_8333,RIfca3328_6879,RIe1672c8_2551,RIe164730_2520,RIe161a30_2488,RIee36cb8_5082,
        RIe15ed30_2456,RIfcc7250_7288,RIe15c030_2424,RIe156630_2360,RIe153930_2328,RIfcc7688_7291,RIe150c30_2296,RIfc8af08_6603,RIe14df30_2264,RIfc9a250_6776,
        RIe14b230_2232,RIe148530_2200,RIe145830_2168,RIfc9aac0_6782,RIfc56bb8_6009,RIfca1ca8_6863,RIfcec960_7714,RIe1406a0_2110,RIdf3e440_2085,RIdf3c280_2061,
        RIdf39f58_2036,RIfc9a958_6781,RIee2f0f8_4994,RIfcdb458_7517,RIee2cf38_4970,RIdf34c60_1977,RIfec2940_8334,RIdf30778_1928,RIdf2e888_1906,RIee2b480_4951,
        RIfec23a0_8330,RIee288e8_4920,RIfec2238_8329,RIdf29b30_1851,RIdf27808_1826,RIdf25a80_1805,RIdf23e60_1785,RIfc55100_5990,RIfcd9f40_7502,RIfc54f98_5989,
        RIfc54cc8_5987,RIfc4b218_5877,RIdf1efa0_1729,RIfcc69e0_7282,RIdf18bc8_1658,RIdf16300_1629,RIdf13600_1597,RIdf10900_1565,RIdf0dc00_1533,RIdf0af00_1501,
        RIdf08200_1469,RIdf05500_1437,RIdf02800_1405,RIdefce00_1341,RIdefa100_1309,RIdef7400_1277,RIdef4700_1245,RIdef1a00_1213,RIdeeed00_1181,RIdeec000_1149,
        RIdee9300_1117,RIfce4ad0_7624,RIfc9e8a0_6826,RIfcc46b8_7257,RIfcd4108_7435,RIdee4440_1061,RIdee2280_1037,RIdee0390_1015,RIdede068_990,RIfcda0a8_7503,
        RIfce54a8_7631,RIfca0790_6848,RIfc50ee8_5943,RIded8d70_931,RIded68e0_905,RIded4888_882,RIded2560_857,RIdecfb30_827,RIdecce30_795,RIdeca130_763,
        RIdec7430_731,RIdeb3930_507,RIde94b98_315,RIe16d538_2621,RIe159330_2392,RIe142b30_2136,RIdf37528_2006,RIdf2bb88_1874,RIdf1c408_1698,RIdeffb00_1373,
        RIdee6600_1085,RIdedb368_958,RIde7aae0_188,RIe19c9c8_3159,RIe199cc8_3127,RIfe8ea28_7967,RIe196fc8_3095,RIfec20d0_8328,RIe1942c8_3063,RIe1915c8_3031,
        RIe18e8c8_2999,RIe188ec8_2935,RIe1861c8_2903,RIfc68228_6207,RIe1834c8_2871,RIfccb5d0_7336,RIe1807c8_2839,RIe17dac8_2807,RIe17adc8_2775,RIf141e18_5209,
        RIf140900_5194,RIf140090_5188,RIe1753c8_2711,RIf13f988_5183,RIf13ece0_5174,RIee3e170_5165,RIee3cf28_5152,RIee3bce0_5139,RIee3ac00_5127,RIee39850_5113,
        RIe172dd0_2684,RIf16fc28_5731,RIf16f0e8_5723,RIf16dd38_5709,RIfce9120_7674,RIfc404a8_5757,RIe222d20_4686,RIf16b8a8_5683,RIe220020_4654,RIf16a930_5672,
        RIe21d320_4622,RIe217920_4558,RIe214c20_4526,RIfc5b910_6064,RIe211f20_4494,RIfe8e8c0_7966,RIe20f220_4462,RIfe8e758_7965,RIe20c520_4430,RIe209820_4398,
        RIe206b20_4366,RIf166b50_5628,RIf165a70_5616,RIfe8dd80_7958,RIfe8dab0_7956,RIf164c60_5606,RIf163e50_5596,RIf162ed8_5585,RIf1616f0_5568,RIf15f800_5546,
        RIf15da78_5525,RIfe8d948_7955,RIfe8dc18_7957,RIf15c560_5510,RIf15b048_5495,RIfc62828_6143,RIf159860_5478,RIf158780_5466,RIf157538_5453,RIfca6e38_6921,
        RIe1f9b00_4218,RIfc61e50_6136,RIfc61748_6131,RIf154130_5416,RIe1f4ad8_4161,RIf152ab0_5400,RIf151700_5386,RIf1501e8_5371,RIe1f27b0_4136,RIfc60ed8_6125,
        RIfc7b620_6426,RIf14d7b8_5341,RIe1ed4b8_4077,RIe1eaa88_4047,RIe1e7d88_4015,RIe1e5088_3983,RIe1e2388_3951,RIe1df688_3919,RIe1dc988_3887,RIe1d9c88_3855,
        RIe1d6f88_3823,RIe1d1588_3759,RIe1ce888_3727,RIe1cbb88_3695,RIe1c8e88_3663,RIe1c6188_3631,RIe1c3488_3599,RIe1c0788_3567,RIe1bda88_3535,RIfca4de0_6898,
        RIfc5ea48_6099,RIe1b8a60_3478,RIe1b6a08_3455,RIfcbd638_7177,RIfc44fa8_5807,RIfe8e5f0_7964,RIfe8e1b8_7961,RIf1488f8_5285,RIf147818_5273,RIfe8e050_7960,
        RIfe8e488_7963,RIf146e40_5266,RIf146030_5256,RIfe8dee8_7959,RIfe8e320_7962,RIe1a7dc8_3287,RIe1a50c8_3255,RIe1a23c8_3223,RIe19f6c8_3191,RIe18bbc8_2967,
        RIe1780c8_2743,RIe225a20_4718,RIe21a620_4590,RIe203e20_4334,RIe1fde80_4266,RIe1f7238_4189,RIe1efd80_4106,RIe1d4288_3791,RIe1bad88_3503,RIe1adc00_3354,
        RIe170238_2653,RIdec45c8_698,RIdec18c8_666,RIfce85e0_7666,RIdebebc8_634,RIfcb8bb0_7124,RIdebbec8_602,RIdeb91c8_570,RIdeb64c8_538,RIfc85d78_6545,
        RIdeb0ac8_474,RIfc85aa8_6543,RIdeaddc8_442,RIfc4d3d8_5901,RIdea8350_410,RIdea1a50_378,RIde9b150_346,RIfc85ee0_6546,RIfc9c9b0_6804,RIfce13f8_7585,
        RIfcb8778_7121,RIfe8d510_7952,RIfe8d3a8_7951,RIde886b8_255,RIde841d0_234,RIde806c0_216,RIfcb8070_7116,RIfce1128_7583,RIfc9c140_6798,RIee38d10_5105,
        RIe16ac70_2592,RIfc850d0_6536,RIe167160_2550,RIe1645c8_2519,RIe1618c8_2487,RIee36b50_5081,RIe15ebc8_2455,RIee35d40_5071,RIe15bec8_2423,RIe1564c8_2359,
        RIe1537c8_2327,RIfc3ef90_5742,RIe150ac8_2295,RIfe8d7e0_7954,RIe14ddc8_2263,RIfce0fc0_7582,RIe14b0c8_2231,RIe1483c8_2199,RIe1456c8_2167,RIee33e50_5049,
        RIee32c08_5036,RIee319c0_5023,RIee30d18_5014,RIfe8cf70_7948,RIfe8ce08_7947,RIfe8d240_7950,RIfe8d0d8_7949,RIfce9dc8_7683,RIee2ef90_4993,RIfce51d8_7629,
        RIee2cdd0_4969,RIdf34af8_1976,RIfe8d678_7953,RIdf30610_1927,RIdf2e720_1905,RIee2b318_4950,RIee29c98_4934,RIee28780_4919,RIee27538_4906,RIdf299c8_1850,
        RIdf276a0_1825,RIdf25918_1804,RIdf23cf8_1784,RIfc83ff0_6524,RIfcb73c8_7107,RIfc51320_5946,RIfcdaa80_7510,RIfc83d20_6522,RIdf1ee38_1728,RIfc51b90_5952,
        RIdf18a60_1657,RIdf16198_1628,RIdf13498_1596,RIdf10798_1564,RIdf0da98_1532,RIdf0ad98_1500,RIdf08098_1468,RIdf05398_1436,RIdf02698_1404,RIdefcc98_1340,
        RIdef9f98_1308,RIdef7298_1276,RIdef4598_1244,RIdef1898_1212,RIdeeeb98_1180,RIdeebe98_1148,RIdee9198_1116,RIee25210_4881,RIee24400_4871,RIee238c0_4863,
        RIee22ee8_4856,RIfe8cca0_7946,RIdee2118_1036,RIfe8cb38_7945,RIdeddf00_989,RIfcc5a68_7271,RIee21f70_4845,RIfcb6cc0_7102,RIee20e90_4833,RIded8c08_930,
        RIded6778_904,RIded4720_881,RIded23f8_856,RIdecf9c8_826,RIdecccc8_794,RIdec9fc8_762,RIdec72c8_730,RIdeb37c8_506,RIde94850_314,RIe16d3d0_2620,
        RIe1591c8_2391,RIe1429c8_2135,RIdf373c0_2005,RIdf2ba20_1873,RIdf1c2a0_1697,RIdeff998_1372,RIdee6498_1084,RIdedb200_957,RIde7a798_187,RIe19c860_3158,
        RIe199b60_3126,RIf145220_5246,RIe196e60_3094,RIf144140_5234,RIe194160_3062,RIe191460_3030,RIe18e760_2998,RIe188d60_2934,RIe186060_2902,RIf1431c8_5223,
        RIe183360_2870,RIf142ac0_5218,RIe180660_2838,RIe17d960_2806,RIe17ac60_2774,RIf141cb0_5208,RIf140798_5193,RIf13ff28_5187,RIfe8be90_7936,RIfceb880_7702,
        RIf13eb78_5173,RIee3e008_5164,RIee3cdc0_5151,RIee3bb78_5138,RIee3aa98_5126,RIee396e8_5112,RIe172c68_2683,RIf16fac0_5730,RIf16ef80_5722,RIf16dbd0_5708,
        RIfcc4af0_7260,RIf16c820_5694,RIe222bb8_4685,RIf16b740_5682,RIe21feb8_4653,RIf16a7c8_5671,RIe21d1b8_4621,RIe2177b8_4557,RIe214ab8_4525,RIfe8c430_7940,
        RIe211db8_4493,RIf1688d8_5649,RIe20f0b8_4461,RIf167960_5638,RIe20c3b8_4429,RIe2096b8_4397,RIe2069b8_4365,RIf1669e8_5627,RIf165908_5615,RIfe8c9d0_7944,
        RIfe8c700_7942,RIfc9c578_6801,RIf163ce8_5595,RIf162d70_5584,RIf161588_5567,RIf15f698_5545,RIf15d910_5524,RIfe8c598_7941,RIfe8c868_7943,RIf15c3f8_5509,
        RIf15aee0_5494,RIf15a0d0_5484,RIf1596f8_5477,RIf158618_5465,RIf1573d0_5452,RIf156b60_5446,RIfec1f68_8327,RIf155eb8_5437,RIf155378_5429,RIf153fc8_5415,
        RIfe8bff8_7937,RIf152948_5399,RIf151598_5385,RIf150080_5370,RIfe8c2c8_7939,RIf14f270_5360,RIfc503a8_5935,RIf14d650_5340,RIfe8c160_7938,RIe1ea920_4046,
        RIe1e7c20_4014,RIe1e4f20_3982,RIe1e2220_3950,RIe1df520_3918,RIe1dc820_3886,RIe1d9b20_3854,RIe1d6e20_3822,RIe1d1420_3758,RIe1ce720_3726,RIe1cba20_3694,
        RIe1c8d20_3662,RIe1c6020_3630,RIe1c3320_3598,RIe1c0620_3566,RIe1bd920_3534,RIf14c2a0_5326,RIf14aef0_5312,RIe1b88f8_3477,RIe1b68a0_3454,RIfcd4db0_7444,
        RIfc4ebc0_5918,RIfec1e00_8326,RIfe8bd28_7935,RIf148790_5284,RIf1476b0_5272,RIfe8ba58_7933,RIfec1b30_8324,RIfc4e788_5915,RIfcb8e80_7126,RIfe8bbc0_7934,
        RIfec1c98_8325,RIe1a7c60_3286,RIe1a4f60_3254,RIe1a2260_3222,RIe19f560_3190,RIe18ba60_2966,RIe177f60_2742,RIe2258b8_4717,RIe21a4b8_4589,RIe203cb8_4333,
        RIe1fdd18_4265,RIe1f70d0_4188,RIe1efc18_4105,RIe1d4120_3790,RIe1bac20_3502,RIe1ada98_3353,RIe1700d0_2652,RIdec4a00_701,RIdec1d00_669,RIfcad7b0_6996,
        RIdebf000_637,RIfc64cb8_6169,RIdebc300_605,RIdeb9600_573,RIdeb6900_541,RIfc6f9b0_6292,RIdeb0f00_477,RIfc657f8_6177,RIdeae200_445,RIfce69c0_7646,
        RIdea8d28_413,RIdea2428_381,RIde9bb28_349,RIfc6fc80_6294,RIee1b760_4771,RIfca8080_6934,RIfe8b8f0_7932,RIde90020_292,RIde8c510_274,RIde89090_258,
        RIde84ba8_237,RIfc65ac8_6179,RIfcad210_6992,RIfcce168_7367,RIfcce2d0_7368,RIfc51488_5947,RIe16af40_2594,RIfc65c30_6180,RIe167598_2553,RIe164a00_2522,
        RIe161d00_2490,RIfc66e78_6193,RIe15f000_2458,RIfc6e498_6277,RIe15c300_2426,RIe156900_2362,RIe153c00_2330,RIfc6e330_6276,RIe150f00_2298,RIfccda60_7362,
        RIe14e200_2266,RIfc6e1c8_6275,RIe14b500_2234,RIe148800_2202,RIe145b00_2170,RIee33fb8_5050,RIee32d70_5037,RIee31c90_5025,RIee30fe8_5016,RIfea8630_8232,
        RIdf3e5a8_2086,RIdf3c550_2063,RIfea8798_8233,RIfc6e060_6274,RIfcac6d0_6984,RIfc56078_6001,RIfc6e600_6278,RIdf34dc8_1978,RIdf32d70_1955,RIfea84c8_8231,
        RIdf2eb58_1908,RIee2b750_4953,RIfc6ee70_6284,RIfc6efd8_6285,RIee27808_4908,RIfe8b788_7931,RIdf27ad8_1828,RIdf25d50_1807,RIdf24130_1787,RIfc66608_6187,
        RIfccde98_7365,RIfc66a40_6190,RIfc668d8_6189,RIfcacf40_6990,RIfeaaef8_8261,RIfc6e8d0_6280,RIdf18d30_1659,RIdf165d0_1631,RIdf138d0_1599,RIdf10bd0_1567,
        RIdf0ded0_1535,RIdf0b1d0_1503,RIdf084d0_1471,RIdf057d0_1439,RIdf02ad0_1407,RIdefd0d0_1343,RIdefa3d0_1311,RIdef76d0_1279,RIdef49d0_1247,RIdef1cd0_1215,
        RIdeeefd0_1183,RIdeec2d0_1151,RIdee95d0_1119,RIfc6dc28_6271,RIfc67c88_6203,RIfccb300_7334,RIfccd4c0_7358,RIfea81f8_8229,RIfea8360_8230,RIdee04f8_1016,
        RIdede338_992,RIfc6def8_6273,RIfcac130_6980,RIfc67b20_6202,RIfc67df0_6204,RIded9040_933,RIded6a48_906,RIded4b58_884,RIded26c8_858,RIdecfe00_829,
        RIdecd100_797,RIdeca400_765,RIdec7700_733,RIdeb3c00_509,RIde95228_317,RIe16d808_2623,RIe159600_2394,RIe142e00_2138,RIdf377f8_2008,RIdf2be58_1876,
        RIdf1c6d8_1700,RIdeffdd0_1375,RIdee68d0_1087,RIdedb638_960,RIde7b170_190,RIe19cc98_3161,RIe199f98_3129,RIfc73088_6331,RIe197298_3097,RIf1442a8_5235,
        RIe194598_3065,RIe191898_3033,RIe18eb98_3001,RIe189198_2937,RIe186498_2905,RIfc72278_6321,RIe183798_2873,RIfc61ce8_6135,RIe180a98_2841,RIe17dd98_2809,
        RIe17b098_2777,RIfcaf268_7015,RIfca6a00_6918,RIfcc9b18_7317,RIe175530_2712,RIfc72818_6325,RIfc726b0_6324,RIfccf7e8_7383,RIfc72548_6323,RIee3be48_5140,
        RIee3ad68_5128,RIfc71fa8_6319,RIe1730a0_2686,RIfcaef98_7013,RIfccf518_7381,RIfc71e40_6318,RIfc62120_6138,RIfe8b350_7928,RIe222ff0_4688,RIfcc9f50_7320,
        RIe2202f0_4656,RIfc4a570_5868,RIe21d5f0_4624,RIe217bf0_4560,RIe214ef0_4528,RIfccf3b0_7380,RIe2121f0_4496,RIf168ba8_5651,RIe20f4f0_4464,RIfc71300_6310,
        RIe20c7f0_4432,RIe209af0_4400,RIe206df0_4368,RIfc718a0_6314,RIfc71a08_6315,RIe202098_4313,RIfe8b1e8_7927,RIfc715d0_6312,RIfce6588_7643,RIfc62c60_6146,
        RIf161858_5569,RIf15fad0_5548,RIf15dbe0_5526,RIe1fc698_4249,RIfe8b4b8_7929,RIfcae5c0_7006,RIfc63098_6149,RIfc63200_6150,RIfc71198_6309,RIf158a50_5468,
        RIf1576a0_5454,RIfcdc808_7531,RIfe8b620_7930,RIfc634d0_6152,RIfcceb40_7374,RIf154400_5418,RIe1f4da8_4163,RIf152c18_5401,RIf151868_5387,RIfc4d108_5899,
        RIe1f2a80_4138,RIfc70a90_6304,RIfc63bd8_6157,RIfca7810_6928,RIe1ed788_4079,RIe1ead58_4049,RIe1e8058_4017,RIe1e5358_3985,RIe1e2658_3953,RIe1df958_3921,
        RIe1dcc58_3889,RIe1d9f58_3857,RIe1d7258_3825,RIe1d1858_3761,RIe1ceb58_3729,RIe1cbe58_3697,RIe1c9158_3665,RIe1c6458_3633,RIe1c3758_3601,RIe1c0a58_3569,
        RIe1bdd58_3537,RIf14c408_5327,RIf14b1c0_5314,RIe1b8d30_3480,RIe1b6cd8_3457,RIfc707c0_6302,RIfca7c48_6931,RIe1b4de8_3435,RIe1b3a38_3421,RIfc70220_6298,
        RIfcce870_7372,RIe1b23b8_3405,RIe1b0630_3384,RIfc645b0_6164,RIfc700b8_6297,RIfeaac28_8259,RIe1aa690_3316,RIe1a8098_3289,RIe1a5398_3257,RIe1a2698_3225,
        RIe19f998_3193,RIe18be98_2969,RIe178398_2745,RIe225cf0_4720,RIe21a8f0_4592,RIe2040f0_4336,RIe1fe150_4268,RIe1f7508_4191,RIe1f0050_4108,RIe1d4558_3793,
        RIe1bb058_3505,RIe1aded0_3356,RIe170508_2655,RIdec4898_700,RIdec1b98_668,RIfc661d0_6184,RIdebee98_636,RIfce6b28_7647,RIdebc198_604,RIdeb9498_572,
        RIdeb6798_540,RIfc40d18_5763,RIdeb0d98_476,RIfcad648_6995,RIdeae098_444,RIfcaa510_6960,RIdea89e0_412,RIdea20e0_380,RIde9b7e0_348,RIfcab320_6970,
        RIfca8350_6936,RIfc6f6e0_6290,RIfcaa240_6958,RIde8fcd8_291,RIfe8aae0_7922,RIde88d48_257,RIde84860_236,RIde80a08_217,RIfc64718_6165,RIfcae020_7002,
        RIfcadeb8_7001,RIee38fe0_5107,RIe16add8_2593,RIe1695f0_2576,RIe167430_2552,RIe164898_2521,RIe161b98_2489,RIfe8a3d8_7917,RIe15ee98_2457,RIfe8a270_7916,
        RIe15c198_2425,RIe156798_2361,RIe153a98_2329,RIfc3f0f8_5743,RIe150d98_2297,RIfcab050_6968,RIe14e098_2265,RIfcca658_7325,RIe14b398_2233,RIe148698_2201,
        RIe145998_2169,RIfe8a810_7920,RIfe8a6a8_7919,RIee31b28_5024,RIee30e80_5015,RIe140808_2111,RIfe8a540_7918,RIdf3c3e8_2062,RIdf3a0c0_2037,RIfc6b1f8_6241,
        RIee2f260_4995,RIfc70d60_6306,RIee2d0a0_4971,RIfe8a978_7921,RIdf32c08_1954,RIdf308e0_1929,RIdf2e9f0_1907,RIee2b5e8_4952,RIee29e00_4935,RIee28a50_4921,
        RIee276a0_4907,RIdf29c98_1852,RIdf27970_1827,RIdf25be8_1806,RIdf23fc8_1786,RIfc6aaf0_6236,RIfc6ac58_6237,RIdf22678_1768,RIfcdd4b0_7540,RIdf21160_1753,
        RIdf1f108_1730,RIdf1ac20_1681,RIfeaa7f0_8256,RIdf16468_1630,RIdf13768_1598,RIdf10a68_1566,RIdf0dd68_1534,RIdf0b068_1502,RIdf08368_1470,RIdf05668_1438,
        RIdf02968_1406,RIdefcf68_1342,RIdefa268_1310,RIdef7568_1278,RIdef4868_1246,RIdef1b68_1214,RIdeeee68_1182,RIdeec168_1150,RIdee9468_1118,RIee25378_4882,
        RIee24568_4872,RIee23a28_4864,RIee23050_4857,RIfe8adb0_7924,RIdee23e8_1038,RIfe8ac48_7923,RIdede1d0_991,RIfca5650_6904,RIee220d8_4846,RIfceeb20_7738,
        RIee20ff8_4834,RIded8ed8_932,RIfe8af18_7925,RIded49f0_883,RIfe8b080_7926,RIdecfc98_828,RIdeccf98_796,RIdeca298_764,RIdec7598_732,RIdeb3a98_508,
        RIde94ee0_316,RIe16d6a0_2622,RIe159498_2393,RIe142c98_2137,RIdf37690_2007,RIdf2bcf0_1875,RIdf1c570_1699,RIdeffc68_1374,RIdee6768_1086,RIdedb4d0_959,
        RIde7ae28_189,RIe19cb30_3160,RIe199e30_3128,RIf145388_5247,RIe197130_3096,RIfe8a108_7915,RIe194430_3064,RIe191730_3032,RIe18ea30_3000,RIe189030_2936,
        RIe186330_2904,RIfc6c878_6257,RIe183630_2872,RIfcabcf8_6977,RIe180930_2840,RIe17dc30_2808,RIe17af30_2776,RIfcccc50_7352,RIfcccdb8_7353,RIe176d18_2729,
        RIfea7af0_8224,RIfe89fa0_7914,RIfe89e38_7913,RIfcdd078_7537,RIfccb738_7337,RIfca9868_6951,RIfcabb90_6976,RIfca99d0_6952,RIe172f38_2685,RIf16fd90_5732,
        RIf16f250_5724,RIfc6c440_6254,RIfcaba28_6975,RIfc40610_5758,RIe222e88_4687,RIfc5d260_6082,RIe220188_4655,RIfcab758_6973,RIe21d488_4623,RIe217a88_4559,
        RIe214d88_4527,RIfe892f8_7905,RIe212088_4495,RIf168a40_5650,RIe20f388_4463,RIf167ac8_5639,RIe20c688_4431,RIe209988_4399,RIe206c88_4367,RIfc6c2d8_6253,
        RIfceec88_7739,RIe201f30_4312,RIe200748_4295,RIf164dc8_5607,RIf163fb8_5597,RIf163040_5586,RIfe895c8_7907,RIf15f968_5547,RIfe89898_7909,RIfe89460_7906,
        RIe1fb5b8_4237,RIf15c6c8_5511,RIfe89730_7908,RIf15a238_5485,RIf1599c8_5479,RIf1588e8_5467,RIfe89cd0_7912,RIfc5ba78_6065,RIe1f9c68_4219,RIfc5bd48_6067,
        RIf1554e0_5430,RIf154298_5417,RIe1f4c40_4162,RIfe89b68_7911,RIfe89a00_7910,RIf150350_5372,RIe1f2918_4137,RIf14f3d8_5361,RIfccc818_7349,RIf14d920_5342,
        RIe1ed620_4078,RIe1eabf0_4048,RIe1e7ef0_4016,RIe1e51f0_3984,RIe1e24f0_3952,RIe1df7f0_3920,RIe1dcaf0_3888,RIe1d9df0_3856,RIe1d70f0_3824,RIe1d16f0_3760,
        RIe1ce9f0_3728,RIe1cbcf0_3696,RIe1c8ff0_3664,RIe1c62f0_3632,RIe1c35f0_3600,RIe1c08f0_3568,RIe1bdbf0_3536,RIfc680c0_6206,RIf14b058_5313,RIe1b8bc8_3479,
        RIe1b6b70_3456,RIfcac298_6981,RIf1499d8_5297,RIfe89190_7904,RIfec19c8_8323,RIf148a60_5286,RIfccdd30_7364,RIe1b2250_3404,RIfec1860_8322,RIfc6e768_6279,
        RIfc54728_5983,RIe1abfe0_3334,RIe1aa528_3315,RIe1a7f30_3288,RIe1a5230_3256,RIe1a2530_3224,RIe19f830_3192,RIe18bd30_2968,RIe178230_2744,RIe225b88_4719,
        RIe21a788_4591,RIe203f88_4335,RIe1fdfe8_4267,RIe1f73a0_4190,RIe1efee8_4107,RIe1d43f0_3792,RIe1baef0_3504,RIe1add68_3355,RIe1703a0_2654,RIdec4cd0_703,
        RIdec1fd0_671,RIfc7b4b8_6425,RIdebf2d0_639,RIfc7b1e8_6423,RIdebc5d0_607,RIdeb98d0_575,RIdeb6bd0_543,RIfe83358_7837,RIdeb11d0_479,RIee1e5c8_4804,
        RIdeae4d0_447,RIfc437c0_5790,RIdea93b8_415,RIdea2ab8_383,RIde9c1b8_351,RIfc90ea8_6671,RIfc7af18_6421,RIfe83088_7835,RIee1a950_4761,RIde906b0_294,
        RIde8cba0_276,RIfe82f20_7834,RIfe82db8_7833,RIee1a248_4756,RIfe831f0_7836,RIfcc2390_7232,RIee195a0_4747,RIfcbe718_7189,RIfea9e18_8249,RIfc43220_5786,
        RIe167868_2555,RIe164cd0_2524,RIe161fd0_2492,RIee36f88_5084,RIe15f2d0_2460,RIee35ea8_5072,RIe15c5d0_2428,RIe156bd0_2364,RIe153ed0_2332,RIfe83628_7839,
        RIe1511d0_2300,RIfebfda8_8303,RIe14e4d0_2268,RIfebfc40_8302,RIe14b7d0_2236,RIe148ad0_2204,RIe145dd0_2172,RIee34120_5051,RIee32ed8_5038,RIee31df8_5026,
        RIfcc1f58_7229,RIe140ad8_2113,RIdf3e878_2088,RIfe834c0_7838,RIdf3a390_2039,RIfc5a6c8_6051,RIfc91e20_6682,RIee2e888_4988,RIfc96a10_6736,RIdf35098_1980,
        RIfeab600_8266,RIdf30bb0_1931,RIfeab768_8267,RIfcbe9e8_7191,RIfc79fa0_6410,RIfc96740_6734,RIfc92258_6685,RIfea7118_8217,RIfea95a8_8243,RIdf26020_1809,
        RIdf24400_1789,RIfc79a00_6406,RIfc5add0_6056,RIfce5d18_7637,RIfc92690_6688,RIfce3018_7605,RIdf1f270_1731,RIfc79730_6404,RIdf19000_1661,RIdf168a0_1633,
        RIdf13ba0_1601,RIdf10ea0_1569,RIdf0e1a0_1537,RIdf0b4a0_1505,RIdf087a0_1473,RIdf05aa0_1441,RIdf02da0_1409,RIdefd3a0_1345,RIdefa6a0_1313,RIdef79a0_1281,
        RIdef4ca0_1249,RIdef1fa0_1217,RIdeef2a0_1185,RIdeec5a0_1153,RIdee98a0_1121,RIfc5b7a8_6063,RIfc5b640_6062,RIfc931d0_6696,RIfcecac8_7715,RIdee4710_1063,
        RIdee26b8_1040,RIdee07c8_1018,RIdede4a0_993,RIfcbf0f0_7196,RIfcbf528_7199,RIfc792f8_6401,RIfc93068_6695,RIded91a8_934,RIded6d18_908,RIded4e28_886,
        RIded2998_860,RIded00d0_831,RIdecd3d0_799,RIdeca6d0_767,RIdec79d0_735,RIdeb3ed0_511,RIde958b8_319,RIe16dad8_2625,RIe1598d0_2396,RIe1430d0_2140,
        RIdf37ac8_2010,RIdf2c128_1878,RIdf1c9a8_1702,RIdf000a0_1377,RIdee6ba0_1089,RIdedb908_962,RIde7b800_192,RIe19cf68_3163,RIe19a268_3131,RIfc8d7d0_6632,
        RIe197568_3099,RIfc561e0_6002,RIe194868_3067,RIe191b68_3035,RIe18ee68_3003,RIe189468_2939,RIe186768_2907,RIf143330_5224,RIe183a68_2875,RIfc7d948_6451,
        RIe180d68_2843,RIe17e068_2811,RIe17b368_2779,RIfc564b0_6004,RIfcd6700_7462,RIfc461f0_5820,RIe175698_2713,RIfc46088_5819,RIfc45f20_5818,RIfc7dc18_6453,
        RIfcd69d0_7464,RIfc98630_6756,RIfcc2a98_7237,RIfc7d510_6448,RIe173208_2687,RIfc8e478_6641,RIfc45ae8_5815,RIfc8e8b0_6644,RIfc45980_5814,RIfe82ae8_7831,
        RIe2232c0_4690,RIf16ba10_5684,RIe2205c0_4658,RIfcd24e8_7415,RIe21d8c0_4626,RIe217ec0_4562,RIe2151c0_4530,RIfebf268_8295,RIe2124c0_4498,RIf168d10_5652,
        RIe20f7c0_4466,RIfc7d240_6446,RIe20cac0_4434,RIe209dc0_4402,RIe2070c0_4370,RIf166e20_5630,RIfebf6a0_8298,RIfebf808_8299,RIfebf538_8297,RIfc8eb80_6646,
        RIf164120_5598,RIfc453e0_5810,RIf161b28_5571,RIf15fc38_5549,RIf15dd48_5527,RIe1fc968_4251,RIe1fb888_4239,RIfebf3d0_8296,RIf15b318_5497,RIfca2518_6869,
        RIfc8f120_6650,RIfebfad8_8301,RIfebf970_8300,RIfc7cca0_6442,RIe1f9dd0_4220,RIfe82c50_7832,RIf155648_5431,RIfc8f288_6651,RIe1f4f10_4164,RIf152d80_5402,
        RIfc8f828_6655,RIfcb3b88_7067,RIe1f2d50_4140,RIfc445d0_5800,RIfc8faf8_6657,RIf14da88_5343,RIe1eda58_4081,RIe1eb028_4051,RIe1e8328_4019,RIe1e5628_3987,
        RIe1e2928_3955,RIe1dfc28_3923,RIe1dcf28_3891,RIe1da228_3859,RIe1d7528_3827,RIe1d1b28_3763,RIe1cee28_3731,RIe1cc128_3699,RIe1c9428_3667,RIe1c6728_3635,
        RIe1c3a28_3603,RIe1c0d28_3571,RIe1be028_3539,RIfc7bff8_6433,RIfc44030_5796,RIe1b9000_3482,RIe1b6fa8_3459,RIfcbdd40_7182,RIfc8ff30_6660,RIe1b50b8_3437,
        RIe1b3d08_3423,RIfcbe178_7185,RIfc43d60_5794,RIe1b2520_3406,RIe1b0798_3385,RIfcdb5c0_7518,RIfc7ba58_6429,RIe1ac148_3335,RIe1aa960_3318,RIe1a8368_3291,
        RIe1a5668_3259,RIe1a2968_3227,RIe19fc68_3195,RIe18c168_2971,RIe178668_2747,RIe225fc0_4722,RIe21abc0_4594,RIe2043c0_4338,RIe1fe420_4270,RIe1f77d8_4193,
        RIe1f0320_4110,RIe1d4828_3795,RIe1bb328_3507,RIe1ae1a0_3358,RIe1707d8_2657,RIdec4b68_702,RIdec1e68_670,RIfc5df08_6091,RIdebf168_638,RIfce6df8_7649,
        RIdebc468_606,RIdeb9768_574,RIdeb6a68_542,RIfc75ef0_6364,RIdeb1068_478,RIfcc12b0_7220,RIdeae368_446,RIfc5e340_6094,RIdea9070_414,RIdea2770_382,
        RIde9be70_350,RIfced4a0_7722,RIfcc1418_7221,RIfc95930_6724,RIfcec0f0_7708,RIde90368_293,RIde8c858_275,RIde893d8_259,RIde84ef0_238,RIde80d50_218,
        RIfc95a98_6725,RIfced068_7719,RIfced1d0_7720,RIfcedfe0_7730,RIe16b0a8_2595,RIe169758_2577,RIe167700_2554,RIe164b68_2523,RIe161e68_2491,RIee36e20_5083,
        RIe15f168_2459,RIfc426e0_5778,RIe15c468_2427,RIe156a68_2363,RIe153d68_2331,RIfe82818_7829,RIe151068_2299,RIee34c60_5059,RIe14e368_2267,RIfc5f9c0_6110,
        RIe14b668_2235,RIe148968_2203,RIe145c68_2171,RIfccfef0_7388,RIfca57b8_6905,RIfc600c8_6115,RIfcafda8_7023,RIe140970_2112,RIdf3e710_2087,RIdf3c6b8_2064,
        RIdf3a228_2038,RIfc5fc90_6112,RIee2f3c8_4996,RIfc742d0_6344,RIee2d208_4972,RIdf34f30_1979,RIfebf100_8294,RIdf30a48_1930,RIdf2ecc0_1909,RIfcb08e8_7031,
        RIfcee418_7733,RIfc95ed0_6728,RIfcdef68_7559,RIdf29e00_1853,RIdf27c40_1829,RIdf25eb8_1808,RIdf24298_1788,RIfc5ed18_6101,RIfcee850_7736,RIdf227e0_1769,
        RIfc5efe8_6103,RIdf212c8_1754,RIfeaa520_8254,RIdf1ad88_1682,RIdf18e98_1660,RIdf16738_1632,RIdf13a38_1600,RIdf10d38_1568,RIdf0e038_1536,RIdf0b338_1504,
        RIdf08638_1472,RIdf05938_1440,RIdf02c38_1408,RIdefd238_1344,RIdefa538_1312,RIdef7838_1280,RIdef4b38_1248,RIdef1e38_1216,RIdeef138_1184,RIdeec438_1152,
        RIdee9738_1120,RIfcc96e0_7314,RIfccfd88_7387,RIfc60aa0_6122,RIfca5ec0_6910,RIdee45a8_1062,RIdee2550_1039,RIdee0660_1017,RIfe826b0_7828,RIfcdeb30_7556,
        RIfc73bc8_6339,RIfca5bf0_6908,RIfc73a60_6338,RIfe82980_7830,RIded6bb0_907,RIded4cc0_885,RIded2830_859,RIdecff68_830,RIdecd268_798,RIdeca568_766,
        RIdec7868_734,RIdeb3d68_510,RIde95570_318,RIe16d970_2624,RIe159768_2395,RIe142f68_2139,RIdf37960_2009,RIdf2bfc0_1877,RIdf1c840_1701,RIdefff38_1376,
        RIdee6a38_1088,RIdedb7a0_961,RIde7b4b8_191,RIe19ce00_3162,RIe19a100_3130,RIfce96c0_7678,RIe197400_3098,RIf144410_5236,RIe194700_3066,RIe191a00_3034,
        RIe18ed00_3002,RIe189300_2938,RIe186600_2906,RIfebee30_8292,RIe183900_2874,RIfcdbcc8_7523,RIe180c00_2842,RIe17df00_2810,RIe17b200_2778,RIf141f80_5210,
        RIfce7398_7653,RIfcb1e00_7046,RIfe82548_7827,RIfca42a0_6890,RIfcbff00_7206,RIfcaaee8_6967,RIee3d090_5153,RIfc5c180_6070,RIfce35b8_7609,RIee399b8_5114,
        RIfea8a68_8235,RIf16fef8_5733,RIfebecc8_8291,RIfc5c450_6072,RIfce9288_7675,RIfc40778_5759,RIe223158_4689,RIfce77d0_7656,RIe220458_4657,RIfce24d8_7597,
        RIe21d758_4625,RIe217d58_4561,RIe215058_4529,RIfce8a18_7669,RIe212358_4497,RIfce1998_7589,RIe20f658_4465,RIfc77840_6382,RIe20c958_4433,RIe209c58_4401,
        RIe206f58_4369,RIf166cb8_5629,RIf165bd8_5617,RIfe81fa8_7823,RIfe81e40_7822,RIfc5c888_6075,RIfceb178_7697,RIf1631a8_5587,RIf1619c0_5570,RIfccf248_7379,
        RIfc77570_6380,RIe1fc800_4250,RIe1fb720_4238,RIf15c830_5512,RIf15b1b0_5496,RIfcd0fd0_7400,RIfccc6b0_7348,RIf158bb8_5469,RIf157808_5455,RIfc5d0f8_6081,
        RIfebef98_8293,RIfcc8a38_7305,RIfcd7ab0_7476,RIfcb1428_7039,RIfeaa0e8_8251,RIfccc548_7347,RIfce3450_7608,RIf1504b8_5373,RIe1f2be8_4139,RIf14f540_5362,
        RIfc772a0_6378,RIfcec258_7709,RIe1ed8f0_4080,RIe1eaec0_4050,RIe1e81c0_4018,RIe1e54c0_3986,RIe1e27c0_3954,RIe1dfac0_3922,RIe1dcdc0_3890,RIe1da0c0_3858,
        RIe1d73c0_3826,RIe1d19c0_3762,RIe1cecc0_3730,RIe1cbfc0_3698,RIe1c92c0_3666,RIe1c65c0_3634,RIe1c38c0_3602,RIe1c0bc0_3570,RIe1bdec0_3538,RIf14c570_5328,
        RIf14b328_5315,RIe1b8e98_3481,RIe1b6e40_3458,RIfc76760_6370,RIfc94b20_6714,RIe1b4f50_3436,RIe1b3ba0_3422,RIfcec3c0_7710,RIfceb010_7696,RIfe823e0_7826,
        RIfe82110_7824,RIfcdd8e8_7543,RIfcc0ba8_7215,RIfe82278_7825,RIe1aa7f8_3317,RIe1a8200_3290,RIe1a5500_3258,RIe1a2800_3226,RIe19fb00_3194,RIe18c000_2970,
        RIe178500_2746,RIe225e58_4721,RIe21aa58_4593,RIe204258_4337,RIe1fe2b8_4269,RIe1f7670_4192,RIe1f01b8_4109,RIe1d46c0_3794,RIe1bb1c0_3506,RIe1ae038_3357,
        RIe170670_2656,RIdec4fa0_705,RIdec22a0_673,RIee1fdb0_4821,RIdebf5a0_641,RIee1f270_4813,RIdebc8a0_609,RIdeb9ba0_577,RIdeb6ea0_545,RIee1ecd0_4809,
        RIdeb14a0_481,RIee1e730_4805,RIdeae7a0_449,RIee1d920_4795,RIdea9a48_417,RIdea3148_385,RIde9c848_353,RIee1cb10_4785,RIee1ba30_4773,RIee1b1c0_4767,
        RIfec04b0_8308,RIfe850e0_7858,RIde8d230_278,RIfea9cb0_8248,RIfe84f78_7857,RIee1a3b0_4757,RIfe853b0_7860,RIee199d8_4750,RIfe85248_7859,RIee39148_5108,
        RIe16b378_2597,RIee38608_5100,RIe167b38_2557,RIe164fa0_2526,RIe1622a0_2494,RIfe85950_7864,RIe15f5a0_2462,RIee36010_5073,RIe15c8a0_2430,RIe156ea0_2366,
        RIe1541a0_2334,RIfe85c20_7866,RIe1514a0_2302,RIee34dc8_5060,RIe14e7a0_2270,RIfc861b0_6548,RIe14baa0_2238,RIe148da0_2206,RIe1460a0_2174,RIee343f0_5053,
        RIfe85518_7861,RIfe857e8_7863,RIfe85680_7862,RIe140c40_2114,RIdf3eb48_2090,RIdf3c820_2065,RIdf3a660_2041,RIfc9d4f0_6812,RIee2f698_4998,RIfc52298_5957,
        RIee2d4d8_4974,RIdf35368_1982,RIdf32ed8_1956,RIdf30e80_1933,RIfe85ab8_7865,RIee2b8b8_4954,RIee29f68_4936,RIee28bb8_4922,RIee27970_4909,RIdf2a0d0_1855,
        RIfe84e10_7856,RIdf262f0_1811,RIfe84ca8_7855,RIee27100_4903,RIee26b60_4899,RIfcd32f8_7425,RIee265c0_4895,RIfc9e300_6822,RIdf1f540_1733,RIee25eb8_4890,
        RIfe84b40_7854,RIdf16b70_1635,RIdf13e70_1603,RIdf11170_1571,RIdf0e470_1539,RIdf0b770_1507,RIdf08a70_1475,RIdf05d70_1443,RIdf03070_1411,RIdefd670_1347,
        RIdefa970_1315,RIdef7c70_1283,RIdef4f70_1251,RIdef2270_1219,RIdeef570_1187,RIdeec870_1155,RIdee9b70_1123,RIfec0348_8307,RIfcb54d8_7085,RIee23cf8_4866,
        RIfc54e30_5988,RIfec0078_8305,RIdee2988_1042,RIfec01e0_8306,RIdede770_995,RIfcd7ee8_7479,RIfcd43d8_7437,RIfc88eb0_6580,RIfc9e5d0_6824,RIded9478_936,
        RIded6fe8_910,RIded50f8_888,RIfeab330_8264,RIded03a0_833,RIdecd6a0_801,RIdeca9a0_769,RIdec7ca0_737,RIdeb41a0_513,RIde95f48_321,RIe16dda8_2627,
        RIe159ba0_2398,RIe1433a0_2142,RIdf37d98_2012,RIdf2c3f8_1880,RIdf1cc78_1704,RIdf00370_1379,RIdee6e70_1091,RIdedbbd8_964,RIde7be90_194,RIe19d238_3165,
        RIe19a538_3133,RIf145658_5249,RIe197838_3101,RIf1446e0_5238,RIe194b38_3069,RIe191e38_3037,RIe18f138_3005,RIe189738_2941,RIe186a38_2909,RIf143600_5226,
        RIe183d38_2877,RIf142c28_5219,RIe181038_2845,RIe17e338_2813,RIe17b638_2781,RIf1420e8_5211,RIf140a68_5195,RIf1401f8_5189,RIfebff10_8304,RIf13faf0_5184,
        RIf13ee48_5175,RIee3e2d8_5166,RIee3d1f8_5154,RIee3c118_5142,RIee3b038_5130,RIee39c88_5116,RIfe838f8_7841,RIf1701c8_5735,RIfc5ab00_6054,RIf16e008_5711,
        RIfcb0e88_7035,RIf16caf0_5696,RIe223590_4692,RIf16bce0_5686,RIe220890_4660,RIf16ac00_5674,RIe21db90_4628,RIe218190_4564,RIe215490_4532,RIf16a228_5667,
        RIe212790_4500,RIf168fe0_5654,RIe20fa90_4468,RIf167d98_5641,RIe20cd90_4436,RIe20a090_4404,RIe207390_4372,RIf1670f0_5632,RIf165ea8_5619,RIe202200_4314,
        RIfe83e98_7845,RIf164f30_5608,RIf1643f0_5600,RIfce8310_7664,RIf161df8_5573,RIf15ff08_5551,RIf15e018_5529,RIfe83d30_7844,RIfe84000_7846,RIf15cb00_5514,
        RIf15b5e8_5499,RIf15a508_5487,RIfc887a8_6575,RIf158d20_5470,RIf157970_5456,RIf156cc8_5447,RIfe84438_7849,RIf156020_5438,RIfc51fc8_5955,RIf154568_5419,
        RIe1f51e0_4166,RIf153050_5404,RIf1519d0_5388,RIf150788_5375,RIfe842d0_7848,RIf14f810_5364,RIf14eb68_5355,RIf14dd58_5345,RIfe84168_7847,RIe1eb2f8_4053,
        RIe1e85f8_4021,RIe1e58f8_3989,RIe1e2bf8_3957,RIe1dfef8_3925,RIe1dd1f8_3893,RIe1da4f8_3861,RIe1d77f8_3829,RIe1d1df8_3765,RIe1cf0f8_3733,RIe1cc3f8_3701,
        RIe1c96f8_3669,RIe1c69f8_3637,RIe1c3cf8_3605,RIe1c0ff8_3573,RIe1be2f8_3541,RIf14c840_5330,RIf14b5f8_5317,RIfe83a60_7842,RIfe849d8_7853,RIfc74168_6343,
        RIf149b40_5298,RIfe83bc8_7843,RIfe84708_7851,RIf148d30_5288,RIf147ae8_5275,RIfe84870_7852,RIe1b0900_3386,RIf146fa8_5267,RIf146300_5258,RIfe845a0_7850,
        RIfe83790_7840,RIe1a8638_3293,RIe1a5938_3261,RIe1a2c38_3229,RIe19ff38_3197,RIe18c438_2973,RIe178938_2749,RIe226290_4724,RIe21ae90_4596,RIe204690_4340,
        RIe1fe6f0_4272,RIe1f7aa8_4195,RIe1f05f0_4112,RIe1d4af8_3797,RIe1bb5f8_3509,RIe1ae470_3360,RIe170aa8_2659,RIdec4e38_704,RIdec2138_672,RIee1fc48_4820,
        RIdebf438_640,RIfc49490_5856,RIdebc738_608,RIdeb9a38_576,RIdeb6d38_544,RIfc48ef0_5852,RIdeb1338_480,RIfcd9b08_7499,RIdeae638_448,RIfc8b610_6608,
        RIdea9700_416,RIdea2e00_384,RIde9c500_352,RIee1c9a8_4784,RIee1b8c8_4772,RIfc80918_6485,RIfcdad50_7512,RIfe86e68_7879,RIde8cee8_277,RIfe86d00_7878,
        RIfec0d20_8314,RIde81098_219,RIfc8b8e0_6610,RIfcd2d58_7421,RIfce4530_7620,RIfc8ba48_6611,RIe16b210_2596,RIe1698c0_2578,RIe1679d0_2556,RIe164e38_2525,
        RIe162138_2493,RIee370f0_5085,RIe15f438_2461,RIfc999e0_6770,RIe15c738_2429,RIe156d38_2365,RIe154038_2333,RIfc3f260_5744,RIe151338_2301,RIfc48518_5845,
        RIe14e638_2269,RIfc99e18_6773,RIe14b938_2237,RIe148c38_2205,RIe145f38_2173,RIee34288_5052,RIee33040_5039,RIee31f60_5027,RIfcd99a0_7498,RIfe86b98_7877,
        RIdf3e9e0_2089,RIfe86a30_7876,RIdf3a4f8_2040,RIfcc3470_7244,RIee2f530_4997,RIfc7fdd8_6477,RIee2d370_4973,RIdf35200_1981,RIfec0ff0_8316,RIdf30d18_1932,
        RIfec0e88_8315,RIfcd2a88_7419,RIfc8c858_6621,RIfc47ca8_5839,RIfcd6430_7460,RIdf29f68_1854,RIdf27da8_1830,RIdf26188_1810,RIdf24568_1790,RIfc8cb28_6623,
        RIfcdb188_7515,RIdf22948_1770,RIfc475a0_5834,RIdf21430_1755,RIdf1f3d8_1732,RIfec0bb8_8313,RIfe868c8_7875,RIdf16a08_1634,RIdf13d08_1602,RIdf11008_1570,
        RIdf0e308_1538,RIdf0b608_1506,RIdf08908_1474,RIdf05c08_1442,RIdf02f08_1410,RIdefd508_1346,RIdefa808_1314,RIdef7b08_1282,RIdef4e08_1250,RIdef2108_1218,
        RIdeef408_1186,RIdeec708_1154,RIdee9a08_1122,RIee254e0_4883,RIee246d0_4873,RIee23b90_4865,RIee231b8_4858,RIfe86fd0_7880,RIdee2820_1041,RIdee0930_1019,
        RIdede608_994,RIfc55da8_5999,RIfc98a68_6759,RIfcc3038_7241,RIfc464c0_5822,RIded9310_935,RIded6e80_909,RIded4f90_887,RIded2b00_861,RIded0238_832,
        RIdecd538_800,RIdeca838_768,RIdec7b38_736,RIdeb4038_512,RIde95c00_320,RIe16dc40_2626,RIe159a38_2397,RIe143238_2141,RIdf37c30_2011,RIdf2c290_1879,
        RIdf1cb10_1703,RIdf00208_1378,RIdee6d08_1090,RIdedba70_963,RIde7bb48_193,RIe19d0d0_3164,RIe19a3d0_3132,RIf1454f0_5248,RIe1976d0_3100,RIf144578_5237,
        RIe1949d0_3068,RIe191cd0_3036,RIe18efd0_3004,RIe1895d0_2940,RIe1868d0_2908,RIf143498_5225,RIe183bd0_2876,RIfc51758_5949,RIe180ed0_2844,RIe17e1d0_2812,
        RIe17b4d0_2780,RIfc9b060_6786,RIfc9ee40_6830,RIe176e80_2730,RIe175800_2714,RIfcb70f8_7105,RIfce0cf0_7580,RIfcc4280_7254,RIfcba7d0_7144,RIee3bfb0_5141,
        RIee3aed0_5129,RIee39b20_5115,RIe173370_2688,RIf170060_5734,RIf16f3b8_5725,RIf16dea0_5710,RIf16d4c8_5703,RIf16c988_5695,RIe223428_4691,RIf16bb78_5685,
        RIe220728_4659,RIf16aa98_5673,RIe21da28_4627,RIe218028_4563,RIe215328_4531,RIf16a0c0_5666,RIe212628_4499,RIf168e78_5653,RIe20f928_4467,RIf167c30_5640,
        RIe20cc28_4435,RIe209f28_4403,RIe207228_4371,RIf166f88_5631,RIf165d40_5618,RIfec0618_8309,RIfe86760_7874,RIfc52b08_5963,RIf164288_5599,RIf163310_5588,
        RIf161c90_5572,RIf15fda0_5550,RIf15deb0_5528,RIfe865f8_7873,RIfe85d88_7867,RIf15c998_5513,RIf15b480_5498,RIf15a3a0_5486,RIf159b30_5480,RIfc83348_6515,
        RIfc4ade0_5874,RIfc89720_6586,RIe1f9f38_4221,RIfc4ac78_5873,RIfc9f110_6832,RIfc4ab10_5872,RIe1f5078_4165,RIf152ee8_5403,RIfc899f0_6588,RIf150620_5374,
        RIe1f2eb8_4141,RIf14f6a8_5363,RIf14ea00_5354,RIf14dbf0_5344,RIe1edbc0_4082,RIe1eb190_4052,RIe1e8490_4020,RIe1e5790_3988,RIe1e2a90_3956,RIe1dfd90_3924,
        RIe1dd090_3892,RIe1da390_3860,RIe1d7690_3828,RIe1d1c90_3764,RIe1cef90_3732,RIe1cc290_3700,RIe1c9590_3668,RIe1c6890_3636,RIe1c3b90_3604,RIe1c0e90_3572,
        RIe1be190_3540,RIf14c6d8_5329,RIf14b490_5316,RIfe85ef0_7868,RIfe86490_7872,RIf14a248_5303,RIfc819f8_6497,RIfec0a50_8312,RIfe861c0_7870,RIf148bc8_5287,
        RIf147980_5274,RIfe86328_7871,RIfec0780_8310,RIfcbb478_7153,RIf146198_5257,RIfe86058_7869,RIfec08e8_8311,RIe1a84d0_3292,RIe1a57d0_3260,RIe1a2ad0_3228,
        RIe19fdd0_3196,RIe18c2d0_2972,RIe1787d0_2748,RIe226128_4723,RIe21ad28_4595,RIe204528_4339,RIe1fe588_4271,RIe1f7940_4194,RIe1f0488_4111,RIe1d4990_3796,
        RIe1bb490_3508,RIe1ae308_3359,RIe170940_2658,RIdec53d8_708,RIdec26d8_676,RIee20080_4823,RIdebf9d8_644,RIee1f3d8_4814,RIdebccd8_612,RIdeb9fd8_580,
        RIdeb72d8_548,RIee1ee38_4810,RIdeb18d8_484,RIee1e898_4806,RIdeaebd8_452,RIee1da88_4796,RIdeaa420_420,RIdea3b20_388,RIde9d220_356,RIee1cde0_4787,
        RIee1bd00_4775,RIee1b490_4769,RIfcd8a28_7487,RIde91088_297,RIde8d8c0_280,RIfe7dac0_7774,RIfe7d958_7773,RIee1a518_4758,RIee19e10_4753,RIee19b40_4751,
        RIfc768c8_6371,RIfcd05f8_7393,RIfe7dd90_7776,RIee38770_5101,RIfe7dc28_7775,RIe1653d8_2529,RIe1626d8_2497,RIee373c0_5087,RIe15f9d8_2465,RIee362e0_5075,
        RIe15ccd8_2433,RIe1572d8_2369,RIe1545d8_2337,RIfe7def8_7777,RIe1518d8_2305,RIfebdeb8_8281,RIe14ebd8_2273,RIfc649e8_6167,RIe14bed8_2241,RIe1491d8_2209,
        RIe1464d8_2177,RIfe7d7f0_7772,RIfe7d688_7771,RIee32230_5029,RIfceb9e8_7703,RIfebdd50_8280,RIfe7d520_7770,RIfebdbe8_8279,RIfe7d3b8_7769,RIfc734c0_6334,
        RIee2f968_5000,RIfccfab8_7385,RIee2d7a8_4976,RIdf357a0_1985,RIdf33310_1959,RIdf312b8_1936,RIdf2f0f8_1912,RIee2bcf0_4957,RIee2a238_4938,RIee28e88_4924,
        RIee27c40_4911,RIfe7ce18_7765,RIfe7ccb0_7764,RIfe7cf80_7766,RIfe7cb48_7763,RIee27268_4904,RIee26e30_4901,RIee26890_4897,RIfcaa0d8_6957,RIee262f0_4893,
        RIfe7d250_7768,RIee26020_4891,RIfe7d0e8_7767,RIdf16fa8_1638,RIdf142a8_1606,RIdf115a8_1574,RIdf0e8a8_1542,RIdf0bba8_1510,RIdf08ea8_1478,RIdf061a8_1446,
        RIdf034a8_1414,RIdefdaa8_1350,RIdefada8_1318,RIdef80a8_1286,RIdef53a8_1254,RIdef26a8_1222,RIdeef9a8_1190,RIdeecca8_1158,RIdee9fa8_1126,RIee25648_4884,
        RIee249a0_4875,RIfebe020_8282,RIee23488_4860,RIfebe2f0_8284,RIfebe188_8283,RIfe7e1c8_7779,RIfe7e060_7778,RIfcbf7f8_7201,RIfc7aae0_6418,RIfc787b8_6393,
        RIfc618b0_6132,RIded98b0_939,RIded72b8_912,RIded5530_891,RIded2dd0_863,RIded07d8_836,RIdecdad8_804,RIdecadd8_772,RIdec80d8_740,RIdeb45d8_516,
        RIde96920_324,RIe16e1e0_2630,RIe159fd8_2401,RIe1437d8_2145,RIdf381d0_2015,RIdf2c830_1883,RIdf1d0b0_1707,RIdf007a8_1382,RIdee72a8_1094,RIdedc010_967,
        RIde7c868_197,RIe19d670_3168,RIe19a970_3136,RIfe7b630_7748,RIe197c70_3104,RIfe7b4c8_7747,RIe194f70_3072,RIe192270_3040,RIe18f570_3008,RIe189b70_2944,
        RIe186e70_2912,RIfe7b360_7746,RIe184170_2880,RIfe7b1f8_7745,RIe181470_2848,RIe17e770_2816,RIe17ba70_2784,RIf1423b8_5213,RIf140ea0_5198,RIf140360_5190,
        RIfe7b798_7749,RIf13fc58_5185,RIf13f280_5178,RIfc79460_6402,RIee3d4c8_5156,RIfe7b090_7744,RIfe7af28_7743,RIee39df0_5117,RIe1737a8_2691,RIfe7adc0_7742,
        RIfe7ac58_7741,RIf16e440_5714,RIfcb20d0_7048,RIfe7bd38_7753,RIe2239c8_4695,RIf16be48_5687,RIe220cc8_4663,RIf16aed0_5676,RIe21dfc8_4631,RIe2185c8_4567,
        RIe2158c8_4535,RIfebd7b0_8276,RIe212bc8_4503,RIfebd648_8275,RIe20fec8_4471,RIfe7b900_7750,RIe20d1c8_4439,RIe20a4c8_4407,RIe2077c8_4375,RIf167258_5633,
        RIf166178_5621,RIe2024d0_4316,RIfe7bbd0_7752,RIf165368_5611,RIf1646c0_5602,RIfcd0a30_7396,RIf1620c8_5575,RIf1601d8_5553,RIf15e2e8_5531,RIfe7ba68_7751,
        RIfe7bea0_7754,RIf15cdd0_5516,RIf15b8b8_5501,RIf15a7d8_5489,RIfca4840_6894,RIf158ff0_5472,RIf157c40_5458,RIf156f98_5449,RIfe7c170_7756,RIf156458_5441,
        RIf155918_5433,RIf1549a0_5422,RIe1f54b0_4168,RIfe7c008_7755,RIf151b38_5389,RIf150bc0_5378,RIe1f32f0_4144,RIf14fae0_5366,RIf14ee38_5357,RIf14e028_5347,
        RIe1edff8_4085,RIe1eb730_4056,RIe1e8a30_4024,RIe1e5d30_3992,RIe1e3030_3960,RIe1e0330_3928,RIe1dd630_3896,RIe1da930_3864,RIe1d7c30_3832,RIe1d2230_3768,
        RIe1cf530_3736,RIe1cc830_3704,RIe1c9b30_3672,RIe1c6e30_3640,RIe1c4130_3608,RIe1c1430_3576,RIe1be730_3544,RIf14cb10_5332,RIf14b8c8_5319,RIfebda80_8278,
        RIfe7c878_7761,RIf14a680_5306,RIfe7c2d8_7757,RIfe7c9e0_7762,RIfe7c440_7758,RIf149000_5290,RIf147db8_5277,RIe1b2688_3407,RIfebd918_8277,RIfe7c5a8_7759,
        RIf146738_5261,RIfe7c710_7760,RIe1aad98_3321,RIe1a8a70_3296,RIe1a5d70_3264,RIe1a3070_3232,RIe1a0370_3200,RIe18c870_2976,RIe178d70_2752,RIe2266c8_4727,
        RIe21b2c8_4599,RIe204ac8_4343,RIe1feb28_4275,RIe1f7ee0_4198,RIe1f0a28_4115,RIe1d4f30_3800,RIe1bba30_3512,RIe1ae8a8_3363,RIe170ee0_2662,RIdec5270_707,
        RIdec2570_675,RIee1ff18_4822,RIdebf870_643,RIfe7f848_7795,RIdebcb70_611,RIdeb9e70_579,RIdeb7170_547,RIfe7fc80_7798,RIdeb1770_483,RIfca5d58_6909,
        RIdeaea70_451,RIfcaf808_7019,RIdeaa0d8_419,RIdea37d8_387,RIde9ced8_355,RIfcdc3d0_7528,RIfcce438_7369,RIfcb0a50_7032,RIfc75680_6358,RIde90d40_296,
        RIfe7f9b0_7796,RIde89720_260,RIde85580_240,RIde81728_221,RIfc52f40_5966,RIfc82100_6502,RIfca7108_6923,RIfe7fb18_7797,RIe16b648_2599,RIe169a28_2579,
        RIe167ca0_2558,RIe165270_2528,RIe162570_2496,RIee37258_5086,RIe15f870_2464,RIee36178_5074,RIe15cb70_2432,RIe157170_2368,RIe154470_2336,RIfc86fc0_6558,
        RIe151770_2304,RIfc4eff8_5921,RIe14ea70_2272,RIfce1290_7584,RIe14bd70_2240,RIe149070_2208,RIe146370_2176,RIee34558_5054,RIee331a8_5040,RIee320c8_5028,
        RIee31150_5017,RIfe800b8_7801,RIfe7ff50_7800,RIdf3caf0_2067,RIfe7fde8_7799,RIfcc8330_7300,RIee2f800_4999,RIfca0d30_6852,RIee2d640_4975,RIdf35638_1984,
        RIdf331a8_1958,RIdf31150_1935,RIdf2ef90_1911,RIee2bb88_4956,RIee2a0d0_4937,RIee28d20_4923,RIfe7f578_7793,RIdf2a238_1856,RIdf27f10_1831,RIfe7f6e0_7794,
        RIdf246d0_1791,RIfcce9d8_7373,RIfc63638_6153,RIdf22c18_1772,RIfc62990_6144,RIdf21700_1757,RIdf1f810_1735,RIfeaa958_8257,RIdf19168_1662,RIdf16e40_1637,
        RIdf14140_1605,RIdf11440_1573,RIdf0e740_1541,RIdf0ba40_1509,RIdf08d40_1477,RIdf06040_1445,RIdf03340_1413,RIdefd940_1349,RIdefac40_1317,RIdef7f40_1285,
        RIdef5240_1253,RIdef2540_1221,RIdeef840_1189,RIdeecb40_1157,RIdee9e40_1125,RIfcb7800_7110,RIee24838_4874,RIfc4cb68_5895,RIee23320_4859,RIfe80388_7803,
        RIdee2c58_1044,RIfe80220_7802,RIdedea40_997,RIfc98900_6758,RIee223a8_4848,RIfcc8600_7302,RIee212c8_4836,RIded9748_938,RIfe804f0_7804,RIded53c8_890,
        RIded2c68_862,RIded0670_835,RIdecd970_803,RIdecac70_771,RIdec7f70_739,RIdeb4470_515,RIde965d8_323,RIe16e078_2629,RIe159e70_2400,RIe143670_2144,
        RIdf38068_2014,RIdf2c6c8_1882,RIdf1cf48_1706,RIdf00640_1381,RIdee7140_1093,RIdedbea8_966,RIde7c520_196,RIe19d508_3167,RIe19a808_3135,RIfe7ee70_7788,
        RIe197b08_3103,RIfe7efd8_7789,RIe194e08_3071,RIe192108_3039,RIe18f408_3007,RIe189a08_2943,RIe186d08_2911,RIf143768_5227,RIe184008_2879,RIfc4bbf0_5884,
        RIe181308_2847,RIe17e608_2815,RIe17b908_2783,RIfe7f410_7792,RIf140d38_5197,RIe176fe8_2731,RIe175ad0_2716,RIfe7f2a8_7791,RIf13f118_5177,RIee3e440_5167,
        RIee3d360_5155,RIee3c280_5143,RIee3b1a0_5131,RIfe7f140_7790,RIe173640_2690,RIf170330_5736,RIf16f520_5726,RIf16e2d8_5713,RIf16d630_5704,RIfe7ea38_7785,
        RIe223860_4694,RIfc9c410_6800,RIe220b60_4662,RIfcb8340_7118,RIe21de60_4630,RIe218460_4566,RIe215760_4534,RIfc9cc80_6806,RIe212a60_4502,RIfc4ddb0_5908,
        RIe20fd60_4470,RIfc873f8_6561,RIe20d060_4438,RIe20a360_4406,RIe207660_4374,RIfc86750_6552,RIfc4e4b8_5913,RIe202368_4315,RIe200a18_4297,RIf165200_5610,
        RIf164558_5601,RIf163478_5589,RIf161f60_5574,RIf160070_5552,RIf15e180_5530,RIe1fcc38_4253,RIe1fb9f0_4240,RIf15cc68_5515,RIf15b750_5500,RIf15a670_5488,
        RIf159c98_5481,RIf158e88_5471,RIf157ad8_5457,RIf156e30_5448,RIfe7e768_7783,RIf1562f0_5440,RIf1557b0_5432,RIf154838_5421,RIfe7e8d0_7784,RIf1531b8_5405,
        RIfc52400_5958,RIf150a58_5377,RIe1f3188_4143,RIf14f978_5365,RIf14ecd0_5356,RIf14dec0_5346,RIe1ede90_4084,RIe1eb5c8_4055,RIe1e88c8_4023,RIe1e5bc8_3991,
        RIe1e2ec8_3959,RIe1e01c8_3927,RIe1dd4c8_3895,RIe1da7c8_3863,RIe1d7ac8_3831,RIe1d20c8_3767,RIe1cf3c8_3735,RIe1cc6c8_3703,RIe1c99c8_3671,RIe1c6cc8_3639,
        RIe1c3fc8_3607,RIe1c12c8_3575,RIe1be5c8_3543,RIf14c9a8_5331,RIf14b760_5318,RIfe7ed08_7787,RIfe7e600_7782,RIf14a518_5305,RIfca1f78_6865,RIfe7eba0_7786,
        RIfe7e498_7781,RIf148e98_5289,RIf147c50_5276,RIfe7e330_7780,RIe1b0a68_3387,RIf147278_5269,RIf1465d0_5260,RIe1ac418_3337,RIe1aac30_3320,RIe1a8908_3295,
        RIe1a5c08_3263,RIe1a2f08_3231,RIe1a0208_3199,RIe18c708_2975,RIe178c08_2751,RIe226560_4726,RIe21b160_4598,RIe204960_4342,RIe1fe9c0_4274,RIe1f7d78_4197,
        RIe1f08c0_4114,RIe1d4dc8_3799,RIe1bb8c8_3511,RIe1ae740_3362,RIe170d78_2661,RIdec56a8_710,RIdec29a8_678,RIfc54020_5978,RIdebfca8_646,RIee1f540_4815,
        RIdebcfa8_614,RIdeba2a8_582,RIdeb75a8_550,RIfc4fe08_5931,RIdeb1ba8_486,RIfc6b630_6244,RIdeaeea8_454,RIfc6a118_6229,RIdeaaab0_422,RIdea41b0_390,
        RIde9d8b0_358,RIfc69ce0_6226,RIee1be68_4776,RIfc653c0_6174,RIee1ac20_4763,RIde91718_299,RIde8df50_282,RIde89db0_262,RIde85c10_242,RIde81db8_223,
        RIfca76a8_6927,RIfcca4f0_7324,RIfc4ce38_5897,RIfc6b360_6242,RIe16b918_2601,RIe169cf8_2581,RIe167f70_2560,RIe1656a8_2531,RIe1629a8_2499,RIee37690_5089,
        RIe15fca8_2467,RIfce93f0_7676,RIe15cfa8_2435,RIe1575a8_2371,RIe1548a8_2339,RIee35908_5068,RIe151ba8_2307,RIee34f30_5061,RIe14eea8_2275,RIfce32e8_7607,
        RIe14c1a8_2243,RIe1494a8_2211,RIe1467a8_2179,RIfcde2c0_7550,RIfc687c8_6211,RIfca9160_6946,RIfcb1590_7040,RIe141078_2117,RIdf3ef80_2093,RIdf3cdc0_2069,
        RIfebeb60_8290,RIfc64448_6163,RIee2fad0_5001,RIfca7978_6929,RIfc676e8_6199,RIdf35a70_1987,RIdf335e0_1961,RIdf31420_1937,RIdf2f3c8_1914,RIfccef78_7377,
        RIfca6fa0_6922,RIfc62558_6141,RIfc61fb8_6137,RIfe81b70_7820,RIdf281e0_1833,RIfe81cd8_7821,RIdf249a0_1793,RIfc44300_5798,RIfcafc40_7022,RIdf22ee8_1774,
        RIfcaac18_6965,RIdf219d0_1759,RIdf1fae0_1737,RIdf1b1c0_1685,RIdf19438_1664,RIdf17278_1640,RIdf14578_1608,RIdf11878_1576,RIdf0eb78_1544,RIdf0be78_1512,
        RIdf09178_1480,RIdf06478_1448,RIdf03778_1416,RIdefdd78_1352,RIdefb078_1320,RIdef8378_1288,RIdef5678_1256,RIdef2978_1224,RIdeefc78_1192,RIdeecf78_1160,
        RIdeea278_1128,RIfc611a8_6127,RIfc61a18_6133,RIfca65c8_6915,RIfca6b68_6919,RIdee4b48_1066,RIdee2dc0_1045,RIdee0c00_1021,RIdedeba8_998,RIfc626c0_6142,
        RIfc738f8_6337,RIfcb31b0_7060,RIee21430_4837,RIded9a18_940,RIded7588_914,RIded5698_892,RIded30a0_865,RIded0aa8_838,RIdecdda8_806,RIdecb0a8_774,
        RIdec83a8_742,RIdeb48a8_518,RIde96fb0_326,RIe16e4b0_2632,RIe15a2a8_2403,RIe143aa8_2147,RIdf384a0_2017,RIdf2cb00_1885,RIdf1d380_1709,RIdf00a78_1384,
        RIdee7578_1096,RIdedc2e0_969,RIde7cef8_199,RIe19d940_3170,RIe19ac40_3138,RIfc64880_6166,RIe197f40_3106,RIf144848_5239,RIe195240_3074,RIe192540_3042,
        RIe18f840_3010,RIe189e40_2946,RIe187140_2914,RIf143a38_5229,RIe184440_2882,RIfc6f140_6286,RIe181740_2850,RIe17ea40_2818,RIe17bd40_2786,RIfc64f88_6171,
        RIf141008_5199,RIe177150_2732,RIfe81738_7817,RIfccabf8_7329,RIf13f3e8_5179,RIfca81e8_6935,RIee3d630_5157,RIfc66068_6183,RIfc6ed08_6283,RIfcdde88_7547,
        RIe173a78_2693,RIfc66338_6185,RIfc6eba0_6282,RIfc664a0_6186,RIfcacdd8_6989,RIfe81468_7815,RIe223c98_4697,RIfc66d10_6192,RIe220f98_4665,RIf16b038_5677,
        RIe21e298_4633,RIe218898_4569,RIe215b98_4537,RIfc3fc38_5751,RIe212e98_4505,RIfc67850_6200,RIe210198_4473,RIf167f00_5642,RIe20d498_4441,RIe20a798_4409,
        RIe207a98_4377,RIfcacb08_6987,RIfcac9a0_6986,RIfea8900_8234,RIfe818a0_7818,RIfca8a58_6941,RIfccad60_7330,RIfcac838_6985,RIfc67418_6197,RIf160340_5554,
        RIf15e450_5532,RIfe81a08_7819,RIfe81300_7814,RIfc6dac0_6270,RIf15ba20_5502,RIfc6d958_6269,RIfc6d7f0_6268,RIfc587d8_6029,RIfc6cf80_6262,RIfc6d3b8_6265,
        RIfe815d0_7816,RIfc6d520_6266,RIfcabe60_6978,RIfc6d0e8_6263,RIe1f5780_4170,RIfc6c5a8_6255,RIfc68d68_6215,RIfc68c00_6214,RIe1f3458_4145,RIfc68a98_6213,
        RIfccb8a0_7338,RIfca9b38_6953,RIe1ee160_4086,RIe1eba00_4058,RIe1e8d00_4026,RIe1e6000_3994,RIe1e3300_3962,RIe1e0600_3930,RIe1dd900_3898,RIe1dac00_3866,
        RIe1d7f00_3834,RIe1d2500_3770,RIe1cf800_3738,RIe1ccb00_3706,RIe1c9e00_3674,RIe1c7100_3642,RIe1c4400_3610,RIe1c1700_3578,RIe1bea00_3546,RIfc6bbd0_6248,
        RIfcdd348_7539,RIe1b9438_3485,RIe1b73e0_3462,RIfcab5f0_6972,RIfccbb70_7340,RIe1b5220_3438,RIe1b3e70_3424,RIfc6c9e0_6258,RIfcab488_6971,RIfea7dc0_8226,
        RIe1b0bd0_3388,RIfc6ce18_6261,RIfcabfc8_6979,RIe1ac580_3338,RIe1aaf00_3322,RIe1a8d40_3298,RIe1a6040_3266,RIe1a3340_3234,RIe1a0640_3202,RIe18cb40_2978,
        RIe179040_2754,RIe226998_4729,RIe21b598_4601,RIe204d98_4345,RIe1fedf8_4277,RIe1f81b0_4200,RIe1f0cf8_4117,RIe1d5200_3802,RIe1bbd00_3514,RIe1aeb78_3365,
        RIe1711b0_2664,RIdec5540_709,RIdec2840_677,RIfcc4dc0_7262,RIdebfb40_645,RIfc9d7c0_6814,RIdebce40_613,RIdeba140_581,RIdeb7440_549,RIfc4d978_5905,
        RIdeb1a40_485,RIfc9dbf8_6817,RIdeaed40_453,RIfcb8610_7120,RIdeaa768_421,RIdea3e68_389,RIde9d568_357,RIfc50678_5937,RIfc507e0_5938,RIfc9dec8_6819,
        RIfc853a0_6538,RIde913d0_298,RIde8dc08_281,RIde89a68_261,RIde858c8_241,RIde81a70_222,RIfc84860_6530,RIfc50948_5939,RIfc84c98_6533,RIfcb7da0_7114,
        RIe16b7b0_2600,RIe169b90_2580,RIe167e08_2559,RIe165540_2530,RIe162840_2498,RIee37528_5088,RIe15fb40_2466,RIfcb5be0_7090,RIe15ce40_2434,RIe157440_2370,
        RIe154740_2338,RIfcd35c8_7427,RIe151a40_2306,RIfc53a80_5974,RIe14ed40_2274,RIfcc6170_7276,RIe14c040_2242,RIe149340_2210,RIe146640_2178,RIfc7f130_6468,
        RIee33310_5041,RIfcb4f38_7081,RIfc47f78_5841,RIe140f10_2116,RIdf3ee18_2092,RIdf3cc58_2068,RIdf3a7c8_2042,RIfc7fc70_6476,RIfcd27b8_7417,RIfca1000_6854,
        RIfcc6b48_7283,RIdf35908_1986,RIdf33478_1960,RIfebe9f8_8289,RIdf2f260_1913,RIfcb7968_7111,RIee2a3a0_4939,RIfc51050_5944,RIfcd3fa0_7434,RIdf2a3a0_1857,
        RIdf28078_1832,RIfe81198_7813,RIdf24838_1792,RIfc84428_6527,RIfce7ed8_7661,RIdf22d80_1773,RIfc515f0_5948,RIdf21868_1758,RIdf1f978_1736,RIdf1b058_1684,
        RIdf192d0_1663,RIdf17110_1639,RIdf14410_1607,RIdf11710_1575,RIdf0ea10_1543,RIdf0bd10_1511,RIdf09010_1479,RIdf06310_1447,RIdf03610_1415,RIdefdc10_1351,
        RIdefaf10_1319,RIdef8210_1287,RIdef5510_1255,RIdef2810_1223,RIdeefb10_1191,RIdeece10_1159,RIdeea110_1127,RIfc7e1b8_6457,RIfca19d8_6861,RIfc7dab0_6452,
        RIfc7e488_6459,RIdee49e0_1065,RIfe80d60_7810,RIfeabba0_8270,RIfe80bf8_7809,RIfcb3750_7064,RIfce9f30_7684,RIfc7e5f0_6460,RIfc56a50_6008,RIfe81030_7812,
        RIded7420_913,RIfe80ec8_7811,RIded2f38_864,RIded0940_837,RIdecdc40_805,RIdecaf40_773,RIdec8240_741,RIdeb4740_517,RIde96c68_325,RIe16e348_2631,
        RIe15a140_2402,RIe143940_2146,RIdf38338_2016,RIdf2c998_1884,RIdf1d218_1708,RIdf00910_1383,RIdee7410_1095,RIdedc178_968,RIde7cbb0_198,RIe19d7d8_3169,
        RIe19aad8_3137,RIfcc2d68_7239,RIe197dd8_3105,RIfc5c5b8_6073,RIe1950d8_3073,RIe1923d8_3041,RIe18f6d8_3009,RIe189cd8_2945,RIe186fd8_2913,RIf1438d0_5228,
        RIe1842d8_2881,RIfc5b370_6060,RIe1815d8_2849,RIe17e8d8_2817,RIe17bbd8_2785,RIfcbb748_7155,RIfc59480_6038,RIfcbbce8_7159,RIe175c38_2717,RIfcdb890_7520,
        RIfc59b88_6043,RIfc8ada0_6602,RIfcb5eb0_7092,RIfc57c98_6021,RIfc57158_6013,RIfc58aa8_6031,RIe173910_2692,RIfcc62d8_7277,RIfc8a968_6599,RIfc57428_6015,
        RIfc56d20_6010,RIfc408e0_5760,RIe223b30_4696,RIfc82970_6508,RIe220e30_4664,RIfcecc30_7716,RIe21e130_4632,RIe218730_4568,RIe215a30_4536,RIfc3fad0_5750,
        RIe212d30_4504,RIf169148_5655,RIe210030_4472,RIfc545c0_5982,RIe20d330_4440,RIe20a630_4408,RIe207930_4376,RIfc88d48_6579,RIfc4bec0_5886,RIe202638_4317,
        RIe200b80_4298,RIfc88910_6576,RIfc4c190_5888,RIfc4c2f8_5889,RIfcba398_7141,RIfcd4270_7436,RIfcba0c8_7139,RIe1fcda0_4254,RIe1fbb58_4241,RIfc53d50_5976,
        RIfc9b768_6791,RIfc537b0_5972,RIfc4c5c8_5891,RIfc9e468_6823,RIf157da8_5459,RIfcb9f60_7138,RIe1fa208_4223,RIfc849c8_6531,RIfc529a0_5962,RIfc9f6b0_6836,
        RIe1f5618_4169,RIf153320_5406,RIfcc4988_7259,RIf150d28_5379,RIfebe458_8285,RIfc87f38_6569,RIfcb7f08_7115,RIf14e190_5348,RIfe80658_7805,RIe1eb898_4057,
        RIe1e8b98_4025,RIe1e5e98_3993,RIe1e3198_3961,RIe1e0498_3929,RIe1dd798_3897,RIe1daa98_3865,RIe1d7d98_3833,RIe1d2398_3769,RIe1cf698_3737,RIe1cc998_3705,
        RIe1c9c98_3673,RIe1c6f98_3641,RIe1c4298_3609,RIe1c1598_3577,RIe1be898_3545,RIf14cc78_5333,RIf14ba30_5320,RIe1b92d0_3484,RIe1b7278_3461,RIf14a7e8_5307,
        RIf149ca8_5299,RIfebe5c0_8286,RIfe807c0_7806,RIfc50510_5936,RIfce4f08_7627,RIfe80a90_7808,RIfebe890_8288,RIfc9cde8_6807,RIfc87560_6562,RIfe80928_7807,
        RIfebe728_8287,RIe1a8bd8_3297,RIe1a5ed8_3265,RIe1a31d8_3233,RIe1a04d8_3201,RIe18c9d8_2977,RIe178ed8_2753,RIe226830_4728,RIe21b430_4600,RIe204c30_4344,
        RIe1fec90_4276,RIe1f8048_4199,RIe1f0b90_4116,RIe1d5098_3801,RIe1bbb98_3513,RIe1aea10_3364,RIe171048_2663,RIdec5978_712,RIdec2c78_680,RIfc8aad0_6600,
        RIdebff78_648,RIfc8ac38_6601,RIdebd278_616,RIdeba578_584,RIdeb7878_552,RIfc40e80_5764,RIdeb1e78_488,RIfcdaeb8_7513,RIdeaf178_456,RIee1dbf0_4797,
        RIdeab140_424,RIdea4840_392,RIde9df40_360,RIfc8b070_6604,RIfcc38a8_7247,RIfc807b0_6484,RIfcbb8b0_7156,RIde91a60_300,RIde8e298_283,RIde8a440_264,
        RIde862a0_244,RIde82100_224,RIfcbbb80_7158,RIfc8c150_6616,RIfcbbfb8_7161,RIfc54458_5981,RIe16bbe8_2603,RIfc8c2b8_6617,RIe168240_2562,RIe165978_2533,
        RIe162c78_2501,RIee37960_5091,RIe15ff78_2469,RIfcd6b38_7465,RIe15d278_2437,RIe157878_2373,RIe154b78_2341,RIfc8e5e0_6642,RIe151e78_2309,RIfcb4290_7072,
        RIe14f178_2277,RIfc56ff0_6012,RIe14c478_2245,RIe149778_2213,RIe146a78_2181,RIee346c0_5055,RIee335e0_5043,RIee32398_5030,RIee31420_5019,RIe141348_2119,
        RIe13f020_2094,RIfec16f8_8321,RIdf3a930_2043,RIfce3e28_7615,RIfc56780_6006,RIfcb4128_7071,RIfce2eb0_7604,RIdf35d40_1989,RIfe88218_7893,RIdf316f0_1939,
        RIdf2f698_1916,RIfc7f9a0_6474,RIfce4260_7618,RIfcd62c8_7459,RIfce9990_7680,RIdf2a670_1859,RIdf284b0_1835,RIdf26728_1814,RIdf24c70_1795,RIfc7ecf8_6465,
        RIfcc31a0_7242,RIfc99008_6763,RIfc46e98_5829,RIfce2a78_7601,RIdf1fdb0_1739,RIfcc6e18_7285,RIdf19708_1666,RIdf17548_1642,RIdf14848_1610,RIdf11b48_1578,
        RIdf0ee48_1546,RIdf0c148_1514,RIdf09448_1482,RIdf06748_1450,RIdf03a48_1418,RIdefe048_1354,RIdefb348_1322,RIdef8648_1290,RIdef5948_1258,RIdef2c48_1226,
        RIdeeff48_1194,RIdeed248_1162,RIdeea548_1130,RIfcd9130_7492,RIfc7cb38_6441,RIfc97af0_6748,RIfcb3e58_7069,RIdee4e18_1068,RIdee3090_1047,RIdee0ed0_1023,
        RIfe88380_7894,RIfc97dc0_6750,RIfcc2930_7236,RIfcd9298_7493,RIfc7c868_6439,RIded9ce8_942,RIded76f0_915,RIded5968_894,RIded3370_867,RIded0d78_840,
        RIdece078_808,RIdecb378_776,RIdec8678_744,RIdeb4b78_520,RIde97640_328,RIe16e780_2634,RIe15a578_2405,RIe143d78_2149,RIdf38770_2019,RIdf2cdd0_1887,
        RIdf1d650_1711,RIdf00d48_1386,RIdee7848_1098,RIdedc5b0_971,RIde7d588_201,RIe19dc10_3172,RIe19af10_3140,RIfec1590_8320,RIe198210_3108,RIfec1428_8319,
        RIe195510_3076,RIe192810_3044,RIe18fb10_3012,RIe18a110_2948,RIe187410_2916,RIfec12c0_8318,RIe184710_2884,RIfc88370_6572,RIe181a10_2852,RIe17ed10_2820,
        RIe17c010_2788,RIfc6ccb0_6260,RIfc5f858_6109,RIfca88f0_6940,RIe175f08_2719,RIfc81020_6490,RIfcc6008_7275,RIfc4ea58_5917,RIfc42140_5774,RIfca3b98_6885,
        RIfc5ac68_6055,RIfc984c8_6755,RIe173d48_2695,RIfc9b330_6788,RIf16f688_5727,RIfc42410_5776,RIfc5f588_6107,RIfe880b0_7892,RIe223f68_4699,RIf16bfb0_5688,
        RIe221268_4667,RIfc86cf0_6556,RIe21e568_4635,RIe218b68_4571,RIe215e68_4539,RIfe87de0_7890,RIe213168_4507,RIf1692b0_5656,RIe210468_4475,RIfcdf670_7564,
        RIe20d768_4443,RIe20aa68_4411,RIe207d68_4379,RIfca6460_6914,RIf1662e0_5622,RIe202908_4319,RIfe87b10_7888,RIfc58c10_6032,RIfc50ab0_5940,RIfccd790_7360,
        RIfccd1f0_7356,RIf160610_5556,RIf15e720_5534,RIfe87c78_7889,RIfe87f48_7891,RIfce7668_7655,RIfc86480_6550,RIfcd2218_7413,RIfcb01e0_7026,RIfc47b40_5838,
        RIfc84158_6525,RIfc4b920_5882,RIe1fa4d8_4225,RIfc4ba88_5883,RIfcb7530_7108,RIfcd58f0_7452,RIe1f5a50_4172,RIf153488_5407,RIf151ca0_5390,RIfc51e60_5954,
        RIe1f3728_4147,RIfc9aef8_6785,RIfcbaaa0_7146,RIfc52130_5956,RIe1ee430_4088,RIe1ebcd0_4060,RIe1e8fd0_4028,RIe1e62d0_3996,RIe1e35d0_3964,RIe1e08d0_3932,
        RIe1ddbd0_3900,RIe1daed0_3868,RIe1d81d0_3836,RIe1d27d0_3772,RIe1cfad0_3740,RIe1ccdd0_3708,RIe1ca0d0_3676,RIe1c73d0_3644,RIe1c46d0_3612,RIe1c19d0_3580,
        RIe1becd0_3548,RIfce0b88_7579,RIfc82808_6507,RIe1b9708_3487,RIe1b76b0_3464,RIfcd5bc0_7454,RIfcb69f0_7100,RIe1b54f0_3440,RIe1b4140_3426,RIfc89f90_6592,
        RIfce9af8_7681,RIe1b2958_3409,RIe1b0ea0_3390,RIfc4a138_5865,RIfc8a260_6594,RIe1ac850_3340,RIe1ab1d0_3324,RIe1a9010_3300,RIe1a6310_3268,RIe1a3610_3236,
        RIe1a0910_3204,RIe18ce10_2980,RIe179310_2756,RIe226c68_4731,RIe21b868_4603,RIe205068_4347,RIe1ff0c8_4279,RIe1f8480_4202,RIe1f0fc8_4119,RIe1d54d0_3804,
        RIe1bbfd0_3516,RIe1aee48_3367,RIe171480_2666,RIdec5810_711,RIdec2b10_679,RIfce6f60_7650,RIdebfe10_647,RIfc95228_6719,RIdebd110_615,RIdeba410_583,
        RIdeb7710_551,RIfe879a8_7887,RIdeb1d10_487,RIfcc16e8_7223,RIdeaf010_455,RIfca4f48_6899,RIdeaadf8_423,RIdea44f8_391,RIde9dbf8_359,RIee1cf48_4788,
        RIee1bfd0_4777,RIfc95660_6722,RIfcee148_7731,RIfe87840_7886,RIfe876d8_7885,RIde8a0f8_263,RIde85f58_243,RIfcb0780_7030,RIfcee9b8_7737,RIfc5f150_6104,
        RIfcdee00_7558,RIfcd8050_7480,RIe16ba80_2602,RIfca5380_6902,RIe1680d8_2561,RIe165810_2532,RIe162b10_2500,RIee377f8_5090,RIe15fe10_2468,RIee36448_5076,
        RIe15d110_2436,RIe157710_2372,RIe154a10_2340,RIfc3f3c8_5745,RIe151d10_2308,RIfcde9c8_7555,RIe14f010_2276,RIfc4a2a0_5866,RIe14c310_2244,RIe149610_2212,
        RIe146910_2180,RIfc62288_6139,RIee33478_5042,RIfc71b70_6316,RIee312b8_5018,RIe1411e0_2118,RIfe87570_7884,RIdf3cf28_2070,RIfe87408_7883,RIfcc99b0_7316,
        RIfccf0e0_7378,RIfcaeb60_7010,RIfcca220_7322,RIdf35bd8_1988,RIdf33748_1962,RIdf31588_1938,RIdf2f530_1915,RIee2be58_4958,RIee2a508_4940,RIee28ff0_4925,
        RIee27da8_4912,RIdf2a508_1858,RIdf28348_1834,RIdf265c0_1813,RIdf24b08_1794,RIfc74708_6347,RIfc42578_5777,RIfc43388_5787,RIfc745a0_6346,RIfcb0078_7025,
        RIdf1fc48_1738,RIfcaff10_7024,RIdf195a0_1665,RIdf173e0_1641,RIdf146e0_1609,RIdf119e0_1577,RIdf0ece0_1545,RIdf0bfe0_1513,RIdf092e0_1481,RIdf065e0_1449,
        RIdf038e0_1417,RIdefdee0_1353,RIdefb1e0_1321,RIdef84e0_1289,RIdef57e0_1257,RIdef2ae0_1225,RIdeefde0_1193,RIdeed0e0_1161,RIdeea3e0_1129,RIee257b0_4885,
        RIfca73d8_6925,RIee23e60_4867,RIfce66f0_7644,RIdee4cb0_1067,RIdee2f28_1046,RIdee0d68_1022,RIdeded10_999,RIfcca388_7323,RIfce6858_7645,RIfcceca8_7375,
        RIfcdc970_7532,RIded9b80_941,RIfeaaac0_8258,RIded5800_893,RIded3208_866,RIded0c10_839,RIdecdf10_807,RIdecb210_775,RIdec8510_743,RIdeb4a10_519,
        RIde972f8_327,RIe16e618_2633,RIe15a410_2404,RIe143c10_2148,RIdf38608_2018,RIdf2cc68_1886,RIdf1d4e8_1710,RIdf00be0_1385,RIdee76e0_1097,RIdedc448_970,
        RIde7d240_200,RIe19daa8_3171,RIe19ada8_3139,RIf1457c0_5250,RIe1980a8_3107,RIf1449b0_5240,RIe1953a8_3075,RIe1926a8_3043,RIe18f9a8_3011,RIe189fa8_2947,
        RIe1872a8_2915,RIf143ba0_5230,RIe1845a8_2883,RIfc912e0_6674,RIe1818a8_2851,RIe17eba8_2819,RIe17bea8_2787,RIfc915b0_6676,RIfcbe5b0_7188,RIfce3b58_7613,
        RIe175da0_2718,RIfceb448_7699,RIfcc7958_7293,RIfc42de8_5783,RIfc96e48_6739,RIfc7a810_6416,RIfc96ce0_6738,RIfcc7ac0_7294,RIe173be0_2694,RIfce39f0_7612,
        RIfc7a540_6414,RIfc91b50_6680,RIfc429b0_5780,RIfea9710_8244,RIe223e00_4698,RIfcd8488_7483,RIe221100_4666,RIfc920f0_6684,RIe21e400_4634,RIe218a00_4570,
        RIe215d00_4538,RIfc79e38_6409,RIe213000_4506,RIfcbee20_7194,RIe210300_4474,RIf168068_5643,RIe20d600_4442,RIe20a900_4410,RIe207c00_4378,RIfc5af38_6057,
        RIfcd73a8_7471,RIe2027a0_4318,RIe200ce8_4299,RIfcb2670_7052,RIfcdf940_7566,RIfc5b208_6059,RIfcbf3c0_7198,RIf1604a8_5555,RIf15e5b8_5533,RIfe872a0_7882,
        RIfe87138_7881,RIfc78920_6394,RIfec1158_8317,RIfc93338_6697,RIfcea368_7687,RIfcb23a0_7050,RIfc5bbe0_6066,RIfcede78_7729,RIe1fa370_4224,RIfcd4c48_7443,
        RIfce1dd0_7592,RIfcbf960_7202,RIe1f58e8_4171,RIfcbfc30_7204,RIfc78380_6390,RIfc93770_6700,RIe1f35c0_4146,RIfcb1f68_7047,RIfce1b00_7590,RIfc93a40_6702,
        RIe1ee2c8_4087,RIe1ebb68_4059,RIe1e8e68_4027,RIe1e6168_3995,RIe1e3468_3963,RIe1e0768_3931,RIe1dda68_3899,RIe1dad68_3867,RIe1d8068_3835,RIe1d2668_3771,
        RIe1cf968_3739,RIe1ccc68_3707,RIe1c9f68_3675,RIe1c7268_3643,RIe1c4568_3611,RIe1c1868_3579,RIe1beb68_3547,RIfcdec98_7557,RIfc94148_6707,RIe1b95a0_3486,
        RIe1b7548_3463,RIfcd12a0_7402,RIfceabd8_7693,RIe1b5388_3439,RIe1b3fd8_3425,RIfc94850_6712,RIfcd7c18_7477,RIe1b27f0_3408,RIe1b0d38_3389,RIfc76a30_6372,
        RIfce2640_7598,RIe1ac6e8_3339,RIe1ab068_3323,RIe1a8ea8_3299,RIe1a61a8_3267,RIe1a34a8_3235,RIe1a07a8_3203,RIe18cca8_2979,RIe1791a8_2755,RIe226b00_4730,
        RIe21b700_4602,RIe204f00_4346,RIe1fef60_4278,RIe1f8318_4201,RIe1f0e60_4118,RIe1d5368_3803,RIe1bbe68_3515,RIe1aece0_3366,RIe171318_2665,RIdec5c48_714,
        RIdec2f48_682,RIfc7c160_6434,RIdec0248_650,RIfcb38b8_7065,RIdebd548_618,RIdeba848_586,RIdeb7b48_554,RIfce7c08_7659,RIdeb2148_490,RIfce7aa0_7658,
        RIdeaf448_458,RIfca38c8_6883,RIdeab7d0_426,RIdea4ed0_394,RIde9e5d0_362,RIfc41e70_5772,RIfc5b0a0_6058,RIfcdbb60_7522,RIfc78650_6392,RIfea92d8_8241,
        RIde8e5e0_284,RIfea0d40_8174,RIfea0bd8_8173,RIfcdf508_7563,RIfcb1b30_7044,RIfc5ccc0_6078,RIfcb16f8_7041,RIfc77b10_6384,RIe16beb8_2605,RIe169e60_2582,
        RIe168510_2564,RIe165c48_2535,RIe162f48_2503,RIfc4f9d0_5928,RIe160248_2471,RIfc4e8f0_5916,RIe15d548_2439,RIe157b48_2375,RIe154e48_2343,RIfc4e1e8_5911,
        RIe152148_2311,RIfc868b8_6553,RIe14f448_2279,RIfc865e8_6551,RIe14c748_2247,RIe149a48_2215,RIe146d48_2183,RIfc9eb70_6828,RIfc9ecd8_6829,RIfcc5630_7268,
        RIfc83bb8_6521,RIe141618_2121,RIfea0ea8_8175,RIdf3d1f8_2072,RIdf3ac00_2045,RIee308e0_5011,RIfcd3cd0_7432,RIfc84e00_6534,RIfc834b0_6516,RIdf36010_1991,
        RIdf33a18_1964,RIdf31858_1940,RIdf2f968_1918,RIee2c128_4960,RIee2a7d8_4942,RIee292c0_4927,RIee28078_4914,RIdf2a940_1861,RIdf28780_1837,RIfea0a70_8172,
        RIfea0908_8171,RIfcd4f18_7445,RIfca0628_6847,RIdf23050_1775,RIfcd3190_7424,RIdf21b38_1760,RIdf20080_1741,RIdf1b328_1686,RIdf199d8_1668,RIdf17818_1644,
        RIdf14b18_1612,RIdf11e18_1580,RIdf0f118_1548,RIdf0c418_1516,RIdf09718_1484,RIdf06a18_1452,RIdf03d18_1420,RIdefe318_1356,RIdefb618_1324,RIdef8918_1292,
        RIdef5c18_1260,RIdef2f18_1228,RIdef0218_1196,RIdeed518_1164,RIdeea818_1132,RIfcdf3a0_7562,RIfca5218_6901,RIfcdc538_7529,RIfcdc6a0_7530,RIdee50e8_1070,
        RIdee3360_1049,RIfea07a0_8170,RIdedefe0_1001,RIfcb0d20_7034,RIfcd4978_7441,RIfca49a8_6895,RIfca1708_6859,RIded9fb8_944,RIded79c0_917,RIded5ad0_895,
        RIfeab498_8265,RIded1048_842,RIdece348_810,RIdecb648_778,RIdec8948_746,RIdeb4e48_522,RIde97cd0_330,RIe16ea50_2636,RIe15a848_2407,RIe144048_2151,
        RIdf38a40_2021,RIdf2d0a0_1889,RIdf1d920_1713,RIdf01018_1388,RIdee7b18_1100,RIdedc880_973,RIde7dc18_203,RIe19dee0_3174,RIe19b1e0_3142,RIfc67580_6198,
        RIe1984e0_3110,RIfccb030_7332,RIe1957e0_3078,RIe192ae0_3046,RIe18fde0_3014,RIe18a3e0_2950,RIe1876e0_2918,RIfc6a550_6232,RIe1849e0_2886,RIfcaa7e0_6962,
        RIe181ce0_2854,RIe17efe0_2822,RIe17c2e0_2790,RIfc65d98_6181,RIfc65690_6176,RIe1772b8_2733,RIfea0638_8169,RIfcca928_7327,RIfc607d0_6120,RIfc65258_6173,
        RIee3d798_5158,RIee3c3e8_5144,RIfca9430_6948,RIee39f58_5118,RIe174018_2697,RIfcecf00_7718,RIfc650f0_6172,RIf16e5a8_5715,RIfc43a90_5792,RIfc65528_6175,
        RIe224238_4701,RIfca9f70_6956,RIe221538_4669,RIfc6b4c8_6243,RIe21e838_4637,RIe218e38_4573,RIe216138_4541,RIfc3fda0_5752,RIe213438_4509,RIfc61310_6128,
        RIe210738_4477,RIfc60c08_6123,RIe20da38_4445,RIe20ad38_4413,RIe208038_4381,RIfc66ba8_6191,RIfccbcd8_7341,RIe202bd8_4321,RIe200fb8_4301,RIfcadbe8_6999,
        RIfccbe40_7342,RIfca7540_6926,RIfc6a3e8_6231,RIfca6898_6917,RIfc73358_6333,RIe1fd070_4256,RIe1fbe28_4243,RIfcc2660_7234,RIfc44468_5799,RIf15a940_5490,
        RIfca7270_6924,RIfc5e070_6092,RIfc5dda0_6090,RIfc7e050_6456,RIe1fa7a8_4227,RIfc5d968_6087,RIfcd9568_7495,RIfc8d668_6631,RIe1f5d20_4174,RIfca4138_6889,
        RIfc8cdf8_6625,RIfcc7c28_7295,RIe1f39f8_4149,RIfc99440_6766,RIfcbc3f0_7164,RIfc5a128_6047,RIe1ee700_4090,RIe1ebfa0_4062,RIe1e92a0_4030,RIe1e65a0_3998,
        RIe1e38a0_3966,RIe1e0ba0_3934,RIe1ddea0_3902,RIe1db1a0_3870,RIe1d84a0_3838,RIe1d2aa0_3774,RIe1cfda0_3742,RIe1cd0a0_3710,RIe1ca3a0_3678,RIe1c76a0_3646,
        RIe1c49a0_3614,RIe1c1ca0_3582,RIe1befa0_3550,RIf14cde0_5334,RIf14bb98_5321,RIe1b99d8_3489,RIe1b7980_3466,RIfc4c460_5890,RIfc9e738_6825,RIe1b5658_3441,
        RIfec54d8_8365,RIf149168_5291,RIf147f20_5278,RIe1b2ac0_3410,RIe1b1170_3392,RIf1473e0_5270,RIf1468a0_5262,RIe1acb20_3342,RIe1ab338_3325,RIe1a92e0_3302,
        RIe1a65e0_3270,RIe1a38e0_3238,RIe1a0be0_3206,RIe18d0e0_2982,RIe1795e0_2758,RIe226f38_4733,RIe21bb38_4605,RIe205338_4349,RIe1ff398_4281,RIe1f8750_4204,
        RIe1f1298_4121,RIe1d57a0_3806,RIe1bc2a0_3518,RIe1af118_3369,RIe171750_2668,RIdec5ae0_713,RIdec2de0_681,RIfc82268_6503,RIdec00e0_649,RIfcb8d18_7125,
        RIdebd3e0_617,RIdeba6e0_585,RIdeb79e0_553,RIfcb9858_7133,RIdeb1fe0_489,RIfc9efa8_6831,RIdeaf2e0_457,RIfce0750_7576,RIdeab488_425,RIdea4b88_393,
        RIde9e288_361,RIee1d0b0_4789,RIee1c138_4778,RIfcd0e68_7399,RIfc76d00_6374,RIfe89028_7903,RIfe88d58_7901,RIfe88ec0_7902,RIfe88bf0_7900,RIfcda7b0_7508,
        RIfc4d810_5904,RIfc52dd8_5965,RIfcde590_7552,RIfc4f868_5927,RIe16bd50_2604,RIfc68930_6212,RIe1683a8_2563,RIe165ae0_2534,RIe162de0_2502,RIfe88a88_7899,
        RIe1600e0_2470,RIfcc9140_7310,RIe15d3e0_2438,RIe1579e0_2374,RIe154ce0_2342,RIfc698a8_6223,RIe151fe0_2310,RIee35098_5062,RIe14f2e0_2278,RIfcc0338_7209,
        RIe14c5e0_2246,RIe1498e0_2214,RIe146be0_2182,RIfc88208_6571,RIfc85670_6540,RIfc81f98_6501,RIfcc4f28_7263,RIe1414b0_2120,RIe13f188_2095,RIdf3d090_2071,
        RIdf3aa98_2044,RIfcd2920_7418,RIfc7d7e0_6450,RIfc49760_5858,RIfce5a48_7635,RIdf35ea8_1990,RIdf338b0_1963,RIfe88920_7898,RIdf2f800_1917,RIee2bfc0_4959,
        RIee2a670_4941,RIee29158_4926,RIee27f10_4913,RIdf2a7d8_1860,RIdf28618_1836,RIdf26890_1815,RIdf24dd8_1796,RIfcad918_6997,RIfc69fb0_6228,RIfc63368_6151,
        RIfc623f0_6140,RIfc60938_6121,RIdf1ff18_1740,RIfcba500_7142,RIdf19870_1667,RIdf176b0_1643,RIdf149b0_1611,RIdf11cb0_1579,RIdf0efb0_1547,RIdf0c2b0_1515,
        RIdf095b0_1483,RIdf068b0_1451,RIdf03bb0_1419,RIdefe1b0_1355,RIdefb4b0_1323,RIdef87b0_1291,RIdef5ab0_1259,RIdef2db0_1227,RIdef00b0_1195,RIdeed3b0_1163,
        RIdeea6b0_1131,RIfcc9848_7315,RIfc69a10_6224,RIfcacc70_6988,RIfccbfa8_7343,RIdee4f80_1069,RIdee31f8_1048,RIdee1038_1024,RIdedee78_1000,RIfc84590_6528,
        RIfc9bba0_6794,RIee21b38_4842,RIfc47168_5831,RIded9e50_943,RIded7858_916,RIfe887b8_7897,RIded34d8_868,RIded0ee0_841,RIdece1e0_809,RIdecb4e0_777,
        RIdec87e0_745,RIdeb4ce0_521,RIde97988_329,RIe16e8e8_2635,RIe15a6e0_2406,RIe143ee0_2150,RIdf388d8_2020,RIdf2cf38_1888,RIdf1d7b8_1712,RIdf00eb0_1387,
        RIdee79b0_1099,RIdedc718_972,RIde7d8d0_202,RIe19dd78_3173,RIe19b078_3141,RIfca1438_6857,RIe198378_3109,RIfca35f8_6881,RIe195678_3077,RIe192978_3045,
        RIe18fc78_3013,RIe18a278_2949,RIe187578_2917,RIfcba230_7140,RIe184878_2885,RIf142d90_5220,RIe181b78_2853,RIe17ee78_2821,RIe17c178_2789,RIfc9be70_6796,
        RIfc9bd08_6795,RIfc4ccd0_5896,RIe176070_2720,RIfc87c68_6567,RIfc87b00_6566,RIfcc4c58_7261,RIfc4fca0_5930,RIfc4f598_5925,RIfc876c8_6563,RIfc4dae0_5906,
        RIe173eb0_2696,RIfcb9420_7130,RIfc4e080_5910,RIfc4e350_5912,RIfc9d388_6811,RIfc40a48_5761,RIe2240d0_4700,RIfc85508_6539,RIe2213d0_4668,RIfc9ba38_6793,
        RIe21e6d0_4636,RIe218cd0_4572,RIe215fd0_4540,RIfc52c70_5964,RIe2132d0_4508,RIfca3760_6882,RIe2105d0_4476,RIfc97988_6747,RIe20d8d0_4444,RIe20abd0_4412,
        RIe207ed0_4380,RIfceb5b0_7700,RIfcddbb8_7545,RIe202a70_4320,RIe200e50_4300,RIfc73d30_6340,RIfcaf100_7014,RIfc71468_6311,RIfcdcad8_7533,RIfcdda50_7544,
        RIfca8620_6938,RIe1fcf08_4255,RIe1fbcc0_4242,RIfc6c008_6251,RIfcdd1e0_7538,RIfca9700_6950,RIfca92c8_6947,RIfcce5a0_7370,RIfc6ba68_6247,RIfc6f410_6288,
        RIe1fa640_4226,RIfcce000_7366,RIfc53918_5973,RIfcce708_7371,RIe1f5bb8_4173,RIf1535f0_5408,RIf151e08_5391,RIfc72db8_6329,RIe1f3890_4148,RIf14fc48_5367,
        RIfc72c50_6328,RIfc73e98_6341,RIe1ee598_4089,RIe1ebe38_4061,RIe1e9138_4029,RIe1e6438_3997,RIe1e3738_3965,RIe1e0a38_3933,RIe1ddd38_3901,RIe1db038_3869,
        RIe1d8338_3837,RIe1d2938_3773,RIe1cfc38_3741,RIe1ccf38_3709,RIe1ca238_3677,RIe1c7538_3645,RIe1c4838_3613,RIe1c1b38_3581,RIe1bee38_3549,RIfcb8a48_7123,
        RIfcb84a8_7119,RIe1b9870_3488,RIe1b7818_3465,RIfc85940_6542,RIfc9e198_6821,RIfeac140_8274,RIe1b42a8_3427,RIfc518c0_5950,RIfc838e8_6519,RIfe884e8_7895,
        RIe1b1008_3391,RIfcc5900_7270,RIfc82ad8_6509,RIe1ac9b8_3341,RIfe88650_7896,RIe1a9178_3301,RIe1a6478_3269,RIe1a3778_3237,RIe1a0a78_3205,RIe18cf78_2981,
        RIe179478_2757,RIe226dd0_4732,RIe21b9d0_4604,RIe2051d0_4348,RIe1ff230_4280,RIe1f85e8_4203,RIe1f1130_4120,RIe1d5638_3805,RIe1bc138_3517,RIe1aefb0_3368,
        RIe1715e8_2667,RIdec5f18_716,RIdec3218_684,RIee20350_4825,RIdec0518_652,RIee1f6a8_4816,RIdebd818_620,RIdebab18_588,RIdeb7e18_556,RIfce4da0_7626,
        RIdeb2418_492,RIfcea908_7691,RIdeaf718_460,RIfce20a0_7594,RIdeabe60_428,RIdea5560_396,RIde9ec60_364,RIfce6420_7642,RIee1c2a0_4779,RIfc75950_6360,
        RIee1ad88_4764,RIde920f0_302,RIfea4148_8211,RIfeaa688_8255,RIfea3fe0_8210,RIde82790_226,RIfc6f848_6291,RIfc5dc38_6089,RIfc76b98_6373,RIfcae2f0_7004,
        RIe16c020_2606,RIe16a130_2584,RIe1687e0_2566,RIe165f18_2537,RIe163218_2505,RIfcadd50_7000,RIe160518_2473,RIfc55268_5991,RIe15d818_2441,RIe157e18_2377,
        RIe155118_2345,RIfc45548_5811,RIe152418_2313,RIfc498c8_5859,RIe14f718_2281,RIfcbda70_7180,RIe14ca18_2249,RIe149d18_2217,RIe147018_2185,RIee34828_5056,
        RIee33748_5044,RIee32668_5032,RIee31588_5020,RIe1418e8_2123,RIe13f458_2097,RIdf3d360_2073,RIdf3aed0_2047,RIfc526d0_5960,RIfc42848_5779,RIfcae9f8_7009,
        RIfcb7260_7106,RIfea42b0_8212,RIdf33ce8_1966,RIdf31b28_1942,RIdf2fc38_1920,RIee2c3f8_4962,RIfc4cfa0_5898,RIfc572c0_6014,RIfc4f430_5924,RIfea3e78_8209,
        RIdf28a50_1839,RIdf26b60_1817,RIdf250a8_1798,RIfc9b600_6790,RIfcb9df8_7137,RIdf23320_1777,RIfc86318_6549,RIfeabfd8_8273,RIdf201e8_1742,RIdf1b5f8_1688,
        RIdf19ca8_1670,RIdf17ae8_1646,RIdf14de8_1614,RIdf120e8_1582,RIdf0f3e8_1550,RIdf0c6e8_1518,RIdf099e8_1486,RIdf06ce8_1454,RIdf03fe8_1422,RIdefe5e8_1358,
        RIdefb8e8_1326,RIdef8be8_1294,RIdef5ee8_1262,RIdef31e8_1230,RIdef04e8_1198,RIdeed7e8_1166,RIdeeaae8_1134,RIfc89018_6581,RIfcc54c8_7267,RIfc89180_6582,
        RIfc4b380_5878,RIdee53b8_1072,RIdee34c8_1050,RIfea3d10_8208,RIdedf148_1002,RIfcae188_7003,RIfc4b0b0_5876,RIfc74870_6348,RIfce4968_7623,RIdeda288_946,
        RIded7c90_919,RIded5da0_897,RIded3640_869,RIded1318_844,RIdece618_812,RIdecb918_780,RIdec8c18_748,RIdeb5118_524,RIde98360_332,RIe16ed20_2638,
        RIe15ab18_2409,RIe144318_2153,RIdf38d10_2023,RIdf2d370_1891,RIdf1dbf0_1715,RIdf012e8_1390,RIdee7de8_1102,RIdedcb50_975,RIde7e2a8_205,RIe19e1b0_3176,
        RIe19b4b0_3144,RIfc9cf50_6808,RIe1987b0_3112,RIfc87290_6560,RIe195ab0_3080,RIe192db0_3048,RIe1900b0_3016,RIe18a6b0_2952,RIe1879b0_2920,RIfc842c0_6526,
        RIe184cb0_2888,RIfc83a50_6520,RIe181fb0_2856,RIe17f2b0_2824,RIe17c5b0_2792,RIfc9d0b8_6809,RIfc9e030_6820,RIe177420_2734,RIe176340_2722,RIfc4f700_5926,
        RIfcc4820_7258,RIfc4fb38_5929,RIfce8040_7662,RIee3c6b8_5146,RIee3b308_5132,RIfc812f0_6492,RIe174180_2698,RIfcd3028_7423,RIfc7f400_6470,RIfc46a60_5826,
        RIfc472d0_5832,RIf16cc58_5697,RIe224508_4703,RIfc7d3a8_6447,RIe221808_4671,RIfc97c58_6749,RIe21eb08_4639,RIe219108_4575,RIe216408_4543,RIfcdbe30_7524,
        RIe213708_4511,RIf169580_5658,RIe210a08_4479,RIfca4570_6892,RIe20dd08_4447,RIe20b008_4415,RIe208308_4383,RIfc7b080_6422,RIfc59cf0_6044,RIfea9b48_8247,
        RIfea4418_8213,RIfc79cd0_6408,RIfcd19a8_7407,RIfcc81c8_7299,RIf162230_5576,RIf160778_5557,RIf15e888_5535,RIfea4580_8214,RIfea46e8_8215,RIfc77f48_6387,
        RIfc41fd8_5773,RIf15aaa8_5491,RIfc7c430_6436,RIf159158_5473,RIf157f10_5460,RIfcae890_7008,RIe1faa78_4229,RIfc4a840_5870,RIfc4ed28_5919,RIfce0e58_7581,
        RIe1f5ff0_4176,RIf153758_5409,RIf151f70_5392,RIfccb468_7335,RIe1f3cc8_4151,RIfc68ed0_6216,RIfc6d250_6264,RIfca9ca0_6954,RIe1ee9d0_4092,RIe1ec270_4064,
        RIe1e9570_4032,RIe1e6870_4000,RIe1e3b70_3968,RIe1e0e70_3936,RIe1de170_3904,RIe1db470_3872,RIe1d8770_3840,RIe1d2d70_3776,RIe1d0070_3744,RIe1cd370_3712,
        RIe1ca670_3680,RIe1c7970_3648,RIe1c4c70_3616,RIe1c1f70_3584,RIe1bf270_3552,RIfc784e8_6391,RIfcbef88_7195,RIe1b9ca8_3491,RIe1b7ae8_3467,RIfcc20c0_7230,
        RIfca6190_6912,RIe1b5928_3443,RIe1b4410_3428,RIfcb81d8_7117,RIfcc5090_7264,RIe1b2d90_3412,RIe1b1440_3394,RIfcd5350_7448,RIfcb9588_7131,RIe1acc88_3343,
        RIe1ab4a0_3326,RIe1a95b0_3304,RIe1a68b0_3272,RIe1a3bb0_3240,RIe1a0eb0_3208,RIe18d3b0_2984,RIe1798b0_2760,RIe227208_4735,RIe21be08_4607,RIe205608_4351,
        RIe1ff668_4283,RIe1f8a20_4206,RIe1f1568_4123,RIe1d5a70_3808,RIe1bc570_3520,RIe1af3e8_3371,RIe171a20_2670,RIdec5db0_715,RIdec30b0_683,RIee201e8_4824,
        RIdec03b0_651,RIfcaf538_7017,RIdebd6b0_619,RIdeba9b0_587,RIdeb7cb0_555,RIfc40fe8_5765,RIdeb22b0_491,RIfcd08c8_7395,RIdeaf5b0_459,RIee1dd58_4798,
        RIdeabb18_427,RIdea5218_395,RIde9e918_363,RIee1d218_4790,RIfcedd10_7728,RIfce62b8_7641,RIfcc92a8_7311,RIde91da8_301,RIde8e928_285,RIde8a788_265,
        RIde865e8_245,RIde82448_225,RIfea1448_8179,RIfc750e0_6354,RIfcc19b8_7225,RIfced8d8_7725,RIfec5eb0_8372,RIe169fc8_2583,RIe168678_2565,RIe165db0_2536,
        RIe1630b0_2504,RIfccfc20_7386,RIe1603b0_2472,RIee365b0_5077,RIe15d6b0_2440,RIe157cb0_2376,RIe154fb0_2344,RIfea1718_8181,RIe1522b0_2312,RIee35200_5063,
        RIe14f5b0_2280,RIfcb0348_7027,RIe14c8b0_2248,RIe149bb0_2216,RIe146eb0_2184,RIfc73790_6336,RIfcdf238_7561,RIee32500_5031,RIfc94f58_6717,RIe141780_2122,
        RIe13f2f0_2096,RIfec5be0_8370,RIdf3ad68_2046,RIfea15b0_8180,RIfc5fb28_6111,RIfcae728_7007,RIfc74438_6345,RIdf36178_1992,RIdf33b80_1965,RIdf319c0_1941,
        RIdf2fad0_1919,RIee2c290_4961,RIee2a940_4943,RIfc70658_6301,RIfc704f0_6300,RIdf2aaa8_1862,RIdf288e8_1838,RIdf269f8_1816,RIdf24f40_1797,RIfc64b50_6168,
        RIfccaa90_7328,RIdf231b8_1776,RIfcad4e0_6994,RIdf21ca0_1761,RIfeaad90_8260,RIdf1b490_1687,RIdf19b40_1669,RIdf17980_1645,RIdf14c80_1613,RIdf11f80_1581,
        RIdf0f280_1549,RIdf0c580_1517,RIdf09880_1485,RIdf06b80_1453,RIdf03e80_1421,RIdefe480_1357,RIdefb780_1325,RIdef8a80_1293,RIdef5d80_1261,RIdef3080_1229,
        RIdef0380_1197,RIdeed680_1165,RIdeea980_1133,RIfc595e8_6039,RIfcac568_6983,RIfcccf20_7354,RIfccd358_7357,RIdee5250_1071,RIfea7f28_8227,RIdee11a0_1025,
        RIfea12e0_8178,RIfc679b8_6201,RIee22510_4849,RIfc6dd90_6272,RIfc6cb48_6259,RIdeda120_945,RIded7b28_918,RIded5c38_896,RIfec5d48_8371,RIded11b0_843,
        RIdece4b0_811,RIdecb7b0_779,RIdec8ab0_747,RIdeb4fb0_523,RIde98018_331,RIe16ebb8_2637,RIe15a9b0_2408,RIe1441b0_2152,RIdf38ba8_2022,RIdf2d208_1890,
        RIdf1da88_1714,RIdf01180_1389,RIdee7c80_1101,RIdedc9e8_974,RIde7df60_204,RIe19e048_3175,RIe19b348_3143,RIfcc3ce0_7250,RIe198648_3111,RIfc7efc8_6467,
        RIe195948_3079,RIe192c48_3047,RIe18ff48_3015,RIe18a548_2951,RIe187848_2919,RIfc46790_5824,RIe184b48_2887,RIfc98d38_6761,RIe181e48_2855,RIe17f148_2823,
        RIe17c448_2791,RIfcb5d48_7091,RIfc995a8_6767,RIfc9a3b8_6777,RIe1761d8_2721,RIfc54188_5979,RIfcd2bf0_7420,RIfc8b778_6609,RIfc7dee8_6455,RIee3c550_5145,
        RIfc8c420_6618,RIee3a0c0_5119,RIfeaba38_8269,RIfc46628_5823,RIfcbc288_7163,RIf16e710_5716,RIfc8fdc8_6659,RIfc48c20_5850,RIe2243a0_4702,RIfca0358_6845,
        RIe2216a0_4670,RIfc9a688_6779,RIe21e9a0_4638,RIe218fa0_4574,RIe2162a0_4542,RIfc456b0_5812,RIe2135a0_4510,RIf169418_5657,RIe2108a0_4478,RIfc8bfe8_6615,
        RIe20dba0_4446,RIe20aea0_4414,RIe2081a0_4382,RIfc8c9c0_6622,RIfc7f568_6471,RIe202d40_4322,RIe201120_4302,RIfce2910_7600,RIfc487e8_5847,RIfc46d30_5828,
        RIfc992d8_6765,RIfca2680_6870,RIfc44a08_5803,RIe1fd1d8_4257,RIe1fbf90_4244,RIfc580d0_6024,RIfcbdbd8_7181,RIfc8dd70_6636,RIfce01b0_7572,RIfc7bbc0_6430,
        RIfc90368_6663,RIfc7b8f0_6428,RIe1fa910_4228,RIfcd8b90_7488,RIfc43ec8_5795,RIfc7b788_6427,RIe1f5e88_4175,RIfc7b350_6424,RIfc90d40_6670,RIfca3490_6880,
        RIe1f3b60_4150,RIfc91010_6672,RIfcdb728_7519,RIfcd8758_7485,RIe1ee868_4091,RIe1ec108_4063,RIe1e9408_4031,RIe1e6708_3999,RIe1e3a08_3967,RIe1e0d08_3935,
        RIe1de008_3903,RIe1db308_3871,RIe1d8608_3839,RIe1d2c08_3775,RIe1cff08_3743,RIe1cd208_3711,RIe1ca508_3679,RIe1c7808_3647,RIe1c4b08_3615,RIe1c1e08_3583,
        RIe1bf108_3551,RIf14cf48_5335,RIfc78d58_6397,RIe1b9b40_3490,RIfec5910_8368,RIfc78a88_6395,RIfcd51e8_7447,RIe1b57c0_3442,RIfea1010_8176,RIf1492d0_5292,
        RIfec5a78_8369,RIe1b2c28_3411,RIe1b12d8_3393,RIfec5640_8366,RIf146a08_5263,RIfec57a8_8367,RIfea1178_8177,RIe1a9448_3303,RIe1a6748_3271,RIe1a3a48_3239,
        RIe1a0d48_3207,RIe18d248_2983,RIe179748_2759,RIe2270a0_4734,RIe21bca0_4606,RIe2054a0_4350,RIe1ff500_4282,RIe1f88b8_4205,RIe1f1400_4122,RIe1d5908_3807,
        RIe1bc408_3519,RIe1af280_3370,RIe1718b8_2669,RIdec6350_719,RIdec3650_687,RIfcaf3d0_7016,RIdec0950_655,RIfc6a280_6230,RIdebdc50_623,RIdebaf50_591,
        RIdeb8250_559,RIfc42f50_5784,RIdeb2850_495,RIfc981f8_6753,RIdeafb50_463,RIfc8c6f0_6620,RIdeac838_431,RIdea5f38_399,RIde9f638_367,RIee1d4e8_4792,
        RIfcda648_7507,RIfcc6440_7278,RIfcd5620_7450,RIde92ac8_305,RIfea34a0_8202,RIfea31d0_8200,RIfea3338_8201,RIfcb6b58_7101,RIfcb6888_7099,RIfc9dd60_6818,
        RIee19708_4748,RIfc50c18_5941,RIe16c458_2609,RIfc80a80_6486,RIfec62e8_8375,RIe166350_2540,RIe163650_2508,RIee37d98_5094,RIe160950_2476,RIfcaa678_6961,
        RIe15dc50_2444,RIe158250_2380,RIe155550_2348,RIfea3ba8_8207,RIe152850_2316,RIee35638_5066,RIe14fb50_2284,RIfc62f30_6148,RIe14ce50_2252,RIe14a150_2220,
        RIe147450_2188,RIfc97f28_6751,RIfc89888_6587,RIfc8f558_6653,RIfc52838_5961,RIe141bb8_2125,RIe13f890_2100,RIdf3d798_2076,RIdf3b308_2050,RIee30a48_5012,
        RIfc568e8_6007,RIee2e9f0_4989,RIee2dbe0_4979,RIdf365b0_1995,RIfea38d8_8205,RIfea3a40_8206,RIdf2ff08_1922,RIee2c6c8_4964,RIee2ac10_4945,RIee29590_4929,
        RIee28348_4916,RIdf2ad78_1864,RIdf28e88_1842,RIfea3608_8203,RIfea3770_8204,RIfcc0d10_7216,RIfc75c20_6362,RIfca50b0_6900,RIfc74e10_6352,RIfcc9410_7312,
        RIdf20620_1745,RIfc73628_6335,RIdf1a0e0_1673,RIdf17f20_1649,RIdf15220_1617,RIdf12520_1585,RIdf0f820_1553,RIdf0cb20_1521,RIdf09e20_1489,RIdf07120_1457,
        RIdf04420_1425,RIdefea20_1361,RIdefbd20_1329,RIdef9020_1297,RIdef6320_1265,RIdef3620_1233,RIdef0920_1201,RIdeedc20_1169,RIdeeaf20_1137,RIfcab8c0_6974,
        RIfc7c598_6437,RIfc5beb0_6068,RIfc58ee0_6034,RIdee5688_1074,RIdee3798_1052,RIdee15d8_1028,RIdedf580_1005,RIfcb3048_7059,RIfc72ae8_6327,RIfca3d00_6886,
        RIfcb6450_7096,RIdeda558_948,RIded7f60_921,RIfea3068_8199,RIded3a78_872,RIded1750_847,RIdecea50_815,RIdecbd50_783,RIdec9050_751,RIdeb5550_527,
        RIde98d38_335,RIe16f158_2641,RIe15af50_2412,RIe144750_2156,RIdf39148_2026,RIdf2d7a8_1894,RIdf1e028_1718,RIdf01720_1393,RIdee8220_1105,RIdedcf88_978,
        RIde7ec80_208,RIe19e5e8_3179,RIe19b8e8_3147,RIfca84b8_6937,RIe198be8_3115,RIfc846f8_6529,RIe195ee8_3083,RIe1931e8_3051,RIe1904e8_3019,RIe18aae8_2955,
        RIe187de8_2923,RIfce2be0_7602,RIe1850e8_2891,RIfc8e310_6640,RIe1823e8_2859,RIe17f6e8_2827,RIe17c9e8_2795,RIfcd1570_7404,RIfccc278_7345,RIf1404c8_5191,
        RIfea2d98_8197,RIfcc1b20_7226,RIfc60398_6117,RIee3e5a8_5168,RIee3da68_5160,RIfc642e0_6162,RIfca7f18_6933,RIee3a228_5120,RIfec6180_8374,RIfca9598_6949,
        RIfc5c720_6074,RIfc6bea0_6250,RIfccaec8_7331,RIfc44cd8_5805,RIe224940_4706,RIfcb6180_7094,RIe221c40_4674,RIfc55ad8_5997,RIe21ef40_4642,RIe219540_4578,
        RIe216840_4546,RIfc4dc48_5907,RIe213b40_4514,RIfcdcf10_7536,RIe210e40_4482,RIfcab1b8_6969,RIe20e140_4450,RIe20b440_4418,RIe208740_4386,RIfce3720_7610,
        RIfc64178_6161,RIe203178_4325,RIe201558_4305,RIfcd2ec0_7422,RIf164828_5603,RIfc7f838_6473,RIf162398_5577,RIfcc9c80_7318,RIfca8bc0_6942,RIfea2ac8_8195,
        RIfea2c30_8196,RIfc59318_6037,RIfc4f160_5922,RIf15ac10_5492,RIfcebf88_7707,RIfcbb040_7150,RIfca1870_6860,RIfc93d10_6704,RIe1faeb0_4232,RIf1565c0_5442,
        RIf155a80_5434,RIfc45c50_5816,RIe1f6428_4179,RIfccdbc8_7363,RIfcccae8_7351,RIfca6cd0_6920,RIfec6018_8373,RIfc64010_6160,RIfc434f0_5788,RIfc4c028_5887,
        RIe1eee08_4095,RIe1ec6a8_4067,RIe1e99a8_4035,RIe1e6ca8_4003,RIe1e3fa8_3971,RIe1e12a8_3939,RIe1de5a8_3907,RIe1db8a8_3875,RIe1d8ba8_3843,RIe1d31a8_3779,
        RIe1d04a8_3747,RIe1cd7a8_3715,RIe1caaa8_3683,RIe1c7da8_3651,RIe1c50a8_3619,RIe1c23a8_3587,RIe1bf6a8_3555,RIfc63908_6155,RIfc6bd38_6249,RIe1ba0e0_3494,
        RIe1b7f20_3470,RIfc66fe0_6194,RIfc92ac8_6691,RIe1b5d60_3446,RIfea2f00_8198,RIfc9bfd8_6797,RIfc50d80_5942,RIe1b31c8_3415,RIe1b1878_3397,RIfc4df18_5909,
        RIfc9d658_6813,RIe1ad0c0_3346,RIe1ab8d8_3329,RIe1a99e8_3307,RIe1a6ce8_3275,RIe1a3fe8_3243,RIe1a12e8_3211,RIe18d7e8_2987,RIe179ce8_2763,RIe227640_4738,
        RIe21c240_4610,RIe205a40_4354,RIe1ffaa0_4286,RIe1f8e58_4209,RIe1f19a0_4126,RIe1d5ea8_3811,RIe1bc9a8_3523,RIe1af820_3374,RIe171e58_2673,RIdec61e8_718,
        RIdec34e8_686,RIee20620_4827,RIdec07e8_654,RIfc4b7b8_5881,RIdebdae8_622,RIdebade8_590,RIdeb80e8_558,RIfc41150_5766,RIdeb26e8_494,RIfc87830_6564,
        RIdeaf9e8_462,RIee1dec0_4799,RIdeac4f0_430,RIdea5bf0_398,RIde9f2f0_366,RIee1d380_4791,RIfc77c78_6385,RIfc84f68_6535,RIfc6ff50_6296,RIde92780_304,
        RIde8efb8_287,RIde8ae18_267,RIde86c78_247,RIee1a680_4759,RIee19f78_4754,RIfcd7240_7470,RIfcbeb50_7192,RIfc76328_6367,RIe16c2f0_2608,RIee388d8_5102,
        RIfea20f0_8188,RIe1661e8_2539,RIe1634e8_2507,RIee37c30_5093,RIe1607e8_2475,RIfce7500_7654,RIe15dae8_2443,RIe1580e8_2379,RIe1553e8_2347,RIfc3f698_5747,
        RIe1526e8_2315,RIee354d0_5065,RIe14f9e8_2283,RIfc83e88_6523,RIe14cce8_2251,RIe149fe8_2219,RIe1472e8_2187,RIfcea4d0_7688,RIfcb7ad0_7112,RIfc695d8_6221,
        RIfc51a28_5951,RIe141a50_2124,RIe13f728_2099,RIdf3d630_2075,RIdf3b1a0_2049,RIfca9e08_6955,RIee2fda0_5003,RIfc88a78_6577,RIee2da78_4978,RIdf36448_1994,
        RIdf33fb8_1968,RIdf31df8_1944,RIfea2258_8189,RIee2c560_4963,RIee2aaa8_4944,RIee29428_4928,RIee281e0_4915,RIdf2ac10_1863,RIdf28d20_1841,RIfea27f8_8193,
        RIfea2960_8194,RIfcdabe8_7511,RIfca08f8_6849,RIfc8b1d8_6605,RIfc49058_5853,RIfca0a60_6850,RIdf204b8_1744,RIfc99cb0_6772,RIdf19f78_1672,RIdf17db8_1648,
        RIdf150b8_1616,RIdf123b8_1584,RIdf0f6b8_1552,RIdf0c9b8_1520,RIdf09cb8_1488,RIdf06fb8_1456,RIdf042b8_1424,RIdefe8b8_1360,RIdefbbb8_1328,RIdef8eb8_1296,
        RIdef61b8_1264,RIdef34b8_1232,RIdef07b8_1200,RIdeedab8_1168,RIdeeadb8_1136,RIfcd1f48_7411,RIfc57f68_6023,RIfcbe2e0_7186,RIfcd8fc8_7491,RIdee5520_1073,
        RIfea2690_8192,RIdee1470_1027,RIdedf418_1004,RIfc57b30_6020,RIfcb35e8_7063,RIfcbd7a0_7178,RIfc91178_6673,RIfea2528_8191,RIded7df8_920,RIfea23c0_8190,
        RIded3910_871,RIded15e8_846,RIdece8e8_814,RIdecbbe8_782,RIdec8ee8_750,RIdeb53e8_526,RIde989f0_334,RIe16eff0_2640,RIe15ade8_2411,RIe1445e8_2155,
        RIdf38fe0_2025,RIdf2d640_1893,RIdf1dec0_1717,RIdf015b8_1392,RIdee80b8_1104,RIdedce20_977,RIde7e938_207,RIe19e480_3178,RIe19b780_3146,RIfccc980_7350,
        RIe198a80_3114,RIfcc1148_7219,RIe195d80_3082,RIe193080_3050,RIe190380_3018,RIe18a980_2954,RIe187c80_2922,RIfcb2ee0_7058,RIe184f80_2890,RIfc615e0_6130,
        RIe182280_2858,RIe17f580_2826,RIe17c880_2794,RIfc69038_6217,RIfc4c898_5893,RIfc6f2a8_6287,RIe1764a8_2723,RIfcad0a8_6991,RIfc6adc0_6238,RIfc70388_6299,
        RIfea1b50_8184,RIfea1f88_8187,RIfc56e88_6011,RIfea1cb8_8185,RIe174450_2700,RIfc60d70_6124,RIfc6a820_6234,RIfea1e20_8186,RIf16d798_5705,RIfc40bb0_5762,
        RIe2247d8_4705,RIfc77138_6377,RIe221ad8_4673,RIfcd7d80_7478,RIe21edd8_4641,RIe2193d8_4577,RIe2166d8_4545,RIfc40070_5754,RIe2139d8_4513,RIf169850_5660,
        RIe210cd8_4481,RIfcc1580_7222,RIe20dfd8_4449,RIe20b2d8_4417,RIe2085d8_4385,RIfcd0058_7389,RIfc749d8_6349,RIe203010_4324,RIe2013f0_4304,RIfc60230_6116,
        RIfc60668_6119,RIfcaf970_7020,RIfc45818_5813,RIf160a48_5559,RIf15eb58_5537,RIfea1880_8182,RIfea19e8_8183,RIfc72110_6320,RIfc49b98_5861,RIfcca0b8_7321,
        RIfc71738_6313,RIfc4ca00_5894,RIfc71030_6308,RIfcde428_7551,RIe1fad48_4231,RIfc70bf8_6305,RIfc63a70_6156,RIfca7db0_6932,RIe1f62c0_4178,RIfcada80_6998,
        RIfc6fde8_6295,RIfc6f578_6289,RIe1f3f98_4153,RIfcde158_7549,RIfcad378_6993,RIfc65f00_6182,RIe1eeca0_4094,RIe1ec540_4066,RIe1e9840_4034,RIe1e6b40_4002,
        RIe1e3e40_3970,RIe1e1140_3938,RIe1de440_3906,RIe1db740_3874,RIe1d8a40_3842,RIe1d3040_3778,RIe1d0340_3746,RIe1cd640_3714,RIe1ca940_3682,RIe1c7c40_3650,
        RIe1c4f40_3618,RIe1c2240_3586,RIe1bf540_3554,RIfc69308_6219,RIfccba08_7339,RIe1b9f78_3493,RIe1b7db8_3469,RIfccd628_7359,RIfc69740_6222,RIe1b5bf8_3445,
        RIe1b4578_3429,RIfccf950_7384,RIf148088_5279,RIe1b3060_3414,RIe1b1710_3396,RIfc9f818_6837,RIfcb9c90_7136,RIe1acf58_3345,RIe1ab770_3328,RIe1a9880_3306,
        RIe1a6b80_3274,RIe1a3e80_3242,RIe1a1180_3210,RIe18d680_2986,RIe179b80_2762,RIe2274d8_4737,RIe21c0d8_4609,RIe2058d8_4353,RIe1ff938_4285,RIe1f8cf0_4208,
        RIe1f1838_4125,RIe1d5d40_3810,RIe1bc840_3522,RIe1af6b8_3373,RIe171cf0_2672;
output R_58_102f1b78,R_59_be1fc68,R_5a_10279198,R_5b_102299e8,R_5c_101d0448,R_5d_f7f82f0,R_5e_be21600,R_5f_f7fa5b8,R_60_1027d530,
        R_61_10205ae8,R_62_10283510,R_63_f82b578,R_64_ace4e68,R_65_f8204e0,R_66_1027a0b0,R_67_1022dc30,R_68_102478a8,R_69_10286f78,R_6a_f7edd80,
        R_6b_101c3628,R_6c_f7fbe00,R_6d_f7ce9f8,R_6e_f7c8830,R_6f_101ffc68,R_70_f7d4000,R_71_acee958,R_72_94046c0,R_73_101ee420,R_74_102eb268,
        R_75_b320c50,R_76_ad80a90,R_77_1027fd48,R_78_f7ce4b8,R_79_ad77048,R_7a_102a6ae0,R_7b_f7e4c78,R_7c_e2a6ce0,R_7d_101e86e0,R_7e_e2a9cc8,
        R_7f_10292be0,R_80_b33cde8,R_81_101e2908,R_82_102e9780,R_83_f8157a0,R_84_f819358,R_85_ace8b70,R_86_be142b0,R_87_f81b770,R_88_b330278,
        R_89_f7fe9f8,R_8a_101cf488,R_8b_f8225c0,R_8c_101d4738,R_8d_101c4000,R_8e_101fe960,R_8f_102a0330,R_90_f7f4bd0,R_91_1023e5a8,R_92_10248da8,
        R_93_be2c938,R_94_f7f5458,R_95_f7c6808,R_96_be316a8,R_97_e2a0328,R_98_be2d850,R_99_10217db0,R_9a_f7ec340,R_9b_be23ec0,R_9c_101d4540,
        R_9d_f800828,R_9e_102970c8,R_9f_10221de0,R_a0_ad8d568,R_a1_be4eb58,R_a2_f7c5500,R_a3_ad88f30,R_a4_f82f088,R_a5_f7dcbc8,R_a6_10292940,
        R_a7_be138d8,R_a8_acee418,R_a9_ad84450,R_aa_be10838,R_ab_be31fd8,R_ac_acdaef0,R_ad_acea908,R_ae_101f8830,R_af_f7dec98,R_b0_101e2c50,
        R_b1_f801b30,R_b2_be16e00,R_b3_102e3cf0,R_b4_10291788;

wire \8308_N$1 , \8309_N$4 , \8310_N$5 , \8311_N$6 , \8312_N$8 , \8313_N$9 , \8314_N$10 , \8315_N$11 , \8316_N$15 ,
         \8317_N$16 , \8318_N$17 , \8319_N$18 , \8320_N$21 , \8321_N$22 , \8322_N$23 , \8323_N$24 , \8324_N$25 , \8325_N$26 , \8326_N$29 ,
         \8327_N$30 , \8328_N$31 , \8329_N$32 , \8330_N$33 , \8331_N$34 , \8332_N$35 , \8333_N$36 , \8334_N$37 , \8335_N$38 , \8336_N$39 ,
         \8337_N$40 , \8338_N$41 , \8339_N$42 , \8340_N$43 , \8341_N$44 , \8342_N$45 , \8343_N$46 , \8344_N$47 , \8345_N$48 , \8346_N$49 ,
         \8347_N$50 , \8348_N$51 , \8349_N$52 , \8350_N$53 , \8351_N$54 , \8352_N$55 , \8353_N$56 , \8354_N$57 , \8355_N$58 , \8356_N$59 ,
         \8357_N$60 , \8358_N$61 , \8359_N$62 , \8360_N$63 , \8361_N$64 , \8362_N$65 , \8363_N$66 , \8364_N$67 , \8365_N$68 , \8366_N$69 ,
         \8367_N$70 , \8368_N$71 , \8369_N$72 , \8370_N$73 , \8371_N$74 , \8372_N$75 , \8373_N$76 , \8374_N$77 , \8375_N$78 , \8376_N$79 ,
         \8377_N$80 , \8378_N$81 , \8379_N$82 , \8380_N$83 , \8381_N$84 , \8382_N$85 , \8383_N$86 , \8384_N$87 , \8385_N$88 , \8386_N$89 ,
         \8387_N$90 , \8388_N$91 , \8389_N$92 , \8390_N$93 , \8391_N$94 , \8392_N$95 , \8393_N$96 , \8394_N$97 , \8395_N$98 , \8396_N$99 ,
         \8397_N$100 , \8398_N$101 , \8399_N$102 , \8400_N$103 , \8401_N$104 , \8402_N$105 , \8403_N$106 , \8404_N$107 , \8405_N$108 , \8406_N$109 ,
         \8407_N$110 , \8408_N$111 , \8409_N$112 , \8410_N$113 , \8411_N$114 , \8412_N$115 , \8413_N$116 , \8414_N$117 , \8415_N$118 , \8416_N$119 ,
         \8417_N$120 , \8418_N$121 , \8419_N$122 , \8420_N$123 , \8421_N$124 , \8422_N$125 , \8423_N$126 , \8424_N$127 , \8425_N$128 , \8426_N$129 ,
         \8427_N$130 , \8428_N$131 , \8429_N$132 , \8430_N$133 , \8431_N$134 , \8432_N$135 , \8433_N$136 , \8434_N$137 , \8435_N$138 , \8436_N$139 ,
         \8437_N$140 , \8438_N$141 , \8439_N$142 , \8440_N$143 , \8441_N$144 , \8442_N$145 , \8443_N$146 , \8444_N$147 , \8445_N$148 , \8446_N$149 ,
         \8447_N$150 , \8448_N$151 , \8449_N$152 , \8450_N$153 , \8451_N$154 , \8452_N$155 , \8453_N$156 , \8454_N$157 , \8455_N$158 , \8456_N$159 ,
         \8457_N$160 , \8458_N$161 , \8459_N$162 , \8460_N$163 , \8461_N$164 , \8462_N$165 , \8463_N$166 , \8464_N$167 , \8465_N$168 , \8466_N$169 ,
         \8467_N$170 , \8468_N$171 , \8469_N$172 , \8470_N$173 , \8471_N$174 , \8472_N$175 , \8473_N$176 , \8474_N$177 , \8475_N$178 , \8476_N$179 ,
         \8477_N$180 , \8478_N$181 , \8479_N$182 , \8480_N$183 , \8481_N$184 , \8482_N$185 , \8483_N$186 , \8484_N$187 , \8485_N$188 , \8486_N$189 ,
         \8487_N$190 , \8488_N$191 , \8489_N$192 , \8490_N$193 , \8491_N$194 , \8492_N$195 , \8493_N$196 , \8494_N$197 , \8495_N$198 , \8496_N$199 ,
         \8497_N$200 , \8498_N$201 , \8499_N$202 , \8500_N$203 , \8501_N$204 , \8502_N$205 , \8503_N$206 , \8504_N$207 , \8505_N$208 , \8506_N$209 ,
         \8507_N$210 , \8508_N$211 , \8509_N$212 , \8510_N$213 , \8511_N$214 , \8512_N$215 , \8513_N$216 , \8514_N$219 , \8515_N$220 , \8516_N$221 ,
         \8517_N$222 , \8518_N$223 , \8519_N$224 , \8520_N$226 , \8521_N$227 , \8522_N$228 , \8523_N$229 , \8524_N$230 , \8525_N$231 , \8526_N$232 ,
         \8527_N$233 , \8528_N$234 , \8529_N$235 , \8530_N$236 , \8531_N$237 , \8532_N$238 , \8533_N$239 , \8534_N$240 , \8535_N$241 , \8536_N$242 ,
         \8537_N$243 , \8538_N$244 , \8539_N$245 , \8540_N$246 , \8541_N$247 , \8542_N$248 , \8543_N$249 , \8544_N$250 , \8545_N$251 , \8546_N$252 ,
         \8547_N$253 , \8548_N$254 , \8549_N$255 , \8550_N$256 , \8551_N$257 , \8552_N$258 , \8553_N$259 , \8554_N$260 , \8555_N$261 , \8556_N$262 ,
         \8557_N$263 , \8558_N$264 , \8559_N$265 , \8560_N$266 , \8561_N$267 , \8562_N$268 , \8563_N$269 , \8564_N$270 , \8565_N$271 , \8566_N$272 ,
         \8567_N$273 , \8568_N$274 , \8569_N$275 , \8570_N$276 , \8571_N$277 , \8572_N$278 , \8573_N$279 , \8574_N$280 , \8575_N$281 , \8576_N$282 ,
         \8577_N$283 , \8578_N$284 , \8579_N$285 , \8580_N$286 , \8581_N$287 , \8582_N$288 , \8583_N$289 , \8584_N$290 , \8585_N$291 , \8586_N$292 ,
         \8587_N$293 , \8588_N$294 , \8589_N$295 , \8590_N$296 , \8591_N$297 , \8592_N$298 , \8593_N$299 , \8594_N$300 , \8595_N$301 , \8596_N$302 ,
         \8597_N$303 , \8598_N$304 , \8599_N$305 , \8600_N$306 , \8601_N$307 , \8602_N$308 , \8603_N$309 , \8604_N$310 , \8605_N$311 , \8606_N$312 ,
         \8607_N$313 , \8608_N$314 , \8609_N$315 , \8610_N$316 , \8611_N$317 , \8612_N$318 , \8613_N$319 , \8614_N$320 , \8615_N$321 , \8616_N$322 ,
         \8617_N$323 , \8618_N$324 , \8619_N$325 , \8620_N$326 , \8621_N$327 , \8622_N$328 , \8623_N$329 , \8624_N$330 , \8625_N$331 , \8626_N$332 ,
         \8627_N$333 , \8628_N$334 , \8629_N$335 , \8630_N$336 , \8631_N$337 , \8632_N$338 , \8633_N$339 , \8634_N$340 , \8635_N$341 , \8636_N$342 ,
         \8637_N$343 , \8638_N$344 , \8639_N$345 , \8640_N$346 , \8641_N$347 , \8642_N$348 , \8643_N$349 , \8644_N$350 , \8645_N$351 , \8646_N$352 ,
         \8647_N$353 , \8648_N$354 , \8649_N$355 , \8650_N$356 , \8651_N$357 , \8652_N$358 , \8653_N$359 , \8654_N$360 , \8655_N$361 , \8656_N$362 ,
         \8657_N$363 , \8658_N$364 , \8659_N$365 , \8660_N$366 , \8661_N$367 , \8662_N$368 , \8663_N$369 , \8664_N$370 , \8665_N$371 , \8666_N$372 ,
         \8667_N$373 , \8668_N$374 , \8669_N$375 , \8670_N$376 , \8671_N$377 , \8672_N$378 , \8673_N$379 , \8674_N$380 , \8675_N$381 , \8676_N$382 ,
         \8677_N$383 , \8678_N$384 , \8679_N$385 , \8680_N$386 , \8681_N$387 , \8682_N$388 , \8683_N$389 , \8684_N$390 , \8685_N$391 , \8686_N$392 ,
         \8687_N$393 , \8688_N$394 , \8689_N$395 , \8690_N$396 , \8691_N$397 , \8692_N$398 , \8693_N$399 , \8694_N$400 , \8695_N$401 , \8696_N$402 ,
         \8697_N$403 , \8698_N$404 , \8699_N$405 , \8700_N$406 , \8701_N$407 , \8702_N$408 , \8703_N$409 , \8704_N$410 , \8705_N$411 , \8706_N$412 ,
         \8707_N$413 , \8708_N$414 , \8709_N$415 , \8710_N$416 , \8711_N$417 , \8712_N$418 , \8713_N$419 , \8714_N$420 , \8715_N$421 , \8716_N$422 ,
         \8717_N$423 , \8718_N$424 , \8719_N$425 , \8720_N$426 , \8721_N$427 , \8722_N$428 , \8723_N$429 , \8724_N$430 , \8725_N$431 , \8726_N$432 ,
         \8727_N$433 , \8728_N$434 , \8729_N$435 , \8730_N$436 , \8731_N$437 , \8732_N$438 , \8733_N$439 , \8734_N$440 , \8735_N$441 , \8736_N$443 ,
         \8737_ZERO , \8738_N$2 , \8739_N$3 , \8740_N$7 , \8741_N$12 , \8742_N$13 , \8743_N$14 , \8744_N$19 , \8745_N$20 , \8746_N$27 ,
         \8747_N$28 , \8748_N$217 , \8749_N$218 , \8750_N$225 , \8751_N$442 , \8752_ONE , \8753_9052 , \8754_9053 , \8755_9054 , \8756_9055 ,
         \8757_9056 , \8758_9057 , \8759_9058 , \8760_9059 , \8761_9060 , \8762_9061 , \8763_9062 , \8764_9063 , \8765_9064 , \8766_9065 ,
         \8767_9066 , \8768_9067 , \8769_9068 , \8770_9069 , \8771_9070 , \8772_9071 , \8773_9072 , \8774_9073 , \8775_9074 , \8776_9075 ,
         \8777_9076 , \8778_9077 , \8779_9078 , \8780_9079 , \8781_9080 , \8782_9081 , \8783_9082 , \8784_9083 , \8785_9084 , \8786_9085 ,
         \8787_9086 , \8788_9087 , \8789_9088 , \8790_9089 , \8791_9090 , \8792_9091 , \8793_9092 , \8794_9093 , \8795_9094 , \8796_9095 ,
         \8797_9096 , \8798_9097 , \8799_9098 , \8800_9099 , \8801_9100 , \8802_9101 , \8803_9102 , \8804_9103 , \8805_9104 , \8806_9105 ,
         \8807_9106 , \8808_9107 , \8809_9108 , \8810_9109 , \8811_9110 , \8812_9111 , \8813_9112 , \8814_9113 , \8815_9114 , \8816_9115 ,
         \8817_9116 , \8818_9117 , \8819_9118 , \8820_9119 , \8821_9120 , \8822_9121 , \8823_9122 , \8824_9123 , \8825_9124 , \8826_9125 ,
         \8827_9126 , \8828_9127 , \8829_9128 , \8830_9129 , \8831_9130 , \8832_9131 , \8833_9132 , \8834_9133 , \8835_9134 , \8836_9135 ,
         \8837_9136 , \8838_9137 , \8839_9138 , \8840_9139 , \8841_9140 , \8842_9141 , \8843_9142 , \8844_9143 , \8845_9144 , \8846_9145 ,
         \8847_9146 , \8848_9147 , \8849_9148 , \8850_9149 , \8851_9150 , \8852_9151 , \8853_9152 , \8854_9153 , \8855_9154 , \8856_9155 ,
         \8857_9156 , \8858_9157 , \8859_9158 , \8860_9159 , \8861_9160 , \8862_9161 , \8863_9162 , \8864_9163 , \8865_9164 , \8866_9165 ,
         \8867_9166 , \8868_9167 , \8869_9168 , \8870_9169 , \8871_9170 , \8872_9171 , \8873_9172 , \8874_9173 , \8875_9174 , \8876_9175 ,
         \8877_9176 , \8878_9177 , \8879_9178 , \8880_9179 , \8881_9180 , \8882_9181 , \8883_9182 , \8884_9183 , \8885_9184 , \8886_9185 ,
         \8887_9186 , \8888_9187 , \8889_9188 , \8890_9189 , \8891_9190 , \8892_9191 , \8893_9192 , \8894_9193 , \8895_9194 , \8896_9195 ,
         \8897_9196 , \8898_9197 , \8899_9198 , \8900_9199 , \8901_9200 , \8902_9201 , \8903_9202 , \8904_9203 , \8905_9204 , \8906_9205 ,
         \8907_9206 , \8908_9207 , \8909_9208 , \8910_9209 , \8911_9210 , \8912_9211 , \8913_9212 , \8914_9213 , \8915_9214 , \8916_9215 ,
         \8917_9216 , \8918_9217 , \8919_9218 , \8920_9219 , \8921_9220 , \8922_9221 , \8923_9222 , \8924_9223 , \8925_9224 , \8926_9225 ,
         \8927_9226 , \8928_9227 , \8929_9228 , \8930_9229 , \8931_9230 , \8932_9231 , \8933_9232 , \8934_9233 , \8935_9234 , \8936_9235 ,
         \8937_9236 , \8938_9237 , \8939_9238 , \8940_9239 , \8941_9240 , \8942_9241 , \8943_9242 , \8944_9243 , \8945_9244 , \8946_9245 ,
         \8947_9246 , \8948_9247 , \8949_9248 , \8950_9249 , \8951_9250 , \8952_9251 , \8953_9252 , \8954_9253 , \8955_9254 , \8956_9255 ,
         \8957_9256 , \8958_9257 , \8959_9258 , \8960_9259 , \8961_9260 , \8962_9261 , \8963_9262 , \8964_9263 , \8965_9264 , \8966_9265 ,
         \8967_9266 , \8968_9267 , \8969_9268 , \8970_9269 , \8971_9270 , \8972_9271 , \8973_9272 , \8974_9273 , \8975_9274 , \8976_9275 ,
         \8977_9276 , \8978_9277 , \8979_9278 , \8980_9279 , \8981_9280 , \8982_9281 , \8983_9282 , \8984_9283 , \8985_9284 , \8986_9285 ,
         \8987_9286 , \8988_9287 , \8989_9288 , \8990_9289 , \8991_9290 , \8992_9291 , \8993_9292 , \8994_9293 , \8995_9294 , \8996_9295 ,
         \8997_9296 , \8998_9297 , \8999_9298 , \9000_9299 , \9001_9300 , \9002_9301 , \9003_9302 , \9004_9303 , \9005_9304 , \9006_9305 ,
         \9007_9306 , \9008_9307 , \9009_9308 , \9010_9309 , \9011_9310 , \9012_9311 , \9013_9312 , \9014_9313 , \9015_9314 , \9016_9315 ,
         \9017_9316 , \9018_9317 , \9019_9318 , \9020_9319 , \9021_9320 , \9022_9321 , \9023_9322 , \9024_9323 , \9025 , \9026_9325 ,
         \9027_9326 , \9028_9327 , \9029_9328 , \9030_9329 , \9031_9330 , \9032_9331 , \9033_9332 , \9034_9333 , \9035_9334 , \9036_9335 ,
         \9037_9336 , \9038_9337 , \9039_9338 , \9040_9339 , \9041_9340 , \9042_9341 , \9043_9342 , \9044_9343 , \9045_9344 , \9046_9345 ,
         \9047_9346 , \9048_9347 , \9049_9348 , \9050_9349 , \9051_9350 , \9052_9351 , \9053_9352 , \9054_9353 , \9055_9354 , \9056_9355 ,
         \9057_9356 , \9058_9357 , \9059_9358 , \9060_9359 , \9061_9360 , \9062_9361 , \9063_9362 , \9064_9363 , \9065_9364 , \9066_9365 ,
         \9067_9366 , \9068_9367 , \9069_9368 , \9070_9369 , \9071_9370 , \9072_9371 , \9073_9372 , \9074_9373 , \9075_9374 , \9076_9375 ,
         \9077_9376 , \9078_9377 , \9079_9378 , \9080_9379 , \9081_9380 , \9082_9381 , \9083_9382 , \9084_9383 , \9085_9384 , \9086_9385 ,
         \9087_9386 , \9088_9387 , \9089_9388 , \9090_9389 , \9091_9390 , \9092_9391 , \9093_9392 , \9094_9393 , \9095_9394 , \9096_9395 ,
         \9097_9396 , \9098_9397 , \9099_9398 , \9100_9399 , \9101_9400 , \9102_9401 , \9103_9402 , \9104_9403 , \9105_9404 , \9106_9405 ,
         \9107_9406 , \9108_9407 , \9109_9408 , \9110_9409 , \9111_9410 , \9112_9411 , \9113_9412 , \9114_9413 , \9115_9414 , \9116_9415 ,
         \9117_9416 , \9118_9417 , \9119_9418 , \9120_9419 , \9121_9420 , \9122_9421 , \9123_9422 , \9124_9423 , \9125_9424 , \9126_9425 ,
         \9127_9426 , \9128_9427 , \9129_9428 , \9130_9429 , \9131_9430 , \9132_9431 , \9133_9432 , \9134_9433 , \9135_9434 , \9136_9435 ,
         \9137_9436 , \9138_9437 , \9139_9438 , \9140_9439 , \9141_9440 , \9142_9441 , \9143_9442 , \9144_9443 , \9145_9444 , \9146_9445 ,
         \9147_9446 , \9148_9447 , \9149_9448 , \9150_9449 , \9151_9450 , \9152_9451 , \9153_9452 , \9154_9453 , \9155_9454 , \9156_9455 ,
         \9157_9456 , \9158_9457 , \9159_9458 , \9160_9459 , \9161_9460 , \9162_9461 , \9163_9462 , \9164_9463 , \9165_9464 , \9166_9465 ,
         \9167_9466 , \9168_9467 , \9169_9468 , \9170_9469 , \9171_9470 , \9172_9471 , \9173_9472 , \9174_9473 , \9175_9474 , \9176_9475 ,
         \9177_9476 , \9178_9477 , \9179_9478 , \9180_9479 , \9181_9480 , \9182_9481 , \9183_9482 , \9184_9483 , \9185_9484 , \9186_9485 ,
         \9187_9486 , \9188_9487 , \9189_9488 , \9190_9489 , \9191_9490 , \9192_9491 , \9193_9492 , \9194_9493 , \9195_9494 , \9196_9495 ,
         \9197_9496 , \9198_9497 , \9199_9498 , \9200_9499 , \9201_9500 , \9202_9501 , \9203_9502 , \9204_9503 , \9205_9504 , \9206_9505 ,
         \9207_9506 , \9208_9507 , \9209_9508 , \9210_9509 , \9211_9510 , \9212_9511 , \9213_9512 , \9214_9513 , \9215_9514 , \9216_9515 ,
         \9217_9516 , \9218_9517 , \9219_9518 , \9220_9519 , \9221_9520 , \9222_9521 , \9223_9522 , \9224_9523 , \9225_9524 , \9226_9525 ,
         \9227_9526 , \9228_9527 , \9229_9528 , \9230_9529 , \9231_9530 , \9232_9531 , \9233_9532 , \9234_9533 , \9235_9534 , \9236_9535 ,
         \9237_9536 , \9238_9537 , \9239_9538 , \9240_9539 , \9241_9540 , \9242_9541 , \9243_9542 , \9244_9543 , \9245_9544 , \9246_9545 ,
         \9247_9546 , \9248_9547 , \9249_9548 , \9250_9549 , \9251_9550 , \9252_9551 , \9253_9552 , \9254_9553 , \9255_9554 , \9256_9555 ,
         \9257_9556 , \9258_9557 , \9259_9558 , \9260_9559 , \9261_9560 , \9262_9561 , \9263_9562 , \9264_9563 , \9265_9564 , \9266_9565 ,
         \9267_9566 , \9268_9567 , \9269_9568 , \9270_9569 , \9271_9570 , \9272_9571 , \9273_9572 , \9274_9573 , \9275_9574 , \9276_9575 ,
         \9277_9576 , \9278_9577 , \9279_9578 , \9280_9579 , \9281_9580 , \9282_9581 , \9283_9582 , \9284_9583 , \9285_9584 , \9286_9585 ,
         \9287_9586 , \9288_9587 , \9289_9588 , \9290_9589 , \9291_9590 , \9292_9591 , \9293_9592 , \9294_9593 , \9295_9594 , \9296_9595 ,
         \9297_9596 , \9298_9597 , \9299 , \9300_9599 , \9301_9600 , \9302_9601 , \9303_9602 , \9304_9603 , \9305_9604 , \9306_9605 ,
         \9307_9606 , \9308_9607 , \9309_9608 , \9310_9609 , \9311_9610 , \9312_9611 , \9313_9612 , \9314_9613 , \9315_9614 , \9316_9615 ,
         \9317_9616 , \9318_9617 , \9319_9618 , \9320_9619 , \9321_9620 , \9322_9621 , \9323_9622 , \9324_9623 , \9325_9624 , \9326_9625 ,
         \9327_9626 , \9328_9627 , \9329_9628 , \9330_9629 , \9331_9630 , \9332_9631 , \9333_9632 , \9334_9633 , \9335_9634 , \9336_9635 ,
         \9337_9636 , \9338_9637 , \9339_9638 , \9340_9639 , \9341_9640 , \9342_9641 , \9343_9642 , \9344_9643 , \9345_9644 , \9346_9645 ,
         \9347_9646 , \9348_9647 , \9349_9648 , \9350_9649 , \9351_9650 , \9352_9651 , \9353_9652 , \9354_9653 , \9355_9654 , \9356_9655 ,
         \9357_9656 , \9358_9657 , \9359_9658 , \9360_9659 , \9361_9660 , \9362_9661 , \9363_9662 , \9364_9663 , \9365_9664 , \9366_9665 ,
         \9367_9666 , \9368_9667 , \9369_9668 , \9370_9669 , \9371_9670 , \9372_9671 , \9373_9672 , \9374_9673 , \9375_9674 , \9376_9675 ,
         \9377_9676 , \9378_9677 , \9379_9678 , \9380_9679 , \9381_9680 , \9382_9681 , \9383_9682 , \9384_9683 , \9385_9684 , \9386_9685 ,
         \9387_9686 , \9388_9687 , \9389_9688 , \9390_9689 , \9391_9690 , \9392_9691 , \9393_9692 , \9394_9693 , \9395_9694 , \9396_9695 ,
         \9397_9696 , \9398_9697 , \9399_9698 , \9400_9699 , \9401_9700 , \9402_9701 , \9403_9702 , \9404_9703 , \9405_9704 , \9406_9705 ,
         \9407_9706 , \9408_9707 , \9409_9708 , \9410_9709 , \9411_9710 , \9412_9711 , \9413_9712 , \9414_9713 , \9415_9714 , \9416_9715 ,
         \9417_9716 , \9418_9717 , \9419_9718 , \9420_9719 , \9421_9720 , \9422_9721 , \9423_9722 , \9424_9723 , \9425_9724 , \9426_9725 ,
         \9427_9726 , \9428_9727 , \9429_9728 , \9430_9729 , \9431_9730 , \9432_9731 , \9433 , \9434_9733 , \9435_9734 , \9436_9735 ,
         \9437_9736 , \9438_9737 , \9439_9738 , \9440_9739 , \9441_9740 , \9442_9741 , \9443_9742 , \9444_9743 , \9445_9744 , \9446_9745 ,
         \9447_9746 , \9448_9747 , \9449_9748 , \9450_9749 , \9451_9750 , \9452_9751 , \9453_9752 , \9454_9753 , \9455_9754 , \9456_9755 ,
         \9457_9756 , \9458_9757 , \9459_9758 , \9460_9759 , \9461_9760 , \9462_9761 , \9463_9762 , \9464_9763 , \9465_9764 , \9466_9765 ,
         \9467_9766 , \9468_9767 , \9469_9768 , \9470_9769 , \9471_9770 , \9472_9771 , \9473_9772 , \9474_9773 , \9475_9774 , \9476_9775 ,
         \9477_9776 , \9478_9777 , \9479_9778 , \9480_9779 , \9481_9780 , \9482_9781 , \9483_9782 , \9484_9783 , \9485_9784 , \9486_9785 ,
         \9487_9786 , \9488_9787 , \9489_9788 , \9490_9789 , \9491_9790 , \9492_9791 , \9493_9792 , \9494_9793 , \9495_9794 , \9496_9795 ,
         \9497_9796 , \9498_9797 , \9499_9798 , \9500_9799 , \9501_9800 , \9502_9801 , \9503_9802 , \9504_9803 , \9505_9804 , \9506_9805 ,
         \9507_9806 , \9508_9807 , \9509_9808 , \9510_9809 , \9511_9810 , \9512_9811 , \9513_9812 , \9514_9813 , \9515_9814 , \9516_9815 ,
         \9517_9816 , \9518_9817 , \9519_9818 , \9520_9819 , \9521_9820 , \9522_9821 , \9523_9822 , \9524_9823 , \9525_9824 , \9526_9825 ,
         \9527_9826 , \9528_9827 , \9529_9828 , \9530_9829 , \9531_9830 , \9532_9831 , \9533_9832 , \9534_9833 , \9535_9834 , \9536_9835 ,
         \9537_9836 , \9538_9837 , \9539_9838 , \9540_9839 , \9541_9840 , \9542_9841 , \9543_9842 , \9544_9843 , \9545_9844 , \9546_9845 ,
         \9547_9846 , \9548_9847 , \9549_9848 , \9550_9849 , \9551_9850 , \9552_9851 , \9553_9852 , \9554_9853 , \9555_9854 , \9556_9855 ,
         \9557_9856 , \9558_9857 , \9559_9858 , \9560_9859 , \9561_9860 , \9562_9861 , \9563_9862 , \9564_9863 , \9565_9864 , \9566 ,
         \9567_9866 , \9568_9867 , \9569_9868 , \9570_9869 , \9571_9870 , \9572_9871 , \9573_9872 , \9574_9873 , \9575_9874 , \9576_9875 ,
         \9577_9876 , \9578_9877 , \9579_9878 , \9580_9879 , \9581_9880 , \9582_9881 , \9583_9882 , \9584_9883 , \9585_9884 , \9586_9885 ,
         \9587_9886 , \9588_9887 , \9589_9888 , \9590_9889 , \9591_9890 , \9592_9891 , \9593_9892 , \9594_9893 , \9595_9894 , \9596_9895 ,
         \9597_9896 , \9598_9897 , \9599_9898 , \9600_9899 , \9601_9900 , \9602_9901 , \9603_9902 , \9604_9903 , \9605_9904 , \9606_9905 ,
         \9607_9906 , \9608_9907 , \9609_9908 , \9610_9909 , \9611_9910 , \9612_9911 , \9613_9912 , \9614_9913 , \9615_9914 , \9616_9915 ,
         \9617_9916 , \9618_9917 , \9619_9918 , \9620_9919 , \9621_9920 , \9622_9921 , \9623_9922 , \9624_9923 , \9625_9924 , \9626_9925 ,
         \9627_9926 , \9628_9927 , \9629_9928 , \9630_9929 , \9631_9930 , \9632_9931 , \9633_9932 , \9634_9933 , \9635_9934 , \9636_9935 ,
         \9637_9936 , \9638_9937 , \9639_9938 , \9640_9939 , \9641_9940 , \9642_9941 , \9643_9942 , \9644_9943 , \9645_9944 , \9646_9945 ,
         \9647_9946 , \9648_9947 , \9649_9948 , \9650_9949 , \9651_9950 , \9652_9951 , \9653_9952 , \9654_9953 , \9655_9954 , \9656_9955 ,
         \9657_9956 , \9658_9957 , \9659_9958 , \9660_9959 , \9661_9960 , \9662_9961 , \9663_9962 , \9664_9963 , \9665_9964 , \9666_9965 ,
         \9667_9966 , \9668_9967 , \9669_9968 , \9670_9969 , \9671_9970 , \9672_9971 , \9673_9972 , \9674_9973 , \9675_9974 , \9676_9975 ,
         \9677_9976 , \9678_9977 , \9679_9978 , \9680_9979 , \9681_9980 , \9682_9981 , \9683_9982 , \9684_9983 , \9685_9984 , \9686_9985 ,
         \9687_9986 , \9688_9987 , \9689_9988 , \9690_9989 , \9691_9990 , \9692_9991 , \9693_9992 , \9694_9993 , \9695_9994 , \9696_9995 ,
         \9697_9996 , \9698_9997 , \9699_9998 , \9700 , \9701_10000 , \9702_10001 , \9703_10002 , \9704_10003 , \9705_10004 , \9706_10005 ,
         \9707_10006 , \9708_10007 , \9709_10008 , \9710_10009 , \9711_10010 , \9712_10011 , \9713_10012 , \9714_10013 , \9715_10014 , \9716_10015 ,
         \9717_10016 , \9718_10017 , \9719_10018 , \9720_10019 , \9721_10020 , \9722_10021 , \9723_10022 , \9724_10023 , \9725_10024 , \9726_10025 ,
         \9727_10026 , \9728_10027 , \9729_10028 , \9730_10029 , \9731_10030 , \9732_10031 , \9733_10032 , \9734_10033 , \9735_10034 , \9736_10035 ,
         \9737_10036 , \9738_10037 , \9739_10038 , \9740_10039 , \9741_10040 , \9742_10041 , \9743_10042 , \9744_10043 , \9745_10044 , \9746_10045 ,
         \9747_10046 , \9748_10047 , \9749_10048 , \9750_10049 , \9751_10050 , \9752_10051 , \9753_10052 , \9754_10053 , \9755_10054 , \9756_10055 ,
         \9757_10056 , \9758_10057 , \9759_10058 , \9760_10059 , \9761_10060 , \9762_10061 , \9763_10062 , \9764_10063 , \9765_10064 , \9766_10065 ,
         \9767_10066 , \9768_10067 , \9769_10068 , \9770_10069 , \9771_10070 , \9772_10071 , \9773_10072 , \9774_10073 , \9775_10074 , \9776_10075 ,
         \9777_10076 , \9778_10077 , \9779_10078 , \9780_10079 , \9781_10080 , \9782_10081 , \9783_10082 , \9784_10083 , \9785_10084 , \9786_10085 ,
         \9787_10086 , \9788_10087 , \9789_10088 , \9790_10089 , \9791_10090 , \9792_10091 , \9793_10092 , \9794_10093 , \9795_10094 , \9796_10095 ,
         \9797_10096 , \9798_10097 , \9799_10098 , \9800_10099 , \9801_10100 , \9802_10101 , \9803_10102 , \9804_10103 , \9805_10104 , \9806_10105 ,
         \9807_10106 , \9808_10107 , \9809_10108 , \9810_10109 , \9811_10110 , \9812_10111 , \9813_10112 , \9814_10113 , \9815_10114 , \9816_10115 ,
         \9817_10116 , \9818_10117 , \9819_10118 , \9820_10119 , \9821_10120 , \9822_10121 , \9823_10122 , \9824_10123 , \9825_10124 , \9826_10125 ,
         \9827_10126 , \9828_10127 , \9829_10128 , \9830_10129 , \9831_10130 , \9832_10131 , \9833 , \9834_10133 , \9835_10134 , \9836_10135 ,
         \9837_10136 , \9838_10137 , \9839_10138 , \9840_10139 , \9841_10140 , \9842_10141 , \9843_10142 , \9844_10143 , \9845_10144 , \9846_10145 ,
         \9847_10146 , \9848_10147 , \9849_10148 , \9850_10149 , \9851_10150 , \9852_10151 , \9853_10152 , \9854_10153 , \9855_10154 , \9856_10155 ,
         \9857_10156 , \9858_10157 , \9859_10158 , \9860_10159 , \9861_10160 , \9862_10161 , \9863_10162 , \9864_10163 , \9865_10164 , \9866_10165 ,
         \9867_10166 , \9868_10167 , \9869_10168 , \9870_10169 , \9871_10170 , \9872_10171 , \9873_10172 , \9874_10173 , \9875_10174 , \9876_10175 ,
         \9877_10176 , \9878_10177 , \9879_10178 , \9880_10179 , \9881_10180 , \9882_10181 , \9883_10182 , \9884_10183 , \9885_10184 , \9886_10185 ,
         \9887_10186 , \9888_10187 , \9889_10188 , \9890_10189 , \9891_10190 , \9892_10191 , \9893_10192 , \9894_10193 , \9895_10194 , \9896_10195 ,
         \9897_10196 , \9898_10197 , \9899_10198 , \9900_10199 , \9901_10200 , \9902_10201 , \9903_10202 , \9904_10203 , \9905_10204 , \9906_10205 ,
         \9907_10206 , \9908_10207 , \9909_10208 , \9910_10209 , \9911_10210 , \9912_10211 , \9913_10212 , \9914_10213 , \9915_10214 , \9916_10215 ,
         \9917_10216 , \9918_10217 , \9919_10218 , \9920_10219 , \9921_10220 , \9922_10221 , \9923_10222 , \9924_10223 , \9925_10224 , \9926_10225 ,
         \9927_10226 , \9928_10227 , \9929_10228 , \9930_10229 , \9931_10230 , \9932_10231 , \9933_10232 , \9934_10233 , \9935_10234 , \9936_10235 ,
         \9937_10236 , \9938_10237 , \9939_10238 , \9940_10239 , \9941_10240 , \9942_10241 , \9943_10242 , \9944_10243 , \9945_10244 , \9946_10245 ,
         \9947_10246 , \9948_10247 , \9949_10248 , \9950_10249 , \9951_10250 , \9952_10251 , \9953_10252 , \9954_10253 , \9955_10254 , \9956_10255 ,
         \9957_10256 , \9958_10257 , \9959_10258 , \9960_10259 , \9961_10260 , \9962_10261 , \9963_10262 , \9964_10263 , \9965_10264 , \9966_10265 ,
         \9967 , \9968_10267 , \9969_10268 , \9970_10269 , \9971_10270 , \9972_10271 , \9973_10272 , \9974_10273 , \9975_10274 , \9976_10275 ,
         \9977_10276 , \9978_10277 , \9979_10278 , \9980_10279 , \9981_10280 , \9982_10281 , \9983_10282 , \9984_10283 , \9985_10284 , \9986_10285 ,
         \9987_10286 , \9988_10287 , \9989_10288 , \9990_10289 , \9991_10290 , \9992_10291 , \9993_10292 , \9994_10293 , \9995_10294 , \9996_10295 ,
         \9997_10296 , \9998_10297 , \9999_10298 , \10000_10299 , \10001_10300 , \10002_10301 , \10003_10302 , \10004_10303 , \10005_10304 , \10006_10305 ,
         \10007_10306 , \10008_10307 , \10009_10308 , \10010_10309 , \10011_10310 , \10012_10311 , \10013_10312 , \10014_10313 , \10015_10314 , \10016_10315 ,
         \10017_10316 , \10018_10317 , \10019_10318 , \10020_10319 , \10021_10320 , \10022_10321 , \10023_10322 , \10024_10323 , \10025_10324 , \10026_10325 ,
         \10027_10326 , \10028_10327 , \10029_10328 , \10030_10329 , \10031_10330 , \10032_10331 , \10033_10332 , \10034_10333 , \10035_10334 , \10036_10335 ,
         \10037_10336 , \10038_10337 , \10039_10338 , \10040_10339 , \10041_10340 , \10042_10341 , \10043_10342 , \10044_10343 , \10045_10344 , \10046_10345 ,
         \10047_10346 , \10048_10347 , \10049_10348 , \10050_10349 , \10051_10350 , \10052_10351 , \10053_10352 , \10054_10353 , \10055_10354 , \10056_10355 ,
         \10057_10356 , \10058_10357 , \10059_10358 , \10060_10359 , \10061_10360 , \10062_10361 , \10063_10362 , \10064_10363 , \10065_10364 , \10066_10365 ,
         \10067_10366 , \10068_10367 , \10069_10368 , \10070_10369 , \10071_10370 , \10072_10371 , \10073_10372 , \10074_10373 , \10075_10374 , \10076_10375 ,
         \10077_10376 , \10078_10377 , \10079_10378 , \10080_10379 , \10081_10380 , \10082_10381 , \10083_10382 , \10084_10383 , \10085_10384 , \10086_10385 ,
         \10087_10386 , \10088_10387 , \10089_10388 , \10090_10389 , \10091_10390 , \10092_10391 , \10093_10392 , \10094_10393 , \10095_10394 , \10096_10395 ,
         \10097_10396 , \10098_10397 , \10099_10398 , \10100 , \10101_10400 , \10102_10401 , \10103_10402 , \10104_10403 , \10105_10404 , \10106_10405 ,
         \10107_10406 , \10108_10407 , \10109_10408 , \10110_10409_nG444e , \10111_10410 , \10112_10411 , \10113_10412_nG4451 , \10114_10413 , \10115_10414 , \10116_10415_nG4454 ,
         \10117_10416 , \10118_10417 , \10119_10418 , \10120_10422 , \10121_10423 , \10122_10424 , \10123_10425 , \10124_10426 , \10125_10427 , \10126_10428 ,
         \10127_10429 , \10128_10430 , \10129_10431 , \10130_10432 , \10131_10433 , \10132_10434 , \10133_10435 , \10134_10436 , \10135_10437 , \10136_10438 ,
         \10137_10439 , \10138_10440 , \10139_10441 , \10140_10442 , \10141_10443 , \10142_10444 , \10143_10445 , \10144_10446 , \10145_10447 , \10146_10448 ,
         \10147_10449 , \10148_10450 , \10149_10451 , \10150_10452 , \10151_10453 , \10152_10454 , \10153_10455 , \10154_10456 , \10155_10457 , \10156_10458 ,
         \10157_10459 , \10158_10460 , \10159_10461 , \10160_10462 , \10161_10463 , \10162_10464 , \10163_10465 , \10164_10466 , \10165_10467 , \10166_10468 ,
         \10167_10469 , \10168_10470 , \10169_10471 , \10170_10472 , \10171_10473 , \10172_10474 , \10173_10475 , \10174_10476 , \10175_10477 , \10176_10478 ,
         \10177_10479 , \10178_10480 , \10179_10481 , \10180_10482 , \10181_10483 , \10182_10484 , \10183_10485 , \10184_10486 , \10185_10487 , \10186_10488 ,
         \10187_10489 , \10188_10490 , \10189_10491 , \10190_10492 , \10191_10493 , \10192_10494 , \10193_10495 , \10194_10496 , \10195_10497 , \10196_10498 ,
         \10197_10499 , \10198_10500 , \10199_10501 , \10200_10502 , \10201_10503 , \10202_10504 , \10203_10505 , \10204_10506 , \10205_10507 , \10206_10508 ,
         \10207_10509 , \10208_10510 , \10209_10511 , \10210_10512 , \10211_10513 , \10212_10514 , \10213_10515 , \10214_10516 , \10215_10517 , \10216_10518 ,
         \10217_10519 , \10218_10520 , \10219_10521 , \10220_10522 , \10221_10523 , \10222_10524 , \10223_10525 , \10224_10526 , \10225_10527 , \10226_10528 ,
         \10227_10529 , \10228_10530 , \10229_10531 , \10230_10532 , \10231_10533 , \10232_10534 , \10233_10535 , \10234_10536 , \10235_10537 , \10236_10538 ,
         \10237_10539 , \10238_10540 , \10239_10541 , \10240_10542 , \10241_10543 , \10242_10544 , \10243_10545 , \10244_10546 , \10245_10547 , \10246_10548 ,
         \10247_10549 , \10248_10550 , \10249_10551 , \10250_10552 , \10251 , \10252_10554 , \10253_10555 , \10254_10556 , \10255_10557 , \10256_10558 ,
         \10257_10559 , \10258_10560 , \10259_10561 , \10260_10562 , \10261_10563 , \10262_10564 , \10263_10565 , \10264_10566 , \10265_10567 , \10266_10568 ,
         \10267_10569 , \10268_10570 , \10269_10571 , \10270_10572 , \10271_10573 , \10272_10574 , \10273_10575 , \10274_10576 , \10275_10577 , \10276_10578 ,
         \10277_10579 , \10278_10580 , \10279_10581 , \10280_10582 , \10281_10583 , \10282_10584 , \10283_10585 , \10284_10586 , \10285_10587 , \10286_10588 ,
         \10287_10589 , \10288_10590 , \10289_10591 , \10290_10592 , \10291_10593 , \10292_10594 , \10293_10595 , \10294_10596 , \10295_10597 , \10296_10598 ,
         \10297_10599 , \10298_10600 , \10299_10601 , \10300_10602 , \10301_10603 , \10302_10604 , \10303_10605 , \10304_10606 , \10305_10607 , \10306_10608 ,
         \10307_10609 , \10308_10610 , \10309_10611 , \10310_10612 , \10311_10613 , \10312_10614 , \10313_10615 , \10314_10616 , \10315_10617 , \10316_10618 ,
         \10317_10619 , \10318_10620 , \10319_10621 , \10320_10622 , \10321_10623 , \10322_10624 , \10323_10625 , \10324_10626 , \10325_10627 , \10326_10628 ,
         \10327_10629 , \10328_10630 , \10329_10631 , \10330_10632 , \10331_10633 , \10332_10634 , \10333_10635 , \10334_10636 , \10335_10637 , \10336_10638 ,
         \10337_10639 , \10338_10640 , \10339_10641 , \10340_10642 , \10341_10643 , \10342_10644 , \10343_10645 , \10344_10646 , \10345_10647 , \10346_10648 ,
         \10347_10649 , \10348_10650 , \10349_10651 , \10350_10652 , \10351_10653 , \10352_10654 , \10353_10655 , \10354_10656 , \10355_10657 , \10356_10658 ,
         \10357_10659 , \10358_10660 , \10359_10661 , \10360_10662 , \10361_10663 , \10362_10664 , \10363_10665 , \10364_10666 , \10365_10667 , \10366_10668 ,
         \10367_10669 , \10368_10670 , \10369_10671 , \10370_10672 , \10371_10673 , \10372_10674 , \10373_10675 , \10374_10676 , \10375_10677 , \10376_10678 ,
         \10377_10679 , \10378_10680 , \10379_10681 , \10380_10682 , \10381_10683 , \10382_10684 , \10383 , \10384_10686_nG6579 , \10385_10687 , \10386 ,
         \10387 , \10388_10690_nG455f , \10389_10691 , \10390_10692 , \10391_10693 , \10392_10694_nG9c0e , \10393_10695 , \10394_10696 , \10395_10697 , \10396_10698 ,
         \10397_10699 , \10398_10700 , \10399_10703 , \10400_10701 , \10401_10702_nG4456 , \10402_10704 , \10403_10708 , \10404_10709 , \10405_10710 , \10406_10711 ,
         \10407_10712 , \10408_10713 , \10409_10705 , \10410_10706 , \10411_10707 , \10412_10714 , \10413_10715 , \10414_10716 , \10415_10717 , \10416_10718 ,
         \10417_10719 , \10418_10720 , \10419_10721 , \10420_10722 , \10421_10723 , \10422_10724 , \10423_10725 , \10424_10726 , \10425_10727 , \10426_10728 ,
         \10427_10729 , \10428_10730 , \10429_10731 , \10430_10732 , \10431_10733 , \10432_10734 , \10433_10735 , \10434_10736 , \10435_10737 , \10436_10738 ,
         \10437_10739 , \10438_10740 , \10439_10741 , \10440_10742 , \10441_10743 , \10442_10744 , \10443_10745 , \10444_10746 , \10445_10747 , \10446_10748 ,
         \10447_10749 , \10448_10750 , \10449_10751 , \10450_10752 , \10451_10753 , \10452_10754 , \10453_10755 , \10454_10756 , \10455_10757 , \10456_10758 ,
         \10457_10759 , \10458_10760 , \10459_10761 , \10460_10762 , \10461_10763 , \10462_10764 , \10463_10765 , \10464_10766 , \10465_10767 , \10466_10768 ,
         \10467_10769 , \10468_10770 , \10469_10771 , \10470_10772 , \10471_10773 , \10472_10774 , \10473_10775 , \10474_10776 , \10475_10777 , \10476_10778 ,
         \10477_10779 , \10478_10780 , \10479_10781 , \10480_10782 , \10481_10783 , \10482_10784 , \10483_10785 , \10484_10786 , \10485_10787 , \10486_10788 ,
         \10487_10789 , \10488_10790 , \10489_10791 , \10490_10792 , \10491_10793 , \10492_10794 , \10493_10795 , \10494_10796 , \10495_10797 , \10496_10798 ,
         \10497_10799 , \10498_10800 , \10499_10801 , \10500_10802 , \10501_10803 , \10502_10804 , \10503_10805 , \10504_10806 , \10505_10807 , \10506_10808 ,
         \10507_10809 , \10508_10810 , \10509_10811 , \10510_10812 , \10511_10813 , \10512_10814 , \10513_10815 , \10514_10816 , \10515_10817 , \10516_10818 ,
         \10517_10819 , \10518_10820 , \10519_10821 , \10520_10822 , \10521_10823 , \10522_10824 , \10523_10825 , \10524_10826 , \10525_10827 , \10526_10828 ,
         \10527_10829 , \10528_10830 , \10529_10831 , \10530_10832 , \10531_10833 , \10532_10834 , \10533_10835 , \10534_10836 , \10535_10837 , \10536_10838 ,
         \10537_10839 , \10538_10840 , \10539_10841 , \10540_10842 , \10541_10843 , \10542_10844 , \10543_10845 , \10544 , \10545_10847 , \10546_10848 ,
         \10547_10849 , \10548_10850 , \10549_10851 , \10550_10852 , \10551_10853 , \10552_10854 , \10553_10855 , \10554_10856 , \10555_10857 , \10556_10858 ,
         \10557_10859 , \10558_10860 , \10559_10861 , \10560_10862 , \10561_10863 , \10562_10864 , \10563_10865 , \10564_10866 , \10565_10867 , \10566_10868 ,
         \10567_10869 , \10568_10870 , \10569_10871 , \10570_10872 , \10571_10873 , \10572_10874 , \10573_10875 , \10574_10876 , \10575_10877 , \10576_10878 ,
         \10577_10879 , \10578_10880 , \10579_10881 , \10580_10882 , \10581_10883 , \10582_10884 , \10583_10885 , \10584_10886 , \10585_10887 , \10586_10888 ,
         \10587_10889 , \10588_10890 , \10589_10891 , \10590_10892 , \10591_10893 , \10592_10894 , \10593_10895 , \10594_10896 , \10595_10897 , \10596_10898 ,
         \10597_10899 , \10598_10900 , \10599_10901 , \10600_10902 , \10601_10903 , \10602_10904 , \10603_10905 , \10604_10906 , \10605_10907 , \10606_10908 ,
         \10607_10909 , \10608_10910 , \10609_10911 , \10610_10912 , \10611_10913 , \10612_10914 , \10613_10915 , \10614_10916 , \10615_10917 , \10616_10918 ,
         \10617_10919 , \10618_10920 , \10619_10921 , \10620_10922 , \10621_10923 , \10622_10924 , \10623_10925 , \10624_10926 , \10625_10927 , \10626_10928 ,
         \10627_10929 , \10628_10930 , \10629_10931 , \10630_10932 , \10631_10933 , \10632_10934 , \10633_10935 , \10634_10936 , \10635_10937 , \10636_10938 ,
         \10637_10939 , \10638_10940 , \10639_10941 , \10640_10942 , \10641_10943 , \10642_10944 , \10643_10945 , \10644_10946 , \10645_10947 , \10646_10948 ,
         \10647_10949 , \10648_10950 , \10649_10951 , \10650_10952 , \10651_10953 , \10652_10954 , \10653_10955 , \10654_10956 , \10655_10957 , \10656_10958 ,
         \10657_10959 , \10658_10960 , \10659_10961 , \10660_10962 , \10661_10963 , \10662_10964 , \10663_10965 , \10664_10966 , \10665_10967 , \10666_10968 ,
         \10667_10969 , \10668_10970 , \10669_10971 , \10670_10972 , \10671_10973 , \10672_10974 , \10673_10975 , \10674_10976 , \10675_10977 , \10676 ,
         \10677_10979_nG4668 , \10678_10980 , \10679_10981 , \10680_10982 , \10681_10983 , \10682_10984 , \10683 , \10684 , \10685_10987_nG657c , \10686_10988 ,
         \10687_10989 , \10688_10990 , \10689_10991 , \10690_10992 , \10691_10993 , \10692_10994 , \10693_10995_nG9c0b , \10694_10996 , \10695_10997 , \10696_10998 ,
         \10697_10999 , \10698_11000 , \10699_11001 , \10700_11002 , \10701_11003 , \10702_11004 , \10703_11005 , \10704_11006 , \10705_11007 , \10706_11008 ,
         \10707_11009 , \10708_11010 , \10709_11011 , \10710_11012 , \10711_11013 , \10712_11014 , \10713_11015 , \10714_11016 , \10715_11017 , \10716_11018 ,
         \10717_11019 , \10718_11020 , \10719_11021 , \10720_11022 , \10721_11023 , \10722_11024 , \10723_11025 , \10724_11026 , \10725_11027 , \10726_11028 ,
         \10727_11029 , \10728_11030 , \10729_11031 , \10730_11032 , \10731_11033 , \10732_11034 , \10733_11035 , \10734_11036 , \10735_11037 , \10736_11038 ,
         \10737_11039 , \10738_11040 , \10739_11041 , \10740_11042 , \10741_11043 , \10742_11044 , \10743_11045 , \10744_11046 , \10745_11047 , \10746_11048 ,
         \10747_11049 , \10748_11050 , \10749_11051 , \10750_11052 , \10751_11053 , \10752_11054 , \10753_11055 , \10754_11056 , \10755_11057 , \10756_11058 ,
         \10757_11059 , \10758_11060 , \10759_11061 , \10760_11062 , \10761_11063 , \10762_11064 , \10763_11065 , \10764_11066 , \10765_11067 , \10766_11068 ,
         \10767_11069 , \10768_11070 , \10769_11071 , \10770_11072 , \10771_11073 , \10772_11074 , \10773_11075 , \10774_11076 , \10775_11077 , \10776_11078 ,
         \10777_11079 , \10778_11080 , \10779_11081 , \10780_11082 , \10781_11083 , \10782_11084 , \10783_11085 , \10784_11086 , \10785_11087 , \10786_11088 ,
         \10787_11089 , \10788_11090 , \10789_11091 , \10790_11092 , \10791_11093 , \10792_11094 , \10793_11095 , \10794_11096 , \10795_11097 , \10796_11098 ,
         \10797_11099 , \10798_11100 , \10799_11101 , \10800_11102 , \10801_11103 , \10802_11104 , \10803_11105 , \10804_11106 , \10805_11107 , \10806_11108 ,
         \10807_11109 , \10808_11110 , \10809_11111 , \10810_11112 , \10811_11113 , \10812_11114 , \10813_11115 , \10814_11116 , \10815_11117 , \10816_11118 ,
         \10817_11119 , \10818_11120 , \10819_11121 , \10820_11122 , \10821_11123 , \10822_11124 , \10823_11125 , \10824_11126 , \10825_11127 , \10826_11128 ,
         \10827_11129 , \10828_11130 , \10829_11131 , \10830_11132 , \10831_11133 , \10832_11134 , \10833_11135 , \10834 , \10835_11137 , \10836_11138 ,
         \10837_11139 , \10838_11140 , \10839_11141 , \10840_11142 , \10841_11143 , \10842_11144 , \10843_11145 , \10844_11146 , \10845_11147 , \10846_11148 ,
         \10847_11149 , \10848_11150 , \10849_11151 , \10850_11152 , \10851_11153 , \10852_11154 , \10853_11155 , \10854_11156 , \10855_11157 , \10856_11158 ,
         \10857_11159 , \10858_11160 , \10859_11161 , \10860_11162 , \10861_11163 , \10862_11164 , \10863_11165 , \10864_11166 , \10865_11167 , \10866_11168 ,
         \10867_11169 , \10868_11170 , \10869_11171 , \10870_11172 , \10871_11173 , \10872_11174 , \10873_11175 , \10874_11176 , \10875_11177 , \10876_11178 ,
         \10877_11179 , \10878_11180 , \10879_11181 , \10880_11182 , \10881_11183 , \10882_11184 , \10883_11185 , \10884_11186 , \10885_11187 , \10886_11188 ,
         \10887_11189 , \10888_11190 , \10889_11191 , \10890_11192 , \10891_11193 , \10892_11194 , \10893_11195 , \10894_11196 , \10895_11197 , \10896_11198 ,
         \10897_11199 , \10898_11200 , \10899_11201 , \10900_11202 , \10901_11203 , \10902_11204 , \10903_11205 , \10904_11206 , \10905_11207 , \10906_11208 ,
         \10907_11209 , \10908_11210 , \10909_11211 , \10910_11212 , \10911_11213 , \10912_11214 , \10913_11215 , \10914_11216 , \10915_11217 , \10916_11218 ,
         \10917_11219 , \10918_11220 , \10919_11221 , \10920_11222 , \10921_11223 , \10922_11224 , \10923_11225 , \10924_11226 , \10925_11227 , \10926_11228 ,
         \10927_11229 , \10928_11230 , \10929_11231 , \10930_11232 , \10931_11233 , \10932_11234 , \10933_11235 , \10934_11236 , \10935_11237 , \10936_11238 ,
         \10937_11239 , \10938_11240 , \10939_11241 , \10940_11242 , \10941_11243 , \10942_11244 , \10943_11245 , \10944_11246 , \10945_11247 , \10946_11248 ,
         \10947_11249 , \10948_11250 , \10949_11251 , \10950_11252 , \10951_11253 , \10952_11254 , \10953_11255 , \10954_11256 , \10955_11257 , \10956_11258 ,
         \10957_11259 , \10958_11260 , \10959_11261 , \10960_11262 , \10961_11263 , \10962_11264 , \10963_11265 , \10964_11266 , \10965_11267 , \10966 ,
         \10967_11269_nG657f , \10968_11270 , \10969_11271 , \10970_11272 , \10971_11273 , \10972 , \10973 , \10974_11276_nG4771 , \10975_11277 , \10976_11278 ,
         \10977_11279 , \10978_11280 , \10979_11281 , \10980_11282 , \10981_11283_nG9c08 , \10982_11284 , \10983_11285 , \10984_11286 , \10985_11287 , \10986_11288 ,
         \10987_11289 , \10988_11290 , \10989_11291 , \10990_11292 , \10991_11293 , \10992_11294 , \10993_11295 , \10994_10419 , \10995_10420 , \10996_10421 ,
         \10997_11296 , \10998_11297 , \10999_11298 , \11000_11299 , \11001_11300 , \11002_11301 , \11003_11302 , \11004_11303 , \11005_11304 , \11006_11305 ,
         \11007_11306 , \11008_11307 , \11009_11308 , \11010_11309 , \11011_11310 , \11012_11311 , \11013_11312 , \11014_11313 , \11015_11314 , \11016_11315 ,
         \11017_11316 , \11018_11317 , \11019_11318 , \11020_11319 , \11021_11320 , \11022_11321 , \11023_11322 , \11024_11323 , \11025_11324 , \11026_11325 ,
         \11027_11326 , \11028_11327 , \11029_11328 , \11030_11329 , \11031_11330 , \11032_11331 , \11033_11332 , \11034_11333 , \11035_11334 , \11036_11335 ,
         \11037_11336 , \11038_11337 , \11039_11338 , \11040_11339 , \11041_11340 , \11042_11341 , \11043_11342 , \11044_11343 , \11045_11344 , \11046_11345 ,
         \11047_11346 , \11048_11347 , \11049_11348 , \11050_11349 , \11051_11350 , \11052_11351 , \11053_11352 , \11054_11353 , \11055_11354 , \11056_11355 ,
         \11057_11356 , \11058_11357 , \11059_11358 , \11060_11359 , \11061_11360 , \11062_11361 , \11063_11362 , \11064_11363 , \11065_11364 , \11066_11365 ,
         \11067_11366 , \11068_11367 , \11069_11368 , \11070_11369 , \11071_11370 , \11072_11371 , \11073_11372 , \11074_11373 , \11075_11374 , \11076_11375 ,
         \11077_11376 , \11078_11377 , \11079_11378 , \11080_11379 , \11081_11380 , \11082_11381 , \11083_11382 , \11084_11383 , \11085_11384 , \11086_11385 ,
         \11087_11386 , \11088_11387 , \11089_11388 , \11090_11389 , \11091_11390 , \11092_11391 , \11093_11392 , \11094_11393 , \11095_11394 , \11096_11395 ,
         \11097_11396 , \11098_11397 , \11099_11398 , \11100_11399 , \11101_11400 , \11102_11401 , \11103_11402 , \11104_11403 , \11105_11404 , \11106_11405 ,
         \11107_11406 , \11108_11407 , \11109_11408 , \11110_11409 , \11111_11410 , \11112_11411 , \11113_11412 , \11114_11413 , \11115_11414 , \11116_11415 ,
         \11117_11416 , \11118_11417 , \11119_11418 , \11120_11419 , \11121_11420 , \11122_11421 , \11123_11422 , \11124_11423 , \11125_11424 , \11126_11425 ,
         \11127_11426 , \11128_11427 , \11129_11428 , \11130_11429 , \11131_11430 , \11132_11431 , \11133_11432 , \11134_11433 , \11135_11434 , \11136_11435 ,
         \11137_11436 , \11138 , \11139_11438 , \11140_11439 , \11141_11440 , \11142_11441 , \11143_11442 , \11144_11443 , \11145_11444 , \11146_11445 ,
         \11147_11446 , \11148_11447 , \11149_11448 , \11150_11449 , \11151_11450 , \11152_11451 , \11153_11452 , \11154_11453 , \11155_11454 , \11156_11455 ,
         \11157_11456 , \11158_11457 , \11159_11458 , \11160_11459 , \11161_11460 , \11162_11461 , \11163_11462 , \11164_11463 , \11165_11464 , \11166_11465 ,
         \11167_11466 , \11168_11467 , \11169_11468 , \11170_11469 , \11171_11470 , \11172_11471 , \11173_11472 , \11174_11473 , \11175_11474 , \11176_11475 ,
         \11177_11476 , \11178_11477 , \11179_11478 , \11180_11479 , \11181_11480 , \11182_11481 , \11183_11482 , \11184_11483 , \11185_11484 , \11186_11485 ,
         \11187_11486 , \11188_11487 , \11189_11488 , \11190_11489 , \11191_11490 , \11192_11491 , \11193_11492 , \11194_11493 , \11195_11494 , \11196_11495 ,
         \11197_11496 , \11198_11497 , \11199_11498 , \11200_11499 , \11201_11500 , \11202_11501 , \11203_11502 , \11204_11503 , \11205_11504 , \11206_11505 ,
         \11207_11506 , \11208_11507 , \11209_11508 , \11210_11509 , \11211_11510 , \11212_11511 , \11213_11512 , \11214_11513 , \11215_11514 , \11216_11515 ,
         \11217_11516 , \11218_11517 , \11219_11518 , \11220_11519 , \11221_11520 , \11222_11521 , \11223_11522 , \11224_11523 , \11225_11524 , \11226_11525 ,
         \11227_11526 , \11228_11527 , \11229_11528 , \11230_11529 , \11231_11530 , \11232_11531 , \11233_11532 , \11234_11533 , \11235_11534 , \11236_11535 ,
         \11237_11536 , \11238_11537 , \11239_11538 , \11240_11539 , \11241_11540 , \11242_11541 , \11243_11542 , \11244_11543 , \11245_11544 , \11246_11545 ,
         \11247_11546 , \11248_11547 , \11249_11548 , \11250_11549 , \11251_11550 , \11252_11551 , \11253_11552 , \11254_11553 , \11255_11554 , \11256_11555 ,
         \11257_11556 , \11258_11557 , \11259_11558 , \11260_11559 , \11261_11560 , \11262_11561 , \11263_11562 , \11264_11563 , \11265_11564 , \11266_11565 ,
         \11267_11566 , \11268_11567 , \11269_11568 , \11270 , \11271_11570_nG487a , \11272_11571 , \11273_11572 , \11274_11573 , \11275_11574 , \11276_11575 ,
         \11277_11576 , \11278_11577 , \11279_11578 , \11280_11579 , \11281_11580 , \11282_11581 , \11283_11582 , \11284 , \11285 , \11286_11585_nG6582 ,
         \11287_11586 , \11288_11587 , \11289_11588 , \11290_11589 , \11291_11590 , \11292_11591 , \11293_11592 , \11294_11593 , \11295_11594 , \11296_11595 ,
         \11297_11596 , \11298_11597 , \11299_11598_nG9c05 , \11300_11599 , \11301_11600 , \11302_11601 , \11303_11602 , \11304_11603 , \11305_11604 , \11306_11605 ,
         \11307_11606 , \11308_11607 , \11309_11608 , \11310_11609 , \11311_11610 , \11312_11611 , \11313_11612 , \11314_11613 , \11315_11614 , \11316_11615 ,
         \11317_11616 , \11318_11617 , \11319_11618 , \11320_11619 , \11321_11620 , \11322_11621 , \11323_11622 , \11324_11623 , \11325_11624 , \11326_11625 ,
         \11327_11626 , \11328_11627 , \11329_11628 , \11330_11629 , \11331_11630 , \11332_11631 , \11333_11632 , \11334_11633 , \11335_11634 , \11336_11635 ,
         \11337_11636 , \11338_11637 , \11339_11638 , \11340_11639 , \11341_11640 , \11342_11641 , \11343_11642 , \11344_11643 , \11345_11644 , \11346_11645 ,
         \11347_11646 , \11348_11647 , \11349_11648 , \11350_11649 , \11351_11650 , \11352_11651 , \11353_11652 , \11354_11653 , \11355_11654 , \11356_11655 ,
         \11357_11656 , \11358_11657 , \11359_11658 , \11360_11659 , \11361_11660 , \11362_11661 , \11363_11662 , \11364_11663 , \11365_11664 , \11366_11665 ,
         \11367_11666 , \11368_11667 , \11369_11668 , \11370_11669 , \11371_11670 , \11372_11671 , \11373_11672 , \11374_11673 , \11375_11674 , \11376_11675 ,
         \11377_11676 , \11378_11677 , \11379_11678 , \11380_11679 , \11381_11680 , \11382_11681 , \11383_11682 , \11384_11683 , \11385_11684 , \11386_11685 ,
         \11387_11686 , \11388_11687 , \11389_11688 , \11390_11689 , \11391_11690 , \11392_11691 , \11393_11692 , \11394_11693 , \11395_11694 , \11396_11695 ,
         \11397_11696 , \11398_11697 , \11399_11698 , \11400_11699 , \11401_11700 , \11402_11701 , \11403_11702 , \11404_11703 , \11405_11704 , \11406_11705 ,
         \11407_11706 , \11408_11707 , \11409_11708 , \11410_11709 , \11411_11710 , \11412_11711 , \11413_11712 , \11414_11713 , \11415_11714 , \11416_11715 ,
         \11417_11716 , \11418_11717 , \11419_11718 , \11420_11719 , \11421_11720 , \11422_11721 , \11423_11722 , \11424_11723 , \11425_11724 , \11426_11725 ,
         \11427_11726 , \11428_11727 , \11429_11728 , \11430_11729 , \11431_11730 , \11432_11731 , \11433_11732 , \11434_11733 , \11435_11734 , \11436_11735 ,
         \11437_11736 , \11438 , \11439_11738 , \11440_11739 , \11441_11740 , \11442_11741 , \11443_11742 , \11444_11743 , \11445_11744 , \11446_11745 ,
         \11447_11746 , \11448_11747 , \11449_11748 , \11450_11749 , \11451_11750 , \11452_11751 , \11453_11752 , \11454_11753 , \11455_11754 , \11456_11755 ,
         \11457_11756 , \11458_11757 , \11459_11758 , \11460_11759 , \11461_11760 , \11462_11761 , \11463_11762 , \11464_11763 , \11465_11764 , \11466_11765 ,
         \11467_11766 , \11468_11767 , \11469_11768 , \11470_11769 , \11471_11770 , \11472_11771 , \11473_11772 , \11474_11773 , \11475_11774 , \11476_11775 ,
         \11477_11776 , \11478_11777 , \11479_11778 , \11480_11779 , \11481_11780 , \11482_11781 , \11483_11782 , \11484_11783 , \11485_11784 , \11486_11785 ,
         \11487_11786 , \11488_11787 , \11489_11788 , \11490_11789 , \11491_11790 , \11492_11791 , \11493_11792 , \11494_11793 , \11495_11794 , \11496_11795 ,
         \11497_11796 , \11498_11797 , \11499_11798 , \11500_11799 , \11501_11800 , \11502_11801 , \11503_11802 , \11504_11803 , \11505_11804 , \11506_11805 ,
         \11507_11806 , \11508_11807 , \11509_11808 , \11510_11809 , \11511_11810 , \11512_11811 , \11513_11812 , \11514_11813 , \11515_11814 , \11516_11815 ,
         \11517_11816 , \11518_11817 , \11519_11818 , \11520_11819 , \11521_11820 , \11522_11821 , \11523_11822 , \11524_11823 , \11525_11824 , \11526_11825 ,
         \11527_11826 , \11528_11827 , \11529_11828 , \11530_11829 , \11531_11830 , \11532_11831 , \11533_11832 , \11534_11833 , \11535_11834 , \11536_11835 ,
         \11537_11836 , \11538_11837 , \11539_11838 , \11540_11839 , \11541_11840 , \11542_11841 , \11543_11842 , \11544_11843 , \11545_11844 , \11546_11845 ,
         \11547_11846 , \11548_11847 , \11549_11848 , \11550_11849 , \11551_11850 , \11552_11851 , \11553_11852 , \11554_11853 , \11555_11854 , \11556_11855 ,
         \11557_11856 , \11558_11857 , \11559_11858 , \11560_11859 , \11561_11860 , \11562_11861 , \11563_11862 , \11564_11863 , \11565_11864 , \11566_11865 ,
         \11567_11866 , \11568_11867 , \11569_11868 , \11570_11869 , \11571 , \11572_11871 , \11573_11872 , \11574_11873 , \11575_11874 , \11576_11875 ,
         \11577_11876 , \11578_11877 , \11579_11878 , \11580_11879 , \11581_11880 , \11582_11881 , \11583_11882 , \11584_11883 , \11585_11884 , \11586_11885 ,
         \11587_11886 , \11588_11887 , \11589_11888 , \11590_11889 , \11591_11890 , \11592_11891 , \11593_11892 , \11594_11893 , \11595_11894 , \11596_11895 ,
         \11597_11896 , \11598_11897 , \11599_11898 , \11600_11899 , \11601_11900 , \11602_11901 , \11603_11902 , \11604_11903 , \11605_11904 , \11606_11905 ,
         \11607_11906 , \11608_11907 , \11609_11908 , \11610_11909 , \11611_11910 , \11612_11911 , \11613_11912 , \11614_11913 , \11615_11914 , \11616_11915 ,
         \11617_11916 , \11618_11917 , \11619_11918 , \11620_11919 , \11621_11920 , \11622_11921 , \11623_11922 , \11624_11923 , \11625_11924 , \11626_11925 ,
         \11627_11926 , \11628_11927 , \11629_11928 , \11630_11929 , \11631_11930 , \11632_11931 , \11633_11932 , \11634_11933 , \11635_11934 , \11636_11935 ,
         \11637_11936 , \11638_11937 , \11639_11938 , \11640_11939 , \11641_11940 , \11642_11941 , \11643_11942 , \11644_11943 , \11645_11944 , \11646_11945 ,
         \11647_11946 , \11648_11947 , \11649_11948 , \11650_11949 , \11651_11950 , \11652_11951 , \11653_11952 , \11654_11953 , \11655_11954 , \11656_11955 ,
         \11657_11956 , \11658_11957 , \11659_11958 , \11660_11959 , \11661_11960 , \11662_11961 , \11663_11962 , \11664_11963 , \11665_11964 , \11666_11965 ,
         \11667_11966 , \11668_11967 , \11669_11968 , \11670_11969 , \11671_11970 , \11672_11971 , \11673_11972 , \11674_11973 , \11675_11974 , \11676_11975 ,
         \11677_11976 , \11678_11977 , \11679_11978 , \11680_11979 , \11681_11980 , \11682_11981 , \11683_11982 , \11684_11983 , \11685_11984 , \11686_11985 ,
         \11687_11986 , \11688_11987 , \11689_11988 , \11690_11989 , \11691_11990 , \11692_11991 , \11693_11992 , \11694_11993 , \11695_11994 , \11696_11995 ,
         \11697_11996 , \11698_11997 , \11699_11998 , \11700_11999 , \11701_12000 , \11702_12001 , \11703_12002 , \11704_12003 , \11705 , \11706_12005 ,
         \11707_12006 , \11708_12007 , \11709_12008 , \11710_12009 , \11711_12010 , \11712_12011 , \11713_12012 , \11714_12013 , \11715_12014 , \11716_12015 ,
         \11717_12016 , \11718_12017 , \11719_12018 , \11720_12019 , \11721_12020 , \11722_12021 , \11723_12022 , \11724_12023 , \11725_12024 , \11726_12025 ,
         \11727_12026 , \11728_12027 , \11729_12028 , \11730_12029 , \11731_12030 , \11732_12031 , \11733_12032 , \11734_12033 , \11735_12034 , \11736_12035 ,
         \11737_12036 , \11738_12037 , \11739_12038 , \11740_12039 , \11741_12040 , \11742_12041 , \11743_12042 , \11744_12043 , \11745_12044 , \11746_12045 ,
         \11747_12046 , \11748_12047 , \11749_12048 , \11750_12049 , \11751_12050 , \11752_12051 , \11753_12052 , \11754_12053 , \11755_12054 , \11756_12055 ,
         \11757_12056 , \11758_12057 , \11759_12058 , \11760_12059 , \11761_12060 , \11762_12061 , \11763_12062 , \11764_12063 , \11765_12064 , \11766_12065 ,
         \11767_12066 , \11768_12067 , \11769_12068 , \11770_12069 , \11771_12070 , \11772_12071 , \11773_12072 , \11774_12073 , \11775_12074 , \11776_12075 ,
         \11777_12076 , \11778_12077 , \11779_12078 , \11780_12079 , \11781_12080 , \11782_12081 , \11783_12082 , \11784_12083 , \11785_12084 , \11786_12085 ,
         \11787_12086 , \11788_12087 , \11789_12088 , \11790_12089 , \11791_12090 , \11792_12091 , \11793_12092 , \11794_12093 , \11795_12094 , \11796_12095 ,
         \11797_12096 , \11798_12097 , \11799_12098 , \11800_12099 , \11801_12100 , \11802_12101 , \11803_12102 , \11804_12103 , \11805_12104 , \11806_12105 ,
         \11807_12106 , \11808_12107 , \11809_12108 , \11810_12109 , \11811_12110 , \11812_12111 , \11813_12112 , \11814_12113 , \11815_12114 , \11816_12115 ,
         \11817_12116 , \11818_12117 , \11819_12118 , \11820_12119 , \11821_12120 , \11822_12121 , \11823_12122 , \11824_12123 , \11825_12124 , \11826_12125 ,
         \11827_12126 , \11828_12127 , \11829_12128 , \11830_12129 , \11831_12130 , \11832_12131 , \11833_12132 , \11834_12133 , \11835_12134 , \11836_12135 ,
         \11837_12136 , \11838 , \11839_12138 , \11840_12139 , \11841_12140 , \11842_12141 , \11843_12142 , \11844_12143 , \11845_12144 , \11846_12145 ,
         \11847_12146 , \11848_12147 , \11849_12148_nG4448 , \11850_12149 , \11851_12150 , \11852_12151_nG444b , \11853_12152 , \11854_12153 , \11855_12154 , \11856_12158 ,
         \11857_12159 , \11858_12160 , \11859_12161 , \11860_12162 , \11861_12163 , \11862_12164 , \11863_12165 , \11864_12166 , \11865_12167 , \11866_12168 ,
         \11867_12169 , \11868_12170 , \11869_12171 , \11870_12172 , \11871_12173 , \11872_12174 , \11873_12175 , \11874_12176 , \11875_12177 , \11876_12178 ,
         \11877_12179 , \11878_12180 , \11879_12181 , \11880_12182 , \11881_12183 , \11882_12184 , \11883_12185 , \11884_12186 , \11885_12187 , \11886_12188 ,
         \11887_12189 , \11888_12190 , \11889_12191 , \11890_12192 , \11891_12193 , \11892_12194 , \11893_12195 , \11894_12196 , \11895_12197 , \11896_12198 ,
         \11897_12199 , \11898_12200 , \11899_12201 , \11900_12202 , \11901_12203 , \11902_12204 , \11903_12205 , \11904_12206 , \11905_12207 , \11906_12208 ,
         \11907_12209 , \11908_12210 , \11909_12211 , \11910_12212 , \11911_12213 , \11912_12214 , \11913_12215 , \11914_12216 , \11915_12217 , \11916_12218 ,
         \11917_12219 , \11918_12220 , \11919_12221 , \11920_12222 , \11921_12223 , \11922_12224 , \11923_12225 , \11924_12226 , \11925_12227 , \11926_12228 ,
         \11927_12229 , \11928_12230 , \11929_12231 , \11930_12232 , \11931_12233 , \11932_12234 , \11933_12235 , \11934_12236 , \11935_12237 , \11936_12238 ,
         \11937_12239 , \11938_12240 , \11939_12241 , \11940_12242 , \11941_12243 , \11942_12244 , \11943_12245 , \11944_12246 , \11945_12247 , \11946_12248 ,
         \11947_12249 , \11948_12250 , \11949_12251 , \11950_12252 , \11951_12253 , \11952_12254 , \11953_12255 , \11954_12256 , \11955_12257 , \11956_12258 ,
         \11957_12259 , \11958_12260 , \11959_12261 , \11960_12262 , \11961_12263 , \11962_12264 , \11963_12265 , \11964_12266 , \11965_12267 , \11966_12268 ,
         \11967_12269 , \11968_12270 , \11969_12271 , \11970_12272 , \11971_12273 , \11972_12274 , \11973_12275 , \11974_12276 , \11975_12277 , \11976_12278 ,
         \11977_12279 , \11978_12280 , \11979_12281 , \11980_12282 , \11981_12283 , \11982_12284 , \11983_12285 , \11984_12286 , \11985_12287 , \11986_12288 ,
         \11987_12289 , \11988_12290 , \11989_12291 , \11990_12292 , \11991_12293 , \11992_12294 , \11993_12295 , \11994_12296 , \11995_12297 , \11996_12298 ,
         \11997_12299 , \11998_12300 , \11999_12301 , \12000_12302 , \12001_12303 , \12002_12304 , \12003_12305 , \12004_12306 , \12005_12307 , \12006_12308 ,
         \12007_12309 , \12008_12310 , \12009_12311 , \12010_12312 , \12011_12313 , \12012 , \12013_12315 , \12014_12316 , \12015_12317 , \12016_12318 ,
         \12017_12319 , \12018_12320 , \12019_12321 , \12020_12322 , \12021_12323 , \12022_12324 , \12023_12325 , \12024_12326 , \12025_12327 , \12026_12328 ,
         \12027_12329 , \12028_12330 , \12029_12331 , \12030_12332 , \12031_12333 , \12032_12334 , \12033_12335 , \12034_12336 , \12035_12337 , \12036_12338 ,
         \12037_12339 , \12038_12340 , \12039_12341 , \12040_12342 , \12041_12343 , \12042_12344 , \12043_12345 , \12044_12346 , \12045_12347 , \12046_12348 ,
         \12047_12349 , \12048_12350 , \12049_12351 , \12050_12352 , \12051_12353 , \12052_12354 , \12053_12355 , \12054_12356 , \12055_12357 , \12056_12358 ,
         \12057_12359 , \12058_12360 , \12059_12361 , \12060_12362 , \12061_12363 , \12062_12364 , \12063_12365 , \12064_12366 , \12065_12367 , \12066_12368 ,
         \12067_12369 , \12068_12370 , \12069_12371 , \12070_12372 , \12071_12373 , \12072_12374 , \12073_12375 , \12074_12376 , \12075_12377 , \12076_12378 ,
         \12077_12379 , \12078_12380 , \12079_12381 , \12080_12382 , \12081_12383 , \12082_12384 , \12083_12385 , \12084_12386 , \12085_12387 , \12086_12388 ,
         \12087_12389 , \12088_12390 , \12089_12391 , \12090_12392 , \12091_12393 , \12092_12394 , \12093_12395 , \12094_12396 , \12095_12397 , \12096_12398 ,
         \12097_12399 , \12098_12400 , \12099_12401 , \12100_12402 , \12101_12403 , \12102_12404 , \12103_12405 , \12104_12406 , \12105_12407 , \12106_12408 ,
         \12107_12409 , \12108_12410 , \12109_12411 , \12110_12412 , \12111_12413 , \12112_12414 , \12113_12415 , \12114_12416 , \12115_12417 , \12116_12418 ,
         \12117_12419 , \12118_12420 , \12119_12421 , \12120_12422 , \12121_12423 , \12122_12424 , \12123_12425 , \12124_12426 , \12125_12427 , \12126_12428 ,
         \12127_12429 , \12128_12430 , \12129_12431 , \12130_12432 , \12131_12433 , \12132_12434 , \12133_12435 , \12134_12436 , \12135_12437 , \12136_12438 ,
         \12137_12439 , \12138_12440 , \12139_12441 , \12140_12442 , \12141_12443 , \12142_12444 , \12143_12445 , \12144 , \12145_12447_nG6585 , \12146_12448 ,
         \12147_12449 , \12148_12450 , \12149_12451 , \12150_12452 , \12151_12453 , \12152_12454 , \12153_12455 , \12154_12456 , \12155 , \12156 ,
         \12157_12459_nG4983 , \12158_12460 , \12159_12461 , \12160_12462 , \12161_12463 , \12162_12464 , \12163_12465 , \12164_12466 , \12165_12467 , \12166_12468 ,
         \12167_12469 , \12168_12470_nG9c02 , \12169_12471 , \12170_12472 , \12171_12473 , \12172_12474 , \12173_12475 , \12174_12476 , \12175_12477 , \12176_12478 ,
         \12177_12479 , \12178_12480 , \12179_12481 , \12180_12482 , \12181_12155 , \12182_12156 , \12183_12157 , \12184_12483 , \12185_12484 , \12186_12485 ,
         \12187_12486 , \12188_12487 , \12189_12488 , \12190_12489 , \12191_12490 , \12192_12491 , \12193_12492 , \12194_12493 , \12195_12494 , \12196_12495 ,
         \12197_12496 , \12198_12497 , \12199_12498 , \12200_12499 , \12201_12500 , \12202_12501 , \12203_12502 , \12204_12503 , \12205_12504 , \12206_12505 ,
         \12207_12506 , \12208_12507 , \12209_12508 , \12210_12509 , \12211_12510 , \12212_12511 , \12213_12512 , \12214_12513 , \12215_12514 , \12216_12515 ,
         \12217_12516 , \12218_12517 , \12219_12518 , \12220_12519 , \12221_12520 , \12222_12521 , \12223_12522 , \12224_12523 , \12225_12524 , \12226_12525 ,
         \12227_12526 , \12228_12527 , \12229_12528 , \12230_12529 , \12231_12530 , \12232_12531 , \12233_12532 , \12234_12533 , \12235_12534 , \12236_12535 ,
         \12237_12536 , \12238_12537 , \12239_12538 , \12240_12539 , \12241_12540 , \12242_12541 , \12243_12542 , \12244_12543 , \12245_12544 , \12246_12545 ,
         \12247_12546 , \12248_12547 , \12249_12548 , \12250_12549 , \12251_12550 , \12252_12551 , \12253_12552 , \12254_12553 , \12255_12554 , \12256_12555 ,
         \12257_12556 , \12258_12557 , \12259_12558 , \12260_12559 , \12261_12560 , \12262_12561 , \12263_12562 , \12264_12563 , \12265_12564 , \12266_12565 ,
         \12267_12566 , \12268_12567 , \12269_12568 , \12270_12569 , \12271_12570 , \12272_12571 , \12273_12572 , \12274_12573 , \12275_12574 , \12276_12575 ,
         \12277_12576 , \12278_12577 , \12279_12578 , \12280_12579 , \12281_12580 , \12282_12581 , \12283_12582 , \12284_12583 , \12285_12584 , \12286_12585 ,
         \12287_12586 , \12288_12587 , \12289_12588 , \12290_12589 , \12291_12590 , \12292_12591 , \12293_12592 , \12294_12593 , \12295_12594 , \12296_12595 ,
         \12297_12596 , \12298_12597 , \12299_12598 , \12300_12599 , \12301_12600 , \12302_12601 , \12303_12602 , \12304_12603 , \12305_12604 , \12306_12605 ,
         \12307_12606 , \12308_12607 , \12309_12608 , \12310_12609 , \12311_12610 , \12312_12611 , \12313_12612 , \12314_12613 , \12315_12614 , \12316_12615 ,
         \12317_12616 , \12318_12617 , \12319_12618 , \12320_12619 , \12321_12620 , \12322_12621 , \12323_12622 , \12324_12623 , \12325_12624 , \12326_12625 ,
         \12327_12626 , \12328_12627 , \12329_12628 , \12330_12629 , \12331_12630 , \12332_12631 , \12333_12632 , \12334_12633 , \12335_12634 , \12336 ,
         \12337_12636 , \12338_12637 , \12339_12638 , \12340_12639 , \12341_12640 , \12342_12641 , \12343_12642 , \12344_12643 , \12345_12644 , \12346_12645 ,
         \12347_12646 , \12348_12647 , \12349_12648 , \12350_12649 , \12351_12650 , \12352_12651 , \12353_12652 , \12354_12653 , \12355_12654 , \12356_12655 ,
         \12357_12656 , \12358_12657 , \12359_12658 , \12360_12659 , \12361_12660 , \12362_12661 , \12363_12662 , \12364_12663 , \12365_12664 , \12366_12665 ,
         \12367_12666 , \12368_12667 , \12369_12668 , \12370_12669 , \12371_12670 , \12372_12671 , \12373_12672 , \12374_12673 , \12375_12674 , \12376_12675 ,
         \12377_12676 , \12378_12677 , \12379_12678 , \12380_12679 , \12381_12680 , \12382_12681 , \12383_12682 , \12384_12683 , \12385_12684 , \12386_12685 ,
         \12387_12686 , \12388_12687 , \12389_12688 , \12390_12689 , \12391_12690 , \12392_12691 , \12393_12692 , \12394_12693 , \12395_12694 , \12396_12695 ,
         \12397_12696 , \12398_12697 , \12399_12698 , \12400_12699 , \12401_12700 , \12402_12701 , \12403_12702 , \12404_12703 , \12405_12704 , \12406_12705 ,
         \12407_12706 , \12408_12707 , \12409_12708 , \12410_12709 , \12411_12710 , \12412_12711 , \12413_12712 , \12414_12713 , \12415_12714 , \12416_12715 ,
         \12417_12716 , \12418_12717 , \12419_12718 , \12420_12719 , \12421_12720 , \12422_12721 , \12423_12722 , \12424_12723 , \12425_12724 , \12426_12725 ,
         \12427_12726 , \12428_12727 , \12429_12728 , \12430_12729 , \12431_12730 , \12432_12731 , \12433_12732 , \12434_12733 , \12435_12734 , \12436_12735 ,
         \12437_12736 , \12438_12737 , \12439_12738 , \12440_12739 , \12441_12740 , \12442_12741 , \12443_12742 , \12444_12743 , \12445_12744 , \12446_12745 ,
         \12447_12746 , \12448_12747 , \12449_12748 , \12450_12749 , \12451_12750 , \12452_12751 , \12453_12752 , \12454_12753 , \12455_12754 , \12456_12755 ,
         \12457_12756 , \12458_12757 , \12459_12758 , \12460_12759 , \12461_12760 , \12462_12761 , \12463_12762 , \12464_12763 , \12465_12764 , \12466_12765 ,
         \12467_12766 , \12468 , \12469_12768_nG6588 , \12470_12769 , \12471_12770 , \12472_12771 , \12473_12772 , \12474_12773 , \12475 , \12476 ,
         \12477_12776_nG4a8c , \12478_12777 , \12479_12778 , \12480_12779 , \12481_12780 , \12482_12781 , \12483_12782 , \12484_12783 , \12485_12784 , \12486_12785 ,
         \12487_12786 , \12488_12787 , \12489_12788 , \12490_12789 , \12491_12790 , \12492_12791 , \12493_12792 , \12494_12793 , \12495_12794 , \12496_12795 ,
         \12497_12796 , \12498_12797 , \12499_12798 , \12500_12799 , \12501_12800 , \12502_12801_nG9bff , \12503_12802 , \12504_12803 , \12505_12804 , \12506_12805 ,
         \12507_12806 , \12508_12807 , \12509_12808 , \12510_12809 , \12511_12810 , \12512_12811 , \12513_12812 , \12514_12813 , \12515_12814 , \12516_12815 ,
         \12517_12816 , \12518_12817 , \12519_12818 , \12520_12819 , \12521_12820 , \12522_12821 , \12523_12822 , \12524_12823 , \12525_12824 , \12526_12825 ,
         \12527_12826 , \12528_12827 , \12529_12828 , \12530_12829 , \12531_12830 , \12532_12831 , \12533_12832 , \12534_12833 , \12535_12834 , \12536_12835 ,
         \12537_12836 , \12538_12837 , \12539_12838 , \12540_12839 , \12541_12840 , \12542_12841 , \12543_12842 , \12544_12843 , \12545_12844 , \12546_12845 ,
         \12547_12846 , \12548_12847 , \12549_12848 , \12550_12849 , \12551_12850 , \12552_12851 , \12553_12852 , \12554_12853 , \12555_12854 , \12556_12855 ,
         \12557_12856 , \12558_12857 , \12559_12858 , \12560_12859 , \12561_12860 , \12562_12861 , \12563_12862 , \12564_12863 , \12565_12864 , \12566_12865 ,
         \12567_12866 , \12568_12867 , \12569_12868 , \12570_12869 , \12571_12870 , \12572_12871 , \12573_12872 , \12574_12873 , \12575_12874 , \12576_12875 ,
         \12577_12876 , \12578_12877 , \12579_12878 , \12580_12879 , \12581_12880 , \12582_12881 , \12583_12882 , \12584_12883 , \12585_12884 , \12586_12885 ,
         \12587_12886 , \12588_12887 , \12589_12888 , \12590_12889 , \12591_12890 , \12592_12891 , \12593_12892 , \12594_12893 , \12595_12894 , \12596_12895 ,
         \12597_12896 , \12598_12897 , \12599_12898 , \12600_12899 , \12601_12900 , \12602_12901 , \12603_12902 , \12604_12903 , \12605_12904 , \12606_12905 ,
         \12607_12906 , \12608_12907 , \12609_12908 , \12610_12909 , \12611_12910 , \12612_12911 , \12613_12912 , \12614_12913 , \12615_12914 , \12616_12915 ,
         \12617_12916 , \12618_12917 , \12619_12918 , \12620_12919 , \12621_12920 , \12622_12921 , \12623_12922 , \12624_12923 , \12625_12924 , \12626_12925 ,
         \12627_12926 , \12628_12927 , \12629_12928 , \12630_12929 , \12631_12930 , \12632_12931 , \12633_12932 , \12634_12933 , \12635_12934 , \12636_12935 ,
         \12637_12936 , \12638_12937 , \12639_12938 , \12640_12939 , \12641_12940 , \12642_12941 , \12643_12942 , \12644_12943 , \12645_12944 , \12646_12945 ,
         \12647_12946 , \12648_12947 , \12649_12948 , \12650_12949 , \12651 , \12652_12951 , \12653_12952 , \12654_12953 , \12655_12954 , \12656_12955 ,
         \12657_12956 , \12658_12957 , \12659_12958 , \12660_12959 , \12661_12960 , \12662_12961 , \12663_12962 , \12664_12963 , \12665_12964 , \12666_12965 ,
         \12667_12966 , \12668_12967 , \12669_12968 , \12670_12969 , \12671_12970 , \12672_12971 , \12673_12972 , \12674_12973 , \12675_12974 , \12676_12975 ,
         \12677_12976 , \12678_12977 , \12679_12978 , \12680_12979 , \12681_12980 , \12682_12981 , \12683_12982 , \12684_12983 , \12685_12984 , \12686_12985 ,
         \12687_12986 , \12688_12987 , \12689_12988 , \12690_12989 , \12691_12990 , \12692_12991 , \12693_12992 , \12694_12993 , \12695_12994 , \12696_12995 ,
         \12697_12996 , \12698_12997 , \12699_12998 , \12700_12999 , \12701_13000 , \12702_13001 , \12703_13002 , \12704_13003 , \12705_13004 , \12706_13005 ,
         \12707_13006 , \12708_13007 , \12709_13008 , \12710_13009 , \12711_13010 , \12712_13011 , \12713_13012 , \12714_13013 , \12715_13014 , \12716_13015 ,
         \12717_13016 , \12718_13017 , \12719_13018 , \12720_13019 , \12721_13020 , \12722_13021 , \12723_13022 , \12724_13023 , \12725_13024 , \12726_13025 ,
         \12727_13026 , \12728_13027 , \12729_13028 , \12730_13029 , \12731_13030 , \12732_13031 , \12733_13032 , \12734_13033 , \12735_13034 , \12736_13035 ,
         \12737_13036 , \12738_13037 , \12739_13038 , \12740_13039 , \12741_13040 , \12742_13041 , \12743_13042 , \12744_13043 , \12745_13044 , \12746_13045 ,
         \12747_13046 , \12748_13047 , \12749_13048 , \12750_13049 , \12751_13050 , \12752_13051 , \12753_13052 , \12754_13053 , \12755_13054 , \12756_13055 ,
         \12757_13056 , \12758_13057 , \12759_13058 , \12760_13059 , \12761_13060 , \12762_13061 , \12763_13062 , \12764_13063 , \12765_13064 , \12766_13065 ,
         \12767_13066 , \12768_13067 , \12769_13068 , \12770_13069 , \12771_13070 , \12772_13071 , \12773_13072 , \12774_13073 , \12775_13074 , \12776_13075 ,
         \12777_13076 , \12778_13077 , \12779_13078 , \12780_13079 , \12781_13080 , \12782_13081 , \12783_13082 , \12784 , \12785_13084 , \12786_13085 ,
         \12787_13086 , \12788_13087 , \12789_13088 , \12790_13089 , \12791_13090 , \12792_13091 , \12793_13092 , \12794_13093 , \12795_13094 , \12796_13095 ,
         \12797_13096 , \12798_13097 , \12799_13098 , \12800_13099 , \12801_13100 , \12802_13101 , \12803_13102 , \12804_13103 , \12805_13104 , \12806_13105 ,
         \12807_13106 , \12808_13107 , \12809_13108 , \12810_13109 , \12811_13110 , \12812_13111 , \12813_13112 , \12814_13113 , \12815_13114 , \12816_13115 ,
         \12817_13116 , \12818_13117 , \12819_13118 , \12820_13119 , \12821_13120 , \12822_13121 , \12823_13122 , \12824_13123 , \12825_13124 , \12826_13125 ,
         \12827_13126 , \12828_13127 , \12829_13128 , \12830_13129 , \12831_13130 , \12832_13131 , \12833_13132 , \12834_13133 , \12835_13134 , \12836_13135 ,
         \12837_13136 , \12838_13137 , \12839_13138 , \12840_13139 , \12841_13140 , \12842_13141 , \12843_13142 , \12844_13143 , \12845_13144 , \12846_13145 ,
         \12847_13146 , \12848_13147 , \12849_13148 , \12850_13149 , \12851_13150 , \12852_13151 , \12853_13152 , \12854_13153 , \12855_13154 , \12856_13155 ,
         \12857_13156 , \12858_13157 , \12859_13158 , \12860_13159 , \12861_13160 , \12862_13161 , \12863_13162 , \12864_13163 , \12865_13164 , \12866_13165 ,
         \12867_13166 , \12868_13167 , \12869_13168 , \12870_13169 , \12871_13170 , \12872_13171 , \12873_13172 , \12874_13173 , \12875_13174 , \12876_13175 ,
         \12877_13176 , \12878_13177 , \12879_13178 , \12880_13179 , \12881_13180 , \12882_13181 , \12883_13182 , \12884_13183 , \12885_13184 , \12886_13185 ,
         \12887_13186 , \12888_13187 , \12889_13188 , \12890_13189 , \12891_13190 , \12892_13191 , \12893_13192 , \12894_13193 , \12895_13194 , \12896_13195 ,
         \12897_13196 , \12898_13197 , \12899_13198 , \12900_13199 , \12901_13200 , \12902_13201 , \12903_13202 , \12904_13203 , \12905_13204 , \12906_13205 ,
         \12907_13206 , \12908_13207 , \12909_13208 , \12910_13209 , \12911_13210 , \12912_13211 , \12913_13212 , \12914_13213 , \12915_13214 , \12916_13215 ,
         \12917_13216 , \12918 , \12919_13218 , \12920_13219 , \12921_13220 , \12922_13221 , \12923_13222 , \12924_13223 , \12925_13224 , \12926_13225 ,
         \12927_13226 , \12928_13227 , \12929_13228 , \12930_13229 , \12931_13230 , \12932_13231 , \12933_13232 , \12934_13233 , \12935_13234 , \12936_13235 ,
         \12937_13236 , \12938_13237 , \12939_13238 , \12940_13239 , \12941_13240 , \12942_13241 , \12943_13242 , \12944_13243 , \12945_13244 , \12946_13245 ,
         \12947_13246 , \12948_13247 , \12949_13248 , \12950_13249 , \12951_13250 , \12952_13251 , \12953_13252 , \12954_13253 , \12955_13254 , \12956_13255 ,
         \12957_13256 , \12958_13257 , \12959_13258 , \12960_13259 , \12961_13260 , \12962_13261 , \12963_13262 , \12964_13263 , \12965_13264 , \12966_13265 ,
         \12967_13266 , \12968_13267 , \12969_13268 , \12970_13269 , \12971_13270 , \12972_13271 , \12973_13272 , \12974_13273 , \12975_13274 , \12976_13275 ,
         \12977_13276 , \12978_13277 , \12979_13278 , \12980_13279 , \12981_13280 , \12982_13281 , \12983_13282 , \12984_13283 , \12985_13284 , \12986_13285 ,
         \12987_13286 , \12988_13287 , \12989_13288 , \12990_13289 , \12991_13290 , \12992_13291 , \12993_13292 , \12994_13293 , \12995_13294 , \12996_13295 ,
         \12997_13296 , \12998_13297 , \12999_13298 , \13000_13299 , \13001_13300 , \13002_13301 , \13003_13302 , \13004_13303 , \13005_13304 , \13006_13305 ,
         \13007_13306 , \13008_13307 , \13009_13308 , \13010_13309 , \13011_13310 , \13012_13311 , \13013_13312 , \13014_13313 , \13015_13314 , \13016_13315 ,
         \13017_13316 , \13018_13317 , \13019_13318 , \13020_13319 , \13021_13320 , \13022_13321 , \13023_13322 , \13024_13323 , \13025_13324 , \13026_13325 ,
         \13027_13326 , \13028_13327 , \13029_13328 , \13030_13329 , \13031_13330 , \13032_13331 , \13033_13332 , \13034_13333 , \13035_13334 , \13036_13335 ,
         \13037_13336 , \13038_13337 , \13039_13338 , \13040_13339 , \13041_13340 , \13042_13341 , \13043_13342 , \13044_13343 , \13045_13344 , \13046_13345 ,
         \13047_13346 , \13048_13347 , \13049_13348 , \13050_13349 , \13051 , \13052_13351 , \13053_13352 , \13054_13353 , \13055_13354 , \13056_13355 ,
         \13057_13356 , \13058_13357 , \13059_13358 , \13060_13359 , \13061_13360 , \13062_13361_nG4442 , \13063_13362 , \13064_13363 , \13065_13364_nG4445 , \13066_13365 ,
         \13067_13366 , \13068_13367 , \13069_13371 , \13070_13372 , \13071_13373 , \13072_13374 , \13073_13375 , \13074_13376 , \13075_13377 , \13076_13378 ,
         \13077_13379 , \13078_13380 , \13079_13381 , \13080_13382 , \13081_13383 , \13082_13384 , \13083_13385 , \13084_13386 , \13085_13387 , \13086_13388 ,
         \13087_13389 , \13088_13390 , \13089_13391 , \13090_13392 , \13091_13393 , \13092_13394 , \13093_13395 , \13094_13396 , \13095_13397 , \13096_13398 ,
         \13097_13399 , \13098_13400 , \13099_13401 , \13100_13402 , \13101_13403 , \13102_13404 , \13103_13405 , \13104_13406 , \13105_13407 , \13106_13408 ,
         \13107_13409 , \13108_13410 , \13109_13411 , \13110_13412 , \13111_13413 , \13112_13414 , \13113_13415 , \13114_13416 , \13115_13417 , \13116_13418 ,
         \13117_13419 , \13118_13420 , \13119_13421 , \13120_13422 , \13121_13423 , \13122_13424 , \13123_13425 , \13124_13426 , \13125_13427 , \13126_13428 ,
         \13127_13429 , \13128_13430 , \13129_13431 , \13130_13432 , \13131_13433 , \13132_13434 , \13133_13435 , \13134_13436 , \13135_13437 , \13136_13438 ,
         \13137_13439 , \13138_13440 , \13139_13441 , \13140_13442 , \13141_13443 , \13142_13444 , \13143_13445 , \13144_13446 , \13145_13447 , \13146_13448 ,
         \13147_13449 , \13148_13450 , \13149_13451 , \13150_13452 , \13151_13453 , \13152_13454 , \13153_13455 , \13154_13456 , \13155_13457 , \13156_13458 ,
         \13157_13459 , \13158_13460 , \13159_13461 , \13160_13462 , \13161_13463 , \13162_13464 , \13163_13465 , \13164_13466 , \13165_13467 , \13166_13468 ,
         \13167_13469 , \13168_13470 , \13169_13471 , \13170_13472 , \13171_13473 , \13172_13474 , \13173_13475 , \13174_13476 , \13175_13477 , \13176_13478 ,
         \13177_13479 , \13178_13480 , \13179_13481 , \13180_13482 , \13181_13483 , \13182_13484 , \13183_13485 , \13184_13486 , \13185_13487 , \13186_13488 ,
         \13187_13489 , \13188_13490 , \13189_13491 , \13190_13492 , \13191_13493 , \13192_13494 , \13193_13495 , \13194_13496 , \13195_13497 , \13196_13498 ,
         \13197_13499 , \13198_13500 , \13199_13501 , \13200_13502 , \13201_13503 , \13202_13504 , \13203_13505 , \13204_13506 , \13205_13507 , \13206_13508 ,
         \13207_13509 , \13208_13510 , \13209_13511 , \13210_13512 , \13211_13513 , \13212_13514 , \13213_13515 , \13214_13516 , \13215_13517 , \13216_13518 ,
         \13217_13519 , \13218_13520 , \13219_13521 , \13220_13522 , \13221_13523 , \13222_13524 , \13223_13525 , \13224_13526 , \13225_13527 , \13226_13528 ,
         \13227_13529 , \13228_13530 , \13229_13531 , \13230_13532 , \13231_13533 , \13232_13534 , \13233_13535 , \13234_13536 , \13235_13537 , \13236_13538 ,
         \13237_13539 , \13238_13540 , \13239_13541 , \13240_13542 , \13241_13543 , \13242_13544 , \13243 , \13244_13546 , \13245_13547 , \13246_13548 ,
         \13247_13549 , \13248_13550 , \13249_13551 , \13250_13552 , \13251_13553 , \13252_13554 , \13253_13555 , \13254_13556 , \13255_13557 , \13256_13558 ,
         \13257_13559 , \13258_13560 , \13259_13561 , \13260_13562 , \13261_13563 , \13262_13564 , \13263_13565 , \13264_13566 , \13265_13567 , \13266_13568 ,
         \13267_13569 , \13268_13570 , \13269_13571 , \13270_13572 , \13271_13573 , \13272_13574 , \13273_13575 , \13274_13576 , \13275_13577 , \13276_13578 ,
         \13277_13579 , \13278_13580 , \13279_13581 , \13280_13582 , \13281_13583 , \13282_13584 , \13283_13585 , \13284_13586 , \13285_13587 , \13286_13588 ,
         \13287_13589 , \13288_13590 , \13289_13591 , \13290_13592 , \13291_13593 , \13292_13594 , \13293_13595 , \13294_13596 , \13295_13597 , \13296_13598 ,
         \13297_13599 , \13298_13600 , \13299_13601 , \13300_13602 , \13301_13603 , \13302_13604 , \13303_13605 , \13304_13606 , \13305_13607 , \13306_13608 ,
         \13307_13609 , \13308_13610 , \13309_13611 , \13310_13612 , \13311_13613 , \13312_13614 , \13313_13615 , \13314_13616 , \13315_13617 , \13316_13618 ,
         \13317_13619 , \13318_13620 , \13319_13621 , \13320_13622 , \13321_13623 , \13322_13624 , \13323_13625 , \13324_13626 , \13325_13627 , \13326_13628 ,
         \13327_13629 , \13328_13630 , \13329_13631 , \13330_13632 , \13331_13633 , \13332_13634 , \13333_13635 , \13334_13636 , \13335_13637 , \13336_13638 ,
         \13337_13639 , \13338_13640 , \13339_13641 , \13340_13642 , \13341_13643 , \13342_13644 , \13343_13645 , \13344_13646 , \13345_13647 , \13346_13648 ,
         \13347_13649 , \13348_13650 , \13349_13651 , \13350_13652 , \13351_13653 , \13352_13654 , \13353_13655 , \13354_13656 , \13355_13657 , \13356_13658 ,
         \13357_13659 , \13358_13660 , \13359_13661 , \13360_13662 , \13361_13663 , \13362_13664 , \13363_13665 , \13364_13666 , \13365_13667 , \13366_13668 ,
         \13367_13669 , \13368_13670 , \13369_13671 , \13370_13672 , \13371_13673 , \13372_13674 , \13373_13675 , \13374_13676 , \13375 , \13376_13678_nG658b ,
         \13377_13679 , \13378_13680 , \13379_13681 , \13380_13682 , \13381_13683 , \13382_13684 , \13383_13685 , \13384_13686 , \13385_13687 , \13386 ,
         \13387 , \13388_13690_nG4b95 , \13389_13691 , \13390_13692 , \13391_13693 , \13392_13694 , \13393_13695 , \13394_13696 , \13395_13697 , \13396_13698 ,
         \13397_13699 , \13398_13700 , \13399_13701 , \13400_13702 , \13401_13703 , \13402_13704 , \13403_13705_nG9bfc , \13404_13706 , \13405_13707 , \13406_13708 ,
         \13407_13709 , \13408_13710 , \13409_13711 , \13410_13712 , \13411_13713 , \13412_13714 , \13413_13715 , \13414_13716 , \13415_13717 , \13416_13718 ,
         \13417_13719 , \13418_13720 , \13419_13721 , \13420_13722 , \13421_13723 , \13422_13724 , \13423_13725 , \13424_13726 , \13425_13727 , \13426_13728 ,
         \13427_13729 , \13428_13730 , \13429_13368 , \13430_13369 , \13431_13370 , \13432_13731 , \13433_13732 , \13434_13733 , \13435_13734 , \13436_13735 ,
         \13437_13736 , \13438_13737 , \13439_13738 , \13440_13739 , \13441_13740 , \13442_13741 , \13443_13742 , \13444_13743 , \13445_13744 , \13446_13745 ,
         \13447_13746 , \13448_13747 , \13449_13748 , \13450_13749 , \13451_13750 , \13452_13751 , \13453_13752 , \13454_13753 , \13455_13754 , \13456_13755 ,
         \13457_13756 , \13458_13757 , \13459_13758 , \13460_13759 , \13461_13760 , \13462_13761 , \13463_13762 , \13464_13763 , \13465_13764 , \13466_13765 ,
         \13467_13766 , \13468_13767 , \13469_13768 , \13470_13769 , \13471_13770 , \13472_13771 , \13473_13772 , \13474_13773 , \13475_13774 , \13476_13775 ,
         \13477_13776 , \13478_13777 , \13479_13778 , \13480_13779 , \13481_13780 , \13482_13781 , \13483_13782 , \13484_13783 , \13485_13784 , \13486_13785 ,
         \13487_13786 , \13488_13787 , \13489_13788 , \13490_13789 , \13491_13790 , \13492_13791 , \13493_13792 , \13494_13793 , \13495_13794 , \13496_13795 ,
         \13497_13796 , \13498_13797 , \13499_13798 , \13500_13799 , \13501_13800 , \13502_13801 , \13503_13802 , \13504_13803 , \13505_13804 , \13506_13805 ,
         \13507_13806 , \13508_13807 , \13509_13808 , \13510_13809 , \13511_13810 , \13512_13811 , \13513_13812 , \13514_13813 , \13515_13814 , \13516_13815 ,
         \13517_13816 , \13518_13817 , \13519_13818 , \13520_13819 , \13521_13820 , \13522_13821 , \13523_13822 , \13524_13823 , \13525_13824 , \13526_13825 ,
         \13527_13826 , \13528_13827 , \13529_13828 , \13530_13829 , \13531_13830 , \13532_13831 , \13533_13832 , \13534_13833 , \13535_13834 , \13536_13835 ,
         \13537_13836 , \13538_13837 , \13539_13838 , \13540_13839 , \13541_13840 , \13542_13841 , \13543_13842 , \13544_13843 , \13545_13844 , \13546_13845 ,
         \13547_13846 , \13548_13847 , \13549_13848 , \13550_13849 , \13551_13850 , \13552_13851 , \13553_13852 , \13554_13853 , \13555_13854 , \13556_13855 ,
         \13557_13856 , \13558_13857 , \13559_13858 , \13560_13859 , \13561_13860 , \13562_13861 , \13563_13862 , \13564_13863 , \13565_13864 , \13566_13865 ,
         \13567_13866 , \13568_13867 , \13569_13868 , \13570_13869 , \13571_13870 , \13572_13871 , \13573_13872 , \13574_13873 , \13575_13874 , \13576_13875 ,
         \13577_13876 , \13578_13877 , \13579_13878 , \13580_13879 , \13581_13880 , \13582_13881 , \13583_13882 , \13584_13883 , \13585_13884 , \13586_13885 ,
         \13587_13886 , \13588_13887 , \13589_13888 , \13590_13889 , \13591 , \13592_13891 , \13593_13892 , \13594_13893 , \13595_13894 , \13596_13895 ,
         \13597_13896 , \13598_13897 , \13599_13898 , \13600_13899 , \13601_13900 , \13602_13901 , \13603_13902 , \13604_13903 , \13605_13904 , \13606_13905 ,
         \13607_13906 , \13608_13907 , \13609_13908 , \13610_13909 , \13611_13910 , \13612_13911 , \13613_13912 , \13614_13913 , \13615_13914 , \13616_13915 ,
         \13617_13916 , \13618_13917 , \13619_13918 , \13620_13919 , \13621_13920 , \13622_13921 , \13623_13922 , \13624_13923 , \13625_13924 , \13626_13925 ,
         \13627_13926 , \13628_13927 , \13629_13928 , \13630_13929 , \13631_13930 , \13632_13931 , \13633_13932 , \13634_13933 , \13635_13934 , \13636_13935 ,
         \13637_13936 , \13638_13937 , \13639_13938 , \13640_13939 , \13641_13940 , \13642_13941 , \13643_13942 , \13644_13943 , \13645_13944 , \13646_13945 ,
         \13647_13946 , \13648_13947 , \13649_13948 , \13650_13949 , \13651_13950 , \13652_13951 , \13653_13952 , \13654_13953 , \13655_13954 , \13656_13955 ,
         \13657_13956 , \13658_13957 , \13659_13958 , \13660_13959 , \13661_13960 , \13662_13961 , \13663_13962 , \13664_13963 , \13665_13964 , \13666_13965 ,
         \13667_13966 , \13668_13967 , \13669_13968 , \13670_13969 , \13671_13970 , \13672_13971 , \13673_13972 , \13674_13973 , \13675_13974 , \13676_13975 ,
         \13677_13976 , \13678_13977 , \13679_13978 , \13680_13979 , \13681_13980 , \13682_13981 , \13683_13982 , \13684_13983 , \13685_13984 , \13686_13985 ,
         \13687_13986 , \13688_13987 , \13689_13988 , \13690_13989 , \13691_13990 , \13692_13991 , \13693_13992 , \13694_13993 , \13695_13994 , \13696_13995 ,
         \13697_13996 , \13698_13997 , \13699_13998 , \13700_13999 , \13701_14000 , \13702_14001 , \13703_14002 , \13704_14003 , \13705_14004 , \13706_14005 ,
         \13707_14006 , \13708_14007 , \13709_14008 , \13710_14009 , \13711_14010 , \13712_14011 , \13713_14012 , \13714_14013 , \13715_14014 , \13716_14015 ,
         \13717_14016 , \13718_14017 , \13719_14018 , \13720_14019 , \13721_14020 , \13722_14021 , \13723 , \13724_14023_nG658e , \13725_14024 , \13726_14025 ,
         \13727_14026 , \13728_14027 , \13729_14028 , \13730 , \13731 , \13732_14031_nG4c9e , \13733_14032 , \13734_14033 , \13735_14034 , \13736_14035 ,
         \13737_14036 , \13738_14037 , \13739_14038 , \13740_14039 , \13741_14040 , \13742_14041 , \13743_14042 , \13744_14043 , \13745_14044 , \13746_14045 ,
         \13747_14046 , \13748_14047 , \13749_14048 , \13750_14049 , \13751_14050 , \13752_14051 , \13753_14052 , \13754_14053 , \13755_14054 , \13756_14055 ,
         \13757_14056 , \13758_14057 , \13759_14058 , \13760_14059 , \13761_14060 , \13762_14061 , \13763_14062 , \13764_14063 , \13765_14064 , \13766_14065 ,
         \13767_14066 , \13768_14067 , \13769_14068 , \13770_14069 , \13771_14070_nG9bf9 , \13772_14071 , \13773_14072 , \13774_14073 , \13775_14074 , \13776_14075 ,
         \13777_14076 , \13778_14077 , \13779_14078 , \13780_14079 , \13781_14080 , \13782_14081 , \13783_14082 , \13784_14083 , \13785_14084 , \13786_14085 ,
         \13787_14086 , \13788_14087 , \13789_14088 , \13790_14089 , \13791_14090 , \13792_14091 , \13793_14092 , \13794_14093 , \13795_14094 , \13796_14095 ,
         \13797_14096 , \13798_14097 , \13799_14098 , \13800_14099 , \13801_14100 , \13802_14101 , \13803_14102 , \13804_14103 , \13805_14104 , \13806_14105 ,
         \13807_14106 , \13808_14107 , \13809_14108 , \13810_14109 , \13811_14110 , \13812_14111 , \13813_14112 , \13814_14113 , \13815_14114 , \13816_14115 ,
         \13817_14116 , \13818_14117 , \13819_14118 , \13820_14119 , \13821_14120 , \13822_14121 , \13823_14122 , \13824_14123 , \13825_14124 , \13826_14125 ,
         \13827_14126 , \13828_14127 , \13829_14128 , \13830_14129 , \13831_14130 , \13832_14131 , \13833_14132 , \13834_14133 , \13835_14134 , \13836_14135 ,
         \13837_14136 , \13838_14137 , \13839_14138 , \13840_14139 , \13841_14140 , \13842_14141 , \13843_14142 , \13844_14143 , \13845_14144 , \13846_14145 ,
         \13847_14146 , \13848_14147 , \13849_14148 , \13850_14149 , \13851_14150 , \13852_14151 , \13853_14152 , \13854_14153 , \13855_14154 , \13856_14155 ,
         \13857_14156 , \13858_14157 , \13859_14158 , \13860_14159 , \13861_14160 , \13862_14161 , \13863_14162 , \13864_14163 , \13865_14164 , \13866_14165 ,
         \13867_14166 , \13868_14167 , \13869_14168 , \13870_14169 , \13871_14170 , \13872_14171 , \13873_14172 , \13874_14173 , \13875_14174 , \13876_14175 ,
         \13877_14176 , \13878_14177 , \13879_14178 , \13880_14179 , \13881_14180 , \13882_14181 , \13883_14182 , \13884_14183 , \13885_14184 , \13886_14185 ,
         \13887_14186 , \13888_14187 , \13889_14188 , \13890_14189 , \13891_14190 , \13892_14191 , \13893_14192 , \13894_14193 , \13895_14194 , \13896_14195 ,
         \13897_14196 , \13898_14197 , \13899_14198 , \13900_14199 , \13901_14200 , \13902_14201 , \13903_14202 , \13904_14203 , \13905_14204 , \13906_14205 ,
         \13907_14206 , \13908_14207 , \13909_14208 , \13910_14209 , \13911_14210 , \13912 , \13913_14212 , \13914_14213 , \13915_14214 , \13916_14215 ,
         \13917_14216 , \13918_14217 , \13919_14218 , \13920_14219 , \13921_14220 , \13922_14221 , \13923_14222 , \13924_14223 , \13925_14224 , \13926_14225 ,
         \13927_14226 , \13928_14227 , \13929_14228 , \13930_14229 , \13931_14230 , \13932_14231 , \13933_14232 , \13934_14233 , \13935_14234 , \13936_14235 ,
         \13937_14236 , \13938_14237 , \13939_14238 , \13940_14239 , \13941_14240 , \13942_14241 , \13943_14242 , \13944_14243 , \13945_14244 , \13946_14245 ,
         \13947_14246 , \13948_14247 , \13949_14248 , \13950_14249 , \13951_14250 , \13952_14251 , \13953_14252 , \13954_14253 , \13955_14254 , \13956_14255 ,
         \13957_14256 , \13958_14257 , \13959_14258 , \13960_14259 , \13961_14260 , \13962_14261 , \13963_14262 , \13964_14263 , \13965_14264 , \13966_14265 ,
         \13967_14266 , \13968_14267 , \13969_14268 , \13970_14269 , \13971_14270 , \13972_14271 , \13973_14272 , \13974_14273 , \13975_14274 , \13976_14275 ,
         \13977_14276 , \13978_14277 , \13979_14278 , \13980_14279 , \13981_14280 , \13982_14281 , \13983_14282 , \13984_14283 , \13985_14284 , \13986_14285 ,
         \13987_14286 , \13988_14287 , \13989_14288 , \13990_14289 , \13991_14290 , \13992_14291 , \13993_14292 , \13994_14293 , \13995_14294 , \13996_14295 ,
         \13997_14296 , \13998_14297 , \13999_14298 , \14000_14299 , \14001_14300 , \14002_14301 , \14003_14302 , \14004_14303 , \14005_14304 , \14006_14305 ,
         \14007_14306 , \14008_14307 , \14009_14308 , \14010_14309 , \14011_14310 , \14012_14311 , \14013_14312 , \14014_14313 , \14015_14314 , \14016_14315 ,
         \14017_14316 , \14018_14317 , \14019_14318 , \14020_14319 , \14021_14320 , \14022_14321 , \14023_14322 , \14024_14323 , \14025_14324 , \14026_14325 ,
         \14027_14326 , \14028_14327 , \14029_14328 , \14030_14329 , \14031_14330 , \14032_14331 , \14033_14332 , \14034_14333 , \14035_14334 , \14036_14335 ,
         \14037_14336 , \14038_14337 , \14039_14338 , \14040_14339 , \14041_14340 , \14042_14341 , \14043_14342 , \14044_14343 , \14045 , \14046_14345 ,
         \14047_14346 , \14048_14347 , \14049_14348 , \14050_14349 , \14051_14350 , \14052_14351 , \14053_14352 , \14054_14353 , \14055_14354 , \14056_14355 ,
         \14057_14356 , \14058_14357 , \14059_14358 , \14060_14359 , \14061_14360 , \14062_14361 , \14063_14362 , \14064_14363 , \14065_14364 , \14066_14365 ,
         \14067_14366 , \14068_14367 , \14069_14368 , \14070_14369 , \14071_14370 , \14072_14371 , \14073_14372 , \14074_14373 , \14075_14374 , \14076_14375 ,
         \14077_14376 , \14078_14377 , \14079_14378 , \14080_14379 , \14081_14380 , \14082_14381 , \14083_14382 , \14084_14383 , \14085_14384 , \14086_14385 ,
         \14087_14386 , \14088_14387 , \14089_14388 , \14090_14389 , \14091_14390 , \14092_14391 , \14093_14392 , \14094_14393 , \14095_14394 , \14096_14395 ,
         \14097_14396 , \14098_14397 , \14099_14398 , \14100_14399 , \14101_14400 , \14102_14401 , \14103_14402 , \14104_14403 , \14105_14404 , \14106_14405 ,
         \14107_14406 , \14108_14407 , \14109_14408 , \14110_14409 , \14111_14410 , \14112_14411 , \14113_14412 , \14114_14413 , \14115_14414 , \14116_14415 ,
         \14117_14416 , \14118_14417 , \14119_14418 , \14120_14419 , \14121_14420 , \14122_14421 , \14123_14422 , \14124_14423 , \14125_14424 , \14126_14425 ,
         \14127_14426 , \14128_14427 , \14129_14428 , \14130_14429 , \14131_14430 , \14132_14431 , \14133_14432 , \14134_14433 , \14135_14434 , \14136_14435 ,
         \14137_14436 , \14138_14437 , \14139_14438 , \14140_14439 , \14141_14440 , \14142_14441 , \14143_14442 , \14144_14443 , \14145_14444 , \14146_14445 ,
         \14147_14446 , \14148_14447 , \14149_14448 , \14150_14449 , \14151_14450 , \14152_14451 , \14153_14452 , \14154_14453 , \14155_14454 , \14156_14455 ,
         \14157_14456 , \14158_14457 , \14159_14458 , \14160_14459 , \14161_14460 , \14162_14461 , \14163_14462 , \14164_14463 , \14165_14464 , \14166_14465 ,
         \14167_14466 , \14168_14467 , \14169_14468 , \14170_14469 , \14171_14470 , \14172_14471 , \14173_14472 , \14174_14473 , \14175_14474 , \14176_14475 ,
         \14177_14476 , \14178_14477 , \14179 , \14180_14479 , \14181_14480 , \14182_14481 , \14183_14482 , \14184_14483 , \14185_14484 , \14186_14485 ,
         \14187_14486 , \14188_14487 , \14189_14488 , \14190_14489 , \14191_14490 , \14192_14491 , \14193_14492 , \14194_14493 , \14195_14494 , \14196_14495 ,
         \14197_14496 , \14198_14497 , \14199_14498 , \14200_14499 , \14201_14500 , \14202_14501 , \14203_14502 , \14204_14503 , \14205_14504 , \14206_14505 ,
         \14207_14506 , \14208_14507 , \14209_14508 , \14210_14509 , \14211_14510 , \14212_14511 , \14213_14512 , \14214_14513 , \14215_14514 , \14216_14515 ,
         \14217_14516 , \14218_14517 , \14219_14518 , \14220_14519 , \14221_14520 , \14222_14521 , \14223_14522 , \14224_14523 , \14225_14524 , \14226_14525 ,
         \14227_14526 , \14228_14527 , \14229_14528 , \14230_14529 , \14231_14530 , \14232_14531 , \14233_14532 , \14234_14533 , \14235_14534 , \14236_14535 ,
         \14237_14536 , \14238_14537 , \14239_14538 , \14240_14539 , \14241_14540 , \14242_14541 , \14243_14542 , \14244_14543 , \14245_14544 , \14246_14545 ,
         \14247_14546 , \14248_14547 , \14249_14548 , \14250_14549 , \14251_14550 , \14252_14551 , \14253_14552 , \14254_14553 , \14255_14554 , \14256_14555 ,
         \14257_14556 , \14258_14557 , \14259_14558 , \14260_14559 , \14261_14560 , \14262_14561 , \14263_14562 , \14264_14563 , \14265_14564 , \14266_14565 ,
         \14267_14566 , \14268_14567 , \14269_14568 , \14270_14569 , \14271_14570 , \14272_14571 , \14273_14572 , \14274_14573 , \14275_14574 , \14276_14575 ,
         \14277_14576 , \14278_14577 , \14279_14578 , \14280_14579 , \14281_14580 , \14282_14581 , \14283_14582 , \14284_14583 , \14285_14584 , \14286_14585 ,
         \14287_14586 , \14288_14587 , \14289_14588 , \14290_14589 , \14291_14590 , \14292_14591 , \14293_14592 , \14294_14593 , \14295_14594 , \14296_14595 ,
         \14297_14596 , \14298_14597 , \14299_14598 , \14300_14599 , \14301_14600 , \14302_14601 , \14303_14602 , \14304_14603 , \14305_14604 , \14306_14605 ,
         \14307_14606 , \14308_14607 , \14309_14608 , \14310_14609 , \14311_14610 , \14312 , \14313_14612 , \14314_14613 , \14315_14614 , \14316_14615 ,
         \14317_14616 , \14318_14617 , \14319_14618 , \14320_14619 , \14321_14620 , \14322_14621 , \14323_14622_nG443c , \14324_14623 , \14325_14624 , \14326_14625_nG443f ,
         \14327_14626 , \14328_14627 , \14329_14628 , \14330_14632 , \14331_14633 , \14332_14634 , \14333_14635 , \14334_14636 , \14335_14637 , \14336_14638 ,
         \14337_14639 , \14338_14640 , \14339_14641 , \14340_14642 , \14341_14643 , \14342_14644 , \14343_14645 , \14344_14646 , \14345_14647 , \14346_14648 ,
         \14347_14649 , \14348_14650 , \14349_14651 , \14350_14652 , \14351_14653 , \14352_14654 , \14353_14655 , \14354_14656 , \14355_14657 , \14356_14658 ,
         \14357_14659 , \14358_14660 , \14359_14661 , \14360_14662 , \14361_14663 , \14362_14664 , \14363_14665 , \14364_14666 , \14365_14667 , \14366_14668 ,
         \14367_14669 , \14368_14670 , \14369_14671 , \14370_14672 , \14371_14673 , \14372_14674 , \14373_14675 , \14374_14676 , \14375_14677 , \14376_14678 ,
         \14377_14679 , \14378_14680 , \14379_14681 , \14380_14682 , \14381_14683 , \14382_14684 , \14383_14685 , \14384_14686 , \14385_14687 , \14386_14688 ,
         \14387_14689 , \14388_14690 , \14389_14691 , \14390_14692 , \14391_14693 , \14392_14694 , \14393_14695 , \14394_14696 , \14395_14697 , \14396_14698 ,
         \14397_14699 , \14398_14700 , \14399_14701 , \14400_14702 , \14401_14703 , \14402_14704 , \14403_14705 , \14404_14706 , \14405_14707 , \14406_14708 ,
         \14407_14709 , \14408_14710 , \14409_14711 , \14410_14712 , \14411_14713 , \14412_14714 , \14413_14715 , \14414_14716 , \14415_14717 , \14416_14718 ,
         \14417_14719 , \14418_14720 , \14419_14721 , \14420_14722 , \14421_14723 , \14422_14724 , \14423_14725 , \14424_14726 , \14425_14727 , \14426_14728 ,
         \14427_14729 , \14428_14730 , \14429_14731 , \14430_14732 , \14431_14733 , \14432_14734 , \14433_14735 , \14434_14736 , \14435_14737 , \14436_14738 ,
         \14437_14739 , \14438_14740 , \14439_14741 , \14440_14742 , \14441_14743 , \14442_14744 , \14443_14745 , \14444_14746 , \14445_14747 , \14446_14748 ,
         \14447_14749 , \14448_14750 , \14449_14751 , \14450_14752 , \14451_14753 , \14452_14754 , \14453_14755 , \14454_14756 , \14455_14757 , \14456_14758 ,
         \14457_14759 , \14458_14760 , \14459_14761 , \14460_14762 , \14461_14763 , \14462_14764 , \14463_14765 , \14464_14766 , \14465_14767 , \14466_14768 ,
         \14467_14769 , \14468_14770 , \14469_14771 , \14470_14772 , \14471_14773 , \14472_14774 , \14473_14775 , \14474_14776 , \14475_14777 , \14476_14778 ,
         \14477_14779 , \14478_14780 , \14479_14781 , \14480_14782 , \14481_14783 , \14482_14784 , \14483_14785 , \14484_14786 , \14485_14787 , \14486_14788 ,
         \14487_14789 , \14488_14790 , \14489_14791 , \14490_14792 , \14491_14793 , \14492_14794 , \14493_14795 , \14494_14796 , \14495_14797 , \14496_14798 ,
         \14497_14799 , \14498_14800 , \14499_14801 , \14500_14802 , \14501_14803 , \14502_14804 , \14503_14805 , \14504_14806 , \14505_14807 , \14506_14808 ,
         \14507_14809 , \14508_14810 , \14509_14811 , \14510_14812 , \14511_14813 , \14512_14814 , \14513_14815 , \14514 , \14515_14817 , \14516_14818 ,
         \14517_14819 , \14518_14820 , \14519_14821 , \14520_14822 , \14521_14823 , \14522_14824 , \14523_14825 , \14524_14826 , \14525_14827 , \14526_14828 ,
         \14527_14829 , \14528_14830 , \14529_14831 , \14530_14832 , \14531_14833 , \14532_14834 , \14533_14835 , \14534_14836 , \14535_14837 , \14536_14838 ,
         \14537_14839 , \14538_14840 , \14539_14841 , \14540_14842 , \14541_14843 , \14542_14844 , \14543_14845 , \14544_14846 , \14545_14847 , \14546_14848 ,
         \14547_14849 , \14548_14850 , \14549_14851 , \14550_14852 , \14551_14853 , \14552_14854 , \14553_14855 , \14554_14856 , \14555_14857 , \14556_14858 ,
         \14557_14859 , \14558_14860 , \14559_14861 , \14560_14862 , \14561_14863 , \14562_14864 , \14563_14865 , \14564_14866 , \14565_14867 , \14566_14868 ,
         \14567_14869 , \14568_14870 , \14569_14871 , \14570_14872 , \14571_14873 , \14572_14874 , \14573_14875 , \14574_14876 , \14575_14877 , \14576_14878 ,
         \14577_14879 , \14578_14880 , \14579_14881 , \14580_14882 , \14581_14883 , \14582_14884 , \14583_14885 , \14584_14886 , \14585_14887 , \14586_14888 ,
         \14587_14889 , \14588_14890 , \14589_14891 , \14590_14892 , \14591_14893 , \14592_14894 , \14593_14895 , \14594_14896 , \14595_14897 , \14596_14898 ,
         \14597_14899 , \14598_14900 , \14599_14901 , \14600_14902 , \14601_14903 , \14602_14904 , \14603_14905 , \14604_14906 , \14605_14907 , \14606_14908 ,
         \14607_14909 , \14608_14910 , \14609_14911 , \14610_14912 , \14611_14913 , \14612_14914 , \14613_14915 , \14614_14916 , \14615_14917 , \14616_14918 ,
         \14617_14919 , \14618_14920 , \14619_14921 , \14620_14922 , \14621_14923 , \14622_14924 , \14623_14925 , \14624_14926 , \14625_14927 , \14626_14928 ,
         \14627_14929 , \14628_14930 , \14629_14931 , \14630_14932 , \14631_14933 , \14632_14934 , \14633_14935 , \14634_14936 , \14635_14937 , \14636_14938 ,
         \14637_14939 , \14638_14940 , \14639_14941 , \14640_14942 , \14641_14943 , \14642_14944 , \14643_14945 , \14644_14946 , \14645_14947 , \14646 ,
         \14647_14949_nG6591 , \14648_14950 , \14649_14951 , \14650_14952 , \14651_14953 , \14652_14954 , \14653_14955 , \14654_14956 , \14655_14957 , \14656_14958 ,
         \14657 , \14658 , \14659_14961_nG4da7 , \14660_14962 , \14661_14963 , \14662_14964 , \14663_14965 , \14664_14966 , \14665_14967 , \14666_14968 ,
         \14667_14969 , \14668_14970 , \14669_14971 , \14670_14972 , \14671_14973 , \14672_14974 , \14673_14975 , \14674_14976 , \14675_14977 , \14676_14978 ,
         \14677_14979 , \14678_14980 , \14679_14981 , \14680_14982 , \14681_14983 , \14682_14984_nG9bf6 , \14683_14985 , \14684_14986 , \14685_14987 , \14686_14988 ,
         \14687_14989 , \14688_14990 , \14689_14991 , \14690_14992 , \14691_14993 , \14692_14994 , \14693_14995 , \14694_14996 , \14695_14997 , \14696_14998 ,
         \14697_14999 , \14698_15000 , \14699_15001 , \14700_15002 , \14701_15003 , \14702_15004 , \14703_15005 , \14704_15006 , \14705_15007 , \14706_15008 ,
         \14707_15009 , \14708_14629 , \14709_14630 , \14710_14631 , \14711_15010 , \14712_15011 , \14713_15012 , \14714_15013 , \14715_15014 , \14716_15015 ,
         \14717_15016 , \14718_15017 , \14719_15018 , \14720_15019 , \14721_15020 , \14722_15021 , \14723_15022 , \14724_15023 , \14725_15024 , \14726_15025 ,
         \14727_15026 , \14728_15027 , \14729_15028 , \14730_15029 , \14731_15030 , \14732_15031 , \14733_15032 , \14734_15033 , \14735_15034 , \14736_15035 ,
         \14737_15036 , \14738_15037 , \14739_15038 , \14740_15039 , \14741_15040 , \14742_15041 , \14743_15042 , \14744_15043 , \14745_15044 , \14746_15045 ,
         \14747_15046 , \14748_15047 , \14749_15048 , \14750_15049 , \14751_15050 , \14752_15051 , \14753_15052 , \14754_15053 , \14755_15054 , \14756_15055 ,
         \14757_15056 , \14758_15057 , \14759_15058 , \14760_15059 , \14761_15060 , \14762_15061 , \14763_15062 , \14764_15063 , \14765_15064 , \14766_15065 ,
         \14767_15066 , \14768_15067 , \14769_15068 , \14770_15069 , \14771_15070 , \14772_15071 , \14773_15072 , \14774_15073 , \14775_15074 , \14776_15075 ,
         \14777_15076 , \14778_15077 , \14779_15078 , \14780_15079 , \14781_15080 , \14782_15081 , \14783_15082 , \14784_15083 , \14785_15084 , \14786_15085 ,
         \14787_15086 , \14788_15087 , \14789_15088 , \14790_15089 , \14791_15090 , \14792_15091 , \14793_15092 , \14794_15093 , \14795_15094 , \14796_15095 ,
         \14797_15096 , \14798_15097 , \14799_15098 , \14800_15099 , \14801_15100 , \14802_15101 , \14803_15102 , \14804_15103 , \14805_15104 , \14806_15105 ,
         \14807_15106 , \14808_15107 , \14809_15108 , \14810_15109 , \14811_15110 , \14812_15111 , \14813_15112 , \14814_15113 , \14815_15114 , \14816_15115 ,
         \14817_15116 , \14818_15117 , \14819_15118 , \14820_15119 , \14821_15120 , \14822_15121 , \14823_15122 , \14824_15123 , \14825_15124 , \14826_15125 ,
         \14827_15126 , \14828_15127 , \14829_15128 , \14830_15129 , \14831_15130 , \14832_15131 , \14833_15132 , \14834_15133 , \14835_15134 , \14836_15135 ,
         \14837_15136 , \14838_15137 , \14839_15138 , \14840_15139 , \14841_15140 , \14842_15141 , \14843_15142 , \14844_15143 , \14845_15144 , \14846_15145 ,
         \14847_15146 , \14848_15147 , \14849_15148 , \14850_15149 , \14851_15150 , \14852_15151 , \14853_15152 , \14854_15153 , \14855_15154 , \14856_15155 ,
         \14857_15156 , \14858_15157 , \14859_15158 , \14860_15159 , \14861_15160 , \14862_15161 , \14863_15162 , \14864_15163 , \14865_15164 , \14866_15165 ,
         \14867_15166 , \14868_15167 , \14869_15168 , \14870_15169 , \14871_15170 , \14872_15171 , \14873_15172 , \14874_15173 , \14875_15174 , \14876_15175 ,
         \14877_15176 , \14878_15177 , \14879_15178 , \14880_15179 , \14881_15180 , \14882_15181 , \14883_15182 , \14884_15183 , \14885_15184 , \14886_15185 ,
         \14887_15186 , \14888 , \14889_15188 , \14890_15189 , \14891_15190 , \14892_15191 , \14893_15192 , \14894_15193 , \14895_15194 , \14896_15195 ,
         \14897_15196 , \14898_15197 , \14899_15198 , \14900_15199 , \14901_15200 , \14902_15201 , \14903_15202 , \14904_15203 , \14905_15204 , \14906_15205 ,
         \14907_15206 , \14908_15207 , \14909_15208 , \14910_15209 , \14911_15210 , \14912_15211 , \14913_15212 , \14914_15213 , \14915_15214 , \14916_15215 ,
         \14917_15216 , \14918_15217 , \14919_15218 , \14920_15219 , \14921_15220 , \14922_15221 , \14923_15222 , \14924_15223 , \14925_15224 , \14926_15225 ,
         \14927_15226 , \14928_15227 , \14929_15228 , \14930_15229 , \14931_15230 , \14932_15231 , \14933_15232 , \14934_15233 , \14935_15234 , \14936_15235 ,
         \14937_15236 , \14938_15237 , \14939_15238 , \14940_15239 , \14941_15240 , \14942_15241 , \14943_15242 , \14944_15243 , \14945_15244 , \14946_15245 ,
         \14947_15246 , \14948_15247 , \14949_15248 , \14950_15249 , \14951_15250 , \14952_15251 , \14953_15252 , \14954_15253 , \14955_15254 , \14956_15255 ,
         \14957_15256 , \14958_15257 , \14959_15258 , \14960_15259 , \14961_15260 , \14962_15261 , \14963_15262 , \14964_15263 , \14965_15264 , \14966_15265 ,
         \14967_15266 , \14968_15267 , \14969_15268 , \14970_15269 , \14971_15270 , \14972_15271 , \14973_15272 , \14974_15273 , \14975_15274 , \14976_15275 ,
         \14977_15276 , \14978_15277 , \14979_15278 , \14980_15279 , \14981_15280 , \14982_15281 , \14983_15282 , \14984_15283 , \14985_15284 , \14986_15285 ,
         \14987_15286 , \14988_15287 , \14989_15288 , \14990_15289 , \14991_15290 , \14992_15291 , \14993_15292 , \14994_15293 , \14995_15294 , \14996_15295 ,
         \14997_15296 , \14998_15297 , \14999_15298 , \15000_15299 , \15001_15300 , \15002_15301 , \15003_15302 , \15004_15303 , \15005_15304 , \15006_15305 ,
         \15007_15306 , \15008_15307 , \15009_15308 , \15010_15309 , \15011_15310 , \15012_15311 , \15013_15312 , \15014_15313 , \15015_15314 , \15016_15315 ,
         \15017_15316 , \15018_15317 , \15019_15318 , \15020 , \15021_15320_nG6594 , \15022_15321 , \15023_15322 , \15024_15323 , \15025_15324 , \15026_15325 ,
         \15027_15326 , \15028_15327 , \15029_15328 , \15030_15329 , \15031 , \15032 , \15033_15332_nG4eb0 , \15034_15333 , \15035_15334 , \15036_15335 ,
         \15037_15336 , \15038_15337 , \15039_15338 , \15040_15339 , \15041_15340 , \15042_15341 , \15043_15342 , \15044_15343 , \15045_15344 , \15046_15345 ,
         \15047_15346 , \15048_15347 , \15049_15348 , \15050_15349 , \15051_15350 , \15052_15351 , \15053_15352 , \15054_15353 , \15055_15354 , \15056_15355 ,
         \15057_15356 , \15058_15357 , \15059_15358 , \15060_15359 , \15061_15360 , \15062_15361 , \15063_15362 , \15064_15363 , \15065_15364 , \15066_15365 ,
         \15067_15366 , \15068_15367 , \15069_15368 , \15070_15369 , \15071_15370 , \15072_15371 , \15073_15372 , \15074_15373_nG9bf3 , \15075_15374 , \15076_15375 ,
         \15077_15376 , \15078_15377 , \15079_15378 , \15080_15379 , \15081_15380 , \15082_15381 , \15083_15382 , \15084_15383 , \15085_15384 , \15086_15385 ,
         \15087_15386 , \15088_15387 , \15089_15388 , \15090_15389 , \15091_15390 , \15092_15391 , \15093_15392 , \15094_15393 , \15095_15394 , \15096_15395 ,
         \15097_15396 , \15098_15397 , \15099_15398 , \15100_15399 , \15101_15400 , \15102_15401 , \15103_15402 , \15104_15403 , \15105_15404 , \15106_15405 ,
         \15107_15406 , \15108_15407 , \15109_15408 , \15110_15409 , \15111_15410 , \15112_15411 , \15113_15412 , \15114_15413 , \15115_15414 , \15116_15415 ,
         \15117_15416 , \15118_15417 , \15119_15418 , \15120_15419 , \15121_15420 , \15122_15421 , \15123_15422 , \15124_15423 , \15125_15424 , \15126_15425 ,
         \15127_15426 , \15128_15427 , \15129_15428 , \15130_15429 , \15131_15430 , \15132_15431 , \15133_15432 , \15134_15433 , \15135_15434 , \15136_15435 ,
         \15137_15436 , \15138_15437 , \15139_15438 , \15140_15439 , \15141_15440 , \15142_15441 , \15143_15442 , \15144_15443 , \15145_15444 , \15146_15445 ,
         \15147_15446 , \15148_15447 , \15149_15448 , \15150_15449 , \15151_15450 , \15152_15451 , \15153_15452 , \15154_15453 , \15155_15454 , \15156_15455 ,
         \15157_15456 , \15158_15457 , \15159_15458 , \15160_15459 , \15161_15460 , \15162_15461 , \15163_15462 , \15164_15463 , \15165_15464 , \15166_15465 ,
         \15167_15466 , \15168_15467 , \15169_15468 , \15170_15469 , \15171_15470 , \15172_15471 , \15173_15472 , \15174_15473 , \15175_15474 , \15176_15475 ,
         \15177_15476 , \15178_15477 , \15179_15478 , \15180_15479 , \15181_15480 , \15182_15481 , \15183_15482 , \15184_15483 , \15185_15484 , \15186_15485 ,
         \15187_15486 , \15188_15487 , \15189_15488 , \15190_15489 , \15191_15490 , \15192_15491 , \15193_15492 , \15194_15493 , \15195_15494 , \15196_15495 ,
         \15197_15496 , \15198_15497 , \15199_15498 , \15200_15499 , \15201_15500 , \15202_15501 , \15203_15502 , \15204_15503 , \15205_15504 , \15206_15505 ,
         \15207_15506 , \15208_15507 , \15209_15508 , \15210_15509 , \15211_15510 , \15212_15511 , \15213_15512 , \15214_15513 , \15215_15514 , \15216_15515 ,
         \15217_15516 , \15218_15517 , \15219_15518 , \15220_15519 , \15221 , \15222_15521 , \15223_15522 , \15224_15523 , \15225_15524 , \15226_15525 ,
         \15227_15526 , \15228_15527 , \15229_15528 , \15230_15529 , \15231_15530 , \15232_15531 , \15233_15532 , \15234_15533 , \15235_15534 , \15236_15535 ,
         \15237_15536 , \15238_15537 , \15239_15538 , \15240_15539 , \15241_15540 , \15242_15541 , \15243_15542 , \15244_15543 , \15245_15544 , \15246_15545 ,
         \15247_15546 , \15248_15547 , \15249_15548 , \15250_15549 , \15251_15550 , \15252_15551 , \15253_15552 , \15254_15553 , \15255_15554 , \15256_15555 ,
         \15257_15556 , \15258_15557 , \15259_15558 , \15260_15559 , \15261_15560 , \15262_15561 , \15263_15562 , \15264_15563 , \15265_15564 , \15266_15565 ,
         \15267_15566 , \15268_15567 , \15269_15568 , \15270_15569 , \15271_15570 , \15272_15571 , \15273_15572 , \15274_15573 , \15275_15574 , \15276_15575 ,
         \15277_15576 , \15278_15577 , \15279_15578 , \15280_15579 , \15281_15580 , \15282_15581 , \15283_15582 , \15284_15583 , \15285_15584 , \15286_15585 ,
         \15287_15586 , \15288_15587 , \15289_15588 , \15290_15589 , \15291_15590 , \15292_15591 , \15293_15592 , \15294_15593 , \15295_15594 , \15296_15595 ,
         \15297_15596 , \15298_15597 , \15299_15598 , \15300_15599 , \15301_15600 , \15302_15601 , \15303_15602 , \15304_15603 , \15305_15604 , \15306_15605 ,
         \15307_15606 , \15308_15607 , \15309_15608 , \15310_15609 , \15311_15610 , \15312_15611 , \15313_15612 , \15314_15613 , \15315_15614 , \15316_15615 ,
         \15317_15616 , \15318_15617 , \15319_15618 , \15320_15619 , \15321_15620 , \15322_15621 , \15323_15622 , \15324_15623 , \15325_15624 , \15326_15625 ,
         \15327_15626 , \15328_15627 , \15329_15628 , \15330_15629 , \15331_15630 , \15332_15631 , \15333_15632 , \15334_15633 , \15335_15634 , \15336_15635 ,
         \15337_15636 , \15338_15637 , \15339_15638 , \15340_15639 , \15341_15640 , \15342_15641 , \15343_15642 , \15344_15643 , \15345_15644 , \15346_15645 ,
         \15347_15646 , \15348_15647 , \15349_15648 , \15350_15649 , \15351_15650 , \15352_15651 , \15353_15652 , \15354 , \15355_15654 , \15356_15655 ,
         \15357_15656 , \15358_15657 , \15359_15658 , \15360_15659 , \15361_15660 , \15362_15661 , \15363_15662 , \15364_15663 , \15365_15664 , \15366_15665 ,
         \15367_15666 , \15368_15667 , \15369_15668 , \15370_15669 , \15371_15670 , \15372_15671 , \15373_15672 , \15374_15673 , \15375_15674 , \15376_15675 ,
         \15377_15676 , \15378_15677 , \15379_15678 , \15380_15679 , \15381_15680 , \15382_15681 , \15383_15682 , \15384_15683 , \15385_15684 , \15386_15685 ,
         \15387_15686 , \15388_15687 , \15389_15688 , \15390_15689 , \15391_15690 , \15392_15691 , \15393_15692 , \15394_15693 , \15395_15694 , \15396_15695 ,
         \15397_15696 , \15398_15697 , \15399_15698 , \15400_15699 , \15401_15700 , \15402_15701 , \15403_15702 , \15404_15703 , \15405_15704 , \15406_15705 ,
         \15407_15706 , \15408_15707 , \15409_15708 , \15410_15709 , \15411_15710 , \15412_15711 , \15413_15712 , \15414_15713 , \15415_15714 , \15416_15715 ,
         \15417_15716 , \15418_15717 , \15419_15718 , \15420_15719 , \15421_15720 , \15422_15721 , \15423_15722 , \15424_15723 , \15425_15724 , \15426_15725 ,
         \15427_15726 , \15428_15727 , \15429_15728 , \15430_15729 , \15431_15730 , \15432_15731 , \15433_15732 , \15434_15733 , \15435_15734 , \15436_15735 ,
         \15437_15736 , \15438_15737 , \15439_15738 , \15440_15739 , \15441_15740 , \15442_15741 , \15443_15742 , \15444_15743 , \15445_15744 , \15446_15745 ,
         \15447_15746 , \15448_15747 , \15449_15748 , \15450_15749 , \15451_15750 , \15452_15751 , \15453_15752 , \15454_15753 , \15455_15754 , \15456_15755 ,
         \15457_15756 , \15458_15757 , \15459_15758 , \15460_15759 , \15461_15760 , \15462_15761 , \15463_15762 , \15464_15763 , \15465_15764 , \15466_15765 ,
         \15467_15766 , \15468_15767 , \15469_15768 , \15470_15769 , \15471_15770 , \15472_15771 , \15473_15772 , \15474_15773 , \15475_15774 , \15476_15775 ,
         \15477_15776 , \15478_15777 , \15479_15778 , \15480_15779 , \15481_15780 , \15482_15781 , \15483_15782 , \15484_15783 , \15485_15784 , \15486_15785 ,
         \15487_15786 , \15488 , \15489_15788 , \15490_15789 , \15491_15790 , \15492_15791 , \15493_15792 , \15494_15793 , \15495_15794 , \15496_15795 ,
         \15497_15796 , \15498_15797 , \15499_15798 , \15500_15799 , \15501_15800 , \15502_15801 , \15503_15802 , \15504_15803 , \15505_15804 , \15506_15805 ,
         \15507_15806 , \15508_15807 , \15509_15808 , \15510_15809 , \15511_15810 , \15512_15811 , \15513_15812 , \15514_15813 , \15515_15814 , \15516_15815 ,
         \15517_15816 , \15518_15817 , \15519_15818 , \15520_15819 , \15521_15820 , \15522_15821 , \15523_15822 , \15524_15823 , \15525_15824 , \15526_15825 ,
         \15527_15826 , \15528_15827 , \15529_15828 , \15530_15829 , \15531_15830 , \15532_15831 , \15533_15832 , \15534_15833 , \15535_15834 , \15536_15835 ,
         \15537_15836 , \15538_15837 , \15539_15838 , \15540_15839 , \15541_15840 , \15542_15841 , \15543_15842 , \15544_15843 , \15545_15844 , \15546_15845 ,
         \15547_15846 , \15548_15847 , \15549_15848 , \15550_15849 , \15551_15850 , \15552_15851 , \15553_15852 , \15554_15853 , \15555_15854 , \15556_15855 ,
         \15557_15856 , \15558_15857 , \15559_15858 , \15560_15859 , \15561_15860 , \15562_15861 , \15563_15862 , \15564_15863 , \15565_15864 , \15566_15865 ,
         \15567_15866 , \15568_15867 , \15569_15868 , \15570_15869 , \15571_15870 , \15572_15871 , \15573_15872 , \15574_15873 , \15575_15874 , \15576_15875 ,
         \15577_15876 , \15578_15877 , \15579_15878 , \15580_15879 , \15581_15880 , \15582_15881 , \15583_15882 , \15584_15883 , \15585_15884 , \15586_15885 ,
         \15587_15886 , \15588_15887 , \15589_15888 , \15590_15889 , \15591_15890 , \15592_15891 , \15593_15892 , \15594_15893 , \15595_15894 , \15596_15895 ,
         \15597_15896 , \15598_15897 , \15599_15898 , \15600_15899 , \15601_15900 , \15602_15901 , \15603_15902 , \15604_15903 , \15605_15904 , \15606_15905 ,
         \15607_15906 , \15608_15907 , \15609_15908 , \15610_15909 , \15611_15910 , \15612_15911 , \15613_15912 , \15614_15913 , \15615_15914 , \15616_15915 ,
         \15617_15916 , \15618_15917 , \15619_15918 , \15620_15919 , \15621 , \15622_15921 , \15623_15922 , \15624_15923 , \15625_15924 , \15626_15925 ,
         \15627_15926 , \15628_15927 , \15629_15928 , \15630_15929 , \15631_15930 , \15632_15931_nG4436 , \15633_15932 , \15634_15933 , \15635_15934_nG4439 , \15636_15935 ,
         \15637_15936 , \15638_15937 , \15639_15941 , \15640_15942 , \15641_15943 , \15642_15944 , \15643_15945 , \15644_15946 , \15645_15947 , \15646_15948 ,
         \15647_15949 , \15648_15950 , \15649_15951 , \15650_15952 , \15651_15953 , \15652_15954 , \15653_15955 , \15654_15956 , \15655_15957 , \15656_15958 ,
         \15657_15959 , \15658_15960 , \15659_15961 , \15660_15962 , \15661_15963 , \15662_15964 , \15663_15965 , \15664_15966 , \15665_15967 , \15666_15968 ,
         \15667_15969 , \15668_15970 , \15669_15971 , \15670_15972 , \15671_15973 , \15672_15974 , \15673_15975 , \15674_15976 , \15675_15977 , \15676_15978 ,
         \15677_15979 , \15678_15980 , \15679_15981 , \15680_15982 , \15681_15983 , \15682_15984 , \15683_15985 , \15684_15986 , \15685_15987 , \15686_15988 ,
         \15687_15989 , \15688_15990 , \15689_15991 , \15690_15992 , \15691_15993 , \15692_15994 , \15693_15995 , \15694_15996 , \15695_15997 , \15696_15998 ,
         \15697_15999 , \15698_16000 , \15699_16001 , \15700_16002 , \15701_16003 , \15702_16004 , \15703_16005 , \15704_16006 , \15705_16007 , \15706_16008 ,
         \15707_16009 , \15708_16010 , \15709_16011 , \15710_16012 , \15711_16013 , \15712_16014 , \15713_16015 , \15714_16016 , \15715_16017 , \15716_16018 ,
         \15717_16019 , \15718_16020 , \15719_16021 , \15720_16022 , \15721_16023 , \15722_16024 , \15723_16025 , \15724_16026 , \15725_16027 , \15726_16028 ,
         \15727_16029 , \15728_16030 , \15729_16031 , \15730_16032 , \15731_16033 , \15732_16034 , \15733_16035 , \15734_16036 , \15735_16037 , \15736_16038 ,
         \15737_16039 , \15738_16040 , \15739_16041 , \15740_16042 , \15741_16043 , \15742_16044 , \15743_16045 , \15744_16046 , \15745_16047 , \15746_16048 ,
         \15747_16049 , \15748_16050 , \15749_16051 , \15750_16052 , \15751_16053 , \15752_16054 , \15753_16055 , \15754_16056 , \15755_16057 , \15756_16058 ,
         \15757_16059 , \15758_16060 , \15759_16061 , \15760_16062 , \15761_16063 , \15762_16064 , \15763_16065 , \15764_16066 , \15765_16067 , \15766_16068 ,
         \15767_16069 , \15768_16070 , \15769_16071 , \15770_16072 , \15771_16073 , \15772_16074 , \15773_16075 , \15774_16076 , \15775_16077 , \15776_16078 ,
         \15777_16079 , \15778_16080 , \15779_16081 , \15780_16082 , \15781_16083 , \15782_16084 , \15783_16085 , \15784_16086 , \15785_16087 , \15786_16088 ,
         \15787_16089 , \15788_16090 , \15789_16091 , \15790_16092 , \15791_16093 , \15792_16094 , \15793_16095 , \15794_16096 , \15795_16097 , \15796_16098 ,
         \15797_16099 , \15798_16100 , \15799_16101 , \15800_16102 , \15801_16103 , \15802_16104 , \15803_16105 , \15804_16106 , \15805_16107 , \15806_16108 ,
         \15807_16109 , \15808_16110 , \15809_16111 , \15810_16112 , \15811_16113 , \15812_16114 , \15813_16115 , \15814_16116 , \15815_16117 , \15816_16118 ,
         \15817_16119 , \15818_16120 , \15819_16121 , \15820_16122 , \15821_16123 , \15822_16124 , \15823_16125 , \15824_16126 , \15825_16127 , \15826_16128 ,
         \15827_16129 , \15828_16130 , \15829_16131 , \15830_16132 , \15831 , \15832_16134 , \15833_16135 , \15834_16136 , \15835_16137 , \15836_16138 ,
         \15837_16139 , \15838_16140 , \15839_16141 , \15840_16142 , \15841_16143 , \15842_16144 , \15843_16145 , \15844_16146 , \15845_16147 , \15846_16148 ,
         \15847_16149 , \15848_16150 , \15849_16151 , \15850_16152 , \15851_16153 , \15852_16154 , \15853_16155 , \15854_16156 , \15855_16157 , \15856_16158 ,
         \15857_16159 , \15858_16160 , \15859_16161 , \15860_16162 , \15861_16163 , \15862_16164 , \15863_16165 , \15864_16166 , \15865_16167 , \15866_16168 ,
         \15867_16169 , \15868_16170 , \15869_16171 , \15870_16172 , \15871_16173 , \15872_16174 , \15873_16175 , \15874_16176 , \15875_16177 , \15876_16178 ,
         \15877_16179 , \15878_16180 , \15879_16181 , \15880_16182 , \15881_16183 , \15882_16184 , \15883_16185 , \15884_16186 , \15885_16187 , \15886_16188 ,
         \15887_16189 , \15888_16190 , \15889_16191 , \15890_16192 , \15891_16193 , \15892_16194 , \15893_16195 , \15894_16196 , \15895_16197 , \15896_16198 ,
         \15897_16199 , \15898_16200 , \15899_16201 , \15900_16202 , \15901_16203 , \15902_16204 , \15903_16205 , \15904_16206 , \15905_16207 , \15906_16208 ,
         \15907_16209 , \15908_16210 , \15909_16211 , \15910_16212 , \15911_16213 , \15912_16214 , \15913_16215 , \15914_16216 , \15915_16217 , \15916_16218 ,
         \15917_16219 , \15918_16220 , \15919_16221 , \15920_16222 , \15921_16223 , \15922_16224 , \15923_16225 , \15924_16226 , \15925_16227 , \15926_16228 ,
         \15927_16229 , \15928_16230 , \15929_16231 , \15930_16232 , \15931_16233 , \15932_16234 , \15933_16235 , \15934_16236 , \15935_16237 , \15936_16238 ,
         \15937_16239 , \15938_16240 , \15939_16241 , \15940_16242 , \15941_16243 , \15942_16244 , \15943_16245 , \15944_16246 , \15945_16247 , \15946_16248 ,
         \15947_16249 , \15948_16250 , \15949_16251 , \15950_16252 , \15951_16253 , \15952_16254 , \15953_16255 , \15954_16256 , \15955_16257 , \15956_16258 ,
         \15957_16259 , \15958_16260 , \15959_16261 , \15960_16262 , \15961_16263 , \15962_16264 , \15963 , \15964_16266_nG6597 , \15965_16267 , \15966_16268 ,
         \15967_16269 , \15968_16270 , \15969_16271 , \15970_16272 , \15971_16273 , \15972_16274 , \15973_16275 , \15974_16276 , \15975_16277 , \15976_16278 ,
         \15977_16279 , \15978_16280 , \15979_16281 , \15980_16282 , \15981_16283 , \15982_16284 , \15983_16285 , \15984_16286 , \15985_16287 , \15986_16288 ,
         \15987_16289 , \15988_16290 , \15989_16291 , \15990_16292 , \15991_16293 , \15992_16294 , \15993_16295 , \15994_16296 , \15995 , \15996 ,
         \15997_16299_nG4fb9 , \15998_16300 , \15999_16301 , \16000_16302 , \16001_16303 , \16002_16304 , \16003_16305 , \16004_16306 , \16005_16307 , \16006_16308 ,
         \16007_16309 , \16008_16310 , \16009_16311 , \16010_16312 , \16011_16313 , \16012_16314 , \16013_16315_nG9bf0 , \16014_16316 , \16015_16317 , \16016_16318 ,
         \16017_16319 , \16018_16320 , \16019_16321 , \16020_16322 , \16021_16323 , \16022_16324 , \16023_16325 , \16024_16326 , \16025_16327 , \16026_16328 ,
         \16027_16329 , \16028_16330 , \16029_16331 , \16030_16332 , \16031_16333 , \16032_16334 , \16033_16335 , \16034_16336 , \16035_16337 , \16036_16338 ,
         \16037_16339 , \16038_16340 , \16039_16341 , \16040_16342 , \16041_16343 , \16042_16344 , \16043_16345 , \16044_16346 , \16045_16347 , \16046_16348 ,
         \16047_16349 , \16048_16350 , \16049_16351 , \16050_16352 , \16051_16353 , \16052_16354 , \16053_16355 , \16054_16356 , \16055_16357 , \16056_16358 ,
         \16057_16359 , \16058_16360 , \16059_16361 , \16060_16362 , \16061_16363 , \16062_16364 , \16063_16365 , \16064_16366 , \16065_16367 , \16066_16368 ,
         \16067_16369 , \16068_16370 , \16069_16371 , \16070_16372 , \16071_16373 , \16072_16374 , \16073_16375 , \16074_16376 , \16075_16377 , \16076_16378 ,
         \16077_16379 , \16078_16380 , \16079_16381 , \16080_16382 , \16081_16383 , \16082_16384 , \16083_16385 , \16084_16386 , \16085_16387 , \16086_16388 ,
         \16087_16389 , \16088_16390 , \16089_16391 , \16090_16392 , \16091_16393 , \16092_16394 , \16093_16395 , \16094_16396 , \16095_16397 , \16096_16398 ,
         \16097_16399 , \16098_16400 , \16099_16401 , \16100_16402 , \16101_16403 , \16102_16404 , \16103_16405 , \16104_16406 , \16105_16407 , \16106_16408 ,
         \16107_16409 , \16108_16410 , \16109_16411 , \16110_16412 , \16111_16413 , \16112_16414 , \16113_16415 , \16114_16416 , \16115_16417 , \16116_16418 ,
         \16117_16419 , \16118_16420 , \16119_16421 , \16120_16422 , \16121_16423 , \16122_16424 , \16123_16425 , \16124_16426 , \16125_16427 , \16126_16428 ,
         \16127_16429 , \16128_16430 , \16129_16431 , \16130_16432 , \16131_16433 , \16132_16434 , \16133_16435 , \16134_16436 , \16135_16437 , \16136_16438 ,
         \16137_16439 , \16138_16440 , \16139_16441 , \16140_16442 , \16141_16443 , \16142_16444 , \16143_16445 , \16144_16446 , \16145_16447 , \16146_16448 ,
         \16147_16449 , \16148_16450 , \16149_16451 , \16150_16452 , \16151_16453 , \16152_16454 , \16153_16455 , \16154_16456 , \16155_16457 , \16156_16458 ,
         \16157_16459 , \16158_16460 , \16159_16461 , \16160_16462 , \16161_16463 , \16162_16464 , \16163_16465 , \16164_16466 , \16165_16467 , \16166_16468 ,
         \16167_16469 , \16168_16470 , \16169_16471 , \16170_16472 , \16171_16473 , \16172_16474 , \16173_16475 , \16174_16476 , \16175_16477 , \16176_16478 ,
         \16177_16479 , \16178_16480 , \16179_16481 , \16180_16482 , \16181_16483 , \16182_16484 , \16183_16485 , \16184_16486 , \16185_16487 , \16186 ,
         \16187_16489 , \16188_16490 , \16189_16491 , \16190_16492 , \16191_16493 , \16192_16494 , \16193_16495 , \16194_16496 , \16195_16497 , \16196_16498 ,
         \16197_16499 , \16198_16500 , \16199_16501 , \16200_16502 , \16201_16503 , \16202_16504 , \16203_16505 , \16204_16506 , \16205_16507 , \16206_16508 ,
         \16207_16509 , \16208_16510 , \16209_16511 , \16210_16512 , \16211_16513 , \16212_16514 , \16213_16515 , \16214_16516 , \16215_16517 , \16216_16518 ,
         \16217_16519 , \16218_16520 , \16219_16521 , \16220_16522 , \16221_16523 , \16222_16524 , \16223_16525 , \16224_16526 , \16225_16527 , \16226_16528 ,
         \16227_16529 , \16228_16530 , \16229_16531 , \16230_16532 , \16231_16533 , \16232_16534 , \16233_16535 , \16234_16536 , \16235_16537 , \16236_16538 ,
         \16237_16539 , \16238_16540 , \16239_16541 , \16240_16542 , \16241_16543 , \16242_16544 , \16243_16545 , \16244_16546 , \16245_16547 , \16246_16548 ,
         \16247_16549 , \16248_16550 , \16249_16551 , \16250_16552 , \16251_16553 , \16252_16554 , \16253_16555 , \16254_16556 , \16255_16557 , \16256_16558 ,
         \16257_16559 , \16258_16560 , \16259_16561 , \16260_16562 , \16261_16563 , \16262_16564 , \16263_16565 , \16264_16566 , \16265_16567 , \16266_16568 ,
         \16267_16569 , \16268_16570 , \16269_16571 , \16270_16572 , \16271_16573 , \16272_16574 , \16273_16575 , \16274_16576 , \16275_16577 , \16276_16578 ,
         \16277_16579 , \16278_16580 , \16279_16581 , \16280_16582 , \16281_16583 , \16282_16584 , \16283_16585 , \16284_16586 , \16285_16587 , \16286_16588 ,
         \16287_16589 , \16288_16590 , \16289_16591 , \16290_16592 , \16291_16593 , \16292_16594 , \16293_16595 , \16294_16596 , \16295_16597 , \16296_16598 ,
         \16297_16599 , \16298_16600 , \16299_16601 , \16300_16602 , \16301_16603 , \16302_16604 , \16303_16605 , \16304_16606 , \16305_16607 , \16306_16608 ,
         \16307_16609 , \16308_16610 , \16309_16611 , \16310_16612 , \16311_16613 , \16312_16614 , \16313_16615 , \16314_16616 , \16315_16617 , \16316_16618 ,
         \16317_16619 , \16318 , \16319_16621_nG50c2 , \16320_16622 , \16321_16623 , \16322_16624 , \16323_16625 , \16324_16626 , \16325_16627 , \16326_16628 ,
         \16327_16629 , \16328_16630 , \16329_16631 , \16330_16632 , \16331_16633 , \16332_16634 , \16333_16635 , \16334_16636 , \16335_16637 , \16336_16638 ,
         \16337_16639 , \16338_16640 , \16339_16641 , \16340_16642 , \16341_16643 , \16342_16644 , \16343_16645 , \16344_16646 , \16345_16647 , \16346_16648 ,
         \16347_16649 , \16348_16650 , \16349_16651 , \16350 , \16351 , \16352_16654_nG659a , \16353_16655 , \16354_16656 , \16355_16657 , \16356_16658 ,
         \16357_16659 , \16358_16660 , \16359_16661 , \16360_16662 , \16361_16663 , \16362_16664 , \16363_16665 , \16364_16666 , \16365_16667 , \16366_16668 ,
         \16367_16669 , \16368_16670 , \16369_16671 , \16370_16672 , \16371_16673 , \16372_16674 , \16373_16675 , \16374_16676 , \16375_16677 , \16376_16678 ,
         \16377_16679 , \16378_16680_nG9bed , \16379_16681 , \16380_16682 , \16381_16683 , \16382_16684 , \16383_16685 , \16384_16686 , \16385_16687 , \16386_16688 ,
         \16387_16689 , \16388_16690 , \16389_16691 , \16390_16692 , \16391_16693 , \16392_16694 , \16393_16695 , \16394_16696 , \16395_16697 , \16396_16698 ,
         \16397_16699 , \16398_16700 , \16399_16701 , \16400_16702 , \16401_16703 , \16402_16704 , \16403_15938 , \16404_15939 , \16405_15940 , \16406_16705 ,
         \16407_16706 , \16408_16707 , \16409_16708 , \16410_16709 , \16411_16710 , \16412_16711 , \16413_16712 , \16414_16713 , \16415_16714 , \16416_16715 ,
         \16417_16716 , \16418_16717 , \16419_16718 , \16420_16719 , \16421_16720 , \16422_16721 , \16423_16722 , \16424_16723 , \16425_16724 , \16426_16725 ,
         \16427_16726 , \16428_16727 , \16429_16728 , \16430_16729 , \16431_16730 , \16432_16731 , \16433_16732 , \16434_16733 , \16435_16734 , \16436_16735 ,
         \16437_16736 , \16438_16737 , \16439_16738 , \16440_16739 , \16441_16740 , \16442_16741 , \16443_16742 , \16444_16743 , \16445_16744 , \16446_16745 ,
         \16447_16746 , \16448_16747 , \16449_16748 , \16450_16749 , \16451_16750 , \16452_16751 , \16453_16752 , \16454_16753 , \16455_16754 , \16456_16755 ,
         \16457_16756 , \16458_16757 , \16459_16758 , \16460_16759 , \16461_16760 , \16462_16761 , \16463_16762 , \16464_16763 , \16465_16764 , \16466_16765 ,
         \16467_16766 , \16468_16767 , \16469_16768 , \16470_16769 , \16471_16770 , \16472_16771 , \16473_16772 , \16474_16773 , \16475_16774 , \16476_16775 ,
         \16477_16776 , \16478_16777 , \16479_16778 , \16480_16779 , \16481_16780 , \16482_16781 , \16483_16782 , \16484_16783 , \16485_16784 , \16486_16785 ,
         \16487_16786 , \16488_16787 , \16489_16788 , \16490_16789 , \16491_16790 , \16492_16791 , \16493_16792 , \16494_16793 , \16495_16794 , \16496_16795 ,
         \16497_16796 , \16498_16797 , \16499_16798 , \16500_16799 , \16501_16800 , \16502_16801 , \16503_16802 , \16504_16803 , \16505_16804 , \16506_16805 ,
         \16507_16806 , \16508_16807 , \16509_16808 , \16510_16809 , \16511_16810 , \16512_16811 , \16513_16812 , \16514_16813 , \16515_16814 , \16516_16815 ,
         \16517_16816 , \16518_16817 , \16519_16818 , \16520_16819 , \16521_16820 , \16522_16821 , \16523_16822 , \16524_16823 , \16525_16824 , \16526_16825 ,
         \16527_16826 , \16528_16827 , \16529_16828 , \16530_16829 , \16531_16830 , \16532_16831 , \16533_16832 , \16534_16833 , \16535_16834 , \16536_16835 ,
         \16537_16836 , \16538_16837 , \16539_16838 , \16540_16839 , \16541_16840 , \16542_16841 , \16543_16842 , \16544_16843 , \16545_16844 , \16546_16845 ,
         \16547_16846 , \16548_16847 , \16549_16848 , \16550_16849 , \16551_16850 , \16552_16851 , \16553_16852 , \16554_16853 , \16555_16854 , \16556_16855 ,
         \16557_16856 , \16558_16857 , \16559_16858 , \16560_16859 , \16561_16860 , \16562_16861 , \16563_16862 , \16564_16863 , \16565_16864 , \16566_16865 ,
         \16567_16866 , \16568_16867 , \16569_16868 , \16570_16869 , \16571_16870 , \16572_16871 , \16573_16872 , \16574_16873 , \16575_16874 , \16576_16875 ,
         \16577_16876 , \16578 , \16579_16878 , \16580_16879 , \16581_16880 , \16582_16881 , \16583_16882 , \16584_16883 , \16585_16884 , \16586_16885 ,
         \16587_16886 , \16588_16887 , \16589_16888 , \16590_16889 , \16591_16890 , \16592_16891 , \16593_16892 , \16594_16893 , \16595_16894 , \16596_16895 ,
         \16597_16896 , \16598_16897 , \16599_16898 , \16600_16899 , \16601_16900 , \16602_16901 , \16603_16902 , \16604_16903 , \16605_16904 , \16606_16905 ,
         \16607_16906 , \16608_16907 , \16609_16908 , \16610_16909 , \16611_16910 , \16612_16911 , \16613_16912 , \16614_16913 , \16615_16914 , \16616_16915 ,
         \16617_16916 , \16618_16917 , \16619_16918 , \16620_16919 , \16621_16920 , \16622_16921 , \16623_16922 , \16624_16923 , \16625_16924 , \16626_16925 ,
         \16627_16926 , \16628_16927 , \16629_16928 , \16630_16929 , \16631_16930 , \16632_16931 , \16633_16932 , \16634_16933 , \16635_16934 , \16636_16935 ,
         \16637_16936 , \16638_16937 , \16639_16938 , \16640_16939 , \16641_16940 , \16642_16941 , \16643_16942 , \16644_16943 , \16645_16944 , \16646_16945 ,
         \16647_16946 , \16648_16947 , \16649_16948 , \16650_16949 , \16651_16950 , \16652_16951 , \16653_16952 , \16654_16953 , \16655_16954 , \16656_16955 ,
         \16657_16956 , \16658_16957 , \16659_16958 , \16660_16959 , \16661_16960 , \16662_16961 , \16663_16962 , \16664_16963 , \16665_16964 , \16666_16965 ,
         \16667_16966 , \16668_16967 , \16669_16968 , \16670_16969 , \16671_16970 , \16672_16971 , \16673_16972 , \16674_16973 , \16675_16974 , \16676_16975 ,
         \16677_16976 , \16678_16977 , \16679_16978 , \16680_16979 , \16681_16980 , \16682_16981 , \16683_16982 , \16684_16983 , \16685_16984 , \16686_16985 ,
         \16687_16986 , \16688_16987 , \16689_16988 , \16690_16989 , \16691_16990 , \16692_16991 , \16693_16992 , \16694_16993 , \16695_16994 , \16696_16995 ,
         \16697_16996 , \16698_16997 , \16699_16998 , \16700_16999 , \16701_17000 , \16702_17001 , \16703_17002 , \16704_17003 , \16705_17004 , \16706_17005 ,
         \16707_17006 , \16708_17007 , \16709_17008 , \16710_17009 , \16711 , \16712_17011 , \16713_17012 , \16714_17013 , \16715_17014 , \16716_17015 ,
         \16717_17016 , \16718_17017 , \16719_17018 , \16720_17019 , \16721_17020 , \16722_17021 , \16723_17022 , \16724_17023 , \16725_17024 , \16726_17025 ,
         \16727_17026 , \16728_17027 , \16729_17028 , \16730_17029 , \16731_17030 , \16732_17031 , \16733_17032 , \16734_17033 , \16735_17034 , \16736_17035 ,
         \16737_17036 , \16738_17037 , \16739_17038 , \16740_17039 , \16741_17040 , \16742_17041 , \16743_17042 , \16744_17043 , \16745_17044 , \16746_17045 ,
         \16747_17046 , \16748_17047 , \16749_17048 , \16750_17049 , \16751_17050 , \16752_17051 , \16753_17052 , \16754_17053 , \16755_17054 , \16756_17055 ,
         \16757_17056 , \16758_17057 , \16759_17058 , \16760_17059 , \16761_17060 , \16762_17061 , \16763_17062 , \16764_17063 , \16765_17064 , \16766_17065 ,
         \16767_17066 , \16768_17067 , \16769_17068 , \16770_17069 , \16771_17070 , \16772_17071 , \16773_17072 , \16774_17073 , \16775_17074 , \16776_17075 ,
         \16777_17076 , \16778_17077 , \16779_17078 , \16780_17079 , \16781_17080 , \16782_17081 , \16783_17082 , \16784_17083 , \16785_17084 , \16786_17085 ,
         \16787_17086 , \16788_17087 , \16789_17088 , \16790_17089 , \16791_17090 , \16792_17091 , \16793_17092 , \16794_17093 , \16795_17094 , \16796_17095 ,
         \16797_17096 , \16798_17097 , \16799_17098 , \16800_17099 , \16801_17100 , \16802_17101 , \16803_17102 , \16804_17103 , \16805_17104 , \16806_17105 ,
         \16807_17106 , \16808_17107 , \16809_17108 , \16810_17109 , \16811_17110 , \16812_17111 , \16813_17112 , \16814_17113 , \16815_17114 , \16816_17115 ,
         \16817_17116 , \16818_17117 , \16819_17118 , \16820_17119 , \16821_17120 , \16822_17121 , \16823_17122 , \16824_17123 , \16825_17124 , \16826_17125 ,
         \16827_17126 , \16828_17127 , \16829_17128 , \16830_17129 , \16831_17130 , \16832_17131 , \16833_17132 , \16834_17133 , \16835_17134 , \16836_17135 ,
         \16837_17136 , \16838_17137 , \16839_17138 , \16840_17139 , \16841_17140 , \16842_17141 , \16843_17142 , \16844_17143 , \16845 , \16846_17145 ,
         \16847_17146 , \16848_17147 , \16849_17148 , \16850_17149 , \16851_17150 , \16852_17151 , \16853_17152 , \16854_17153 , \16855_17154 , \16856_17155 ,
         \16857_17156 , \16858_17157 , \16859_17158 , \16860_17159 , \16861_17160 , \16862_17161 , \16863_17162 , \16864_17163 , \16865_17164 , \16866_17165 ,
         \16867_17166 , \16868_17167 , \16869_17168 , \16870_17169 , \16871_17170 , \16872_17171 , \16873_17172 , \16874_17173 , \16875_17174 , \16876_17175 ,
         \16877_17176 , \16878_17177 , \16879_17178 , \16880_17179 , \16881_17180 , \16882_17181 , \16883_17182 , \16884_17183 , \16885_17184 , \16886_17185 ,
         \16887_17186 , \16888_17187 , \16889_17188 , \16890_17189 , \16891_17190 , \16892_17191 , \16893_17192 , \16894_17193 , \16895_17194 , \16896_17195 ,
         \16897_17196 , \16898_17197 , \16899_17198 , \16900_17199 , \16901_17200 , \16902_17201 , \16903_17202 , \16904_17203 , \16905_17204 , \16906_17205 ,
         \16907_17206 , \16908_17207 , \16909_17208 , \16910_17209 , \16911_17210 , \16912_17211 , \16913_17212 , \16914_17213 , \16915_17214 , \16916_17215 ,
         \16917_17216 , \16918_17217 , \16919_17218 , \16920_17219 , \16921_17220 , \16922_17221 , \16923_17222 , \16924_17223 , \16925_17224 , \16926_17225 ,
         \16927_17226 , \16928_17227 , \16929_17228 , \16930_17229 , \16931_17230 , \16932_17231 , \16933_17232 , \16934_17233 , \16935_17234 , \16936_17235 ,
         \16937_17236 , \16938_17237 , \16939_17238 , \16940_17239 , \16941_17240 , \16942_17241 , \16943_17242 , \16944_17243 , \16945_17244 , \16946_17245 ,
         \16947_17246 , \16948_17247 , \16949_17248 , \16950_17249 , \16951_17250 , \16952_17251 , \16953_17252 , \16954_17253 , \16955_17254 , \16956_17255 ,
         \16957_17256 , \16958_17257 , \16959_17258 , \16960_17259 , \16961_17260 , \16962_17261 , \16963_17262 , \16964_17263 , \16965_17264 , \16966_17265 ,
         \16967_17266 , \16968_17267 , \16969_17268 , \16970_17269 , \16971_17270 , \16972_17271 , \16973_17272 , \16974_17273 , \16975_17274 , \16976_17275 ,
         \16977_17276 , \16978 , \16979_17278 , \16980_17279 , \16981_17280 , \16982_17281 , \16983_17282 , \16984_17283 , \16985_17284 , \16986_17285 ,
         \16987_17286 , \16988_17287 , \16989_17288_nG4430 , \16990_17289 , \16991_17290 , \16992_17291_nG4433 , \16993_17292 , \16994_17293 , \16995_17294 , \16996_17298 ,
         \16997_17299 , \16998_17300 , \16999_17301 , \17000_17302 , \17001_17303 , \17002_17304 , \17003_17305 , \17004_17306 , \17005_17307 , \17006_17308 ,
         \17007_17309 , \17008_17310 , \17009_17311 , \17010_17312 , \17011_17313 , \17012_17314 , \17013_17315 , \17014_17316 , \17015_17317 , \17016_17318 ,
         \17017_17319 , \17018_17320 , \17019_17321 , \17020_17322 , \17021_17323 , \17022_17324 , \17023_17325 , \17024_17326 , \17025_17327 , \17026_17328 ,
         \17027_17329 , \17028_17330 , \17029_17331 , \17030_17332 , \17031_17333 , \17032_17334 , \17033_17335 , \17034_17336 , \17035_17337 , \17036_17338 ,
         \17037_17339 , \17038_17340 , \17039_17341 , \17040_17342 , \17041_17343 , \17042_17344 , \17043_17345 , \17044_17346 , \17045_17347 , \17046_17348 ,
         \17047_17349 , \17048_17350 , \17049_17351 , \17050_17352 , \17051_17353 , \17052_17354 , \17053_17355 , \17054_17356 , \17055_17357 , \17056_17358 ,
         \17057_17359 , \17058_17360 , \17059_17361 , \17060_17362 , \17061_17363 , \17062_17364 , \17063_17365 , \17064_17366 , \17065_17367 , \17066_17368 ,
         \17067_17369 , \17068_17370 , \17069_17371 , \17070_17372 , \17071_17373 , \17072_17374 , \17073_17375 , \17074_17376 , \17075_17377 , \17076_17378 ,
         \17077_17379 , \17078_17380 , \17079_17381 , \17080_17382 , \17081_17383 , \17082_17384 , \17083_17385 , \17084_17386 , \17085_17387 , \17086_17388 ,
         \17087_17389 , \17088_17390 , \17089_17391 , \17090_17392 , \17091_17393 , \17092_17394 , \17093_17395 , \17094_17396 , \17095_17397 , \17096_17398 ,
         \17097_17399 , \17098_17400 , \17099_17401 , \17100_17402 , \17101_17403 , \17102_17404 , \17103_17405 , \17104_17406 , \17105_17407 , \17106_17408 ,
         \17107_17409 , \17108_17410 , \17109_17411 , \17110_17412 , \17111_17413 , \17112_17414 , \17113_17415 , \17114_17416 , \17115_17417 , \17116_17418 ,
         \17117_17419 , \17118_17420 , \17119_17421 , \17120_17422 , \17121_17423 , \17122_17424 , \17123_17425 , \17124_17426 , \17125_17427 , \17126_17428 ,
         \17127_17429 , \17128_17430 , \17129_17431 , \17130_17432 , \17131_17433 , \17132_17434 , \17133_17435 , \17134_17436 , \17135_17437 , \17136_17438 ,
         \17137_17439 , \17138_17440 , \17139_17441 , \17140_17442 , \17141_17443 , \17142_17444 , \17143_17445 , \17144_17446 , \17145_17447 , \17146_17448 ,
         \17147_17449 , \17148_17450 , \17149_17451 , \17150_17452 , \17151_17453 , \17152_17454 , \17153_17455 , \17154_17456 , \17155_17457 , \17156_17458 ,
         \17157_17459 , \17158_17460 , \17159_17461 , \17160_17462 , \17161_17463 , \17162_17464 , \17163_17465 , \17164_17466 , \17165_17467 , \17166_17468 ,
         \17167_17469 , \17168_17470 , \17169_17471 , \17170_17472 , \17171_17473 , \17172_17474 , \17173_17475 , \17174_17476 , \17175_17477 , \17176_17478 ,
         \17177_17479 , \17178_17480 , \17179_17481 , \17180_17482 , \17181_17483 , \17182_17484 , \17183_17485 , \17184_17486 , \17185_17487 , \17186_17488 ,
         \17187_17489 , \17188_17490 , \17189_17491 , \17190_17492 , \17191 , \17192_17494 , \17193_17495 , \17194_17496 , \17195_17497 , \17196_17498 ,
         \17197_17499 , \17198_17500 , \17199_17501 , \17200_17502 , \17201_17503 , \17202_17504 , \17203_17505 , \17204_17506 , \17205_17507 , \17206_17508 ,
         \17207_17509 , \17208_17510 , \17209_17511 , \17210_17512 , \17211_17513 , \17212_17514 , \17213_17515 , \17214_17516 , \17215_17517 , \17216_17518 ,
         \17217_17519 , \17218_17520 , \17219_17521 , \17220_17522 , \17221_17523 , \17222_17524 , \17223_17525 , \17224_17526 , \17225_17527 , \17226_17528 ,
         \17227_17529 , \17228_17530 , \17229_17531 , \17230_17532 , \17231_17533 , \17232_17534 , \17233_17535 , \17234_17536 , \17235_17537 , \17236_17538 ,
         \17237_17539 , \17238_17540 , \17239_17541 , \17240_17542 , \17241_17543 , \17242_17544 , \17243_17545 , \17244_17546 , \17245_17547 , \17246_17548 ,
         \17247_17549 , \17248_17550 , \17249_17551 , \17250_17552 , \17251_17553 , \17252_17554 , \17253_17555 , \17254_17556 , \17255_17557 , \17256_17558 ,
         \17257_17559 , \17258_17560 , \17259_17561 , \17260_17562 , \17261_17563 , \17262_17564 , \17263_17565 , \17264_17566 , \17265_17567 , \17266_17568 ,
         \17267_17569 , \17268_17570 , \17269_17571 , \17270_17572 , \17271_17573 , \17272_17574 , \17273_17575 , \17274_17576 , \17275_17577 , \17276_17578 ,
         \17277_17579 , \17278_17580 , \17279_17581 , \17280_17582 , \17281_17583 , \17282_17584 , \17283_17585 , \17284_17586 , \17285_17587 , \17286_17588 ,
         \17287_17589 , \17288_17590 , \17289_17591 , \17290_17592 , \17291_17593 , \17292_17594 , \17293_17595 , \17294_17596 , \17295_17597 , \17296_17598 ,
         \17297_17599 , \17298_17600 , \17299_17601 , \17300_17602 , \17301_17603 , \17302_17604 , \17303_17605 , \17304_17606 , \17305_17607 , \17306_17608 ,
         \17307_17609 , \17308_17610 , \17309_17611 , \17310_17612 , \17311_17613 , \17312_17614 , \17313_17615 , \17314_17616 , \17315_17617 , \17316_17618 ,
         \17317_17619 , \17318_17620 , \17319_17621 , \17320_17622 , \17321_17623 , \17322_17624 , \17323 , \17324_17626_nG659d , \17325_17627 , \17326_17628 ,
         \17327_17629 , \17328_17630 , \17329_17631 , \17330_17632 , \17331_17633 , \17332_17634 , \17333_17635 , \17334_17636 , \17335_17637 , \17336_17638 ,
         \17337_17639 , \17338_17640 , \17339_17641 , \17340_17642 , \17341_17643 , \17342_17644 , \17343_17645 , \17344_17646 , \17345_17647 , \17346_17648 ,
         \17347_17649 , \17348_17650 , \17349 , \17350 , \17351_17653_nG51cb , \17352_17654 , \17353_17655 , \17354_17656 , \17355_17657 , \17356_17658 ,
         \17357_17659 , \17358_17660 , \17359_17661 , \17360_17662 , \17361_17663 , \17362_17664 , \17363_17665_nG9bea , \17364_17666 , \17365_17667 , \17366_17668 ,
         \17367_17669 , \17368_17670 , \17369_17671 , \17370_17672 , \17371_17673 , \17372_17674 , \17373_17675 , \17374_17676 , \17375_17677 , \17376_17678 ,
         \17377_17679 , \17378_17680 , \17379_17681 , \17380_17682 , \17381_17683 , \17382_17684 , \17383_17685 , \17384_17686 , \17385_17687 , \17386_17688 ,
         \17387_17689 , \17388_17690 , \17389_17691 , \17390_17692 , \17391_17693 , \17392_17694 , \17393_17695 , \17394_17696 , \17395_17697 , \17396_17698 ,
         \17397_17699 , \17398_17700 , \17399_17701 , \17400_17702 , \17401_17703 , \17402_17704 , \17403_17705 , \17404_17706 , \17405_17707 , \17406_17708 ,
         \17407_17709 , \17408_17710 , \17409_17711 , \17410_17712 , \17411_17713 , \17412_17714 , \17413_17715 , \17414_17716 , \17415_17717 , \17416_17718 ,
         \17417_17719 , \17418_17720 , \17419_17721 , \17420_17722 , \17421_17723 , \17422_17724 , \17423_17725 , \17424_17726 , \17425_17727 , \17426_17728 ,
         \17427_17729 , \17428_17730 , \17429_17731 , \17430_17732 , \17431_17733 , \17432_17734 , \17433_17735 , \17434_17736 , \17435_17295 , \17436_17296 ,
         \17437_17297 , \17438_17737 , \17439_17738 , \17440_17739 , \17441_17740 , \17442_17741 , \17443_17742 , \17444_17743 , \17445_17744 , \17446_17745 ,
         \17447_17746 , \17448_17747 , \17449_17748 , \17450_17749 , \17451_17750 , \17452_17751 , \17453_17752 , \17454_17753 , \17455_17754 , \17456_17755 ,
         \17457_17756 , \17458_17757 , \17459_17758 , \17460_17759 , \17461_17760 , \17462_17761 , \17463_17762 , \17464_17763 , \17465_17764 , \17466_17765 ,
         \17467_17766 , \17468_17767 , \17469_17768 , \17470_17769 , \17471_17770 , \17472_17771 , \17473_17772 , \17474_17773 , \17475_17774 , \17476_17775 ,
         \17477_17776 , \17478_17777 , \17479_17778 , \17480_17779 , \17481_17780 , \17482_17781 , \17483_17782 , \17484_17783 , \17485_17784 , \17486_17785 ,
         \17487_17786 , \17488_17787 , \17489_17788 , \17490_17789 , \17491_17790 , \17492_17791 , \17493_17792 , \17494_17793 , \17495_17794 , \17496_17795 ,
         \17497_17796 , \17498_17797 , \17499_17798 , \17500_17799 , \17501_17800 , \17502_17801 , \17503_17802 , \17504_17803 , \17505_17804 , \17506_17805 ,
         \17507_17806 , \17508_17807 , \17509_17808 , \17510_17809 , \17511_17810 , \17512_17811 , \17513_17812 , \17514_17813 , \17515_17814 , \17516_17815 ,
         \17517_17816 , \17518_17817 , \17519_17818 , \17520_17819 , \17521_17820 , \17522_17821 , \17523_17822 , \17524_17823 , \17525_17824 , \17526_17825 ,
         \17527_17826 , \17528_17827 , \17529_17828 , \17530_17829 , \17531_17830 , \17532_17831 , \17533_17832 , \17534_17833 , \17535_17834 , \17536_17835 ,
         \17537_17836 , \17538_17837 , \17539_17838 , \17540_17839 , \17541_17840 , \17542_17841 , \17543_17842 , \17544_17843 , \17545_17844 , \17546_17845 ,
         \17547_17846 , \17548_17847 , \17549_17848 , \17550_17849 , \17551_17850 , \17552_17851 , \17553_17852 , \17554_17853 , \17555_17854 , \17556_17855 ,
         \17557_17856 , \17558_17857 , \17559_17858 , \17560_17859 , \17561_17860 , \17562_17861 , \17563_17862 , \17564_17863 , \17565_17864 , \17566_17865 ,
         \17567_17866 , \17568_17867 , \17569_17868 , \17570_17869 , \17571_17870 , \17572_17871 , \17573_17872 , \17574_17873 , \17575_17874 , \17576_17875 ,
         \17577_17876 , \17578_17877 , \17579_17878 , \17580_17879 , \17581_17880 , \17582_17881 , \17583_17882 , \17584_17883 , \17585_17884 , \17586_17885 ,
         \17587_17886 , \17588_17887 , \17589_17888 , \17590_17889 , \17591_17890 , \17592_17891 , \17593_17892 , \17594_17893 , \17595_17894 , \17596_17895 ,
         \17597_17896 , \17598_17897 , \17599_17898 , \17600_17899 , \17601_17900 , \17602 , \17603_17902 , \17604_17903 , \17605_17904 , \17606_17905 ,
         \17607_17906 , \17608_17907 , \17609_17908 , \17610_17909 , \17611_17910 , \17612_17911 , \17613_17912 , \17614_17913 , \17615_17914 , \17616_17915 ,
         \17617_17916 , \17618_17917 , \17619_17918 , \17620_17919 , \17621_17920 , \17622_17921 , \17623_17922 , \17624_17923 , \17625_17924 , \17626_17925 ,
         \17627_17926 , \17628_17927 , \17629_17928 , \17630_17929 , \17631_17930 , \17632_17931 , \17633_17932 , \17634_17933 , \17635_17934 , \17636_17935 ,
         \17637_17936 , \17638_17937 , \17639_17938 , \17640_17939 , \17641_17940 , \17642_17941 , \17643_17942 , \17644_17943 , \17645_17944 , \17646_17945 ,
         \17647_17946 , \17648_17947 , \17649_17948 , \17650_17949 , \17651_17950 , \17652_17951 , \17653_17952 , \17654_17953 , \17655_17954 , \17656_17955 ,
         \17657_17956 , \17658_17957 , \17659_17958 , \17660_17959 , \17661_17960 , \17662_17961 , \17663_17962 , \17664_17963 , \17665_17964 , \17666_17965 ,
         \17667_17966 , \17668_17967 , \17669_17968 , \17670_17969 , \17671_17970 , \17672_17971 , \17673_17972 , \17674_17973 , \17675_17974 , \17676_17975 ,
         \17677_17976 , \17678_17977 , \17679_17978 , \17680_17979 , \17681_17980 , \17682_17981 , \17683_17982 , \17684_17983 , \17685_17984 , \17686_17985 ,
         \17687_17986 , \17688_17987 , \17689_17988 , \17690_17989 , \17691_17990 , \17692_17991 , \17693_17992 , \17694_17993 , \17695_17994 , \17696_17995 ,
         \17697_17996 , \17698_17997 , \17699_17998 , \17700_17999 , \17701_18000 , \17702_18001 , \17703_18002 , \17704_18003 , \17705_18004 , \17706_18005 ,
         \17707_18006 , \17708_18007 , \17709_18008 , \17710_18009 , \17711_18010 , \17712_18011 , \17713_18012 , \17714_18013 , \17715_18014 , \17716_18015 ,
         \17717_18016 , \17718_18017 , \17719_18018 , \17720_18019 , \17721_18020 , \17722_18021 , \17723_18022 , \17724_18023 , \17725_18024 , \17726_18025 ,
         \17727_18026 , \17728_18027 , \17729_18028 , \17730_18029 , \17731_18030 , \17732_18031 , \17733_18032 , \17734 , \17735_18034_nG65a0 , \17736_18035 ,
         \17737_18036 , \17738_18037 , \17739_18038 , \17740_18039 , \17741 , \17742 , \17743_18042_nG52d4 , \17744_18043 , \17745_18044 , \17746_18045 ,
         \17747_18046 , \17748_18047 , \17749_18048 , \17750_18049 , \17751_18050 , \17752_18051 , \17753_18052 , \17754_18053 , \17755_18054 , \17756_18055 ,
         \17757_18056 , \17758_18057 , \17759_18058 , \17760_18059 , \17761_18060 , \17762_18061 , \17763_18062 , \17764_18063 , \17765_18064 , \17766_18065 ,
         \17767_18066 , \17768_18067 , \17769_18068 , \17770_18069 , \17771_18070 , \17772_18071 , \17773_18072 , \17774_18073 , \17775_18074 , \17776_18075 ,
         \17777_18076 , \17778_18077 , \17779_18078 , \17780_18079 , \17781_18080 , \17782_18081 , \17783_18082 , \17784_18083 , \17785_18084 , \17786_18085 ,
         \17787_18086 , \17788_18087 , \17789_18088 , \17790_18089 , \17791_18090 , \17792_18091 , \17793_18092 , \17794_18093 , \17795_18094 , \17796_18095 ,
         \17797_18096 , \17798_18097 , \17799_18098 , \17800_18099 , \17801_18100 , \17802_18101 , \17803_18102 , \17804_18103 , \17805_18104 , \17806_18105 ,
         \17807_18106 , \17808_18107_nG9be7 , \17809_18108 , \17810_18109 , \17811_18110 , \17812_18111 , \17813_18112 , \17814_18113 , \17815_18114 , \17816_18115 ,
         \17817_18116 , \17818_18117 , \17819_18118 , \17820_18119 , \17821_18120 , \17822_18121 , \17823_18122 , \17824_18123 , \17825_18124 , \17826_18125 ,
         \17827_18126 , \17828_18127 , \17829_18128 , \17830_18129 , \17831_18130 , \17832_18131 , \17833_18132 , \17834_18133 , \17835_18134 , \17836_18135 ,
         \17837_18136 , \17838_18137 , \17839_18138 , \17840_18139 , \17841_18140 , \17842_18141 , \17843_18142 , \17844_18143 , \17845_18144 , \17846_18145 ,
         \17847_18146 , \17848_18147 , \17849_18148 , \17850_18149 , \17851_18150 , \17852_18151 , \17853_18152 , \17854_18153 , \17855_18154 , \17856_18155 ,
         \17857_18156 , \17858_18157 , \17859_18158 , \17860_18159 , \17861_18160 , \17862_18161 , \17863_18162 , \17864_18163 , \17865_18164 , \17866_18165 ,
         \17867_18166 , \17868_18167 , \17869_18168 , \17870_18169 , \17871_18170 , \17872_18171 , \17873_18172 , \17874_18173 , \17875_18174 , \17876_18175 ,
         \17877_18176 , \17878_18177 , \17879_18178 , \17880_18179 , \17881_18180 , \17882_18181 , \17883_18182 , \17884_18183 , \17885_18184 , \17886_18185 ,
         \17887_18186 , \17888_18187 , \17889_18188 , \17890_18189 , \17891_18190 , \17892_18191 , \17893_18192 , \17894_18193 , \17895_18194 , \17896_18195 ,
         \17897_18196 , \17898_18197 , \17899_18198 , \17900_18199 , \17901_18200 , \17902_18201 , \17903_18202 , \17904_18203 , \17905_18204 , \17906_18205 ,
         \17907_18206 , \17908_18207 , \17909_18208 , \17910_18209 , \17911_18210 , \17912_18211 , \17913_18212 , \17914_18213 , \17915_18214 , \17916_18215 ,
         \17917_18216 , \17918_18217 , \17919_18218 , \17920_18219 , \17921_18220 , \17922_18221 , \17923_18222 , \17924_18223 , \17925_18224 , \17926_18225 ,
         \17927_18226 , \17928_18227 , \17929_18228 , \17930_18229 , \17931_18230 , \17932_18231 , \17933_18232 , \17934_18233 , \17935_18234 , \17936_18235 ,
         \17937_18236 , \17938_18237 , \17939_18238 , \17940_18239 , \17941_18240 , \17942_18241 , \17943_18242 , \17944_18243 , \17945_18244 , \17946_18245 ,
         \17947_18246 , \17948_18247 , \17949_18248 , \17950_18249 , \17951_18250 , \17952_18251 , \17953_18252 , \17954_18253 , \17955_18254 , \17956_18255 ,
         \17957_18256 , \17958_18257 , \17959_18258 , \17960_18259 , \17961_18260 , \17962_18261 , \17963_18262 , \17964_18263 , \17965_18264 , \17966_18265 ,
         \17967_18266 , \17968_18267 , \17969_18268 , \17970_18269 , \17971_18270 , \17972_18271 , \17973_18272 , \17974_18273 , \17975_18274 , \17976_18275 ,
         \17977_18276 , \17978_18277 , \17979_18278 , \17980_18279 , \17981_18280 , \17982_18281 , \17983 , \17984_18283 , \17985_18284 , \17986_18285 ,
         \17987_18286 , \17988_18287 , \17989_18288 , \17990_18289 , \17991_18290 , \17992_18291 , \17993_18292 , \17994_18293 , \17995_18294 , \17996_18295 ,
         \17997_18296 , \17998_18297 , \17999_18298 , \18000_18299 , \18001_18300 , \18002_18301 , \18003_18302 , \18004_18303 , \18005_18304 , \18006_18305 ,
         \18007_18306 , \18008_18307 , \18009_18308 , \18010_18309 , \18011_18310 , \18012_18311 , \18013_18312 , \18014_18313 , \18015_18314 , \18016_18315 ,
         \18017_18316 , \18018_18317 , \18019_18318 , \18020_18319 , \18021_18320 , \18022_18321 , \18023_18322 , \18024_18323 , \18025_18324 , \18026_18325 ,
         \18027_18326 , \18028_18327 , \18029_18328 , \18030_18329 , \18031_18330 , \18032_18331 , \18033_18332 , \18034_18333 , \18035_18334 , \18036_18335 ,
         \18037_18336 , \18038_18337 , \18039_18338 , \18040_18339 , \18041_18340 , \18042_18341 , \18043_18342 , \18044_18343 , \18045_18344 , \18046_18345 ,
         \18047_18346 , \18048_18347 , \18049_18348 , \18050_18349 , \18051_18350 , \18052_18351 , \18053_18352 , \18054_18353 , \18055_18354 , \18056_18355 ,
         \18057_18356 , \18058_18357 , \18059_18358 , \18060_18359 , \18061_18360 , \18062_18361 , \18063_18362 , \18064_18363 , \18065_18364 , \18066_18365 ,
         \18067_18366 , \18068_18367 , \18069_18368 , \18070_18369 , \18071_18370 , \18072_18371 , \18073_18372 , \18074_18373 , \18075_18374 , \18076_18375 ,
         \18077_18376 , \18078_18377 , \18079_18378 , \18080_18379 , \18081_18380 , \18082_18381 , \18083_18382 , \18084_18383 , \18085_18384 , \18086_18385 ,
         \18087_18386 , \18088_18387 , \18089_18388 , \18090_18389 , \18091_18390 , \18092_18391 , \18093_18392 , \18094_18393 , \18095_18394 , \18096_18395 ,
         \18097_18396 , \18098_18397 , \18099_18398 , \18100_18399 , \18101_18400 , \18102_18401 , \18103_18402 , \18104_18403 , \18105_18404 , \18106_18405 ,
         \18107_18406 , \18108_18407 , \18109_18408 , \18110_18409 , \18111_18410 , \18112_18411 , \18113_18412 , \18114_18413 , \18115_18414 , \18116 ,
         \18117_18416 , \18118_18417 , \18119_18418 , \18120_18419 , \18121_18420 , \18122_18421 , \18123_18422 , \18124_18423 , \18125_18424 , \18126_18425 ,
         \18127_18426 , \18128_18427 , \18129_18428 , \18130_18429 , \18131_18430 , \18132_18431 , \18133_18432 , \18134_18433 , \18135_18434 , \18136_18435 ,
         \18137_18436 , \18138_18437 , \18139_18438 , \18140_18439 , \18141_18440 , \18142_18441 , \18143_18442 , \18144_18443 , \18145_18444 , \18146_18445 ,
         \18147_18446 , \18148_18447 , \18149_18448 , \18150_18449 , \18151_18450 , \18152_18451 , \18153_18452 , \18154_18453 , \18155_18454 , \18156_18455 ,
         \18157_18456 , \18158_18457 , \18159_18458 , \18160_18459 , \18161_18460 , \18162_18461 , \18163_18462 , \18164_18463 , \18165_18464 , \18166_18465 ,
         \18167_18466 , \18168_18467 , \18169_18468 , \18170_18469 , \18171_18470 , \18172_18471 , \18173_18472 , \18174_18473 , \18175_18474 , \18176_18475 ,
         \18177_18476 , \18178_18477 , \18179_18478 , \18180_18479 , \18181_18480 , \18182_18481 , \18183_18482 , \18184_18483 , \18185_18484 , \18186_18485 ,
         \18187_18486 , \18188_18487 , \18189_18488 , \18190_18489 , \18191_18490 , \18192_18491 , \18193_18492 , \18194_18493 , \18195_18494 , \18196_18495 ,
         \18197_18496 , \18198_18497 , \18199_18498 , \18200_18499 , \18201_18500 , \18202_18501 , \18203_18502 , \18204_18503 , \18205_18504 , \18206_18505 ,
         \18207_18506 , \18208_18507 , \18209_18508 , \18210_18509 , \18211_18510 , \18212_18511 , \18213_18512 , \18214_18513 , \18215_18514 , \18216_18515 ,
         \18217_18516 , \18218_18517 , \18219_18518 , \18220_18519 , \18221_18520 , \18222_18521 , \18223_18522 , \18224_18523 , \18225_18524 , \18226_18525 ,
         \18227_18526 , \18228_18527 , \18229_18528 , \18230_18529 , \18231_18530 , \18232_18531 , \18233_18532 , \18234_18533 , \18235_18534 , \18236_18535 ,
         \18237_18536 , \18238_18537 , \18239_18538 , \18240_18539 , \18241_18540 , \18242_18541 , \18243_18542 , \18244_18543 , \18245_18544 , \18246_18545 ,
         \18247_18546 , \18248_18547 , \18249_18548 , \18250 , \18251_18550 , \18252_18551 , \18253_18552 , \18254_18553 , \18255_18554 , \18256_18555 ,
         \18257_18556 , \18258_18557 , \18259_18558 , \18260_18559 , \18261_18560 , \18262_18561 , \18263_18562 , \18264_18563 , \18265_18564 , \18266_18565 ,
         \18267_18566 , \18268_18567 , \18269_18568 , \18270_18569 , \18271_18570 , \18272_18571 , \18273_18572 , \18274_18573 , \18275_18574 , \18276_18575 ,
         \18277_18576 , \18278_18577 , \18279_18578 , \18280_18579 , \18281_18580 , \18282_18581 , \18283_18582 , \18284_18583 , \18285_18584 , \18286_18585 ,
         \18287_18586 , \18288_18587 , \18289_18588 , \18290_18589 , \18291_18590 , \18292_18591 , \18293_18592 , \18294_18593 , \18295_18594 , \18296_18595 ,
         \18297_18596 , \18298_18597 , \18299_18598 , \18300_18599 , \18301_18600 , \18302_18601 , \18303_18602 , \18304_18603 , \18305_18604 , \18306_18605 ,
         \18307_18606 , \18308_18607 , \18309_18608 , \18310_18609 , \18311_18610 , \18312_18611 , \18313_18612 , \18314_18613 , \18315_18614 , \18316_18615 ,
         \18317_18616 , \18318_18617 , \18319_18618 , \18320_18619 , \18321_18620 , \18322_18621 , \18323_18622 , \18324_18623 , \18325_18624 , \18326_18625 ,
         \18327_18626 , \18328_18627 , \18329_18628 , \18330_18629 , \18331_18630 , \18332_18631 , \18333_18632 , \18334_18633 , \18335_18634 , \18336_18635 ,
         \18337_18636 , \18338_18637 , \18339_18638 , \18340_18639 , \18341_18640 , \18342_18641 , \18343_18642 , \18344_18643 , \18345_18644 , \18346_18645 ,
         \18347_18646 , \18348_18647 , \18349_18648 , \18350_18649 , \18351_18650 , \18352_18651 , \18353_18652 , \18354_18653 , \18355_18654 , \18356_18655 ,
         \18357_18656 , \18358_18657 , \18359_18658 , \18360_18659 , \18361_18660 , \18362_18661 , \18363_18662 , \18364_18663 , \18365_18664 , \18366_18665 ,
         \18367_18666 , \18368_18667 , \18369_18668 , \18370_18669 , \18371_18670 , \18372_18671 , \18373_18672 , \18374_18673 , \18375_18674 , \18376_18675 ,
         \18377_18676 , \18378_18677 , \18379_18678 , \18380_18679 , \18381_18680 , \18382_18681 , \18383 , \18384_18683 , \18385_18684 , \18386_18685 ,
         \18387_18686 , \18388_18687 , \18389_18688 , \18390_18689 , \18391_18690 , \18392_18691 , \18393_18692 , \18394_18693_nG442a , \18395_18694 , \18396_18695 ,
         \18397_18696_nG442d , \18398_18697 , \18399_18698 , \18400_18699 , \18401_18703 , \18402_18704 , \18403_18705 , \18404_18706 , \18405_18707 , \18406_18708 ,
         \18407_18709 , \18408_18710 , \18409_18711 , \18410_18712 , \18411_18713 , \18412_18714 , \18413_18715 , \18414_18716 , \18415_18717 , \18416_18718 ,
         \18417_18719 , \18418_18720 , \18419_18721 , \18420_18722 , \18421_18723 , \18422_18724 , \18423_18725 , \18424_18726 , \18425_18727 , \18426_18728 ,
         \18427_18729 , \18428_18730 , \18429_18731 , \18430_18732 , \18431_18733 , \18432_18734 , \18433_18735 , \18434_18736 , \18435_18737 , \18436_18738 ,
         \18437_18739 , \18438_18740 , \18439_18741 , \18440_18742 , \18441_18743 , \18442_18744 , \18443_18745 , \18444_18746 , \18445_18747 , \18446_18748 ,
         \18447_18749 , \18448_18750 , \18449_18751 , \18450_18752 , \18451_18753 , \18452_18754 , \18453_18755 , \18454_18756 , \18455_18757 , \18456_18758 ,
         \18457_18759 , \18458_18760 , \18459_18761 , \18460_18762 , \18461_18763 , \18462_18764 , \18463_18765 , \18464_18766 , \18465_18767 , \18466_18768 ,
         \18467_18769 , \18468_18770 , \18469_18771 , \18470_18772 , \18471_18773 , \18472_18774 , \18473_18775 , \18474_18776 , \18475_18777 , \18476_18778 ,
         \18477_18779 , \18478_18780 , \18479_18781 , \18480_18782 , \18481_18783 , \18482_18784 , \18483_18785 , \18484_18786 , \18485_18787 , \18486_18788 ,
         \18487_18789 , \18488_18790 , \18489_18791 , \18490_18792 , \18491_18793 , \18492_18794 , \18493_18795 , \18494_18796 , \18495_18797 , \18496_18798 ,
         \18497_18799 , \18498_18800 , \18499_18801 , \18500_18802 , \18501_18803 , \18502_18804 , \18503_18805 , \18504_18806 , \18505_18807 , \18506_18808 ,
         \18507_18809 , \18508_18810 , \18509_18811 , \18510_18812 , \18511_18813 , \18512_18814 , \18513_18815 , \18514_18816 , \18515_18817 , \18516_18818 ,
         \18517_18819 , \18518_18820 , \18519_18821 , \18520_18822 , \18521_18823 , \18522_18824 , \18523_18825 , \18524_18826 , \18525_18827 , \18526_18828 ,
         \18527_18829 , \18528_18830 , \18529_18831 , \18530_18832 , \18531_18833 , \18532_18834 , \18533_18835 , \18534_18836 , \18535_18837 , \18536_18838 ,
         \18537_18839 , \18538_18840 , \18539_18841 , \18540_18842 , \18541_18843 , \18542_18844 , \18543_18845 , \18544_18846 , \18545_18847 , \18546_18848 ,
         \18547_18849 , \18548_18850 , \18549_18851 , \18550_18852 , \18551_18853 , \18552_18854 , \18553_18855 , \18554_18856 , \18555_18857 , \18556_18858 ,
         \18557_18859 , \18558_18860 , \18559_18861 , \18560_18862 , \18561_18863 , \18562_18864 , \18563_18865 , \18564_18866 , \18565_18867 , \18566_18868 ,
         \18567_18869 , \18568_18870 , \18569_18871 , \18570_18872 , \18571_18873 , \18572_18874 , \18573_18875 , \18574_18876 , \18575_18877 , \18576_18878 ,
         \18577_18879 , \18578_18880 , \18579_18881 , \18580_18882 , \18581_18883 , \18582_18884 , \18583_18885 , \18584_18886 , \18585_18887 , \18586_18888 ,
         \18587_18889 , \18588_18890 , \18589_18891 , \18590_18892 , \18591_18893 , \18592_18894 , \18593_18895 , \18594_18896 , \18595_18897 , \18596 ,
         \18597_18899 , \18598_18900 , \18599_18901 , \18600_18902 , \18601_18903 , \18602_18904 , \18603_18905 , \18604_18906 , \18605_18907 , \18606_18908 ,
         \18607_18909 , \18608_18910 , \18609_18911 , \18610_18912 , \18611_18913 , \18612_18914 , \18613_18915 , \18614_18916 , \18615_18917 , \18616_18918 ,
         \18617_18919 , \18618_18920 , \18619_18921 , \18620_18922 , \18621_18923 , \18622_18924 , \18623_18925 , \18624_18926 , \18625_18927 , \18626_18928 ,
         \18627_18929 , \18628_18930 , \18629_18931 , \18630_18932 , \18631_18933 , \18632_18934 , \18633_18935 , \18634_18936 , \18635_18937 , \18636_18938 ,
         \18637_18939 , \18638_18940 , \18639_18941 , \18640_18942 , \18641_18943 , \18642_18944 , \18643_18945 , \18644_18946 , \18645_18947 , \18646_18948 ,
         \18647_18949 , \18648_18950 , \18649_18951 , \18650_18952 , \18651_18953 , \18652_18954 , \18653_18955 , \18654_18956 , \18655_18957 , \18656_18958 ,
         \18657_18959 , \18658_18960 , \18659_18961 , \18660_18962 , \18661_18963 , \18662_18964 , \18663_18965 , \18664_18966 , \18665_18967 , \18666_18968 ,
         \18667_18969 , \18668_18970 , \18669_18971 , \18670_18972 , \18671_18973 , \18672_18974 , \18673_18975 , \18674_18976 , \18675_18977 , \18676_18978 ,
         \18677_18979 , \18678_18980 , \18679_18981 , \18680_18982 , \18681_18983 , \18682_18984 , \18683_18985 , \18684_18986 , \18685_18987 , \18686_18988 ,
         \18687_18989 , \18688_18990 , \18689_18991 , \18690_18992 , \18691_18993 , \18692_18994 , \18693_18995 , \18694_18996 , \18695_18997 , \18696_18998 ,
         \18697_18999 , \18698_19000 , \18699_19001 , \18700_19002 , \18701_19003 , \18702_19004 , \18703_19005 , \18704_19006 , \18705_19007 , \18706_19008 ,
         \18707_19009 , \18708_19010 , \18709_19011 , \18710_19012 , \18711_19013 , \18712_19014 , \18713_19015 , \18714_19016 , \18715_19017 , \18716_19018 ,
         \18717_19019 , \18718_19020 , \18719_19021 , \18720_19022 , \18721_19023 , \18722_19024 , \18723_19025 , \18724_19026 , \18725_19027 , \18726_19028 ,
         \18727_19029 , \18728 , \18729_19031_nG65a3 , \18730_19032 , \18731_19033 , \18732_19034 , \18733_19035 , \18734_19036 , \18735_19037 , \18736_19038 ,
         \18737_19039 , \18738_19040 , \18739 , \18740 , \18741_19043_nG53dd , \18742_19044 , \18743_19045 , \18744_19046 , \18745_19047 , \18746_19048 ,
         \18747_19049 , \18748_19050 , \18749_19051 , \18750_19052 , \18751_19053 , \18752_19054 , \18753_19055 , \18754_19056 , \18755_19057 , \18756_19058 ,
         \18757_19059 , \18758_19060 , \18759_19061 , \18760_19062 , \18761_19063 , \18762_19064 , \18763_19065 , \18764_19066 , \18765_19067 , \18766_19068 ,
         \18767_19069 , \18768_19070 , \18769_19071 , \18770_19072 , \18771_19073 , \18772_19074 , \18773_19075 , \18774_19076 , \18775_19077 , \18776_19078 ,
         \18777_19079 , \18778_19080 , \18779_19081 , \18780_19082 , \18781_19083 , \18782_19084 , \18783_19085 , \18784_19086 , \18785_19087 , \18786_19088 ,
         \18787_19089 , \18788_19090 , \18789_19091_nG9be4 , \18790_19092 , \18791_19093 , \18792_19094 , \18793_19095 , \18794_19096 , \18795_19097 , \18796_19098 ,
         \18797_19099 , \18798_19100 , \18799_19101 , \18800_19102 , \18801_19103 , \18802_19104 , \18803_19105 , \18804_19106 , \18805_19107 , \18806_19108 ,
         \18807_19109 , \18808_19110 , \18809_19111 , \18810_19112 , \18811_19113 , \18812_19114 , \18813_19115 , \18814_19116 , \18815_19117 , \18816_19118 ,
         \18817_19119 , \18818_19120 , \18819_19121 , \18820_19122 , \18821_19123 , \18822_19124 , \18823_19125 , \18824_19126 , \18825_19127 , \18826_19128 ,
         \18827_19129 , \18828_19130 , \18829_19131 , \18830_19132 , \18831_19133 , \18832_19134 , \18833_19135 , \18834_19136 , \18835_19137 , \18836_19138 ,
         \18837_19139 , \18838_19140 , \18839_19141 , \18840_19142 , \18841_19143 , \18842_19144 , \18843_19145 , \18844_19146 , \18845_19147 , \18846_19148 ,
         \18847_19149 , \18848_19150 , \18849_19151 , \18850_19152 , \18851_19153 , \18852_19154 , \18853_19155 , \18854_19156 , \18855_19157 , \18856_19158 ,
         \18857_19159 , \18858_19160 , \18859_19161 , \18860_19162 , \18861_19163 , \18862_19164 , \18863_19165 , \18864_19166 , \18865_19167 , \18866_19168 ,
         \18867_19169 , \18868_19170 , \18869_19171 , \18870_19172 , \18871_19173 , \18872_19174 , \18873_19175 , \18874_19176 , \18875_19177 , \18876_19178 ,
         \18877_19179 , \18878_19180 , \18879_19181 , \18880_19182 , \18881_19183 , \18882_19184 , \18883_19185 , \18884_19186 , \18885_19187 , \18886_19188 ,
         \18887_19189 , \18888_19190 , \18889_19191 , \18890_19192 , \18891_19193 , \18892_19194 , \18893_19195 , \18894_19196 , \18895_19197 , \18896_19198 ,
         \18897_19199 , \18898_19200 , \18899_19201 , \18900_19202 , \18901_19203 , \18902_19204 , \18903_19205 , \18904_19206 , \18905_19207 , \18906_18700 ,
         \18907_18701 , \18908_18702 , \18909_19208 , \18910_19209 , \18911_19210 , \18912_19211 , \18913_19212 , \18914_19213 , \18915_19214 , \18916_19215 ,
         \18917_19216 , \18918_19217 , \18919_19218 , \18920_19219 , \18921_19220 , \18922_19221 , \18923_19222 , \18924_19223 , \18925_19224 , \18926_19225 ,
         \18927_19226 , \18928_19227 , \18929_19228 , \18930_19229 , \18931_19230 , \18932_19231 , \18933_19232 , \18934_19233 , \18935_19234 , \18936_19235 ,
         \18937_19236 , \18938_19237 , \18939_19238 , \18940_19239 , \18941_19240 , \18942_19241 , \18943_19242 , \18944_19243 , \18945_19244 , \18946_19245 ,
         \18947_19246 , \18948_19247 , \18949_19248 , \18950_19249 , \18951_19250 , \18952_19251 , \18953_19252 , \18954_19253 , \18955_19254 , \18956_19255 ,
         \18957_19256 , \18958_19257 , \18959_19258 , \18960_19259 , \18961_19260 , \18962_19261 , \18963_19262 , \18964_19263 , \18965_19264 , \18966_19265 ,
         \18967_19266 , \18968_19267 , \18969_19268 , \18970_19269 , \18971_19270 , \18972_19271 , \18973_19272 , \18974_19273 , \18975_19274 , \18976_19275 ,
         \18977_19276 , \18978_19277 , \18979_19278 , \18980_19279 , \18981_19280 , \18982_19281 , \18983_19282 , \18984_19283 , \18985_19284 , \18986_19285 ,
         \18987_19286 , \18988_19287 , \18989_19288 , \18990_19289 , \18991_19290 , \18992_19291 , \18993_19292 , \18994_19293 , \18995_19294 , \18996_19295 ,
         \18997_19296 , \18998_19297 , \18999_19298 , \19000_19299 , \19001_19300 , \19002_19301 , \19003_19302 , \19004_19303 , \19005_19304 , \19006_19305 ,
         \19007_19306 , \19008_19307 , \19009_19308 , \19010_19309 , \19011_19310 , \19012_19311 , \19013_19312 , \19014_19313 , \19015_19314 , \19016_19315 ,
         \19017_19316 , \19018_19317 , \19019_19318 , \19020_19319 , \19021_19320 , \19022_19321 , \19023_19322 , \19024_19323 , \19025_19324 , \19026_19325 ,
         \19027_19326 , \19028_19327 , \19029_19328 , \19030_19329 , \19031_19330 , \19032_19331 , \19033_19332 , \19034_19333 , \19035_19334 , \19036_19335 ,
         \19037_19336 , \19038_19337 , \19039_19338 , \19040_19339 , \19041_19340 , \19042_19341 , \19043_19342 , \19044_19343 , \19045_19344 , \19046_19345 ,
         \19047_19346 , \19048_19347 , \19049_19348 , \19050_19349 , \19051_19350 , \19052_19351 , \19053_19352 , \19054_19353 , \19055_19354 , \19056_19355 ,
         \19057_19356 , \19058_19357 , \19059_19358 , \19060_19359 , \19061_19360 , \19062_19361 , \19063_19362 , \19064_19363 , \19065_19364 , \19066_19365 ,
         \19067_19366 , \19068_19367 , \19069_19368 , \19070_19369 , \19071_19370 , \19072_19371 , \19073_19372 , \19074_19373 , \19075_19374 , \19076_19375 ,
         \19077_19376 , \19078_19377 , \19079_19378 , \19080_19379 , \19081_19380 , \19082_19381 , \19083_19382 , \19084_19383 , \19085_19384 , \19086_19385 ,
         \19087_19386 , \19088_19387 , \19089_19388 , \19090_19389 , \19091_19390 , \19092_19391 , \19093_19392 , \19094_19393 , \19095_19394 , \19096_19395 ,
         \19097_19396 , \19098 , \19099_19398 , \19100_19399 , \19101_19400 , \19102_19401 , \19103_19402 , \19104_19403 , \19105_19404 , \19106_19405 ,
         \19107_19406 , \19108_19407 , \19109_19408 , \19110_19409 , \19111_19410 , \19112_19411 , \19113_19412 , \19114_19413 , \19115_19414 , \19116_19415 ,
         \19117_19416 , \19118_19417 , \19119_19418 , \19120_19419 , \19121_19420 , \19122_19421 , \19123_19422 , \19124_19423 , \19125_19424 , \19126_19425 ,
         \19127_19426 , \19128_19427 , \19129_19428 , \19130_19429 , \19131_19430 , \19132_19431 , \19133_19432 , \19134_19433 , \19135_19434 , \19136_19435 ,
         \19137_19436 , \19138_19437 , \19139_19438 , \19140_19439 , \19141_19440 , \19142_19441 , \19143_19442 , \19144_19443 , \19145_19444 , \19146_19445 ,
         \19147_19446 , \19148_19447 , \19149_19448 , \19150_19449 , \19151_19450 , \19152_19451 , \19153_19452 , \19154_19453 , \19155_19454 , \19156_19455 ,
         \19157_19456 , \19158_19457 , \19159_19458 , \19160_19459 , \19161_19460 , \19162_19461 , \19163_19462 , \19164_19463 , \19165_19464 , \19166_19465 ,
         \19167_19466 , \19168_19467 , \19169_19468 , \19170_19469 , \19171_19470 , \19172_19471 , \19173_19472 , \19174_19473 , \19175_19474 , \19176_19475 ,
         \19177_19476 , \19178_19477 , \19179_19478 , \19180_19479 , \19181_19480 , \19182_19481 , \19183_19482 , \19184_19483 , \19185_19484 , \19186_19485 ,
         \19187_19486 , \19188_19487 , \19189_19488 , \19190_19489 , \19191_19490 , \19192_19491 , \19193_19492 , \19194_19493 , \19195_19494 , \19196_19495 ,
         \19197_19496 , \19198_19497 , \19199_19498 , \19200_19499 , \19201_19500 , \19202_19501 , \19203_19502 , \19204_19503 , \19205_19504 , \19206_19505 ,
         \19207_19506 , \19208_19507 , \19209_19508 , \19210_19509 , \19211_19510 , \19212_19511 , \19213_19512 , \19214_19513 , \19215_19514 , \19216_19515 ,
         \19217_19516 , \19218_19517 , \19219_19518 , \19220_19519 , \19221_19520 , \19222_19521 , \19223_19522 , \19224_19523 , \19225_19524 , \19226_19525 ,
         \19227_19526 , \19228_19527 , \19229_19528 , \19230 , \19231_19530_nG54e6 , \19232_19531 , \19233_19532 , \19234_19533 , \19235_19534 , \19236_19535 ,
         \19237_19536 , \19238_19537 , \19239_19538 , \19240_19539 , \19241_19540 , \19242_19541 , \19243_19542 , \19244_19543 , \19245_19544 , \19246_19545 ,
         \19247_19546 , \19248_19547 , \19249_19548 , \19250_19549 , \19251_19550 , \19252_19551 , \19253_19552 , \19254_19553 , \19255_19554 , \19256 ,
         \19257 , \19258_19557_nG65a6 , \19259_19558 , \19260_19559 , \19261_19560 , \19262_19561 , \19263_19562 , \19264_19563 , \19265_19564 , \19266_19565 ,
         \19267_19566 , \19268_19567 , \19269_19568 , \19270_19569 , \19271_19570 , \19272_19571 , \19273_19572 , \19274_19573 , \19275_19574 , \19276_19575 ,
         \19277_19576 , \19278_19577 , \19279_19578 , \19280_19579 , \19281_19580 , \19282_19581 , \19283_19582 , \19284_19583 , \19285_19584 , \19286_19585 ,
         \19287_19586_nG9be1 , \19288_19587 , \19289_19588 , \19290_19589 , \19291_19590 , \19292_19591 , \19293_19592 , \19294_19593 , \19295_19594 , \19296_19595 ,
         \19297_19596 , \19298_19597 , \19299_19598 , \19300_19599 , \19301_19600 , \19302_19601 , \19303_19602 , \19304_19603 , \19305_19604 , \19306_19605 ,
         \19307_19606 , \19308_19607 , \19309_19608 , \19310_19609 , \19311_19610 , \19312_19611 , \19313_19612 , \19314_19613 , \19315_19614 , \19316_19615 ,
         \19317_19616 , \19318_19617 , \19319_19618 , \19320_19619 , \19321_19620 , \19322_19621 , \19323_19622 , \19324_19623 , \19325_19624 , \19326_19625 ,
         \19327_19626 , \19328_19627 , \19329_19628 , \19330_19629 , \19331_19630 , \19332_19631 , \19333_19632 , \19334_19633 , \19335_19634 , \19336_19635 ,
         \19337_19636 , \19338_19637 , \19339_19638 , \19340_19639 , \19341_19640 , \19342_19641 , \19343_19642 , \19344_19643 , \19345_19644 , \19346_19645 ,
         \19347_19646 , \19348_19647 , \19349_19648 , \19350_19649 , \19351_19650 , \19352_19651 , \19353_19652 , \19354_19653 , \19355_19654 , \19356_19655 ,
         \19357_19656 , \19358_19657 , \19359_19658 , \19360_19659 , \19361_19660 , \19362_19661 , \19363_19662 , \19364_19663 , \19365_19664 , \19366_19665 ,
         \19367_19666 , \19368_19667 , \19369_19668 , \19370_19669 , \19371_19670 , \19372_19671 , \19373_19672 , \19374_19673 , \19375_19674 , \19376_19675 ,
         \19377_19676 , \19378_19677 , \19379_19678 , \19380_19679 , \19381_19680 , \19382_19681 , \19383_19682 , \19384_19683 , \19385_19684 , \19386_19685 ,
         \19387_19686 , \19388_19687 , \19389_19688 , \19390_19689 , \19391_19690 , \19392_19691 , \19393_19692 , \19394_19693 , \19395_19694 , \19396_19695 ,
         \19397_19696 , \19398_19697 , \19399_19698 , \19400_19699 , \19401_19700 , \19402_19701 , \19403_19702 , \19404_19703 , \19405_19704 , \19406_19705 ,
         \19407_19706 , \19408_19707 , \19409_19708 , \19410_19709 , \19411_19710 , \19412_19711 , \19413_19712 , \19414_19713 , \19415_19714 , \19416_19715 ,
         \19417_19716 , \19418_19717 , \19419_19718 , \19420_19719 , \19421_19720 , \19422_19721 , \19423_19722 , \19424_19723 , \19425_19724 , \19426_19725 ,
         \19427_19726 , \19428_19727 , \19429_19728 , \19430_19729 , \19431_19730 , \19432_19731 , \19433_19732 , \19434_19733 , \19435_19734 , \19436 ,
         \19437_19736 , \19438_19737 , \19439_19738 , \19440_19739 , \19441_19740 , \19442_19741 , \19443_19742 , \19444_19743 , \19445_19744 , \19446_19745 ,
         \19447_19746 , \19448_19747 , \19449_19748 , \19450_19749 , \19451_19750 , \19452_19751 , \19453_19752 , \19454_19753 , \19455_19754 , \19456_19755 ,
         \19457_19756 , \19458_19757 , \19459_19758 , \19460_19759 , \19461_19760 , \19462_19761 , \19463_19762 , \19464_19763 , \19465_19764 , \19466_19765 ,
         \19467_19766 , \19468_19767 , \19469_19768 , \19470_19769 , \19471_19770 , \19472_19771 , \19473_19772 , \19474_19773 , \19475_19774 , \19476_19775 ,
         \19477_19776 , \19478_19777 , \19479_19778 , \19480_19779 , \19481_19780 , \19482_19781 , \19483_19782 , \19484_19783 , \19485_19784 , \19486_19785 ,
         \19487_19786 , \19488_19787 , \19489_19788 , \19490_19789 , \19491_19790 , \19492_19791 , \19493_19792 , \19494_19793 , \19495_19794 , \19496_19795 ,
         \19497_19796 , \19498_19797 , \19499_19798 , \19500_19799 , \19501_19800 , \19502_19801 , \19503_19802 , \19504_19803 , \19505_19804 , \19506_19805 ,
         \19507_19806 , \19508_19807 , \19509_19808 , \19510_19809 , \19511_19810 , \19512_19811 , \19513_19812 , \19514_19813 , \19515_19814 , \19516_19815 ,
         \19517_19816 , \19518_19817 , \19519_19818 , \19520_19819 , \19521_19820 , \19522_19821 , \19523_19822 , \19524_19823 , \19525_19824 , \19526_19825 ,
         \19527_19826 , \19528_19827 , \19529_19828 , \19530_19829 , \19531_19830 , \19532_19831 , \19533_19832 , \19534_19833 , \19535_19834 , \19536_19835 ,
         \19537_19836 , \19538_19837 , \19539_19838 , \19540_19839 , \19541_19840 , \19542_19841 , \19543_19842 , \19544_19843 , \19545_19844 , \19546_19845 ,
         \19547_19846 , \19548_19847 , \19549_19848 , \19550_19849 , \19551_19850 , \19552_19851 , \19553_19852 , \19554_19853 , \19555_19854 , \19556_19855 ,
         \19557_19856 , \19558_19857 , \19559_19858 , \19560_19859 , \19561_19860 , \19562_19861 , \19563_19862 , \19564_19863 , \19565_19864 , \19566_19865 ,
         \19567_19866 , \19568_19867 , \19569 , \19570_19869 , \19571_19870 , \19572_19871 , \19573_19872 , \19574_19873 , \19575_19874 , \19576_19875 ,
         \19577_19876 , \19578_19877 , \19579_19878 , \19580_19879 , \19581_19880 , \19582_19881 , \19583_19882 , \19584_19883 , \19585_19884 , \19586_19885 ,
         \19587_19886 , \19588_19887 , \19589_19888 , \19590_19889 , \19591_19890 , \19592_19891 , \19593_19892 , \19594_19893 , \19595_19894 , \19596_19895 ,
         \19597_19896 , \19598_19897 , \19599_19898 , \19600_19899 , \19601_19900 , \19602_19901 , \19603_19902 , \19604_19903 , \19605_19904 , \19606_19905 ,
         \19607_19906 , \19608_19907 , \19609_19908 , \19610_19909 , \19611_19910 , \19612_19911 , \19613_19912 , \19614_19913 , \19615_19914 , \19616_19915 ,
         \19617_19916 , \19618_19917 , \19619_19918 , \19620_19919 , \19621_19920 , \19622_19921 , \19623_19922 , \19624_19923 , \19625_19924 , \19626_19925 ,
         \19627_19926 , \19628_19927 , \19629_19928 , \19630_19929 , \19631_19930 , \19632_19931 , \19633_19932 , \19634_19933 , \19635_19934 , \19636_19935 ,
         \19637_19936 , \19638_19937 , \19639_19938 , \19640_19939 , \19641_19940 , \19642_19941 , \19643_19942 , \19644_19943 , \19645_19944 , \19646_19945 ,
         \19647_19946 , \19648_19947 , \19649_19948 , \19650_19949 , \19651_19950 , \19652_19951 , \19653_19952 , \19654_19953 , \19655_19954 , \19656_19955 ,
         \19657_19956 , \19658_19957 , \19659_19958 , \19660_19959 , \19661_19960 , \19662_19961 , \19663_19962 , \19664_19963 , \19665_19964 , \19666_19965 ,
         \19667_19966 , \19668_19967 , \19669_19968 , \19670_19969 , \19671_19970 , \19672_19971 , \19673_19972 , \19674_19973 , \19675_19974 , \19676_19975 ,
         \19677_19976 , \19678_19977 , \19679_19978 , \19680_19979 , \19681_19980 , \19682_19981 , \19683_19982 , \19684_19983 , \19685_19984 , \19686_19985 ,
         \19687_19986 , \19688_19987 , \19689_19988 , \19690_19989 , \19691_19990 , \19692_19991 , \19693_19992 , \19694_19993 , \19695_19994 , \19696_19995 ,
         \19697_19996 , \19698_19997 , \19699_19998 , \19700_19999 , \19701_20000 , \19702_20001 , \19703 , \19704_20003 , \19705_20004 , \19706_20005 ,
         \19707_20006 , \19708_20007 , \19709_20008 , \19710_20009 , \19711_20010 , \19712_20011 , \19713_20012 , \19714_20013 , \19715_20014 , \19716_20015 ,
         \19717_20016 , \19718_20017 , \19719_20018 , \19720_20019 , \19721_20020 , \19722_20021 , \19723_20022 , \19724_20023 , \19725_20024 , \19726_20025 ,
         \19727_20026 , \19728_20027 , \19729_20028 , \19730_20029 , \19731_20030 , \19732_20031 , \19733_20032 , \19734_20033 , \19735_20034 , \19736_20035 ,
         \19737_20036 , \19738_20037 , \19739_20038 , \19740_20039 , \19741_20040 , \19742_20041 , \19743_20042 , \19744_20043 , \19745_20044 , \19746_20045 ,
         \19747_20046 , \19748_20047 , \19749_20048 , \19750_20049 , \19751_20050 , \19752_20051 , \19753_20052 , \19754_20053 , \19755_20054 , \19756_20055 ,
         \19757_20056 , \19758_20057 , \19759_20058 , \19760_20059 , \19761_20060 , \19762_20061 , \19763_20062 , \19764_20063 , \19765_20064 , \19766_20065 ,
         \19767_20066 , \19768_20067 , \19769_20068 , \19770_20069 , \19771_20070 , \19772_20071 , \19773_20072 , \19774_20073 , \19775_20074 , \19776_20075 ,
         \19777_20076 , \19778_20077 , \19779_20078 , \19780_20079 , \19781_20080 , \19782_20081 , \19783_20082 , \19784_20083 , \19785_20084 , \19786_20085 ,
         \19787_20086 , \19788_20087 , \19789_20088 , \19790_20089 , \19791_20090 , \19792_20091 , \19793_20092 , \19794_20093 , \19795_20094 , \19796_20095 ,
         \19797_20096 , \19798_20097 , \19799_20098 , \19800_20099 , \19801_20100 , \19802_20101 , \19803_20102 , \19804_20103 , \19805_20104 , \19806_20105 ,
         \19807_20106 , \19808_20107 , \19809_20108 , \19810_20109 , \19811_20110 , \19812_20111 , \19813_20112 , \19814_20113 , \19815_20114 , \19816_20115 ,
         \19817_20116 , \19818_20117 , \19819_20118 , \19820_20119 , \19821_20120 , \19822_20121 , \19823_20122 , \19824_20123 , \19825_20124 , \19826_20125 ,
         \19827_20126 , \19828_20127 , \19829_20128 , \19830_20129 , \19831_20130 , \19832_20131 , \19833_20132 , \19834_20133 , \19835_20134 , \19836 ,
         \19837_20136 , \19838_20137 , \19839_20138 , \19840_20139 , \19841_20140 , \19842_20141 , \19843_20142 , \19844_20143 , \19845_20144 , \19846_20145 ,
         \19847_20146_nG4424 , \19848_20147 , \19849_20148 , \19850_20149_nG4427 , \19851_20150 , \19852_20151 , \19853_20152 , \19854_20156 , \19855_20157 , \19856_20158 ,
         \19857_20159 , \19858_20160 , \19859_20161 , \19860_20162 , \19861_20163 , \19862_20164 , \19863_20165 , \19864_20166 , \19865_20167 , \19866_20168 ,
         \19867_20169 , \19868_20170 , \19869_20171 , \19870_20172 , \19871_20173 , \19872_20174 , \19873_20175 , \19874_20176 , \19875_20177 , \19876_20178 ,
         \19877_20179 , \19878_20180 , \19879_20181 , \19880_20182 , \19881_20183 , \19882_20184 , \19883_20185 , \19884_20186 , \19885_20187 , \19886_20188 ,
         \19887_20189 , \19888_20190 , \19889_20191 , \19890_20192 , \19891_20193 , \19892_20194 , \19893_20195 , \19894_20196 , \19895_20197 , \19896_20198 ,
         \19897_20199 , \19898_20200 , \19899_20201 , \19900_20202 , \19901_20203 , \19902_20204 , \19903_20205 , \19904_20206 , \19905_20207 , \19906_20208 ,
         \19907_20209 , \19908_20210 , \19909_20211 , \19910_20212 , \19911_20213 , \19912_20214 , \19913_20215 , \19914_20216 , \19915_20217 , \19916_20218 ,
         \19917_20219 , \19918_20220 , \19919_20221 , \19920_20222 , \19921_20223 , \19922_20224 , \19923_20225 , \19924_20226 , \19925_20227 , \19926_20228 ,
         \19927_20229 , \19928_20230 , \19929_20231 , \19930_20232 , \19931_20233 , \19932_20234 , \19933_20235 , \19934_20236 , \19935_20237 , \19936_20238 ,
         \19937_20239 , \19938_20240 , \19939_20241 , \19940_20242 , \19941_20243 , \19942_20244 , \19943_20245 , \19944_20246 , \19945_20247 , \19946_20248 ,
         \19947_20249 , \19948_20250 , \19949_20251 , \19950_20252 , \19951_20253 , \19952_20254 , \19953_20255 , \19954_20256 , \19955_20257 , \19956_20258 ,
         \19957_20259 , \19958_20260 , \19959_20261 , \19960_20262 , \19961_20263 , \19962_20264 , \19963_20265 , \19964_20266 , \19965_20267 , \19966_20268 ,
         \19967_20269 , \19968_20270 , \19969_20271 , \19970_20272 , \19971_20273 , \19972_20274 , \19973_20275 , \19974_20276 , \19975_20277 , \19976_20278 ,
         \19977_20279 , \19978_20280 , \19979_20281 , \19980_20282 , \19981_20283 , \19982_20284 , \19983_20285 , \19984_20286 , \19985_20287 , \19986_20288 ,
         \19987_20289 , \19988_20290 , \19989_20291 , \19990_20292 , \19991_20293 , \19992_20294 , \19993_20295 , \19994_20296 , \19995_20297 , \19996_20298 ,
         \19997_20299 , \19998_20300 , \19999_20301 , \20000_20302 , \20001_20303 , \20002_20304 , \20003_20305 , \20004_20306 , \20005_20307 , \20006_20308 ,
         \20007_20309 , \20008_20310 , \20009_20311 , \20010_20312 , \20011_20313 , \20012_20314 , \20013_20315 , \20014_20316 , \20015_20317 , \20016_20318 ,
         \20017_20319 , \20018_20320 , \20019_20321 , \20020_20322 , \20021_20323 , \20022_20324 , \20023_20325 , \20024_20326 , \20025_20327 , \20026_20328 ,
         \20027_20329 , \20028_20330 , \20029_20331 , \20030_20332 , \20031_20333 , \20032_20334 , \20033_20335 , \20034_20336 , \20035_20337 , \20036_20338 ,
         \20037_20339 , \20038_20340 , \20039_20341 , \20040_20342 , \20041_20343 , \20042_20344 , \20043_20345 , \20044_20346 , \20045_20347 , \20046_20348 ,
         \20047_20349 , \20048_20350 , \20049_20351 , \20050_20352 , \20051_20353 , \20052_20354 , \20053_20355 , \20054_20356 , \20055_20357 , \20056_20358 ,
         \20057_20359 , \20058_20360 , \20059_20361 , \20060_20362 , \20061_20363 , \20062_20364 , \20063_20365 , \20064_20366 , \20065_20367 , \20066_20368 ,
         \20067_20369 , \20068_20370 , \20069_20371 , \20070_20372 , \20071_20373 , \20072_20374 , \20073_20375 , \20074_20376 , \20075_20377 , \20076_20378 ,
         \20077_20379 , \20078_20380 , \20079_20381 , \20080_20382 , \20081_20383 , \20082_20384 , \20083_20385 , \20084_20386 , \20085_20387 , \20086_20388 ,
         \20087_20389 , \20088_20390 , \20089_20391 , \20090_20392 , \20091_20393 , \20092_20394 , \20093_20395 , \20094_20396 , \20095_20397 , \20096_20398 ,
         \20097_20399 , \20098_20400 , \20099_20401 , \20100_20402 , \20101_20403 , \20102_20404 , \20103_20405 , \20104_20406 , \20105_20407 , \20106_20408 ,
         \20107_20409 , \20108 , \20109_20411 , \20110_20412 , \20111_20413 , \20112_20414 , \20113_20415 , \20114_20416 , \20115_20417 , \20116_20418 ,
         \20117_20419 , \20118_20420 , \20119_20421 , \20120_20422 , \20121_20423 , \20122_20424 , \20123_20425 , \20124_20426 , \20125_20427 , \20126_20428 ,
         \20127_20429 , \20128_20430 , \20129_20431 , \20130_20432 , \20131_20433 , \20132_20434 , \20133_20435 , \20134_20436 , \20135_20437 , \20136_20438 ,
         \20137_20439 , \20138_20440 , \20139_20441 , \20140_20442 , \20141_20443 , \20142_20444 , \20143_20445 , \20144_20446 , \20145_20447 , \20146_20448 ,
         \20147_20449 , \20148_20450 , \20149_20451 , \20150_20452 , \20151_20453 , \20152_20454 , \20153_20455 , \20154_20456 , \20155_20457 , \20156_20458 ,
         \20157_20459 , \20158_20460 , \20159_20461 , \20160_20462 , \20161_20463 , \20162_20464 , \20163_20465 , \20164_20466 , \20165_20467 , \20166_20468 ,
         \20167_20469 , \20168_20470 , \20169_20471 , \20170_20472 , \20171_20473 , \20172_20474 , \20173_20475 , \20174_20476 , \20175_20477 , \20176_20478 ,
         \20177_20479 , \20178_20480 , \20179_20481 , \20180_20482 , \20181_20483 , \20182_20484 , \20183_20485 , \20184_20486 , \20185_20487 , \20186_20488 ,
         \20187_20489 , \20188_20490 , \20189_20491 , \20190_20492 , \20191_20493 , \20192_20494 , \20193_20495 , \20194_20496 , \20195_20497 , \20196_20498 ,
         \20197_20499 , \20198_20500 , \20199_20501 , \20200_20502 , \20201_20503 , \20202_20504 , \20203_20505 , \20204_20506 , \20205_20507 , \20206_20508 ,
         \20207_20509 , \20208_20510 , \20209_20511 , \20210_20512 , \20211_20513 , \20212_20514 , \20213_20515 , \20214_20516 , \20215_20517 , \20216_20518 ,
         \20217_20519 , \20218_20520 , \20219_20521 , \20220_20522 , \20221_20523 , \20222_20524 , \20223_20525 , \20224_20526 , \20225_20527 , \20226_20528 ,
         \20227_20529 , \20228_20530 , \20229_20531 , \20230_20532 , \20231_20533 , \20232_20534 , \20233_20535 , \20234_20536 , \20235_20537 , \20236_20538 ,
         \20237_20539 , \20238_20540 , \20239_20541 , \20240 , \20241_20543_nG65a9 , \20242_20544 , \20243_20545 , \20244_20546 , \20245_20547 , \20246_20548 ,
         \20247_20549 , \20248_20550 , \20249_20551 , \20250_20552 , \20251 , \20252 , \20253_20555_nG55ef , \20254_20556 , \20255_20557 , \20256_20558 ,
         \20257_20559 , \20258_20560 , \20259_20561 , \20260_20562 , \20261_20563 , \20262_20564 , \20263_20565 , \20264_20566 , \20265_20567 , \20266_20568 ,
         \20267_20569 , \20268_20570 , \20269_20571 , \20270_20572 , \20271_20573 , \20272_20574 , \20273_20575 , \20274_20576 , \20275_20577 , \20276_20578 ,
         \20277_20579 , \20278_20580 , \20279_20581 , \20280_20582 , \20281_20583 , \20282_20584 , \20283_20585 , \20284_20586 , \20285_20587 , \20286_20588 ,
         \20287_20589 , \20288_20590 , \20289_20591 , \20290_20592 , \20291_20593 , \20292_20594 , \20293_20595 , \20294_20596 , \20295_20597 , \20296_20598 ,
         \20297_20599 , \20298_20600 , \20299_20601 , \20300_20602 , \20301_20603 , \20302_20604 , \20303_20605 , \20304_20606 , \20305_20607 , \20306_20608_nG9bde ,
         \20307_20609 , \20308_20610 , \20309_20611 , \20310_20612 , \20311_20613 , \20312_20614 , \20313_20615 , \20314_20616 , \20315_20617 , \20316_20618 ,
         \20317_20619 , \20318_20620 , \20319_20621 , \20320_20622 , \20321_20623 , \20322_20624 , \20323_20625 , \20324_20626 , \20325_20627 , \20326_20628 ,
         \20327_20629 , \20328_20630 , \20329_20631 , \20330_20632 , \20331_20633 , \20332_20634 , \20333_20635 , \20334_20636 , \20335_20637 , \20336_20638 ,
         \20337_20639 , \20338_20640 , \20339_20641 , \20340_20642 , \20341_20643 , \20342_20644 , \20343_20645 , \20344_20646 , \20345_20647 , \20346_20648 ,
         \20347_20649 , \20348_20650 , \20349_20651 , \20350_20652 , \20351_20153 , \20352_20154 , \20353_20155 , \20354_20653 , \20355_20654 , \20356_20655 ,
         \20357_20656 , \20358_20657 , \20359_20658 , \20360_20659 , \20361_20660 , \20362_20661 , \20363_20662 , \20364_20663 , \20365_20664 , \20366_20665 ,
         \20367_20666 , \20368_20667 , \20369_20668 , \20370_20669 , \20371_20670 , \20372_20671 , \20373_20672 , \20374_20673 , \20375_20674 , \20376_20675 ,
         \20377_20676 , \20378_20677 , \20379_20678 , \20380_20679 , \20381_20680 , \20382_20681 , \20383_20682 , \20384_20683 , \20385_20684 , \20386_20685 ,
         \20387_20686 , \20388_20687 , \20389_20688 , \20390_20689 , \20391_20690 , \20392_20691 , \20393_20692 , \20394_20693 , \20395_20694 , \20396_20695 ,
         \20397_20696 , \20398_20697 , \20399_20698 , \20400_20699 , \20401_20700 , \20402_20701 , \20403_20702 , \20404_20703 , \20405_20704 , \20406_20705 ,
         \20407_20706 , \20408_20707 , \20409_20708 , \20410_20709 , \20411_20710 , \20412_20711 , \20413_20712 , \20414_20713 , \20415_20714 , \20416_20715 ,
         \20417_20716 , \20418_20717 , \20419_20718 , \20420_20719 , \20421_20720 , \20422_20721 , \20423_20722 , \20424_20723 , \20425_20724 , \20426_20725 ,
         \20427_20726 , \20428_20727 , \20429_20728 , \20430_20729 , \20431_20730 , \20432_20731 , \20433_20732 , \20434_20733 , \20435_20734 , \20436_20735 ,
         \20437_20736 , \20438_20737 , \20439_20738 , \20440_20739 , \20441_20740 , \20442_20741 , \20443_20742 , \20444_20743 , \20445_20744 , \20446_20745 ,
         \20447_20746 , \20448_20747 , \20449_20748 , \20450_20749 , \20451_20750 , \20452_20751 , \20453_20752 , \20454_20753 , \20455_20754 , \20456_20755 ,
         \20457_20756 , \20458_20757 , \20459_20758 , \20460_20759 , \20461_20760 , \20462_20761 , \20463_20762 , \20464_20763 , \20465_20764 , \20466_20765 ,
         \20467_20766 , \20468_20767 , \20469_20768 , \20470_20769 , \20471_20770 , \20472_20771 , \20473_20772 , \20474_20773 , \20475_20774 , \20476_20775 ,
         \20477_20776 , \20478_20777 , \20479_20778 , \20480_20779 , \20481_20780 , \20482_20781 , \20483_20782 , \20484_20783 , \20485_20784 , \20486_20785 ,
         \20487_20786 , \20488_20787 , \20489_20788 , \20490_20789 , \20491_20790 , \20492_20791 , \20493_20792 , \20494_20793 , \20495_20794 , \20496_20795 ,
         \20497_20796 , \20498_20797 , \20499_20798 , \20500_20799 , \20501_20800 , \20502_20801 , \20503_20802 , \20504_20803 , \20505_20804 , \20506_20805 ,
         \20507_20806 , \20508_20807 , \20509_20808 , \20510_20809 , \20511_20810 , \20512_20811 , \20513_20812 , \20514_20813 , \20515_20814 , \20516_20815 ,
         \20517_20816 , \20518_20817 , \20519_20818 , \20520_20819 , \20521_20820 , \20522_20821 , \20523_20822 , \20524_20823 , \20525_20824 , \20526_20825 ,
         \20527_20826 , \20528_20827 , \20529_20828 , \20530_20829 , \20531_20830 , \20532_20831 , \20533_20832 , \20534_20833 , \20535_20834 , \20536_20835 ,
         \20537_20836 , \20538_20837 , \20539_20838 , \20540_20839 , \20541_20840 , \20542_20841 , \20543_20842 , \20544_20843 , \20545_20844 , \20546_20845 ,
         \20547_20846 , \20548_20847 , \20549_20848 , \20550_20849 , \20551_20850 , \20552_20851 , \20553_20852 , \20554_20853 , \20555_20854 , \20556_20855 ,
         \20557_20856 , \20558_20857 , \20559_20858 , \20560_20859 , \20561_20860 , \20562_20861 , \20563_20862 , \20564_20863 , \20565_20864 , \20566_20865 ,
         \20567_20866 , \20568_20867 , \20569 , \20570_20869 , \20571_20870 , \20572_20871 , \20573_20872 , \20574_20873 , \20575_20874 , \20576_20875 ,
         \20577_20876 , \20578_20877 , \20579_20878 , \20580_20879 , \20581_20880 , \20582_20881 , \20583_20882 , \20584_20883 , \20585_20884 , \20586_20885 ,
         \20587_20886 , \20588_20887 , \20589_20888 , \20590_20889 , \20591_20890 , \20592_20891 , \20593_20892 , \20594_20893 , \20595_20894 , \20596_20895 ,
         \20597_20896 , \20598_20897 , \20599_20898 , \20600_20899 , \20601_20900 , \20602_20901 , \20603_20902 , \20604_20903 , \20605_20904 , \20606_20905 ,
         \20607_20906 , \20608_20907 , \20609_20908 , \20610_20909 , \20611_20910 , \20612_20911 , \20613_20912 , \20614_20913 , \20615_20914 , \20616_20915 ,
         \20617_20916 , \20618_20917 , \20619_20918 , \20620_20919 , \20621_20920 , \20622_20921 , \20623_20922 , \20624_20923 , \20625_20924 , \20626_20925 ,
         \20627_20926 , \20628_20927 , \20629_20928 , \20630_20929 , \20631_20930 , \20632_20931 , \20633_20932 , \20634_20933 , \20635_20934 , \20636_20935 ,
         \20637_20936 , \20638_20937 , \20639_20938 , \20640_20939 , \20641_20940 , \20642_20941 , \20643_20942 , \20644_20943 , \20645_20944 , \20646_20945 ,
         \20647_20946 , \20648_20947 , \20649_20948 , \20650_20949 , \20651_20950 , \20652_20951 , \20653_20952 , \20654_20953 , \20655_20954 , \20656_20955 ,
         \20657_20956 , \20658_20957 , \20659_20958 , \20660_20959 , \20661_20960 , \20662_20961 , \20663_20962 , \20664_20963 , \20665_20964 , \20666_20965 ,
         \20667_20966 , \20668_20967 , \20669_20968 , \20670_20969 , \20671_20970 , \20672_20971 , \20673_20972 , \20674_20973 , \20675_20974 , \20676_20975 ,
         \20677_20976 , \20678_20977 , \20679_20978 , \20680_20979 , \20681_20980 , \20682_20981 , \20683_20982 , \20684_20983 , \20685_20984 , \20686_20985 ,
         \20687_20986 , \20688_20987 , \20689_20988 , \20690_20989 , \20691_20990 , \20692_20991 , \20693_20992 , \20694_20993 , \20695_20994 , \20696_20995 ,
         \20697_20996 , \20698_20997 , \20699_20998 , \20700_20999 , \20701 , \20702_21001_nG56f8 , \20703_21002 , \20704_21003 , \20705_21004 , \20706_21005 ,
         \20707_21006 , \20708_21007 , \20709_21008 , \20710_21009 , \20711_21010 , \20712_21011 , \20713_21012 , \20714_21013 , \20715_21014 , \20716_21015 ,
         \20717_21016 , \20718_21017 , \20719_21018 , \20720_21019 , \20721_21020 , \20722_21021 , \20723_21022 , \20724_21023 , \20725_21024 , \20726_21025 ,
         \20727_21026 , \20728_21027 , \20729_21028 , \20730_21029 , \20731 , \20732 , \20733_21032_nG65ac , \20734_21033 , \20735_21034 , \20736_21035 ,
         \20737_21036 , \20738_21037 , \20739_21038 , \20740_21039 , \20741_21040 , \20742_21041 , \20743_21042 , \20744_21043 , \20745_21044 , \20746_21045 ,
         \20747_21046 , \20748_21047 , \20749_21048 , \20750_21049 , \20751_21050 , \20752_21051 , \20753_21052 , \20754_21053 , \20755_21054 , \20756_21055 ,
         \20757_21056 , \20758_21057 , \20759_21058 , \20760_21059 , \20761_21060 , \20762_21061 , \20763_21062 , \20764_21063 , \20765_21064 , \20766_21065 ,
         \20767_21066 , \20768_21067 , \20769_21068 , \20770_21069 , \20771_21070 , \20772_21071 , \20773_21072 , \20774_21073 , \20775_21074 , \20776_21075 ,
         \20777_21076 , \20778_21077 , \20779_21078 , \20780_21079 , \20781_21080 , \20782_21081 , \20783_21082 , \20784_21083 , \20785_21084 , \20786_21085 ,
         \20787_21086_nG9bdb , \20788_21087 , \20789_21088 , \20790_21089 , \20791_21090 , \20792_21091 , \20793_21092 , \20794_21093 , \20795_21094 , \20796_21095 ,
         \20797_21096 , \20798_21097 , \20799_21098 , \20800_21099 , \20801_21100 , \20802_21101 , \20803_21102 , \20804_21103 , \20805_21104 , \20806_21105 ,
         \20807_21106 , \20808_21107 , \20809_21108 , \20810_21109 , \20811_21110 , \20812_21111 , \20813_21112 , \20814_21113 , \20815_21114 , \20816_21115 ,
         \20817_21116 , \20818_21117 , \20819_21118 , \20820_21119 , \20821_21120 , \20822_21121 , \20823_21122 , \20824_21123 , \20825_21124 , \20826_21125 ,
         \20827_21126 , \20828_21127 , \20829_21128 , \20830_21129 , \20831_21130 , \20832_21131 , \20833_21132 , \20834_21133 , \20835_21134 , \20836_21135 ,
         \20837_21136 , \20838_21137 , \20839_21138 , \20840_21139 , \20841_21140 , \20842_21141 , \20843_21142 , \20844_21143 , \20845_21144 , \20846_21145 ,
         \20847_21146 , \20848_21147 , \20849_21148 , \20850_21149 , \20851_21150 , \20852_21151 , \20853_21152 , \20854_21153 , \20855_21154 , \20856_21155 ,
         \20857_21156 , \20858_21157 , \20859_21158 , \20860_21159 , \20861_21160 , \20862_21161 , \20863_21162 , \20864_21163 , \20865_21164 , \20866_21165 ,
         \20867_21166 , \20868_21167 , \20869_21168 , \20870_21169 , \20871_21170 , \20872_21171 , \20873_21172 , \20874_21173 , \20875_21174 , \20876_21175 ,
         \20877_21176 , \20878_21177 , \20879_21178 , \20880_21179 , \20881_21180 , \20882_21181 , \20883_21182 , \20884_21183 , \20885_21184 , \20886_21185 ,
         \20887_21186 , \20888_21187 , \20889_21188 , \20890_21189 , \20891_21190 , \20892_21191 , \20893_21192 , \20894_21193 , \20895_21194 , \20896_21195 ,
         \20897_21196 , \20898_21197 , \20899_21198 , \20900_21199 , \20901_21200 , \20902_21201 , \20903_21202 , \20904_21203 , \20905_21204 , \20906_21205 ,
         \20907_21206 , \20908_21207 , \20909_21208 , \20910_21209 , \20911_21210 , \20912_21211 , \20913_21212 , \20914_21213 , \20915_21214 , \20916_21215 ,
         \20917_21216 , \20918_21217 , \20919_21218 , \20920_21219 , \20921_21220 , \20922_21221 , \20923_21222 , \20924_21223 , \20925_21224 , \20926_21225 ,
         \20927_21226 , \20928_21227 , \20929_21228 , \20930_21229 , \20931_21230 , \20932_21231 , \20933_21232 , \20934_21233 , \20935_21234 , \20936_21235 ,
         \20937_21236 , \20938_21237 , \20939 , \20940_21239 , \20941_21240 , \20942_21241 , \20943_21242 , \20944_21243 , \20945_21244 , \20946_21245 ,
         \20947_21246 , \20948_21247 , \20949_21248 , \20950_21249 , \20951_21250 , \20952_21251 , \20953_21252 , \20954_21253 , \20955_21254 , \20956_21255 ,
         \20957_21256 , \20958_21257 , \20959_21258 , \20960_21259 , \20961_21260 , \20962_21261 , \20963_21262 , \20964_21263 , \20965_21264 , \20966_21265 ,
         \20967_21266 , \20968_21267 , \20969_21268 , \20970_21269 , \20971_21270 , \20972_21271 , \20973_21272 , \20974_21273 , \20975_21274 , \20976_21275 ,
         \20977_21276 , \20978_21277 , \20979_21278 , \20980_21279 , \20981_21280 , \20982_21281 , \20983_21282 , \20984_21283 , \20985_21284 , \20986_21285 ,
         \20987_21286 , \20988_21287 , \20989_21288 , \20990_21289 , \20991_21290 , \20992_21291 , \20993_21292 , \20994_21293 , \20995_21294 , \20996_21295 ,
         \20997_21296 , \20998_21297 , \20999_21298 , \21000_21299 , \21001_21300 , \21002_21301 , \21003_21302 , \21004_21303 , \21005_21304 , \21006_21305 ,
         \21007_21306 , \21008_21307 , \21009_21308 , \21010_21309 , \21011_21310 , \21012_21311 , \21013_21312 , \21014_21313 , \21015_21314 , \21016_21315 ,
         \21017_21316 , \21018_21317 , \21019_21318 , \21020_21319 , \21021_21320 , \21022_21321 , \21023_21322 , \21024_21323 , \21025_21324 , \21026_21325 ,
         \21027_21326 , \21028_21327 , \21029_21328 , \21030_21329 , \21031_21330 , \21032_21331 , \21033_21332 , \21034_21333 , \21035_21334 , \21036_21335 ,
         \21037_21336 , \21038_21337 , \21039_21338 , \21040_21339 , \21041_21340 , \21042_21341 , \21043_21342 , \21044_21343 , \21045_21344 , \21046_21345 ,
         \21047_21346 , \21048_21347 , \21049_21348 , \21050_21349 , \21051_21350 , \21052_21351 , \21053_21352 , \21054_21353 , \21055_21354 , \21056_21355 ,
         \21057_21356 , \21058_21357 , \21059_21358 , \21060_21359 , \21061_21360 , \21062_21361 , \21063_21362 , \21064_21363 , \21065_21364 , \21066_21365 ,
         \21067_21366 , \21068_21367 , \21069_21368 , \21070_21369 , \21071_21370 , \21072 , \21073_21372 , \21074_21373 , \21075_21374 , \21076_21375 ,
         \21077_21376 , \21078_21377 , \21079_21378 , \21080_21379 , \21081_21380 , \21082_21381 , \21083_21382 , \21084_21383 , \21085_21384 , \21086_21385 ,
         \21087_21386 , \21088_21387 , \21089_21388 , \21090_21389 , \21091_21390 , \21092_21391 , \21093_21392 , \21094_21393 , \21095_21394 , \21096_21395 ,
         \21097_21396 , \21098_21397 , \21099_21398 , \21100_21399 , \21101_21400 , \21102_21401 , \21103_21402 , \21104_21403 , \21105_21404 , \21106_21405 ,
         \21107_21406 , \21108_21407 , \21109_21408 , \21110_21409 , \21111_21410 , \21112_21411 , \21113_21412 , \21114_21413 , \21115_21414 , \21116_21415 ,
         \21117_21416 , \21118_21417 , \21119_21418 , \21120_21419 , \21121_21420 , \21122_21421 , \21123_21422 , \21124_21423 , \21125_21424 , \21126_21425 ,
         \21127_21426 , \21128_21427 , \21129_21428 , \21130_21429 , \21131_21430 , \21132_21431 , \21133_21432 , \21134_21433 , \21135_21434 , \21136_21435 ,
         \21137_21436 , \21138_21437 , \21139_21438 , \21140_21439 , \21141_21440 , \21142_21441 , \21143_21442 , \21144_21443 , \21145_21444 , \21146_21445 ,
         \21147_21446 , \21148_21447 , \21149_21448 , \21150_21449 , \21151_21450 , \21152_21451 , \21153_21452 , \21154_21453 , \21155_21454 , \21156_21455 ,
         \21157_21456 , \21158_21457 , \21159_21458 , \21160_21459 , \21161_21460 , \21162_21461 , \21163_21462 , \21164_21463 , \21165_21464 , \21166_21465 ,
         \21167_21466 , \21168_21467 , \21169_21468 , \21170_21469 , \21171_21470 , \21172_21471 , \21173_21472 , \21174_21473 , \21175_21474 , \21176_21475 ,
         \21177_21476 , \21178_21477 , \21179_21478 , \21180_21479 , \21181_21480 , \21182_21481 , \21183_21482 , \21184_21483 , \21185_21484 , \21186_21485 ,
         \21187_21486 , \21188_21487 , \21189_21488 , \21190_21489 , \21191_21490 , \21192_21491 , \21193_21492 , \21194_21493 , \21195_21494 , \21196_21495 ,
         \21197_21496 , \21198_21497 , \21199_21498 , \21200_21499 , \21201_21500 , \21202_21501 , \21203_21502 , \21204_21503 , \21205_21504 , \21206 ,
         \21207_21506 , \21208_21507 , \21209_21508 , \21210_21509 , \21211_21510 , \21212_21511 , \21213_21512 , \21214_21513 , \21215_21514 , \21216_21515 ,
         \21217_21516 , \21218_21517 , \21219_21518 , \21220_21519 , \21221_21520 , \21222_21521 , \21223_21522 , \21224_21523 , \21225_21524 , \21226_21525 ,
         \21227_21526 , \21228_21527 , \21229_21528 , \21230_21529 , \21231_21530 , \21232_21531 , \21233_21532 , \21234_21533 , \21235_21534 , \21236_21535 ,
         \21237_21536 , \21238_21537 , \21239_21538 , \21240_21539 , \21241_21540 , \21242_21541 , \21243_21542 , \21244_21543 , \21245_21544 , \21246_21545 ,
         \21247_21546 , \21248_21547 , \21249_21548 , \21250_21549 , \21251_21550 , \21252_21551 , \21253_21552 , \21254_21553 , \21255_21554 , \21256_21555 ,
         \21257_21556 , \21258_21557 , \21259_21558 , \21260_21559 , \21261_21560 , \21262_21561 , \21263_21562 , \21264_21563 , \21265_21564 , \21266_21565 ,
         \21267_21566 , \21268_21567 , \21269_21568 , \21270_21569 , \21271_21570 , \21272_21571 , \21273_21572 , \21274_21573 , \21275_21574 , \21276_21575 ,
         \21277_21576 , \21278_21577 , \21279_21578 , \21280_21579 , \21281_21580 , \21282_21581 , \21283_21582 , \21284_21583 , \21285_21584 , \21286_21585 ,
         \21287_21586 , \21288_21587 , \21289_21588 , \21290_21589 , \21291_21590 , \21292_21591 , \21293_21592 , \21294_21593 , \21295_21594 , \21296_21595 ,
         \21297_21596 , \21298_21597 , \21299_21598 , \21300_21599 , \21301_21600 , \21302_21601 , \21303_21602 , \21304_21603 , \21305_21604 , \21306_21605 ,
         \21307_21606 , \21308_21607 , \21309_21608 , \21310_21609 , \21311_21610 , \21312_21611 , \21313_21612 , \21314_21613 , \21315_21614 , \21316_21615 ,
         \21317_21616 , \21318_21617 , \21319_21618 , \21320_21619 , \21321_21620 , \21322_21621 , \21323_21622 , \21324_21623 , \21325_21624 , \21326_21625 ,
         \21327_21626 , \21328_21627 , \21329_21628 , \21330_21629 , \21331_21630 , \21332_21631 , \21333_21632 , \21334_21633 , \21335_21634 , \21336_21635 ,
         \21337_21636 , \21338_21637 , \21339 , \21340_21639 , \21341_21640 , \21342_21641 , \21343_21642 , \21344_21643 , \21345_21644 , \21346_21645 ,
         \21347_21646 , \21348_21647 , \21349_21648 , \21350_21649_nG441e , \21351_21650 , \21352_21651 , \21353_21652_nG4421 , \21354_21653 , \21355_21654 , \21356_21655 ,
         \21357_21659 , \21358_21660 , \21359_21661 , \21360_21662 , \21361_21663 , \21362_21664 , \21363_21665 , \21364_21666 , \21365_21667 , \21366_21668 ,
         \21367_21669 , \21368_21670 , \21369_21671 , \21370_21672 , \21371_21673 , \21372_21674 , \21373_21675 , \21374_21676 , \21375_21677 , \21376_21678 ,
         \21377_21679 , \21378_21680 , \21379_21681 , \21380_21682 , \21381_21683 , \21382_21684 , \21383_21685 , \21384_21686 , \21385_21687 , \21386_21688 ,
         \21387_21689 , \21388_21690 , \21389_21691 , \21390_21692 , \21391_21693 , \21392_21694 , \21393_21695 , \21394_21696 , \21395_21697 , \21396_21698 ,
         \21397_21699 , \21398_21700 , \21399_21701 , \21400_21702 , \21401_21703 , \21402_21704 , \21403_21705 , \21404_21706 , \21405_21707 , \21406_21708 ,
         \21407_21709 , \21408_21710 , \21409_21711 , \21410_21712 , \21411_21713 , \21412_21714 , \21413_21715 , \21414_21716 , \21415_21717 , \21416_21718 ,
         \21417_21719 , \21418_21720 , \21419_21721 , \21420_21722 , \21421_21723 , \21422_21724 , \21423_21725 , \21424_21726 , \21425_21727 , \21426_21728 ,
         \21427_21729 , \21428_21730 , \21429_21731 , \21430_21732 , \21431_21733 , \21432_21734 , \21433_21735 , \21434_21736 , \21435_21737 , \21436_21738 ,
         \21437_21739 , \21438_21740 , \21439_21741 , \21440_21742 , \21441_21743 , \21442_21744 , \21443_21745 , \21444_21746 , \21445_21747 , \21446_21748 ,
         \21447_21749 , \21448_21750 , \21449_21751 , \21450_21752 , \21451_21753 , \21452_21754 , \21453_21755 , \21454_21756 , \21455_21757 , \21456_21758 ,
         \21457_21759 , \21458_21760 , \21459_21761 , \21460_21762 , \21461_21763 , \21462_21764 , \21463_21765 , \21464_21766 , \21465_21767 , \21466_21768 ,
         \21467_21769 , \21468_21770 , \21469_21771 , \21470_21772 , \21471_21773 , \21472_21774 , \21473_21775 , \21474_21776 , \21475_21777 , \21476_21778 ,
         \21477_21779 , \21478_21780 , \21479_21781 , \21480_21782 , \21481_21783 , \21482_21784 , \21483_21785 , \21484_21786 , \21485_21787 , \21486_21788 ,
         \21487_21789 , \21488_21790 , \21489_21791 , \21490_21792 , \21491_21793 , \21492_21794 , \21493_21795 , \21494_21796 , \21495_21797 , \21496_21798 ,
         \21497_21799 , \21498_21800 , \21499_21801 , \21500_21802 , \21501_21803 , \21502_21804 , \21503_21805 , \21504_21806 , \21505_21807 , \21506_21808 ,
         \21507_21809 , \21508_21810 , \21509_21811 , \21510_21812 , \21511_21813 , \21512_21814 , \21513_21815 , \21514_21816 , \21515_21817 , \21516_21818 ,
         \21517_21819 , \21518_21820 , \21519_21821 , \21520_21822 , \21521_21823 , \21522_21824 , \21523_21825 , \21524_21826 , \21525_21827 , \21526_21828 ,
         \21527_21829 , \21528_21830 , \21529_21831 , \21530_21832 , \21531_21833 , \21532_21834 , \21533_21835 , \21534_21836 , \21535_21837 , \21536_21838 ,
         \21537_21839 , \21538_21840 , \21539_21841 , \21540_21842 , \21541_21843 , \21542_21844 , \21543_21845 , \21544_21846 , \21545_21847 , \21546_21848 ,
         \21547_21849 , \21548_21850 , \21549_21851 , \21550_21852 , \21551_21853 , \21552_21854 , \21553_21855 , \21554_21856 , \21555_21857 , \21556_21858 ,
         \21557_21859 , \21558_21860 , \21559_21861 , \21560_21862 , \21561_21863 , \21562_21864 , \21563_21865 , \21564_21866 , \21565_21867 , \21566_21868 ,
         \21567_21869 , \21568_21870 , \21569_21871 , \21570_21872 , \21571_21873 , \21572_21874 , \21573_21875 , \21574_21876 , \21575_21877 , \21576_21878 ,
         \21577_21879 , \21578_21880 , \21579_21881 , \21580_21882 , \21581_21883 , \21582_21884 , \21583_21885 , \21584_21886 , \21585_21887 , \21586_21888 ,
         \21587_21889 , \21588_21890 , \21589_21891 , \21590_21892 , \21591_21893 , \21592_21894 , \21593_21895 , \21594_21896 , \21595_21897 , \21596_21898 ,
         \21597_21899 , \21598_21900 , \21599_21901 , \21600_21902 , \21601_21903 , \21602_21904 , \21603_21905 , \21604_21906 , \21605_21907 , \21606_21908 ,
         \21607_21909 , \21608_21910 , \21609_21911 , \21610_21912 , \21611_21913 , \21612_21914 , \21613_21915 , \21614_21916 , \21615_21917 , \21616_21918 ,
         \21617_21919 , \21618_21920 , \21619_21921 , \21620_21922 , \21621_21923 , \21622_21924 , \21623_21925 , \21624_21926 , \21625_21927 , \21626_21928 ,
         \21627_21929 , \21628_21930 , \21629_21931 , \21630_21932 , \21631_21933 , \21632_21934 , \21633_21935 , \21634_21936 , \21635_21937 , \21636_21938 ,
         \21637_21939 , \21638_21940 , \21639_21941 , \21640_21942 , \21641_21943 , \21642_21944 , \21643_21945 , \21644_21946 , \21645_21947 , \21646_21948 ,
         \21647_21949 , \21648_21950 , \21649_21951 , \21650_21952 , \21651_21953 , \21652_21954 , \21653_21955 , \21654 , \21655_21957 , \21656_21958 ,
         \21657_21959 , \21658_21960 , \21659_21961 , \21660_21962 , \21661_21963 , \21662_21964 , \21663_21965 , \21664_21966 , \21665_21967 , \21666_21968 ,
         \21667_21969 , \21668_21970 , \21669_21971 , \21670_21972 , \21671_21973 , \21672_21974 , \21673_21975 , \21674_21976 , \21675_21977 , \21676_21978 ,
         \21677_21979 , \21678_21980 , \21679_21981 , \21680_21982 , \21681_21983 , \21682_21984 , \21683_21985 , \21684_21986 , \21685_21987 , \21686_21988 ,
         \21687_21989 , \21688_21990 , \21689_21991 , \21690_21992 , \21691_21993 , \21692_21994 , \21693_21995 , \21694_21996 , \21695_21997 , \21696_21998 ,
         \21697_21999 , \21698_22000 , \21699_22001 , \21700_22002 , \21701_22003 , \21702_22004 , \21703_22005 , \21704_22006 , \21705_22007 , \21706_22008 ,
         \21707_22009 , \21708_22010 , \21709_22011 , \21710_22012 , \21711_22013 , \21712_22014 , \21713_22015 , \21714_22016 , \21715_22017 , \21716_22018 ,
         \21717_22019 , \21718_22020 , \21719_22021 , \21720_22022 , \21721_22023 , \21722_22024 , \21723_22025 , \21724_22026 , \21725_22027 , \21726_22028 ,
         \21727_22029 , \21728_22030 , \21729_22031 , \21730_22032 , \21731_22033 , \21732_22034 , \21733_22035 , \21734_22036 , \21735_22037 , \21736_22038 ,
         \21737_22039 , \21738_22040 , \21739_22041 , \21740_22042 , \21741_22043 , \21742_22044 , \21743_22045 , \21744_22046 , \21745_22047 , \21746_22048 ,
         \21747_22049 , \21748_22050 , \21749_22051 , \21750_22052 , \21751_22053 , \21752_22054 , \21753_22055 , \21754_22056 , \21755_22057 , \21756_22058 ,
         \21757_22059 , \21758_22060 , \21759_22061 , \21760_22062 , \21761_22063 , \21762_22064 , \21763_22065 , \21764_22066 , \21765_22067 , \21766_22068 ,
         \21767_22069 , \21768_22070 , \21769_22071 , \21770_22072 , \21771_22073 , \21772_22074 , \21773_22075 , \21774_22076 , \21775_22077 , \21776_22078 ,
         \21777_22079 , \21778_22080 , \21779_22081 , \21780_22082 , \21781_22083 , \21782_22084 , \21783_22085 , \21784_22086 , \21785_22087 , \21786 ,
         \21787_22089_nG65af , \21788_22090 , \21789_22091 , \21790_22092 , \21791_22093 , \21792_22094 , \21793_22095 , \21794_22096 , \21795_22097 , \21796_22098 ,
         \21797 , \21798 , \21799_22101_nG5801 , \21800_22102 , \21801_22103 , \21802_22104 , \21803_22105 , \21804_22106 , \21805_22107 , \21806_22108 ,
         \21807_22109 , \21808_22110 , \21809_22111 , \21810_22112 , \21811_22113 , \21812_22114 , \21813_22115 , \21814_22116 , \21815_22117 , \21816_22118 ,
         \21817_22119 , \21818_22120 , \21819_22121 , \21820_22122 , \21821_22123 , \21822_22124 , \21823_22125 , \21824_22126 , \21825_22127 , \21826_22128 ,
         \21827_22129_nG9bd8 , \21828_22130 , \21829_22131 , \21830_22132 , \21831_22133 , \21832_22134 , \21833_22135 , \21834_22136 , \21835_22137 , \21836_22138 ,
         \21837_22139 , \21838_22140 , \21839_22141 , \21840_22142 , \21841_22143 , \21842_22144 , \21843_22145 , \21844_22146 , \21845_22147 , \21846_22148 ,
         \21847_22149 , \21848_22150 , \21849_22151 , \21850_22152 , \21851_22153 , \21852_22154 , \21853_22155 , \21854_22156 , \21855_22157 , \21856_22158 ,
         \21857_22159 , \21858_22160 , \21859_22161 , \21860_22162 , \21861_22163 , \21862_22164 , \21863_22165 , \21864_22166 , \21865_22167 , \21866_22168 ,
         \21867_22169 , \21868_22170 , \21869_22171 , \21870_22172 , \21871_22173 , \21872_22174 , \21873_22175 , \21874_22176 , \21875_22177 , \21876_22178 ,
         \21877_22179 , \21878_22180 , \21879_22181 , \21880_22182 , \21881_22183 , \21882_22184 , \21883_22185 , \21884_22186 , \21885_22187 , \21886_22188 ,
         \21887_22189 , \21888_22190 , \21889_22191 , \21890_22192 , \21891_22193 , \21892_22194 , \21893_22195 , \21894_22196 , \21895_22197 , \21896_22198 ,
         \21897_22199 , \21898_22200 , \21899_22201 , \21900_22202 , \21901_22203 , \21902_22204 , \21903_22205 , \21904_22206 , \21905_22207 , \21906_21656 ,
         \21907_21657 , \21908_21658 , \21909_22208 , \21910_22209 , \21911_22210 , \21912_22211 , \21913_22212 , \21914_22213 , \21915_22214 , \21916_22215 ,
         \21917_22216 , \21918_22217 , \21919_22218 , \21920_22219 , \21921_22220 , \21922_22221 , \21923_22222 , \21924_22223 , \21925_22224 , \21926_22225 ,
         \21927_22226 , \21928_22227 , \21929_22228 , \21930_22229 , \21931_22230 , \21932_22231 , \21933_22232 , \21934_22233 , \21935_22234 , \21936_22235 ,
         \21937_22236 , \21938_22237 , \21939_22238 , \21940_22239 , \21941_22240 , \21942_22241 , \21943_22242 , \21944_22243 , \21945_22244 , \21946_22245 ,
         \21947_22246 , \21948_22247 , \21949_22248 , \21950_22249 , \21951_22250 , \21952_22251 , \21953_22252 , \21954_22253 , \21955_22254 , \21956_22255 ,
         \21957_22256 , \21958_22257 , \21959_22258 , \21960_22259 , \21961_22260 , \21962_22261 , \21963_22262 , \21964_22263 , \21965_22264 , \21966_22265 ,
         \21967_22266 , \21968_22267 , \21969_22268 , \21970_22269 , \21971_22270 , \21972_22271 , \21973_22272 , \21974_22273 , \21975_22274 , \21976_22275 ,
         \21977_22276 , \21978_22277 , \21979_22278 , \21980_22279 , \21981_22280 , \21982_22281 , \21983_22282 , \21984_22283 , \21985_22284 , \21986_22285 ,
         \21987_22286 , \21988_22287 , \21989_22288 , \21990_22289 , \21991_22290 , \21992_22291 , \21993_22292 , \21994_22293 , \21995_22294 , \21996_22295 ,
         \21997_22296 , \21998_22297 , \21999_22298 , \22000_22299 , \22001_22300 , \22002_22301 , \22003_22302 , \22004_22303 , \22005_22304 , \22006_22305 ,
         \22007_22306 , \22008_22307 , \22009_22308 , \22010_22309 , \22011_22310 , \22012_22311 , \22013_22312 , \22014_22313 , \22015_22314 , \22016_22315 ,
         \22017_22316 , \22018_22317 , \22019_22318 , \22020_22319 , \22021_22320 , \22022_22321 , \22023_22322 , \22024_22323 , \22025_22324 , \22026_22325 ,
         \22027_22326 , \22028_22327 , \22029_22328 , \22030_22329 , \22031_22330 , \22032_22331 , \22033_22332 , \22034_22333 , \22035_22334 , \22036_22335 ,
         \22037_22336 , \22038_22337 , \22039_22338 , \22040_22339 , \22041_22340 , \22042_22341 , \22043_22342 , \22044_22343 , \22045_22344 , \22046_22345 ,
         \22047_22346 , \22048_22347 , \22049_22348 , \22050_22349 , \22051_22350 , \22052_22351 , \22053_22352 , \22054_22353 , \22055_22354 , \22056_22355 ,
         \22057_22356 , \22058_22357 , \22059_22358 , \22060_22359 , \22061_22360 , \22062_22361 , \22063_22362 , \22064_22363 , \22065_22364 , \22066_22365 ,
         \22067_22366 , \22068_22367 , \22069_22368 , \22070_22369 , \22071_22370 , \22072_22371 , \22073_22372 , \22074_22373 , \22075_22374 , \22076_22375 ,
         \22077_22376 , \22078_22377 , \22079_22378 , \22080_22379 , \22081_22380 , \22082_22381 , \22083_22382 , \22084_22383 , \22085_22384 , \22086_22385 ,
         \22087_22386 , \22088_22387 , \22089_22388 , \22090_22389 , \22091_22390 , \22092_22391 , \22093_22392 , \22094_22393 , \22095_22394 , \22096_22395 ,
         \22097_22396 , \22098_22397 , \22099_22398 , \22100_22399 , \22101_22400 , \22102_22401 , \22103_22402 , \22104_22403 , \22105_22404 , \22106 ,
         \22107_22406 , \22108_22407 , \22109_22408 , \22110_22409 , \22111_22410 , \22112_22411 , \22113_22412 , \22114_22413 , \22115_22414 , \22116_22415 ,
         \22117_22416 , \22118_22417 , \22119_22418 , \22120_22419 , \22121_22420 , \22122_22421 , \22123_22422 , \22124_22423 , \22125_22424 , \22126_22425 ,
         \22127_22426 , \22128_22427 , \22129_22428 , \22130_22429 , \22131_22430 , \22132_22431 , \22133_22432 , \22134_22433 , \22135_22434 , \22136_22435 ,
         \22137_22436 , \22138_22437 , \22139_22438 , \22140_22439 , \22141_22440 , \22142_22441 , \22143_22442 , \22144_22443 , \22145_22444 , \22146_22445 ,
         \22147_22446 , \22148_22447 , \22149_22448 , \22150_22449 , \22151_22450 , \22152_22451 , \22153_22452 , \22154_22453 , \22155_22454 , \22156_22455 ,
         \22157_22456 , \22158_22457 , \22159_22458 , \22160_22459 , \22161_22460 , \22162_22461 , \22163_22462 , \22164_22463 , \22165_22464 , \22166_22465 ,
         \22167_22466 , \22168_22467 , \22169_22468 , \22170_22469 , \22171_22470 , \22172_22471 , \22173_22472 , \22174_22473 , \22175_22474 , \22176_22475 ,
         \22177_22476 , \22178_22477 , \22179_22478 , \22180_22479 , \22181_22480 , \22182_22481 , \22183_22482 , \22184_22483 , \22185_22484 , \22186_22485 ,
         \22187_22486 , \22188_22487 , \22189_22488 , \22190_22489 , \22191_22490 , \22192_22491 , \22193_22492 , \22194_22493 , \22195_22494 , \22196_22495 ,
         \22197_22496 , \22198_22497 , \22199_22498 , \22200_22499 , \22201_22500 , \22202_22501 , \22203_22502 , \22204_22503 , \22205_22504 , \22206_22505 ,
         \22207_22506 , \22208_22507 , \22209_22508 , \22210_22509 , \22211_22510 , \22212_22511 , \22213_22512 , \22214_22513 , \22215_22514 , \22216_22515 ,
         \22217_22516 , \22218_22517 , \22219_22518 , \22220_22519 , \22221_22520 , \22222_22521 , \22223_22522 , \22224_22523 , \22225_22524 , \22226_22525 ,
         \22227_22526 , \22228_22527 , \22229_22528 , \22230_22529 , \22231_22530 , \22232_22531 , \22233_22532 , \22234_22533 , \22235_22534 , \22236_22535 ,
         \22237_22536 , \22238 , \22239_22538_nG590a , \22240_22539 , \22241_22540 , \22242_22541 , \22243_22542 , \22244_22543 , \22245_22544 , \22246_22545 ,
         \22247_22546 , \22248_22547 , \22249_22548 , \22250_22549 , \22251_22550 , \22252_22551 , \22253_22552 , \22254 , \22255 , \22256_22555_nG65b2 ,
         \22257_22556 , \22258_22557 , \22259_22558 , \22260_22559 , \22261_22560 , \22262_22561 , \22263_22562 , \22264_22563 , \22265_22564 , \22266_22565 ,
         \22267_22566 , \22268_22567 , \22269_22568 , \22270_22569 , \22271_22570 , \22272_22571 , \22273_22572 , \22274_22573 , \22275_22574 , \22276_22575 ,
         \22277_22576 , \22278_22577 , \22279_22578 , \22280_22579 , \22281_22580 , \22282_22581 , \22283_22582 , \22284_22583 , \22285_22584 , \22286_22585 ,
         \22287_22586 , \22288_22587 , \22289_22588 , \22290_22589 , \22291_22590 , \22292_22591 , \22293_22592 , \22294_22593 , \22295_22594 , \22296_22595 ,
         \22297_22596 , \22298_22597 , \22299_22598 , \22300_22599 , \22301_22600 , \22302_22601 , \22303_22602 , \22304_22603 , \22305_22604 , \22306_22605 ,
         \22307_22606 , \22308_22607 , \22309_22608 , \22310_22609 , \22311_22610 , \22312_22611 , \22313_22612 , \22314_22613 , \22315_22614 , \22316_22615 ,
         \22317_22616 , \22318_22617 , \22319_22618 , \22320_22619 , \22321_22620 , \22322_22621 , \22323_22622 , \22324_22623 , \22325_22624 , \22326_22625 ,
         \22327_22626 , \22328_22627 , \22329_22628 , \22330_22629_nG9bd5 , \22331_22630 , \22332_22631 , \22333_22632 , \22334_22633 , \22335_22634 , \22336_22635 ,
         \22337_22636 , \22338_22637 , \22339_22638 , \22340_22639 , \22341_22640 , \22342_22641 , \22343_22642 , \22344_22643 , \22345_22644 , \22346_22645 ,
         \22347_22646 , \22348_22647 , \22349_22648 , \22350_22649 , \22351_22650 , \22352_22651 , \22353_22652 , \22354_22653 , \22355_22654 , \22356_22655 ,
         \22357_22656 , \22358_22657 , \22359_22658 , \22360_22659 , \22361_22660 , \22362_22661 , \22363_22662 , \22364_22663 , \22365_22664 , \22366_22665 ,
         \22367_22666 , \22368_22667 , \22369_22668 , \22370_22669 , \22371_22670 , \22372_22671 , \22373_22672 , \22374_22673 , \22375_22674 , \22376_22675 ,
         \22377_22676 , \22378_22677 , \22379_22678 , \22380_22679 , \22381_22680 , \22382_22681 , \22383_22682 , \22384_22683 , \22385_22684 , \22386_22685 ,
         \22387_22686 , \22388_22687 , \22389_22688 , \22390_22689 , \22391_22690 , \22392_22691 , \22393_22692 , \22394_22693 , \22395_22694 , \22396_22695 ,
         \22397_22696 , \22398_22697 , \22399_22698 , \22400_22699 , \22401_22700 , \22402_22701 , \22403_22702 , \22404_22703 , \22405_22704 , \22406_22705 ,
         \22407_22706 , \22408_22707 , \22409_22708 , \22410_22709 , \22411_22710 , \22412_22711 , \22413_22712 , \22414_22713 , \22415_22714 , \22416_22715 ,
         \22417_22716 , \22418_22717 , \22419_22718 , \22420_22719 , \22421_22720 , \22422_22721 , \22423_22722 , \22424_22723 , \22425_22724 , \22426_22725 ,
         \22427_22726 , \22428_22727 , \22429_22728 , \22430_22729 , \22431_22730 , \22432_22731 , \22433_22732 , \22434_22733 , \22435_22734 , \22436_22735 ,
         \22437_22736 , \22438_22737 , \22439_22738 , \22440_22739 , \22441_22740 , \22442_22741 , \22443_22742 , \22444_22743 , \22445_22744 , \22446_22745 ,
         \22447_22746 , \22448_22747 , \22449_22748 , \22450_22749 , \22451_22750 , \22452_22751 , \22453_22752 , \22454_22753 , \22455_22754 , \22456_22755 ,
         \22457_22756 , \22458_22757 , \22459_22758 , \22460_22759 , \22461_22760 , \22462_22761 , \22463_22762 , \22464_22763 , \22465_22764 , \22466_22765 ,
         \22467_22766 , \22468_22767 , \22469_22768 , \22470_22769 , \22471_22770 , \22472_22771 , \22473_22772 , \22474_22773 , \22475_22774 , \22476_22775 ,
         \22477_22776 , \22478_22777 , \22479_22778 , \22480_22779 , \22481_22780 , \22482 , \22483_22782 , \22484_22783 , \22485_22784 , \22486_22785 ,
         \22487_22786 , \22488_22787 , \22489_22788 , \22490_22789 , \22491_22790 , \22492_22791 , \22493_22792 , \22494_22793 , \22495_22794 , \22496_22795 ,
         \22497_22796 , \22498_22797 , \22499_22798 , \22500_22799 , \22501_22800 , \22502_22801 , \22503_22802 , \22504_22803 , \22505_22804 , \22506_22805 ,
         \22507_22806 , \22508_22807 , \22509_22808 , \22510_22809 , \22511_22810 , \22512_22811 , \22513_22812 , \22514_22813 , \22515_22814 , \22516_22815 ,
         \22517_22816 , \22518_22817 , \22519_22818 , \22520_22819 , \22521_22820 , \22522_22821 , \22523_22822 , \22524_22823 , \22525_22824 , \22526_22825 ,
         \22527_22826 , \22528_22827 , \22529_22828 , \22530_22829 , \22531_22830 , \22532_22831 , \22533_22832 , \22534_22833 , \22535_22834 , \22536_22835 ,
         \22537_22836 , \22538_22837 , \22539_22838 , \22540_22839 , \22541_22840 , \22542_22841 , \22543_22842 , \22544_22843 , \22545_22844 , \22546_22845 ,
         \22547_22846 , \22548_22847 , \22549_22848 , \22550_22849 , \22551_22850 , \22552_22851 , \22553_22852 , \22554_22853 , \22555_22854 , \22556_22855 ,
         \22557_22856 , \22558_22857 , \22559_22858 , \22560_22859 , \22561_22860 , \22562_22861 , \22563_22862 , \22564_22863 , \22565_22864 , \22566_22865 ,
         \22567_22866 , \22568_22867 , \22569_22868 , \22570_22869 , \22571_22870 , \22572_22871 , \22573_22872 , \22574_22873 , \22575_22874 , \22576_22875 ,
         \22577_22876 , \22578_22877 , \22579_22878 , \22580_22879 , \22581_22880 , \22582_22881 , \22583_22882 , \22584_22883 , \22585_22884 , \22586_22885 ,
         \22587_22886 , \22588_22887 , \22589_22888 , \22590_22889 , \22591_22890 , \22592_22891 , \22593_22892 , \22594_22893 , \22595_22894 , \22596_22895 ,
         \22597_22896 , \22598_22897 , \22599_22898 , \22600_22899 , \22601_22900 , \22602_22901 , \22603_22902 , \22604_22903 , \22605_22904 , \22606_22905 ,
         \22607_22906 , \22608_22907 , \22609_22908 , \22610_22909 , \22611_22910 , \22612_22911 , \22613_22912 , \22614_22913 , \22615 , \22616_22915 ,
         \22617_22916 , \22618_22917 , \22619_22918 , \22620_22919 , \22621_22920 , \22622_22921 , \22623_22922 , \22624_22923 , \22625_22924 , \22626_22925 ,
         \22627_22926 , \22628_22927 , \22629_22928 , \22630_22929 , \22631_22930 , \22632_22931 , \22633_22932 , \22634_22933 , \22635_22934 , \22636_22935 ,
         \22637_22936 , \22638_22937 , \22639_22938 , \22640_22939 , \22641_22940 , \22642_22941 , \22643_22942 , \22644_22943 , \22645_22944 , \22646_22945 ,
         \22647_22946 , \22648_22947 , \22649_22948 , \22650_22949 , \22651_22950 , \22652_22951 , \22653_22952 , \22654_22953 , \22655_22954 , \22656_22955 ,
         \22657_22956 , \22658_22957 , \22659_22958 , \22660_22959 , \22661_22960 , \22662_22961 , \22663_22962 , \22664_22963 , \22665_22964 , \22666_22965 ,
         \22667_22966 , \22668_22967 , \22669_22968 , \22670_22969 , \22671_22970 , \22672_22971 , \22673_22972 , \22674_22973 , \22675_22974 , \22676_22975 ,
         \22677_22976 , \22678_22977 , \22679_22978 , \22680_22979 , \22681_22980 , \22682_22981 , \22683_22982 , \22684_22983 , \22685_22984 , \22686_22985 ,
         \22687_22986 , \22688_22987 , \22689_22988 , \22690_22989 , \22691_22990 , \22692_22991 , \22693_22992 , \22694_22993 , \22695_22994 , \22696_22995 ,
         \22697_22996 , \22698_22997 , \22699_22998 , \22700_22999 , \22701_23000 , \22702_23001 , \22703_23002 , \22704_23003 , \22705_23004 , \22706_23005 ,
         \22707_23006 , \22708_23007 , \22709_23008 , \22710_23009 , \22711_23010 , \22712_23011 , \22713_23012 , \22714_23013 , \22715_23014 , \22716_23015 ,
         \22717_23016 , \22718_23017 , \22719_23018 , \22720_23019 , \22721_23020 , \22722_23021 , \22723_23022 , \22724_23023 , \22725_23024 , \22726_23025 ,
         \22727_23026 , \22728_23027 , \22729_23028 , \22730_23029 , \22731_23030 , \22732_23031 , \22733_23032 , \22734_23033 , \22735_23034 , \22736_23035 ,
         \22737_23036 , \22738_23037 , \22739_23038 , \22740_23039 , \22741_23040 , \22742_23041 , \22743_23042 , \22744_23043 , \22745_23044 , \22746_23045 ,
         \22747_23046 , \22748_23047 , \22749 , \22750_23049 , \22751_23050 , \22752_23051 , \22753_23052 , \22754_23053 , \22755_23054 , \22756_23055 ,
         \22757_23056 , \22758_23057 , \22759_23058 , \22760_23059 , \22761_23060 , \22762_23061 , \22763_23062 , \22764_23063 , \22765_23064 , \22766_23065 ,
         \22767_23066 , \22768_23067 , \22769_23068 , \22770_23069 , \22771_23070 , \22772_23071 , \22773_23072 , \22774_23073 , \22775_23074 , \22776_23075 ,
         \22777_23076 , \22778_23077 , \22779_23078 , \22780_23079 , \22781_23080 , \22782_23081 , \22783_23082 , \22784_23083 , \22785_23084 , \22786_23085 ,
         \22787_23086 , \22788_23087 , \22789_23088 , \22790_23089 , \22791_23090 , \22792_23091 , \22793_23092 , \22794_23093 , \22795_23094 , \22796_23095 ,
         \22797_23096 , \22798_23097 , \22799_23098 , \22800_23099 , \22801_23100 , \22802_23101 , \22803_23102 , \22804_23103 , \22805_23104 , \22806_23105 ,
         \22807_23106 , \22808_23107 , \22809_23108 , \22810_23109 , \22811_23110 , \22812_23111 , \22813_23112 , \22814_23113 , \22815_23114 , \22816_23115 ,
         \22817_23116 , \22818_23117 , \22819_23118 , \22820_23119 , \22821_23120 , \22822_23121 , \22823_23122 , \22824_23123 , \22825_23124 , \22826_23125 ,
         \22827_23126 , \22828_23127 , \22829_23128 , \22830_23129 , \22831_23130 , \22832_23131 , \22833_23132 , \22834_23133 , \22835_23134 , \22836_23135 ,
         \22837_23136 , \22838_23137 , \22839_23138 , \22840_23139 , \22841_23140 , \22842_23141 , \22843_23142 , \22844_23143 , \22845_23144 , \22846_23145 ,
         \22847_23146 , \22848_23147 , \22849_23148 , \22850_23149 , \22851_23150 , \22852_23151 , \22853_23152 , \22854_23153 , \22855_23154 , \22856_23155 ,
         \22857_23156 , \22858_23157 , \22859_23158 , \22860_23159 , \22861_23160 , \22862_23161 , \22863_23162 , \22864_23163 , \22865_23164 , \22866_23165 ,
         \22867_23166 , \22868_23167 , \22869_23168 , \22870_23169 , \22871_23170 , \22872_23171 , \22873_23172 , \22874_23173 , \22875_23174 , \22876_23175 ,
         \22877_23176 , \22878_23177 , \22879_23178 , \22880_23179 , \22881_23180 , \22882 , \22883_23182 , \22884_23183 , \22885_23184 , \22886_23185 ,
         \22887_23186 , \22888_23187 , \22889_23188 , \22890_23189 , \22891_23190 , \22892_23191 , \22893_23192_nG4418 , \22894_23193 , \22895_23194 , \22896_23195_nG441b ,
         \22897_23196 , \22898_23197 , \22899_23198 , \22900_23202 , \22901_23203 , \22902_23204 , \22903_23205 , \22904_23206 , \22905_23207 , \22906_23208 ,
         \22907_23209 , \22908_23210 , \22909_23211 , \22910_23212 , \22911_23213 , \22912_23214 , \22913_23215 , \22914_23216 , \22915_23217 , \22916_23218 ,
         \22917_23219 , \22918_23220 , \22919_23221 , \22920_23222 , \22921_23223 , \22922_23224 , \22923_23225 , \22924_23226 , \22925_23227 , \22926_23228 ,
         \22927_23229 , \22928_23230 , \22929_23231 , \22930_23232 , \22931_23233 , \22932_23234 , \22933_23235 , \22934_23236 , \22935_23237 , \22936_23238 ,
         \22937_23239 , \22938_23240 , \22939_23241 , \22940_23242 , \22941_23243 , \22942_23244 , \22943_23245 , \22944_23246 , \22945_23247 , \22946_23248 ,
         \22947_23249 , \22948_23250 , \22949_23251 , \22950_23252 , \22951_23253 , \22952_23254 , \22953_23255 , \22954_23256 , \22955_23257 , \22956_23258 ,
         \22957_23259 , \22958_23260 , \22959_23261 , \22960_23262 , \22961_23263 , \22962_23264 , \22963_23265 , \22964_23266 , \22965_23267 , \22966_23268 ,
         \22967_23269 , \22968_23270 , \22969_23271 , \22970_23272 , \22971_23273 , \22972_23274 , \22973_23275 , \22974_23276 , \22975_23277 , \22976_23278 ,
         \22977_23279 , \22978_23280 , \22979_23281 , \22980_23282 , \22981_23283 , \22982_23284 , \22983_23285 , \22984_23286 , \22985_23287 , \22986_23288 ,
         \22987_23289 , \22988_23290 , \22989_23291 , \22990_23292 , \22991_23293 , \22992_23294 , \22993_23295 , \22994_23296 , \22995_23297 , \22996_23298 ,
         \22997_23299 , \22998_23300 , \22999_23301 , \23000_23302 , \23001_23303 , \23002_23304 , \23003_23305 , \23004_23306 , \23005_23307 , \23006_23308 ,
         \23007_23309 , \23008_23310 , \23009_23311 , \23010_23312 , \23011_23313 , \23012_23314 , \23013_23315 , \23014_23316 , \23015_23317 , \23016_23318 ,
         \23017_23319 , \23018_23320 , \23019_23321 , \23020_23322 , \23021_23323 , \23022_23324 , \23023_23325 , \23024_23326 , \23025_23327 , \23026_23328 ,
         \23027_23329 , \23028_23330 , \23029_23331 , \23030_23332 , \23031_23333 , \23032_23334 , \23033_23335 , \23034_23336 , \23035_23337 , \23036_23338 ,
         \23037_23339 , \23038_23340 , \23039_23341 , \23040_23342 , \23041_23343 , \23042_23344 , \23043_23345 , \23044_23346 , \23045_23347 , \23046_23348 ,
         \23047_23349 , \23048_23350 , \23049_23351 , \23050_23352 , \23051_23353 , \23052_23354 , \23053_23355 , \23054_23356 , \23055_23357 , \23056_23358 ,
         \23057_23359 , \23058_23360 , \23059_23361 , \23060_23362 , \23061_23363 , \23062_23364 , \23063_23365 , \23064_23366 , \23065_23367 , \23066_23368 ,
         \23067_23369 , \23068_23370 , \23069_23371 , \23070_23372 , \23071_23373 , \23072_23374 , \23073_23375 , \23074_23376 , \23075_23377 , \23076_23378 ,
         \23077_23379 , \23078_23380 , \23079_23381 , \23080_23382 , \23081_23383 , \23082_23384 , \23083_23385 , \23084_23386 , \23085_23387 , \23086_23388 ,
         \23087_23389 , \23088_23390 , \23089_23391 , \23090_23392 , \23091_23393 , \23092_23394 , \23093_23395 , \23094_23396 , \23095_23397 , \23096_23398 ,
         \23097_23399 , \23098_23400 , \23099_23401 , \23100_23402 , \23101_23403 , \23102_23404 , \23103_23405 , \23104_23406 , \23105_23407 , \23106_23408 ,
         \23107_23409 , \23108_23410 , \23109_23411 , \23110_23412 , \23111_23413 , \23112_23414 , \23113_23415 , \23114_23416 , \23115_23417 , \23116_23418 ,
         \23117_23419 , \23118_23420 , \23119_23421 , \23120_23422 , \23121_23423 , \23122_23424 , \23123_23425 , \23124_23426 , \23125_23427 , \23126_23428 ,
         \23127_23429 , \23128_23430 , \23129_23431 , \23130_23432 , \23131_23433 , \23132_23434 , \23133_23435 , \23134_23436 , \23135_23437 , \23136_23438 ,
         \23137_23439 , \23138_23440 , \23139_23441 , \23140_23442 , \23141_23443 , \23142_23444 , \23143_23445 , \23144_23446 , \23145_23447 , \23146_23448 ,
         \23147_23449 , \23148_23450 , \23149_23451 , \23150_23452 , \23151_23453 , \23152_23454 , \23153_23455 , \23154_23456 , \23155_23457 , \23156_23458 ,
         \23157_23459 , \23158_23460 , \23159_23461 , \23160_23462 , \23161_23463 , \23162_23464 , \23163_23465 , \23164_23466 , \23165_23467 , \23166_23468 ,
         \23167_23469 , \23168_23470 , \23169_23471 , \23170_23472 , \23171_23473 , \23172_23474 , \23173_23475 , \23174_23476 , \23175_23477 , \23176_23478 ,
         \23177_23479 , \23178_23480 , \23179_23481 , \23180_23482 , \23181 , \23182_23484 , \23183_23485 , \23184_23486 , \23185_23487 , \23186_23488 ,
         \23187_23489 , \23188_23490 , \23189_23491 , \23190_23492 , \23191_23493 , \23192_23494 , \23193_23495 , \23194_23496 , \23195_23497 , \23196_23498 ,
         \23197_23499 , \23198_23500 , \23199_23501 , \23200_23502 , \23201_23503 , \23202_23504 , \23203_23505 , \23204_23506 , \23205_23507 , \23206_23508 ,
         \23207_23509 , \23208_23510 , \23209_23511 , \23210_23512 , \23211_23513 , \23212_23514 , \23213_23515 , \23214_23516 , \23215_23517 , \23216_23518 ,
         \23217_23519 , \23218_23520 , \23219_23521 , \23220_23522 , \23221_23523 , \23222_23524 , \23223_23525 , \23224_23526 , \23225_23527 , \23226_23528 ,
         \23227_23529 , \23228_23530 , \23229_23531 , \23230_23532 , \23231_23533 , \23232_23534 , \23233_23535 , \23234_23536 , \23235_23537 , \23236_23538 ,
         \23237_23539 , \23238_23540 , \23239_23541 , \23240_23542 , \23241_23543 , \23242_23544 , \23243_23545 , \23244_23546 , \23245_23547 , \23246_23548 ,
         \23247_23549 , \23248_23550 , \23249_23551 , \23250_23552 , \23251_23553 , \23252_23554 , \23253_23555 , \23254_23556 , \23255_23557 , \23256_23558 ,
         \23257_23559 , \23258_23560 , \23259_23561 , \23260_23562 , \23261_23563 , \23262_23564 , \23263_23565 , \23264_23566 , \23265_23567 , \23266_23568 ,
         \23267_23569 , \23268_23570 , \23269_23571 , \23270_23572 , \23271_23573 , \23272_23574 , \23273_23575 , \23274_23576 , \23275_23577 , \23276_23578 ,
         \23277_23579 , \23278_23580 , \23279_23581 , \23280_23582 , \23281_23583 , \23282_23584 , \23283_23585 , \23284_23586 , \23285_23587 , \23286_23588 ,
         \23287_23589 , \23288_23590 , \23289_23591 , \23290_23592 , \23291_23593 , \23292_23594 , \23293_23595 , \23294_23596 , \23295_23597 , \23296_23598 ,
         \23297_23599 , \23298_23600 , \23299_23601 , \23300_23602 , \23301_23603 , \23302_23604 , \23303_23605 , \23304_23606 , \23305_23607 , \23306_23608 ,
         \23307_23609 , \23308_23610 , \23309_23611 , \23310_23612 , \23311_23613 , \23312_23614 , \23313 , \23314_23616_nG65b5 , \23315_23617 , \23316_23618 ,
         \23317_23619 , \23318_23620 , \23319_23621 , \23320_23622 , \23321_23623 , \23322_23624 , \23323_23625 , \23324 , \23325 , \23326_23628_nG5a13 ,
         \23327_23629 , \23328_23630 , \23329_23631 , \23330_23632 , \23331_23633 , \23332_23634 , \23333_23635 , \23334_23636 , \23335_23637 , \23336_23638 ,
         \23337_23639 , \23338_23640 , \23339_23641 , \23340_23642 , \23341_23643 , \23342_23644 , \23343_23645 , \23344_23646 , \23345_23647 , \23346_23648 ,
         \23347_23649 , \23348_23650 , \23349_23651 , \23350_23652 , \23351_23653 , \23352_23654 , \23353_23655 , \23354_23656 , \23355_23657 , \23356_23658 ,
         \23357_23659 , \23358_23660 , \23359_23661 , \23360_23662 , \23361_23663 , \23362_23664 , \23363_23665 , \23364_23666 , \23365_23667 , \23366_23668 ,
         \23367_23669 , \23368_23670 , \23369_23671 , \23370_23672 , \23371_23673 , \23372_23674 , \23373_23675 , \23374_23676 , \23375_23677 , \23376_23678 ,
         \23377_23679 , \23378_23680 , \23379_23681 , \23380_23682 , \23381_23683 , \23382_23684 , \23383_23685 , \23384_23686 , \23385_23687 , \23386_23688 ,
         \23387_23689 , \23388_23690 , \23389_23691 , \23390_23692 , \23391_23693 , \23392_23694 , \23393_23695 , \23394_23696_nG9bd2 , \23395_23697 , \23396_23698 ,
         \23397_23699 , \23398_23700 , \23399_23701 , \23400_23702 , \23401_23703 , \23402_23704 , \23403_23705 , \23404_23706 , \23405_23707 , \23406_23708 ,
         \23407_23709 , \23408_23710 , \23409_23711 , \23410_23712 , \23411_23713 , \23412_23714 , \23413_23715 , \23414_23716 , \23415_23717 , \23416_23718 ,
         \23417_23719 , \23418_23720 , \23419_23721 , \23420_23722 , \23421_23723 , \23422_23724 , \23423_23725 , \23424_23726 , \23425_23727 , \23426_23728 ,
         \23427_23729 , \23428_23730 , \23429_23731 , \23430_23732 , \23431_23733 , \23432_23734 , \23433_23735 , \23434_23736 , \23435_23737 , \23436_23738 ,
         \23437_23739 , \23438_23740 , \23439_23741 , \23440_23742 , \23441_23743 , \23442_23744 , \23443_23745 , \23444_23746 , \23445_23747 , \23446_23748 ,
         \23447_23749 , \23448_23750 , \23449_23751 , \23450_23752 , \23451_23753 , \23452_23754 , \23453_23755 , \23454_23756 , \23455_23757 , \23456_23758 ,
         \23457_23759 , \23458_23760 , \23459_23761 , \23460_23762 , \23461_23763 , \23462_23764 , \23463_23765 , \23464_23766 , \23465_23767 , \23466_23768 ,
         \23467_23769 , \23468_23770 , \23469_23771 , \23470_23772 , \23471_23773 , \23472_23774 , \23473_23775 , \23474_23776 , \23475_23777 , \23476_23778 ,
         \23477_23779 , \23478_23780 , \23479_23781 , \23480_23782 , \23481_23783 , \23482_23784 , \23483_23785 , \23484_23786 , \23485_23787 , \23486_23788 ,
         \23487_23789 , \23488_23790 , \23489_23791 , \23490_23792 , \23491_23793 , \23492_23794 , \23493_23199 , \23494_23200 , \23495_23201 , \23496_23795 ,
         \23497_23796 , \23498_23797 , \23499_23798 , \23500_23799 , \23501_23800 , \23502_23801 , \23503_23802 , \23504_23803 , \23505_23804 , \23506_23805 ,
         \23507_23806 , \23508_23807 , \23509_23808 , \23510_23809 , \23511_23810 , \23512_23811 , \23513_23812 , \23514_23813 , \23515_23814 , \23516_23815 ,
         \23517_23816 , \23518_23817 , \23519_23818 , \23520_23819 , \23521_23820 , \23522_23821 , \23523_23822 , \23524_23823 , \23525_23824 , \23526_23825 ,
         \23527_23826 , \23528_23827 , \23529_23828 , \23530_23829 , \23531_23830 , \23532_23831 , \23533_23832 , \23534_23833 , \23535_23834 , \23536_23835 ,
         \23537_23836 , \23538_23837 , \23539_23838 , \23540_23839 , \23541_23840 , \23542_23841 , \23543_23842 , \23544_23843 , \23545_23844 , \23546_23845 ,
         \23547_23846 , \23548_23847 , \23549_23848 , \23550_23849 , \23551_23850 , \23552_23851 , \23553_23852 , \23554_23853 , \23555_23854 , \23556_23855 ,
         \23557_23856 , \23558_23857 , \23559_23858 , \23560_23859 , \23561_23860 , \23562_23861 , \23563_23862 , \23564_23863 , \23565_23864 , \23566_23865 ,
         \23567_23866 , \23568_23867 , \23569_23868 , \23570_23869 , \23571_23870 , \23572_23871 , \23573_23872 , \23574_23873 , \23575_23874 , \23576_23875 ,
         \23577_23876 , \23578_23877 , \23579_23878 , \23580_23879 , \23581_23880 , \23582_23881 , \23583_23882 , \23584_23883 , \23585_23884 , \23586_23885 ,
         \23587_23886 , \23588_23887 , \23589_23888 , \23590_23889 , \23591_23890 , \23592_23891 , \23593_23892 , \23594_23893 , \23595_23894 , \23596_23895 ,
         \23597_23896 , \23598_23897 , \23599_23898 , \23600_23899 , \23601_23900 , \23602_23901 , \23603_23902 , \23604_23903 , \23605_23904 , \23606_23905 ,
         \23607_23906 , \23608_23907 , \23609_23908 , \23610_23909 , \23611_23910 , \23612_23911 , \23613_23912 , \23614_23913 , \23615_23914 , \23616_23915 ,
         \23617_23916 , \23618_23917 , \23619_23918 , \23620_23919 , \23621_23920 , \23622_23921 , \23623_23922 , \23624_23923 , \23625_23924 , \23626_23925 ,
         \23627_23926 , \23628_23927 , \23629_23928 , \23630_23929 , \23631_23930 , \23632_23931 , \23633_23932 , \23634_23933 , \23635_23934 , \23636_23935 ,
         \23637_23936 , \23638_23937 , \23639_23938 , \23640_23939 , \23641_23940 , \23642_23941 , \23643_23942 , \23644_23943 , \23645_23944 , \23646_23945 ,
         \23647_23946 , \23648_23947 , \23649_23948 , \23650_23949 , \23651_23950 , \23652_23951 , \23653_23952 , \23654_23953 , \23655_23954 , \23656_23955 ,
         \23657_23956 , \23658_23957 , \23659_23958 , \23660_23959 , \23661_23960 , \23662_23961 , \23663_23962 , \23664_23963 , \23665_23964 , \23666_23965 ,
         \23667_23966 , \23668_23967 , \23669_23968 , \23670_23969 , \23671_23970 , \23672_23971 , \23673_23972 , \23674_23973 , \23675_23974 , \23676_23975 ,
         \23677_23976 , \23678_23977 , \23679_23978 , \23680_23979 , \23681_23980 , \23682_23981 , \23683_23982 , \23684_23983 , \23685_23984 , \23686_23985 ,
         \23687_23986 , \23688_23987 , \23689_23988 , \23690_23989 , \23691_23990 , \23692_23991 , \23693_23992 , \23694_23993 , \23695_23994 , \23696_23995 ,
         \23697_23996 , \23698_23997 , \23699_23998 , \23700_23999 , \23701_24000 , \23702 , \23703_24002 , \23704_24003 , \23705_24004 , \23706_24005 ,
         \23707_24006 , \23708_24007 , \23709_24008 , \23710_24009 , \23711_24010 , \23712_24011 , \23713_24012 , \23714_24013 , \23715_24014 , \23716_24015 ,
         \23717_24016 , \23718_24017 , \23719_24018 , \23720_24019 , \23721_24020 , \23722_24021 , \23723_24022 , \23724_24023 , \23725_24024 , \23726_24025 ,
         \23727_24026 , \23728_24027 , \23729_24028 , \23730_24029 , \23731_24030 , \23732_24031 , \23733_24032 , \23734_24033 , \23735_24034 , \23736_24035 ,
         \23737_24036 , \23738_24037 , \23739_24038 , \23740_24039 , \23741_24040 , \23742_24041 , \23743_24042 , \23744_24043 , \23745_24044 , \23746_24045 ,
         \23747_24046 , \23748_24047 , \23749_24048 , \23750_24049 , \23751_24050 , \23752_24051 , \23753_24052 , \23754_24053 , \23755_24054 , \23756_24055 ,
         \23757_24056 , \23758_24057 , \23759_24058 , \23760_24059 , \23761_24060 , \23762_24061 , \23763_24062 , \23764_24063 , \23765_24064 , \23766_24065 ,
         \23767_24066 , \23768_24067 , \23769_24068 , \23770_24069 , \23771_24070 , \23772_24071 , \23773_24072 , \23774_24073 , \23775_24074 , \23776_24075 ,
         \23777_24076 , \23778_24077 , \23779_24078 , \23780_24079 , \23781_24080 , \23782_24081 , \23783_24082 , \23784_24083 , \23785_24084 , \23786_24085 ,
         \23787_24086 , \23788_24087 , \23789_24088 , \23790_24089 , \23791_24090 , \23792_24091 , \23793_24092 , \23794_24093 , \23795_24094 , \23796_24095 ,
         \23797_24096 , \23798_24097 , \23799_24098 , \23800_24099 , \23801_24100 , \23802_24101 , \23803_24102 , \23804_24103 , \23805_24104 , \23806_24105 ,
         \23807_24106 , \23808_24107 , \23809_24108 , \23810_24109 , \23811_24110 , \23812_24111 , \23813_24112 , \23814_24113 , \23815_24114 , \23816_24115 ,
         \23817_24116 , \23818_24117 , \23819_24118 , \23820_24119 , \23821_24120 , \23822_24121 , \23823_24122 , \23824_24123 , \23825_24124 , \23826_24125 ,
         \23827_24126 , \23828_24127 , \23829_24128 , \23830_24129 , \23831_24130 , \23832_24131 , \23833_24132 , \23834 , \23835_24134_nG5b1c , \23836_24135 ,
         \23837_24136 , \23838_24137 , \23839_24138 , \23840_24139 , \23841_24140 , \23842_24141 , \23843_24142 , \23844_24143 , \23845_24144 , \23846_24145 ,
         \23847_24146 , \23848_24147 , \23849_24148 , \23850_24149 , \23851_24150 , \23852_24151 , \23853_24152 , \23854_24153 , \23855_24154 , \23856_24155 ,
         \23857_24156 , \23858_24157 , \23859_24158 , \23860_24159 , \23861_24160 , \23862_24161 , \23863_24162 , \23864_24163 , \23865_24164 , \23866_24165 ,
         \23867_24166 , \23868_24167 , \23869_24168 , \23870_24169 , \23871_24170 , \23872_24171 , \23873_24172 , \23874_24173 , \23875_24174 , \23876_24175 ,
         \23877_24176 , \23878_24177 , \23879_24178 , \23880_24179 , \23881_24180 , \23882_24181 , \23883_24182 , \23884_24183 , \23885_24184 , \23886_24185 ,
         \23887_24186 , \23888_24187 , \23889_24188 , \23890_24189 , \23891_24190 , \23892_24191 , \23893_24192 , \23894_24193 , \23895_24194 , \23896_24195 ,
         \23897 , \23898 , \23899_24198_nG65b8 , \23900_24199 , \23901_24200 , \23902_24201 , \23903_24202 , \23904_24203 , \23905_24204 , \23906_24205 ,
         \23907_24206 , \23908_24207 , \23909_24208 , \23910_24209 , \23911_24210 , \23912_24211 , \23913_24212 , \23914_24213 , \23915_24214 , \23916_24215 ,
         \23917_24216 , \23918_24217 , \23919_24218 , \23920_24219 , \23921_24220 , \23922_24221 , \23923_24222 , \23924_24223 , \23925_24224 , \23926_24225 ,
         \23927_24226_nG9bcf , \23928_24227 , \23929_24228 , \23930_24229 , \23931_24230 , \23932_24231 , \23933_24232 , \23934_24233 , \23935_24234 , \23936_24235 ,
         \23937_24236 , \23938_24237 , \23939_24238 , \23940_24239 , \23941_24240 , \23942_24241 , \23943_24242 , \23944_24243 , \23945_24244 , \23946_24245 ,
         \23947_24246 , \23948_24247 , \23949_24248 , \23950_24249 , \23951_24250 , \23952_24251 , \23953_24252 , \23954_24253 , \23955_24254 , \23956_24255 ,
         \23957_24256 , \23958_24257 , \23959_24258 , \23960_24259 , \23961_24260 , \23962_24261 , \23963_24262 , \23964_24263 , \23965_24264 , \23966_24265 ,
         \23967_24266 , \23968_24267 , \23969_24268 , \23970_24269 , \23971_24270 , \23972_24271 , \23973_24272 , \23974_24273 , \23975_24274 , \23976_24275 ,
         \23977_24276 , \23978_24277 , \23979_24278 , \23980_24279 , \23981_24280 , \23982_24281 , \23983_24282 , \23984_24283 , \23985_24284 , \23986_24285 ,
         \23987_24286 , \23988_24287 , \23989_24288 , \23990_24289 , \23991_24290 , \23992_24291 , \23993_24292 , \23994_24293 , \23995_24294 , \23996_24295 ,
         \23997_24296 , \23998_24297 , \23999_24298 , \24000_24299 , \24001_24300 , \24002_24301 , \24003_24302 , \24004_24303 , \24005_24304 , \24006_24305 ,
         \24007_24306 , \24008_24307 , \24009_24308 , \24010_24309 , \24011_24310 , \24012_24311 , \24013_24312 , \24014_24313 , \24015_24314 , \24016_24315 ,
         \24017_24316 , \24018_24317 , \24019_24318 , \24020_24319 , \24021_24320 , \24022_24321 , \24023_24322 , \24024_24323 , \24025_24324 , \24026_24325 ,
         \24027_24326 , \24028_24327 , \24029_24328 , \24030_24329 , \24031_24330 , \24032_24331 , \24033_24332 , \24034_24333 , \24035_24334 , \24036_24335 ,
         \24037_24336 , \24038_24337 , \24039_24338 , \24040_24339 , \24041_24340 , \24042_24341 , \24043_24342 , \24044_24343 , \24045_24344 , \24046_24345 ,
         \24047_24346 , \24048_24347 , \24049_24348 , \24050_24349 , \24051_24350 , \24052_24351 , \24053_24352 , \24054_24353 , \24055_24354 , \24056_24355 ,
         \24057_24356 , \24058_24357 , \24059_24358 , \24060_24359 , \24061_24360 , \24062_24361 , \24063_24362 , \24064_24363 , \24065_24364 , \24066_24365 ,
         \24067_24366 , \24068_24367 , \24069_24368 , \24070_24369 , \24071_24370 , \24072_24371 , \24073 , \24074_24373 , \24075_24374 , \24076_24375 ,
         \24077_24376 , \24078_24377 , \24079_24378 , \24080_24379 , \24081_24380 , \24082_24381 , \24083_24382 , \24084_24383 , \24085_24384 , \24086_24385 ,
         \24087_24386 , \24088_24387 , \24089_24388 , \24090_24389 , \24091_24390 , \24092_24391 , \24093_24392 , \24094_24393 , \24095_24394 , \24096_24395 ,
         \24097_24396 , \24098_24397 , \24099_24398 , \24100_24399 , \24101_24400 , \24102_24401 , \24103_24402 , \24104_24403 , \24105_24404 , \24106_24405 ,
         \24107_24406 , \24108_24407 , \24109_24408 , \24110_24409 , \24111_24410 , \24112_24411 , \24113_24412 , \24114_24413 , \24115_24414 , \24116_24415 ,
         \24117_24416 , \24118_24417 , \24119_24418 , \24120_24419 , \24121_24420 , \24122_24421 , \24123_24422 , \24124_24423 , \24125_24424 , \24126_24425 ,
         \24127_24426 , \24128_24427 , \24129_24428 , \24130_24429 , \24131_24430 , \24132_24431 , \24133_24432 , \24134_24433 , \24135_24434 , \24136_24435 ,
         \24137_24436 , \24138_24437 , \24139_24438 , \24140_24439 , \24141_24440 , \24142_24441 , \24143_24442 , \24144_24443 , \24145_24444 , \24146_24445 ,
         \24147_24446 , \24148_24447 , \24149_24448 , \24150_24449 , \24151_24450 , \24152_24451 , \24153_24452 , \24154_24453 , \24155_24454 , \24156_24455 ,
         \24157_24456 , \24158_24457 , \24159_24458 , \24160_24459 , \24161_24460 , \24162_24461 , \24163_24462 , \24164_24463 , \24165_24464 , \24166_24465 ,
         \24167_24466 , \24168_24467 , \24169_24468 , \24170_24469 , \24171_24470 , \24172_24471 , \24173_24472 , \24174_24473 , \24175_24474 , \24176_24475 ,
         \24177_24476 , \24178_24477 , \24179_24478 , \24180_24479 , \24181_24480 , \24182_24481 , \24183_24482 , \24184_24483 , \24185_24484 , \24186_24485 ,
         \24187_24486 , \24188_24487 , \24189_24488 , \24190_24489 , \24191_24490 , \24192_24491 , \24193_24492 , \24194_24493 , \24195_24494 , \24196_24495 ,
         \24197_24496 , \24198_24497 , \24199_24498 , \24200_24499 , \24201_24500 , \24202_24501 , \24203_24502 , \24204_24503 , \24205_24504 , \24206 ,
         \24207_24506 , \24208_24507 , \24209_24508 , \24210_24509 , \24211_24510 , \24212_24511 , \24213_24512 , \24214_24513 , \24215_24514 , \24216_24515 ,
         \24217_24516 , \24218_24517 , \24219_24518 , \24220_24519 , \24221_24520 , \24222_24521 , \24223_24522 , \24224_24523 , \24225_24524 , \24226_24525 ,
         \24227_24526 , \24228_24527 , \24229_24528 , \24230_24529 , \24231_24530 , \24232_24531 , \24233_24532 , \24234_24533 , \24235_24534 , \24236_24535 ,
         \24237_24536 , \24238_24537 , \24239_24538 , \24240_24539 , \24241_24540 , \24242_24541 , \24243_24542 , \24244_24543 , \24245_24544 , \24246_24545 ,
         \24247_24546 , \24248_24547 , \24249_24548 , \24250_24549 , \24251_24550 , \24252_24551 , \24253_24552 , \24254_24553 , \24255_24554 , \24256_24555 ,
         \24257_24556 , \24258_24557 , \24259_24558 , \24260_24559 , \24261_24560 , \24262_24561 , \24263_24562 , \24264_24563 , \24265_24564 , \24266_24565 ,
         \24267_24566 , \24268_24567 , \24269_24568 , \24270_24569 , \24271_24570 , \24272_24571 , \24273_24572 , \24274_24573 , \24275_24574 , \24276_24575 ,
         \24277_24576 , \24278_24577 , \24279_24578 , \24280_24579 , \24281_24580 , \24282_24581 , \24283_24582 , \24284_24583 , \24285_24584 , \24286_24585 ,
         \24287_24586 , \24288_24587 , \24289_24588 , \24290_24589 , \24291_24590 , \24292_24591 , \24293_24592 , \24294_24593 , \24295_24594 , \24296_24595 ,
         \24297_24596 , \24298_24597 , \24299_24598 , \24300_24599 , \24301_24600 , \24302_24601 , \24303_24602 , \24304_24603 , \24305_24604 , \24306_24605 ,
         \24307_24606 , \24308_24607 , \24309_24608 , \24310_24609 , \24311_24610 , \24312_24611 , \24313_24612 , \24314_24613 , \24315_24614 , \24316_24615 ,
         \24317_24616 , \24318_24617 , \24319_24618 , \24320_24619 , \24321_24620 , \24322_24621 , \24323_24622 , \24324_24623 , \24325_24624 , \24326_24625 ,
         \24327_24626 , \24328_24627 , \24329_24628 , \24330_24629 , \24331_24630 , \24332_24631 , \24333_24632 , \24334_24633 , \24335_24634 , \24336_24635 ,
         \24337_24636 , \24338_24637 , \24339_24638 , \24340 , \24341_24640 , \24342_24641 , \24343_24642 , \24344_24643 , \24345_24644 , \24346_24645 ,
         \24347_24646 , \24348_24647 , \24349_24648 , \24350_24649 , \24351_24650 , \24352_24651 , \24353_24652 , \24354_24653 , \24355_24654 , \24356_24655 ,
         \24357_24656 , \24358_24657 , \24359_24658 , \24360_24659 , \24361_24660 , \24362_24661 , \24363_24662 , \24364_24663 , \24365_24664 , \24366_24665 ,
         \24367_24666 , \24368_24667 , \24369_24668 , \24370_24669 , \24371_24670 , \24372_24671 , \24373_24672 , \24374_24673 , \24375_24674 , \24376_24675 ,
         \24377_24676 , \24378_24677 , \24379_24678 , \24380_24679 , \24381_24680 , \24382_24681 , \24383_24682 , \24384_24683 , \24385_24684 , \24386_24685 ,
         \24387_24686 , \24388_24687 , \24389_24688 , \24390_24689 , \24391_24690 , \24392_24691 , \24393_24692 , \24394_24693 , \24395_24694 , \24396_24695 ,
         \24397_24696 , \24398_24697 , \24399_24698 , \24400_24699 , \24401_24700 , \24402_24701 , \24403_24702 , \24404_24703 , \24405_24704 , \24406_24705 ,
         \24407_24706 , \24408_24707 , \24409_24708 , \24410_24709 , \24411_24710 , \24412_24711 , \24413_24712 , \24414_24713 , \24415_24714 , \24416_24715 ,
         \24417_24716 , \24418_24717 , \24419_24718 , \24420_24719 , \24421_24720 , \24422_24721 , \24423_24722 , \24424_24723 , \24425_24724 , \24426_24725 ,
         \24427_24726 , \24428_24727 , \24429_24728 , \24430_24729 , \24431_24730 , \24432_24731 , \24433_24732 , \24434_24733 , \24435_24734 , \24436_24735 ,
         \24437_24736 , \24438_24737 , \24439_24738 , \24440_24739 , \24441_24740 , \24442_24741 , \24443_24742 , \24444_24743 , \24445_24744 , \24446_24745 ,
         \24447_24746 , \24448_24747 , \24449_24748 , \24450_24749 , \24451_24750 , \24452_24751 , \24453_24752 , \24454_24753 , \24455_24754 , \24456_24755 ,
         \24457_24756 , \24458_24757 , \24459_24758 , \24460_24759 , \24461_24760 , \24462_24761 , \24463_24762 , \24464_24763 , \24465_24764 , \24466_24765 ,
         \24467_24766 , \24468_24767 , \24469_24768 , \24470_24769 , \24471_24770 , \24472_24771 , \24473 , \24474_24773 , \24475_24774 , \24476_24775 ,
         \24477_24776 , \24478_24777 , \24479_24778 , \24480_24779 , \24481_24780 , \24482_24781 , \24483_24782 , \24484_24783_nG4412 , \24485_24784 , \24486_24785 ,
         \24487_24786_nG4415 , \24488_24787 , \24489_24788 , \24490_24789 , \24491_24793 , \24492_24794 , \24493_24795 , \24494_24796 , \24495_24797 , \24496_24798 ,
         \24497_24799 , \24498_24800 , \24499_24801 , \24500_24802 , \24501_24803 , \24502_24804 , \24503_24805 , \24504_24806 , \24505_24807 , \24506_24808 ,
         \24507_24809 , \24508_24810 , \24509_24811 , \24510_24812 , \24511_24813 , \24512_24814 , \24513_24815 , \24514_24816 , \24515_24817 , \24516_24818 ,
         \24517_24819 , \24518_24820 , \24519_24821 , \24520_24822 , \24521_24823 , \24522_24824 , \24523_24825 , \24524_24826 , \24525_24827 , \24526_24828 ,
         \24527_24829 , \24528_24830 , \24529_24831 , \24530_24832 , \24531_24833 , \24532_24834 , \24533_24835 , \24534_24836 , \24535_24837 , \24536_24838 ,
         \24537_24839 , \24538_24840 , \24539_24841 , \24540_24842 , \24541_24843 , \24542_24844 , \24543_24845 , \24544_24846 , \24545_24847 , \24546_24848 ,
         \24547_24849 , \24548_24850 , \24549_24851 , \24550_24852 , \24551_24853 , \24552_24854 , \24553_24855 , \24554_24856 , \24555_24857 , \24556_24858 ,
         \24557_24859 , \24558_24860 , \24559_24861 , \24560_24862 , \24561_24863 , \24562_24864 , \24563_24865 , \24564_24866 , \24565_24867 , \24566_24868 ,
         \24567_24869 , \24568_24870 , \24569_24871 , \24570_24872 , \24571_24873 , \24572_24874 , \24573_24875 , \24574_24876 , \24575_24877 , \24576_24878 ,
         \24577_24879 , \24578_24880 , \24579_24881 , \24580_24882 , \24581_24883 , \24582_24884 , \24583_24885 , \24584_24886 , \24585_24887 , \24586_24888 ,
         \24587_24889 , \24588_24890 , \24589_24891 , \24590_24892 , \24591_24893 , \24592_24894 , \24593_24895 , \24594_24896 , \24595_24897 , \24596_24898 ,
         \24597_24899 , \24598_24900 , \24599_24901 , \24600_24902 , \24601_24903 , \24602_24904 , \24603_24905 , \24604_24906 , \24605_24907 , \24606_24908 ,
         \24607_24909 , \24608_24910 , \24609_24911 , \24610_24912 , \24611_24913 , \24612_24914 , \24613_24915 , \24614_24916 , \24615_24917 , \24616_24918 ,
         \24617_24919 , \24618_24920 , \24619_24921 , \24620_24922 , \24621_24923 , \24622_24924 , \24623_24925 , \24624_24926 , \24625_24927 , \24626_24928 ,
         \24627_24929 , \24628_24930 , \24629_24931 , \24630_24932 , \24631_24933 , \24632_24934 , \24633_24935 , \24634_24936 , \24635_24937 , \24636_24938 ,
         \24637_24939 , \24638_24940 , \24639_24941 , \24640_24942 , \24641_24943 , \24642_24944 , \24643_24945 , \24644_24946 , \24645_24947 , \24646_24948 ,
         \24647_24949 , \24648_24950 , \24649_24951 , \24650_24952 , \24651_24953 , \24652_24954 , \24653_24955 , \24654_24956 , \24655_24957 , \24656_24958 ,
         \24657_24959 , \24658_24960 , \24659_24961 , \24660_24962 , \24661_24963 , \24662_24964 , \24663_24965 , \24664_24966 , \24665_24967 , \24666_24968 ,
         \24667_24969 , \24668_24970 , \24669_24971 , \24670_24972 , \24671_24973 , \24672_24974 , \24673_24975 , \24674_24976 , \24675_24977 , \24676_24978 ,
         \24677_24979 , \24678_24980 , \24679_24981 , \24680_24982 , \24681_24983 , \24682_24984 , \24683_24985 , \24684_24986 , \24685_24987 , \24686_24988 ,
         \24687_24989 , \24688_24990 , \24689_24991 , \24690_24992 , \24691_24993 , \24692_24994 , \24693_24995 , \24694_24996 , \24695_24997 , \24696_24998 ,
         \24697_24999 , \24698_25000 , \24699_25001 , \24700_25002 , \24701_25003 , \24702_25004 , \24703_25005 , \24704_25006 , \24705_25007 , \24706_25008 ,
         \24707_25009 , \24708_25010 , \24709_25011 , \24710_25012 , \24711_25013 , \24712_25014 , \24713_25015 , \24714_25016 , \24715_25017 , \24716_25018 ,
         \24717_25019 , \24718_25020 , \24719_25021 , \24720_25022 , \24721_25023 , \24722_25024 , \24723_25025 , \24724_25026 , \24725_25027 , \24726_25028 ,
         \24727_25029 , \24728_25030 , \24729_25031 , \24730_25032 , \24731_25033 , \24732_25034 , \24733_25035 , \24734_25036 , \24735_25037 , \24736_25038 ,
         \24737_25039 , \24738_25040 , \24739_25041 , \24740_25042 , \24741_25043 , \24742_25044 , \24743_25045 , \24744_25046 , \24745_25047 , \24746_25048 ,
         \24747_25049 , \24748_25050 , \24749_25051 , \24750_25052 , \24751_25053 , \24752_25054 , \24753_25055 , \24754_25056 , \24755_25057 , \24756_25058 ,
         \24757_25059 , \24758_25060 , \24759_25061 , \24760_25062 , \24761_25063 , \24762_25064 , \24763_25065 , \24764_25066 , \24765_25067 , \24766_25068 ,
         \24767_25069 , \24768_25070 , \24769_25071 , \24770_25072 , \24771_25073 , \24772_25074 , \24773_25075 , \24774_25076 , \24775_25077 , \24776_25078 ,
         \24777_25079 , \24778_25080 , \24779_25081 , \24780_25082 , \24781_25083 , \24782_25084 , \24783_25085 , \24784_25086 , \24785_25087 , \24786_25088 ,
         \24787_25089 , \24788_25090 , \24789_25091 , \24790_25092 , \24791_25093 , \24792_25094 , \24793_25095 , \24794_25096 , \24795_25097 , \24796_25098 ,
         \24797_25099 , \24798_25100 , \24799_25101 , \24800_25102 , \24801_25103 , \24802_25104 , \24803_25105 , \24804_25106 , \24805_25107 , \24806_25108 ,
         \24807_25109 , \24808_25110 , \24809_25111 , \24810_25112 , \24811_25113 , \24812_25114 , \24813_25115 , \24814_25116 , \24815_25117 , \24816_25118 ,
         \24817_25119 , \24818_25120 , \24819_25121 , \24820_25122 , \24821_25123 , \24822_25124 , \24823_25125 , \24824_25126 , \24825_25127 , \24826_25128 ,
         \24827 , \24828_25130 , \24829_25131 , \24830_25132 , \24831_25133 , \24832_25134 , \24833_25135 , \24834_25136 , \24835_25137 , \24836_25138 ,
         \24837_25139 , \24838_25140 , \24839_25141 , \24840_25142 , \24841_25143 , \24842_25144 , \24843_25145 , \24844_25146 , \24845_25147 , \24846_25148 ,
         \24847_25149 , \24848_25150 , \24849_25151 , \24850_25152 , \24851_25153 , \24852_25154 , \24853_25155 , \24854_25156 , \24855_25157 , \24856_25158 ,
         \24857_25159 , \24858_25160 , \24859_25161 , \24860_25162 , \24861_25163 , \24862_25164 , \24863_25165 , \24864_25166 , \24865_25167 , \24866_25168 ,
         \24867_25169 , \24868_25170 , \24869_25171 , \24870_25172 , \24871_25173 , \24872_25174 , \24873_25175 , \24874_25176 , \24875_25177 , \24876_25178 ,
         \24877_25179 , \24878_25180 , \24879_25181 , \24880_25182 , \24881_25183 , \24882_25184 , \24883_25185 , \24884_25186 , \24885_25187 , \24886_25188 ,
         \24887_25189 , \24888_25190 , \24889_25191 , \24890_25192 , \24891_25193 , \24892_25194 , \24893_25195 , \24894_25196 , \24895_25197 , \24896_25198 ,
         \24897_25199 , \24898_25200 , \24899_25201 , \24900_25202 , \24901_25203 , \24902_25204 , \24903_25205 , \24904_25206 , \24905_25207 , \24906_25208 ,
         \24907_25209 , \24908_25210 , \24909_25211 , \24910_25212 , \24911_25213 , \24912_25214 , \24913_25215 , \24914_25216 , \24915_25217 , \24916_25218 ,
         \24917_25219 , \24918_25220 , \24919_25221 , \24920_25222 , \24921_25223 , \24922_25224 , \24923_25225 , \24924_25226 , \24925_25227 , \24926_25228 ,
         \24927_25229 , \24928_25230 , \24929_25231 , \24930_25232 , \24931_25233 , \24932_25234 , \24933_25235 , \24934_25236 , \24935_25237 , \24936_25238 ,
         \24937_25239 , \24938_25240 , \24939_25241 , \24940_25242 , \24941_25243 , \24942_25244 , \24943_25245 , \24944_25246 , \24945_25247 , \24946_25248 ,
         \24947_25249 , \24948_25250 , \24949_25251 , \24950_25252 , \24951_25253 , \24952_25254 , \24953_25255 , \24954_25256 , \24955_25257 , \24956_25258 ,
         \24957_25259 , \24958_25260 , \24959 , \24960_25262_nG5c25 , \24961_25263 , \24962_25264 , \24963_25265 , \24964_25266 , \24965_25267 , \24966_25268 ,
         \24967 , \24968 , \24969_25271_nG65bb , \24970_25272 , \24971_25273 , \24972_25274 , \24973_25275 , \24974_25276 , \24975_25277 , \24976_25278 ,
         \24977_25279 , \24978_25280 , \24979_25281 , \24980_25282 , \24981_25283 , \24982_25284 , \24983_25285 , \24984_25286 , \24985_25287 , \24986_25288 ,
         \24987_25289 , \24988_25290 , \24989_25291 , \24990_25292 , \24991_25293 , \24992_25294 , \24993_25295 , \24994_25296 , \24995_25297 , \24996_25298_nG9bcc ,
         \24997_25299 , \24998_25300 , \24999_25301 , \25000_25302 , \25001_25303 , \25002_25304 , \25003_25305 , \25004_25306 , \25005_25307 , \25006_25308 ,
         \25007_25309 , \25008_25310 , \25009_25311 , \25010_25312 , \25011_25313 , \25012_25314 , \25013_25315 , \25014_25316 , \25015_25317 , \25016_25318 ,
         \25017_25319 , \25018_25320 , \25019_25321 , \25020_25322 , \25021_25323 , \25022_25324 , \25023_25325 , \25024_25326 , \25025_25327 , \25026_25328 ,
         \25027_25329 , \25028_25330 , \25029_25331 , \25030_25332 , \25031_25333 , \25032_25334 , \25033_25335 , \25034_25336 , \25035_25337 , \25036_25338 ,
         \25037_25339 , \25038_25340 , \25039_25341 , \25040_25342 , \25041_25343 , \25042_24790 , \25043_24791 , \25044_24792 , \25045_25344 , \25046_25345 ,
         \25047_25346 , \25048_25347 , \25049_25348 , \25050_25349 , \25051_25350 , \25052_25351 , \25053_25352 , \25054_25353 , \25055_25354 , \25056_25355 ,
         \25057_25356 , \25058_25357 , \25059_25358 , \25060_25359 , \25061_25360 , \25062_25361 , \25063_25362 , \25064_25363 , \25065_25364 , \25066_25365 ,
         \25067_25366 , \25068_25367 , \25069_25368 , \25070_25369 , \25071_25370 , \25072_25371 , \25073_25372 , \25074_25373 , \25075_25374 , \25076_25375 ,
         \25077_25376 , \25078_25377 , \25079_25378 , \25080_25379 , \25081_25380 , \25082_25381 , \25083_25382 , \25084_25383 , \25085_25384 , \25086_25385 ,
         \25087_25386 , \25088_25387 , \25089_25388 , \25090_25389 , \25091_25390 , \25092_25391 , \25093_25392 , \25094_25393 , \25095_25394 , \25096_25395 ,
         \25097_25396 , \25098_25397 , \25099_25398 , \25100_25399 , \25101_25400 , \25102_25401 , \25103_25402 , \25104_25403 , \25105_25404 , \25106_25405 ,
         \25107_25406 , \25108_25407 , \25109_25408 , \25110_25409 , \25111_25410 , \25112_25411 , \25113_25412 , \25114_25413 , \25115_25414 , \25116_25415 ,
         \25117_25416 , \25118_25417 , \25119_25418 , \25120_25419 , \25121_25420 , \25122_25421 , \25123_25422 , \25124_25423 , \25125_25424 , \25126_25425 ,
         \25127_25426 , \25128_25427 , \25129_25428 , \25130_25429 , \25131_25430 , \25132_25431 , \25133_25432 , \25134_25433 , \25135_25434 , \25136_25435 ,
         \25137_25436 , \25138_25437 , \25139_25438 , \25140_25439 , \25141_25440 , \25142_25441 , \25143_25442 , \25144_25443 , \25145_25444 , \25146_25445 ,
         \25147_25446 , \25148_25447 , \25149_25448 , \25150_25449 , \25151_25450 , \25152_25451 , \25153_25452 , \25154_25453 , \25155_25454 , \25156_25455 ,
         \25157_25456 , \25158_25457 , \25159_25458 , \25160_25459 , \25161_25460 , \25162_25461 , \25163_25462 , \25164_25463 , \25165_25464 , \25166_25465 ,
         \25167_25466 , \25168_25467 , \25169_25468 , \25170_25469 , \25171_25470 , \25172_25471 , \25173_25472 , \25174_25473 , \25175_25474 , \25176_25475 ,
         \25177_25476 , \25178_25477 , \25179_25478 , \25180_25479 , \25181_25480 , \25182_25481 , \25183_25482 , \25184_25483 , \25185_25484 , \25186_25485 ,
         \25187_25486 , \25188_25487 , \25189_25488 , \25190_25489 , \25191_25490 , \25192_25491 , \25193_25492 , \25194_25493 , \25195_25494 , \25196_25495 ,
         \25197_25496 , \25198_25497 , \25199_25498 , \25200_25499 , \25201_25500 , \25202_25501 , \25203_25502 , \25204_25503 , \25205_25504 , \25206_25505 ,
         \25207_25506 , \25208_25507 , \25209_25508 , \25210_25509 , \25211_25510 , \25212_25511 , \25213_25512 , \25214_25513 , \25215_25514 , \25216_25515 ,
         \25217_25516 , \25218_25517 , \25219_25518 , \25220_25519 , \25221_25520 , \25222_25521 , \25223_25522 , \25224_25523 , \25225_25524 , \25226_25525 ,
         \25227_25526 , \25228_25527 , \25229_25528 , \25230_25529 , \25231_25530 , \25232_25531 , \25233_25532 , \25234_25533 , \25235_25534 , \25236_25535 ,
         \25237_25536 , \25238_25537 , \25239_25538 , \25240_25539 , \25241_25540 , \25242_25541 , \25243_25542 , \25244_25543 , \25245_25544 , \25246_25545 ,
         \25247_25546 , \25248_25547 , \25249_25548 , \25250_25549 , \25251_25550 , \25252_25551 , \25253_25552 , \25254_25553 , \25255_25554 , \25256_25555 ,
         \25257_25556 , \25258_25557 , \25259_25558 , \25260_25559 , \25261_25560 , \25262_25561 , \25263_25562 , \25264_25563 , \25265_25564 , \25266_25565 ,
         \25267_25566 , \25268_25567 , \25269_25568 , \25270_25569 , \25271_25570 , \25272_25571 , \25273_25572 , \25274_25573 , \25275_25574 , \25276_25575 ,
         \25277_25576 , \25278_25577 , \25279_25578 , \25280_25579 , \25281_25580 , \25282_25581 , \25283_25582 , \25284_25583 , \25285_25584 , \25286_25585 ,
         \25287_25586 , \25288_25587 , \25289_25588 , \25290_25589 , \25291_25590 , \25292_25591 , \25293_25592 , \25294_25593 , \25295_25594 , \25296_25595 ,
         \25297_25596 , \25298_25597 , \25299_25598 , \25300_25599 , \25301_25600 , \25302_25601 , \25303_25602 , \25304_25603 , \25305_25604 , \25306_25605 ,
         \25307_25606 , \25308_25607 , \25309_25608 , \25310_25609 , \25311_25610 , \25312_25611 , \25313_25612 , \25314_25613 , \25315_25614 , \25316_25615 ,
         \25317_25616 , \25318_25617 , \25319_25618 , \25320_25619 , \25321_25620 , \25322_25621 , \25323_25622 , \25324_25623 , \25325_25624 , \25326_25625 ,
         \25327_25626 , \25328_25627 , \25329_25628 , \25330_25629 , \25331_25630 , \25332_25631 , \25333_25632 , \25334_25633 , \25335_25634 , \25336_25635 ,
         \25337 , \25338_25637 , \25339_25638 , \25340_25639 , \25341_25640 , \25342_25641 , \25343_25642 , \25344_25643 , \25345_25644 , \25346_25645 ,
         \25347_25646 , \25348_25647 , \25349_25648 , \25350_25649 , \25351_25650 , \25352_25651 , \25353_25652 , \25354_25653 , \25355_25654 , \25356_25655 ,
         \25357_25656 , \25358_25657 , \25359_25658 , \25360_25659 , \25361_25660 , \25362_25661 , \25363_25662 , \25364_25663 , \25365_25664 , \25366_25665 ,
         \25367_25666 , \25368_25667 , \25369_25668 , \25370_25669 , \25371_25670 , \25372_25671 , \25373_25672 , \25374_25673 , \25375_25674 , \25376_25675 ,
         \25377_25676 , \25378_25677 , \25379_25678 , \25380_25679 , \25381_25680 , \25382_25681 , \25383_25682 , \25384_25683 , \25385_25684 , \25386_25685 ,
         \25387_25686 , \25388_25687 , \25389_25688 , \25390_25689 , \25391_25690 , \25392_25691 , \25393_25692 , \25394_25693 , \25395_25694 , \25396_25695 ,
         \25397_25696 , \25398_25697 , \25399_25698 , \25400_25699 , \25401_25700 , \25402_25701 , \25403_25702 , \25404_25703 , \25405_25704 , \25406_25705 ,
         \25407_25706 , \25408_25707 , \25409_25708 , \25410_25709 , \25411_25710 , \25412_25711 , \25413_25712 , \25414_25713 , \25415_25714 , \25416_25715 ,
         \25417_25716 , \25418_25717 , \25419_25718 , \25420_25719 , \25421_25720 , \25422_25721 , \25423_25722 , \25424_25723 , \25425_25724 , \25426_25725 ,
         \25427_25726 , \25428_25727 , \25429_25728 , \25430_25729 , \25431_25730 , \25432_25731 , \25433_25732 , \25434_25733 , \25435_25734 , \25436_25735 ,
         \25437_25736 , \25438_25737 , \25439_25738 , \25440_25739 , \25441_25740 , \25442_25741 , \25443_25742 , \25444_25743 , \25445_25744 , \25446_25745 ,
         \25447_25746 , \25448_25747 , \25449_25748 , \25450_25749 , \25451_25750 , \25452_25751 , \25453_25752 , \25454_25753 , \25455_25754 , \25456_25755 ,
         \25457_25756 , \25458_25757 , \25459_25758 , \25460_25759 , \25461_25760 , \25462_25761 , \25463_25762 , \25464_25763 , \25465_25764 , \25466_25765 ,
         \25467_25766 , \25468_25767 , \25469 , \25470_25769_nG5d2e , \25471_25770 , \25472_25771 , \25473_25772 , \25474_25773 , \25475_25774 , \25476_25775 ,
         \25477_25776 , \25478_25777 , \25479_25778 , \25480_25779 , \25481_25780 , \25482_25781 , \25483_25782 , \25484_25783 , \25485_25784 , \25486_25785 ,
         \25487_25786 , \25488_25787 , \25489_25788 , \25490_25789 , \25491_25790 , \25492_25791 , \25493_25792 , \25494_25793 , \25495_25794 , \25496_25795 ,
         \25497_25796 , \25498_25797 , \25499_25798 , \25500_25799 , \25501_25800 , \25502_25801 , \25503_25802 , \25504_25803 , \25505_25804 , \25506_25805 ,
         \25507_25806 , \25508_25807 , \25509_25808 , \25510_25809 , \25511_25810 , \25512_25811 , \25513 , \25514 , \25515_25814_nG65be , \25516_25815 ,
         \25517_25816 , \25518_25817 , \25519_25818 , \25520_25819 , \25521_25820 , \25522_25821 , \25523_25822 , \25524_25823 , \25525_25824 , \25526_25825 ,
         \25527_25826 , \25528_25827 , \25529_25828 , \25530_25829 , \25531_25830 , \25532_25831 , \25533_25832 , \25534_25833 , \25535_25834 , \25536_25835 ,
         \25537_25836 , \25538_25837 , \25539_25838 , \25540_25839 , \25541_25840 , \25542_25841 , \25543_25842 , \25544_25843 , \25545_25844 , \25546_25845 ,
         \25547_25846 , \25548_25847 , \25549_25848 , \25550_25849 , \25551_25850 , \25552_25851 , \25553_25852 , \25554_25853 , \25555_25854 , \25556_25855 ,
         \25557_25856 , \25558_25857 , \25559_25858 , \25560_25859 , \25561_25860_nG9bc9 , \25562_25861 , \25563_25862 , \25564_25863 , \25565_25864 , \25566_25865 ,
         \25567_25866 , \25568_25867 , \25569_25868 , \25570_25869 , \25571_25870 , \25572_25871 , \25573_25872 , \25574_25873 , \25575_25874 , \25576_25875 ,
         \25577_25876 , \25578_25877 , \25579_25878 , \25580_25879 , \25581_25880 , \25582_25881 , \25583_25882 , \25584_25883 , \25585_25884 , \25586_25885 ,
         \25587_25886 , \25588_25887 , \25589_25888 , \25590_25889 , \25591_25890 , \25592_25891 , \25593_25892 , \25594_25893 , \25595_25894 , \25596_25895 ,
         \25597_25896 , \25598_25897 , \25599_25898 , \25600_25899 , \25601_25900 , \25602_25901 , \25603_25902 , \25604_25903 , \25605_25904 , \25606_25905 ,
         \25607_25906 , \25608_25907 , \25609_25908 , \25610_25909 , \25611_25910 , \25612_25911 , \25613_25912 , \25614_25913 , \25615_25914 , \25616_25915 ,
         \25617_25916 , \25618_25917 , \25619_25918 , \25620_25919 , \25621_25920 , \25622_25921 , \25623_25922 , \25624_25923 , \25625_25924 , \25626_25925 ,
         \25627_25926 , \25628_25927 , \25629_25928 , \25630_25929 , \25631_25930 , \25632_25931 , \25633_25932 , \25634_25933 , \25635_25934 , \25636_25935 ,
         \25637_25936 , \25638_25937 , \25639_25938 , \25640_25939 , \25641_25940 , \25642_25941 , \25643_25942 , \25644_25943 , \25645_25944 , \25646_25945 ,
         \25647_25946 , \25648_25947 , \25649_25948 , \25650_25949 , \25651_25950 , \25652_25951 , \25653_25952 , \25654_25953 , \25655_25954 , \25656_25955 ,
         \25657_25956 , \25658_25957 , \25659_25958 , \25660_25959 , \25661_25960 , \25662_25961 , \25663_25962 , \25664_25963 , \25665_25964 , \25666_25965 ,
         \25667_25966 , \25668_25967 , \25669_25968 , \25670_25969 , \25671_25970 , \25672_25971 , \25673_25972 , \25674_25973 , \25675_25974 , \25676_25975 ,
         \25677_25976 , \25678_25977 , \25679_25978 , \25680_25979 , \25681_25980 , \25682_25981 , \25683_25982 , \25684_25983 , \25685_25984 , \25686_25985 ,
         \25687_25986 , \25688_25987 , \25689_25988 , \25690_25989 , \25691_25990 , \25692_25991 , \25693_25992 , \25694_25993 , \25695_25994 , \25696_25995 ,
         \25697_25996 , \25698_25997 , \25699_25998 , \25700_25999 , \25701_26000 , \25702_26001 , \25703_26002 , \25704_26003 , \25705_26004 , \25706_26005 ,
         \25707_26006 , \25708_26007 , \25709_26008 , \25710_26009 , \25711_26010 , \25712 , \25713_26012 , \25714_26013 , \25715_26014 , \25716_26015 ,
         \25717_26016 , \25718_26017 , \25719_26018 , \25720_26019 , \25721_26020 , \25722_26021 , \25723_26022 , \25724_26023 , \25725_26024 , \25726_26025 ,
         \25727_26026 , \25728_26027 , \25729_26028 , \25730_26029 , \25731_26030 , \25732_26031 , \25733_26032 , \25734_26033 , \25735_26034 , \25736_26035 ,
         \25737_26036 , \25738_26037 , \25739_26038 , \25740_26039 , \25741_26040 , \25742_26041 , \25743_26042 , \25744_26043 , \25745_26044 , \25746_26045 ,
         \25747_26046 , \25748_26047 , \25749_26048 , \25750_26049 , \25751_26050 , \25752_26051 , \25753_26052 , \25754_26053 , \25755_26054 , \25756_26055 ,
         \25757_26056 , \25758_26057 , \25759_26058 , \25760_26059 , \25761_26060 , \25762_26061 , \25763_26062 , \25764_26063 , \25765_26064 , \25766_26065 ,
         \25767_26066 , \25768_26067 , \25769_26068 , \25770_26069 , \25771_26070 , \25772_26071 , \25773_26072 , \25774_26073 , \25775_26074 , \25776_26075 ,
         \25777_26076 , \25778_26077 , \25779_26078 , \25780_26079 , \25781_26080 , \25782_26081 , \25783_26082 , \25784_26083 , \25785_26084 , \25786_26085 ,
         \25787_26086 , \25788_26087 , \25789_26088 , \25790_26089 , \25791_26090 , \25792_26091 , \25793_26092 , \25794_26093 , \25795_26094 , \25796_26095 ,
         \25797_26096 , \25798_26097 , \25799_26098 , \25800_26099 , \25801_26100 , \25802_26101 , \25803_26102 , \25804_26103 , \25805_26104 , \25806_26105 ,
         \25807_26106 , \25808_26107 , \25809_26108 , \25810_26109 , \25811_26110 , \25812_26111 , \25813_26112 , \25814_26113 , \25815_26114 , \25816_26115 ,
         \25817_26116 , \25818_26117 , \25819_26118 , \25820_26119 , \25821_26120 , \25822_26121 , \25823_26122 , \25824_26123 , \25825_26124 , \25826_26125 ,
         \25827_26126 , \25828_26127 , \25829_26128 , \25830_26129 , \25831_26130 , \25832_26131 , \25833_26132 , \25834_26133 , \25835_26134 , \25836_26135 ,
         \25837_26136 , \25838_26137 , \25839_26138 , \25840_26139 , \25841_26140 , \25842_26141 , \25843_26142 , \25844_26143 , \25845 , \25846_26145 ,
         \25847_26146 , \25848_26147 , \25849_26148 , \25850_26149 , \25851_26150 , \25852_26151 , \25853_26152 , \25854_26153 , \25855_26154 , \25856_26155 ,
         \25857_26156 , \25858_26157 , \25859_26158 , \25860_26159 , \25861_26160 , \25862_26161 , \25863_26162 , \25864_26163 , \25865_26164 , \25866_26165 ,
         \25867_26166 , \25868_26167 , \25869_26168 , \25870_26169 , \25871_26170 , \25872_26171 , \25873_26172 , \25874_26173 , \25875_26174 , \25876_26175 ,
         \25877_26176 , \25878_26177 , \25879_26178 , \25880_26179 , \25881_26180 , \25882_26181 , \25883_26182 , \25884_26183 , \25885_26184 , \25886_26185 ,
         \25887_26186 , \25888_26187 , \25889_26188 , \25890_26189 , \25891_26190 , \25892_26191 , \25893_26192 , \25894_26193 , \25895_26194 , \25896_26195 ,
         \25897_26196 , \25898_26197 , \25899_26198 , \25900_26199 , \25901_26200 , \25902_26201 , \25903_26202 , \25904_26203 , \25905_26204 , \25906_26205 ,
         \25907_26206 , \25908_26207 , \25909_26208 , \25910_26209 , \25911_26210 , \25912_26211 , \25913_26212 , \25914_26213 , \25915_26214 , \25916_26215 ,
         \25917_26216 , \25918_26217 , \25919_26218 , \25920_26219 , \25921_26220 , \25922_26221 , \25923_26222 , \25924_26223 , \25925_26224 , \25926_26225 ,
         \25927_26226 , \25928_26227 , \25929_26228 , \25930_26229 , \25931_26230 , \25932_26231 , \25933_26232 , \25934_26233 , \25935_26234 , \25936_26235 ,
         \25937_26236 , \25938_26237 , \25939_26238 , \25940_26239 , \25941_26240 , \25942_26241 , \25943_26242 , \25944_26243 , \25945_26244 , \25946_26245 ,
         \25947_26246 , \25948_26247 , \25949_26248 , \25950_26249 , \25951_26250 , \25952_26251 , \25953_26252 , \25954_26253 , \25955_26254 , \25956_26255 ,
         \25957_26256 , \25958_26257 , \25959_26258 , \25960_26259 , \25961_26260 , \25962_26261 , \25963_26262 , \25964_26263 , \25965_26264 , \25966_26265 ,
         \25967_26266 , \25968_26267 , \25969_26268 , \25970_26269 , \25971_26270 , \25972_26271 , \25973_26272 , \25974_26273 , \25975_26274 , \25976_26275 ,
         \25977_26276 , \25978_26277 , \25979 , \25980_26279 , \25981_26280 , \25982_26281 , \25983_26282 , \25984_26283 , \25985_26284 , \25986_26285 ,
         \25987_26286 , \25988_26287 , \25989_26288 , \25990_26289 , \25991_26290 , \25992_26291 , \25993_26292 , \25994_26293 , \25995_26294 , \25996_26295 ,
         \25997_26296 , \25998_26297 , \25999_26298 , \26000_26299 , \26001_26300 , \26002_26301 , \26003_26302 , \26004_26303 , \26005_26304 , \26006_26305 ,
         \26007_26306 , \26008_26307 , \26009_26308 , \26010_26309 , \26011_26310 , \26012_26311 , \26013_26312 , \26014_26313 , \26015_26314 , \26016_26315 ,
         \26017_26316 , \26018_26317 , \26019_26318 , \26020_26319 , \26021_26320 , \26022_26321 , \26023_26322 , \26024_26323 , \26025_26324 , \26026_26325 ,
         \26027_26326 , \26028_26327 , \26029_26328 , \26030_26329 , \26031_26330 , \26032_26331 , \26033_26332 , \26034_26333 , \26035_26334 , \26036_26335 ,
         \26037_26336 , \26038_26337 , \26039_26338 , \26040_26339 , \26041_26340 , \26042_26341 , \26043_26342 , \26044_26343 , \26045_26344 , \26046_26345 ,
         \26047_26346 , \26048_26347 , \26049_26348 , \26050_26349 , \26051_26350 , \26052_26351 , \26053_26352 , \26054_26353 , \26055_26354 , \26056_26355 ,
         \26057_26356 , \26058_26357 , \26059_26358 , \26060_26359 , \26061_26360 , \26062_26361 , \26063_26362 , \26064_26363 , \26065_26364 , \26066_26365 ,
         \26067_26366 , \26068_26367 , \26069_26368 , \26070_26369 , \26071_26370 , \26072_26371 , \26073_26372 , \26074_26373 , \26075_26374 , \26076_26375 ,
         \26077_26376 , \26078_26377 , \26079_26378 , \26080_26379 , \26081_26380 , \26082_26381 , \26083_26382 , \26084_26383 , \26085_26384 , \26086_26385 ,
         \26087_26386 , \26088_26387 , \26089_26388 , \26090_26389 , \26091_26390 , \26092_26391 , \26093_26392 , \26094_26393 , \26095_26394 , \26096_26395 ,
         \26097_26396 , \26098_26397 , \26099_26398 , \26100_26399 , \26101_26400 , \26102_26401 , \26103_26402 , \26104_26403 , \26105_26404 , \26106_26405 ,
         \26107_26406 , \26108_26407 , \26109_26408 , \26110_26409 , \26111_26410 , \26112 , \26113_26412 , \26114_26413 , \26115_26414 , \26116_26415 ,
         \26117_26416 , \26118_26417 , \26119_26418 , \26120_26419 , \26121_26420 , \26122_26421 , \26123_26422_nG440c , \26124_26423 , \26125_26424 , \26126_26425_nG440f ,
         \26127_26426 , \26128_26427 , \26129_26428 , \26130_26432 , \26131_26433 , \26132_26434 , \26133_26435 , \26134_26436 , \26135_26437 , \26136_26438 ,
         \26137_26439 , \26138_26440 , \26139_26441 , \26140_26442 , \26141_26443 , \26142_26444 , \26143_26445 , \26144_26446 , \26145_26447 , \26146_26448 ,
         \26147_26449 , \26148_26450 , \26149_26451 , \26150_26452 , \26151_26453 , \26152_26454 , \26153_26455 , \26154_26456 , \26155_26457 , \26156_26458 ,
         \26157_26459 , \26158_26460 , \26159_26461 , \26160_26462 , \26161_26463 , \26162_26464 , \26163_26465 , \26164_26466 , \26165_26467 , \26166_26468 ,
         \26167_26469 , \26168_26470 , \26169_26471 , \26170_26472 , \26171_26473 , \26172_26474 , \26173_26475 , \26174_26476 , \26175_26477 , \26176_26478 ,
         \26177_26479 , \26178_26480 , \26179_26481 , \26180_26482 , \26181_26483 , \26182_26484 , \26183_26485 , \26184_26486 , \26185_26487 , \26186_26488 ,
         \26187_26489 , \26188_26490 , \26189_26491 , \26190_26492 , \26191_26493 , \26192_26494 , \26193_26495 , \26194_26496 , \26195_26497 , \26196_26498 ,
         \26197_26499 , \26198_26500 , \26199_26501 , \26200_26502 , \26201_26503 , \26202_26504 , \26203_26505 , \26204_26506 , \26205_26507 , \26206_26508 ,
         \26207_26509 , \26208_26510 , \26209_26511 , \26210_26512 , \26211_26513 , \26212_26514 , \26213_26515 , \26214_26516 , \26215_26517 , \26216_26518 ,
         \26217_26519 , \26218_26520 , \26219_26521 , \26220_26522 , \26221_26523 , \26222_26524 , \26223_26525 , \26224_26526 , \26225_26527 , \26226_26528 ,
         \26227_26529 , \26228_26530 , \26229_26531 , \26230_26532 , \26231_26533 , \26232_26534 , \26233_26535 , \26234_26536 , \26235_26537 , \26236_26538 ,
         \26237_26539 , \26238_26540 , \26239_26541 , \26240_26542 , \26241_26543 , \26242_26544 , \26243_26545 , \26244_26546 , \26245_26547 , \26246_26548 ,
         \26247_26549 , \26248_26550 , \26249_26551 , \26250_26552 , \26251_26553 , \26252_26554 , \26253_26555 , \26254_26556 , \26255_26557 , \26256_26558 ,
         \26257_26559 , \26258_26560 , \26259_26561 , \26260_26562 , \26261_26563 , \26262_26564 , \26263_26565 , \26264_26566 , \26265_26567 , \26266_26568 ,
         \26267_26569 , \26268_26570 , \26269_26571 , \26270_26572 , \26271_26573 , \26272_26574 , \26273_26575 , \26274_26576 , \26275_26577 , \26276_26578 ,
         \26277_26579 , \26278_26580 , \26279_26581 , \26280_26582 , \26281_26583 , \26282_26584 , \26283_26585 , \26284_26586 , \26285_26587 , \26286_26588 ,
         \26287_26589 , \26288_26590 , \26289_26591 , \26290_26592 , \26291_26593 , \26292_26594 , \26293_26595 , \26294_26596 , \26295_26597 , \26296_26598 ,
         \26297_26599 , \26298_26600 , \26299_26601 , \26300_26602 , \26301_26603 , \26302_26604 , \26303_26605 , \26304_26606 , \26305_26607 , \26306_26608 ,
         \26307_26609 , \26308_26610 , \26309_26611 , \26310_26612 , \26311_26613 , \26312_26614 , \26313_26615 , \26314_26616 , \26315_26617 , \26316_26618 ,
         \26317_26619 , \26318_26620 , \26319_26621 , \26320_26622 , \26321_26623 , \26322_26624 , \26323_26625 , \26324_26626 , \26325_26627 , \26326_26628 ,
         \26327_26629 , \26328_26630 , \26329_26631 , \26330_26632 , \26331_26633 , \26332_26634 , \26333_26635 , \26334_26636 , \26335_26637 , \26336_26638 ,
         \26337_26639 , \26338_26640 , \26339_26641 , \26340_26642 , \26341_26643 , \26342_26644 , \26343_26645 , \26344_26646 , \26345_26647 , \26346_26648 ,
         \26347_26649 , \26348_26650 , \26349_26651 , \26350_26652 , \26351_26653 , \26352_26654 , \26353_26655 , \26354_26656 , \26355_26657 , \26356_26658 ,
         \26357_26659 , \26358_26660 , \26359_26661 , \26360_26662 , \26361_26663 , \26362_26664 , \26363_26665 , \26364_26666 , \26365_26667 , \26366_26668 ,
         \26367_26669 , \26368_26670 , \26369_26671 , \26370 , \26371_26673 , \26372_26674 , \26373_26675 , \26374_26676 , \26375_26677 , \26376_26678 ,
         \26377_26679 , \26378_26680 , \26379_26681 , \26380_26682 , \26381_26683 , \26382_26684 , \26383_26685 , \26384_26686 , \26385_26687 , \26386_26688 ,
         \26387_26689 , \26388_26690 , \26389_26691 , \26390_26692 , \26391_26693 , \26392_26694 , \26393_26695 , \26394_26696 , \26395_26697 , \26396_26698 ,
         \26397_26699 , \26398_26700 , \26399_26701 , \26400_26702 , \26401_26703 , \26402_26704 , \26403_26705 , \26404_26706 , \26405_26707 , \26406_26708 ,
         \26407_26709 , \26408_26710 , \26409_26711 , \26410_26712 , \26411_26713 , \26412_26714 , \26413_26715 , \26414_26716 , \26415_26717 , \26416_26718 ,
         \26417_26719 , \26418_26720 , \26419_26721 , \26420_26722 , \26421_26723 , \26422_26724 , \26423_26725 , \26424_26726 , \26425_26727 , \26426_26728 ,
         \26427_26729 , \26428_26730 , \26429_26731 , \26430_26732 , \26431_26733 , \26432_26734 , \26433_26735 , \26434_26736 , \26435_26737 , \26436_26738 ,
         \26437_26739 , \26438_26740 , \26439_26741 , \26440_26742 , \26441_26743 , \26442_26744 , \26443_26745 , \26444_26746 , \26445_26747 , \26446_26748 ,
         \26447_26749 , \26448_26750 , \26449_26751 , \26450_26752 , \26451_26753 , \26452_26754 , \26453_26755 , \26454_26756 , \26455_26757 , \26456_26758 ,
         \26457_26759 , \26458_26760 , \26459_26761 , \26460_26762 , \26461_26763 , \26462_26764 , \26463_26765 , \26464_26766 , \26465_26767 , \26466_26768 ,
         \26467_26769 , \26468_26770 , \26469_26771 , \26470_26772 , \26471_26773 , \26472_26774 , \26473_26775 , \26474_26776 , \26475_26777 , \26476_26778 ,
         \26477_26779 , \26478_26780 , \26479_26781 , \26480_26782 , \26481_26783 , \26482_26784 , \26483_26785 , \26484_26786 , \26485_26787 , \26486_26788 ,
         \26487_26789 , \26488_26790 , \26489_26791 , \26490_26792 , \26491_26793 , \26492_26794 , \26493_26795 , \26494_26796 , \26495_26797 , \26496_26798 ,
         \26497_26799 , \26498_26800 , \26499_26801 , \26500_26802 , \26501_26803 , \26502 , \26503_26805_nG5e37 , \26504_26806 , \26505_26807 , \26506_26808 ,
         \26507_26809 , \26508_26810 , \26509_26811 , \26510_26812 , \26511_26813 , \26512_26814 , \26513_26815 , \26514_26816 , \26515_26817 , \26516_26818 ,
         \26517_26819 , \26518_26820 , \26519_26821 , \26520_26822 , \26521_26823 , \26522_26824 , \26523_26825 , \26524 , \26525 , \26526_26828_nG65c1 ,
         \26527_26829 , \26528_26830 , \26529_26831 , \26530_26832 , \26531_26833 , \26532_26834 , \26533_26835 , \26534_26836 , \26535_26837 , \26536_26838 ,
         \26537_26839 , \26538_26840 , \26539_26841 , \26540_26842 , \26541_26843 , \26542_26844 , \26543_26845 , \26544_26846 , \26545_26847 , \26546_26848 ,
         \26547_26849 , \26548_26850 , \26549_26851 , \26550_26852 , \26551_26853 , \26552_26854 , \26553_26855 , \26554_26856 , \26555_26857 , \26556_26858 ,
         \26557_26859 , \26558_26860 , \26559_26861 , \26560_26862 , \26561_26863 , \26562_26864 , \26563_26865 , \26564_26866 , \26565_26867 , \26566_26868 ,
         \26567_26869 , \26568_26870 , \26569_26871 , \26570_26872 , \26571_26873 , \26572_26874 , \26573_26875 , \26574_26876 , \26575_26877 , \26576_26878 ,
         \26577_26879 , \26578_26880 , \26579_26881 , \26580_26882 , \26581_26883 , \26582_26884 , \26583_26885 , \26584_26886 , \26585_26887_nG9bc6 , \26586_26888 ,
         \26587_26889 , \26588_26890 , \26589_26891 , \26590_26892 , \26591_26893 , \26592_26894 , \26593_26895 , \26594_26896 , \26595_26897 , \26596_26898 ,
         \26597_26899 , \26598_26900 , \26599_26901 , \26600_26902 , \26601_26903 , \26602_26904 , \26603_26905 , \26604_26906 , \26605_26907 , \26606_26908 ,
         \26607_26909 , \26608_26910 , \26609_26911 , \26610_26912 , \26611_26913 , \26612_26914 , \26613_26915 , \26614_26916 , \26615_26917 , \26616_26918 ,
         \26617_26919 , \26618_26920 , \26619_26921 , \26620_26922 , \26621_26923 , \26622_26924 , \26623_26925 , \26624_26926 , \26625_26927 , \26626_26928 ,
         \26627_26929 , \26628_26930 , \26629_26931 , \26630_26932 , \26631_26933 , \26632_26934 , \26633_26935 , \26634_26936 , \26635_26937 , \26636_26938 ,
         \26637_26939 , \26638_26940 , \26639_26941 , \26640_26942 , \26641_26943 , \26642_26944 , \26643_26945 , \26644_26946 , \26645_26947 , \26646_26948 ,
         \26647_26949 , \26648_26950 , \26649_26951 , \26650_26952 , \26651_26953 , \26652_26954 , \26653_26955 , \26654_26956 , \26655_26957 , \26656_26958 ,
         \26657_26959 , \26658_26960 , \26659_26961 , \26660_26962 , \26661_26963 , \26662_26964 , \26663_26965 , \26664_26966 , \26665_26967 , \26666_26968 ,
         \26667_26969 , \26668_26970 , \26669_26971 , \26670_26972 , \26671_26973 , \26672_26974 , \26673_26975 , \26674_26976 , \26675_26977 , \26676_26978 ,
         \26677_26979 , \26678_26980 , \26679_26981 , \26680_26982 , \26681_26983 , \26682_26984 , \26683_26985 , \26684_26986 , \26685_26987 , \26686_26988 ,
         \26687_26989 , \26688_26990 , \26689_26991 , \26690_26992 , \26691_26993 , \26692_26994 , \26693_26995 , \26694_26996 , \26695_26997 , \26696_26998 ,
         \26697_26999 , \26698_27000 , \26699_27001 , \26700_27002 , \26701_27003 , \26702_27004 , \26703_27005 , \26704_27006 , \26705_27007 , \26706_27008 ,
         \26707_27009 , \26708_27010 , \26709_27011 , \26710_27012 , \26711_27013 , \26712_27014 , \26713_27015 , \26714_27016 , \26715_27017 , \26716_27018 ,
         \26717_27019 , \26718_27020 , \26719_27021 , \26720_27022 , \26721_27023 , \26722_27024 , \26723_27025 , \26724_27026 , \26725_27027 , \26726_27028 ,
         \26727_27029 , \26728_27030 , \26729_27031 , \26730_27032 , \26731_27033 , \26732_27034 , \26733_27035 , \26734_27036 , \26735_27037 , \26736_27038 ,
         \26737_27039 , \26738_27040 , \26739_27041 , \26740_27042 , \26741_27043 , \26742_27044 , \26743_27045 , \26744_27046 , \26745_27047 , \26746_27048 ,
         \26747_27049 , \26748_27050 , \26749_27051 , \26750_27052 , \26751_27053 , \26752_27054 , \26753_27055 , \26754_27056 , \26755_27057 , \26756_27058 ,
         \26757_27059 , \26758_27060 , \26759_27061 , \26760_27062 , \26761_27063 , \26762_27064 , \26763_27065 , \26764_27066 , \26765_27067 , \26766_27068 ,
         \26767_27069 , \26768_27070 , \26769_27071 , \26770_27072 , \26771_27073 , \26772_27074 , \26773_27075 , \26774_27076 , \26775_27077 , \26776_27078 ,
         \26777_27079 , \26778_27080 , \26779_27081 , \26780_27082 , \26781_27083 , \26782_27084 , \26783_27085 , \26784_27086 , \26785_27087 , \26786_27088 ,
         \26787_27089 , \26788_27090 , \26789_27091 , \26790_27092 , \26791_27093 , \26792_27094 , \26793_27095 , \26794_27096 , \26795_27097 , \26796_27098 ,
         \26797_27099 , \26798_27100 , \26799_27101 , \26800_27102 , \26801_27103 , \26802_27104 , \26803_27105 , \26804_27106 , \26805_27107 , \26806_27108 ,
         \26807_27109 , \26808_27110 , \26809_27111 , \26810_27112 , \26811_27113 , \26812_27114 , \26813_27115 , \26814_27116 , \26815_27117 , \26816_27118 ,
         \26817_27119 , \26818_27120 , \26819_27121 , \26820_27122 , \26821_27123 , \26822_27124 , \26823_27125 , \26824_27126 , \26825_27127 , \26826_27128 ,
         \26827_27129 , \26828_27130 , \26829_27131 , \26830_27132 , \26831_27133 , \26832_27134 , \26833_27135 , \26834_27136 , \26835_27137 , \26836_27138 ,
         \26837_27139 , \26838_27140 , \26839_27141 , \26840_27142 , \26841_27143 , \26842_27144 , \26843_27145 , \26844_27146 , \26845_27147 , \26846_27148 ,
         \26847_27149 , \26848_27150 , \26849_27151 , \26850_27152 , \26851_27153 , \26852_27154 , \26853_27155 , \26854_27156 , \26855_27157 , \26856 ,
         \26857_27159 , \26858_27160 , \26859_27161 , \26860_27162 , \26861_27163 , \26862_27164 , \26863_27165 , \26864_27166 , \26865_27167 , \26866_27168 ,
         \26867_27169 , \26868_27170 , \26869_27171 , \26870_27172 , \26871_27173 , \26872_27174 , \26873_27175 , \26874_27176 , \26875_27177 , \26876_27178 ,
         \26877_27179 , \26878_27180 , \26879_27181 , \26880_27182 , \26881_27183 , \26882_27184 , \26883_27185 , \26884_27186 , \26885_27187 , \26886_27188 ,
         \26887_27189 , \26888_27190 , \26889_27191 , \26890_27192 , \26891_27193 , \26892_27194 , \26893_27195 , \26894_27196 , \26895_27197 , \26896_27198 ,
         \26897_27199 , \26898_27200 , \26899_27201 , \26900_27202 , \26901_27203 , \26902_27204 , \26903_27205 , \26904_27206 , \26905_27207 , \26906_27208 ,
         \26907_27209 , \26908_27210 , \26909_27211 , \26910_27212 , \26911_27213 , \26912_27214 , \26913_27215 , \26914_27216 , \26915_27217 , \26916_27218 ,
         \26917_27219 , \26918_27220 , \26919_27221 , \26920_27222 , \26921_27223 , \26922_27224 , \26923_27225 , \26924_27226 , \26925_27227 , \26926_27228 ,
         \26927_27229 , \26928_27230 , \26929_27231 , \26930_27232 , \26931_27233 , \26932_27234 , \26933_27235 , \26934_27236 , \26935_27237 , \26936_27238 ,
         \26937_27239 , \26938_27240 , \26939_27241 , \26940_27242 , \26941_27243 , \26942_27244 , \26943_27245 , \26944_27246 , \26945_27247 , \26946_27248 ,
         \26947_27249 , \26948_27250 , \26949_27251 , \26950_27252 , \26951_27253 , \26952_27254 , \26953_27255 , \26954_27256 , \26955_27257 , \26956_27258 ,
         \26957_27259 , \26958_27260 , \26959_27261 , \26960_27262 , \26961_27263 , \26962_27264 , \26963_27265 , \26964_27266 , \26965_27267 , \26966_27268 ,
         \26967_27269 , \26968_27270 , \26969_27271 , \26970_27272 , \26971_27273 , \26972_27274 , \26973_27275 , \26974_27276 , \26975_27277 , \26976_27278 ,
         \26977_27279 , \26978_27280 , \26979_27281 , \26980_27282 , \26981_27283 , \26982_27284 , \26983_27285 , \26984_27286 , \26985_27287 , \26986_27288 ,
         \26987_27289 , \26988 , \26989_27291_nG5f40 , \26990_27292 , \26991_27293 , \26992_27294 , \26993_27295 , \26994_27296 , \26995_27297 , \26996_27298 ,
         \26997_27299 , \26998_27300 , \26999_27301 , \27000_27302 , \27001_27303 , \27002_27304 , \27003_27305 , \27004_27306 , \27005_27307 , \27006_27308 ,
         \27007_27309 , \27008 , \27009 , \27010_27312_nG65c4 , \27011_27313 , \27012_27314 , \27013_27315 , \27014_27316 , \27015_27317 , \27016_27318 ,
         \27017_27319 , \27018_27320 , \27019_27321 , \27020_27322 , \27021_27323 , \27022_27324 , \27023_27325 , \27024_27326 , \27025_27327 , \27026_27328 ,
         \27027_27329 , \27028_27330 , \27029_27331 , \27030_27332 , \27031_27333 , \27032_27334 , \27033_27335 , \27034_27336 , \27035_27337 , \27036_27338 ,
         \27037_27339 , \27038_27340 , \27039_27341 , \27040_27342 , \27041_27343 , \27042_27344 , \27043_27345 , \27044_27346 , \27045_27347 , \27046_27348 ,
         \27047_27349 , \27048_27350 , \27049_27351 , \27050_27352 , \27051_27353 , \27052_27354 , \27053_27355 , \27054_27356 , \27055_27357 , \27056_27358 ,
         \27057_27359 , \27058_27360 , \27059_27361 , \27060_27362 , \27061_27363 , \27062_27364 , \27063_27365 , \27064_27366 , \27065_27367 , \27066_27368 ,
         \27067_27369 , \27068_27370 , \27069_27371 , \27070_27372 , \27071_27373 , \27072_27374 , \27073_27375 , \27074_27376 , \27075_27377 , \27076_27378 ,
         \27077_27379 , \27078_27380 , \27079_27381 , \27080_27382 , \27081_27383 , \27082_27384 , \27083_27385 , \27084_27386 , \27085_27387 , \27086_27388 ,
         \27087_27389 , \27088_27390 , \27089_27391 , \27090_27392 , \27091_27393 , \27092_27394 , \27093_27395 , \27094_27396 , \27095_27397 , \27096_27398 ,
         \27097_27399 , \27098_27400 , \27099_27401 , \27100_27402 , \27101_27403 , \27102_27404 , \27103_27405 , \27104_27406 , \27105_27407 , \27106_27408 ,
         \27107_27409 , \27108_27410 , \27109_27411 , \27110_27412 , \27111_27413 , \27112_27414 , \27113_27415 , \27114_27416_nG9bc3 , \27115_27417 , \27116_27418 ,
         \27117_27419 , \27118_27420 , \27119_27421 , \27120_27422 , \27121_27423 , \27122_27424 , \27123_27425 , \27124_27426 , \27125_27427 , \27126_27428 ,
         \27127_27429 , \27128_27430 , \27129_27431 , \27130_27432 , \27131_27433 , \27132_27434 , \27133_27435 , \27134_27436 , \27135_27437 , \27136_27438 ,
         \27137_27439 , \27138_27440 , \27139_26429 , \27140_26430 , \27141_26431 , \27142_27441 , \27143_27442 , \27144_27443 , \27145_27444 , \27146_27445 ,
         \27147_27446 , \27148_27447 , \27149_27448 , \27150_27449 , \27151_27450 , \27152_27451 , \27153_27452 , \27154_27453 , \27155_27454 , \27156_27455 ,
         \27157_27456 , \27158_27457 , \27159_27458 , \27160_27459 , \27161_27460 , \27162_27461 , \27163_27462 , \27164_27463 , \27165_27464 , \27166_27465 ,
         \27167_27466 , \27168_27467 , \27169_27468 , \27170_27469 , \27171_27470 , \27172_27471 , \27173_27472 , \27174_27473 , \27175_27474 , \27176_27475 ,
         \27177_27476 , \27178_27477 , \27179_27478 , \27180_27479 , \27181_27480 , \27182_27481 , \27183_27482 , \27184_27483 , \27185_27484 , \27186_27485 ,
         \27187_27486 , \27188_27487 , \27189_27488 , \27190_27489 , \27191_27490 , \27192_27491 , \27193_27492 , \27194_27493 , \27195_27494 , \27196_27495 ,
         \27197_27496 , \27198_27497 , \27199_27498 , \27200_27499 , \27201_27500 , \27202_27501 , \27203_27502 , \27204_27503 , \27205_27504 , \27206_27505 ,
         \27207_27506 , \27208_27507 , \27209_27508 , \27210_27509 , \27211_27510 , \27212_27511 , \27213_27512 , \27214_27513 , \27215_27514 , \27216_27515 ,
         \27217_27516 , \27218_27517 , \27219_27518 , \27220_27519 , \27221_27520 , \27222_27521 , \27223_27522 , \27224_27523 , \27225_27524 , \27226_27525 ,
         \27227_27526 , \27228_27527 , \27229_27528 , \27230_27529 , \27231_27530 , \27232_27531 , \27233_27532 , \27234_27533 , \27235_27534 , \27236_27535 ,
         \27237_27536 , \27238_27537 , \27239_27538 , \27240_27539 , \27241_27540 , \27242_27541 , \27243_27542 , \27244_27543 , \27245_27544 , \27246_27545 ,
         \27247_27546 , \27248_27547 , \27249_27548 , \27250_27549 , \27251_27550 , \27252_27551 , \27253_27552 , \27254_27553 , \27255_27554 , \27256_27555 ,
         \27257_27556 , \27258_27557 , \27259_27558 , \27260_27559 , \27261_27560 , \27262_27561 , \27263_27562 , \27264_27563 , \27265_27564 , \27266_27565 ,
         \27267_27566 , \27268_27567 , \27269_27568 , \27270_27569 , \27271_27570 , \27272_27571 , \27273_27572 , \27274_27573 , \27275_27574 , \27276_27575 ,
         \27277_27576 , \27278_27577 , \27279_27578 , \27280_27579 , \27281_27580 , \27282_27581 , \27283_27582 , \27284_27583 , \27285_27584 , \27286_27585 ,
         \27287_27586 , \27288_27587 , \27289_27588 , \27290_27589 , \27291_27590 , \27292_27591 , \27293_27592 , \27294_27593 , \27295_27594 , \27296_27595 ,
         \27297_27596 , \27298_27597 , \27299_27598 , \27300_27599 , \27301_27600 , \27302_27601 , \27303_27602 , \27304_27603 , \27305_27604 , \27306_27605 ,
         \27307_27606 , \27308_27607 , \27309_27608 , \27310_27609 , \27311_27610 , \27312_27611 , \27313_27612 , \27314_27613 , \27315_27614 , \27316_27615 ,
         \27317_27616 , \27318_27617 , \27319_27618 , \27320_27619 , \27321_27620 , \27322_27621 , \27323_27622 , \27324_27623 , \27325_27624 , \27326_27625 ,
         \27327_27626 , \27328_27627 , \27329_27628 , \27330_27629 , \27331_27630 , \27332_27631 , \27333_27632 , \27334_27633 , \27335_27634 , \27336_27635 ,
         \27337_27636 , \27338_27637 , \27339_27638 , \27340_27639 , \27341_27640 , \27342_27641 , \27343_27642 , \27344_27643 , \27345_27644 , \27346_27645 ,
         \27347_27646 , \27348_27647 , \27349_27648 , \27350_27649 , \27351_27650 , \27352_27651 , \27353_27652 , \27354_27653 , \27355_27654 , \27356_27655 ,
         \27357_27656 , \27358_27657 , \27359_27658 , \27360_27659 , \27361_27660 , \27362_27661 , \27363_27662 , \27364_27663 , \27365_27664 , \27366_27665 ,
         \27367_27666 , \27368_27667 , \27369_27668 , \27370_27669 , \27371_27670 , \27372_27671 , \27373_27672 , \27374_27673 , \27375_27674 , \27376_27675 ,
         \27377_27676 , \27378_27677 , \27379_27678 , \27380_27679 , \27381_27680 , \27382_27681 , \27383_27682 , \27384_27683 , \27385_27684 , \27386_27685 ,
         \27387_27686 , \27388_27687 , \27389_27688 , \27390_27689 , \27391_27690 , \27392_27691 , \27393_27692 , \27394_27693 , \27395_27694 , \27396_27695 ,
         \27397_27696 , \27398_27697 , \27399 , \27400_27699 , \27401_27700 , \27402_27701 , \27403_27702 , \27404_27703 , \27405_27704 , \27406_27705 ,
         \27407_27706 , \27408_27707 , \27409_27708 , \27410_27709 , \27411_27710 , \27412_27711 , \27413_27712 , \27414_27713 , \27415_27714 , \27416_27715 ,
         \27417_27716 , \27418_27717 , \27419_27718 , \27420_27719 , \27421_27720 , \27422_27721 , \27423_27722 , \27424_27723 , \27425_27724 , \27426_27725 ,
         \27427_27726 , \27428_27727 , \27429_27728 , \27430_27729 , \27431_27730 , \27432_27731 , \27433_27732 , \27434_27733 , \27435_27734 , \27436_27735 ,
         \27437_27736 , \27438_27737 , \27439_27738 , \27440_27739 , \27441_27740 , \27442_27741 , \27443_27742 , \27444_27743 , \27445_27744 , \27446_27745 ,
         \27447_27746 , \27448_27747 , \27449_27748 , \27450_27749 , \27451_27750 , \27452_27751 , \27453_27752 , \27454_27753 , \27455_27754 , \27456_27755 ,
         \27457_27756 , \27458_27757 , \27459_27758 , \27460_27759 , \27461_27760 , \27462_27761 , \27463_27762 , \27464_27763 , \27465_27764 , \27466_27765 ,
         \27467_27766 , \27468_27767 , \27469_27768 , \27470_27769 , \27471_27770 , \27472_27771 , \27473_27772 , \27474_27773 , \27475_27774 , \27476_27775 ,
         \27477_27776 , \27478_27777 , \27479_27778 , \27480_27779 , \27481_27780 , \27482_27781 , \27483_27782 , \27484_27783 , \27485_27784 , \27486_27785 ,
         \27487_27786 , \27488_27787 , \27489_27788 , \27490_27789 , \27491_27790 , \27492_27791 , \27493_27792 , \27494_27793 , \27495_27794 , \27496_27795 ,
         \27497_27796 , \27498_27797 , \27499_27798 , \27500_27799 , \27501_27800 , \27502_27801 , \27503_27802 , \27504_27803 , \27505_27804 , \27506_27805 ,
         \27507_27806 , \27508_27807 , \27509_27808 , \27510_27809 , \27511_27810 , \27512_27811 , \27513_27812 , \27514_27813 , \27515_27814 , \27516_27815 ,
         \27517_27816 , \27518_27817 , \27519_27818 , \27520_27819 , \27521_27820 , \27522_27821 , \27523_27822 , \27524_27823 , \27525_27824 , \27526_27825 ,
         \27527_27826 , \27528_27827 , \27529_27828 , \27530_27829 , \27531_27830 , \27532 , \27533_27832 , \27534_27833 , \27535_27834 , \27536_27835 ,
         \27537_27836 , \27538_27837 , \27539_27838 , \27540_27839 , \27541_27840 , \27542_27841 , \27543_27842 , \27544_27843 , \27545_27844 , \27546_27845 ,
         \27547_27846 , \27548_27847 , \27549_27848 , \27550_27849 , \27551_27850 , \27552_27851 , \27553_27852 , \27554_27853 , \27555_27854 , \27556_27855 ,
         \27557_27856 , \27558_27857 , \27559_27858 , \27560_27859 , \27561_27860 , \27562_27861 , \27563_27862 , \27564_27863 , \27565_27864 , \27566_27865 ,
         \27567_27866 , \27568_27867 , \27569_27868 , \27570_27869 , \27571_27870 , \27572_27871 , \27573_27872 , \27574_27873 , \27575_27874 , \27576_27875 ,
         \27577_27876 , \27578_27877 , \27579_27878 , \27580_27879 , \27581_27880 , \27582_27881 , \27583_27882 , \27584_27883 , \27585_27884 , \27586_27885 ,
         \27587_27886 , \27588_27887 , \27589_27888 , \27590_27889 , \27591_27890 , \27592_27891 , \27593_27892 , \27594_27893 , \27595_27894 , \27596_27895 ,
         \27597_27896 , \27598_27897 , \27599_27898 , \27600_27899 , \27601_27900 , \27602_27901 , \27603_27902 , \27604_27903 , \27605_27904 , \27606_27905 ,
         \27607_27906 , \27608_27907 , \27609_27908 , \27610_27909 , \27611_27910 , \27612_27911 , \27613_27912 , \27614_27913 , \27615_27914 , \27616_27915 ,
         \27617_27916 , \27618_27917 , \27619_27918 , \27620_27919 , \27621_27920 , \27622_27921 , \27623_27922 , \27624_27923 , \27625_27924 , \27626_27925 ,
         \27627_27926 , \27628_27927 , \27629_27928 , \27630_27929 , \27631_27930 , \27632_27931 , \27633_27932 , \27634_27933 , \27635_27934 , \27636_27935 ,
         \27637_27936 , \27638_27937 , \27639_27938 , \27640_27939 , \27641_27940 , \27642_27941 , \27643_27942 , \27644_27943 , \27645_27944 , \27646_27945 ,
         \27647_27946 , \27648_27947 , \27649_27948 , \27650_27949 , \27651_27950 , \27652_27951 , \27653_27952 , \27654_27953 , \27655_27954 , \27656_27955 ,
         \27657_27956 , \27658_27957 , \27659_27958 , \27660_27959 , \27661_27960 , \27662_27961 , \27663_27962 , \27664_27963 , \27665_27964 , \27666 ,
         \27667_27966 , \27668_27967 , \27669_27968 , \27670_27969 , \27671_27970 , \27672_27971 , \27673_27972 , \27674_27973 , \27675_27974 , \27676_27975 ,
         \27677_27976 , \27678_27977 , \27679_27978 , \27680_27979 , \27681_27980 , \27682_27981 , \27683_27982 , \27684_27983 , \27685_27984 , \27686_27985 ,
         \27687_27986 , \27688_27987 , \27689_27988 , \27690_27989 , \27691_27990 , \27692_27991 , \27693_27992 , \27694_27993 , \27695_27994 , \27696_27995 ,
         \27697_27996 , \27698_27997 , \27699_27998 , \27700_27999 , \27701_28000 , \27702_28001 , \27703_28002 , \27704_28003 , \27705_28004 , \27706_28005 ,
         \27707_28006 , \27708_28007 , \27709_28008 , \27710_28009 , \27711_28010 , \27712_28011 , \27713_28012 , \27714_28013 , \27715_28014 , \27716_28015 ,
         \27717_28016 , \27718_28017 , \27719_28018 , \27720_28019 , \27721_28020 , \27722_28021 , \27723_28022 , \27724_28023 , \27725_28024 , \27726_28025 ,
         \27727_28026 , \27728_28027 , \27729_28028 , \27730_28029 , \27731_28030 , \27732_28031 , \27733_28032 , \27734_28033 , \27735_28034 , \27736_28035 ,
         \27737_28036 , \27738_28037 , \27739_28038 , \27740_28039 , \27741_28040 , \27742_28041 , \27743_28042 , \27744_28043 , \27745_28044 , \27746_28045 ,
         \27747_28046 , \27748_28047 , \27749_28048 , \27750_28049 , \27751_28050 , \27752_28051 , \27753_28052 , \27754_28053 , \27755_28054 , \27756_28055 ,
         \27757_28056 , \27758_28057 , \27759_28058 , \27760_28059 , \27761_28060 , \27762_28061 , \27763_28062 , \27764_28063 , \27765_28064 , \27766_28065 ,
         \27767_28066 , \27768_28067 , \27769_28068 , \27770_28069 , \27771_28070 , \27772_28071 , \27773_28072 , \27774_28073 , \27775_28074 , \27776_28075 ,
         \27777_28076 , \27778_28077 , \27779_28078 , \27780_28079 , \27781_28080 , \27782_28081 , \27783_28082 , \27784_28083 , \27785_28084 , \27786_28085 ,
         \27787_28086 , \27788_28087 , \27789_28088 , \27790_28089 , \27791_28090 , \27792_28091 , \27793_28092 , \27794_28093 , \27795_28094 , \27796_28095 ,
         \27797_28096 , \27798_28097 , \27799 , \27800_28099 , \27801_28100 , \27802_28101 , \27803_28102 , \27804_28103 , \27805_28104 , \27806_28105 ,
         \27807_28106 , \27808_28107 , \27809_28108 , \27810_28109_nG4406 , \27811_28110 , \27812_28111 , \27813_28112_nG4409 , \27814_28113 , \27815_28114 , \27816_28115 ,
         \27817_28119 , \27818_28120 , \27819_28121 , \27820_28122 , \27821_28123 , \27822_28124 , \27823_28125 , \27824_28126 , \27825_28127 , \27826_28128 ,
         \27827_28129 , \27828_28130 , \27829_28131 , \27830_28132 , \27831_28133 , \27832_28134 , \27833_28135 , \27834_28136 , \27835_28137 , \27836_28138 ,
         \27837_28139 , \27838_28140 , \27839_28141 , \27840_28142 , \27841_28143 , \27842_28144 , \27843_28145 , \27844_28146 , \27845_28147 , \27846_28148 ,
         \27847_28149 , \27848_28150 , \27849_28151 , \27850_28152 , \27851_28153 , \27852_28154 , \27853_28155 , \27854_28156 , \27855_28157 , \27856_28158 ,
         \27857_28159 , \27858_28160 , \27859_28161 , \27860_28162 , \27861_28163 , \27862_28164 , \27863_28165 , \27864_28166 , \27865_28167 , \27866_28168 ,
         \27867_28169 , \27868_28170 , \27869_28171 , \27870_28172 , \27871_28173 , \27872_28174 , \27873_28175 , \27874_28176 , \27875_28177 , \27876_28178 ,
         \27877_28179 , \27878_28180 , \27879_28181 , \27880_28182 , \27881_28183 , \27882_28184 , \27883_28185 , \27884_28186 , \27885_28187 , \27886_28188 ,
         \27887_28189 , \27888_28190 , \27889_28191 , \27890_28192 , \27891_28193 , \27892_28194 , \27893_28195 , \27894_28196 , \27895_28197 , \27896_28198 ,
         \27897_28199 , \27898_28200 , \27899_28201 , \27900_28202 , \27901_28203 , \27902_28204 , \27903_28205 , \27904_28206 , \27905_28207 , \27906_28208 ,
         \27907_28209 , \27908_28210 , \27909_28211 , \27910_28212 , \27911_28213 , \27912_28214 , \27913_28215 , \27914_28216 , \27915_28217 , \27916_28218 ,
         \27917_28219 , \27918_28220 , \27919_28221 , \27920_28222 , \27921_28223 , \27922_28224 , \27923_28225 , \27924_28226 , \27925_28227 , \27926_28228 ,
         \27927_28229 , \27928_28230 , \27929_28231 , \27930_28232 , \27931_28233 , \27932_28234 , \27933_28235 , \27934_28236 , \27935_28237 , \27936_28238 ,
         \27937_28239 , \27938_28240 , \27939_28241 , \27940_28242 , \27941_28243 , \27942_28244 , \27943_28245 , \27944_28246 , \27945_28247 , \27946_28248 ,
         \27947_28249 , \27948_28250 , \27949_28251 , \27950_28252 , \27951_28253 , \27952_28254 , \27953_28255 , \27954_28256 , \27955_28257 , \27956_28258 ,
         \27957_28259 , \27958_28260 , \27959_28261 , \27960_28262 , \27961_28263 , \27962_28264 , \27963_28265 , \27964_28266 , \27965_28267 , \27966_28268 ,
         \27967_28269 , \27968_28270 , \27969_28271 , \27970_28272 , \27971_28273 , \27972_28274 , \27973_28275 , \27974_28276 , \27975_28277 , \27976_28278 ,
         \27977_28279 , \27978_28280 , \27979_28281 , \27980_28282 , \27981_28283 , \27982_28284 , \27983_28285 , \27984_28286 , \27985_28287 , \27986_28288 ,
         \27987_28289 , \27988_28290 , \27989_28291 , \27990_28292 , \27991_28293 , \27992_28294 , \27993_28295 , \27994_28296 , \27995_28297 , \27996_28298 ,
         \27997_28299 , \27998_28300 , \27999_28301 , \28000_28302 , \28001_28303 , \28002_28304 , \28003_28305 , \28004_28306 , \28005_28307 , \28006_28308 ,
         \28007_28309 , \28008_28310 , \28009_28311 , \28010_28312 , \28011_28313 , \28012_28314 , \28013_28315 , \28014_28316 , \28015_28317 , \28016_28318 ,
         \28017_28319 , \28018_28320 , \28019_28321 , \28020_28322 , \28021_28323 , \28022_28324 , \28023_28325 , \28024_28326 , \28025_28327 , \28026_28328 ,
         \28027_28329 , \28028_28330 , \28029_28331 , \28030_28332 , \28031_28333 , \28032_28334 , \28033_28335 , \28034_28336 , \28035_28337 , \28036_28338 ,
         \28037_28339 , \28038_28340 , \28039_28341 , \28040_28342 , \28041_28343 , \28042_28344 , \28043_28345 , \28044_28346 , \28045_28347 , \28046_28348 ,
         \28047_28349 , \28048_28350 , \28049_28351 , \28050_28352 , \28051_28353 , \28052_28354 , \28053_28355 , \28054_28356 , \28055_28357 , \28056_28358 ,
         \28057_28359 , \28058_28360 , \28059_28361 , \28060_28362 , \28061_28363 , \28062_28364 , \28063_28365 , \28064_28366 , \28065_28367 , \28066_28368 ,
         \28067_28369 , \28068_28370 , \28069_28371 , \28070_28372 , \28071_28373 , \28072_28374 , \28073_28375 , \28074_28376 , \28075_28377 , \28076_28378 ,
         \28077_28379 , \28078_28380 , \28079_28381 , \28080_28382 , \28081_28383 , \28082_28384 , \28083_28385 , \28084_28386 , \28085_28387 , \28086_28388 ,
         \28087_28389 , \28088_28390 , \28089 , \28090_28392 , \28091_28393 , \28092_28394 , \28093_28395 , \28094_28396 , \28095_28397 , \28096_28398 ,
         \28097_28399 , \28098_28400 , \28099_28401 , \28100_28402 , \28101_28403 , \28102_28404 , \28103_28405 , \28104_28406 , \28105_28407 , \28106_28408 ,
         \28107_28409 , \28108_28410 , \28109_28411 , \28110_28412 , \28111_28413 , \28112_28414 , \28113_28415 , \28114_28416 , \28115_28417 , \28116_28418 ,
         \28117_28419 , \28118_28420 , \28119_28421 , \28120_28422 , \28121_28423 , \28122_28424 , \28123_28425 , \28124_28426 , \28125_28427 , \28126_28428 ,
         \28127_28429 , \28128_28430 , \28129_28431 , \28130_28432 , \28131_28433 , \28132_28434 , \28133_28435 , \28134_28436 , \28135_28437 , \28136_28438 ,
         \28137_28439 , \28138_28440 , \28139_28441 , \28140_28442 , \28141_28443 , \28142_28444 , \28143_28445 , \28144_28446 , \28145_28447 , \28146_28448 ,
         \28147_28449 , \28148_28450 , \28149_28451 , \28150_28452 , \28151_28453 , \28152_28454 , \28153_28455 , \28154_28456 , \28155_28457 , \28156_28458 ,
         \28157_28459 , \28158_28460 , \28159_28461 , \28160_28462 , \28161_28463 , \28162_28464 , \28163_28465 , \28164_28466 , \28165_28467 , \28166_28468 ,
         \28167_28469 , \28168_28470 , \28169_28471 , \28170_28472 , \28171_28473 , \28172_28474 , \28173_28475 , \28174_28476 , \28175_28477 , \28176_28478 ,
         \28177_28479 , \28178_28480 , \28179_28481 , \28180_28482 , \28181_28483 , \28182_28484 , \28183_28485 , \28184_28486 , \28185_28487 , \28186_28488 ,
         \28187_28489 , \28188_28490 , \28189_28491 , \28190_28492 , \28191_28493 , \28192_28494 , \28193_28495 , \28194_28496 , \28195_28497 , \28196_28498 ,
         \28197_28499 , \28198_28500 , \28199_28501 , \28200_28502 , \28201_28503 , \28202_28504 , \28203_28505 , \28204_28506 , \28205_28507 , \28206_28508 ,
         \28207_28509 , \28208_28510 , \28209_28511 , \28210_28512 , \28211_28513 , \28212_28514 , \28213_28515 , \28214_28516 , \28215_28517 , \28216_28518 ,
         \28217_28519 , \28218_28520 , \28219_28521 , \28220_28522 , \28221 , \28222_28524_nG6049 , \28223_28525 , \28224_28526 , \28225_28527 , \28226_28528 ,
         \28227_28529 , \28228_28530 , \28229 , \28230 , \28231_28533_nG65c7 , \28232_28534 , \28233_28535 , \28234_28536 , \28235_28537 , \28236_28538 ,
         \28237_28539 , \28238_28540 , \28239_28541 , \28240_28542 , \28241_28543 , \28242_28544 , \28243_28545 , \28244_28546 , \28245_28547 , \28246_28548 ,
         \28247_28549 , \28248_28550 , \28249_28551 , \28250_28552 , \28251_28553 , \28252_28554 , \28253_28555 , \28254_28556 , \28255_28557 , \28256_28558 ,
         \28257_28559 , \28258_28560 , \28259_28561 , \28260_28562 , \28261_28563 , \28262_28564 , \28263_28565 , \28264_28566 , \28265_28567 , \28266_28568 ,
         \28267_28569 , \28268_28570 , \28269_28571 , \28270_28572 , \28271_28573 , \28272_28574 , \28273_28575 , \28274_28576 , \28275_28577 , \28276_28578 ,
         \28277_28579 , \28278_28580 , \28279_28581 , \28280_28582 , \28281_28583 , \28282_28584 , \28283_28585 , \28284_28586 , \28285_28587 , \28286_28588 ,
         \28287_28589 , \28288_28590 , \28289_28591 , \28290_28592 , \28291_28593 , \28292_28594 , \28293_28595 , \28294_28596 , \28295_28597 , \28296_28598 ,
         \28297_28599 , \28298_28600 , \28299_28601 , \28300_28602_nG9bc0 , \28301_28603 , \28302_28604 , \28303_28605 , \28304_28606 , \28305_28607 , \28306_28608 ,
         \28307_28609 , \28308_28610 , \28309_28611 , \28310_28612 , \28311_28613 , \28312_28614 , \28313_28615 , \28314_28616 , \28315_28617 , \28316_28618 ,
         \28317_28619 , \28318_28620 , \28319_28621 , \28320_28622 , \28321_28623 , \28322_28624 , \28323_28625 , \28324_28626 , \28325_28627 , \28326_28628 ,
         \28327_28629 , \28328_28630 , \28329_28631 , \28330_28632 , \28331_28633 , \28332_28634 , \28333_28635 , \28334_28636 , \28335_28637 , \28336_28638 ,
         \28337_28639 , \28338_28640 , \28339_28641 , \28340_28642 , \28341_28643 , \28342_28644 , \28343_28645 , \28344_28646 , \28345_28647 , \28346_28648 ,
         \28347_28649 , \28348_28650 , \28349_28651 , \28350_28652 , \28351_28653 , \28352_28654 , \28353_28655 , \28354_28656 , \28355_28657 , \28356_28658 ,
         \28357_28659 , \28358_28660 , \28359_28661 , \28360_28662 , \28361_28663 , \28362_28664 , \28363_28665 , \28364_28666 , \28365_28667 , \28366_28668 ,
         \28367_28669 , \28368_28670 , \28369_28671 , \28370_28672 , \28371_28673 , \28372_28674 , \28373_28675 , \28374_28676 , \28375_28677 , \28376_28678 ,
         \28377_28679 , \28378_28680 , \28379_28681 , \28380_28682 , \28381_28683 , \28382_28684 , \28383_28685 , \28384_28686 , \28385_28687 , \28386_28688 ,
         \28387_28689 , \28388_28690 , \28389_28691 , \28390_28692 , \28391_28693 , \28392_28694 , \28393_28695 , \28394_28696 , \28395_28697 , \28396_28698 ,
         \28397_28699 , \28398_28700 , \28399_28701 , \28400_28702 , \28401_28703 , \28402_28704 , \28403_28705 , \28404_28706 , \28405_28707 , \28406_28708 ,
         \28407_28709 , \28408_28710 , \28409_28711 , \28410_28712 , \28411_28713 , \28412_28714 , \28413_28715 , \28414_28716 , \28415_28717 , \28416_28718 ,
         \28417_28719 , \28418_28720 , \28419_28721 , \28420_28722 , \28421_28723 , \28422_28724 , \28423_28725 , \28424_28726 , \28425_28727 , \28426_28728 ,
         \28427_28729 , \28428_28730 , \28429_28731 , \28430_28732 , \28431_28733 , \28432_28734 , \28433_28735 , \28434_28736 , \28435_28737 , \28436_28738 ,
         \28437_28739 , \28438_28740 , \28439_28741 , \28440_28742 , \28441_28743 , \28442_28744 , \28443_28745 , \28444_28746 , \28445_28747 , \28446_28748 ,
         \28447_28749 , \28448_28750 , \28449_28751 , \28450_28752 , \28451_28753 , \28452_28754 , \28453_28755 , \28454_28756 , \28455_28757 , \28456_28758 ,
         \28457_28759 , \28458_28760 , \28459_28761 , \28460_28762 , \28461_28763 , \28462_28764 , \28463_28765 , \28464_28766 , \28465_28767 , \28466_28768 ,
         \28467_28769 , \28468_28770 , \28469_28771 , \28470_28772 , \28471_28773 , \28472_28774 , \28473_28775 , \28474_28776 , \28475_28777 , \28476_28778 ,
         \28477_28779 , \28478_28780 , \28479_28781 , \28480_28782 , \28481_28783 , \28482_28784 , \28483_28785 , \28484_28786 , \28485_28787 , \28486_28788 ,
         \28487_28789 , \28488_28790 , \28489_28791 , \28490_28792 , \28491_28793 , \28492_28794 , \28493_28795 , \28494_28796 , \28495_28797 , \28496_28798 ,
         \28497_28799 , \28498_28800 , \28499_28801 , \28500_28802 , \28501_28803 , \28502_28804 , \28503_28805 , \28504_28806 , \28505_28807 , \28506_28808 ,
         \28507_28809 , \28508_28810 , \28509_28811 , \28510_28812 , \28511_28813 , \28512_28814 , \28513_28815 , \28514_28816 , \28515_28817 , \28516_28818 ,
         \28517_28819 , \28518_28820 , \28519_28821 , \28520_28822 , \28521_28823 , \28522_28824 , \28523_28825 , \28524_28826 , \28525_28827 , \28526_28828 ,
         \28527_28829 , \28528_28830 , \28529_28831 , \28530_28832 , \28531_28833 , \28532_28834 , \28533_28835 , \28534_28836 , \28535_28837 , \28536_28838 ,
         \28537_28839 , \28538_28840 , \28539_28841 , \28540_28842 , \28541_28843 , \28542_28844 , \28543_28845 , \28544_28846 , \28545_28847 , \28546_28848 ,
         \28547_28849 , \28548_28850 , \28549_28851 , \28550_28852 , \28551_28853 , \28552_28854 , \28553_28855 , \28554_28856 , \28555_28857 , \28556_28858 ,
         \28557_28859 , \28558_28860 , \28559_28861 , \28560_28862 , \28561_28863 , \28562_28864 , \28563_28865 , \28564_28866 , \28565_28867 , \28566_28868 ,
         \28567_28869 , \28568_28870 , \28569_28871 , \28570_28872 , \28571_28873 , \28572_28874 , \28573_28875 , \28574_28876 , \28575_28877 , \28576_28878 ,
         \28577_28879 , \28578_28880 , \28579_28881 , \28580_28882 , \28581_28883 , \28582_28884 , \28583_28885 , \28584_28886 , \28585_28887 , \28586_28888 ,
         \28587_28889 , \28588_28890 , \28589_28891 , \28590_28892 , \28591_28893 , \28592_28894 , \28593_28895 , \28594_28896 , \28595_28897 , \28596_28898 ,
         \28597_28899 , \28598_28900 , \28599_28901 , \28600_28902 , \28601_28903 , \28602_28904 , \28603_28905 , \28604_28906 , \28605_28907 , \28606_28908 ,
         \28607_28909 , \28608_28910 , \28609_28911 , \28610_28912 , \28611_28913 , \28612_28914 , \28613_28915 , \28614_28916 , \28615_28917 , \28616_28918 ,
         \28617_28919 , \28618_28920 , \28619_28921 , \28620_28922 , \28621_28923 , \28622_28924 , \28623_28925 , \28624_28926 , \28625_28927 , \28626_28928 ,
         \28627_28929 , \28628_28930 , \28629_28931 , \28630_28932 , \28631 , \28632_28934 , \28633_28935 , \28634_28936 , \28635_28937 , \28636_28938 ,
         \28637_28939 , \28638_28940 , \28639_28941 , \28640_28942 , \28641_28943 , \28642_28944 , \28643_28945 , \28644_28946 , \28645_28947 , \28646_28948 ,
         \28647_28949 , \28648_28950 , \28649_28951 , \28650_28952 , \28651_28953 , \28652_28954 , \28653_28955 , \28654_28956 , \28655_28957 , \28656_28958 ,
         \28657_28959 , \28658_28960 , \28659_28961 , \28660_28962 , \28661_28963 , \28662_28964 , \28663_28965 , \28664_28966 , \28665_28967 , \28666_28968 ,
         \28667_28969 , \28668_28970 , \28669_28971 , \28670_28972 , \28671_28973 , \28672_28974 , \28673_28975 , \28674_28976 , \28675_28977 , \28676_28978 ,
         \28677_28979 , \28678_28980 , \28679_28981 , \28680_28982 , \28681_28983 , \28682_28984 , \28683_28985 , \28684_28986 , \28685_28987 , \28686_28988 ,
         \28687_28989 , \28688_28990 , \28689_28991 , \28690_28992 , \28691_28993 , \28692_28994 , \28693_28995 , \28694_28996 , \28695_28997 , \28696_28998 ,
         \28697_28999 , \28698_29000 , \28699_29001 , \28700_29002 , \28701_29003 , \28702_29004 , \28703_29005 , \28704_29006 , \28705_29007 , \28706_29008 ,
         \28707_29009 , \28708_29010 , \28709_29011 , \28710_29012 , \28711_29013 , \28712_29014 , \28713_29015 , \28714_29016 , \28715_29017 , \28716_29018 ,
         \28717_29019 , \28718_29020 , \28719_29021 , \28720_29022 , \28721_29023 , \28722_29024 , \28723_29025 , \28724_29026 , \28725_29027 , \28726_29028 ,
         \28727_29029 , \28728_29030 , \28729_29031 , \28730_29032 , \28731_29033 , \28732_29034 , \28733_29035 , \28734_29036 , \28735_29037 , \28736_29038 ,
         \28737_29039 , \28738_29040 , \28739_29041 , \28740_29042 , \28741_29043 , \28742_29044 , \28743_29045 , \28744_29046 , \28745_29047 , \28746_29048 ,
         \28747_29049 , \28748_29050 , \28749_29051 , \28750_29052 , \28751_29053 , \28752_29054 , \28753_29055 , \28754_29056 , \28755_29057 , \28756_29058 ,
         \28757_29059 , \28758_29060 , \28759_29061 , \28760_29062 , \28761_29063 , \28762_29064 , \28763 , \28764_29066_nG6152 , \28765_29067 , \28766_29068 ,
         \28767_29069 , \28768_29070 , \28769_29071 , \28770_29072 , \28771_29073 , \28772_29074 , \28773_29075 , \28774_29076 , \28775_29077 , \28776_29078 ,
         \28777_29079 , \28778_29080 , \28779 , \28780 , \28781_29083_nG65ca , \28782_29084 , \28783_29085 , \28784_29086 , \28785_29087 , \28786_29088 ,
         \28787_29089 , \28788_29090 , \28789_29091 , \28790_29092 , \28791_29093 , \28792_29094 , \28793_29095 , \28794_29096 , \28795_29097 , \28796_29098 ,
         \28797_29099 , \28798_29100 , \28799_29101 , \28800_29102 , \28801_29103 , \28802_29104 , \28803_29105 , \28804_29106 , \28805_29107 , \28806_29108 ,
         \28807_29109 , \28808_29110 , \28809_29111 , \28810_29112 , \28811_29113 , \28812_29114 , \28813_29115 , \28814_29116 , \28815_29117 , \28816_29118 ,
         \28817_29119 , \28818_29120 , \28819_29121 , \28820_29122 , \28821_29123 , \28822_29124 , \28823_29125 , \28824_29126 , \28825_29127 , \28826_29128 ,
         \28827_29129 , \28828_29130 , \28829_29131 , \28830_29132 , \28831_29133 , \28832_29134 , \28833_29135 , \28834_29136 , \28835_29137 , \28836_29138 ,
         \28837_29139 , \28838_29140 , \28839_29141 , \28840_29142 , \28841_29143 , \28842_29144 , \28843_29145 , \28844_29146 , \28845_29147 , \28846_29148 ,
         \28847_29149 , \28848_29150 , \28849_29151 , \28850_29152 , \28851_29153 , \28852_29154 , \28853_29155 , \28854_29156 , \28855_29157 , \28856_29158 ,
         \28857_29159 , \28858_29160 , \28859_29161 , \28860_29162 , \28861_29163 , \28862_29164 , \28863_29165 , \28864_29166 , \28865_29167 , \28866_29168 ,
         \28867_29169 , \28868_29170 , \28869_29171 , \28870_29172 , \28871_29173 , \28872_29174 , \28873_29175 , \28874_29176 , \28875_29177 , \28876_29178 ,
         \28877_29179_nG9bbd , \28878_29180 , \28879_29181 , \28880_29182 , \28881_29183 , \28882_29184 , \28883_29185 , \28884_29186 , \28885_29187 , \28886_29188 ,
         \28887_29189 , \28888_29190 , \28889_29191 , \28890_29192 , \28891_29193 , \28892_29194 , \28893_29195 , \28894_29196 , \28895_29197 , \28896_29198 ,
         \28897_29199 , \28898_29200 , \28899_29201 , \28900_29202 , \28901_29203 , \28902_29204 , \28903_29205 , \28904_29206 , \28905_29207 , \28906_29208 ,
         \28907_29209 , \28908_29210 , \28909_29211 , \28910_29212 , \28911_29213 , \28912_29214 , \28913_29215 , \28914_29216 , \28915_29217 , \28916_29218 ,
         \28917_29219 , \28918_29220 , \28919_29221 , \28920_29222 , \28921_29223 , \28922_29224 , \28923_29225 , \28924_29226 , \28925_29227 , \28926_29228 ,
         \28927_29229 , \28928_29230 , \28929_29231 , \28930_29232 , \28931_29233 , \28932_29234 , \28933_29235 , \28934_29236 , \28935_29237 , \28936_29238 ,
         \28937_29239 , \28938_29240 , \28939_29241 , \28940_29242 , \28941_29243 , \28942_29244 , \28943_29245 , \28944_28116 , \28945_28117 , \28946_28118 ,
         \28947_29246 , \28948_29247 , \28949_29248 , \28950_29249 , \28951_29250 , \28952_29251 , \28953_29252 , \28954_29253 , \28955_29254 , \28956_29255 ,
         \28957_29256 , \28958_29257 , \28959_29258 , \28960_29259 , \28961_29260 , \28962_29261 , \28963_29262 , \28964_29263 , \28965_29264 , \28966_29265 ,
         \28967_29266 , \28968_29267 , \28969_29268 , \28970_29269 , \28971_29270 , \28972_29271 , \28973_29272 , \28974_29273 , \28975_29274 , \28976_29275 ,
         \28977_29276 , \28978_29277 , \28979_29278 , \28980_29279 , \28981_29280 , \28982_29281 , \28983_29282 , \28984_29283 , \28985_29284 , \28986_29285 ,
         \28987_29286 , \28988_29287 , \28989_29288 , \28990_29289 , \28991_29290 , \28992_29291 , \28993_29292 , \28994_29293 , \28995_29294 , \28996_29295 ,
         \28997_29296 , \28998_29297 , \28999_29298 , \29000_29299 , \29001_29300 , \29002_29301 , \29003_29302 , \29004_29303 , \29005_29304 , \29006_29305 ,
         \29007_29306 , \29008_29307 , \29009_29308 , \29010_29309 , \29011_29310 , \29012_29311 , \29013_29312 , \29014_29313 , \29015_29314 , \29016_29315 ,
         \29017_29316 , \29018_29317 , \29019_29318 , \29020_29319 , \29021_29320 , \29022_29321 , \29023_29322 , \29024_29323 , \29025_29324 , \29026_29325 ,
         \29027_29326 , \29028_29327 , \29029_29328 , \29030_29329 , \29031_29330 , \29032_29331 , \29033_29332 , \29034_29333 , \29035_29334 , \29036_29335 ,
         \29037_29336 , \29038_29337 , \29039_29338 , \29040_29339 , \29041_29340 , \29042_29341 , \29043_29342 , \29044_29343 , \29045_29344 , \29046_29345 ,
         \29047_29346 , \29048_29347 , \29049_29348 , \29050_29349 , \29051_29350 , \29052_29351 , \29053_29352 , \29054_29353 , \29055_29354 , \29056_29355 ,
         \29057_29356 , \29058_29357 , \29059_29358 , \29060_29359 , \29061_29360 , \29062_29361 , \29063_29362 , \29064_29363 , \29065_29364 , \29066_29365 ,
         \29067_29366 , \29068_29367 , \29069_29368 , \29070_29369 , \29071_29370 , \29072_29371 , \29073_29372 , \29074_29373 , \29075_29374 , \29076_29375 ,
         \29077_29376 , \29078_29377 , \29079_29378 , \29080_29379 , \29081_29380 , \29082_29381 , \29083_29382 , \29084_29383 , \29085_29384 , \29086_29385 ,
         \29087_29386 , \29088_29387 , \29089_29388 , \29090_29389 , \29091_29390 , \29092_29391 , \29093_29392 , \29094_29393 , \29095_29394 , \29096_29395 ,
         \29097_29396 , \29098_29397 , \29099_29398 , \29100_29399 , \29101_29400 , \29102_29401 , \29103_29402 , \29104_29403 , \29105_29404 , \29106_29405 ,
         \29107_29406 , \29108_29407 , \29109_29408 , \29110_29409 , \29111_29410 , \29112_29411 , \29113_29412 , \29114_29413 , \29115_29414 , \29116_29415 ,
         \29117_29416 , \29118_29417 , \29119_29418 , \29120_29419 , \29121_29420 , \29122_29421 , \29123_29422 , \29124_29423 , \29125_29424 , \29126_29425 ,
         \29127_29426 , \29128_29427 , \29129_29428 , \29130_29429 , \29131_29430 , \29132_29431 , \29133_29432 , \29134 , \29135_29434 , \29136_29435 ,
         \29137_29436 , \29138_29437 , \29139_29438 , \29140_29439 , \29141_29440 , \29142_29441 , \29143_29442 , \29144_29443 , \29145_29444 , \29146_29445 ,
         \29147_29446 , \29148_29447 , \29149_29448 , \29150_29449 , \29151_29450 , \29152_29451 , \29153_29452 , \29154_29453 , \29155_29454 , \29156_29455 ,
         \29157_29456 , \29158_29457 , \29159_29458 , \29160_29459 , \29161_29460 , \29162_29461 , \29163_29462 , \29164_29463 , \29165_29464 , \29166_29465 ,
         \29167_29466 , \29168_29467 , \29169_29468 , \29170_29469 , \29171_29470 , \29172_29471 , \29173_29472 , \29174_29473 , \29175_29474 , \29176_29475 ,
         \29177_29476 , \29178_29477 , \29179_29478 , \29180_29479 , \29181_29480 , \29182_29481 , \29183_29482 , \29184_29483 , \29185_29484 , \29186_29485 ,
         \29187_29486 , \29188_29487 , \29189_29488 , \29190_29489 , \29191_29490 , \29192_29491 , \29193_29492 , \29194_29493 , \29195_29494 , \29196_29495 ,
         \29197_29496 , \29198_29497 , \29199_29498 , \29200_29499 , \29201_29500 , \29202_29501 , \29203_29502 , \29204_29503 , \29205_29504 , \29206_29505 ,
         \29207_29506 , \29208_29507 , \29209_29508 , \29210_29509 , \29211_29510 , \29212_29511 , \29213_29512 , \29214_29513 , \29215_29514 , \29216_29515 ,
         \29217_29516 , \29218_29517 , \29219_29518 , \29220_29519 , \29221_29520 , \29222_29521 , \29223_29522 , \29224_29523 , \29225_29524 , \29226_29525 ,
         \29227_29526 , \29228_29527 , \29229_29528 , \29230_29529 , \29231_29530 , \29232_29531 , \29233_29532 , \29234_29533 , \29235_29534 , \29236_29535 ,
         \29237_29536 , \29238_29537 , \29239_29538 , \29240_29539 , \29241_29540 , \29242_29541 , \29243_29542 , \29244_29543 , \29245_29544 , \29246_29545 ,
         \29247_29546 , \29248_29547 , \29249_29548 , \29250_29549 , \29251_29550 , \29252_29551 , \29253_29552 , \29254_29553 , \29255_29554 , \29256_29555 ,
         \29257_29556 , \29258_29557 , \29259_29558 , \29260_29559 , \29261_29560 , \29262_29561 , \29263_29562 , \29264_29563 , \29265_29564 , \29266_29565 ,
         \29267 , \29268_29567 , \29269_29568 , \29270_29569 , \29271_29570 , \29272_29571 , \29273_29572 , \29274_29573 , \29275_29574 , \29276_29575 ,
         \29277_29576 , \29278_29577 , \29279_29578 , \29280_29579 , \29281_29580 , \29282_29581 , \29283_29582 , \29284_29583 , \29285_29584 , \29286_29585 ,
         \29287_29586 , \29288_29587 , \29289_29588 , \29290_29589 , \29291_29590 , \29292_29591 , \29293_29592 , \29294_29593 , \29295_29594 , \29296_29595 ,
         \29297_29596 , \29298_29597 , \29299_29598 , \29300_29599 , \29301_29600 , \29302_29601 , \29303_29602 , \29304_29603 , \29305_29604 , \29306_29605 ,
         \29307_29606 , \29308_29607 , \29309_29608 , \29310_29609 , \29311_29610 , \29312_29611 , \29313_29612 , \29314_29613 , \29315_29614 , \29316_29615 ,
         \29317_29616 , \29318_29617 , \29319_29618 , \29320_29619 , \29321_29620 , \29322_29621 , \29323_29622 , \29324_29623 , \29325_29624 , \29326_29625 ,
         \29327_29626 , \29328_29627 , \29329_29628 , \29330_29629 , \29331_29630 , \29332_29631 , \29333_29632 , \29334_29633 , \29335_29634 , \29336_29635 ,
         \29337_29636 , \29338_29637 , \29339_29638 , \29340_29639 , \29341_29640 , \29342_29641 , \29343_29642 , \29344_29643 , \29345_29644 , \29346_29645 ,
         \29347_29646 , \29348_29647 , \29349_29648 , \29350_29649 , \29351_29650 , \29352_29651 , \29353_29652 , \29354_29653 , \29355_29654 , \29356_29655 ,
         \29357_29656 , \29358_29657 , \29359_29658 , \29360_29659 , \29361_29660 , \29362_29661 , \29363_29662 , \29364_29663 , \29365_29664 , \29366_29665 ,
         \29367_29666 , \29368_29667 , \29369_29668 , \29370_29669 , \29371_29670 , \29372_29671 , \29373_29672 , \29374_29673 , \29375_29674 , \29376_29675 ,
         \29377_29676 , \29378_29677 , \29379_29678 , \29380_29679 , \29381_29680 , \29382_29681 , \29383_29682 , \29384_29683 , \29385_29684 , \29386_29685 ,
         \29387_29686 , \29388_29687 , \29389_29688 , \29390_29689 , \29391_29690 , \29392_29691 , \29393_29692 , \29394_29693 , \29395_29694 , \29396_29695 ,
         \29397_29696 , \29398_29697 , \29399_29698 , \29400_29699 , \29401 , \29402_29701 , \29403_29702 , \29404_29703 , \29405_29704 , \29406_29705 ,
         \29407_29706 , \29408_29707 , \29409_29708 , \29410_29709 , \29411_29710 , \29412_29711 , \29413_29712 , \29414_29713 , \29415_29714 , \29416_29715 ,
         \29417_29716 , \29418_29717 , \29419_29718 , \29420_29719 , \29421_29720 , \29422_29721 , \29423_29722 , \29424_29723 , \29425_29724 , \29426_29725 ,
         \29427_29726 , \29428_29727 , \29429_29728 , \29430_29729 , \29431_29730 , \29432_29731 , \29433_29732 , \29434_29733 , \29435_29734 , \29436_29735 ,
         \29437_29736 , \29438_29737 , \29439_29738 , \29440_29739 , \29441_29740 , \29442_29741 , \29443_29742 , \29444_29743 , \29445_29744 , \29446_29745 ,
         \29447_29746 , \29448_29747 , \29449_29748 , \29450_29749 , \29451_29750 , \29452_29751 , \29453_29752 , \29454_29753 , \29455_29754 , \29456_29755 ,
         \29457_29756 , \29458_29757 , \29459_29758 , \29460_29759 , \29461_29760 , \29462_29761 , \29463_29762 , \29464_29763 , \29465_29764 , \29466_29765 ,
         \29467_29766 , \29468_29767 , \29469_29768 , \29470_29769 , \29471_29770 , \29472_29771 , \29473_29772 , \29474_29773 , \29475_29774 , \29476_29775 ,
         \29477_29776 , \29478_29777 , \29479_29778 , \29480_29779 , \29481_29780 , \29482_29781 , \29483_29782 , \29484_29783 , \29485_29784 , \29486_29785 ,
         \29487_29786 , \29488_29787 , \29489_29788 , \29490_29789 , \29491_29790 , \29492_29791 , \29493_29792 , \29494_29793 , \29495_29794 , \29496_29795 ,
         \29497_29796 , \29498_29797 , \29499_29798 , \29500_29799 , \29501_29800 , \29502_29801 , \29503_29802 , \29504_29803 , \29505_29804 , \29506_29805 ,
         \29507_29806 , \29508_29807 , \29509_29808 , \29510_29809 , \29511_29810 , \29512_29811 , \29513_29812 , \29514_29813 , \29515_29814 , \29516_29815 ,
         \29517_29816 , \29518_29817 , \29519_29818 , \29520_29819 , \29521_29820 , \29522_29821 , \29523_29822 , \29524_29823 , \29525_29824 , \29526_29825 ,
         \29527_29826 , \29528_29827 , \29529_29828 , \29530_29829 , \29531_29830 , \29532_29831 , \29533_29832 , \29534 , \29535_29834 , \29536_29835 ,
         \29537_29836 , \29538_29837 , \29539_29838 , \29540_29839 , \29541_29840 , \29542_29841 , \29543_29842 , \29544_29843 , \29545_29844_nG4400 , \29546_29845 ,
         \29547_29846 , \29548_29847_nG4403 , \29549_29848 , \29550_29849 , \29551_29850 , \29552_29854 , \29553_29855 , \29554_29856 , \29555_29857 , \29556_29858 ,
         \29557_29859 , \29558_29860 , \29559_29861 , \29560_29862 , \29561_29863 , \29562_29864 , \29563_29865 , \29564_29866 , \29565_29867 , \29566_29868 ,
         \29567_29869 , \29568_29870 , \29569_29871 , \29570_29872 , \29571_29873 , \29572_29874 , \29573_29875 , \29574_29876 , \29575_29877 , \29576_29878 ,
         \29577_29879 , \29578_29880 , \29579_29881 , \29580_29882 , \29581_29883 , \29582_29884 , \29583_29885 , \29584_29886 , \29585_29887 , \29586_29888 ,
         \29587_29889 , \29588_29890 , \29589_29891 , \29590_29892 , \29591_29893 , \29592_29894 , \29593_29895 , \29594_29896 , \29595_29897 , \29596_29898 ,
         \29597_29899 , \29598_29900 , \29599_29901 , \29600_29902 , \29601_29903 , \29602_29904 , \29603_29905 , \29604_29906 , \29605_29907 , \29606_29908 ,
         \29607_29909 , \29608_29910 , \29609_29911 , \29610_29912 , \29611_29913 , \29612_29914 , \29613_29915 , \29614_29916 , \29615_29917 , \29616_29918 ,
         \29617_29919 , \29618_29920 , \29619_29921 , \29620_29922 , \29621_29923 , \29622_29924 , \29623_29925 , \29624_29926 , \29625_29927 , \29626_29928 ,
         \29627_29929 , \29628_29930 , \29629_29931 , \29630_29932 , \29631_29933 , \29632_29934 , \29633_29935 , \29634_29936 , \29635_29937 , \29636_29938 ,
         \29637_29939 , \29638_29940 , \29639_29941 , \29640_29942 , \29641_29943 , \29642_29944 , \29643_29945 , \29644_29946 , \29645_29947 , \29646_29948 ,
         \29647_29949 , \29648_29950 , \29649_29951 , \29650_29952 , \29651_29953 , \29652_29954 , \29653_29955 , \29654_29956 , \29655_29957 , \29656_29958 ,
         \29657_29959 , \29658_29960 , \29659_29961 , \29660_29962 , \29661_29963 , \29662_29964 , \29663_29965 , \29664_29966 , \29665_29967 , \29666_29968 ,
         \29667_29969 , \29668_29970 , \29669_29971 , \29670_29972 , \29671_29973 , \29672_29974 , \29673_29975 , \29674_29976 , \29675_29977 , \29676_29978 ,
         \29677_29979 , \29678_29980 , \29679_29981 , \29680_29982 , \29681_29983 , \29682_29984 , \29683_29985 , \29684_29986 , \29685_29987 , \29686_29988 ,
         \29687_29989 , \29688_29990 , \29689_29991 , \29690_29992 , \29691_29993 , \29692_29994 , \29693_29995 , \29694_29996 , \29695_29997 , \29696_29998 ,
         \29697_29999 , \29698_30000 , \29699_30001 , \29700_30002 , \29701_30003 , \29702_30004 , \29703_30005 , \29704_30006 , \29705_30007 , \29706_30008 ,
         \29707_30009 , \29708_30010 , \29709_30011 , \29710_30012 , \29711_30013 , \29712_30014 , \29713_30015 , \29714_30016 , \29715_30017 , \29716_30018 ,
         \29717_30019 , \29718_30020 , \29719_30021 , \29720_30022 , \29721_30023 , \29722_30024 , \29723_30025 , \29724_30026 , \29725_30027 , \29726_30028 ,
         \29727_30029 , \29728_30030 , \29729_30031 , \29730_30032 , \29731_30033 , \29732_30034 , \29733_30035 , \29734_30036 , \29735_30037 , \29736_30038 ,
         \29737_30039 , \29738_30040 , \29739_30041 , \29740_30042 , \29741_30043 , \29742_30044 , \29743_30045 , \29744_30046 , \29745_30047 , \29746_30048 ,
         \29747_30049 , \29748_30050 , \29749_30051 , \29750_30052 , \29751_30053 , \29752_30054 , \29753_30055 , \29754_30056 , \29755_30057 , \29756_30058 ,
         \29757_30059 , \29758_30060 , \29759_30061 , \29760_30062 , \29761_30063 , \29762_30064 , \29763_30065 , \29764_30066 , \29765_30067 , \29766_30068 ,
         \29767_30069 , \29768_30070 , \29769_30071 , \29770_30072 , \29771_30073 , \29772_30074 , \29773_30075 , \29774_30076 , \29775_30077 , \29776_30078 ,
         \29777_30079 , \29778_30080 , \29779_30081 , \29780_30082 , \29781_30083 , \29782_30084 , \29783_30085 , \29784_30086 , \29785_30087 , \29786_30088 ,
         \29787_30089 , \29788_30090 , \29789_30091 , \29790_30092 , \29791_30093 , \29792_30094 , \29793_30095 , \29794_30096 , \29795_30097 , \29796_30098 ,
         \29797_30099 , \29798_30100 , \29799_30101 , \29800_30102 , \29801_30103 , \29802_30104 , \29803_30105 , \29804_30106 , \29805_30107 , \29806_30108 ,
         \29807_30109 , \29808_30110 , \29809 , \29810_30112 , \29811_30113 , \29812_30114 , \29813_30115 , \29814_30116 , \29815_30117 , \29816_30118 ,
         \29817_30119 , \29818_30120 , \29819_30121 , \29820_30122 , \29821_30123 , \29822_30124 , \29823_30125 , \29824_30126 , \29825_30127 , \29826_30128 ,
         \29827_30129 , \29828_30130 , \29829_30131 , \29830_30132 , \29831_30133 , \29832_30134 , \29833_30135 , \29834_30136 , \29835_30137 , \29836_30138 ,
         \29837_30139 , \29838_30140 , \29839_30141 , \29840_30142 , \29841_30143 , \29842_30144 , \29843_30145 , \29844_30146 , \29845_30147 , \29846_30148 ,
         \29847_30149 , \29848_30150 , \29849_30151 , \29850_30152 , \29851_30153 , \29852_30154 , \29853_30155 , \29854_30156 , \29855_30157 , \29856_30158 ,
         \29857_30159 , \29858_30160 , \29859_30161 , \29860_30162 , \29861_30163 , \29862_30164 , \29863_30165 , \29864_30166 , \29865_30167 , \29866_30168 ,
         \29867_30169 , \29868_30170 , \29869_30171 , \29870_30172 , \29871_30173 , \29872_30174 , \29873_30175 , \29874_30176 , \29875_30177 , \29876_30178 ,
         \29877_30179 , \29878_30180 , \29879_30181 , \29880_30182 , \29881_30183 , \29882_30184 , \29883_30185 , \29884_30186 , \29885_30187 , \29886_30188 ,
         \29887_30189 , \29888_30190 , \29889_30191 , \29890_30192 , \29891_30193 , \29892_30194 , \29893_30195 , \29894_30196 , \29895_30197 , \29896_30198 ,
         \29897_30199 , \29898_30200 , \29899_30201 , \29900_30202 , \29901_30203 , \29902_30204 , \29903_30205 , \29904_30206 , \29905_30207 , \29906_30208 ,
         \29907_30209 , \29908_30210 , \29909_30211 , \29910_30212 , \29911_30213 , \29912_30214 , \29913_30215 , \29914_30216 , \29915_30217 , \29916_30218 ,
         \29917_30219 , \29918_30220 , \29919_30221 , \29920_30222 , \29921_30223 , \29922_30224 , \29923_30225 , \29924_30226 , \29925_30227 , \29926_30228 ,
         \29927_30229 , \29928_30230 , \29929_30231 , \29930_30232 , \29931_30233 , \29932_30234 , \29933_30235 , \29934_30236 , \29935_30237 , \29936_30238 ,
         \29937_30239 , \29938_30240 , \29939_30241 , \29940_30242 , \29941 , \29942_30244_nG625b , \29943_30245 , \29944_30246 , \29945_30247 , \29946_30248 ,
         \29947_30249 , \29948_30250 , \29949_30251 , \29950_30252 , \29951_30253 , \29952_30254 , \29953_30255 , \29954_30256 , \29955_30257 , \29956_30258 ,
         \29957_30259 , \29958_30260 , \29959_30261 , \29960_30262 , \29961_30263 , \29962_30264 , \29963 , \29964 , \29965_30267_nG65cd , \29966_30268 ,
         \29967_30269 , \29968_30270 , \29969_30271 , \29970_30272 , \29971_30273 , \29972_30274 , \29973_30275 , \29974_30276 , \29975_30277 , \29976_30278 ,
         \29977_30279 , \29978_30280 , \29979_30281 , \29980_30282 , \29981_30283 , \29982_30284 , \29983_30285 , \29984_30286 , \29985_30287 , \29986_30288 ,
         \29987_30289 , \29988_30290 , \29989_30291 , \29990_30292 , \29991_30293 , \29992_30294 , \29993_30295 , \29994_30296 , \29995_30297 , \29996_30298 ,
         \29997_30299 , \29998_30300 , \29999_30301 , \30000_30302 , \30001_30303 , \30002_30304 , \30003_30305 , \30004_30306 , \30005_30307 , \30006_30308 ,
         \30007_30309 , \30008_30310 , \30009_30311 , \30010_30312 , \30011_30313 , \30012_30314 , \30013_30315 , \30014_30316 , \30015_30317 , \30016_30318 ,
         \30017_30319 , \30018_30320 , \30019_30321 , \30020_30322 , \30021_30323 , \30022_30324 , \30023_30325 , \30024_30326 , \30025_30327 , \30026_30328 ,
         \30027_30329 , \30028_30330 , \30029_30331 , \30030_30332 , \30031_30333 , \30032_30334 , \30033_30335 , \30034_30336 , \30035_30337 , \30036_30338 ,
         \30037_30339 , \30038_30340 , \30039_30341 , \30040_30342 , \30041_30343 , \30042_30344 , \30043_30345 , \30044_30346 , \30045_30347 , \30046_30348 ,
         \30047_30349 , \30048_30350 , \30049_30351 , \30050_30352 , \30051_30353 , \30052_30354 , \30053_30355 , \30054_30356 , \30055_30357 , \30056_30358 ,
         \30057_30359 , \30058_30360 , \30059_30361 , \30060_30362 , \30061_30363 , \30062_30364 , \30063_30365 , \30064_30366_nG9bba , \30065_30367 , \30066_30368 ,
         \30067_30369 , \30068_30370 , \30069_30371 , \30070_30372 , \30071_30373 , \30072_30374 , \30073_30375 , \30074_30376 , \30075_30377 , \30076_30378 ,
         \30077_30379 , \30078_30380 , \30079_30381 , \30080_30382 , \30081_30383 , \30082_30384 , \30083_30385 , \30084_30386 , \30085_30387 , \30086_30388 ,
         \30087_30389 , \30088_30390 , \30089_30391 , \30090_30392 , \30091_30393 , \30092_30394 , \30093_30395 , \30094_30396 , \30095_30397 , \30096_30398 ,
         \30097_30399 , \30098_30400 , \30099_30401 , \30100_30402 , \30101_30403 , \30102_30404 , \30103_30405 , \30104_30406 , \30105_30407 , \30106_30408 ,
         \30107_30409 , \30108_30410 , \30109_30411 , \30110_30412 , \30111_30413 , \30112_30414 , \30113_30415 , \30114_30416 , \30115_30417 , \30116_30418 ,
         \30117_30419 , \30118_30420 , \30119_30421 , \30120_30422 , \30121_30423 , \30122_30424 , \30123_30425 , \30124_30426 , \30125_30427 , \30126_30428 ,
         \30127_30429 , \30128_30430 , \30129_30431 , \30130_30432 , \30131_30433 , \30132_30434 , \30133_30435 , \30134_30436 , \30135_30437 , \30136_30438 ,
         \30137_30439 , \30138_30440 , \30139_30441 , \30140_30442 , \30141_30443 , \30142_30444 , \30143_30445 , \30144_30446 , \30145_30447 , \30146_30448 ,
         \30147_30449 , \30148_30450 , \30149_30451 , \30150_30452 , \30151_30453 , \30152_30454 , \30153_30455 , \30154_30456 , \30155_30457 , \30156_30458 ,
         \30157_30459 , \30158_30460 , \30159_30461 , \30160_30462 , \30161_30463 , \30162_30464 , \30163_30465 , \30164_30466 , \30165_30467 , \30166_30468 ,
         \30167_30469 , \30168_30470 , \30169_30471 , \30170_30472 , \30171_30473 , \30172_30474 , \30173_30475 , \30174_30476 , \30175_30477 , \30176_30478 ,
         \30177_30479 , \30178_30480 , \30179_30481 , \30180_30482 , \30181_30483 , \30182_30484 , \30183_30485 , \30184_30486 , \30185_30487 , \30186_30488 ,
         \30187_30489 , \30188_30490 , \30189_30491 , \30190_30492 , \30191_30493 , \30192_30494 , \30193_30495 , \30194_30496 , \30195_30497 , \30196_30498 ,
         \30197_30499 , \30198_30500 , \30199_30501 , \30200_30502 , \30201_30503 , \30202_30504 , \30203_30505 , \30204_30506 , \30205_30507 , \30206_30508 ,
         \30207_30509 , \30208_30510 , \30209_30511 , \30210_30512 , \30211_30513 , \30212_30514 , \30213_30515 , \30214_30516 , \30215_30517 , \30216_30518 ,
         \30217_30519 , \30218_30520 , \30219_30521 , \30220_30522 , \30221_30523 , \30222_30524 , \30223_30525 , \30224_30526 , \30225_30527 , \30226_30528 ,
         \30227_30529 , \30228_30530 , \30229_30531 , \30230_30532 , \30231_30533 , \30232_30534 , \30233_30535 , \30234_30536 , \30235_30537 , \30236_30538 ,
         \30237_30539 , \30238_30540 , \30239_30541 , \30240_30542 , \30241_30543 , \30242_30544 , \30243_30545 , \30244_30546 , \30245_30547 , \30246_30548 ,
         \30247_30549 , \30248_30550 , \30249_30551 , \30250_30552 , \30251_30553 , \30252_30554 , \30253_30555 , \30254_30556 , \30255_30557 , \30256_30558 ,
         \30257_30559 , \30258_30560 , \30259_30561 , \30260_30562 , \30261_30563 , \30262_30564 , \30263_30565 , \30264_30566 , \30265_30567 , \30266_30568 ,
         \30267_30569 , \30268_30570 , \30269_30571 , \30270_30572 , \30271_30573 , \30272_30574 , \30273_30575 , \30274_30576 , \30275_30577 , \30276_30578 ,
         \30277_30579 , \30278_30580 , \30279_30581 , \30280_30582 , \30281_30583 , \30282_30584 , \30283_30585 , \30284_30586 , \30285_30587 , \30286_30588 ,
         \30287_30589 , \30288_30590 , \30289_30591 , \30290_30592 , \30291_30593 , \30292_30594 , \30293_30595 , \30294_30596 , \30295_30597 , \30296_30598 ,
         \30297_30599 , \30298_30600 , \30299_30601 , \30300_30602 , \30301_30603 , \30302_30604 , \30303_30605 , \30304_30606 , \30305_30607 , \30306_30608 ,
         \30307_30609 , \30308_30610 , \30309_30611 , \30310_30612 , \30311_30613 , \30312_30614 , \30313_30615 , \30314_30616 , \30315_30617 , \30316_30618 ,
         \30317_30619 , \30318_30620 , \30319_30621 , \30320_30622 , \30321_30623 , \30322_30624 , \30323_30625 , \30324_30626 , \30325_30627 , \30326_30628 ,
         \30327_30629 , \30328_30630 , \30329_30631 , \30330_30632 , \30331_30633 , \30332_30634 , \30333_30635 , \30334_30636 , \30335_30637 , \30336_30638 ,
         \30337_30639 , \30338_30640 , \30339_30641 , \30340_30642 , \30341_30643 , \30342_30644 , \30343_30645 , \30344_30646 , \30345_30647 , \30346_30648 ,
         \30347_30649 , \30348_30650 , \30349_30651 , \30350_30652 , \30351_30653 , \30352_30654 , \30353_30655 , \30354_30656 , \30355_30657 , \30356_30658 ,
         \30357_30659 , \30358_30660 , \30359_30661 , \30360_30662 , \30361_30663 , \30362_30664 , \30363_30665 , \30364_30666 , \30365_30667 , \30366 ,
         \30367_30669 , \30368_30670 , \30369_30671 , \30370_30672 , \30371_30673 , \30372_30674 , \30373_30675 , \30374_30676 , \30375_30677 , \30376_30678 ,
         \30377_30679 , \30378_30680 , \30379_30681 , \30380_30682 , \30381_30683 , \30382_30684 , \30383_30685 , \30384_30686 , \30385_30687 , \30386_30688 ,
         \30387_30689 , \30388_30690 , \30389_30691 , \30390_30692 , \30391_30693 , \30392_30694 , \30393_30695 , \30394_30696 , \30395_30697 , \30396_30698 ,
         \30397_30699 , \30398_30700 , \30399_30701 , \30400_30702 , \30401_30703 , \30402_30704 , \30403_30705 , \30404_30706 , \30405_30707 , \30406_30708 ,
         \30407_30709 , \30408_30710 , \30409_30711 , \30410_30712 , \30411_30713 , \30412_30714 , \30413_30715 , \30414_30716 , \30415_30717 , \30416_30718 ,
         \30417_30719 , \30418_30720 , \30419_30721 , \30420_30722 , \30421_30723 , \30422_30724 , \30423_30725 , \30424_30726 , \30425_30727 , \30426_30728 ,
         \30427_30729 , \30428_30730 , \30429_30731 , \30430_30732 , \30431_30733 , \30432_30734 , \30433_30735 , \30434_30736 , \30435_30737 , \30436_30738 ,
         \30437_30739 , \30438_30740 , \30439_30741 , \30440_30742 , \30441_30743 , \30442_30744 , \30443_30745 , \30444_30746 , \30445_30747 , \30446_30748 ,
         \30447_30749 , \30448_30750 , \30449_30751 , \30450_30752 , \30451_30753 , \30452_30754 , \30453_30755 , \30454_30756 , \30455_30757 , \30456_30758 ,
         \30457_30759 , \30458_30760 , \30459_30761 , \30460_30762 , \30461_30763 , \30462_30764 , \30463_30765 , \30464_30766 , \30465_30767 , \30466_30768 ,
         \30467_30769 , \30468_30770 , \30469_30771 , \30470_30772 , \30471_30773 , \30472_30774 , \30473_30775 , \30474_30776 , \30475_30777 , \30476_30778 ,
         \30477_30779 , \30478_30780 , \30479_30781 , \30480_30782 , \30481_30783 , \30482_30784 , \30483_30785 , \30484_30786 , \30485_30787 , \30486_30788 ,
         \30487_30789 , \30488_30790 , \30489_30791 , \30490_30792 , \30491_30793 , \30492_30794 , \30493_30795 , \30494_30796 , \30495_30797 , \30496_30798 ,
         \30497_30799 , \30498 , \30499_30801_nG65d0 , \30500_30802 , \30501_30803 , \30502_30804 , \30503_30805 , \30504_30806 , \30505 , \30506 ,
         \30507_30809_nG6364 , \30508_30810 , \30509_30811 , \30510_30812 , \30511_30813 , \30512_30814 , \30513_30815 , \30514_30816 , \30515_30817 , \30516_30818 ,
         \30517_30819 , \30518_30820 , \30519_30821 , \30520_30822 , \30521_30823 , \30522_30824 , \30523_30825 , \30524_30826 , \30525_30827 , \30526_30828 ,
         \30527_30829 , \30528_30830 , \30529_30831 , \30530_30832 , \30531_30833 , \30532_30834 , \30533_30835 , \30534_30836 , \30535_30837 , \30536_30838 ,
         \30537_30839 , \30538_30840 , \30539_30841 , \30540_30842 , \30541_30843 , \30542_30844 , \30543_30845 , \30544_30846 , \30545_30847 , \30546_30848 ,
         \30547_30849 , \30548_30850 , \30549_30851 , \30550_30852 , \30551_30853 , \30552_30854 , \30553_30855 , \30554_30856 , \30555_30857 , \30556_30858 ,
         \30557_30859 , \30558_30860 , \30559_30861 , \30560_30862 , \30561_30863 , \30562_30864 , \30563_30865 , \30564_30866 , \30565_30867 , \30566_30868 ,
         \30567_30869 , \30568_30870 , \30569_30871 , \30570_30872 , \30571_30873 , \30572_30874 , \30573_30875 , \30574_30876 , \30575_30877 , \30576_30878 ,
         \30577_30879 , \30578_30880 , \30579_30881 , \30580_30882 , \30581_30883 , \30582_30884 , \30583_30885 , \30584_30886 , \30585_30887 , \30586_30888 ,
         \30587_30889 , \30588_30890 , \30589_30891 , \30590_30892 , \30591_30893 , \30592_30894 , \30593_30895 , \30594_30896 , \30595_30897 , \30596_30898 ,
         \30597_30899 , \30598_30900 , \30599_30901 , \30600_30902 , \30601_30903 , \30602_30904 , \30603_30905 , \30604_30906 , \30605_30907 , \30606_30908 ,
         \30607_30909 , \30608_30910 , \30609_30911 , \30610_30912 , \30611_30913 , \30612_30914 , \30613_30915 , \30614_30916 , \30615_30917 , \30616_30918 ,
         \30617_30919 , \30618_30920 , \30619_30921 , \30620_30922 , \30621_30923 , \30622_30924 , \30623_30925 , \30624_30926 , \30625_30927 , \30626_30928 ,
         \30627_30929 , \30628_30930 , \30629_30931 , \30630_30932 , \30631_30933 , \30632_30934 , \30633_30935 , \30634_30936 , \30635_30937 , \30636_30938 ,
         \30637_30939 , \30638_30940_nG9bb7 , \30639_30941 , \30640_30942 , \30641_30943 , \30642_30944 , \30643_30945 , \30644_30946 , \30645_30947 , \30646_30948 ,
         \30647_30949 , \30648_30950 , \30649_30951 , \30650_30952 , \30651_30953 , \30652_30954 , \30653_30955 , \30654_30956 , \30655_30957 , \30656_30958 ,
         \30657_30959 , \30658_30960 , \30659_30961 , \30660_30962 , \30661_30963 , \30662_30964 , \30663_30965 , \30664_30966 , \30665_30967 , \30666_30968 ,
         \30667_30969 , \30668_29851 , \30669_29852 , \30670_29853 , \30671_30970 , \30672_30971 , \30673_30972 , \30674_30973 , \30675_30974 , \30676_30975 ,
         \30677_30976 , \30678_30977 , \30679_30978 , \30680_30979 , \30681_30980 , \30682_30981 , \30683_30982 , \30684_30983 , \30685_30984 , \30686_30985 ,
         \30687_30986 , \30688_30987 , \30689_30988 , \30690_30989 , \30691_30990 , \30692_30991 , \30693_30992 , \30694_30993 , \30695_30994 , \30696_30995 ,
         \30697_30996 , \30698_30997 , \30699_30998 , \30700_30999 , \30701_31000 , \30702_31001 , \30703_31002 , \30704_31003 , \30705_31004 , \30706_31005 ,
         \30707_31006 , \30708_31007 , \30709_31008 , \30710_31009 , \30711_31010 , \30712_31011 , \30713_31012 , \30714_31013 , \30715_31014 , \30716_31015 ,
         \30717_31016 , \30718_31017 , \30719_31018 , \30720_31019 , \30721_31020 , \30722_31021 , \30723_31022 , \30724_31023 , \30725_31024 , \30726_31025 ,
         \30727_31026 , \30728_31027 , \30729_31028 , \30730_31029 , \30731_31030 , \30732_31031 , \30733_31032 , \30734_31033 , \30735_31034 , \30736_31035 ,
         \30737_31036 , \30738_31037 , \30739_31038 , \30740_31039 , \30741_31040 , \30742_31041 , \30743_31042 , \30744_31043 , \30745_31044 , \30746_31045 ,
         \30747_31046 , \30748_31047 , \30749_31048 , \30750_31049 , \30751_31050 , \30752_31051 , \30753_31052 , \30754_31053 , \30755_31054 , \30756_31055 ,
         \30757_31056 , \30758_31057 , \30759_31058 , \30760_31059 , \30761_31060 , \30762_31061 , \30763_31062 , \30764_31063 , \30765_31064 , \30766_31065 ,
         \30767_31066 , \30768_31067 , \30769_31068 , \30770_31069 , \30771_31070 , \30772_31071 , \30773_31072 , \30774_31073 , \30775_31074 , \30776_31075 ,
         \30777_31076 , \30778_31077 , \30779_31078 , \30780_31079 , \30781_31080 , \30782_31081 , \30783_31082 , \30784_31083 , \30785_31084 , \30786_31085 ,
         \30787_31086 , \30788_31087 , \30789_31088 , \30790_31089 , \30791_31090 , \30792_31091 , \30793_31092 , \30794_31093 , \30795_31094 , \30796_31095 ,
         \30797_31096 , \30798_31097 , \30799_31098 , \30800_31099 , \30801_31100 , \30802_31101 , \30803_31102 , \30804_31103 , \30805_31104 , \30806_31105 ,
         \30807_31106 , \30808_31107 , \30809_31108 , \30810_31109 , \30811_31110 , \30812_31111 , \30813_31112 , \30814_31113 , \30815_31114 , \30816_31115 ,
         \30817_31116 , \30818_31117 , \30819_31118 , \30820_31119 , \30821_31120 , \30822_31121 , \30823_31122 , \30824_31123 , \30825_31124 , \30826_31125 ,
         \30827_31126 , \30828_31127 , \30829_31128 , \30830_31129 , \30831_31130 , \30832_31131 , \30833_31132 , \30834_31133 , \30835_31134 , \30836_31135 ,
         \30837_31136 , \30838_31137 , \30839_31138 , \30840_31139 , \30841_31140 , \30842_31141 , \30843_31142 , \30844_31143 , \30845_31144 , \30846_31145 ,
         \30847_31146 , \30848_31147 , \30849_31148 , \30850_31149 , \30851_31150 , \30852_31151 , \30853_31152 , \30854_31153 , \30855_31154 , \30856_31155 ,
         \30857_31156 , \30858_31157 , \30859_31158 , \30860_31159 , \30861_31160 , \30862_31161 , \30863_31162 , \30864_31163 , \30865_31164 , \30866_31165 ,
         \30867_31166 , \30868_31167 , \30869_31168 , \30870_31169 , \30871_31170 , \30872_31171 , \30873_31172 , \30874_31173 , \30875_31174 , \30876_31175 ,
         \30877_31176 , \30878_31177 , \30879_31178 , \30880_31179 , \30881_31180 , \30882_31181 , \30883_31182 , \30884_31183 , \30885_31184 , \30886_31185 ,
         \30887_31186 , \30888_31187 , \30889_31188 , \30890_31189 , \30891_31190 , \30892_31191 , \30893_31192 , \30894_31193 , \30895_31194 , \30896_31195 ,
         \30897_31196 , \30898_31197 , \30899_31198 , \30900_31199 , \30901_31200 , \30902_31201 , \30903_31202 , \30904_31203 , \30905_31204 , \30906_31205 ,
         \30907_31206 , \30908_31207 , \30909_31208 , \30910_31209 , \30911_31210 , \30912_31211 , \30913_31212 , \30914_31213 , \30915_31214 , \30916_31215 ,
         \30917 , \30918_31217 , \30919_31218 , \30920_31219 , \30921_31220 , \30922_31221 , \30923_31222 , \30924_31223 , \30925_31224 , \30926_31225 ,
         \30927_31226 , \30928_31227 , \30929_31228 , \30930_31229 , \30931_31230 , \30932_31231 , \30933_31232 , \30934_31233 , \30935_31234 , \30936_31235 ,
         \30937_31236 , \30938_31237 , \30939_31238 , \30940_31239 , \30941_31240 , \30942_31241 , \30943_31242 , \30944_31243 , \30945_31244 , \30946_31245 ,
         \30947_31246 , \30948_31247 , \30949_31248 , \30950_31249 , \30951_31250 , \30952_31251 , \30953_31252 , \30954_31253 , \30955_31254 , \30956_31255 ,
         \30957_31256 , \30958_31257 , \30959_31258 , \30960_31259 , \30961_31260 , \30962_31261 , \30963_31262 , \30964_31263 , \30965_31264 , \30966_31265 ,
         \30967_31266 , \30968_31267 , \30969_31268 , \30970_31269 , \30971_31270 , \30972_31271 , \30973_31272 , \30974_31273 , \30975_31274 , \30976_31275 ,
         \30977_31276 , \30978_31277 , \30979_31278 , \30980_31279 , \30981_31280 , \30982_31281 , \30983_31282 , \30984_31283 , \30985_31284 , \30986_31285 ,
         \30987_31286 , \30988_31287 , \30989_31288 , \30990_31289 , \30991_31290 , \30992_31291 , \30993_31292 , \30994_31293 , \30995_31294 , \30996_31295 ,
         \30997_31296 , \30998_31297 , \30999_31298 , \31000_31299 , \31001_31300 , \31002_31301 , \31003_31302 , \31004_31303 , \31005_31304 , \31006_31305 ,
         \31007_31306 , \31008_31307 , \31009_31308 , \31010_31309 , \31011_31310 , \31012_31311 , \31013_31312 , \31014_31313 , \31015_31314 , \31016_31315 ,
         \31017_31316 , \31018_31317 , \31019_31318 , \31020_31319 , \31021_31320 , \31022_31321 , \31023_31322 , \31024_31323 , \31025_31324 , \31026_31325 ,
         \31027_31326 , \31028_31327 , \31029_31328 , \31030_31329 , \31031_31330 , \31032_31331 , \31033_31332 , \31034_31333 , \31035_31334 , \31036_31335 ,
         \31037_31336 , \31038_31337 , \31039_31338 , \31040_31339 , \31041_31340 , \31042_31341 , \31043_31342 , \31044_31343 , \31045_31344 , \31046_31345 ,
         \31047_31346 , \31048_31347 , \31049_31348 , \31050 , \31051_31350 , \31052_31351 , \31053_31352 , \31054_31353 , \31055_31354 , \31056_31355 ,
         \31057_31356 , \31058_31357 , \31059_31358 , \31060_31359 , \31061_31360 , \31062_31361 , \31063_31362 , \31064_31363 , \31065_31364 , \31066_31365 ,
         \31067_31366 , \31068_31367 , \31069_31368 , \31070_31369 , \31071_31370 , \31072_31371 , \31073_31372 , \31074_31373 , \31075_31374 , \31076_31375 ,
         \31077_31376 , \31078_31377 , \31079_31378 , \31080_31379 , \31081_31380 , \31082_31381 , \31083_31382 , \31084_31383 , \31085_31384 , \31086_31385 ,
         \31087_31386 , \31088_31387 , \31089_31388 , \31090_31389 , \31091_31390 , \31092_31391 , \31093_31392 , \31094_31393 , \31095_31394 , \31096_31395 ,
         \31097_31396 , \31098_31397 , \31099_31398 , \31100_31399 , \31101_31400 , \31102_31401 , \31103_31402 , \31104_31403 , \31105_31404 , \31106_31405 ,
         \31107_31406 , \31108_31407 , \31109_31408 , \31110_31409 , \31111_31410 , \31112_31411 , \31113_31412 , \31114_31413 , \31115_31414 , \31116_31415 ,
         \31117_31416 , \31118_31417 , \31119_31418 , \31120_31419 , \31121_31420 , \31122_31421 , \31123_31422 , \31124_31423 , \31125_31424 , \31126_31425 ,
         \31127_31426 , \31128_31427 , \31129_31428 , \31130_31429 , \31131_31430 , \31132_31431 , \31133_31432 , \31134_31433 , \31135_31434 , \31136_31435 ,
         \31137_31436 , \31138_31437 , \31139_31438 , \31140_31439 , \31141_31440 , \31142_31441 , \31143_31442 , \31144_31443 , \31145_31444 , \31146_31445 ,
         \31147_31446 , \31148_31447 , \31149_31448 , \31150_31449 , \31151_31450 , \31152_31451 , \31153_31452 , \31154_31453 , \31155_31454 , \31156_31455 ,
         \31157_31456 , \31158_31457 , \31159_31458 , \31160_31459 , \31161_31460 , \31162_31461 , \31163_31462 , \31164_31463 , \31165_31464 , \31166_31465 ,
         \31167_31466 , \31168_31467 , \31169_31468 , \31170_31469 , \31171_31470 , \31172_31471 , \31173_31472 , \31174_31473 , \31175_31474 , \31176_31475 ,
         \31177_31476 , \31178_31477 , \31179_31478 , \31180_31479 , \31181_31480 , \31182_31481 , \31183_31482 , \31184 , \31185_31484 , \31186_31485 ,
         \31187_31486 , \31188_31487 , \31189_31488 , \31190_31489 , \31191_31490 , \31192_31491 , \31193_31492 , \31194_31493 , \31195_31494 , \31196_31495 ,
         \31197_31496 , \31198_31497 , \31199_31498 , \31200_31499 , \31201_31500 , \31202_31501 , \31203_31502 , \31204_31503 , \31205_31504 , \31206_31505 ,
         \31207_31506 , \31208_31507 , \31209_31508 , \31210_31509 , \31211_31510 , \31212_31511 , \31213_31512 , \31214_31513 , \31215_31514 , \31216_31515 ,
         \31217_31516 , \31218_31517 , \31219_31518 , \31220_31519 , \31221_31520 , \31222_31521 , \31223_31522 , \31224_31523 , \31225_31524 , \31226_31525 ,
         \31227_31526 , \31228_31527 , \31229_31528 , \31230_31529 , \31231_31530 , \31232_31531 , \31233_31532 , \31234_31533 , \31235_31534 , \31236_31535 ,
         \31237_31536 , \31238_31537 , \31239_31538 , \31240_31539 , \31241_31540 , \31242_31541 , \31243_31542 , \31244_31543 , \31245_31544 , \31246_31545 ,
         \31247_31546 , \31248_31547 , \31249_31548 , \31250_31549 , \31251_31550 , \31252_31551 , \31253_31552 , \31254_31553 , \31255_31554 , \31256_31555 ,
         \31257_31556 , \31258_31557 , \31259_31558 , \31260_31559 , \31261_31560 , \31262_31561 , \31263_31562 , \31264_31563 , \31265_31564 , \31266_31565 ,
         \31267_31566 , \31268_31567 , \31269_31568 , \31270_31569 , \31271_31570 , \31272_31571 , \31273_31572 , \31274_31573 , \31275_31574 , \31276_31575 ,
         \31277_31576 , \31278_31577 , \31279_31578 , \31280_31579 , \31281_31580 , \31282_31581 , \31283_31582 , \31284_31583 , \31285_31584 , \31286_31585 ,
         \31287_31586 , \31288_31587 , \31289_31588 , \31290_31589 , \31291_31590 , \31292_31591 , \31293_31592 , \31294_31593 , \31295_31594 , \31296_31595 ,
         \31297_31596 , \31298_31597 , \31299_31598 , \31300_31599 , \31301_31600 , \31302_31601 , \31303_31602 , \31304_31603 , \31305_31604 , \31306_31605 ,
         \31307_31606 , \31308_31607 , \31309_31608 , \31310_31609 , \31311_31610 , \31312_31611 , \31313_31612 , \31314_31613 , \31315_31614 , \31316_31615 ,
         \31317 , \31318_31617 , \31319_31618 , \31320_31619 , \31321_31620 , \31322_31621 , \31323_31622 , \31324_31623 , \31325_31624 , \31326_31625 ,
         \31327_31626 , \31328_31627_nG43fa , \31329_31628 , \31330_31629 , \31331_31630_nG43fd , \31332_31631 , \31333_31632 , \31334_31633 , \31335_31637 , \31336_31638 ,
         \31337_31639 , \31338_31640 , \31339_31641 , \31340_31642 , \31341_31643 , \31342_31644 , \31343_31645 , \31344_31646 , \31345_31647 , \31346_31648 ,
         \31347_31649 , \31348_31650 , \31349_31651 , \31350_31652 , \31351_31653 , \31352_31654 , \31353_31655 , \31354_31656 , \31355_31657 , \31356_31658 ,
         \31357_31659 , \31358_31660 , \31359_31661 , \31360_31662 , \31361_31663 , \31362_31664 , \31363_31665 , \31364_31666 , \31365_31667 , \31366_31668 ,
         \31367_31669 , \31368_31670 , \31369_31671 , \31370_31672 , \31371_31673 , \31372_31674 , \31373_31675 , \31374_31676 , \31375_31677 , \31376_31678 ,
         \31377_31679 , \31378_31680 , \31379_31681 , \31380_31682 , \31381_31683 , \31382_31684 , \31383_31685 , \31384_31686 , \31385_31687 , \31386_31688 ,
         \31387_31689 , \31388_31690 , \31389_31691 , \31390_31692 , \31391_31693 , \31392_31694 , \31393_31695 , \31394_31696 , \31395_31697 , \31396_31698 ,
         \31397_31699 , \31398_31700 , \31399_31701 , \31400_31702 , \31401_31703 , \31402_31704 , \31403_31705 , \31404_31706 , \31405_31707 , \31406_31708 ,
         \31407_31709 , \31408_31710 , \31409_31711 , \31410_31712 , \31411_31713 , \31412_31714 , \31413_31715 , \31414_31716 , \31415_31717 , \31416_31718 ,
         \31417_31719 , \31418_31720 , \31419_31721 , \31420_31722 , \31421_31723 , \31422_31724 , \31423_31725 , \31424_31726 , \31425_31727 , \31426_31728 ,
         \31427_31729 , \31428_31730 , \31429_31731 , \31430_31732 , \31431_31733 , \31432_31734 , \31433_31735 , \31434_31736 , \31435_31737 , \31436_31738 ,
         \31437_31739 , \31438_31740 , \31439_31741 , \31440_31742 , \31441_31743 , \31442_31744 , \31443_31745 , \31444_31746 , \31445_31747 , \31446_31748 ,
         \31447_31749 , \31448_31750 , \31449_31751 , \31450_31752 , \31451_31753 , \31452_31754 , \31453_31755 , \31454_31756 , \31455_31757 , \31456_31758 ,
         \31457_31759 , \31458_31760 , \31459_31761 , \31460_31762 , \31461_31763 , \31462_31764 , \31463_31765 , \31464_31766 , \31465_31767 , \31466_31768 ,
         \31467_31769 , \31468_31770 , \31469_31771 , \31470_31772 , \31471_31773 , \31472_31774 , \31473_31775 , \31474_31776 , \31475_31777 , \31476_31778 ,
         \31477_31779 , \31478_31780 , \31479_31781 , \31480_31782 , \31481_31783 , \31482_31784 , \31483_31785 , \31484_31786 , \31485_31787 , \31486_31788 ,
         \31487_31789 , \31488_31790 , \31489_31791 , \31490_31792 , \31491_31793 , \31492_31794 , \31493_31795 , \31494_31796 , \31495_31797 , \31496_31798 ,
         \31497_31799 , \31498_31800 , \31499_31801 , \31500_31802 , \31501_31803 , \31502_31804 , \31503_31805 , \31504_31806 , \31505_31807 , \31506_31808 ,
         \31507_31809 , \31508_31810 , \31509_31811 , \31510_31812 , \31511_31813 , \31512_31814 , \31513_31815 , \31514_31816 , \31515_31817 , \31516_31818 ,
         \31517_31819 , \31518_31820 , \31519_31821 , \31520_31822 , \31521_31823 , \31522_31824 , \31523_31825 , \31524_31826 , \31525_31827 , \31526_31828 ,
         \31527_31829 , \31528_31830 , \31529_31831 , \31530_31832 , \31531_31833 , \31532_31834 , \31533_31835 , \31534_31836 , \31535_31837 , \31536_31838 ,
         \31537_31839 , \31538_31840 , \31539_31841 , \31540_31842 , \31541_31843 , \31542_31844 , \31543_31845 , \31544_31846 , \31545_31847 , \31546_31848 ,
         \31547_31849 , \31548_31850 , \31549_31851 , \31550_31852 , \31551_31853 , \31552_31854 , \31553_31855 , \31554_31856 , \31555_31857 , \31556_31858 ,
         \31557_31859 , \31558_31860 , \31559_31861 , \31560_31862 , \31561_31863 , \31562_31864 , \31563_31865 , \31564_31866 , \31565_31867 , \31566_31868 ,
         \31567_31869 , \31568_31870 , \31569_31871 , \31570_31872 , \31571_31873 , \31572_31874 , \31573_31875 , \31574_31876 , \31575_31877 , \31576_31878 ,
         \31577_31879 , \31578_31880 , \31579_31881 , \31580_31882 , \31581_31883 , \31582_31884 , \31583_31885 , \31584_31886 , \31585_31887 , \31586_31888 ,
         \31587_31889 , \31588_31890 , \31589_31891 , \31590_31892 , \31591_31893 , \31592_31894 , \31593_31895 , \31594_31896 , \31595_31897 , \31596_31898 ,
         \31597_31899 , \31598_31900 , \31599_31901 , \31600_31902 , \31601_31903 , \31602_31904 , \31603_31905 , \31604_31906 , \31605_31907 , \31606_31908 ,
         \31607_31909 , \31608_31910 , \31609_31911 , \31610_31912 , \31611_31913 , \31612_31914 , \31613_31915 , \31614_31916 , \31615_31917 , \31616_31918 ,
         \31617_31919 , \31618 , \31619_31921 , \31620_31922 , \31621_31923 , \31622_31924 , \31623_31925 , \31624_31926 , \31625_31927 , \31626_31928 ,
         \31627_31929 , \31628_31930 , \31629_31931 , \31630_31932 , \31631_31933 , \31632_31934 , \31633_31935 , \31634_31936 , \31635_31937 , \31636_31938 ,
         \31637_31939 , \31638_31940 , \31639_31941 , \31640_31942 , \31641_31943 , \31642_31944 , \31643_31945 , \31644_31946 , \31645_31947 , \31646_31948 ,
         \31647_31949 , \31648_31950 , \31649_31951 , \31650_31952 , \31651_31953 , \31652_31954 , \31653_31955 , \31654_31956 , \31655_31957 , \31656_31958 ,
         \31657_31959 , \31658_31960 , \31659_31961 , \31660_31962 , \31661_31963 , \31662_31964 , \31663_31965 , \31664_31966 , \31665_31967 , \31666_31968 ,
         \31667_31969 , \31668_31970 , \31669_31971 , \31670_31972 , \31671_31973 , \31672_31974 , \31673_31975 , \31674_31976 , \31675_31977 , \31676_31978 ,
         \31677_31979 , \31678_31980 , \31679_31981 , \31680_31982 , \31681_31983 , \31682_31984 , \31683_31985 , \31684_31986 , \31685_31987 , \31686_31988 ,
         \31687_31989 , \31688_31990 , \31689_31991 , \31690_31992 , \31691_31993 , \31692_31994 , \31693_31995 , \31694_31996 , \31695_31997 , \31696_31998 ,
         \31697_31999 , \31698_32000 , \31699_32001 , \31700_32002 , \31701_32003 , \31702_32004 , \31703_32005 , \31704_32006 , \31705_32007 , \31706_32008 ,
         \31707_32009 , \31708_32010 , \31709_32011 , \31710_32012 , \31711_32013 , \31712_32014 , \31713_32015 , \31714_32016 , \31715_32017 , \31716_32018 ,
         \31717_32019 , \31718_32020 , \31719_32021 , \31720_32022 , \31721_32023 , \31722_32024 , \31723_32025 , \31724_32026 , \31725_32027 , \31726_32028 ,
         \31727_32029 , \31728_32030 , \31729_32031 , \31730_32032 , \31731_32033 , \31732_32034 , \31733_32035 , \31734_32036 , \31735_32037 , \31736_32038 ,
         \31737_32039 , \31738_32040 , \31739_32041 , \31740_32042 , \31741_32043 , \31742_32044 , \31743_32045 , \31744_32046 , \31745_32047 , \31746_32048 ,
         \31747_32049 , \31748_32050 , \31749_32051 , \31750 , \31751_32053_nG65d3 , \31752_32054 , \31753_32055 , \31754_32056 , \31755_32057 , \31756_32058 ,
         \31757_32059 , \31758_32060 , \31759_32061 , \31760_32062 , \31761 , \31762 , \31763_32065_nG646d , \31764_32066 , \31765_32067 , \31766_32068 ,
         \31767_32069 , \31768_32070 , \31769_32071 , \31770_32072 , \31771_32073 , \31772_32074 , \31773_32075 , \31774_32076 , \31775_32077 , \31776_32078 ,
         \31777_32079 , \31778_32080 , \31779_32081 , \31780_32082 , \31781_32083 , \31782_32084 , \31783_32085 , \31784_32086 , \31785_32087 , \31786_32088 ,
         \31787_32089 , \31788_32090 , \31789_32091 , \31790_32092 , \31791_32093 , \31792_32094 , \31793_32095 , \31794_32096 , \31795_32097 , \31796_32098 ,
         \31797_32099 , \31798_32100 , \31799_32101 , \31800_32102 , \31801_32103 , \31802_32104 , \31803_32105 , \31804_32106 , \31805_32107 , \31806_32108 ,
         \31807_32109 , \31808_32110 , \31809_32111 , \31810_32112 , \31811_32113 , \31812_32114 , \31813_32115 , \31814_32116 , \31815_32117 , \31816_32118 ,
         \31817_32119 , \31818_32120 , \31819_32121 , \31820_32122 , \31821_32123 , \31822_32124 , \31823_32125 , \31824_32126 , \31825_32127 , \31826_32128 ,
         \31827_32129 , \31828_32130 , \31829_32131 , \31830_32132 , \31831_32133 , \31832_32134 , \31833_32135 , \31834_32136 , \31835_32137 , \31836_32138 ,
         \31837_32139 , \31838_32140 , \31839_32141 , \31840_32142 , \31841_32143 , \31842_32144 , \31843_32145 , \31844_32146 , \31845_32147 , \31846_32148 ,
         \31847_32149 , \31848_32150 , \31849_32151 , \31850_32152 , \31851_32153 , \31852_32154 , \31853_32155 , \31854_32156 , \31855_32157 , \31856_32158 ,
         \31857_32159 , \31858_32160 , \31859_32161 , \31860_32162 , \31861_32163 , \31862_32164 , \31863_32165 , \31864_32166 , \31865_32167 , \31866_32168 ,
         \31867_32169 , \31868_32170 , \31869_32171 , \31870_32172 , \31871_32173 , \31872_32174 , \31873_32175 , \31874_32176 , \31875_32177 , \31876_32178 ,
         \31877_32179_nG9bb4 , \31878_32180 , \31879_32181 , \31880_32182 , \31881_32183 , \31882_32184 , \31883_32185 , \31884_32186 , \31885_32187 , \31886_32188 ,
         \31887_32189 , \31888_32190 , \31889_32191 , \31890_32192 , \31891_32193 , \31892_32194 , \31893_32195 , \31894_32196 , \31895_32197 , \31896_32198 ,
         \31897_32199 , \31898_32200 , \31899_32201 , \31900_32202 , \31901_32203 , \31902_32204 , \31903_32205 , \31904_32206 , \31905_32207 , \31906_32208 ,
         \31907_32209 , \31908_32210 , \31909_32211 , \31910_32212 , \31911_32213 , \31912_32214 , \31913_32215 , \31914_32216 , \31915_32217 , \31916_32218 ,
         \31917_32219 , \31918_32220 , \31919_32221 , \31920_32222 , \31921_32223 , \31922_32224 , \31923_32225 , \31924_32226 , \31925_32227 , \31926_32228 ,
         \31927_32229 , \31928_32230 , \31929_32231 , \31930_32232 , \31931_32233 , \31932_32234 , \31933_32235 , \31934_32236 , \31935_32237 , \31936_32238 ,
         \31937_32239 , \31938_32240 , \31939_32241 , \31940_32242 , \31941_32243 , \31942_32244 , \31943_32245 , \31944_32246 , \31945_32247 , \31946_32248 ,
         \31947_32249 , \31948_32250 , \31949_32251 , \31950_32252 , \31951_32253 , \31952_32254 , \31953_32255 , \31954_32256 , \31955_32257 , \31956_32258 ,
         \31957_32259 , \31958_32260 , \31959_32261 , \31960_32262 , \31961_32263 , \31962_32264 , \31963_32265 , \31964_32266 , \31965_32267 , \31966_32268 ,
         \31967_32269 , \31968_32270 , \31969_32271 , \31970_32272 , \31971_32273 , \31972_32274 , \31973_32275 , \31974_32276 , \31975_32277 , \31976_32278 ,
         \31977_32279 , \31978_32280 , \31979_32281 , \31980_32282 , \31981_32283 , \31982_32284 , \31983_32285 , \31984_32286 , \31985_32287 , \31986_32288 ,
         \31987_31634 , \31988_31635 , \31989_31636 , \31990_32289 , \31991_32290 , \31992_32291 , \31993_32292 , \31994_32293 , \31995_32294 , \31996_32295 ,
         \31997_32296 , \31998_32297 , \31999_32298 , \32000_32299 , \32001_32300 , \32002_32301 , \32003_32302 , \32004_32303 , \32005_32304 , \32006_32305 ,
         \32007_32306 , \32008_32307 , \32009_32308 , \32010_32309 , \32011_32310 , \32012_32311 , \32013_32312 , \32014_32313 , \32015_32314 , \32016_32315 ,
         \32017_32316 , \32018_32317 , \32019_32318 , \32020_32319 , \32021_32320 , \32022_32321 , \32023_32322 , \32024_32323 , \32025_32324 , \32026_32325 ,
         \32027_32326 , \32028_32327 , \32029_32328 , \32030_32329 , \32031_32330 , \32032_32331 , \32033_32332 , \32034_32333 , \32035_32334 , \32036_32335 ,
         \32037_32336 , \32038_32337 , \32039_32338 , \32040_32339 , \32041_32340 , \32042_32341 , \32043_32342 , \32044_32343 , \32045_32344 , \32046_32345 ,
         \32047_32346 , \32048_32347 , \32049_32348 , \32050_32349 , \32051_32350 , \32052_32351 , \32053_32352 , \32054_32353 , \32055_32354 , \32056_32355 ,
         \32057_32356 , \32058_32357 , \32059_32358 , \32060_32359 , \32061_32360 , \32062_32361 , \32063_32362 , \32064_32363 , \32065_32364 , \32066_32365 ,
         \32067_32366 , \32068_32367 , \32069_32368 , \32070_32369 , \32071_32370 , \32072_32371 , \32073_32372 , \32074_32373 , \32075_32374 , \32076_32375 ,
         \32077_32376 , \32078_32377 , \32079_32378 , \32080_32379 , \32081_32380 , \32082_32381 , \32083_32382 , \32084_32383 , \32085_32384 , \32086_32385 ,
         \32087_32386 , \32088_32387 , \32089_32388 , \32090_32389 , \32091_32390 , \32092_32391 , \32093_32392 , \32094_32393 , \32095_32394 , \32096_32395 ,
         \32097_32396 , \32098_32397 , \32099_32398 , \32100_32399 , \32101_32400 , \32102_32401 , \32103_32402 , \32104_32403 , \32105_32404 , \32106_32405 ,
         \32107_32406 , \32108_32407 , \32109_32408 , \32110_32409 , \32111_32410 , \32112_32411 , \32113_32412 , \32114_32413 , \32115_32414 , \32116_32415 ,
         \32117_32416 , \32118_32417 , \32119_32418 , \32120_32419 , \32121_32420 , \32122_32421 , \32123_32422 , \32124_32423 , \32125_32424 , \32126_32425 ,
         \32127_32426 , \32128_32427 , \32129_32428 , \32130_32429 , \32131_32430 , \32132_32431 , \32133_32432 , \32134_32433 , \32135_32434 , \32136_32435 ,
         \32137_32436 , \32138_32437 , \32139_32438 , \32140_32439 , \32141_32440 , \32142_32441 , \32143_32442 , \32144_32443 , \32145_32444 , \32146_32445 ,
         \32147_32446 , \32148_32447 , \32149_32448 , \32150_32449 , \32151_32450 , \32152_32451 , \32153_32452 , \32154_32453 , \32155_32454 , \32156_32455 ,
         \32157_32456 , \32158_32457 , \32159_32458 , \32160_32459 , \32161_32460 , \32162_32461 , \32163_32462 , \32164_32463 , \32165_32464 , \32166_32465 ,
         \32167_32466 , \32168_32467 , \32169_32468 , \32170_32469 , \32171_32470 , \32172_32471 , \32173_32472 , \32174_32473 , \32175_32474 , \32176_32475 ,
         \32177_32476 , \32178_32477 , \32179_32478 , \32180_32479 , \32181_32480 , \32182_32481 , \32183_32482 , \32184_32483 , \32185_32484 , \32186_32485 ,
         \32187_32486 , \32188_32487 , \32189_32488 , \32190_32489 , \32191_32490 , \32192_32491 , \32193_32492 , \32194_32493 , \32195_32494 , \32196_32495 ,
         \32197_32496 , \32198_32497 , \32199_32498 , \32200_32499 , \32201_32500 , \32202_32501 , \32203_32502 , \32204_32503 , \32205_32504 , \32206_32505 ,
         \32207_32506 , \32208_32507 , \32209_32508 , \32210_32509 , \32211_32510 , \32212_32511 , \32213_32512 , \32214_32513 , \32215_32514 , \32216_32515 ,
         \32217_32516 , \32218_32517 , \32219_32518 , \32220_32519 , \32221_32520 , \32222_32521 , \32223_32522 , \32224_32523 , \32225_32524 , \32226_32525 ,
         \32227_32526 , \32228_32527 , \32229_32528 , \32230_32529 , \32231_32530 , \32232_32531 , \32233_32532 , \32234_32533 , \32235_32534 , \32236_32535 ,
         \32237_32536 , \32238_32537 , \32239_32538 , \32240_32539 , \32241_32540 , \32242_32541 , \32243_32542 , \32244_32543 , \32245_32544 , \32246_32545 ,
         \32247_32546 , \32248_32547 , \32249_32548 , \32250_32549 , \32251_32550 , \32252_32551 , \32253_32552 , \32254_32553 , \32255_32554 , \32256_32555 ,
         \32257_32556 , \32258_32557 , \32259_32558 , \32260_32559 , \32261_32560 , \32262_32561 , \32263_32562 , \32264_32563 , \32265_32564 , \32266_32565 ,
         \32267_32566 , \32268_32567 , \32269_32568 , \32270_32569 , \32271_32570 , \32272_32571 , \32273_32572 , \32274_32573 , \32275_32574 , \32276_32575 ,
         \32277_32576 , \32278_32577 , \32279_32578 , \32280_32579 , \32281_32580 , \32282_32581 , \32283_32582 , \32284_32583 , \32285_32584 , \32286_32585 ,
         \32287_32586 , \32288_32587 , \32289_32588 , \32290_32589 , \32291_32590 , \32292_32591 , \32293_32592 , \32294_32593 , \32295_32594 , \32296_32595 ,
         \32297_32596 , \32298_32597 , \32299_32598 , \32300_32599 , \32301_32600 , \32302_32601 , \32303_32602 , \32304_32603 , \32305_32604 , \32306_32605 ,
         \32307_32606 , \32308_32607 , \32309_32608 , \32310_32609 , \32311_32610 , \32312_32611 , \32313_32612 , \32314_32613 , \32315_32614 , \32316_32615 ,
         \32317_32616 , \32318_32617 , \32319_32618 , \32320_32619 , \32321_32620 , \32322_32621 , \32323_32622 , \32324_32623 , \32325_32624 , \32326_32625 ,
         \32327_32626 , \32328_32627 , \32329_32628 , \32330_32629 , \32331_32630 , \32332_32631 , \32333_32632 , \32334_32633 , \32335_32634 , \32336_32635 ,
         \32337_32636 , \32338_32637 , \32339_32638 , \32340_32639 , \32341_32640 , \32342_32641 , \32343_32642 , \32344_32643 , \32345_32644 , \32346_32645 ,
         \32347_32646 , \32348_32647 , \32349_32648 , \32350_32649 , \32351_32650 , \32352_32651 , \32353_32652 , \32354_32653 , \32355_32654 , \32356_32655 ,
         \32357_32656 , \32358_32657 , \32359_32658 , \32360_32659 , \32361 , \32362_32661 , \32363_32662 , \32364_32663 , \32365_32664 , \32366_32665 ,
         \32367_32666 , \32368_32667 , \32369_32668 , \32370_32669 , \32371_32670 , \32372_32671 , \32373_32672 , \32374_32673 , \32375_32674 , \32376_32675 ,
         \32377_32676 , \32378_32677 , \32379_32678 , \32380_32679 , \32381_32680 , \32382_32681 , \32383_32682 , \32384_32683 , \32385_32684 , \32386_32685 ,
         \32387_32686 , \32388_32687 , \32389_32688 , \32390_32689 , \32391_32690 , \32392_32691 , \32393_32692 , \32394_32693 , \32395_32694 , \32396_32695 ,
         \32397_32696 , \32398_32697 , \32399_32698 , \32400_32699 , \32401_32700 , \32402_32701 , \32403_32702 , \32404_32703 , \32405_32704 , \32406_32705 ,
         \32407_32706 , \32408_32707 , \32409_32708 , \32410_32709 , \32411_32710 , \32412_32711 , \32413_32712 , \32414_32713 , \32415_32714 , \32416_32715 ,
         \32417_32716 , \32418_32717 , \32419_32718 , \32420_32719 , \32421_32720 , \32422_32721 , \32423_32722 , \32424_32723 , \32425_32724 , \32426_32725 ,
         \32427_32726 , \32428_32727 , \32429_32728 , \32430_32729 , \32431_32730 , \32432_32731 , \32433_32732 , \32434_32733 , \32435_32734 , \32436_32735 ,
         \32437_32736 , \32438_32737 , \32439_32738 , \32440_32739 , \32441_32740 , \32442_32741 , \32443_32742 , \32444_32743 , \32445_32744 , \32446_32745 ,
         \32447_32746 , \32448_32747 , \32449_32748 , \32450_32749 , \32451_32750 , \32452_32751 , \32453_32752 , \32454_32753 , \32455_32754 , \32456_32755 ,
         \32457_32756 , \32458_32757 , \32459_32758 , \32460_32759 , \32461_32760 , \32462_32761 , \32463_32762 , \32464_32763 , \32465_32764 , \32466_32765 ,
         \32467_32766 , \32468_32767 , \32469_32768 , \32470_32769 , \32471_32770 , \32472_32771 , \32473_32772 , \32474_32773 , \32475_32774 , \32476_32775 ,
         \32477_32776 , \32478_32777 , \32479_32778 , \32480_32779 , \32481_32780 , \32482_32781 , \32483_32782 , \32484_32783 , \32485_32784 , \32486_32785 ,
         \32487_32786 , \32488_32787 , \32489_32788 , \32490_32789 , \32491_32790 , \32492_32791 , \32493 , \32494_32793_nG65d6 , \32495_32794 , \32496_32795 ,
         \32497_32796 , \32498_32797 , \32499_32798 , \32500 , \32501 , \32502_32801_nG6576 , \32503_32802 , \32504_32803 , \32505_32804 , \32506_32805 ,
         \32507_32806 , \32508_32807 , \32509_32808 , \32510_32809 , \32511_32810 , \32512_32811 , \32513_32812 , \32514_32813 , \32515_32814 , \32516_32815 ,
         \32517_32816 , \32518_32817 , \32519_32818 , \32520_32819 , \32521_32820 , \32522_32821 , \32523_32822 , \32524_32823 , \32525_32824 , \32526_32825 ,
         \32527_32826 , \32528_32827 , \32529_32828 , \32530_32829 , \32531_32830 , \32532_32831 , \32533_32832 , \32534_32833 , \32535_32834 , \32536_32835 ,
         \32537_32836 , \32538_32837 , \32539_32838 , \32540_32839 , \32541_32840 , \32542_32841 , \32543_32842 , \32544_32843 , \32545_32844 , \32546_32845 ,
         \32547_32846 , \32548_32847 , \32549_32848 , \32550_32849 , \32551_32850 , \32552_32851 , \32553_32852 , \32554_32853 , \32555_32854 , \32556_32855 ,
         \32557_32856 , \32558_32857 , \32559_32858 , \32560_32859 , \32561_32860 , \32562_32861 , \32563_32862 , \32564_32863 , \32565_32864 , \32566_32865 ,
         \32567_32866 , \32568_32867 , \32569_32868 , \32570_32869 , \32571_32870 , \32572_32871 , \32573_32872 , \32574_32873 , \32575_32874 , \32576_32875 ,
         \32577_32876 , \32578_32877 , \32579_32878 , \32580_32879 , \32581_32880 , \32582_32881 , \32583_32882 , \32584_32883 , \32585_32884 , \32586_32885 ,
         \32587_32886 , \32588_32887 , \32589_32888_nG9bb1 , \32590_32889 , \32591_32890 , \32592_32891 , \32593_32892 , \32594_32893 , \32595_32894 , \32596_32895 ,
         \32597_32896 , \32598_32897 , \32599_32898 , \32600_32899 , \32601_32900 , \32602_32901 , \32603_32902 , \32604_32903 , \32605_32904 , \32606_32905 ,
         \32607_32906 , \32608_32907 , \32609_32908 , \32610_32909 , \32611_32910 , \32612_32911 , \32613_32912 , \32614_32913 , \32615_32914 , \32616_32915 ,
         \32617_32916 , \32618_32918 , \32619_32919 , \32620_32920 , \32621_32921 , \32622_32922 , \32623_32923 , \32624_32924 , \32625_32925 , \32626_32926 ,
         \32627_32927 , \32628_32928 , \32629_32929 , \32630_32930 , \32631_32931 , \32632_32932 , \32633_32933 , \32634_32934 , \32635_32935 , \32636_32936 ,
         \32637_32937 , \32638_32938 , \32639_32939 , \32640_32940 , \32641_32941 , \32642_32942 , \32643_32943 , \32644_32944 , \32645_32945 , \32646_32946 ,
         \32647_32947 , \32648_32948 , \32649_32949 , \32650_32950 , \32651_32951 , \32652_32952 , \32653_32953 , \32654_32954 , \32655_32955 , \32656_32956 ,
         \32657_32957 , \32658_32958 , \32659_32959 , \32660_32960 , \32661_32961 , \32662_32962 , \32663_32963 , \32664_32964 , \32665_32965 , \32666_32966 ,
         \32667_32967 , \32668_32968 , \32669_32969 , \32670_32970 , \32671_32971 , \32672_32972 , \32673_32973 , \32674_32974 , \32675_32975 , \32676_32976 ,
         \32677_32977 , \32678_32978 , \32679_32979 , \32680_32980 , \32681_32981 , \32682_32982 , \32683_32983 , \32684_32984 , \32685_32985 , \32686_32986 ,
         \32687_32987 , \32688_32988 , \32689_32989 , \32690_32990 , \32691_32991 , \32692_32992 , \32693_32993 , \32694_32994 , \32695_32995 , \32696_32996 ,
         \32697_32997 , \32698_32998 , \32699_32999 , \32700_33000 , \32701_33001 , \32702_33002 , \32703_33003 , \32704_33004 , \32705_33005 , \32706_33006 ,
         \32707_33007 , \32708_33008 , \32709_33009 , \32710_33010 , \32711_33011 , \32712_33012 , \32713_33013 , \32714_33014 , \32715_33015 , \32716_33016 ,
         \32717_33017 , \32718_33018 , \32719_33019 , \32720_33020 , \32721_33021 , \32722_33022 , \32723_33023 , \32724_33024 , \32725_33025 , \32726_33026 ,
         \32727_33027 , \32728_33028 , \32729_33029 , \32730_33030 , \32731_33031 , \32732_33032 , \32733_33033 , \32734_33034 , \32735_33035 , \32736_33036 ,
         \32737_33037 , \32738_33038 , \32739_33039 , \32740_33040 , \32741_33041 , \32742_33042 , \32743_33043 , \32744_33044 , \32745_33045 , \32746_33046 ,
         \32747_33047 , \32748_33048 , \32749_33049 , \32750_33050 , \32751_33051 , \32752_33052 , \32753_33053 , \32754_33054 , \32755_33055 , \32756_33056 ,
         \32757_33057 , \32758_33058 , \32759_33059 , \32760_33060 , \32761_33061 , \32762_33062 , \32763_33063 , \32764_33064 , \32765_33065 , \32766_33066 ,
         \32767_33067 , \32768_33068 , \32769_33069 , \32770_33070 , \32771_33071 , \32772_33072 , \32773_33073 , \32774_33074 , \32775_33075 , \32776_33076 ,
         \32777_33077 , \32778_33078 , \32779_33079 , \32780_33080 , \32781_33081 , \32782_33082 , \32783_33083 , \32784_33084 , \32785_33085 , \32786_33086 ,
         \32787_33087 , \32788_33088 , \32789_33089 , \32790_33090 , \32791_33091 , \32792_33092 , \32793_33093 , \32794_33094 , \32795_33095 , \32796_33096 ,
         \32797_33097 , \32798_33098 , \32799_33099 , \32800_33100 , \32801_33101 , \32802_33102 , \32803_33103 , \32804_33104 , \32805_33105 , \32806_33106 ,
         \32807_33107 , \32808_33108 , \32809_33109 , \32810_33110 , \32811_33111 , \32812_33112 , \32813_33113 , \32814_33114 , \32815_33115 , \32816_33116 ,
         \32817_33117 , \32818_33118 , \32819_33119 , \32820_33120 , \32821_33121 , \32822_33122 , \32823_33123 , \32824_33124 , \32825_33125 , \32826_33126 ,
         \32827_33127 , \32828_33128 , \32829_33129 , \32830_33130 , \32831_33131 , \32832_33132 , \32833_33133 , \32834_33134 , \32835_33135 , \32836_33136 ,
         \32837_33137 , \32838_33138 , \32839_33139 , \32840_33140 , \32841_33141 , \32842_33142 , \32843_33143 , \32844_33144 , \32845_33145 , \32846_33146 ,
         \32847_33147 , \32848_33148 , \32849_33149 , \32850_33150 , \32851_33151 , \32852_33152 , \32853_33153 , \32854_33154 , \32855_33155 , \32856_33156 ,
         \32857_33157 , \32858_33158 , \32859_33159 , \32860_33160 , \32861_33161 , \32862_33162 , \32863_33163 , \32864_33164 , \32865_33165 , \32866_33166 ,
         \32867_33167 , \32868_33168 , \32869_33169 , \32870_33170 , \32871_33171 , \32872_33172 , \32873_33173 , \32874_33174 , \32875_33175 , \32876_33176 ,
         \32877_33177 , \32878_33178 , \32879_33179 , \32880_33180 , \32881_33181_nG9bae , \32882_33182 , \32883_33183 , \32884_33184 , \32885_33185 , \32886_33186 ,
         \32887_33187 , \32888_33188 , \32889_33189 , \32890_33190 , \32891_33191 , \32892_33192 , \32893_33193 , \32894_33194 , \32895_33195 , \32896_33196 ,
         \32897_33197 , \32898_33198 , \32899_33199 , \32900_33200 , \32901_33201 , \32902_33202 , \32903_33203 , \32904_33204 , \32905_33205 , \32906_33206 ,
         \32907_33207 , \32908_33208 , \32909_33209 , \32910_33210 , \32911_33211 , \32912_33212 , \32913_33213 , \32914_33214 , \32915_33215 , \32916_33216 ,
         \32917_33217 , \32918_33218 , \32919_33219 , \32920_33220 , \32921_33221 , \32922_33222 , \32923_33223 , \32924_33224 , \32925_33225 , \32926_33226 ,
         \32927_33227 , \32928_33228 , \32929_33229 , \32930_33230 , \32931_33231 , \32932_33232 , \32933_33233 , \32934_33234 , \32935_33235 , \32936_33236 ,
         \32937_33237 , \32938_33238 , \32939_33239 , \32940_33240 , \32941_33241 , \32942_33242 , \32943_33243 , \32944_33244 , \32945_33245 , \32946_33246 ,
         \32947_33247 , \32948_33248 , \32949_33249 , \32950_33250 , \32951_33251 , \32952_33252 , \32953_33253 , \32954_33254 , \32955_33255 , \32956_33256 ,
         \32957_33257 , \32958_33258 , \32959_33259 , \32960_33260 , \32961_33261 , \32962_33262 , \32963_33263 , \32964_33264 , \32965_33265 , \32966_33266 ,
         \32967_33267 , \32968_33268 , \32969_33269 , \32970_33270 , \32971_33271 , \32972_33272 , \32973_33273 , \32974_33274 , \32975_33275 , \32976_33276 ,
         \32977_33277 , \32978_33278 , \32979_33279 , \32980_33280 , \32981_33281 , \32982_33282 , \32983_33283 , \32984_33284 , \32985_33285 , \32986_33286 ,
         \32987_33287 , \32988_33288 , \32989_33289 , \32990_33290 , \32991_33291 , \32992_33292 , \32993_33293 , \32994_33294 , \32995_33295 , \32996_33296 ,
         \32997_33297 , \32998_33298 , \32999_33299 , \33000_33300 , \33001_33301 , \33002_33302 , \33003_33303 , \33004_33304 , \33005_33305 , \33006_33306 ,
         \33007_33307 , \33008_33308 , \33009_33309 , \33010_33310 , \33011_33311 , \33012_33312 , \33013_33313 , \33014_33314 , \33015_33315 , \33016_33316 ,
         \33017_33317 , \33018_33318 , \33019_33319 , \33020_33320 , \33021_33321 , \33022_33322 , \33023_33323 , \33024_33324 , \33025_33325 , \33026_33326 ,
         \33027_33327 , \33028_33328 , \33029_33329 , \33030_33330 , \33031_33331 , \33032_33332 , \33033_33333 , \33034_33334 , \33035_33335 , \33036_33336 ,
         \33037_33337 , \33038_33338 , \33039_33339 , \33040_33340 , \33041_33341 , \33042_33342 , \33043_33343 , \33044_33344 , \33045_33345 , \33046_33346 ,
         \33047_33347 , \33048_33348 , \33049_33349 , \33050_33350 , \33051_33351 , \33052_33352 , \33053_33353 , \33054_33354 , \33055_33355 , \33056_33356 ,
         \33057_33357 , \33058_33358 , \33059_33359 , \33060_33360 , \33061_33361 , \33062_33362 , \33063_33363 , \33064_33364 , \33065_33365 , \33066_33366 ,
         \33067_33367 , \33068_33368 , \33069_33369 , \33070_33370 , \33071_33371 , \33072_33372 , \33073_33373 , \33074_33374 , \33075_33375 , \33076_33376 ,
         \33077_33377 , \33078_33378 , \33079_33379 , \33080_33380 , \33081_33381 , \33082_33382 , \33083_33383 , \33084_33384 , \33085_33385 , \33086_33386 ,
         \33087_33387 , \33088_33388 , \33089_33389 , \33090_33390 , \33091_33391 , \33092_33392 , \33093_33393 , \33094_33394 , \33095_33395 , \33096_33396 ,
         \33097_33397 , \33098_33398 , \33099_33399 , \33100_33400 , \33101_33401 , \33102_33402 , \33103_33403 , \33104_33404 , \33105_33405 , \33106_33406 ,
         \33107_33407 , \33108_33408 , \33109_33409 , \33110_33410 , \33111_33411 , \33112_33412 , \33113_33413 , \33114_33414 , \33115_33415 , \33116_33416 ,
         \33117_33417 , \33118_33418 , \33119_33419 , \33120_33420 , \33121_33421 , \33122_33422 , \33123_33423 , \33124_33424 , \33125_33425 , \33126_33426 ,
         \33127_33427 , \33128_33428 , \33129_33429 , \33130_33430 , \33131_33431 , \33132_33432 , \33133_33433 , \33134_33434 , \33135_33435 , \33136_33436 ,
         \33137_33437 , \33138_33438 , \33139_33439 , \33140_33440 , \33141_33441 , \33142_33442 , \33143_33443 , \33144_33444 , \33145_33445 , \33146_33446 ,
         \33147_33447 , \33148_33448 , \33149_33449 , \33150_33450 , \33151_33451 , \33152_33452 , \33153_33453 , \33154_33454 , \33155_33455 , \33156_33456 ,
         \33157_33457 , \33158_33458 , \33159_33459 , \33160_33460 , \33161_33461 , \33162_33462 , \33163_33463 , \33164_33464 , \33165_33465 , \33166_33466 ,
         \33167_33467 , \33168_33468 , \33169_33469 , \33170_33470 , \33171_33471 , \33172_33472 , \33173_33473 , \33174_33474 , \33175_33475 , \33176_33476 ,
         \33177_33477 , \33178_33478 , \33179_33479 , \33180_33480 , \33181_33481 , \33182_33482 , \33183_33483 , \33184_33484 , \33185_33485 , \33186_33486 ,
         \33187_33487 , \33188_33488 , \33189_33489 , \33190_33490 , \33191_33491 , \33192_33492 , \33193_33493 , \33194_33494 , \33195_33495 , \33196_33496 ,
         \33197_33497 , \33198_33498 , \33199_33499 , \33200_33500 , \33201_33501 , \33202_33502 , \33203_33503 , \33204_33504 , \33205_33505 , \33206_33506 ,
         \33207_33507 , \33208_33508 , \33209_33509 , \33210_33510 , \33211_33511 , \33212_33512 , \33213_33513 , \33214_33514 , \33215_33515 , \33216_33516 ,
         \33217_33517 , \33218_33518 , \33219_33519 , \33220_33520 , \33221_33521 , \33222_33522 , \33223_33523 , \33224_33524 , \33225_33525 , \33226_33526 ,
         \33227_33527 , \33228_33528 , \33229_33529 , \33230_33530 , \33231_33531 , \33232_33532 , \33233_33533 , \33234_33534 , \33235_33535 , \33236_33536 ,
         \33237_33537 , \33238_33538 , \33239_33539 , \33240_33540 , \33241_33541 , \33242_33542 , \33243_33543 , \33244_33544 , \33245_33545 , \33246_33546 ,
         \33247_33547 , \33248_33548 , \33249_33549 , \33250_33550 , \33251_33551 , \33252_33552 , \33253_33553 , \33254_33554 , \33255_33555 , \33256_33556 ,
         \33257_33557 , \33258_33558 , \33259_33559 , \33260_33560 , \33261_33561 , \33262_33562 , \33263_33563 , \33264_33564 , \33265_33565 , \33266_33566 ,
         \33267_33567 , \33268_33568 , \33269_33569 , \33270_33570 , \33271_33571 , \33272_33572 , \33273_33573 , \33274_33574 , \33275_33575 , \33276_33576 ,
         \33277_33577 , \33278_33578 , \33279_33579 , \33280_33580 , \33281_33581 , \33282_33582 , \33283_33583 , \33284_33584 , \33285_33585 , \33286_33586 ,
         \33287_33587 , \33288_33588 , \33289_33589 , \33290_33590 , \33291_33591 , \33292_33592 , \33293_33593 , \33294_33594 , \33295_33595 , \33296_33596 ,
         \33297_33597 , \33298_33598 , \33299_33599 , \33300_33600 , \33301_33601 , \33302_33602 , \33303_33603 , \33304_33604 , \33305_33605 , \33306_33606 ,
         \33307_33607 , \33308_33608 , \33309_33609 , \33310_33610 , \33311_33611 , \33312_33612 , \33313_33613_nG9bab , \33314_33614 , \33315_33615 , \33316_33616 ,
         \33317_33617 , \33318_33618 , \33319_33619 , \33320_33620 , \33321_33621 , \33322_33622 , \33323_33623 , \33324_33624 , \33325_33625 , \33326_33626 ,
         \33327_33627 , \33328_33628 , \33329_33629 , \33330_33630 , \33331_33631 , \33332_33632 , \33333_33633 , \33334_33634 , \33335_33635 , \33336_33636 ,
         \33337_33637 , \33338_33638 , \33339_33639 , \33340_33640 , \33341_33641 , \33342_33642 , \33343_33643 , \33344_33644 , \33345_33645 , \33346_33646 ,
         \33347_33647 , \33348_33648 , \33349_33649 , \33350_33650 , \33351_33651 , \33352_33652 , \33353_33653 , \33354_33654 , \33355_33655 , \33356_33656 ,
         \33357_33657 , \33358_33658 , \33359_33659 , \33360_33660 , \33361_33661 , \33362_33662 , \33363_33663 , \33364_33664 , \33365_33665 , \33366_33666 ,
         \33367_33667 , \33368_33668 , \33369_33669 , \33370_33670 , \33371_33671 , \33372_33672 , \33373_33673 , \33374_33674 , \33375_33675 , \33376_33676 ,
         \33377_33677 , \33378_33678 , \33379_33679 , \33380_33680 , \33381_33681 , \33382_33682 , \33383_33683 , \33384_33684 , \33385_33685 , \33386_33686 ,
         \33387_33687 , \33388_33688 , \33389_33689 , \33390_33690 , \33391_33691 , \33392_33692 , \33393_33693 , \33394_33694 , \33395_33695 , \33396_33696 ,
         \33397_33697 , \33398_33698 , \33399_33699 , \33400_33700 , \33401_33701 , \33402_33702 , \33403_33703 , \33404_33704 , \33405_33705 , \33406_33706 ,
         \33407_33707 , \33408_33708 , \33409_33709 , \33410_33710 , \33411_33711 , \33412_33712 , \33413_33713 , \33414_33714 , \33415_33715 , \33416_33716 ,
         \33417_33717 , \33418_33718 , \33419_33719 , \33420_33720 , \33421_33721 , \33422_33722 , \33423_33723 , \33424_33724 , \33425_33725 , \33426_33726 ,
         \33427_33727 , \33428_33728 , \33429_33729 , \33430_33730 , \33431_33731 , \33432_33732 , \33433_33733 , \33434_33734 , \33435_33735 , \33436_33736 ,
         \33437_33737 , \33438_33738 , \33439_33739 , \33440_33740 , \33441_33741 , \33442_33742 , \33443_33743 , \33444_33744 , \33445_33745 , \33446_33746 ,
         \33447_33747 , \33448_33748 , \33449_33749 , \33450_33750 , \33451_33751 , \33452_33752 , \33453_33753 , \33454_33754 , \33455_33755 , \33456_33756 ,
         \33457_33757 , \33458_33758 , \33459_33759 , \33460_33760 , \33461_33761 , \33462_33762 , \33463_33763 , \33464_33764 , \33465_33765 , \33466_33766 ,
         \33467_33767 , \33468_33768 , \33469_33769 , \33470_33770 , \33471_33771 , \33472_33772 , \33473_33773 , \33474_33774 , \33475_33775 , \33476_33776 ,
         \33477_33777 , \33478_33778 , \33479_33779 , \33480_33780 , \33481_33781 , \33482_33782 , \33483_33783 , \33484_33784 , \33485_33785 , \33486_33786 ,
         \33487_33787 , \33488_33788 , \33489_33789 , \33490_33790 , \33491_33791 , \33492_33792 , \33493_33793 , \33494_33794 , \33495_33795 , \33496_33796 ,
         \33497_33797 , \33498_33798 , \33499_33799 , \33500_33800 , \33501_33801 , \33502_33802 , \33503_33803 , \33504_33804 , \33505_33805 , \33506_33806 ,
         \33507_33807 , \33508_33808 , \33509_33809 , \33510_33810 , \33511_33811 , \33512_33812 , \33513_33813 , \33514_33814 , \33515_33815 , \33516_33816 ,
         \33517_33817 , \33518_33818 , \33519_33819 , \33520_33820 , \33521_33821 , \33522_33822 , \33523_33823 , \33524_33824 , \33525_33825 , \33526_33826 ,
         \33527_33827 , \33528_33828 , \33529_33829 , \33530_33830 , \33531_33831 , \33532_33832 , \33533_33833 , \33534_33834 , \33535_33835 , \33536_33836 ,
         \33537_33837 , \33538_33838 , \33539_33839 , \33540_33840 , \33541_33841 , \33542_33842 , \33543_33843 , \33544_33844 , \33545_33845 , \33546_33846 ,
         \33547_33847 , \33548_33848 , \33549_33849 , \33550_33850 , \33551_33851 , \33552_33852 , \33553_33853 , \33554_33854 , \33555_33855 , \33556_33856 ,
         \33557_33857 , \33558_33858 , \33559_33859 , \33560_33860 , \33561_33861 , \33562_33862 , \33563_33863 , \33564_33864 , \33565_33865 , \33566_33866 ,
         \33567_33867 , \33568_33868 , \33569_33869 , \33570_33870 , \33571_33871 , \33572_33872 , \33573_33873 , \33574_33874 , \33575_33875 , \33576_33876 ,
         \33577_33877 , \33578_33878 , \33579_33879 , \33580_33880 , \33581_33881 , \33582_33882 , \33583_33883 , \33584_33884 , \33585_33885 , \33586_33886 ,
         \33587_33887 , \33588_33888 , \33589_33889 , \33590_33890 , \33591_33891 , \33592_33892 , \33593_33893 , \33594_33894 , \33595_33895 , \33596_33896 ,
         \33597_33897 , \33598_33898 , \33599_33899 , \33600_33900 , \33601_33901 , \33602_33902 , \33603_33903 , \33604_33904 , \33605_33905 , \33606_33906 ,
         \33607_33907 , \33608_33908 , \33609_33909 , \33610_33910 , \33611_33911 , \33612_33912 , \33613_33913 , \33614_33914 , \33615_33915 , \33616_33916 ,
         \33617_33917 , \33618_33918 , \33619_33919 , \33620_33920 , \33621_33921 , \33622_33922 , \33623_33923 , \33624_33924 , \33625_33925 , \33626_33926 ,
         \33627_33927 , \33628_33928 , \33629_33929 , \33630_33930 , \33631_33931 , \33632_33932 , \33633_33933 , \33634_33934 , \33635_33935 , \33636_33936 ,
         \33637_33937 , \33638_33938 , \33639_33939 , \33640_33940 , \33641_33941 , \33642_33942 , \33643_33943 , \33644_33944 , \33645_33945 , \33646_33946 ,
         \33647_33947 , \33648_33948 , \33649_33949 , \33650_33950 , \33651_33951 , \33652_33952 , \33653_33953 , \33654_33954 , \33655_33955 , \33656_33956 ,
         \33657_33957 , \33658_33958 , \33659_33959 , \33660_33960 , \33661_33961 , \33662_33962 , \33663_33963 , \33664_33964 , \33665_33965 , \33666_33966 ,
         \33667_33967 , \33668_33968 , \33669_33969 , \33670_33970 , \33671_33971 , \33672_33972 , \33673_33973 , \33674_33974 , \33675_33975 , \33676_33976 ,
         \33677_33977 , \33678_33978 , \33679_33979 , \33680_33980 , \33681_33981 , \33682_33982 , \33683_33983 , \33684_33984 , \33685_33985 , \33686_33986 ,
         \33687_33987 , \33688_33988 , \33689_33989 , \33690_33990 , \33691_33991 , \33692_33992 , \33693_33993 , \33694_33994 , \33695_33995 , \33696_33996 ,
         \33697_33997 , \33698_33998 , \33699_33999 , \33700_34000 , \33701_34001 , \33702_34002 , \33703_34003 , \33704_34004 , \33705_34005 , \33706_34006 ,
         \33707_34007 , \33708_34008 , \33709_34009 , \33710_34010 , \33711_34011 , \33712_34012 , \33713_34013 , \33714_34014 , \33715_34015 , \33716_34016 ,
         \33717_34017 , \33718_34018 , \33719_34019 , \33720_34020 , \33721_34021 , \33722_34022 , \33723_34023 , \33724_34024 , \33725_34025 , \33726_34026 ,
         \33727_34027 , \33728_34028 , \33729_34029 , \33730_34030 , \33731_34031 , \33732_34032 , \33733_34033 , \33734_34034 , \33735_34035 , \33736_34036 ,
         \33737_34037 , \33738_34038 , \33739_34039 , \33740_34040 , \33741_34041_nG9ba8 , \33742_34042 , \33743_34043 , \33744_34044 , \33745_34045 , \33746_34046 ,
         \33747_34047 , \33748_34048 , \33749_34049 , \33750_34050 , \33751_34051 , \33752_34052 , \33753_34053 , \33754_34054 , \33755_34055 , \33756_34056 ,
         \33757_34057 , \33758_34058 , \33759_34059 , \33760_34060 , \33761_34061 , \33762_34062 , \33763_34063 , \33764_34064 , \33765_34065 , \33766_34066 ,
         \33767_34067 , \33768_34068 , \33769_34069 , \33770_34070 , \33771_34071 , \33772_34072 , \33773_34073 , \33774_34074 , \33775_34075 , \33776_34076 ,
         \33777_34077 , \33778_34078 , \33779_34079 , \33780_34080 , \33781_34081 , \33782_34082 , \33783_34083 , \33784_34084 , \33785_34085 , \33786_34086 ,
         \33787_34087 , \33788_34088 , \33789_34089 , \33790_34090 , \33791_34091 , \33792_34092 , \33793_34093 , \33794_34094 , \33795_34095 , \33796_34096 ,
         \33797_34097 , \33798_34098 , \33799_34099 , \33800_34100 , \33801_34101 , \33802_34102 , \33803_34103 , \33804_34104 , \33805_34105 , \33806_34106 ,
         \33807_34107 , \33808_34108 , \33809_34109 , \33810_34110 , \33811_34111 , \33812_34112 , \33813_34113 , \33814_34114 , \33815_34115 , \33816_34116 ,
         \33817_34117 , \33818_34118 , \33819_34119 , \33820_34120 , \33821_34121 , \33822_34122 , \33823_34123 , \33824_34124 , \33825_34125 , \33826_34126 ,
         \33827_34127 , \33828_34128 , \33829_34129 , \33830_34130 , \33831_34131 , \33832_34132 , \33833_34133 , \33834_34134 , \33835_34135 , \33836_34136 ,
         \33837_34137 , \33838_34138 , \33839_34139 , \33840_34140 , \33841_34141 , \33842_34142 , \33843_34143 , \33844_34144 , \33845_34145 , \33846_34146 ,
         \33847_34147 , \33848_34148 , \33849_34149 , \33850_34150 , \33851_34151 , \33852_34152 , \33853_34153 , \33854_34154 , \33855_34155 , \33856_34156 ,
         \33857_34157 , \33858_34158 , \33859_34159 , \33860_34160 , \33861_34161 , \33862_34162 , \33863_34163 , \33864_34164 , \33865_34165 , \33866_34166 ,
         \33867_34167 , \33868_34168 , \33869_34169 , \33870_34170 , \33871_34171 , \33872_34172 , \33873_34173 , \33874_34174 , \33875_34175 , \33876_34176 ,
         \33877_34177 , \33878_34178 , \33879_34179 , \33880_34180 , \33881_34181 , \33882_34182 , \33883_34183 , \33884_34184 , \33885_34185 , \33886_34186 ,
         \33887_34187 , \33888_34188 , \33889_34189 , \33890_34190 , \33891_34191 , \33892_34192 , \33893_34193 , \33894_34194 , \33895_34195 , \33896_34196 ,
         \33897_34197 , \33898_34198 , \33899_34199 , \33900_34200 , \33901_34201 , \33902_34202 , \33903_34203 , \33904_34204 , \33905_34205 , \33906_34206 ,
         \33907_34207 , \33908_34208 , \33909_34209 , \33910_34210 , \33911_34211 , \33912_34212 , \33913_34213 , \33914_34214 , \33915_34215 , \33916_34216 ,
         \33917_34217 , \33918_34218 , \33919_34219 , \33920_34220 , \33921_34221 , \33922_34222 , \33923_34223 , \33924_34224 , \33925_34225 , \33926_34226 ,
         \33927_34227 , \33928_34228 , \33929_34229 , \33930_34230 , \33931_34231 , \33932_34232 , \33933_34233 , \33934_34234 , \33935_34235 , \33936_34236 ,
         \33937_34237 , \33938_34238 , \33939_34239 , \33940_34240 , \33941_34241 , \33942_34242 , \33943_34243 , \33944_34244 , \33945_34245 , \33946_34246 ,
         \33947_34247 , \33948_34248 , \33949_34249 , \33950_34250 , \33951_34251 , \33952_34252 , \33953_34253 , \33954_34254 , \33955_34255 , \33956_34256 ,
         \33957_34257 , \33958_34258 , \33959_34259 , \33960_34260 , \33961_34261 , \33962_34262 , \33963_34263 , \33964_34264 , \33965_34265 , \33966_34266 ,
         \33967_34267 , \33968_34268 , \33969_34269 , \33970_34270 , \33971_34271 , \33972_34272 , \33973_34273 , \33974_34274 , \33975_34275 , \33976_34276 ,
         \33977_34277 , \33978_34278 , \33979_34279 , \33980_34280 , \33981_34281 , \33982_34282 , \33983_34283 , \33984_34284 , \33985_34285 , \33986_34286 ,
         \33987_34287 , \33988_34288 , \33989_34289 , \33990_34290 , \33991_34291 , \33992_34292 , \33993_34293 , \33994_34294_nG9ba5 , \33995_34295 , \33996_34296 ,
         \33997_34297 , \33998_34298 , \33999_34299 , \34000_34300 , \34001_34301 , \34002_34302 , \34003_34303 , \34004_34304 , \34005_34305 , \34006_34306 ,
         \34007_34307 , \34008_34308 , \34009_34309 , \34010_34310 , \34011_34311 , \34012_34312 , \34013_34313 , \34014_34314 , \34015_34315 , \34016_34316 ,
         \34017_34317 , \34018_34318 , \34019_34319 , \34020_34320 , \34021_34321 , \34022_34322 , \34023_34323 , \34024_34324 , \34025_34325 , \34026_34326 ,
         \34027_34327 , \34028_34328 , \34029_34329 , \34030_34330 , \34031_34331 , \34032_34332 , \34033_34333 , \34034_34334 , \34035_34335 , \34036_34336 ,
         \34037_34337 , \34038_34338 , \34039_34339 , \34040_34340 , \34041_34341 , \34042_34342 , \34043_34343 , \34044_34344 , \34045_34345 , \34046_34346 ,
         \34047_34347 , \34048_34348 , \34049_34349 , \34050_34350 , \34051_34351 , \34052_34352 , \34053_34353 , \34054_34354 , \34055_34355 , \34056_34356 ,
         \34057_34357 , \34058_34358 , \34059_34359 , \34060_34360 , \34061_34361 , \34062_34362 , \34063_34363 , \34064_34364 , \34065_34365 , \34066_34366 ,
         \34067_34367 , \34068_34368 , \34069_34369 , \34070_34370 , \34071_34371 , \34072_34372 , \34073_34373 , \34074_34374 , \34075_34375 , \34076_34376 ,
         \34077_34377 , \34078_34378 , \34079_34379 , \34080_34380 , \34081_34381 , \34082_34382 , \34083_34383 , \34084_34384 , \34085_34385 , \34086_34386 ,
         \34087_34387 , \34088_34388 , \34089_34389 , \34090_34390 , \34091_34391 , \34092_34392 , \34093_34393 , \34094_34394 , \34095_34395 , \34096_34396 ,
         \34097_34397 , \34098_34398 , \34099_34399 , \34100_34400 , \34101_34401 , \34102_34402 , \34103_34403 , \34104_34404 , \34105_34405 , \34106_34406 ,
         \34107_34407 , \34108_34408 , \34109_34409 , \34110_34410 , \34111_34411 , \34112_34412 , \34113_34413 , \34114_34414 , \34115_34415 , \34116_34416 ,
         \34117_34417 , \34118_34418 , \34119_34419 , \34120_34420 , \34121_34421 , \34122_34422 , \34123_34423 , \34124_34424 , \34125_34425 , \34126_34426 ,
         \34127_34427 , \34128_34428 , \34129_34429 , \34130_34430 , \34131_34431 , \34132_34432 , \34133_34433 , \34134_34434 , \34135_34435 , \34136_34436 ,
         \34137_34437 , \34138_34438 , \34139_34439 , \34140_34440 , \34141_34441 , \34142_34442 , \34143_34443 , \34144_34444 , \34145_34445 , \34146_34446 ,
         \34147_34447 , \34148_34448 , \34149_34449 , \34150_34450 , \34151_34451 , \34152_34452 , \34153_34453 , \34154_34454 , \34155_34455 , \34156_34456 ,
         \34157_34457 , \34158_34458 , \34159_34459 , \34160_34460 , \34161_34461 , \34162_34462 , \34163_34463 , \34164_34464 , \34165_34465 , \34166_34466 ,
         \34167_34467 , \34168_34468 , \34169_34469 , \34170_34470 , \34171_34471 , \34172_34472 , \34173_34473 , \34174_34474 , \34175_34475 , \34176_34476 ,
         \34177_34477 , \34178_34478 , \34179_34479 , \34180_34480 , \34181_34481 , \34182_34482 , \34183_34483 , \34184_34484 , \34185_34485 , \34186_34486 ,
         \34187_34487 , \34188_34488 , \34189_34489 , \34190_34490 , \34191_34491 , \34192_34492 , \34193_34493 , \34194_34494 , \34195_34495 , \34196_34496 ,
         \34197_34497 , \34198_34498 , \34199_34499 , \34200_34500 , \34201_34501 , \34202_34502 , \34203_34503 , \34204_34504 , \34205_34505 , \34206_34506 ,
         \34207_34507 , \34208_34508 , \34209_34509 , \34210_34510 , \34211_34511 , \34212_34512 , \34213_34513 , \34214_34514 , \34215_34515 , \34216_34516 ,
         \34217_34517 , \34218_34518 , \34219_34519 , \34220_34520 , \34221_34521 , \34222_34522 , \34223_34523 , \34224_34524 , \34225_34525 , \34226_34526 ,
         \34227_34527 , \34228_34528 , \34229_34529 , \34230_34530 , \34231_34531 , \34232_34532 , \34233_34533 , \34234_34534 , \34235_34535 , \34236_34536 ,
         \34237_34537 , \34238_34538 , \34239_34539 , \34240_34540 , \34241_34541 , \34242_34542 , \34243_34543 , \34244_34544 , \34245_34545 , \34246_34546 ,
         \34247_34547 , \34248_34548 , \34249_34549 , \34250_34550 , \34251_34551 , \34252_34552 , \34253_34553 , \34254_34554 , \34255_34555 , \34256_34556 ,
         \34257_34557 , \34258_34558 , \34259_34559 , \34260_34560 , \34261_34561 , \34262_34562 , \34263_34563 , \34264_34564 , \34265_34565 , \34266_34566 ,
         \34267_34567 , \34268_34568 , \34269_34569 , \34270_34570 , \34271_34571 , \34272_34572 , \34273_34573 , \34274_34574 , \34275_34575 , \34276_34576 ,
         \34277_34577 , \34278_34578 , \34279_34579 , \34280_34580 , \34281_34581 , \34282_34582 , \34283_34583 , \34284_34584 , \34285_34585 , \34286_34586 ,
         \34287_34587 , \34288_34588 , \34289_34589 , \34290_34590 , \34291_34591 , \34292_34592 , \34293_34593 , \34294_34594 , \34295_34595 , \34296_34596 ,
         \34297_34597 , \34298_34598 , \34299_34599 , \34300_34600 , \34301_34601 , \34302_34602 , \34303_34603 , \34304_34604 , \34305_34605 , \34306_34606 ,
         \34307_34607 , \34308_34608 , \34309_34609 , \34310_34610 , \34311_34611 , \34312_34612 , \34313_34613 , \34314_34614 , \34315_34615 , \34316_34616 ,
         \34317_34617 , \34318_34618 , \34319_34619 , \34320_34620 , \34321_34621 , \34322_34622 , \34323_34623 , \34324_34624 , \34325_34625 , \34326_34626 ,
         \34327_34627 , \34328_34628 , \34329_34629 , \34330_34630 , \34331_34631 , \34332_34632 , \34333_34633 , \34334_34634 , \34335_34635 , \34336_34636 ,
         \34337_34637 , \34338_34638 , \34339_34639 , \34340_34640 , \34341_34641 , \34342_34642 , \34343_34643_nG9ba2 , \34344_34644 , \34345_34645 , \34346_34646 ,
         \34347_34647 , \34348_34648 , \34349_34649 , \34350_34650 , \34351_34651 , \34352_34652 , \34353_34653 , \34354_34654 , \34355_34655 , \34356_34656 ,
         \34357_34657 , \34358_34658 , \34359_34659 , \34360_34660 , \34361_34661 , \34362_34662 , \34363_34663 , \34364_34664 , \34365_34665 , \34366_34666 ,
         \34367_34667 , \34368_34668 , \34369_34669 , \34370_34670 , \34371_34671 , \34372_34672 , \34373_34673 , \34374_34674 , \34375_34675 , \34376_34676 ,
         \34377_34677 , \34378_34678 , \34379_34679 , \34380_34680 , \34381_34681 , \34382_34682 , \34383_34683 , \34384_34684 , \34385_34685 , \34386_34686 ,
         \34387_34687 , \34388_34688 , \34389_34689 , \34390_34690 , \34391_34691 , \34392_34692 , \34393_34693 , \34394_34694 , \34395_34695 , \34396_34696 ,
         \34397_34697 , \34398_34698 , \34399_34699 , \34400_34700 , \34401_34701 , \34402_34702 , \34403_34703 , \34404_34704 , \34405_34705 , \34406_34706 ,
         \34407_34707 , \34408_34708 , \34409_34709 , \34410_34710 , \34411_34711 , \34412_34712 , \34413_34713 , \34414_34714 , \34415_34715 , \34416_34716 ,
         \34417_34717 , \34418_34718 , \34419_34719 , \34420_34720 , \34421_34721 , \34422_34722 , \34423_34723 , \34424_34724 , \34425_34725 , \34426_34726 ,
         \34427_34727 , \34428_34728 , \34429_34729 , \34430_34730 , \34431_34731 , \34432_34732 , \34433_34733 , \34434_34734 , \34435_34735 , \34436_34736 ,
         \34437_34737 , \34438_34738 , \34439_34739 , \34440_34740 , \34441_34741 , \34442_34742 , \34443_34743 , \34444_34744 , \34445_34745 , \34446_34746 ,
         \34447_34747 , \34448_34748 , \34449_34749 , \34450_34750 , \34451_34751 , \34452_34752 , \34453_34753 , \34454_34754 , \34455_34755 , \34456_34756 ,
         \34457_34757 , \34458_34758 , \34459_34759 , \34460_34760 , \34461_34761 , \34462_34762 , \34463_34763 , \34464_34764 , \34465_34765 , \34466_34766 ,
         \34467_34767 , \34468_34768 , \34469_34769 , \34470_34770 , \34471_34771 , \34472_34772 , \34473_34773 , \34474_34774 , \34475_34775 , \34476_34776 ,
         \34477_34777 , \34478_34778 , \34479_34779 , \34480_34780 , \34481_34781 , \34482_34782 , \34483_34783 , \34484_34784 , \34485_34785 , \34486_34786 ,
         \34487_34787 , \34488_34788 , \34489_34789 , \34490_34790 , \34491_34791 , \34492_34792 , \34493_34793 , \34494_34794 , \34495_34795 , \34496_34796 ,
         \34497_34797 , \34498_34798 , \34499_34799 , \34500_34800 , \34501_34801 , \34502_34802 , \34503_34803 , \34504_34804 , \34505_34805 , \34506_34806 ,
         \34507_34807 , \34508_34808 , \34509_34809 , \34510_34810 , \34511_34811 , \34512_34812 , \34513_34813 , \34514_34814 , \34515_34815 , \34516_34816 ,
         \34517_34817 , \34518_34818 , \34519_34819 , \34520_34820 , \34521_34821 , \34522_34822 , \34523_34823 , \34524_34824 , \34525_34825 , \34526_34826 ,
         \34527_34827 , \34528_34828 , \34529_34829 , \34530_34830 , \34531_34831 , \34532_34832 , \34533_34833 , \34534_34834 , \34535_34835 , \34536_34836 ,
         \34537_34837 , \34538_34838 , \34539_34839 , \34540_34840 , \34541_34841 , \34542_34842 , \34543_34843 , \34544_34844 , \34545_34845 , \34546_34846 ,
         \34547_34847 , \34548_34848 , \34549_34849 , \34550_34850 , \34551_34851 , \34552_34852 , \34553_34853 , \34554_34854 , \34555_34855 , \34556_34856 ,
         \34557_34857 , \34558_34858 , \34559_34859 , \34560_34860 , \34561_34861 , \34562_34862 , \34563_34863 , \34564_34864 , \34565_34865 , \34566_34866 ,
         \34567_34867 , \34568_34868 , \34569_34869 , \34570_34870 , \34571_34871 , \34572_34872 , \34573_34873 , \34574_34874 , \34575_34875 , \34576_34876 ,
         \34577_34877 , \34578_34878 , \34579_34879 , \34580_34880 , \34581_34881 , \34582_34882 , \34583_34883 , \34584_34884 , \34585_34885 , \34586_34886 ,
         \34587_34887 , \34588_34888 , \34589_34889 , \34590_34890 , \34591_34891 , \34592_34892 , \34593_34893 , \34594_34894 , \34595_34895 , \34596_34896 ,
         \34597_34897 , \34598_34898 , \34599_34899 , \34600_34900 , \34601_34901 , \34602_34902 , \34603_34903 , \34604_34904 , \34605_34905 , \34606_34906 ,
         \34607_34907 , \34608_34908 , \34609_34909 , \34610_34910 , \34611_34911 , \34612_34912 , \34613_34913 , \34614_34914 , \34615_34915 , \34616_34916 ,
         \34617_34917 , \34618_34918 , \34619_34919 , \34620_34920 , \34621_34921 , \34622_34922 , \34623_34923 , \34624_34924 , \34625_34925 , \34626_34926 ,
         \34627_34927 , \34628_34928 , \34629_34929 , \34630_34930 , \34631_34931 , \34632_34932 , \34633_34933 , \34634_34934 , \34635_34935 , \34636_34936 ,
         \34637_34937 , \34638_34938 , \34639_34939 , \34640_34940 , \34641_34941 , \34642_34942 , \34643_34943 , \34644_34944 , \34645_34945 , \34646_34946 ,
         \34647_34947 , \34648_34948 , \34649_34949 , \34650_34950 , \34651_34951 , \34652_34952 , \34653_34953 , \34654_34954 , \34655_34955 , \34656_34956 ,
         \34657_34957 , \34658_34958 , \34659_34959 , \34660_34960 , \34661_34961 , \34662_34962 , \34663_34963 , \34664_34964 , \34665_34965 , \34666_34966 ,
         \34667_34967 , \34668_34968 , \34669_34969 , \34670_34970 , \34671_34971 , \34672_34972 , \34673_34973 , \34674_34974 , \34675_34975 , \34676_34976 ,
         \34677_34977 , \34678_34978 , \34679_34979 , \34680_34980 , \34681_34981 , \34682_34982 , \34683_34983 , \34684_34984 , \34685_34985 , \34686_34986 ,
         \34687_34987 , \34688_34988 , \34689_34989 , \34690_34990 , \34691_34991 , \34692_34992 , \34693_34993 , \34694_34994 , \34695_34995 , \34696_34996 ,
         \34697_34997 , \34698_34998 , \34699_34999 , \34700_35000 , \34701_35001 , \34702_35002 , \34703_35003 , \34704_35004 , \34705_35005 , \34706_35006 ,
         \34707_35007 , \34708_35008 , \34709_35009 , \34710_35010 , \34711_35011 , \34712_35012 , \34713_35013 , \34714_35014 , \34715_35015 , \34716_35016 ,
         \34717_35017 , \34718_35018 , \34719_35019 , \34720_35020 , \34721_35021 , \34722_35022 , \34723_35023 , \34724_35024 , \34725_35025 , \34726_35026 ,
         \34727_35027 , \34728_35028 , \34729_35029 , \34730_35030 , \34731_35031 , \34732_35032 , \34733_35033 , \34734_35034 , \34735_35035 , \34736_35036 ,
         \34737_35037 , \34738_35038 , \34739_35039 , \34740_35040 , \34741_35041 , \34742_35042 , \34743_35043 , \34744_35044 , \34745_35045 , \34746_35046 ,
         \34747_35047 , \34748_35048 , \34749_35049 , \34750_35050 , \34751_35051 , \34752_35052 , \34753_35053 , \34754_35054 , \34755_35055 , \34756_35056 ,
         \34757_35057 , \34758_35058 , \34759_35059 , \34760_35060 , \34761_35061 , \34762_35062 , \34763_35063 , \34764_35064 , \34765_35065 , \34766_35066 ,
         \34767_35067 , \34768_35068 , \34769_35069 , \34770_35070 , \34771_35071 , \34772_35072 , \34773_35073 , \34774_35074 , \34775_35075 , \34776_35076 ,
         \34777_35077 , \34778_35078 , \34779_35079 , \34780_35080 , \34781_35081 , \34782_35082 , \34783_35083 , \34784_35084 , \34785_35085 , \34786_35086 ,
         \34787_35087 , \34788_35088 , \34789_35089 , \34790_35090 , \34791_35091 , \34792_35092 , \34793_35093 , \34794_35094_nG9b9f , \34795_35095 , \34796_35096 ,
         \34797_35097 , \34798_35098 , \34799_35099 , \34800_35100 , \34801_35101 , \34802_35102 , \34803_35103 , \34804_35104 , \34805_35105 , \34806_35106 ,
         \34807_35107 , \34808_35108 , \34809_35109 , \34810_35110 , \34811_35111 , \34812_35112 , \34813_35113 , \34814_35114 , \34815_35115 , \34816_35116 ,
         \34817_35117 , \34818_35118 , \34819_35119 , \34820_35120 , \34821_35121 , \34822_35122 , \34823_35123 , \34824_35124 , \34825_35125 , \34826_35126 ,
         \34827_35127 , \34828_35128 , \34829_35129 , \34830_35130 , \34831_35131 , \34832_35132 , \34833_35133 , \34834_35134 , \34835_35135 , \34836_35136 ,
         \34837_35137 , \34838_35138 , \34839_35139 , \34840_35140 , \34841_35141 , \34842_35142 , \34843_35143 , \34844_35144 , \34845_35145 , \34846_35146 ,
         \34847_35147 , \34848_35148 , \34849_35149 , \34850_35150 , \34851_35151 , \34852_35152 , \34853_35153 , \34854_35154 , \34855_35155 , \34856_35156 ,
         \34857_35157 , \34858_35158 , \34859_35159 , \34860_35160 , \34861_35161 , \34862_35162 , \34863_35163 , \34864_35164 , \34865_35165 , \34866_35166 ,
         \34867_35167 , \34868_35168 , \34869_35169 , \34870_35170 , \34871_35171 , \34872_35172 , \34873_35173 , \34874_35174 , \34875_35175 , \34876_35176 ,
         \34877_35177 , \34878_35178 , \34879_35179 , \34880_35180 , \34881_35181 , \34882_35182 , \34883_35183 , \34884_35184 , \34885_35185 , \34886_35186 ,
         \34887_35187 , \34888_35188 , \34889_35189 , \34890_35190 , \34891_35191 , \34892_35192 , \34893_35193 , \34894_35194 , \34895_35195 , \34896_35196 ,
         \34897_35197 , \34898_35198 , \34899_35199 , \34900_35200 , \34901_35201 , \34902_35202 , \34903_35203 , \34904_35204 , \34905_35205 , \34906_35206 ,
         \34907_35207 , \34908_35208 , \34909_35209 , \34910_35210 , \34911_35211 , \34912_35212 , \34913_35213 , \34914_35214 , \34915_35215 , \34916_35216 ,
         \34917_35217 , \34918_35218 , \34919_35219 , \34920_35220 , \34921_35221 , \34922_35222 , \34923_35223 , \34924_35224 , \34925_35225 , \34926_35226 ,
         \34927_35227 , \34928_35228 , \34929_35229 , \34930_35230 , \34931_35231 , \34932_35232 , \34933_35233 , \34934_35234 , \34935_35235 , \34936_35236 ,
         \34937_35237 , \34938_35238 , \34939_35239 , \34940_35240 , \34941_35241 , \34942_35242 , \34943_35243 , \34944_35244 , \34945_35245 , \34946_35246 ,
         \34947_35247 , \34948_35248 , \34949_35249 , \34950_35250 , \34951_35251 , \34952_35252 , \34953_35253 , \34954_35254 , \34955_35255 , \34956_35256 ,
         \34957_35257 , \34958_35258 , \34959_35259 , \34960_35260 , \34961_35261 , \34962_35262 , \34963_35263 , \34964_35264 , \34965_35265 , \34966_35266 ,
         \34967_35267 , \34968_35268 , \34969_35269 , \34970_35270 , \34971_35271 , \34972_35272 , \34973_35273 , \34974_35274 , \34975_35275 , \34976_35276 ,
         \34977_35277 , \34978_35278 , \34979_35279 , \34980_35280 , \34981_35281 , \34982_35282 , \34983_35283 , \34984_35284 , \34985_35285 , \34986_35286 ,
         \34987_35287 , \34988_35288 , \34989_35289 , \34990_35290 , \34991_35291 , \34992_35292 , \34993_35293 , \34994_35294 , \34995_35295 , \34996_35296 ,
         \34997_35297 , \34998_35298 , \34999_35299 , \35000_35300 , \35001_35301 , \35002_35302 , \35003_35303 , \35004_35304 , \35005_35305 , \35006_35306 ,
         \35007_35307 , \35008_35308 , \35009_35309 , \35010_35310 , \35011_35311 , \35012_35312 , \35013_35313 , \35014_35314 , \35015_35315 , \35016_35316 ,
         \35017_35317 , \35018_35318 , \35019_35319 , \35020_35320 , \35021_35321 , \35022_35322 , \35023_35323 , \35024_35324 , \35025_35325 , \35026_35326 ,
         \35027_35327 , \35028_35328 , \35029_35329 , \35030_35330 , \35031_35331 , \35032_35332 , \35033_35333 , \35034_35334 , \35035_35335 , \35036_35336 ,
         \35037_35337 , \35038_35338 , \35039_35339 , \35040_35340 , \35041_35341 , \35042_35342 , \35043_35343 , \35044_35344 , \35045_35345 , \35046_35346 ,
         \35047_35347 , \35048_35348 , \35049_35349 , \35050_35350 , \35051_35351 , \35052_35352 , \35053_35353 , \35054_35354 , \35055_35355 , \35056_35356 ,
         \35057_35357 , \35058_35358 , \35059_35359 , \35060_35360 , \35061_35361 , \35062_35362 , \35063_35363 , \35064_35364 , \35065_35365 , \35066_35366 ,
         \35067_35367 , \35068_35368 , \35069_35369 , \35070_35370 , \35071_35371 , \35072_35372 , \35073_35373 , \35074_35374 , \35075_35375 , \35076_35376 ,
         \35077_35377 , \35078_35378 , \35079_35379 , \35080_35380 , \35081_35381 , \35082_35382 , \35083_35383 , \35084_35384 , \35085_35385 , \35086_35386 ,
         \35087_35387 , \35088_35388 , \35089_35389 , \35090_35390 , \35091_35391 , \35092_35392 , \35093_35393 , \35094_35394 , \35095_35395 , \35096_35396 ,
         \35097_35397 , \35098_35398 , \35099_35399 , \35100_35400 , \35101_35401 , \35102_35402 , \35103_35403 , \35104_35404 , \35105_35405 , \35106_35406 ,
         \35107_35407 , \35108_35408 , \35109_35409 , \35110_35410 , \35111_35411 , \35112_35412 , \35113_35413 , \35114_35414 , \35115_35415 , \35116_35416 ,
         \35117_35417 , \35118_35418 , \35119_35419 , \35120_35420 , \35121_35421 , \35122_35422 , \35123_35423 , \35124_35424 , \35125_35425 , \35126_35426 ,
         \35127_35427 , \35128_35428 , \35129_35429 , \35130_35430 , \35131_35431 , \35132_35432 , \35133_35433 , \35134_35434 , \35135_35435 , \35136_35436 ,
         \35137_35437 , \35138_35438 , \35139_35439 , \35140_35440 , \35141_35441 , \35142_35442 , \35143_35443 , \35144_35444 , \35145_35445 , \35146_35446 ,
         \35147_35447 , \35148_35448 , \35149_35449 , \35150_35450 , \35151_35451 , \35152_35452 , \35153_35453 , \35154_35454 , \35155_35455 , \35156_35456 ,
         \35157_35457 , \35158_35458 , \35159_35459 , \35160_35460 , \35161_35461 , \35162_35462 , \35163_35463 , \35164_35464 , \35165_35465 , \35166_35466 ,
         \35167_35467 , \35168_35468 , \35169_35469 , \35170_35470 , \35171_35471 , \35172_35472 , \35173_35473 , \35174_35474 , \35175_35475 , \35176_35476 ,
         \35177_35477 , \35178_35478 , \35179_35479 , \35180_35480 , \35181_35481 , \35182_35482 , \35183_35483 , \35184_35484 , \35185_35485 , \35186_35486 ,
         \35187_35487 , \35188_35488 , \35189_35489 , \35190_35490 , \35191_35491 , \35192_35492 , \35193_35493 , \35194_35494 , \35195_35495 , \35196_35496 ,
         \35197_35497 , \35198_35498 , \35199_35499 , \35200_35500 , \35201_35501 , \35202_35502 , \35203_35503 , \35204_35504 , \35205_35505 , \35206_35506 ,
         \35207_35507 , \35208_35508 , \35209_35509 , \35210_35510 , \35211_35511 , \35212_35512 , \35213_35513 , \35214_35514 , \35215_35515 , \35216_35516 ,
         \35217_35517 , \35218_35518 , \35219_35519 , \35220_35520 , \35221_35521 , \35222_35522 , \35223_35523 , \35224_35524 , \35225_35525 , \35226_35526 ,
         \35227_35527 , \35228_35528 , \35229_35529 , \35230_35530 , \35231_35531 , \35232_35532 , \35233_35533 , \35234_35534 , \35235_35535 , \35236_35536 ,
         \35237_35537 , \35238_35538 , \35239_35539 , \35240_35540 , \35241_35541 , \35242_35542 , \35243_35543 , \35244_35544 , \35245_35545 , \35246_35546 ,
         \35247_35547 , \35248_35548 , \35249_35549 , \35250_35550 , \35251_35551 , \35252_35552 , \35253_35553 , \35254_35554 , \35255_35555 , \35256_35556 ,
         \35257_35557 , \35258_35558 , \35259_35559 , \35260_35560 , \35261_35561 , \35262_35562 , \35263_35563 , \35264_35564 , \35265_35565 , \35266_35566 ,
         \35267_35567 , \35268_35568 , \35269_35569 , \35270_35570_nG9b9c , \35271_35571 , \35272_35572 , \35273_35573 , \35274_35574 , \35275_35575 , \35276_35576 ,
         \35277_35577 , \35278_35578 , \35279_35579 , \35280_35580 , \35281_35581 , \35282_35582 , \35283_35583 , \35284_35584 , \35285_35585 , \35286_35586 ,
         \35287_35587 , \35288_35588 , \35289_35589 , \35290_35590 , \35291_35591 , \35292_35592 , \35293_35593 , \35294_35594 , \35295_35595 , \35296_35596 ,
         \35297_35597 , \35298_35598 , \35299_35599 , \35300_35600 , \35301_35601 , \35302_35602 , \35303_35603 , \35304_35604 , \35305_35605 , \35306_35606 ,
         \35307_35607 , \35308_35608 , \35309_35609 , \35310_35610 , \35311_35611 , \35312_35612 , \35313_35613 , \35314_35614 , \35315_35615 , \35316_35616 ,
         \35317_35617 , \35318_35618 , \35319_35619 , \35320_35620 , \35321_35621 , \35322_35622 , \35323_35623 , \35324_35624 , \35325_35625 , \35326_35626 ,
         \35327_35627 , \35328_35628 , \35329_35629 , \35330_35630 , \35331_35631 , \35332_35632 , \35333_35633 , \35334_35634 , \35335_35635 , \35336_35636 ,
         \35337_35637 , \35338_35638 , \35339_35639 , \35340_35640 , \35341_35641 , \35342_35642 , \35343_35643 , \35344_35644 , \35345_35645 , \35346_35646 ,
         \35347_35647 , \35348_35648 , \35349_35649 , \35350_35650 , \35351_35651 , \35352_35652 , \35353_35653 , \35354_35654 , \35355_35655 , \35356_35656 ,
         \35357_35657 , \35358_35658 , \35359_35659 , \35360_35660 , \35361_35661 , \35362_35662 , \35363_35663 , \35364_35664 , \35365_35665 , \35366_35666 ,
         \35367_35667 , \35368_35668 , \35369_35669 , \35370_35670 , \35371_35671 , \35372_35672 , \35373_35673 , \35374_35674 , \35375_35675 , \35376_35676 ,
         \35377_35677 , \35378_35678 , \35379_35679 , \35380_35680 , \35381_35681 , \35382_35682 , \35383_35683 , \35384_35684 , \35385_35685 , \35386_35686 ,
         \35387_35687 , \35388_35688 , \35389_35689 , \35390_35690 , \35391_35691 , \35392_35692 , \35393_35693 , \35394_35694 , \35395_35695 , \35396_35696 ,
         \35397_35697 , \35398_35698 , \35399_35699 , \35400_35700 , \35401_35701 , \35402_35702 , \35403_35703 , \35404_35704 , \35405_35705 , \35406_35706 ,
         \35407_35707 , \35408_35708 , \35409_35709 , \35410_35710 , \35411_35711 , \35412_35712 , \35413_35713 , \35414_35714 , \35415_35715 , \35416_35716 ,
         \35417_35717 , \35418_35718 , \35419_35719 , \35420_35720 , \35421_35721 , \35422_35722 , \35423_35723 , \35424_35724 , \35425_35725 , \35426_35726 ,
         \35427_35727 , \35428_35728 , \35429_35729 , \35430_35730 , \35431_35731 , \35432_35732 , \35433_35733 , \35434_35734 , \35435_35735 , \35436_35736 ,
         \35437_35737 , \35438_35738 , \35439_35739 , \35440_35740 , \35441_35741 , \35442_35742 , \35443_35743 , \35444_35744 , \35445_35745 , \35446_35746 ,
         \35447_35747 , \35448_35748 , \35449_35749 , \35450_35750 , \35451_35751 , \35452_35752 , \35453_35753 , \35454_35754 , \35455_35755 , \35456_35756 ,
         \35457_35757 , \35458_35758 , \35459_35759 , \35460_35760 , \35461_35761 , \35462_35762 , \35463_35763 , \35464_35764 , \35465_35765 , \35466_35766 ,
         \35467_35767 , \35468_35768 , \35469_35769 , \35470_35770 , \35471_35771 , \35472_35772 , \35473_35773 , \35474_35774 , \35475_35775 , \35476_35776 ,
         \35477_35777 , \35478_35778 , \35479_35779 , \35480_35780 , \35481_35781 , \35482_35782 , \35483_35783 , \35484_35784 , \35485_35785 , \35486_35786 ,
         \35487_35787 , \35488_35788 , \35489_35789 , \35490_35790 , \35491_35791 , \35492_35792 , \35493_35793 , \35494_35794 , \35495_35795 , \35496_35796 ,
         \35497_35797 , \35498_35798 , \35499_35799 , \35500_35800 , \35501_35801_nG9b99 , \35502_35802 , \35503_35803 , \35504_35804 , \35505_35805 , \35506_35806 ,
         \35507_35807 , \35508_35808 , \35509_35809 , \35510_35810 , \35511_35811 , \35512_35812 , \35513_35813 , \35514_35814 , \35515_35815 , \35516_35816 ,
         \35517_35817 , \35518_35818 , \35519_35819 , \35520_35820 , \35521_35821 , \35522_35822 , \35523_35823 , \35524_35824 , \35525_35825 , \35526_35826 ,
         \35527_35827 , \35528_35828 , \35529_35829 , \35530_35830 , \35531_35831 , \35532_35832 , \35533_35833 , \35534_35834 , \35535_35835 , \35536_35836 ,
         \35537_35837 , \35538_35838 , \35539_35839 , \35540_35840 , \35541_35841 , \35542_35842 , \35543_35843 , \35544_35844 , \35545_35845 , \35546_35846 ,
         \35547_35847 , \35548_35848 , \35549_35849 , \35550_35850 , \35551_35851 , \35552_35852 , \35553_35853 , \35554_35854 , \35555_35855 , \35556_35856 ,
         \35557_35857 , \35558_35858 , \35559_35859 , \35560_35860 , \35561_35861 , \35562_35862 , \35563_35863 , \35564_35864 , \35565_35865 , \35566_35866 ,
         \35567_35867 , \35568_35868 , \35569_35869 , \35570_35870 , \35571_35871 , \35572_35872 , \35573_35873 , \35574_35874 , \35575_35875 , \35576_35876 ,
         \35577_35877 , \35578_35878 , \35579_35879 , \35580_35880 , \35581_35881 , \35582_35882 , \35583_35883 , \35584_35884 , \35585_35885 , \35586_35886 ,
         \35587_35887 , \35588_35888 , \35589_35889 , \35590_35890 , \35591_35891 , \35592_35892 , \35593_35893 , \35594_35894 , \35595_35895 , \35596_35896 ,
         \35597_35897 , \35598_35898 , \35599_35899 , \35600_35900 , \35601_35901 , \35602_35902 , \35603_35903 , \35604_35904 , \35605_35905 , \35606_35906 ,
         \35607_35907 , \35608_35908 , \35609_35909 , \35610_35910 , \35611_35911 , \35612_35912 , \35613_35913 , \35614_35914 , \35615_35915 , \35616_35916 ,
         \35617_35917 , \35618_35918 , \35619_35919 , \35620_35920 , \35621_35921 , \35622_35922 , \35623_35923 , \35624_35924 , \35625_35925 , \35626_35926 ,
         \35627_35927 , \35628_35928 , \35629_35929 , \35630_35930 , \35631_35931 , \35632_35932 , \35633_35933 , \35634_35934 , \35635_35935 , \35636_35936 ,
         \35637_35937 , \35638_35938 , \35639_35939 , \35640_35940 , \35641_35941 , \35642_35942 , \35643_35943 , \35644_35944 , \35645_35945 , \35646_35946 ,
         \35647_35947 , \35648_35948 , \35649_35949 , \35650_35950 , \35651_35951 , \35652_35952 , \35653_35953 , \35654_35954 , \35655_35955 , \35656_35956 ,
         \35657_35957 , \35658_35958 , \35659_35959 , \35660_35960 , \35661_35961 , \35662_35962 , \35663_35963 , \35664_35964 , \35665_35965 , \35666_35966 ,
         \35667_35967 , \35668_35968 , \35669_35969 , \35670_35970 , \35671_35971 , \35672_35972 , \35673_35973 , \35674_35974 , \35675_35975 , \35676_35976 ,
         \35677_35977 , \35678_35978 , \35679_35979 , \35680_35980 , \35681_35981 , \35682_35982 , \35683_35983 , \35684_35984 , \35685_35985 , \35686_35986 ,
         \35687_35987 , \35688_35988 , \35689_35989 , \35690_35990 , \35691_35991 , \35692_35992 , \35693_35993 , \35694_35994 , \35695_35995 , \35696_35996 ,
         \35697_35997 , \35698_35998 , \35699_35999 , \35700_36000 , \35701_36001 , \35702_36002 , \35703_36003 , \35704_36004 , \35705_36005 , \35706_36006 ,
         \35707_36007 , \35708_36008 , \35709_36009 , \35710_36010 , \35711_36011 , \35712_36012 , \35713_36013 , \35714_36014 , \35715_36015 , \35716_36016 ,
         \35717_36017 , \35718_36018 , \35719_36019 , \35720_36020 , \35721_36021 , \35722_36022 , \35723_36023 , \35724_36024 , \35725_36025 , \35726_36026 ,
         \35727_36027 , \35728_36028 , \35729_36029 , \35730_36030 , \35731_36031 , \35732_36032 , \35733_36033 , \35734_36034 , \35735_36035 , \35736_36036 ,
         \35737_36037 , \35738_36038 , \35739_36039 , \35740_36040 , \35741_36041 , \35742_36042 , \35743_36043 , \35744_36044 , \35745_36045 , \35746_36046 ,
         \35747_36047 , \35748_36048 , \35749_36049 , \35750_36050 , \35751_36051 , \35752_36052 , \35753_36053 , \35754_36054 , \35755_36055 , \35756_36056 ,
         \35757_36057 , \35758_36058 , \35759_36059 , \35760_36060 , \35761_36061 , \35762_36062 , \35763_36063 , \35764_36064 , \35765_36065 , \35766_36066 ,
         \35767_36067 , \35768_36068 , \35769_36069 , \35770_36070 , \35771_36071 , \35772_36072 , \35773_36073 , \35774_36074 , \35775_36075 , \35776_36076 ,
         \35777_36077 , \35778_36078 , \35779_36079 , \35780_36080 , \35781_36081 , \35782_36082 , \35783_36083 , \35784_36084 , \35785_36085 , \35786_36086 ,
         \35787_36087 , \35788_36088 , \35789_36089 , \35790_36090 , \35791_36091 , \35792_36092 , \35793_36093 , \35794_36094 , \35795_36095 , \35796_36096 ,
         \35797_36097 , \35798_36098 , \35799_36099 , \35800_36100 , \35801_36101 , \35802_36102 , \35803_36103 , \35804_36104 , \35805_36105 , \35806_36106 ,
         \35807_36107 , \35808_36108 , \35809_36109 , \35810_36110 , \35811_36111 , \35812_36112 , \35813_36113 , \35814_36114 , \35815_36115 , \35816_36116 ,
         \35817_36117 , \35818_36118 , \35819_36119 , \35820_36120 , \35821_36121 , \35822_36122 , \35823_36123 , \35824_36124 , \35825_36125 , \35826_36126 ,
         \35827_36127 , \35828_36128 , \35829_36129 , \35830_36130 , \35831_36131 , \35832_36132 , \35833_36133 , \35834_36134 , \35835_36135 , \35836_36136 ,
         \35837_36137 , \35838_36138 , \35839_36139 , \35840_36140 , \35841_36141 , \35842_36142 , \35843_36143 , \35844_36144 , \35845_36145 , \35846_36146 ,
         \35847_36147 , \35848_36148 , \35849_36149 , \35850_36150 , \35851_36151 , \35852_36152 , \35853_36153 , \35854_36154 , \35855_36155 , \35856_36156 ,
         \35857_36157 , \35858_36158 , \35859_36159 , \35860_36160 , \35861_36161 , \35862_36162 , \35863_36163 , \35864_36164 , \35865_36165 , \35866_36166 ,
         \35867_36167 , \35868_36168 , \35869_36169 , \35870_36170 , \35871_36171 , \35872_36172_nG9b96 , \35873_36173 , \35874_36174 , \35875_36175 , \35876_36176 ,
         \35877_36177 , \35878_36178 , \35879_36179 , \35880_36180 , \35881_36181 , \35882_36182 , \35883_36183 , \35884_36184 , \35885_36185 , \35886_36186 ,
         \35887_36187 , \35888_36188 , \35889_36189 , \35890_36190 , \35891_36191 , \35892_36192 , \35893_36193 , \35894_36194 , \35895_36195 , \35896_36196 ,
         \35897_36197 , \35898_36198 , \35899_36199 , \35900_36200 , \35901_36201 , \35902_36202 , \35903_36203 , \35904_36204 , \35905_36205 , \35906_36206 ,
         \35907_36207 , \35908_36208 , \35909_36209 , \35910_36210 , \35911_36211 , \35912_36212 , \35913_36213 , \35914_36214 , \35915_36215 , \35916_36216 ,
         \35917_36217 , \35918_36218 , \35919_36219 , \35920_36220 , \35921_36221 , \35922_36222 , \35923_36223 , \35924_36224 , \35925_36225 , \35926_36226 ,
         \35927_36227 , \35928_36228 , \35929_36229 , \35930_36230 , \35931_36231 , \35932_36232 , \35933_36233 , \35934_36234 , \35935_36235 , \35936_36236 ,
         \35937_36237 , \35938_36238 , \35939_36239 , \35940_36240 , \35941_36241 , \35942_36242 , \35943_36243 , \35944_36244 , \35945_36245 , \35946_36246 ,
         \35947_36247 , \35948_36248 , \35949_36249 , \35950_36250 , \35951_36251 , \35952_36252 , \35953_36253 , \35954_36254 , \35955_36255 , \35956_36256 ,
         \35957_36257 , \35958_36258 , \35959_36259 , \35960_36260 , \35961_36261 , \35962_36262 , \35963_36263 , \35964_36264 , \35965_36265 , \35966_36266 ,
         \35967_36267 , \35968_36268 , \35969_36269 , \35970_36270 , \35971_36271 , \35972_36272 , \35973_36273 , \35974_36274 , \35975_36275 , \35976_36276 ,
         \35977_36277 , \35978_36278 , \35979_36279 , \35980_36280 , \35981_36281 , \35982_36282 , \35983_36283 , \35984_36284 , \35985_36285 , \35986_36286 ,
         \35987_36287 , \35988_36288 , \35989_36289 , \35990_36290 , \35991_36291 , \35992_36292 , \35993_36293 , \35994_36294 , \35995_36295 , \35996_36296 ,
         \35997_36297 , \35998_36298 , \35999_36299 , \36000_36300 , \36001_36301 , \36002_36302 , \36003_36303 , \36004_36304 , \36005_36305 , \36006_36306 ,
         \36007_36307 , \36008_36308 , \36009_36309 , \36010_36310 , \36011_36311 , \36012_36312 , \36013_36313 , \36014_36314 , \36015_36315 , \36016_36316 ,
         \36017_36317 , \36018_36318 , \36019_36319 , \36020_36320 , \36021_36321 , \36022_36322 , \36023_36323 , \36024_36324 , \36025_36325 , \36026_36326 ,
         \36027_36327 , \36028_36328 , \36029_36329 , \36030_36330 , \36031_36331 , \36032_36332 , \36033_36333 , \36034_36334 , \36035_36335 , \36036_36336 ,
         \36037_36337 , \36038_36338 , \36039_36339 , \36040_36340 , \36041_36341 , \36042_36342 , \36043_36343 , \36044_36344 , \36045_36345 , \36046_36346 ,
         \36047_36347 , \36048_36348 , \36049_36349 , \36050_36350 , \36051_36351 , \36052_36352 , \36053_36353 , \36054_36354 , \36055_36355 , \36056_36356 ,
         \36057_36357 , \36058_36358 , \36059_36359 , \36060_36360 , \36061_36361 , \36062_36362 , \36063_36363 , \36064_36364 , \36065_36365 , \36066_36366 ,
         \36067_36367 , \36068_36368 , \36069_36369 , \36070_36370 , \36071_36371 , \36072_36372 , \36073_36373 , \36074_36374 , \36075_36375 , \36076_36376 ,
         \36077_36377 , \36078_36378 , \36079_36379 , \36080_36380 , \36081_36381 , \36082_36382 , \36083_36383 , \36084_36384 , \36085_36385 , \36086_36386 ,
         \36087_36387 , \36088_36388 , \36089_36389 , \36090_36390 , \36091_36391 , \36092_36392 , \36093_36393 , \36094_36394 , \36095_36395 , \36096_36396 ,
         \36097_36397 , \36098_36398 , \36099_36399 , \36100_36400 , \36101_36401 , \36102_36402 , \36103_36403 , \36104_36404 , \36105_36405 , \36106_36406 ,
         \36107_36407 , \36108_36408 , \36109_36409 , \36110_36410 , \36111_36411 , \36112_36412 , \36113_36413 , \36114_36414 , \36115_36415 , \36116_36416 ,
         \36117_36417 , \36118_36418 , \36119_36419 , \36120_36420 , \36121_36421 , \36122_36422 , \36123_36423 , \36124_36424 , \36125_36425 , \36126_36426 ,
         \36127_36427 , \36128_36428 , \36129_36429 , \36130_36430 , \36131_36431 , \36132_36432 , \36133_36433 , \36134_36434 , \36135_36435 , \36136_36436 ,
         \36137_36437 , \36138_36438 , \36139_36439 , \36140_36440 , \36141_36441 , \36142_36442 , \36143_36443 , \36144_36444 , \36145_36445 , \36146_36446 ,
         \36147_36447 , \36148_36448 , \36149_36449 , \36150_36450 , \36151_36451 , \36152_36452 , \36153_36453 , \36154_36454 , \36155_36455 , \36156_36456 ,
         \36157_36457 , \36158_36458 , \36159_36459 , \36160_36460 , \36161_36461 , \36162_36462 , \36163_36463 , \36164_36464 , \36165_36465 , \36166_36466 ,
         \36167_36467 , \36168_36468 , \36169_36469 , \36170_36470 , \36171_36471 , \36172_36472 , \36173_36473 , \36174_36474 , \36175_36475 , \36176_36476 ,
         \36177_36477 , \36178_36478 , \36179_36479 , \36180_36480 , \36181_36481 , \36182_36482 , \36183_36483 , \36184_36484 , \36185_36485 , \36186_36486 ,
         \36187_36487 , \36188_36488 , \36189_36489 , \36190_36490 , \36191_36491 , \36192_36492 , \36193_36493 , \36194_36494 , \36195_36495 , \36196_36496 ,
         \36197_36497 , \36198_36498 , \36199_36499 , \36200_36500 , \36201_36501 , \36202_36502 , \36203_36503 , \36204_36504 , \36205_36505 , \36206_36506 ,
         \36207_36507 , \36208_36508 , \36209_36509 , \36210_36510 , \36211_36511 , \36212_36512 , \36213_36513 , \36214_36514 , \36215_36515 , \36216_36516 ,
         \36217_36517 , \36218_36518 , \36219_36519 , \36220_36520 , \36221_36521 , \36222_36522 , \36223_36523 , \36224_36524 , \36225_36525 , \36226_36526 ,
         \36227_36527 , \36228_36528 , \36229_36529 , \36230_36530 , \36231_36531 , \36232_36532 , \36233_36533 , \36234_36534 , \36235_36535 , \36236_36536 ,
         \36237_36537 , \36238_36538 , \36239_36539 , \36240_36540 , \36241_36541 , \36242_36542 , \36243_36543 , \36244_36544 , \36245_36545 , \36246_36546 ,
         \36247_36547 , \36248_36548 , \36249_36549 , \36250_36550 , \36251_36551 , \36252_36552 , \36253_36553 , \36254_36554 , \36255_36555 , \36256_36556 ,
         \36257_36557 , \36258_36558 , \36259_36559 , \36260_36560 , \36261_36561 , \36262_36562 , \36263_36563 , \36264_36564 , \36265_36565 , \36266_36566 ,
         \36267_36567 , \36268_36568 , \36269_36569 , \36270_36570 , \36271_36571 , \36272_36572 , \36273_36573 , \36274_36574 , \36275_36575 , \36276_36576 ,
         \36277_36577 , \36278_36578 , \36279_36579 , \36280_36580 , \36281_36581 , \36282_36582 , \36283_36583 , \36284_36584 , \36285_36585 , \36286_36586 ,
         \36287_36587 , \36288_36588 , \36289_36589_nG9b93 , \36290_36590 , \36291_36591 , \36292_36592 , \36293_36593 , \36294_36594 , \36295_36595 , \36296_36596 ,
         \36297_36597 , \36298_36598 , \36299_36599 , \36300_36600 , \36301_36601 , \36302_36602 , \36303_36603 , \36304_36604 , \36305_36605 , \36306_36606 ,
         \36307_36607 , \36308_36608 , \36309_36609 , \36310_36610 , \36311_36611 , \36312_36612 , \36313_36613 , \36314_36614 , \36315_36615 , \36316_36616 ,
         \36317_36617 , \36318_36618 , \36319_36619 , \36320_36620 , \36321_36621 , \36322_36622 , \36323_36623 , \36324_36624 , \36325_36625 , \36326_36626 ,
         \36327_36627 , \36328_36628 , \36329_36629 , \36330_36630 , \36331_36631 , \36332_36632 , \36333_36633 , \36334_36634 , \36335_36635 , \36336_36636 ,
         \36337_36637 , \36338_36638 , \36339_36639 , \36340_36640 , \36341_36641 , \36342_36642 , \36343_36643 , \36344_36644 , \36345_36645 , \36346_36646 ,
         \36347_36647 , \36348_36648 , \36349_36649 , \36350_36650 , \36351_36651 , \36352_36652 , \36353_36653 , \36354_36654 , \36355_36655 , \36356_36656 ,
         \36357_36657 , \36358_36658 , \36359_36659 , \36360_36660 , \36361_36661 , \36362_36662 , \36363_36663 , \36364_36664 , \36365_36665 , \36366_36666 ,
         \36367_36667 , \36368_36668 , \36369_36669 , \36370_36670 , \36371_36671 , \36372_36672 , \36373_36673 , \36374_36674 , \36375_36675 , \36376_36676 ,
         \36377_36677 , \36378_36678 , \36379_36679 , \36380_36680 , \36381_36681 , \36382_36682 , \36383_36683 , \36384_36684 , \36385_36685 , \36386_36686 ,
         \36387_36687 , \36388_36688 , \36389_36689 , \36390_36690 , \36391_36691 , \36392_36692 , \36393_36693 , \36394_36694 , \36395_36695 , \36396_36696 ,
         \36397_36697 , \36398_36698 , \36399_36699 , \36400_36700 , \36401_36701 , \36402_36702 , \36403_36703 , \36404_36704 , \36405_36705 , \36406_36706 ,
         \36407_36707 , \36408_36708 , \36409_36709 , \36410_36710 , \36411_36711 , \36412_36712 , \36413_36713 , \36414_36714 , \36415_36715 , \36416_36716 ,
         \36417_36717 , \36418_36718 , \36419_36719 , \36420_36720 , \36421_36721 , \36422_36722 , \36423_36723 , \36424_36724 , \36425_36725 , \36426_36726 ,
         \36427_36727 , \36428_36728 , \36429_36729 , \36430_36730 , \36431_36731 , \36432_36732 , \36433_36733 , \36434_36734 , \36435_36735 , \36436_36736 ,
         \36437_36737 , \36438_36738 , \36439_36739 , \36440_36740 , \36441_36741 , \36442_36742 , \36443_36743 , \36444_36744 , \36445_36745 , \36446_36746 ,
         \36447_36747 , \36448_36748 , \36449_36749 , \36450_36750 , \36451_36751 , \36452_36752 , \36453_36753 , \36454_36754 , \36455_36755 , \36456_36756 ,
         \36457_36757 , \36458_36758 , \36459_36759 , \36460_36760 , \36461_36761 , \36462_36762 , \36463_36763 , \36464_36764 , \36465_36765 , \36466_36766 ,
         \36467_36767 , \36468_36768 , \36469_36769 , \36470_36770 , \36471_36771 , \36472_36772 , \36473_36773 , \36474_36774 , \36475_36775 , \36476_36776 ,
         \36477_36777 , \36478_36778 , \36479_36779 , \36480_36780 , \36481_36781 , \36482_36782 , \36483_36783 , \36484_36784 , \36485_36785 , \36486_36786 ,
         \36487_36787 , \36488_36788 , \36489_36789 , \36490_36790 , \36491_36791 , \36492_36792 , \36493_36793 , \36494_36794 , \36495_36795 , \36496_36796 ,
         \36497_36797 , \36498_36798 , \36499_36799 , \36500_36800 , \36501_36801 , \36502_36802 , \36503_36803 , \36504_36804 , \36505_36805 , \36506_36806 ,
         \36507_36807 , \36508_36808 , \36509_36809 , \36510_36810 , \36511_36811 , \36512_36812 , \36513_36813 , \36514_36814 , \36515_36815 , \36516_36816 ,
         \36517_36817 , \36518_36818 , \36519_36819 , \36520_36820 , \36521_36821 , \36522_36822 , \36523_36823 , \36524_36824 , \36525_36825 , \36526_36826 ,
         \36527_36827 , \36528_36828 , \36529_36829 , \36530_36830 , \36531_36831 , \36532_36832 , \36533_36833 , \36534_36834 , \36535_36835 , \36536_36836 ,
         \36537_36837 , \36538_36838 , \36539_36839 , \36540_36840 , \36541_36841 , \36542_36842 , \36543_36843 , \36544_36844 , \36545_36845 , \36546_36846 ,
         \36547_36847 , \36548_36848 , \36549_36849 , \36550_36850 , \36551_36851 , \36552_36852 , \36553_36853 , \36554_36854 , \36555_36855 , \36556_36856 ,
         \36557_36857 , \36558_36858 , \36559_36859 , \36560_36860 , \36561_36861 , \36562_36862 , \36563_36863 , \36564_36864 , \36565_36865 , \36566_36866 ,
         \36567_36867 , \36568_36868 , \36569_36869 , \36570_36870 , \36571_36871 , \36572_36872 , \36573_36873 , \36574_36874 , \36575_36875 , \36576_36876 ,
         \36577_36877 , \36578_36878 , \36579_36879 , \36580_36880 , \36581_36881 , \36582_36882 , \36583_36883 , \36584_36884 , \36585_36885 , \36586_36886 ,
         \36587_36887 , \36588_36888 , \36589_36889 , \36590_36890 , \36591_36891 , \36592_36892 , \36593_36893 , \36594_36894 , \36595_36895 , \36596_36896 ,
         \36597_36897 , \36598_36898 , \36599_36899 , \36600_36900 , \36601_36901 , \36602_36902 , \36603_36903 , \36604_36904 , \36605_36905 , \36606_36906 ,
         \36607_36907 , \36608_36908 , \36609_36909 , \36610_36910 , \36611_36911 , \36612_36912 , \36613_36913 , \36614_36914 , \36615_36915 , \36616_36916 ,
         \36617_36917 , \36618_36918 , \36619_36919 , \36620_36920 , \36621_36921 , \36622_36922 , \36623_36923 , \36624_36924 , \36625_36925 , \36626_36926 ,
         \36627_36927 , \36628_36928 , \36629_36929 , \36630_36930 , \36631_36931 , \36632_36932 , \36633_36933 , \36634_36934 , \36635_36935 , \36636_36936 ,
         \36637_36937 , \36638_36938 , \36639_36939 , \36640_36940 , \36641_36941 , \36642_36942 , \36643_36943 , \36644_36944 , \36645_36945 , \36646_36946 ,
         \36647_36947 , \36648_36948 , \36649_36949 , \36650_36950 , \36651_36951 , \36652_36952 , \36653_36953 , \36654_36954 , \36655_36955 , \36656_36956 ,
         \36657_36957 , \36658_36958 , \36659_36959 , \36660_36960 , \36661_36961 , \36662_36962 , \36663_36963 , \36664_36964 , \36665_36965 , \36666_36966 ,
         \36667_36967 , \36668_36968 , \36669_36969 , \36670_36970 , \36671_36971 , \36672_36972 , \36673_36973 , \36674_36974 , \36675_36975 , \36676_36976 ,
         \36677_36977 , \36678_36978 , \36679_36979 , \36680_36980 , \36681_36981 , \36682_36982 , \36683_36983 , \36684_36984 , \36685_36985 , \36686_36986_nG9b90 ,
         \36687_36987 , \36688_36988 , \36689_36989 , \36690_36990 , \36691_36991 , \36692_36992 , \36693_36993 , \36694_36994 , \36695_36995 , \36696_36996 ,
         \36697_36997 , \36698_36998 , \36699_36999 , \36700_37000 , \36701_37001 , \36702_37002 , \36703_37003 , \36704_37004 , \36705_37005 , \36706_37006 ,
         \36707_37007 , \36708_37008 , \36709_37009 , \36710_37010 , \36711_37011 , \36712_37012 , \36713_37013 , \36714_37014 , \36715_37015 , \36716_37016 ,
         \36717_37017 , \36718_37018 , \36719_37019 , \36720_37020 , \36721_37021 , \36722_37022 , \36723_37023 , \36724_37024 , \36725_37025 , \36726_37026 ,
         \36727_37027 , \36728_37028 , \36729_37029 , \36730_37030 , \36731_37031 , \36732_37032 , \36733_37033 , \36734_37034 , \36735_37035 , \36736_37036 ,
         \36737_37037 , \36738_37038 , \36739_37039 , \36740_37040 , \36741_37041 , \36742_37042 , \36743_37043 , \36744_37044 , \36745_37045 , \36746_37046 ,
         \36747_37047 , \36748_37048 , \36749_37049 , \36750_37050 , \36751_37051 , \36752_37052 , \36753_37053 , \36754_37054 , \36755_37055 , \36756_37056 ,
         \36757_37057 , \36758_37058 , \36759_37059 , \36760_37060 , \36761_37061 , \36762_37062 , \36763_37063 , \36764_37064 , \36765_37065 , \36766_37066 ,
         \36767_37067 , \36768_37068 , \36769_37069 , \36770_37070 , \36771_37071 , \36772_37072 , \36773_37073 , \36774_37074 , \36775_37075 , \36776_37076 ,
         \36777_37077 , \36778_37078 , \36779_37079 , \36780_37080 , \36781_37081 , \36782_37082 , \36783_37083 , \36784_37084 , \36785_37085 , \36786_37086 ,
         \36787_37087 , \36788_37088 , \36789_37089 , \36790_37090 , \36791_37091 , \36792_37092 , \36793_37093 , \36794_37094 , \36795_37095 , \36796_37096 ,
         \36797_37097 , \36798_37098 , \36799_37099 , \36800_37100 , \36801_37101 , \36802_37102 , \36803_37103 , \36804_37104 , \36805_37105 , \36806_37106 ,
         \36807_37107 , \36808_37108 , \36809_37109 , \36810_37110 , \36811_37111 , \36812_37112 , \36813_37113 , \36814_37114 , \36815_37115 , \36816_37116 ,
         \36817_37117 , \36818_37118 , \36819_37119 , \36820_37120 , \36821_37121 , \36822_37122 , \36823_37123 , \36824_37124 , \36825_37125 , \36826_37126 ,
         \36827_37127 , \36828_37128 , \36829_37129 , \36830_37130 , \36831_37131 , \36832_37132 , \36833_37133 , \36834_37134 , \36835_37135 , \36836_37136 ,
         \36837_37137 , \36838_37138 , \36839_37139 , \36840_37140 , \36841_37141 , \36842_37142 , \36843_37143 , \36844_37144 , \36845_37145 , \36846_37146 ,
         \36847_37147 , \36848_37148 , \36849_37149 , \36850_37150 , \36851_37151 , \36852_37152 , \36853_37153 , \36854_37154 , \36855_37155 , \36856_37156 ,
         \36857_37157 , \36858_37158 , \36859_37159 , \36860_37160 , \36861_37161 , \36862_37162 , \36863_37163 , \36864_37164 , \36865_37165 , \36866_37166 ,
         \36867_37167 , \36868_37168 , \36869_37169 , \36870_37170 , \36871_37171 , \36872_37172 , \36873_37173 , \36874_37174 , \36875_37175 , \36876_37176 ,
         \36877_37177 , \36878_37178 , \36879_37179 , \36880_37180 , \36881_37181 , \36882_37182 , \36883_37183 , \36884_37184 , \36885_37185 , \36886_37186 ,
         \36887_37187 , \36888_37188 , \36889_37189 , \36890_37190 , \36891_37191 , \36892_37192 , \36893_37193 , \36894_37194 , \36895_37195 , \36896_37196 ,
         \36897_37197 , \36898_37198 , \36899_37199 , \36900_37200 , \36901_37201 , \36902_37202 , \36903_37203 , \36904_37204 , \36905_37205 , \36906_37206 ,
         \36907_37207 , \36908_37208 , \36909_37209 , \36910_37210 , \36911_37211 , \36912_37212 , \36913_37213 , \36914_37214 , \36915_37215 , \36916_37216 ,
         \36917_37217 , \36918_37218 , \36919_37219 , \36920_37220 , \36921_37221 , \36922_37222 , \36923_37223 , \36924_37224 , \36925_37225 , \36926_37226 ,
         \36927_37227 , \36928_37228 , \36929_37229 , \36930_37230 , \36931_37231 , \36932_37232 , \36933_37233 , \36934_37234 , \36935_37235 , \36936_37236 ,
         \36937_37237 , \36938_37238 , \36939_37239 , \36940_37240 , \36941_37241 , \36942_37242 , \36943_37243 , \36944_37244 , \36945_37245 , \36946_37246 ,
         \36947_37247 , \36948_37248 , \36949_37249 , \36950_37250_nG9b8d , \36951_37251 , \36952_37252 , \36953_37253 , \36954_37254 , \36955_37255 , \36956_37256 ,
         \36957_37257 , \36958_37258 , \36959_37259 , \36960_37260 , \36961_37261 , \36962_37262 , \36963_37263 , \36964_37264 , \36965_37265 , \36966_37266 ,
         \36967_37267 , \36968_37268 , \36969_37269 , \36970_37270 , \36971_37271 , \36972_37272 , \36973_37273 , \36974_37274 , \36975_37275 , \36976_37276 ,
         \36977_37277 , \36978_37278 , \36979_37279 , \36980_37280 , \36981_37281 , \36982_37282 , \36983_37283 , \36984_37284 , \36985_37285 , \36986_37286 ,
         \36987_37287 , \36988_37288 , \36989_37289 , \36990_37290 , \36991_37291 , \36992_37292 , \36993_37293 , \36994_37294 , \36995_37295 , \36996_37296 ,
         \36997_37297 , \36998_37298 , \36999_37299 , \37000_37300 , \37001_37301 , \37002_37302 , \37003_37303 , \37004_37304 , \37005_37305 , \37006_37306 ,
         \37007_37307 , \37008_37308 , \37009_37309 , \37010_37310 , \37011_37311 , \37012_37312 , \37013_37313 , \37014_37314 , \37015_37315 , \37016_37316 ,
         \37017_37317 , \37018_37318 , \37019_37319 , \37020_37320 , \37021_37321 , \37022_37322 , \37023_37323 , \37024_37324 , \37025_37325 , \37026_37326 ,
         \37027_37327 , \37028_37328 , \37029_37329 , \37030_37330 , \37031_37331 , \37032_37332 , \37033_37333 , \37034_37334 , \37035_37335 , \37036_37336 ,
         \37037_37337 , \37038_37338 , \37039_37339 , \37040_37340 , \37041_37341 , \37042_37342 , \37043_37343 , \37044_37344 , \37045_37345 , \37046_37346 ,
         \37047_37347 , \37048_37348 , \37049_37349 , \37050_37350 , \37051_37351 , \37052_37352 , \37053_37353 , \37054_37354 , \37055_37355 , \37056_37356 ,
         \37057_37357 , \37058_37358 , \37059_37359 , \37060_37360 , \37061_37361 , \37062_37362 , \37063_37363 , \37064_37364 , \37065_37365 , \37066_37366 ,
         \37067_37367 , \37068_37368 , \37069_37369 , \37070_37370 , \37071_37371 , \37072_37372 , \37073_37373 , \37074_37374 , \37075_37375 , \37076_37376 ,
         \37077_37377 , \37078_37378 , \37079_37379 , \37080_37380 , \37081_37381 , \37082_37382 , \37083_37383 , \37084_37384 , \37085_37385 , \37086_37386 ,
         \37087_37387 , \37088_37388 , \37089_37389 , \37090_37390 , \37091_37391 , \37092_37392 , \37093_37393 , \37094_37394 , \37095_37395 , \37096_37396 ,
         \37097_37397 , \37098_37398 , \37099_37399 , \37100_37400 , \37101_37401 , \37102_37402 , \37103_37403 , \37104_37404 , \37105_37405 , \37106_37406 ,
         \37107_37407 , \37108_37408 , \37109_37409 , \37110_37410 , \37111_37411 , \37112_37412 , \37113_37413 , \37114_37414 , \37115_37415 , \37116_37416 ,
         \37117_37417 , \37118_37418 , \37119_37419 , \37120_37420 , \37121_37421 , \37122_37422 , \37123_37423 , \37124_37424 , \37125_37425 , \37126_37426 ,
         \37127_37427 , \37128_37428 , \37129_37429 , \37130_37430 , \37131_37431 , \37132_37432 , \37133_37433 , \37134_37434 , \37135_37435 , \37136_37436 ,
         \37137_37437 , \37138_37438 , \37139_37439 , \37140_37440 , \37141_37441 , \37142_37442 , \37143_37443 , \37144_37444 , \37145_37445 , \37146_37446 ,
         \37147_37447 , \37148_37448 , \37149_37449 , \37150_37450 , \37151_37451 , \37152_37452 , \37153_37453 , \37154_37454 , \37155_37455 , \37156_37456 ,
         \37157_37457 , \37158_37458 , \37159_37459 , \37160_37460 , \37161_37461 , \37162_37462 , \37163_37463 , \37164_37464 , \37165_37465 , \37166_37466 ,
         \37167_37467 , \37168_37468 , \37169_37469 , \37170_37470 , \37171_37471 , \37172_37472 , \37173_37473 , \37174_37474 , \37175_37475 , \37176_37476 ,
         \37177_37477 , \37178_37478 , \37179_37479 , \37180_37480 , \37181_37481 , \37182_37482 , \37183_37483 , \37184_37484 , \37185_37485 , \37186_37486 ,
         \37187_37487 , \37188_37488 , \37189_37489 , \37190_37490 , \37191_37491 , \37192_37492 , \37193_37493 , \37194_37494 , \37195_37495 , \37196_37496 ,
         \37197_37497 , \37198_37498 , \37199_37499 , \37200_37500 , \37201_37501 , \37202_37502 , \37203_37503 , \37204_37504 , \37205_37505 , \37206_37506 ,
         \37207_37507 , \37208_37508 , \37209_37509 , \37210_37510 , \37211_37511 , \37212_37512 , \37213_37513 , \37214_37514 , \37215_37515 , \37216_37516 ,
         \37217_37517 , \37218_37518 , \37219_37519 , \37220_37520 , \37221_37521 , \37222_37522 , \37223_37523 , \37224_37524 , \37225_37525 , \37226_37526 ,
         \37227_37527 , \37228_37528 , \37229_37529 , \37230_37530 , \37231_37531 , \37232_37532 , \37233_37533 , \37234_37534 , \37235_37535 , \37236_37536 ,
         \37237_37537 , \37238_37538 , \37239_37539 , \37240_37540 , \37241_37541 , \37242_37542 , \37243_37543 , \37244_37544 , \37245_37545 , \37246_37546 ,
         \37247_37547 , \37248_37548 , \37249_37549 , \37250_37550 , \37251_37551 , \37252_37552 , \37253_37553 , \37254_37554 , \37255_37555 , \37256_37556 ,
         \37257_37557 , \37258_37558 , \37259_37559 , \37260_37560 , \37261_37561 , \37262_37562 , \37263_37563 , \37264_37564 , \37265_37565 , \37266_37566 ,
         \37267_37567 , \37268_37568 , \37269_37569 , \37270_37570 , \37271_37571 , \37272_37572 , \37273_37573 , \37274_37574 , \37275_37575 , \37276_37576 ,
         \37277_37577 , \37278_37578 , \37279_37579 , \37280_37580 , \37281_37581 , \37282_37582 , \37283_37583 , \37284_37584 , \37285_37585 , \37286_37586 ,
         \37287_37587 , \37288_37588 , \37289_37589 , \37290_37590 , \37291_37591 , \37292_37592 , \37293_37593 , \37294_37594 , \37295_37595 , \37296_37596 ,
         \37297_37597 , \37298_37598 , \37299_37599 , \37300_37600 , \37301_37601 , \37302_37602 , \37303_37603 , \37304_37604 , \37305_37605 , \37306_37606 ,
         \37307_37607_nG9b8a , \37308_37608 , \37309_37609 , \37310_37610 , \37311_37611 , \37312_37612 , \37313_37613 , \37314_37614 , \37315_37615 , \37316_37616 ,
         \37317_37617 , \37318_37618 , \37319_37619 , \37320_37620 , \37321_37621 , \37322_37622 , \37323_37623 , \37324_37624 , \37325_37625 , \37326_37626 ,
         \37327_37627 , \37328_37628 , \37329_37629 , \37330_37630 , \37331_37631 , \37332_37632 , \37333_37633 , \37334_37634 , \37335_37635 , \37336_37636 ,
         \37337_37637 , \37338_37638 , \37339_37639 , \37340_37640 , \37341_37641 , \37342_37642 , \37343_37643 , \37344_37644 , \37345_37645 , \37346_37646 ,
         \37347_37647 , \37348_37648 , \37349_37649 , \37350_37650 , \37351_37651 , \37352_37652 , \37353_37653 , \37354_37654 , \37355_37655 , \37356_37656 ,
         \37357_37657 , \37358_37658 , \37359_37659 , \37360_37660 , \37361_37661 , \37362_37662 , \37363_37663 , \37364_37664 , \37365_37665 , \37366_37666 ,
         \37367_37667 , \37368_37668 , \37369_37669 , \37370_37670 , \37371_37671 , \37372_37672 , \37373_37673 , \37374_37674 , \37375_37675 , \37376_37676 ,
         \37377_37677 , \37378_37678 , \37379_37679 , \37380_37680 , \37381_37681 , \37382_37682 , \37383_37683 , \37384_37684 , \37385_37685 , \37386_37686 ,
         \37387_37687 , \37388_37688 , \37389_37689 , \37390_37690 , \37391_37691 , \37392_37692 , \37393_37693 , \37394_37694 , \37395_37695 , \37396_37696 ,
         \37397_37697 , \37398_37698 , \37399_37699 , \37400_37700 , \37401_37701 , \37402_37702 , \37403_37703 , \37404_37704 , \37405_37705 , \37406_37706 ,
         \37407_37707 , \37408_37708 , \37409_37709 , \37410_37710 , \37411_37711 , \37412_37712 , \37413_37713 , \37414_37714 , \37415_37715 , \37416_37716 ,
         \37417_37717 , \37418_37718 , \37419_37719 , \37420_37720 , \37421_37721 , \37422_37722 , \37423_37723 , \37424_37724 , \37425_37725 , \37426_37726 ,
         \37427_37727 , \37428_37728 , \37429_37729 , \37430_37730 , \37431_37731 , \37432_37732 , \37433_37733 , \37434_37734 , \37435_37735 , \37436_37736 ,
         \37437_37737 , \37438_37738 , \37439_37739 , \37440_37740 , \37441_37741 , \37442_37742 , \37443_37743 , \37444_37744 , \37445_37745 , \37446_37746 ,
         \37447_37747 , \37448_37748 , \37449_37749 , \37450_37750 , \37451_37751 , \37452_37752 , \37453_37753 , \37454_37754 , \37455_37755 , \37456_37756 ,
         \37457_37757 , \37458_37758 , \37459_37759 , \37460_37760 , \37461_37761 , \37462_37762 , \37463_37763 , \37464_37764 , \37465_37765 , \37466_37766 ,
         \37467_37767 , \37468_37768 , \37469_37769 , \37470_37770 , \37471_37771 , \37472_37772 , \37473_37773 , \37474_37774 , \37475_37775 , \37476_37776 ,
         \37477_37777 , \37478_37778 , \37479_37779 , \37480_37780 , \37481_37781 , \37482_37782 , \37483_37783 , \37484_37784 , \37485_37785 , \37486_37786 ,
         \37487_37787 , \37488_37788 , \37489_37789 , \37490_37790 , \37491_37791 , \37492_37792 , \37493_37793 , \37494_37794 , \37495_37795 , \37496_37796 ,
         \37497_37797 , \37498_37798 , \37499_37799 , \37500_37800 , \37501_37801 , \37502_37802 , \37503_37803 , \37504_37804 , \37505_37805 , \37506_37806 ,
         \37507_37807 , \37508_37808 , \37509_37809 , \37510_37810 , \37511_37811 , \37512_37812 , \37513_37813 , \37514_37814 , \37515_37815 , \37516_37816 ,
         \37517_37817 , \37518_37818 , \37519_37819 , \37520_37820 , \37521_37821 , \37522_37822 , \37523_37823 , \37524_37824 , \37525_37825 , \37526_37826 ,
         \37527_37827 , \37528_37828 , \37529_37829 , \37530_37830 , \37531_37831 , \37532_37832 , \37533_37833 , \37534_37834 , \37535_37835 , \37536_37836 ,
         \37537_37837 , \37538_37838 , \37539_37839 , \37540_37840 , \37541_37841 , \37542_37842 , \37543_37843 , \37544_37844 , \37545_37845 , \37546_37846 ,
         \37547_37847 , \37548_37848 , \37549_37849 , \37550_37850 , \37551_37851 , \37552_37852 , \37553_37853 , \37554_37854 , \37555_37855 , \37556_37856 ,
         \37557_37857 , \37558_37858 , \37559_37859 , \37560_37860 , \37561_37861 , \37562_37862 , \37563_37863 , \37564_37864 , \37565_37865 , \37566_37866 ,
         \37567_37867 , \37568_37868 , \37569_37869 , \37570_37870 , \37571_37871 , \37572_37872 , \37573_37873 , \37574_37874 , \37575_37875 , \37576_37876 ,
         \37577_37877 , \37578_37878 , \37579_37879 , \37580_37880 , \37581_37881 , \37582_37882 , \37583_37883 , \37584_37884 , \37585_37885 , \37586_37886 ,
         \37587_37887 , \37588_37888 , \37589_37889 , \37590_37890 , \37591_37891 , \37592_37892 , \37593_37893 , \37594_37894 , \37595_37895 , \37596_37896 ,
         \37597_37897 , \37598_37898 , \37599_37899 , \37600_37900 , \37601_37901 , \37602_37902 , \37603_37903 , \37604_37904 , \37605_37905 , \37606_37906 ,
         \37607_37907 , \37608_37908 , \37609_37909 , \37610_37910 , \37611_37911 , \37612_37912 , \37613_37913 , \37614_37914 , \37615_37915 , \37616_37916 ,
         \37617_37917 , \37618_37918 , \37619_37919 , \37620_37920 , \37621_37921 , \37622_37922 , \37623_37923 , \37624_37924 , \37625_37925 , \37626_37926 ,
         \37627_37927 , \37628_37928 , \37629_37929 , \37630_37930 , \37631_37931 , \37632_37932 , \37633_37933 , \37634_37934 , \37635_37935 , \37636_37936 ,
         \37637_37937 , \37638_37938 , \37639_37939 , \37640_37940 , \37641_37941 , \37642_37942 , \37643_37943 , \37644_37944 , \37645_37945 , \37646_37946 ,
         \37647_37947 , \37648_37948 , \37649_37949 , \37650_37950 , \37651_37951 , \37652_37952 , \37653_37953 , \37654_37954 , \37655_37955 , \37656_37956 ,
         \37657_37957 , \37658_37958 , \37659_37959 , \37660_37960 , \37661_37961 , \37662_37962 , \37663_37963 , \37664_37964 , \37665_37965 , \37666_37966 ,
         \37667_37967 , \37668_37968 , \37669_37969 , \37670_37970 , \37671_37971 , \37672_37972 , \37673_37973 , \37674_37974_nG9b87 , \37675_37975 , \37676_37976 ,
         \37677_37977 , \37678_37978 , \37679_37979 , \37680_37980 , \37681_37981 , \37682_37982 , \37683_37983 , \37684_37984 , \37685_37985 , \37686_37986 ,
         \37687_37987 , \37688_37988 , \37689_37989 , \37690_37990 , \37691_37991 , \37692_37992 , \37693_37993 , \37694_37994 , \37695_37995 , \37696_37996 ,
         \37697_37997 , \37698_37998 , \37699_37999 , \37700_38000 , \37701_38001 , \37702_38002 , \37703_38003 , \37704_38004 , \37705_38005 , \37706_38006 ,
         \37707_38007 , \37708_38008 , \37709_38009 , \37710_38010 , \37711_38011 , \37712_38012 , \37713_38013 , \37714_38014 , \37715_38015 , \37716_38016 ,
         \37717_38017 , \37718_38018 , \37719_38019 , \37720_38020 , \37721_38021 , \37722_38022 , \37723_38023 , \37724_38024 , \37725_38025 , \37726_38026 ,
         \37727_38027 , \37728_38028 , \37729_38029 , \37730_38030 , \37731_38031 , \37732_38032 , \37733_38033 , \37734_38034 , \37735_38035 , \37736_38036 ,
         \37737_38037 , \37738_38038 , \37739_38039 , \37740_38040 , \37741_38041 , \37742_38042 , \37743_38043 , \37744_38044 , \37745_38045 , \37746_38046 ,
         \37747_38047 , \37748_38048 , \37749_38049 , \37750_38050 , \37751_38051 , \37752_38052 , \37753_38053 , \37754_38054 , \37755_38055 , \37756_38056 ,
         \37757_38057 , \37758_38058 , \37759_38059 , \37760_38060 , \37761_38061 , \37762_38062 , \37763_38063 , \37764_38064 , \37765_38065 , \37766_38066 ,
         \37767_38067 , \37768_38068 , \37769_38069 , \37770_38070 , \37771_38071 , \37772_38072 , \37773_38073 , \37774_38074 , \37775_38075 , \37776_38076 ,
         \37777_38077 , \37778_38078 , \37779_38079 , \37780_38080 , \37781_38081 , \37782_38082 , \37783_38083 , \37784_38084 , \37785_38085 , \37786_38086 ,
         \37787_38087 , \37788_38088 , \37789_38089 , \37790_38090 , \37791_38091 , \37792_38092 , \37793_38093 , \37794_38094 , \37795_38095 , \37796_38096 ,
         \37797_38097 , \37798_38098 , \37799_38099 , \37800_38100 , \37801_38101 , \37802_38102 , \37803_38103 , \37804_38104 , \37805_38105 , \37806_38106 ,
         \37807_38107 , \37808_38108 , \37809_38109 , \37810_38110 , \37811_38111 , \37812_38112 , \37813_38113 , \37814_38114 , \37815_38115 , \37816_38116 ,
         \37817_38117 , \37818_38118 , \37819_38119 , \37820_38120 , \37821_38121 , \37822_38122 , \37823_38123 , \37824_38124 , \37825_38125 , \37826_38126 ,
         \37827_38127 , \37828_38128 , \37829_38129 , \37830_38130 , \37831_38131 , \37832_38132 , \37833_38133 , \37834_38134 , \37835_38135 , \37836_38136 ,
         \37837_38137 , \37838_38138 , \37839_38139 , \37840_38140 , \37841_38141 , \37842_38142 , \37843_38143 , \37844_38144 , \37845_38145 , \37846_38146 ,
         \37847_38147 , \37848_38148 , \37849_38149 , \37850_38150 , \37851_38151 , \37852_38152 , \37853_38153 , \37854_38154 , \37855_38155 , \37856_38156 ,
         \37857_38157 , \37858_38158 , \37859_38159 , \37860_38160 , \37861_38161 , \37862_38162 , \37863_38163 , \37864_38164 , \37865_38165 , \37866_38166 ,
         \37867_38167 , \37868_38168 , \37869_38169 , \37870_38170 , \37871_38171 , \37872_38172 , \37873_38173 , \37874_38174 , \37875_38175 , \37876_38176 ,
         \37877_38177 , \37878_38178 , \37879_38179 , \37880_38180 , \37881_38181 , \37882_38182 , \37883_38183 , \37884_38184 , \37885_38185 , \37886_38186 ,
         \37887_38187 , \37888_38188 , \37889_38189 , \37890_38190 , \37891_38191 , \37892_38192 , \37893_38193 , \37894_38194 , \37895_38195 , \37896_38196 ,
         \37897_38197 , \37898_38198 , \37899_38199 , \37900_38200 , \37901_38201 , \37902_38202 , \37903_38203 , \37904_38204 , \37905_38205 , \37906_38206 ,
         \37907_38207 , \37908_38208 , \37909_38209 , \37910_38210 , \37911_38211 , \37912_38212 , \37913_38213 , \37914_38214 , \37915_38215 , \37916_38216 ,
         \37917_38217 , \37918_38218 , \37919_38219 , \37920_38220 , \37921_38221 , \37922_38222 , \37923_38223 , \37924_38224 , \37925_38225 , \37926_38226 ,
         \37927_38227 , \37928_38228 , \37929_38229 , \37930_38230 , \37931_38231 , \37932_38232 , \37933_38233 , \37934_38234 , \37935_38235 , \37936_38236 ,
         \37937_38237 , \37938_38238 , \37939_38239 , \37940_38240 , \37941_38241 , \37942_38242 , \37943_38243 , \37944_38244 , \37945_38245 , \37946_38246 ,
         \37947_38247 , \37948_38248 , \37949_38249 , \37950_38250 , \37951_38251 , \37952_38252 , \37953_38253 , \37954_38254 , \37955_38255 , \37956_38256 ,
         \37957_38257 , \37958_38258 , \37959_38259 , \37960_38260 , \37961_38261 , \37962_38262 , \37963_38263 , \37964_38264 , \37965_38265 , \37966_38266 ,
         \37967_38267 , \37968_38268 , \37969_38269 , \37970_38270 , \37971_38271 , \37972_38272 , \37973_38273 , \37974_38274 , \37975_38275 , \37976_38276 ,
         \37977_38277 , \37978_38278 , \37979_38279 , \37980_38280 , \37981_38281 , \37982_38282 , \37983_38283 , \37984_38284 , \37985_38285 , \37986_38286 ,
         \37987_38287 , \37988_38288 , \37989_38289 , \37990_38290 , \37991_38291 , \37992_38292 , \37993_38293 , \37994_38294 , \37995_38295 , \37996_38296 ,
         \37997_38297 , \37998_38298 , \37999_38299 , \38000_38300 , \38001_38301 , \38002_38302 , \38003_38303 , \38004_38304 , \38005_38305 , \38006_38306 ,
         \38007_38307 , \38008_38308 , \38009_38309 , \38010_38310 , \38011_38311 , \38012_38312 , \38013_38313 , \38014_38314 , \38015_38315 , \38016_38316 ,
         \38017_38317 , \38018_38318 , \38019_38319 , \38020_38320 , \38021_38321 , \38022_38322 , \38023_38323 , \38024_38324 , \38025_38325 , \38026_38326 ,
         \38027_38327 , \38028_38328 , \38029_38329 , \38030_38330 , \38031_38331 , \38032_38332 , \38033_38333 , \38034_38334 , \38035_38335 , \38036_38336 ,
         \38037_38337_nG9b84 , \38038_38338 , \38039_38339 , \38040_38340 , \38041_38341 , \38042_38342 , \38043_38343 , \38044_38344 , \38045_38345 , \38046_38346 ,
         \38047_38347 , \38048_38348 , \38049_38349 , \38050_38350 , \38051_38351 , \38052_38352 , \38053_38353 , \38054_38354 , \38055_38355 , \38056_38356 ,
         \38057_38357 , \38058_38358 , \38059_38359 , \38060_38360 , \38061_38361 , \38062_38362 , \38063_38363 , \38064_38364 , \38065_38365 , \38066_38366 ,
         \38067_38367 , \38068_38368 , \38069_38369 , \38070_38370 , \38071_38371 , \38072_38372 , \38073_38373 , \38074_38374 , \38075_38375 , \38076_38376 ,
         \38077_38377 , \38078_38378 , \38079_38379 , \38080_38380 , \38081_38381 , \38082_38382 , \38083_38383 , \38084_38384 , \38085_38385 , \38086_38386 ,
         \38087_38387 , \38088_38388 , \38089_38389 , \38090_38390 , \38091_38391 , \38092_38392 , \38093_38393 , \38094_38394 , \38095_38395 , \38096_38396 ,
         \38097_38397 , \38098_38398 , \38099_38399 , \38100_38400 , \38101_38401 , \38102_38402 , \38103_38403 , \38104_38404 , \38105_38405 , \38106_38406 ,
         \38107_38407 , \38108_38408 , \38109_38409 , \38110_38410 , \38111_38411 , \38112_38412 , \38113_38413 , \38114_38414 , \38115_38415 , \38116_38416 ,
         \38117_38417 , \38118_38418 , \38119_38419 , \38120_38420 , \38121_38421 , \38122_38422 , \38123_38423 , \38124_38424 , \38125_38425 , \38126_38426 ,
         \38127_38427 , \38128_38428 , \38129_38429 , \38130_38430 , \38131_38431 , \38132_38432 , \38133_38433 , \38134_38434 , \38135_38435 , \38136_38436 ,
         \38137_38437 , \38138_38438 , \38139_38439 , \38140_38440 , \38141_38441 , \38142_38442 , \38143_38443 , \38144_38444 , \38145_38445 , \38146_38446 ,
         \38147_38447 , \38148_38448 , \38149_38449 , \38150_38450 , \38151_38451 , \38152_38452 , \38153_38453 , \38154_38454 , \38155_38455 , \38156_38456 ,
         \38157_38457 , \38158_38458 , \38159_38459 , \38160_38460 , \38161_38461 , \38162_38462 , \38163_38463 , \38164_38464 , \38165_38465 , \38166_38466 ,
         \38167_38467 , \38168_38468 , \38169_38469 , \38170_38470 , \38171_38471 , \38172_38472 , \38173_38473 , \38174_38474 , \38175_38475 , \38176_38476 ,
         \38177_38477 , \38178_38478 , \38179_38479 , \38180_38480 , \38181_38481 , \38182_38482 , \38183_38483 , \38184_38484 , \38185_38485 , \38186_38486 ,
         \38187_38487 , \38188_38488 , \38189_38489 , \38190_38490 , \38191_38491 , \38192_38492 , \38193_38493 , \38194_38494 , \38195_38495 , \38196_38496 ,
         \38197_38497 , \38198_38498 , \38199_38499 , \38200_38500 , \38201_38501 , \38202_38502 , \38203_38503 , \38204_38504 , \38205_38505 , \38206_38506 ,
         \38207_38507 , \38208_38508 , \38209_38509 , \38210_38510 , \38211_38511 , \38212_38512 , \38213_38513 , \38214_38514 , \38215_38515 , \38216_38516 ,
         \38217_38517 , \38218_38518 , \38219_38519 , \38220_38520 , \38221_38521 , \38222_38522 , \38223_38523 , \38224_38524 , \38225_38525 , \38226_38526 ,
         \38227_38527 , \38228_38528 , \38229_38529 , \38230_38530 , \38231_38531 , \38232_38532 , \38233_38533 , \38234_38534 , \38235_38535 , \38236_38536 ,
         \38237_38537 , \38238_38538 , \38239_38539 , \38240_38540 , \38241_38541 , \38242_38542 , \38243_38543 , \38244_38544 , \38245_38545 , \38246_38546 ,
         \38247_38547 , \38248_38548 , \38249_38549 , \38250_38550 , \38251_38551 , \38252_38552 , \38253_38553 , \38254_38554 , \38255_38555 , \38256_38556 ,
         \38257_38557 , \38258_38558 , \38259_38559 , \38260_38560 , \38261_38561 , \38262_38562 , \38263_38563 , \38264_38564 , \38265_38565 , \38266_38566 ,
         \38267_38567 , \38268_38568 , \38269_38569 , \38270_38570 , \38271_38571 , \38272_38572 , \38273_38573 , \38274_38574 , \38275_38575 , \38276_38576 ,
         \38277_38577 , \38278_38578 , \38279_38579 , \38280_38580 , \38281_38581 , \38282_38582 , \38283_38583 , \38284_38584 , \38285_38585 , \38286_38586 ,
         \38287_38587 , \38288_38588 , \38289_38589 , \38290_38590 , \38291_38591 , \38292_38592 , \38293_38593 , \38294_38594 , \38295_38595 , \38296_38596 ,
         \38297_38597 , \38298_38598 , \38299_38599 , \38300_38600 , \38301_38601 , \38302_38602 , \38303_38603 , \38304_38604 , \38305_38605 , \38306_38606 ,
         \38307_38607 , \38308_38608 , \38309_38609 , \38310_38610 , \38311_38611 , \38312_38612 , \38313_38613 , \38314_38614 , \38315_38615 , \38316_38616 ,
         \38317_38617 , \38318_38618 , \38319_38619 , \38320_38620 , \38321_38621 , \38322_38622 , \38323_38623 , \38324_38624 , \38325_38625 , \38326_38626 ,
         \38327_38627 , \38328_38628 , \38329_38629 , \38330_38630 , \38331_38631 , \38332_38632 , \38333_38633 , \38334_38634 , \38335_38635 , \38336_38636 ,
         \38337_38637 , \38338_38638 , \38339_38639 , \38340_38640 , \38341_38641 , \38342_38642 , \38343_38643 , \38344_38644 , \38345_38645 , \38346_38646 ,
         \38347_38647 , \38348_38648 , \38349_38649 , \38350_38650 , \38351_38651 , \38352_38652 , \38353_38653 , \38354_38654 , \38355_38655 , \38356_38656 ,
         \38357_38657 , \38358_38658 , \38359_38659 , \38360_38660 , \38361_38661 , \38362_38662 , \38363_38663_nG9b81 , \38364_38664 , \38365_38665 , \38366_38666 ,
         \38367_38667 , \38368_38668 , \38369_38669 , \38370_38670 , \38371_38671 , \38372_38672 , \38373_38673 , \38374_38674 , \38375_38675 , \38376_38676 ,
         \38377_38677 , \38378_38678 , \38379_38679 , \38380_38680 , \38381_38681 , \38382_38682 , \38383_38683 , \38384_38684 , \38385_38685 , \38386_38686 ,
         \38387_38687 , \38388_38688 , \38389_38689 , \38390_38690 , \38391_38691 , \38392_38692 , \38393_38693 , \38394_38694 , \38395_38695 , \38396_38696 ,
         \38397_38697 , \38398_38698 , \38399_38699 , \38400_38700 , \38401_38701 , \38402_38702 , \38403_38703 , \38404_38704 , \38405_38705 , \38406_38706 ,
         \38407_38707 , \38408_38708 , \38409_38709 , \38410_38710 , \38411_38711 , \38412_38712 , \38413_38713 , \38414_38714 , \38415_38715 , \38416_38716 ,
         \38417_38717 , \38418_38718 , \38419_38719 , \38420_38720 , \38421_38721 , \38422_38722 , \38423_38723 , \38424_38724 , \38425_38725 , \38426_38726 ,
         \38427_38727 , \38428_38728 , \38429_38729 , \38430_38730 , \38431_38731 , \38432_38732 , \38433_38733 , \38434_38734 , \38435_38735 , \38436_38736 ,
         \38437_38737 , \38438_38738 , \38439_38739 , \38440_38740 , \38441_38741 , \38442_38742 , \38443_38743 , \38444_38744 , \38445_38745 , \38446_38746 ,
         \38447_38747 , \38448_38748 , \38449_38749 , \38450_38750 , \38451_38751 , \38452_38752 , \38453_38753 , \38454_38754 , \38455_38755 , \38456_38756 ,
         \38457_38757 , \38458_38758 , \38459_38759 , \38460_38760 , \38461_38761 , \38462_38762 , \38463_38763 , \38464_38764 , \38465_38765 , \38466_38766 ,
         \38467_38767 , \38468_38768 , \38469_38769 , \38470_38770 , \38471_38771 , \38472_38772 , \38473_38773 , \38474_38774 , \38475_38775 , \38476_38776 ,
         \38477_38777 , \38478_38778 , \38479_38779 , \38480_38780 , \38481_38781 , \38482_38782 , \38483_38783 , \38484_38784 , \38485_38785 , \38486_38786 ,
         \38487_38787 , \38488_38788 , \38489_38789 , \38490_38790 , \38491_38791 , \38492_38792 , \38493_38793 , \38494_38794 , \38495_38795 , \38496_38796 ,
         \38497_38797 , \38498_38798 , \38499_38799 , \38500_38800 , \38501_38801 , \38502_38802 , \38503_38803 , \38504_38804 , \38505_38805 , \38506_38806 ,
         \38507_38807 , \38508_38808 , \38509_38809 , \38510_38810 , \38511_38811 , \38512_38812 , \38513_38813 , \38514_38814 , \38515_38815 , \38516_38816 ,
         \38517_38817 , \38518_38818 , \38519_38819 , \38520_38820 , \38521_38821 , \38522_38822 , \38523_38823 , \38524_38824 , \38525_38825 , \38526_38826 ,
         \38527_38827 , \38528_38828 , \38529_38829 , \38530_38830 , \38531_38831 , \38532_38832 , \38533_38833 , \38534_38834 , \38535_38835 , \38536_38836 ,
         \38537_38837 , \38538_38838 , \38539_38839 , \38540_38840 , \38541_38841 , \38542_38842 , \38543_38843 , \38544_38844 , \38545_38845 , \38546_38846 ,
         \38547_38847 , \38548_38848 , \38549_38849 , \38550_38850 , \38551_38851 , \38552_38852 , \38553_38853 , \38554_38854 , \38555_38855 , \38556_38856 ,
         \38557_38857 , \38558_38858 , \38559_38859 , \38560_38860 , \38561_38861 , \38562_38862 , \38563_38863 , \38564_38864 , \38565_38865 , \38566_38866 ,
         \38567_38867 , \38568_38868 , \38569_38869 , \38570_38870 , \38571_38871 , \38572_38872 , \38573_38873 , \38574_38874 , \38575_38875 , \38576_38876 ,
         \38577_38877 , \38578_38878 , \38579_38879 , \38580_38880 , \38581_38881 , \38582_38882 , \38583_38883 , \38584_38884 , \38585_38885 , \38586_38886 ,
         \38587_38887 , \38588_38888 , \38589_38889 , \38590_38890 , \38591_38891 , \38592_38892 , \38593_38893 , \38594_38894 , \38595_38895 , \38596_38896 ,
         \38597_38897 , \38598_38898 , \38599_38899 , \38600_38900 , \38601_38901 , \38602_38902 , \38603_38903 , \38604_38904 , \38605_38905 , \38606_38906 ,
         \38607_38907 , \38608_38908 , \38609_38909 , \38610_38910 , \38611_38911 , \38612_38912 , \38613_38913 , \38614_38914 , \38615_38915 , \38616_38916 ,
         \38617_38917 , \38618_38918 , \38619_38919 , \38620_38920 , \38621_38921 , \38622_38922 , \38623_38923 , \38624_38924 , \38625_38925 , \38626_38926 ,
         \38627_38927 , \38628_38928 , \38629_38929 , \38630_38930 , \38631_38931 , \38632_38932 , \38633_38933 , \38634_38934 , \38635_38935 , \38636_38936 ,
         \38637_38937 , \38638_38938 , \38639_38939 , \38640_38940 , \38641_38941 , \38642_38942 , \38643_38943 , \38644_38944 , \38645_38945 , \38646_38946 ,
         \38647_38947 , \38648_38948 , \38649_38949 , \38650_38950 , \38651_38951 , \38652_38952 , \38653_38953 , \38654_38954 , \38655_38955 , \38656_38956 ,
         \38657_38957 , \38658_38958 , \38659_38959 , \38660_38960 , \38661_38961 , \38662_38962 , \38663_38963 , \38664_38964 , \38665_38965 , \38666_38966 ,
         \38667_38967 , \38668_38968_nG9b7e , \38669_38969 , \38670_38970 , \38671_38971 , \38672_38972 , \38673_38973 , \38674_38974 , \38675_38975 , \38676_38976 ,
         \38677_38977 , \38678_38978 , \38679_38979 , \38680_38980 , \38681_38981 , \38682_38982 , \38683_38983 , \38684_38984 , \38685_38985 , \38686_38986 ,
         \38687_38987 , \38688_38988 , \38689_38989 , \38690_38990 , \38691_38991 , \38692_38992 , \38693_38993 , \38694_38994 , \38695_38995 , \38696_38996 ,
         \38697_38997 , \38698_38998 , \38699_38999 , \38700_39000 , \38701_39001 , \38702_39002 , \38703_39003 , \38704_39004 , \38705_39005 , \38706_39006 ,
         \38707_39007 , \38708_39008 , \38709_39009 , \38710_39010 , \38711_39011 , \38712_39012 , \38713_39013 , \38714_39014 , \38715_39015 , \38716_39016 ,
         \38717_39017 , \38718_39018 , \38719_39019 , \38720_39020 , \38721_39021 , \38722_39022 , \38723_39023 , \38724_39024 , \38725_39025 , \38726_39026 ,
         \38727_39027 , \38728_39028 , \38729_39029 , \38730_39030 , \38731_39031 , \38732_39032 , \38733_39033 , \38734_39034 , \38735_39035 , \38736_39036 ,
         \38737_39037 , \38738_39038 , \38739_39039 , \38740_39040 , \38741_39041 , \38742_39042 , \38743_39043 , \38744_39044 , \38745_39045 , \38746_39046 ,
         \38747_39047 , \38748_39048 , \38749_39049 , \38750_39050 , \38751_39051 , \38752_39052 , \38753_39053 , \38754_39054 , \38755_39055 , \38756_39056 ,
         \38757_39057 , \38758_39058 , \38759_39059 , \38760_39060 , \38761_39061 , \38762_39062 , \38763_39063 , \38764_39064 , \38765_39065 , \38766_39066 ,
         \38767_39067 , \38768_39068 , \38769_39069 , \38770_39070 , \38771_39071 , \38772_39072 , \38773_39073 , \38774_39074 , \38775_39075 , \38776_39076 ,
         \38777_39077 , \38778_39078 , \38779_39079 , \38780_39080 , \38781_39081 , \38782_39082 , \38783_39083 , \38784_39084 , \38785_39085 , \38786_39086 ,
         \38787_39087 , \38788_39088 , \38789_39089 , \38790_39090 , \38791_39091 , \38792_39092 , \38793_39093 , \38794_39094 , \38795_39095 , \38796_39096 ,
         \38797_39097 , \38798_39098 , \38799_39099 , \38800_39100 , \38801_39101 , \38802_39102 , \38803_39103 , \38804_39104 , \38805_39105 , \38806_39106 ,
         \38807_39107 , \38808_39108 , \38809_39109 , \38810_39110 , \38811_39111 , \38812_39112 , \38813_39113 , \38814_39114 , \38815_39115 , \38816_39116 ,
         \38817_39117 , \38818_39118 , \38819_39119 , \38820_39120 , \38821_39121 , \38822_39122 , \38823_39123 , \38824_39124 , \38825_39125 , \38826_39126 ,
         \38827_39127 , \38828_39128 , \38829_39129 , \38830_39130 , \38831_39131 , \38832_39132 , \38833_39133 , \38834_39134 , \38835_39135 , \38836_39136 ,
         \38837_39137 , \38838_39138 , \38839_39139 , \38840_39140 , \38841_39141 , \38842_39142 , \38843_39143 , \38844_39144 , \38845_39145 , \38846_39146 ,
         \38847_39147 , \38848_39148 , \38849_39149 , \38850_39150 , \38851_39151 , \38852_39152 , \38853_39153 , \38854_39154 , \38855_39155 , \38856_39156 ,
         \38857_39157 , \38858_39158 , \38859_39159 , \38860_39160 , \38861_39161 , \38862_39162 , \38863_39163 , \38864_39164 , \38865_39165 , \38866_39166 ,
         \38867_39167 , \38868_39168 , \38869_39169 , \38870_39170 , \38871_39171 , \38872_39172 , \38873_39173 , \38874_39174 , \38875_39175 , \38876_39176 ,
         \38877_39177 , \38878_39178 , \38879_39179 , \38880_39180 , \38881_39181 , \38882_39182 , \38883_39183 , \38884_39184 , \38885_39185 , \38886_39186 ,
         \38887_39187 , \38888_39188 , \38889_39189 , \38890_39190 , \38891_39191 , \38892_39192 , \38893_39193 , \38894_39194 , \38895_39195 , \38896_39196 ,
         \38897_39197 , \38898_39198 , \38899_39199 , \38900_39200 , \38901_39201 , \38902_39202 , \38903_39203 , \38904_39204 , \38905_39205 , \38906_39206 ,
         \38907_39207 , \38908_39208 , \38909_39209 , \38910_39210 , \38911_39211 , \38912_39212 , \38913_39213 , \38914_39214 , \38915_39215 , \38916_39216 ,
         \38917_39217 , \38918_39218 , \38919_39219 , \38920_39220 , \38921_39221 , \38922_39222 , \38923_39223 , \38924_39224 , \38925_39225 , \38926_39226 ,
         \38927_39227 , \38928_39228 , \38929_39229 , \38930_39230 , \38931_39231 , \38932_39232 , \38933_39233 , \38934_39234 , \38935_39235 , \38936_39236 ,
         \38937_39237 , \38938_39238 , \38939_39239 , \38940_39240 , \38941_39241 , \38942_39242 , \38943_39243 , \38944_39244 , \38945_39245 , \38946_39246 ,
         \38947_39247 , \38948_39248 , \38949_39249 , \38950_39250 , \38951_39251 , \38952_39252 , \38953_39253 , \38954_39254 , \38955_39255 , \38956_39256 ,
         \38957_39257 , \38958_39258 , \38959_39259 , \38960_39260 , \38961_39261 , \38962_39262 , \38963_39263 , \38964_39264 , \38965_39265 , \38966_39266 ,
         \38967_39267 , \38968_39268 , \38969_39269 , \38970_39270 , \38971_39271 , \38972_39272 , \38973_39273 , \38974_39274 , \38975_39275 , \38976_39276 ,
         \38977_39277 , \38978_39278 , \38979_39279 , \38980_39280 , \38981_39281 , \38982_39282 , \38983_39283 , \38984_39284 , \38985_39285 , \38986_39286 ,
         \38987_39287 , \38988_39288 , \38989_39289 , \38990_39290 , \38991_39291 , \38992_39292 , \38993_39293 , \38994_39294 , \38995_39295 , \38996_39296 ,
         \38997_39297 , \38998_39298 , \38999_39299 , \39000_39300 , \39001_39301 , \39002_39302 , \39003_39303 , \39004_39304 , \39005_39305 , \39006_39306 ,
         \39007_39307 , \39008_39308 , \39009_39309 , \39010_39310 , \39011_39311 , \39012_39312 , \39013_39313 , \39014_39314 , \39015_39315 , \39016_39316 ,
         \39017_39317 , \39018_39318 , \39019_39319 , \39020_39320 , \39021_39321 , \39022_39322 , \39023_39323 , \39024_39324 , \39025_39325 , \39026_39326 ,
         \39027_39327 , \39028_39328 , \39029_39329 , \39030_39330 , \39031_39331 , \39032_39332 , \39033_39333 , \39034_39334_nG9b7b , \39035_39335 , \39036_39336 ,
         \39037_39337 , \39038_39338 , \39039_39339 , \39040_39340 , \39041_39341 , \39042_39342 , \39043_39343 , \39044_39344 , \39045_39345 , \39046_39346 ,
         \39047_39347 , \39048_39348 , \39049_39349 , \39050_39350 , \39051_39351 , \39052_39352 , \39053_39353 , \39054_39354 , \39055_39355 , \39056_39356 ,
         \39057_39357 , \39058_39358 , \39059_39359 , \39060_39360 , \39061_39361 , \39062_39362 , \39063_39363 , \39064_39364 , \39065_39365 , \39066_39366 ,
         \39067_39367 , \39068_39368 , \39069_39369 , \39070_39370 , \39071_39371 , \39072_39372 , \39073_39373 , \39074_39374 , \39075_39375 , \39076_39376 ,
         \39077_39377 , \39078_39378 , \39079_39379 , \39080_39380 , \39081_39381 , \39082_39382 , \39083_39383 , \39084_39384 , \39085_39385 , \39086_39386 ,
         \39087_39387 , \39088_39388 , \39089_39389 , \39090_39390 , \39091_39391 , \39092_39392 , \39093_39393 , \39094_39394 , \39095_39395 , \39096_39396 ,
         \39097_39397 , \39098_39398 , \39099_39399 , \39100_39400 , \39101_39401 , \39102_39402 , \39103_39403 , \39104_39404 , \39105_39405 , \39106_39406 ,
         \39107_39407 , \39108_39408 , \39109_39409 , \39110_39410 , \39111_39411 , \39112_39412 , \39113_39413 , \39114_39414 , \39115_39415 , \39116_39416 ,
         \39117_39417 , \39118_39418 , \39119_39419 , \39120_39420 , \39121_39421 , \39122_39422 , \39123_39423 , \39124_39424 , \39125_39425 , \39126_39426 ,
         \39127_39427 , \39128_39428 , \39129_39429 , \39130_39430 , \39131_39431 , \39132_39432 , \39133_39433 , \39134_39434 , \39135_39435 , \39136_39436 ,
         \39137_39437 , \39138_39438 , \39139_39439 , \39140_39440 , \39141_39441 , \39142_39442 , \39143_39443 , \39144_39444 , \39145_39445 , \39146_39446 ,
         \39147_39447 , \39148_39448 , \39149_39449 , \39150_39450 , \39151_39451 , \39152_39452 , \39153_39453 , \39154_39454 , \39155_39455 , \39156_39456 ,
         \39157_39457 , \39158_39458 , \39159_39459 , \39160_39460 , \39161_39461 , \39162_39462 , \39163_39463 , \39164_39464 , \39165_39465 , \39166_39466 ,
         \39167_39467 , \39168_39468 , \39169_39469 , \39170_39470 , \39171_39471 , \39172_39472 , \39173_39473 , \39174_39474 , \39175_39475 , \39176_39476 ,
         \39177_39477 , \39178_39478 , \39179_39479 , \39180_39480 , \39181_39481 , \39182_39482 , \39183_39483 , \39184_39484 , \39185_39485 , \39186_39486 ,
         \39187_39487 , \39188_39488 , \39189_39489 , \39190_39490 , \39191_39491 , \39192_39492 , \39193_39493 , \39194_39494 , \39195_39495 , \39196_39496 ,
         \39197_39497 , \39198_39498 , \39199_39499 , \39200_39500 , \39201_39501 , \39202_39502 , \39203_39503 , \39204_39504 , \39205_39505 , \39206_39506 ,
         \39207_39507 , \39208_39508 , \39209_39509 , \39210_39510 , \39211_39511 , \39212_39512 , \39213_39513 , \39214_39514 , \39215_39515 , \39216_39516 ,
         \39217_39517 , \39218_39518 , \39219_39519 , \39220_39520 , \39221_39521 , \39222_39522 , \39223_39523 , \39224_39524 , \39225_39525 , \39226_39526 ,
         \39227_39527 , \39228_39528 , \39229_39529 , \39230_39530 , \39231_39531 , \39232_39532 , \39233_39533 , \39234_39534 , \39235_39535 , \39236_39536 ,
         \39237_39537 , \39238_39538 , \39239_39539 , \39240_39540 , \39241_39541 , \39242_39542 , \39243_39543 , \39244_39544 , \39245_39545 , \39246_39546 ,
         \39247_39547 , \39248_39548 , \39249_39549 , \39250_39550 , \39251_39551 , \39252_39552 , \39253_39553 , \39254_39554 , \39255_39555 , \39256_39556 ,
         \39257_39557 , \39258_39558 , \39259_39559 , \39260_39560 , \39261_39561 , \39262_39562 , \39263_39563 , \39264_39564 , \39265_39565 , \39266_39566 ,
         \39267_39567 , \39268_39568 , \39269_39569 , \39270_39570 , \39271_39571 , \39272_39572 , \39273_39573 , \39274_39574 , \39275_39575 , \39276_39576 ,
         \39277_39577 , \39278_39578 , \39279_39579 , \39280_39580 , \39281_39581 , \39282_39582 , \39283_39583 , \39284_39584 , \39285_39585 , \39286_39586 ,
         \39287_39587 , \39288_39588 , \39289_39589 , \39290_39590 , \39291_39591_nG9b78 , \39292_39592 , \39293_39593 , \39294_39594 , \39295_39595 , \39296_39596 ,
         \39297_39597 , \39298_39598 , \39299_39599 , \39300_39600 , \39301_39601 , \39302_39602 , \39303_39603 , \39304_39604 , \39305_39605 , \39306_39606 ,
         \39307_39607 , \39308_39608 , \39309_39609 , \39310_39610 , \39311_39611 , \39312_39612 , \39313_39613 , \39314_39614 , \39315_39615 , \39316_39616 ,
         \39317_39617 , \39318_39618 , \39319_39619 , \39320_39620 , \39321_39621 , \39322_39622 , \39323_39623 , \39324_39624 , \39325_39625 , \39326_39626 ,
         \39327_39627 , \39328_39628 , \39329_39629 , \39330_39630 , \39331_39631 , \39332_39632 , \39333_39633 , \39334_39634 , \39335_39635 , \39336_39636 ,
         \39337_39637 , \39338_39638 , \39339_39639 , \39340_39640 , \39341_39641 , \39342_39642 , \39343_39643 , \39344_39644 , \39345_39645 , \39346_39646 ,
         \39347_39647 , \39348_39648 , \39349_39649 , \39350_39650 , \39351_39651 , \39352_39652 , \39353_39653 , \39354_39654 , \39355_39655 , \39356_39656 ,
         \39357_39657 , \39358_39658 , \39359_39659 , \39360_39660 , \39361_39661 , \39362_39662 , \39363_39663 , \39364_39664 , \39365_39665 , \39366_39666 ,
         \39367_39667 , \39368_39668 , \39369_39669 , \39370_39670 , \39371_39671 , \39372_39672 , \39373_39673 , \39374_39674 , \39375_39675 , \39376_39676 ,
         \39377_39677 , \39378_39678 , \39379_39679 , \39380_39680 , \39381_39681 , \39382_39682 , \39383_39683 , \39384_39684 , \39385_39685 , \39386_39686 ,
         \39387_39687 , \39388_39688 , \39389_39689 , \39390_39690 , \39391_39691 , \39392_39692 , \39393_39693 , \39394_39694 , \39395_39695 , \39396_39696 ,
         \39397_39697 , \39398_39698 , \39399_39699 , \39400_39700 , \39401_39701 , \39402_39702 , \39403_39703 , \39404_39704 , \39405_39705 , \39406_39706 ,
         \39407_39707 , \39408_39708 , \39409_39709 , \39410_39710 , \39411_39711 , \39412_39712 , \39413_39713 , \39414_39714 , \39415_39715 , \39416_39716 ,
         \39417_39717 , \39418_39718 , \39419_39719 , \39420_39720 , \39421_39721 , \39422_39722 , \39423_39723 , \39424_39724 , \39425_39725 , \39426_39726 ,
         \39427_39727 , \39428_39728 , \39429_39729 , \39430_39730 , \39431_39731 , \39432_39732 , \39433_39733 , \39434_39734 , \39435_39735 , \39436_39736 ,
         \39437_39737 , \39438_39738 , \39439_39739 , \39440_39740 , \39441_39741 , \39442_39742 , \39443_39743 , \39444_39744 , \39445_39745 , \39446_39746 ,
         \39447_39747 , \39448_39748 , \39449_39749 , \39450_39750 , \39451_39751 , \39452_39752 , \39453_39753 , \39454_39754 , \39455_39755 , \39456_39756 ,
         \39457_39757 , \39458_39758 , \39459_39759 , \39460_39760 , \39461_39761 , \39462_39762 , \39463_39763 , \39464_39764 , \39465_39765 , \39466_39766 ,
         \39467_39767 , \39468_39768 , \39469_39769 , \39470_39770 , \39471_39771 , \39472_39772 , \39473_39773 , \39474_39774 , \39475_39775 , \39476_39776 ,
         \39477_39777 , \39478_39778 , \39479_39779 , \39480_39780 , \39481_39781 , \39482_39782 , \39483_39783 , \39484_39784 , \39485_39785 , \39486_39786 ,
         \39487_39787 , \39488_39788 , \39489_39789 , \39490_39790 , \39491_39791 , \39492_39792 , \39493_39793 , \39494_39794 , \39495_39795 , \39496_39796 ,
         \39497_39797 , \39498_39798 , \39499_39799 , \39500_39800 , \39501_39801 , \39502_39802 , \39503_39803 , \39504_39804 , \39505_39805 , \39506_39806 ,
         \39507_39807 , \39508_39808 , \39509_39809 , \39510_39810 , \39511_39811 , \39512_39812 , \39513_39813 , \39514_39814 , \39515_39815 , \39516_39816 ,
         \39517_39817 , \39518_39818 , \39519_39819 , \39520_39820 , \39521_39821 , \39522_39822 , \39523_39823 , \39524_39824 , \39525_39825 , \39526_39826 ,
         \39527_39827 , \39528_39828 , \39529_39829 , \39530_39830 , \39531_39831 , \39532_39832 , \39533_39833 , \39534_39834 , \39535_39835 , \39536_39836 ,
         \39537_39837 , \39538_39838 , \39539_39839 , \39540_39840 , \39541_39841 , \39542_39842 , \39543_39843 , \39544_39844 , \39545_39845 , \39546_39846 ,
         \39547_39847 , \39548_39848 , \39549_39849 , \39550_39850 , \39551_39851 , \39552_39852 , \39553_39853 , \39554_39854 , \39555_39855 , \39556_39856 ,
         \39557_39857 , \39558_39858 , \39559_39859 , \39560_39860 , \39561_39861 , \39562_39862 , \39563_39863 , \39564_39864 , \39565_39865 , \39566_39866 ,
         \39567_39867 , \39568_39868 , \39569_39869 , \39570_39870 , \39571_39871 , \39572_39872 , \39573_39873 , \39574_39874 , \39575_39875 , \39576_39876 ,
         \39577_39877 , \39578_39878 , \39579_39879 , \39580_39880 , \39581_39881 , \39582_39882 , \39583_39883 , \39584_39884 , \39585_39885 , \39586_39886 ,
         \39587_39887 , \39588_39888 , \39589_39889 , \39590_39890 , \39591_39891 , \39592_39892 , \39593_39893 , \39594_39894 , \39595_39895 , \39596_39896 ,
         \39597_39897 , \39598_39898 , \39599_39899 , \39600_39900 , \39601_39901 , \39602_39902 , \39603_39903 , \39604_39904 , \39605_39905 , \39606_39906 ,
         \39607_39907 , \39608_39908 , \39609_39909 , \39610_39910 , \39611_39911 , \39612_39912 , \39613_39913 , \39614_39914 , \39615_39915 , \39616_39916 ,
         \39617_39917 , \39618_39918 , \39619_39919 , \39620_39920 , \39621_39921 , \39622_39922 , \39623_39923 , \39624_39924 , \39625_39925 , \39626_39926 ,
         \39627_39927 , \39628_39928 , \39629_39929 , \39630_39930 , \39631_39931 , \39632_39932 , \39633_39933 , \39634_39934 , \39635_39935 , \39636_39936 ,
         \39637_39937 , \39638_39938 , \39639_39939 , \39640_39940 , \39641_39941 , \39642_39942 , \39643_39943 , \39644_39944 , \39645_39945 , \39646_39946 ,
         \39647_39947 , \39648_39948 , \39649_39949 , \39650_39950 , \39651_39951 , \39652_39952 , \39653_39953 , \39654_39954 , \39655_39955 , \39656_39956 ,
         \39657_39957 , \39658_39958 , \39659_39959 , \39660_39960 , \39661_39961 , \39662_39962 , \39663_39963_nG9b75 , \39664_39964 , \39665_39965 , \39666_39966 ,
         \39667_39967 , \39668_39968 , \39669_39969 , \39670_39970 , \39671_39971 , \39672_39972 , \39673_39973 , \39674_39974 , \39675_39975 , \39676_39976 ,
         \39677_39977 , \39678_39978 , \39679_39979 , \39680_39980 , \39681_39981 , \39682_39982 , \39683_39983 , \39684_39984 , \39685_39985 , \39686_39986 ,
         \39687_39987 , \39688_39988 , \39689_39989 , \39690_39990 , \39691_39991 , \39692_39992 , \39693_39993 , \39694_39994 , \39695_39995 , \39696_39996 ,
         \39697_39997 , \39698_39998 , \39699_39999 , \39700_40000 , \39701_40001 , \39702_40002 , \39703_40003 , \39704_40004 , \39705_40005 , \39706_40006 ,
         \39707_40007 , \39708_40008 , \39709_40009 , \39710_40010 , \39711_40011 , \39712_40012 , \39713_40013 , \39714_40014 , \39715_40015 , \39716_40016 ,
         \39717_40017 , \39718_40018 , \39719_40019 , \39720_40020 , \39721_40021 , \39722_40022 , \39723_40023 , \39724_40024 , \39725_40025 , \39726_40026 ,
         \39727_40027 , \39728_40028 , \39729_40029 , \39730_40030 , \39731_40031 , \39732_40032 , \39733_40033 , \39734_40034 , \39735_40035 , \39736_40036 ,
         \39737_40037 , \39738_40038 , \39739_40039 , \39740_40040 , \39741_40041 , \39742_40042 , \39743_40043 , \39744_40044 , \39745_40045 , \39746_40046 ,
         \39747_40047 , \39748_40048 , \39749_40049 , \39750_40050 , \39751_40051 , \39752_40052 , \39753_40053 , \39754_40054 , \39755_40055 , \39756_40056 ,
         \39757_40057 , \39758_40058 , \39759_40059 , \39760_40060 , \39761_40061 , \39762_40062 , \39763_40063 , \39764_40064 , \39765_40065 , \39766_40066 ,
         \39767_40067 , \39768_40068 , \39769_40069 , \39770_40070 , \39771_40071 , \39772_40072 , \39773_40073 , \39774_40074 , \39775_40075 , \39776_40076 ,
         \39777_40077 , \39778_40078 , \39779_40079 , \39780_40080 , \39781_40081 , \39782_40082 , \39783_40083 , \39784_40084 , \39785_40085 , \39786_40086 ,
         \39787_40087 , \39788_40088 , \39789_40089 , \39790_40090 , \39791_40091 , \39792_40092 , \39793_40093 , \39794_40094 , \39795_40095 , \39796_40096 ,
         \39797_40097 , \39798_40098 , \39799_40099 , \39800_40100 , \39801_40101 , \39802_40102 , \39803_40103 , \39804_40104 , \39805_40105 , \39806_40106 ,
         \39807_40107 , \39808_40108 , \39809_40109 , \39810_40110 , \39811_40111 , \39812_40112 , \39813_40113 , \39814_40114 , \39815_40115 , \39816_40116 ,
         \39817_40117 , \39818_40118 , \39819_40119 , \39820_40120 , \39821_40121 , \39822_40122 , \39823_40123 , \39824_40124 , \39825_40125 , \39826_40126 ,
         \39827_40127 , \39828_40128 , \39829_40129 , \39830_40130 , \39831_40131 , \39832_40132 , \39833_40133 , \39834_40134 , \39835_40135 , \39836_40136 ,
         \39837_40137 , \39838_40138 , \39839_40139 , \39840_40140 , \39841_40141 , \39842_40142 , \39843_40143 , \39844_40144 , \39845_40145 , \39846_40146 ,
         \39847_40147 , \39848_40148 , \39849_40149 , \39850_40150 , \39851_40151 , \39852_40152 , \39853_40153 , \39854_40154 , \39855_40155 , \39856_40156 ,
         \39857_40157 , \39858_40158 , \39859_40159 , \39860_40160 , \39861_40161 , \39862_40162 , \39863_40163 , \39864_40164 , \39865_40165 , \39866_40166 ,
         \39867_40167 , \39868_40168 , \39869_40169 , \39870_40170 , \39871_40171 , \39872_40172 , \39873_40173 , \39874_40174 , \39875_40175 , \39876_40176 ,
         \39877_40177 , \39878_40178 , \39879_40179 , \39880_40180 , \39881_40181 , \39882_40182 , \39883_40183 , \39884_40184 , \39885_40185 , \39886_40186 ,
         \39887_40187 , \39888_40188 , \39889_40189 , \39890_40190 , \39891_40191 , \39892_40192 , \39893_40193 , \39894_40194 , \39895_40195 , \39896_40196 ,
         \39897_40197 , \39898_40198 , \39899_40199 , \39900_40200 , \39901_40201 , \39902_40202 , \39903_40203 , \39904_40204_nG9b72 , \39905_40205 , \39906_40206 ,
         \39907_40207 , \39908_40208 , \39909_40209 , \39910_40210 , \39911_40211 , \39912_40212 , \39913_40213 , \39914_40214 , \39915_40215 , \39916_40216 ,
         \39917_40217 , \39918_40218 , \39919_40219 , \39920_40220 , \39921_40221 , \39922_40222 , \39923_40223 , \39924_40224 , \39925_40225 , \39926_40226 ,
         \39927_40227 , \39928_40228 , \39929_40229 , \39930_40230 , \39931_40231 , \39932_40232 , \39933_40233 , \39934_40234 , \39935_40235 , \39936_40236 ,
         \39937_40237 , \39938_40238 , \39939_40239 , \39940_40240 , \39941_40241 , \39942_40242 , \39943_40243 , \39944_40244 , \39945_40245 , \39946_40246 ,
         \39947_40247 , \39948_40248 , \39949_40249 , \39950_40250 , \39951_40251 , \39952_40252 , \39953_40253 , \39954_40254 , \39955_40255 , \39956_40256 ,
         \39957_40257 , \39958_40258 , \39959_40259 , \39960_40260 , \39961_40261 , \39962_40262 , \39963_40263 , \39964_40264 , \39965_40265 , \39966_40266 ,
         \39967_40267 , \39968_40268 , \39969_40269 , \39970_40270 , \39971_40271 , \39972_40272 , \39973_40273 , \39974_40274 , \39975_40275 , \39976_40276 ,
         \39977_40277 , \39978_40278 , \39979_40279 , \39980_40280 , \39981_40281 , \39982_40282 , \39983_40283 , \39984_40284 , \39985_40285 , \39986_40286 ,
         \39987_40287 , \39988_40288 , \39989_40289 , \39990_40290 , \39991_40291 , \39992_40292 , \39993_40293 , \39994_40294 , \39995_40295 , \39996_40296 ,
         \39997_40297 , \39998_40298 , \39999_40299 , \40000_40300 , \40001_40301 , \40002_40302 , \40003_40303 , \40004_40304 , \40005_40305 , \40006_40306 ,
         \40007_40307 , \40008_40308 , \40009_40309 , \40010_40310 , \40011_40311 , \40012_40312 , \40013_40313 , \40014_40314 , \40015_40315 , \40016_40316 ,
         \40017_40317 , \40018_40318 , \40019_40319 , \40020_40320 , \40021_40321 , \40022_40322 , \40023_40323 , \40024_40324 , \40025_40325 , \40026_40326 ,
         \40027_40327 , \40028_40328 , \40029_40329 , \40030_40330 , \40031_40331 , \40032_40332 , \40033_40333 , \40034_40334 , \40035_40335 , \40036_40336 ,
         \40037_40337 , \40038_40338 , \40039_40339 , \40040_40340 , \40041_40341 , \40042_40342 , \40043_40343 , \40044_40344 , \40045_40345 , \40046_40346 ,
         \40047_40347 , \40048_40348 , \40049_40349 , \40050_40350 , \40051_40351 , \40052_40352 , \40053_40353 , \40054_40354 , \40055_40355 , \40056_40356 ,
         \40057_40357 , \40058_40358 , \40059_40359 , \40060_40360 , \40061_40361 , \40062_40362 , \40063_40363 , \40064_40364 , \40065_40365 , \40066_40366 ,
         \40067_40367 , \40068_40368 , \40069_40369 , \40070_40370 , \40071_40371 , \40072_40372 , \40073_40373 , \40074_40374 , \40075_40375 , \40076_40376 ,
         \40077_40377 , \40078_40378 , \40079_40379 , \40080_40380 , \40081_40381 , \40082_40382 , \40083_40383 , \40084_40384 , \40085_40385 , \40086_40386 ,
         \40087_40387 , \40088_40388 , \40089_40389 , \40090_40390 , \40091_40391 , \40092_40392 , \40093_40393 , \40094_40394 , \40095_40395 , \40096_40396 ,
         \40097_40397 , \40098_40398 , \40099_40399 , \40100_40400 , \40101_40401 , \40102_40402 , \40103_40403 , \40104_40404 , \40105_40405 , \40106_40406 ,
         \40107_40407 , \40108_40408 , \40109_40409 , \40110_40410 , \40111_40411 , \40112_40412 , \40113_40413 , \40114_40414 , \40115_40415 , \40116_40416 ,
         \40117_40417 , \40118_40418 , \40119_40419 , \40120_40420 , \40121_40421 , \40122_40422 , \40123_40423 , \40124_40424 , \40125_40425 , \40126_40426 ,
         \40127_40427 , \40128_40428 , \40129_40429 , \40130_40430 , \40131_40431 , \40132_40432 , \40133_40433 , \40134_40434 , \40135_40435 , \40136_40436 ,
         \40137_40437 , \40138_40438 , \40139_40439 , \40140_40440 , \40141_40441 , \40142_40442 , \40143_40443 , \40144_40444 , \40145_40445 , \40146_40446 ,
         \40147_40447 , \40148_40448 , \40149_40449 , \40150_40450 , \40151_40451 , \40152_40452_nG9b6f , \40153_40453 , \40154_40454 , \40155_40455 , \40156_40456 ,
         \40157_40457 , \40158_40458 , \40159_40459 , \40160_40460 , \40161_40461 , \40162_40462 , \40163_40463 , \40164_40464 , \40165_40465 , \40166_40466 ,
         \40167_40467 , \40168_40468 , \40169_40469 , \40170_40470 , \40171_40471 , \40172_40472 , \40173_40473 , \40174_40474 , \40175_40475 , \40176_40476 ,
         \40177_40477 , \40178_40478 , \40179_40479 , \40180_40480 , \40181_40481 , \40182_40482 , \40183_40483 , \40184_40484 , \40185_40485 , \40186_40486 ,
         \40187_40487 , \40188_40488 , \40189_40489 , \40190_40490 , \40191_40491 , \40192_40492 , \40193_40493 , \40194_40494 , \40195_40495 , \40196_40496 ,
         \40197_40497 , \40198_40498 , \40199_40499 , \40200_40500 , \40201_40501 , \40202_40502 , \40203_40503 , \40204_40504 , \40205_40505 , \40206_40506 ,
         \40207_40507 , \40208_40508 , \40209_40509 , \40210_40510 , \40211_40511 , \40212_40512 , \40213_40513 , \40214_40514 , \40215_40515 , \40216_40516 ,
         \40217_40517 , \40218_40518 , \40219_40519 , \40220_40520 , \40221_40521 , \40222_40522 , \40223_40523 , \40224_40524 , \40225_40525 , \40226_40526 ,
         \40227_40527 , \40228_40528 , \40229_40529 , \40230_40530 , \40231_40531 , \40232_40532 , \40233_40533 , \40234_40534 , \40235_40535 , \40236_40536 ,
         \40237_40537 , \40238_40538 , \40239_40539 , \40240_40540 , \40241_40541 , \40242_40542 , \40243_40543 , \40244_40544 , \40245_40545 , \40246_40546 ,
         \40247_40547 , \40248_40548 , \40249_40549 , \40250_40550 , \40251_40551 , \40252_40552 , \40253_40553 , \40254_40554 , \40255_40555 , \40256_40556 ,
         \40257_40557 , \40258_40558 , \40259_40559 , \40260_40560 , \40261_40561 , \40262_40562 , \40263_40563 , \40264_40564 , \40265_40565 , \40266_40566 ,
         \40267_40567 , \40268_40568 , \40269_40569 , \40270_40570 , \40271_40571 , \40272_40572 , \40273_40573 , \40274_40574 , \40275_40575 , \40276_40576 ,
         \40277_40577 , \40278_40578 , \40279_40579 , \40280_40580 , \40281_40581 , \40282_40582 , \40283_40583 , \40284_40584 , \40285_40585 , \40286_40586 ,
         \40287_40587 , \40288_40588 , \40289_40589 , \40290_40590 , \40291_40591 , \40292_40592 , \40293_40593 , \40294_40594 , \40295_40595 , \40296_40596 ,
         \40297_40597 , \40298_40598 , \40299_40599 , \40300_40600 , \40301_40601 , \40302_40602 , \40303_40603 , \40304_40604 , \40305_40605 , \40306_40606 ,
         \40307_40607 , \40308_40608 , \40309_40609 , \40310_40610 , \40311_40611 , \40312_40612 , \40313_40613 , \40314_40614 , \40315_40615 , \40316_40616 ,
         \40317_40617 , \40318_40618 , \40319_40619 , \40320_40620 , \40321_40621 , \40322_40622 , \40323_40623 , \40324_40624 , \40325_40625 , \40326_40626 ,
         \40327_40627 , \40328_40628 , \40329_40629 , \40330_40630 , \40331_40631 , \40332_40632 , \40333_40633 , \40334_40634 , \40335_40635 , \40336_40636 ,
         \40337_40637 , \40338_40638 , \40339_40639 , \40340_40640 , \40341_40641 , \40342_40642 , \40343_40643 , \40344_40644 , \40345_40645 , \40346_40646 ,
         \40347_40647 , \40348_40648 , \40349_40649 , \40350_40650 , \40351_40651 , \40352_40652 , \40353_40653 , \40354_40654 , \40355_40655 , \40356_40656 ,
         \40357_40657 , \40358_40658 , \40359_40659 , \40360_40660 , \40361_40661 , \40362_40662 , \40363_40663 , \40364_40664 , \40365_40665 , \40366_40666 ,
         \40367_40667 , \40368_40668 , \40369_40669 , \40370_40670 , \40371_40671 , \40372_40672 , \40373_40673 , \40374_40674 , \40375_40675 , \40376_40676 ,
         \40377_40677 , \40378_40678 , \40379_40679 , \40380_40680 , \40381_40681 , \40382_40682 , \40383_40683 , \40384_40684 , \40385_40685 , \40386_40686 ,
         \40387_40687 , \40388_40688 , \40389_40689 , \40390_40690 , \40391_40691 , \40392_40692 , \40393_40693 , \40394_40694 , \40395_40695 , \40396_40696 ,
         \40397_40697 , \40398_40698 , \40399_40699 , \40400_40700 , \40401_40701 , \40402_40702 , \40403_40703 , \40404_40704 , \40405_40705 , \40406_40706 ,
         \40407_40707 , \40408_40708 , \40409_40709 , \40410_40710 , \40411_40711 , \40412_40712 , \40413_40713 , \40414_40714 , \40415_40715 , \40416_40716 ,
         \40417_40717 , \40418_40718 , \40419_40719 , \40420_40720 , \40421_40721 , \40422_40722 , \40423_40723 , \40424_40724 , \40425_40725 , \40426_40726 ,
         \40427_40727 , \40428_40728 , \40429_40729 , \40430_40730 , \40431_40731 , \40432_40732 , \40433_40733 , \40434_40734 , \40435_40735 , \40436_40736 ,
         \40437_40737 , \40438_40738 , \40439_40739 , \40440_40740 , \40441_40741 , \40442_40742 , \40443_40743 , \40444_40744 , \40445_40745 , \40446_40746 ,
         \40447_40747 , \40448_40748 , \40449_40749 , \40450_40750 , \40451_40751 , \40452_40752 , \40453_40753 , \40454_40754 , \40455_40755 , \40456_40756 ,
         \40457_40757 , \40458_40758 , \40459_40759 , \40460_40760 , \40461_40761 , \40462_40762 , \40463_40763 , \40464_40764 , \40465_40765 , \40466_40766 ,
         \40467_40767 , \40468_40768 , \40469_40769 , \40470_40770 , \40471_40771 , \40472_40772 , \40473_40773 , \40474_40774 , \40475_40775 , \40476_40776 ,
         \40477_40777 , \40478_40778 , \40479_40779 , \40480_40780 , \40481_40781 , \40482_40782 , \40483_40783 , \40484_40784 , \40485_40785 , \40486_40786 ,
         \40487_40787 , \40488_40788 , \40489_40789 , \40490_40790 , \40491_40791 , \40492_40792 , \40493_40793 , \40494_40794 , \40495_40795 , \40496_40796 ,
         \40497_40797 , \40498_40798 , \40499_40799 , \40500_40800 , \40501_40801 , \40502_40802 , \40503_40803 , \40504_40804 , \40505_40805 , \40506_40806 ,
         \40507_40807 , \40508_40808 , \40509_40809 , \40510_40810 , \40511_40811 , \40512_40812 , \40513_40813 , \40514_40814 , \40515_40815 , \40516_40816 ,
         \40517_40817 , \40518_40818 , \40519_40819 , \40520_40820 , \40521_40821 , \40522_40822 , \40523_40823 , \40524_40824 , \40525_40825 , \40526_40826 ,
         \40527_40827 , \40528_40828 , \40529_40829 , \40530_40830 , \40531_40831 , \40532_40832 , \40533_40833 , \40534_40834 , \40535_40835 , \40536_40836 ,
         \40537_40837 , \40538_40838 , \40539_40839 , \40540_40840 , \40541_40841 , \40542_40842 , \40543_40843_nG9b6c , \40544_40844 , \40545_40845 , \40546_40846 ,
         \40547_40847 , \40548_40848 , \40549_40849 , \40550_40850 , \40551_40851 , \40552_40852 , \40553_40853 , \40554_40854 , \40555_40855 , \40556_40856 ,
         \40557_40857 , \40558_40858 , \40559_40859 , \40560_40860 , \40561_40861 , \40562_40862 , \40563_40863 , \40564_40864 , \40565_40865 , \40566_40866 ,
         \40567_40867 , \40568_40868 , \40569_40869 , \40570_40870 , \40571_40871 , \40572_40872 , \40573_40873 , \40574_40874 , \40575_40875 , \40576_40876 ,
         \40577_40877 , \40578_40878 , \40579_40879 , \40580_40880 , \40581_40881 , \40582_40882 , \40583_40883 , \40584_40884 , \40585_40885 , \40586_40886 ,
         \40587_40887 , \40588_40888 , \40589_40889 , \40590_40890 , \40591_40891 , \40592_40892 , \40593_40893 , \40594_40894 , \40595_40895 , \40596_40896 ,
         \40597_40897 , \40598_40898 , \40599_40899 , \40600_40900 , \40601_40901 , \40602_40902 , \40603_40903 , \40604_40904 , \40605_40905 , \40606_40906 ,
         \40607_40907 , \40608_40908 , \40609_40909 , \40610_40910 , \40611_40911 , \40612_40912 , \40613_40913 , \40614_40914 , \40615_40915 , \40616_40916 ,
         \40617_40917 , \40618_40918 , \40619_40919 , \40620_40920 , \40621_40921 , \40622_40922 , \40623_40923 , \40624_40924 , \40625_40925 , \40626_40926 ,
         \40627_40927 , \40628_40928 , \40629_40929 , \40630_40930 , \40631_40931 , \40632_40932 , \40633_40933 , \40634_40934 , \40635_40935 , \40636_40936 ,
         \40637_40937 , \40638_40938 , \40639_40939 , \40640_40940 , \40641_40941 , \40642_40942 , \40643_40943 , \40644_40944 , \40645_40945 , \40646_40946 ,
         \40647_40947 , \40648_40948 , \40649_40949 , \40650_40950 , \40651_40951 , \40652_40952 , \40653_40953 , \40654_40954 , \40655_40955 , \40656_40956 ,
         \40657_40957 , \40658_40958 , \40659_40959 , \40660_40960 , \40661_40961 , \40662_40962 , \40663_40963 , \40664_40964 , \40665_40965 , \40666_40966 ,
         \40667_40967 , \40668_40968 , \40669_40969 , \40670_40970 , \40671_40971 , \40672_40972 , \40673_40973 , \40674_40974 , \40675_40975 , \40676_40976 ,
         \40677_40977 , \40678_40978 , \40679_40979 , \40680_40980 , \40681_40981 , \40682_40982 , \40683_40983 , \40684_40984 , \40685_40985 , \40686_40986 ,
         \40687_40987 , \40688_40988 , \40689_40989 , \40690_40990 , \40691_40991 , \40692_40992 , \40693_40993 , \40694_40994 , \40695_40995 , \40696_40996 ,
         \40697_40997 , \40698_40998 , \40699_40999 , \40700_41000 , \40701_41001 , \40702_41002 , \40703_41003 , \40704_41004 , \40705_41005 , \40706_41006 ,
         \40707_41007 , \40708_41008 , \40709_41009 , \40710_41010 , \40711_41011 , \40712_41012 , \40713_41013 , \40714_41014 , \40715_41015 , \40716_41016 ,
         \40717_41017 , \40718_41018 , \40719_41019 , \40720_41020 , \40721_41021 , \40722_41022 , \40723_41023 , \40724_41024 , \40725_41025 , \40726_41026 ,
         \40727_41027 , \40728_41028 , \40729_41029 , \40730_41030 , \40731_41031 , \40732_41032 , \40733_41033 , \40734_41034 , \40735_41035 , \40736_41036 ,
         \40737_41037 , \40738_41038 , \40739_41039 , \40740_41040_nG9b69 , \40741_41041 , \40742_41042 , \40743_41043 , \40744_41044 , \40745_41045 , \40746_41046 ,
         \40747_41047 , \40748_41048 , \40749_41049 , \40750_41050 , \40751_41051 , \40752_41052 , \40753_41053 , \40754_41054 , \40755_41055 , \40756_41056 ,
         \40757_41057 , \40758_41058 , \40759_41059 , \40760_41060 , \40761_41061 , \40762_41062 , \40763_41063 , \40764_41064 , \40765_41065 , \40766_41066 ,
         \40767_41067 , \40768_41068 , \40769_41069 , \40770_41070 , \40771_41071 , \40772_41072 , \40773_41073 , \40774_41074 , \40775_41075 , \40776_41076 ,
         \40777_41077 , \40778_41078 , \40779_41079 , \40780_41080 , \40781_41081 , \40782_41082 , \40783_41083 , \40784_41084 , \40785_41085 , \40786_41086 ,
         \40787_41087 , \40788_41088 , \40789_41089 , \40790_41090 , \40791_41091 , \40792_41092 , \40793_41093 , \40794_41094 , \40795_41095 , \40796_41096 ,
         \40797_41097 , \40798_41098 , \40799_41099 , \40800_41100 , \40801_41101 , \40802_41102 , \40803_41103 , \40804_41104 , \40805_41105 , \40806_41106 ,
         \40807_41107 , \40808_41108 , \40809_41109 , \40810_41110 , \40811_41111 , \40812_41112 , \40813_41113 , \40814_41114 , \40815_41115 , \40816_41116 ,
         \40817_41117 , \40818_41118 , \40819_41119 , \40820_41120 , \40821_41121 , \40822_41122 , \40823_41123 , \40824_41124 , \40825_41125 , \40826_41126 ,
         \40827_41127 , \40828_41128 , \40829_41129 , \40830_41130 , \40831_41131 , \40832_41132 , \40833_41133 , \40834_41134 , \40835_41135 , \40836_41136 ,
         \40837_41137 , \40838_41138 , \40839_41139 , \40840_41140 , \40841_41141 , \40842_41142 , \40843_41143 , \40844_41144 , \40845_41145 , \40846_41146 ,
         \40847_41147 , \40848_41148 , \40849_41149 , \40850_41150 , \40851_41151 , \40852_41152 , \40853_41153 , \40854_41154 , \40855_41155 , \40856_41156 ,
         \40857_41157 , \40858_41158 , \40859_41159 , \40860_41160 , \40861_41161 , \40862_41162 , \40863_41163 , \40864_41164 , \40865_41165 , \40866_41166 ,
         \40867_41167 , \40868_41168 , \40869_41169 , \40870_41170 , \40871_41171 , \40872_41172 , \40873_41173 , \40874_41174 , \40875_41175 , \40876_41176 ,
         \40877_41177 , \40878_41178 , \40879_41179 , \40880_41180 , \40881_41181 , \40882_41182 , \40883_41183 , \40884_41184 , \40885_41185 , \40886_41186 ,
         \40887_41187 , \40888_41188 , \40889_41189 , \40890_41190 , \40891_41191 , \40892_41192 , \40893_41193 , \40894_41194 , \40895_41195 , \40896_41196 ,
         \40897_41197 , \40898_41198 , \40899_41199 , \40900_41200 , \40901_41201 , \40902_41202 , \40903_41203 , \40904_41204 , \40905_41205 , \40906_41206 ,
         \40907_41207 , \40908_41208 , \40909_41209 , \40910_41210 , \40911_41211 , \40912_41212 , \40913_41213 , \40914_41214 , \40915_41215 , \40916_41216 ,
         \40917_41217 , \40918_41218 , \40919_41219 , \40920_41220 , \40921_41221 , \40922_41222 , \40923_41223 , \40924_41224 , \40925_41225 , \40926_41226 ,
         \40927_41227 , \40928_41228 , \40929_41229 , \40930_41230 , \40931_41231 , \40932_41232 , \40933_41233 , \40934_41234 , \40935_41235 , \40936_41236 ,
         \40937_41237 , \40938_41238 , \40939_41239 , \40940_41240 , \40941_41241 , \40942_41242 , \40943_41243 , \40944_41244 , \40945_41245 , \40946_41246 ,
         \40947_41247 , \40948_41248 , \40949_41249 , \40950_41250 , \40951_41251 , \40952_41252 , \40953_41253 , \40954_41254 , \40955_41255 , \40956_41256 ,
         \40957_41257 , \40958_41258 , \40959_41259 , \40960_41260 , \40961_41261 , \40962_41262 , \40963_41263 , \40964_41264 , \40965_41265 , \40966_41266 ,
         \40967_41267 , \40968_41268 , \40969_41269 , \40970_41270 , \40971_41271 , \40972_41272 , \40973_41273 , \40974_41274 , \40975_41275 , \40976_41276 ,
         \40977_41277 , \40978_41278 , \40979_41279 , \40980_41280 , \40981_41281 , \40982_41282 , \40983_41283 , \40984_41284 , \40985_41285 , \40986_41286 ,
         \40987_41287 , \40988_41288 , \40989_41289 , \40990_41290 , \40991_41291 , \40992_41292 , \40993_41293 , \40994_41294 , \40995_41295 , \40996_41296 ,
         \40997_41297 , \40998_41298 , \40999_41299 , \41000_41300 , \41001_41301 , \41002_41302 , \41003_41303 , \41004_41304 , \41005_41305 , \41006_41306 ,
         \41007_41307 , \41008_41308 , \41009_41309 , \41010_41310 , \41011_41311 , \41012_41312 , \41013_41313 , \41014_41314 , \41015_41315 , \41016_41316 ,
         \41017_41317 , \41018_41318 , \41019_41319 , \41020_41320 , \41021_41321 , \41022_41322 , \41023_41323 , \41024_41324 , \41025_41325 , \41026_41326 ,
         \41027_41327 , \41028_41328 , \41029_41329 , \41030_41330 , \41031_41331 , \41032_41332 , \41033_41333 , \41034_41334 , \41035_41335 , \41036_41336 ,
         \41037_41337 , \41038_41338 , \41039_41339 , \41040_41340 , \41041_41341 , \41042_41342 , \41043_41343 , \41044_41344 , \41045_41345 , \41046_41346 ,
         \41047_41347 , \41048_41348 , \41049_41349 , \41050_41350 , \41051_41351 , \41052_41352 , \41053_41353 , \41054_41354 , \41055_41355 , \41056_41356 ,
         \41057_41357 , \41058_41358 , \41059_41359 , \41060_41360 , \41061_41361 , \41062_41362 , \41063_41363 , \41064_41364 , \41065_41365 , \41066_41366 ,
         \41067_41367 , \41068_41368 , \41069_41369 , \41070_41370 , \41071_41371 , \41072_41372 , \41073_41373 , \41074_41374 , \41075_41375 , \41076_41376 ,
         \41077_41377 , \41078_41378 , \41079_41379 , \41080_41380 , \41081_41381_nG9b66 , \41082_41382 , \41083_41383 , \41084_41384 , \41085_41385 , \41086_41386 ,
         \41087_41387 , \41088_41388 , \41089_41389 , \41090_41390 , \41091_41391 , \41092_41392 , \41093_41393 , \41094_41394 , \41095_41395 , \41096_41396 ,
         \41097_41397 , \41098_41398 , \41099_41399 , \41100_41400 , \41101_41401 , \41102_41402 , \41103_41403 , \41104_41404 , \41105_41405 , \41106_41406 ,
         \41107_41407 , \41108_41408 , \41109_41409 , \41110_41410 , \41111_41411 , \41112_41412 , \41113_41413 , \41114_41414 , \41115_41415 , \41116_41416 ,
         \41117_41417 , \41118_41418 , \41119_41419 , \41120_41420 , \41121_41421 , \41122_41422 , \41123_41423 , \41124_41424 , \41125_41425 , \41126_41426 ,
         \41127_41427 , \41128_41428 , \41129_41429 , \41130_41430 , \41131_41431 , \41132_41432 , \41133_41433 , \41134_41434 , \41135_41435 , \41136_41436 ,
         \41137_41437 , \41138_41438 , \41139_41439 , \41140_41440 , \41141_41441 , \41142_41442 , \41143_41443 , \41144_41444 , \41145_41445 , \41146_41446 ,
         \41147_41447 , \41148_41448 , \41149_41449 , \41150_41450 , \41151_41451 , \41152_41452 , \41153_41453 , \41154_41454 , \41155_41455 , \41156_41456 ,
         \41157_41457 , \41158_41458 , \41159_41459 , \41160_41460 , \41161_41461 , \41162_41462 , \41163_41463 , \41164_41464 , \41165_41465 , \41166_41466 ,
         \41167_41467 , \41168_41468 , \41169_41469 , \41170_41470 , \41171_41471 , \41172_41472 , \41173_41473 , \41174_41474 , \41175_41475 , \41176_41476 ,
         \41177_41477 , \41178_41478 , \41179_41479 , \41180_41480 , \41181_41481 , \41182_41482 , \41183_41483 , \41184_41484 , \41185_41485 , \41186_41486 ,
         \41187_41487 , \41188_41488 , \41189_41489 , \41190_41490 , \41191_41491 , \41192_41492 , \41193_41493 , \41194_41494 , \41195_41495 , \41196_41496 ,
         \41197_41497 , \41198_41498 , \41199_41499 , \41200_41500 , \41201_41501 , \41202_41502 , \41203_41503 , \41204_41504 , \41205_41505 , \41206_41506 ,
         \41207_41507 , \41208_41508 , \41209_41509 , \41210_41510 , \41211_41511 , \41212_41512 , \41213_41513 , \41214_41514 , \41215_41515 , \41216_41516 ,
         \41217_41517 , \41218_41518 , \41219_41519 , \41220_41520 , \41221_41521 , \41222_41522 , \41223_41523 , \41224_41524 , \41225_41525 , \41226_41526 ,
         \41227_41527 , \41228_41528 , \41229_41529 , \41230_41530 , \41231_41531 , \41232_41532 , \41233_41533 , \41234_41534 , \41235_41535 , \41236_41536 ,
         \41237_41537 , \41238_41538 , \41239_41539 , \41240_41540 , \41241_41541 , \41242_41542 , \41243_41543 , \41244_41544 , \41245_41545 , \41246_41546 ,
         \41247_41547 , \41248_41548 , \41249_41549 , \41250_41550 , \41251_41551 , \41252_41552 , \41253_41553 , \41254_41554 , \41255_41555 , \41256_41556 ,
         \41257_41557 , \41258_41558 , \41259_41559 , \41260_41560 , \41261_41561 , \41262_41562 , \41263_41563 , \41264_41564 , \41265_41565 , \41266_41566 ,
         \41267_41567 , \41268_41568 , \41269_41569 , \41270_41570 , \41271_41571 , \41272_41572 , \41273_41573 , \41274_41574 , \41275_41575 , \41276_41576 ,
         \41277_41577 , \41278_41578 , \41279_41579 , \41280_41580 , \41281_41581 , \41282_41582 , \41283_41583 , \41284_41584 , \41285_41585 , \41286_41586 ,
         \41287_41587 , \41288_41588 , \41289_41589 , \41290_41590 , \41291_41591 , \41292_41592 , \41293_41593 , \41294_41594 , \41295_41595 , \41296_41596 ,
         \41297_41597 , \41298_41598 , \41299_41599 , \41300_41600 , \41301_41601 , \41302_41602 , \41303_41603 , \41304_41604 , \41305_41605 , \41306_41606 ,
         \41307_41607 , \41308_41608 , \41309_41609 , \41310_41610 , \41311_41611 , \41312_41612 , \41313_41613 , \41314_41614 , \41315_41615 , \41316_41616 ,
         \41317_41617 , \41318_41618 , \41319_41619 , \41320_41620 , \41321_41621 , \41322_41622 , \41323_41623 , \41324_41624 , \41325_41625 , \41326_41626 ,
         \41327_41627 , \41328_41628 , \41329_41629 , \41330_41630 , \41331_41631 , \41332_41632 , \41333_41633 , \41334_41634 , \41335_41635 , \41336_41636 ,
         \41337_41637 , \41338_41638 , \41339_41639 , \41340_41640 , \41341_41641 , \41342_41642 , \41343_41643 , \41344_41644 , \41345_41645 , \41346_41646 ,
         \41347_41647 , \41348_41648 , \41349_41649 , \41350_41650 , \41351_41651 , \41352_41652 , \41353_41653 , \41354_41654 , \41355_41655 , \41356_41656 ,
         \41357_41657 , \41358_41658 , \41359_41659 , \41360_41660 , \41361_41661 , \41362_41662 , \41363_41663 , \41364_41664 , \41365_41665 , \41366_41666 ,
         \41367_41667 , \41368_41668 , \41369_41669 , \41370_41670 , \41371_41671 , \41372_41672 , \41373_41673 , \41374_41674 , \41375_41675 , \41376_41676 ,
         \41377_41677 , \41378_41678 , \41379_41679 , \41380_41680 , \41381_41681 , \41382_41682 , \41383_41683 , \41384_41684 , \41385_41685_nG9b63 , \41386_41686 ,
         \41387_41687 , \41388_41688 , \41389_41689 , \41390_41690 , \41391_41691 , \41392_41692 , \41393_41693 , \41394_41694 , \41395_41695 , \41396_41696 ,
         \41397_41697 , \41398_41698 , \41399_41699 , \41400_41700 , \41401_41701 , \41402_41702 , \41403_41703 , \41404_41704 , \41405_41705 , \41406_41706 ,
         \41407_41707 , \41408_41708 , \41409_41709 , \41410_41710 , \41411_41711 , \41412_41712 , \41413_41713 , \41414_41714 , \41415_41715 , \41416_41716 ,
         \41417_41717 , \41418_41718 , \41419_41719 , \41420_41720 , \41421_41721 , \41422_41722 , \41423_41723 , \41424_41724 , \41425_41725 , \41426_41726 ,
         \41427_41727 , \41428_41728 , \41429_41729 , \41430_41730 , \41431_41731 , \41432_41732 , \41433_41733 , \41434_41734 , \41435_41735 , \41436_41736 ,
         \41437_41737 , \41438_41738 , \41439_41739 , \41440_41740 , \41441_41741 , \41442_41742 , \41443_41743 , \41444_41744 , \41445_41745 , \41446_41746 ,
         \41447_41747 , \41448_41748 , \41449_41749 , \41450_41750 , \41451_41751 , \41452_41752 , \41453_41753 , \41454_41754 , \41455_41755 , \41456_41756 ,
         \41457_41757 , \41458_41758 , \41459_41759 , \41460_41760 , \41461_41761 , \41462_41762 , \41463_41763 , \41464_41764 , \41465_41765 , \41466_41766 ,
         \41467_41767 , \41468_41768 , \41469_41769 , \41470_41770 , \41471_41771 , \41472_41772 , \41473_41773 , \41474_41774 , \41475_41775 , \41476_41776 ,
         \41477_41777 , \41478_41778 , \41479_41779 , \41480_41780 , \41481_41781 , \41482_41782 , \41483_41783 , \41484_41784 , \41485_41785 , \41486_41786 ,
         \41487_41787 , \41488_41788 , \41489_41789 , \41490_41790 , \41491_41791 , \41492_41792 , \41493_41793 , \41494_41794 , \41495_41795 , \41496_41796 ,
         \41497_41797 , \41498_41798 , \41499_41799 , \41500_41800 , \41501_41801 , \41502_41802 , \41503_41803 , \41504_41804 , \41505_41805 , \41506_41806 ,
         \41507_41807 , \41508_41808 , \41509_41809 , \41510_41810 , \41511_41811 , \41512_41812 , \41513_41813 , \41514_41814 , \41515_41815 , \41516_41816 ,
         \41517_41817 , \41518_41818 , \41519_41819 , \41520_41820 , \41521_41821 , \41522_41822 , \41523_41823 , \41524_41824 , \41525_41825 , \41526_41826 ,
         \41527_41827 , \41528_41828 , \41529_41829 , \41530_41830 , \41531_41831 , \41532_41832 , \41533_41833 , \41534_41834 , \41535_41835 , \41536_41836 ,
         \41537_41837 , \41538_41838 , \41539_41839 , \41540_41840 , \41541_41841 , \41542_41842 , \41543_41843 , \41544_41844 , \41545_41845 , \41546_41846 ,
         \41547_41847 , \41548_41848 , \41549_41849 , \41550_41850 , \41551_41851 , \41552_41852 , \41553_41853 , \41554_41854 , \41555_41855 , \41556_41856 ,
         \41557_41857 , \41558_41858 , \41559_41859 , \41560_41860 , \41561_41861 , \41562_41862 , \41563_41863 , \41564_41864 , \41565_41865 , \41566_41866 ,
         \41567_41867 , \41568_41868 , \41569_41869 , \41570_41870 , \41571_41871 , \41572_41872 , \41573_41873 , \41574_41874 , \41575_41875 , \41576_41876 ,
         \41577_41877 , \41578_41878 , \41579_41879 , \41580_41880 , \41581_41881 , \41582_41882 , \41583_41883 , \41584_41884 , \41585_41885 , \41586_41886 ,
         \41587_41887 , \41588_41888 , \41589_41889 , \41590_41890 , \41591_41891 , \41592_41892 , \41593_41893 , \41594_41894 , \41595_41895 , \41596_41896 ,
         \41597_41897 , \41598_41898 , \41599_41899 , \41600_41900 , \41601_41901 , \41602_41902 , \41603_41903 , \41604_41904 , \41605_41905 , \41606_41906 ,
         \41607_41907 , \41608_41908 , \41609_41909 , \41610_41910 , \41611_41911 , \41612_41912 , \41613_41913 , \41614_41914 , \41615_41915 , \41616_41916 ,
         \41617_41917 , \41618_41918 , \41619_41919 , \41620_41920 , \41621_41921 , \41622_41922 , \41623_41923 , \41624_41924 , \41625_41925 , \41626_41926 ,
         \41627_41927 , \41628_41928 , \41629_41929 , \41630_41930 , \41631_41931 , \41632_41932 , \41633_41933 , \41634_41934 , \41635_41935 , \41636_41936 ,
         \41637_41937 , \41638_41938 , \41639_41939 , \41640_41940 , \41641_41941 , \41642_41942 , \41643_41943 , \41644_41944 , \41645_41945 , \41646_41946 ,
         \41647_41947 , \41648_41948 , \41649_41949 , \41650_41950 , \41651_41951 , \41652_41952 , \41653_41953 , \41654_41954 , \41655_41955 , \41656_41956 ,
         \41657_41957 , \41658_41958 , \41659_41959 , \41660_41960 , \41661_41961 , \41662_41962 , \41663_41963_nG9b60 , \41664_41964 , \41665_41965 , \41666_41966 ,
         \41667_41967 , \41668_41968 , \41669_41969 , \41670_41970 , \41671_41971 , \41672_41972 , \41673_41973 , \41674_41974 , \41675_41975 , \41676_41976 ,
         \41677_41977 , \41678_41978 , \41679_41979 , \41680_41980 , \41681_41981 , \41682_41982 , \41683_41983 , \41684_41984 , \41685_41985 , \41686_41986 ,
         \41687_41987 , \41688_41988 , \41689_41989 , \41690_41990 , \41691_41991 , \41692_41992 , \41693_41993 , \41694_41994 , \41695_41995 , \41696_41996 ,
         \41697_41997 , \41698_41998 , \41699_41999 , \41700_42000 , \41701_42001 , \41702_42002 , \41703_42003 , \41704_42004 , \41705_42005 , \41706_42006 ,
         \41707_42007 , \41708_42008 , \41709_42009 , \41710_42010 , \41711_42011 , \41712_42012 , \41713_42013 , \41714_42014 , \41715_42015 , \41716_42016 ,
         \41717_42017 , \41718_42018 , \41719_42019 , \41720_42020 , \41721_42021 , \41722_42022 , \41723_42023 , \41724_42024 , \41725_42025 , \41726_42026 ,
         \41727_42027 , \41728_42028 , \41729_42029 , \41730_42030 , \41731_42031 , \41732_42032 , \41733_42033 , \41734_42034 , \41735_42035 , \41736_42036 ,
         \41737_42037 , \41738_42038 , \41739_42039 , \41740_42040 , \41741_42041 , \41742_42042 , \41743_42043 , \41744_42044 , \41745_42045 , \41746_42046 ,
         \41747_42047 , \41748_42048 , \41749_42049 , \41750_42050 , \41751_42051 , \41752_42052 , \41753_42053 , \41754_42054 , \41755_42055 , \41756_42056 ,
         \41757_42057 , \41758_42058 , \41759_42059 , \41760_42060 , \41761_42061 , \41762_42062 , \41763_42063 , \41764_42064 , \41765_42065 , \41766_42066 ,
         \41767_42067 , \41768_42068 , \41769_42069 , \41770_42070 , \41771_42071 , \41772_42072 , \41773_42073 , \41774_42074 , \41775_42075 , \41776_42076 ,
         \41777_42077 , \41778_42078 , \41779_42079 , \41780_42080 , \41781_42081 , \41782_42082 , \41783_42083 , \41784_42084 , \41785_42085 , \41786_42086 ,
         \41787_42087 , \41788_42088 , \41789_42089 , \41790_42090 , \41791_42091 , \41792_42092 , \41793_42093 , \41794_42094 , \41795_42095 , \41796_42096 ,
         \41797_42097 , \41798_42098 , \41799_42099 , \41800_42100 , \41801_42101 , \41802_42102 , \41803_42103 , \41804_42104 , \41805_42105 , \41806_42106 ,
         \41807_42107 , \41808_42108 , \41809_42109 , \41810_42110 , \41811_42111 , \41812_42112 , \41813_42113 , \41814_42114 , \41815_42115 , \41816_42116 ,
         \41817_42117 , \41818_42118 , \41819_42119 , \41820_42120 , \41821_42121 , \41822_42122 , \41823_42123 , \41824_42124 , \41825_42125 , \41826_42126 ,
         \41827_42127 , \41828_42128 , \41829_42129 , \41830_42130 , \41831_42131 , \41832_42132 , \41833_42133 , \41834_42134 , \41835_42135 , \41836_42136 ,
         \41837_42137 , \41838_42138 , \41839_42139 , \41840_42140 , \41841_42141 , \41842_42142 , \41843_42143 , \41844_42144 , \41845_42145 , \41846_42146 ,
         \41847_42147 , \41848_42148 , \41849_42149 , \41850_42150 , \41851_42151 , \41852_42152 , \41853_42153 , \41854_42154 , \41855_42155 , \41856_42156 ,
         \41857_42157 , \41858_42158 , \41859_42159 , \41860_42160 , \41861_42161 , \41862_42162 , \41863_42163 , \41864_42164 , \41865_42165 , \41866_42166 ,
         \41867_42167 , \41868_42168 , \41869_42169 , \41870_42170 , \41871_42171 , \41872_42172 , \41873_42173 , \41874_42174 , \41875_42175 , \41876_42176 ,
         \41877_42177 , \41878_42178 , \41879_42179 , \41880_42180 , \41881_42181 , \41882_42182 , \41883_42183 , \41884_42184 , \41885_42185 , \41886_42186 ,
         \41887_42187 , \41888_42188 , \41889_42189 , \41890_42190 , \41891_42191 , \41892_42192 , \41893_42193 , \41894_42194 , \41895_42195 , \41896_42196 ,
         \41897_42197 , \41898_42198 , \41899_42199 , \41900_42200 , \41901_42201_nG9b5d , \41902_42202 , \41903_42203 , \41904_42204 , \41905_42205 , \41906_42206 ,
         \41907_42207 , \41908_42208 , \41909_42209 , \41910_42210 , \41911_42211 , \41912_42212 , \41913_42213 , \41914_42214 , \41915_42215 , \41916_42216 ,
         \41917_42217 , \41918_42218 , \41919_42219 , \41920_42220 , \41921_42221 , \41922_42222 , \41923_42223 , \41924_42224 , \41925_42225 , \41926_42226 ,
         \41927_42227 , \41928_42228 , \41929_42229 , \41930_42230 , \41931_42231 , \41932_42232 , \41933_42233 , \41934_42234 , \41935_42235 , \41936_42236 ,
         \41937_42237 , \41938_42238 , \41939_42239 , \41940_42240 , \41941_42241 , \41942_42242 , \41943_42243 , \41944_42244 , \41945_42245 , \41946_42246 ,
         \41947_42247 , \41948_42248 , \41949_42249 , \41950_42250 , \41951_42251 , \41952_42252 , \41953_42253 , \41954_42254 , \41955_42255 , \41956_42256 ,
         \41957_42257 , \41958_42258 , \41959_42259 , \41960_42260 , \41961_42261 , \41962_42262 , \41963_42263 , \41964_42264 , \41965_42265 , \41966_42266 ,
         \41967_42267 , \41968_42268 , \41969_42269 , \41970_42270 , \41971_42271 , \41972_42272 , \41973_42273 , \41974_42274 , \41975_42275 , \41976_42276 ,
         \41977_42277 , \41978_42278 , \41979_42279 , \41980_42280 , \41981_42281 , \41982_42282 , \41983_42283 , \41984_42284 , \41985_42285 , \41986_42286 ,
         \41987_42287 , \41988_42288 , \41989_42289 , \41990_42290 , \41991_42291 , \41992_42292 , \41993_42293 , \41994_42294 , \41995_42295 , \41996_42296 ,
         \41997_42297 , \41998_42298 , \41999_42299 , \42000_42300 , \42001_42301 , \42002_42302 , \42003_42303 , \42004_42304 , \42005_42305 , \42006_42306 ,
         \42007_42307 , \42008_42308 , \42009_42309 , \42010_42310 , \42011_42311 , \42012_42312 , \42013_42313 , \42014_42314 , \42015_42315 , \42016_42316 ,
         \42017_42317 , \42018_42318 , \42019_42319 , \42020_42320 , \42021_42321 , \42022_42322 , \42023_42323 , \42024_42324 , \42025_42325 , \42026_42326 ,
         \42027_42327 , \42028_42328 , \42029_42329 , \42030_42330 , \42031_42331 , \42032_42332 , \42033_42333 , \42034_42334 , \42035_42335 , \42036_42336 ,
         \42037_42337 , \42038_42338 , \42039_42339 , \42040_42340 , \42041_42341 , \42042_42342 , \42043_42343 , \42044_42344 , \42045_42345 , \42046_42346 ,
         \42047_42347 , \42048_42348 , \42049_42349 , \42050_42350 , \42051_42351 , \42052_42352 , \42053_42353 , \42054_42354 , \42055_42355 , \42056_42356 ,
         \42057_42357 , \42058_42358 , \42059_42359 , \42060_42360 , \42061_42361 , \42062_42362 , \42063_42363 , \42064_42364 , \42065_42365 , \42066_42366 ,
         \42067_42367 , \42068_42368 , \42069_42369 , \42070_42370 , \42071_42371 , \42072_42372 , \42073_42373 , \42074_42374 , \42075_42375 , \42076_42376 ,
         \42077_42377 , \42078_42378 , \42079_42379 , \42080_42380 , \42081_42381 , \42082_42382 , \42083_42383 , \42084_42384 , \42085_42385 , \42086_42386 ,
         \42087_42387 , \42088_42388 , \42089_42389 , \42090_42390 , \42091_42391 , \42092_42392 , \42093_42393 , \42094_42394 , \42095_42395 , \42096_42396 ,
         \42097_42397 , \42098_42398 , \42099_42399 , \42100_42400 , \42101_42401 , \42102_42402 , \42103_42403 , \42104_42404 , \42105_42405 , \42106_42406 ,
         \42107_42407 , \42108_42408 , \42109_42409 , \42110_42410 , \42111_42411 , \42112_42412 , \42113_42413 , \42114_42414 , \42115_42415 , \42116_42416 ,
         \42117_42417 , \42118_42418 , \42119_42419 , \42120_42420 , \42121_42421 , \42122_42422 , \42123_42423 , \42124_42424 , \42125_42425 , \42126_42426 ,
         \42127_42427 , \42128_42428 , \42129_42429 , \42130_42430 , \42131_42431 , \42132_42432 , \42133_42433_nG9b5a , \42134_42434 , \42135_42435 , \42136_42436 ,
         \42137_42437 , \42138_42438 , \42139_42439 , \42140_42440 , \42141_42441 , \42142_42442 , \42143_42443 , \42144_42444 , \42145_42445 , \42146_42446 ,
         \42147_42447 , \42148_42448 , \42149_42449 , \42150_42450 , \42151_42451 , \42152_42452 , \42153_42453 , \42154_42454 , \42155_42455 , \42156_42456 ,
         \42157_42457 , \42158_42458 , \42159_42459 , \42160_42460 , \42161_42461 , \42162_42462 , \42163_42463 , \42164_42464 , \42165_42465 , \42166_42466 ,
         \42167_42467 , \42168_42468 , \42169_42469 , \42170_42470 , \42171_42471 , \42172_42472 , \42173_42473 , \42174_42474 , \42175_42475 , \42176_42476 ,
         \42177_42477 , \42178_42478 , \42179_42479 , \42180_42480 , \42181_42481 , \42182_42482 , \42183_42483 , \42184_42484 , \42185_42485 , \42186_42486 ,
         \42187_42487 , \42188_42488 , \42189_42489 , \42190_42490 , \42191_42491 , \42192_42492 , \42193_42493 , \42194_42494 , \42195_42495 , \42196_42496 ,
         \42197_42497 , \42198_42498 , \42199_42499 , \42200_42500 , \42201_42501 , \42202_42502 , \42203_42503 , \42204_42504 , \42205_42505 , \42206_42506 ,
         \42207_42507 , \42208_42508 , \42209_42509 , \42210_42510 , \42211_42511 , \42212_42512 , \42213_42513 , \42214_42514 , \42215_42515 , \42216_42516 ,
         \42217_42517 , \42218_42518 , \42219_42519 , \42220_42520 , \42221_42521 , \42222_42522 , \42223_42523 , \42224_42524 , \42225_42525 , \42226_42526 ,
         \42227_42527 , \42228_42528 , \42229_42529 , \42230_42530 , \42231_42531 , \42232_42532 , \42233_42533 , \42234_42534 , \42235_42535 , \42236_42536 ,
         \42237_42537 , \42238_42538 , \42239_42539 , \42240_42540 , \42241_42541 , \42242_42542 , \42243_42543 , \42244_42544 , \42245_42545 , \42246_42546 ,
         \42247_42547 , \42248_42548 , \42249_42549 , \42250_42550 , \42251_42551 , \42252_42552 , \42253_42553 , \42254_42554 , \42255_42555 , \42256_42556 ,
         \42257_42557 , \42258_42558 , \42259_42559 , \42260_42560 , \42261_42561 , \42262_42562 , \42263_42563 , \42264_42564 , \42265_42565 , \42266_42566 ,
         \42267_42567 , \42268_42568 , \42269_42569 , \42270_42570 , \42271_42571 , \42272_42572 , \42273_42573 , \42274_42574 , \42275_42575 , \42276_42576 ,
         \42277_42577 , \42278_42578 , \42279_42579 , \42280_42580 , \42281_42581 , \42282_42582 , \42283_42583 , \42284_42584 , \42285_42585 , \42286_42586 ,
         \42287_42587 , \42288_42588 , \42289_42589 , \42290_42590 , \42291_42591 , \42292_42592 , \42293_42593 , \42294_42594 , \42295_42595 , \42296_42596 ,
         \42297_42597 , \42298_42598 , \42299_42599 , \42300_42600 , \42301_42601 , \42302_42602 , \42303_42603 , \42304_42604 , \42305_42605 , \42306_42606 ,
         \42307_42607 , \42308_42608 , \42309_42609 , \42310_42610 , \42311_42611 , \42312_42612 , \42313_42613 , \42314_42614 , \42315_42615 , \42316_42616 ,
         \42317_42617 , \42318_42618 , \42319_42619 , \42320_42620 , \42321_42621 , \42322_42622 , \42323_42623 , \42324_42624 , \42325_42625 , \42326_42626 ,
         \42327_42627 , \42328_42628 , \42329_42629 , \42330_42630 , \42331_42631 , \42332_42632 , \42333_42633 , \42334_42634 , \42335_42635 , \42336_42636 ,
         \42337_42637 , \42338_42638 , \42339_42639 , \42340_42640 , \42341_42641 , \42342_42642 , \42343_42643 , \42344_42644 , \42345_42645 , \42346_42646 ,
         \42347_42647 , \42348_42648 , \42349_42649 , \42350_42650 , \42351_42651 , \42352_42652 , \42353_42653 , \42354_42654 , \42355_42655 , \42356_42656 ,
         \42357_42657 , \42358_42658 , \42359_42659 , \42360_42660 , \42361_42661 , \42362_42662 , \42363_42663 , \42364_42664 , \42365_42665 , \42366_42666 ,
         \42367_42667 , \42368_42668 , \42369_42669 , \42370_42670 , \42371_42671 , \42372_42672 , \42373_42673 , \42374_42674 , \42375_42675 , \42376_42676 ,
         \42377_42677 , \42378_42678 , \42379_42679 , \42380_42680 , \42381_42681 , \42382_42682 , \42383_42683 , \42384_42684 , \42385_42685 , \42386_42686 ,
         \42387_42687 , \42388_42688 , \42389_42689 , \42390_42690 , \42391_42691 , \42392_42692 , \42393_42693 , \42394_42694 , \42395_42695 , \42396_42696 ,
         \42397_42697 , \42398_42698 , \42399_42699 , \42400_42700 , \42401_42701 , \42402_42702 , \42403_42703 , \42404_42704 , \42405_42705 , \42406_42706 ,
         \42407_42707 , \42408_42708 , \42409_42709 , \42410_42710 , \42411_42711 , \42412_42712 , \42413_42713 , \42414_42714 , \42415_42715 , \42416_42716 ,
         \42417_42717 , \42418_42718 , \42419_42719 , \42420_42720 , \42421_42721 , \42422_42722 , \42423_42723 , \42424_42724 , \42425_42725 , \42426_42726 ,
         \42427_42727 , \42428_42728 , \42429_42729 , \42430_42730 , \42431_42731 , \42432_42732 , \42433_42733 , \42434_42734 , \42435_42735 , \42436_42736 ,
         \42437_42737 , \42438_42738 , \42439_42739 , \42440_42740 , \42441_42741 , \42442_42742 , \42443_42743 , \42444_42744 , \42445_42745 , \42446_42746 ,
         \42447_42747 , \42448_42748 , \42449_42749 , \42450_42750 , \42451_42751 , \42452_42752 , \42453_42753 , \42454_42754 , \42455_42755 , \42456_42756 ,
         \42457_42757 , \42458_42758 , \42459_42759 , \42460_42760 , \42461_42761 , \42462_42762 , \42463_42763 , \42464_42764 , \42465_42765 , \42466_42766_nG9b57 ,
         \42467_42767 , \42468_42768 , \42469_42769 , \42470_42770 , \42471_42771 , \42472_42772 , \42473_42773 , \42474_42774 , \42475_42775 , \42476_42776 ,
         \42477_42777 , \42478_42778 , \42479_42779 , \42480_42780 , \42481_42781 , \42482_42782 , \42483_42783 , \42484_42784 , \42485_42785 , \42486_42786 ,
         \42487_42787 , \42488_42788 , \42489_42789 , \42490_42790 , \42491_42791 , \42492_42792 , \42493_42793 , \42494_42794 , \42495_42795 , \42496_42796 ,
         \42497_42797 , \42498_42798 , \42499_42799 , \42500_42800 , \42501_42801 , \42502_42802 , \42503_42803 , \42504_42804 , \42505_42805 , \42506_42806 ,
         \42507_42807 , \42508_42808 , \42509_42809 , \42510_42810 , \42511_42811 , \42512_42812 , \42513_42813 , \42514_42814 , \42515_42815 , \42516_42816 ,
         \42517_42817 , \42518_42818 , \42519_42819 , \42520_42820 , \42521_42821 , \42522_42822 , \42523_42823 , \42524_42824 , \42525_42825 , \42526_42826 ,
         \42527_42827 , \42528_42828 , \42529_42829 , \42530_42830 , \42531_42831 , \42532_42832 , \42533_42833 , \42534_42834 , \42535_42835 , \42536_42836 ,
         \42537_42837 , \42538_42838 , \42539_42839 , \42540_42840 , \42541_42841 , \42542_42842 , \42543_42843 , \42544_42844 , \42545_42845 , \42546_42846 ,
         \42547_42847 , \42548_42848_nG9b54 , \42549_42849 , \42550_42850 , \42551_42851 , \42552_42852 , \42553_42853 , \42554_42854 , \42555_42855 , \42556_42856 ,
         \42557_42857 , \42558_42858 , \42559_42859 , \42560_42860 , \42561_42861 , \42562_42862 , \42563_42863 , \42564_42864 , \42565_42865 , \42566_42866 ,
         \42567_42867 , \42568_42868 , \42569_42869 , \42570_42870 , \42571_42871 , \42572_42872 , \42573_42873 , \42574_42874 , \42575_42875 , \42576_42876 ,
         \42577_42877 , \42578_42878 , \42579_42879 , \42580_42880 , \42581_42881 , \42582_42882 , \42583_42883 , \42584_42884 , \42585_42885 , \42586_42886 ,
         \42587_42887 , \42588_42888 , \42589_42889 , \42590_42890 , \42591_42891 , \42592_42892 , \42593_42893 , \42594_42894 , \42595_42895 , \42596_42896 ,
         \42597_42897 , \42598_42898 , \42599_42899 , \42600_42900 , \42601_42901 , \42602_42902 , \42603_42903 , \42604_42904 , \42605_42905 , \42606_42906 ,
         \42607_42907 , \42608_42908 , \42609_42909 , \42610_42910 , \42611_42911 , \42612_42912 , \42613_42913 , \42614_42914 , \42615_42915 , \42616_42916 ,
         \42617_42917 , \42618_42918 , \42619_42919 , \42620_42920 , \42621_42921 , \42622_42922 , \42623_42923 , \42624_42924 , \42625_42925 , \42626_42926 ,
         \42627_42927 , \42628_42928 , \42629_42929 , \42630_42930 , \42631_42931 , \42632_42932 , \42633_42933 , \42634_42934 , \42635_42935 , \42636_42936 ,
         \42637_42937 , \42638_42938 , \42639_42939 , \42640_42940 , \42641_42941 , \42642_42942 , \42643_42943 , \42644_42944 , \42645_42945 , \42646_42946 ,
         \42647_42947 , \42648_42948 , \42649_42949 , \42650_42950 , \42651_42951 , \42652_42952 , \42653_42953 , \42654_42954 , \42655_42955 , \42656_42956 ,
         \42657_42957 , \42658_42958 , \42659_42959 , \42660_42960 , \42661_42961 , \42662_42962 , \42663_42963 , \42664_42964 , \42665_42965 , \42666_42966 ,
         \42667_42967 , \42668_42968 , \42669_42969 , \42670_42970 , \42671_42971 , \42672_42972 , \42673_42973 , \42674_42974 , \42675_42975 , \42676_42976 ,
         \42677_42977 , \42678_42978 , \42679_42979 , \42680_42980 , \42681_42981 , \42682_42982 , \42683_42983 , \42684_42984 , \42685_42985 , \42686_42986 ,
         \42687_42987 , \42688_42988 , \42689_42989 , \42690_42990 , \42691_42991 , \42692_42992 , \42693_42993 , \42694_42994 , \42695_42995 , \42696_42996 ,
         \42697_42997 , \42698_42998 , \42699_42999 , \42700_43000 , \42701_43001 , \42702_43002 , \42703_43003 , \42704_43004 , \42705_43005 , \42706_43006 ,
         \42707_43007 , \42708_43008 , \42709_43009 , \42710_43010 , \42711_43011 , \42712_43012 , \42713_43013 , \42714_43014 , \42715_43015 , \42716_43016 ,
         \42717_43017 , \42718_43018 , \42719_43019 , \42720_43020 , \42721_43021 , \42722_43022 , \42723_43023 , \42724_43024 , \42725_43025 , \42726_43026 ,
         \42727_43027 , \42728_43028 , \42729_43029 , \42730_43030 , \42731_43031 , \42732_43032 , \42733_43033 , \42734_43034 , \42735_43035 , \42736_43036 ,
         \42737_43037 , \42738_43038 , \42739_43039 , \42740_43040 , \42741_43041 , \42742_43042 , \42743_43043 , \42744_43044 , \42745_43045 , \42746_43046 ,
         \42747_43047 , \42748_43048 , \42749_43049 , \42750_43050 , \42751_43051 , \42752_43052 , \42753_43053 , \42754_43054 , \42755_43055 , \42756_43056 ,
         \42757_43057 , \42758_43058 , \42759_43059 , \42760_43060 , \42761_43061 , \42762_43062 , \42763_43063 , \42764_43064 , \42765_43065 , \42766_43066 ,
         \42767_43067 , \42768_43068 , \42769_43069 , \42770_43070 , \42771_43071 , \42772_43072 , \42773_43073 , \42774_43074 , \42775_43075 , \42776_43076 ,
         \42777_43077 , \42778_43078 , \42779_43079 , \42780_43080 , \42781_43081 , \42782_43082 , \42783_43083 , \42784_43084 , \42785_43085 , \42786_43086 ,
         \42787_43087 , \42788_43088 , \42789_43089 , \42790_43090 , \42791_43091 , \42792_43092 , \42793_43093 , \42794_43094 , \42795_43095 , \42796_43096 ,
         \42797_43097 , \42798_43098 , \42799_43099 , \42800_43100 , \42801_43101 , \42802_43102 , \42803_43103 , \42804_43104 , \42805_43105 , \42806_43106 ,
         \42807_43107 , \42808_43108 , \42809_43109 , \42810_43110 , \42811_43111 , \42812_43112 , \42813_43113 , \42814_43114 , \42815_43115 , \42816_43116 ,
         \42817_43117 , \42818_43118 , \42819_43119 , \42820_43120 , \42821_43121 , \42822_43122 , \42823_43123 , \42824_43124 , \42825_43125 , \42826_43126 ,
         \42827_43127 , \42828_43128 , \42829_43129 , \42830_43130 , \42831_43131 , \42832_43132 , \42833_43133 , \42834_43134 , \42835_43135 , \42836_43136 ,
         \42837_43137 , \42838_43138 , \42839_43139 , \42840_43140 , \42841_43141 , \42842_43142 , \42843_43143 , \42844_43144 , \42845_43145 , \42846_43146 ,
         \42847_43147 , \42848_43148 , \42849_43149 , \42850_43150 , \42851_43151 , \42852_43152 , \42853_43153 , \42854_43154 , \42855_43155 , \42856_43156 ,
         \42857_43157 , \42858_43158 , \42859_43159 , \42860_43160 , \42861_43161 , \42862_43162 , \42863_43163 , \42864_43164 , \42865_43165 , \42866_43166 ,
         \42867_43167 , \42868_43168 , \42869_43169 , \42870_43170 , \42871_43171 , \42872_43172 , \42873_43173 , \42874_43174 , \42875_43175 , \42876_43176 ,
         \42877_43177 , \42878_43178 , \42879_43179_nG9b51 , \42880_43180 , \42881_43181 , \42882_43182 , \42883_43183 , \42884_43184 , \42885_43185 , \42886_43186 ,
         \42887_43187 , \42888_43188 , \42889_43189 , \42890_43190 , \42891_43191 , \42892_43192 , \42893_43193 , \42894_43194 , \42895_43195 , \42896_43196 ,
         \42897_43197 , \42898_43198 , \42899_43199 , \42900_43200 , \42901_43201 , \42902_43202 , \42903_43203 , \42904_43204 , \42905_43205 , \42906_43206 ,
         \42907_43207 , \42908_43208 , \42909_43209 , \42910_43210 , \42911_43211 , \42912_43212 , \42913_43213 , \42914_43214 , \42915_43215 , \42916_43216 ,
         \42917_43217 , \42918_43218 , \42919_43219 , \42920_43220 , \42921_43221 , \42922_43222 , \42923_43223 , \42924_43224 , \42925_43225 , \42926_43226 ,
         \42927_43227 , \42928_43228 , \42929_43229 , \42930_43230 , \42931_43231 , \42932_43232 , \42933_43233 , \42934_43234 , \42935_43235 , \42936_43236 ,
         \42937_43237 , \42938_43238 , \42939_43239 , \42940_43240 , \42941_43241 , \42942_43242 , \42943_43243 , \42944_43244 , \42945_43245 , \42946_43246 ,
         \42947_43247 , \42948_43248 , \42949_43249 , \42950_43250 , \42951_43251 , \42952_43252 , \42953_43253 , \42954_43254 , \42955_43255 , \42956_43256 ,
         \42957_43257 , \42958_43258 , \42959_43259 , \42960_43260 , \42961_43261 , \42962_43262 , \42963_43263 , \42964_43264 , \42965_43265 , \42966_43266 ,
         \42967_43267 , \42968_43268 , \42969_43269 , \42970_43270 , \42971_43271 , \42972_43272 , \42973_43273 , \42974_43274 , \42975_43275 , \42976_43276 ,
         \42977_43277 , \42978_43278 , \42979_43279 , \42980_43280 , \42981_43281 , \42982_43282 , \42983_43283 , \42984_43284 , \42985_43285 , \42986_43286 ,
         \42987_43287 , \42988_43288 , \42989_43289 , \42990_43290 , \42991_43291 , \42992_43292 , \42993_43293 , \42994_43294 , \42995_43295 , \42996_43296 ,
         \42997_43297 , \42998_43298 , \42999_43299 , \43000_43300 , \43001_43301 , \43002_43302 , \43003_43303 , \43004_43304 , \43005_43305 , \43006_43306 ,
         \43007_43307 , \43008_43308 , \43009_43309 , \43010_43310 , \43011_43311 , \43012_43312 , \43013_43313 , \43014_43314 , \43015_43315 , \43016_43316 ,
         \43017_43317 , \43018_43318 , \43019_43319 , \43020_43320 , \43021_43321 , \43022_43322 , \43023_43323 , \43024_43324 , \43025_43325 , \43026_43326 ,
         \43027_43327 , \43028_43328 , \43029_43329 , \43030_43330 , \43031_43331 , \43032_43332 , \43033_43333 , \43034_43334 , \43035_43335 , \43036_43336 ,
         \43037_43337 , \43038_43338 , \43039_43339 , \43040_43340 , \43041_43341 , \43042_43342 , \43043_43343 , \43044_43344 , \43045_43345 , \43046_43346 ,
         \43047_43347 , \43048_43348 , \43049_43349 , \43050_43350 , \43051_43351 , \43052_43352 , \43053_43353 , \43054_43354 , \43055_43355 , \43056_43356 ,
         \43057_43357 , \43058_43358 , \43059_43359 , \43060_43360 , \43061_43361 , \43062_43362 , \43063_43363 , \43064_43364 , \43065_43365 , \43066_43366 ,
         \43067_43367 , \43068_43368 , \43069_43369 , \43070_43370 , \43071_43371 , \43072_43372 , \43073_43373 , \43074_43374 , \43075_43375 , \43076_43376 ,
         \43077_43377 , \43078_43378 , \43079_43379 , \43080_43380 , \43081_43381 , \43082_43382 , \43083_43383 , \43084_43384 , \43085_43385 , \43086_43386 ,
         \43087_43387 , \43088_43388 , \43089_43389 , \43090_43390 , \43091_43391 , \43092_43392 , \43093_43393 , \43094_43394 , \43095_43395 , \43096_43396 ,
         \43097_43397 , \43098_43398 , \43099_43399 , \43100_43400 , \43101_43401 , \43102_43402 , \43103_43403 , \43104_43404 , \43105_43405 , \43106_43406 ,
         \43107_43407 , \43108_43408 , \43109_43409 , \43110_43410 , \43111_43411 , \43112_43412 , \43113_43413 , \43114_43414 , \43115_43415 , \43116_43416 ,
         \43117_43417 , \43118_43418 , \43119_43419 , \43120_43420 , \43121_43421 , \43122_43422 , \43123_43423 , \43124_43424 , \43125_43425 , \43126_43426 ,
         \43127_43427 , \43128_43428 , \43129_43429 , \43130_43430 , \43131_43431 , \43132_43432 , \43133_43433 , \43134_43434 , \43135_43435 , \43136_43436 ,
         \43137_43437 , \43138_43438 , \43139_43439 , \43140_43440 , \43141_43441 , \43142_43442 , \43143_43443 , \43144_43444 , \43145_43445 , \43146_43446 ,
         \43147_43447 , \43148_43448 , \43149_43449 , \43150_43450 , \43151_43451 , \43152_43452 , \43153_43453 , \43154_43454 , \43155_43455 , \43156_43456 ,
         \43157_43457 , \43158_43458 , \43159_43459 , \43160_43460 , \43161_43461 , \43162_43462 , \43163_43463 , \43164_43464 , \43165_43465 , \43166_43466 ,
         \43167_43467 , \43168_43468 , \43169_43469 , \43170_43470 , \43171_43471 , \43172_43472 , \43173_43473 , \43174_43474 , \43175_43475 , \43176_43476 ,
         \43177_43477 , \43178_43478 , \43179_43479 , \43180_43480 , \43181_43481 , \43182_43482 , \43183_43483 , \43184_43484 , \43185_43485 , \43186_43486 ,
         \43187_43487 , \43188_43488 , \43189_43489 , \43190_43490 , \43191_43491 , \43192_43492 , \43193_43493 , \43194_43494 , \43195_43495 , \43196_43496 ,
         \43197_43497 , \43198_43498 , \43199_43499 , \43200_43500 , \43201_43501 , \43202_43502 , \43203_43503 , \43204_43504 , \43205_43505 , \43206_43506 ,
         \43207_43507 , \43208_43508 , \43209_43509 , \43210_43510 , \43211_43511 , \43212_43512 , \43213_43513 , \43214_43514 , \43215_43515 , \43216_43516 ,
         \43217_43517 , \43218_43518 , \43219_43519 , \43220_43520 , \43221_43521 , \43222_43522 , \43223_43523 , \43224_43524 , \43225_43525 , \43226_43526 ,
         \43227_43527 , \43228_43528 , \43229_43529 , \43230_43530 , \43231_43531 , \43232_43532 , \43233_43533 , \43234_43534 , \43235_43535 , \43236_43536 ,
         \43237_43537 , \43238_43538 , \43239_43539 , \43240_43540 , \43241_43541 , \43242_43542 , \43243_43543 , \43244_43544 , \43245_43545 , \43246_43546 ,
         \43247_43547 , \43248_43548 , \43249_43549 , \43250_43550 , \43251_43551 , \43252_43552 , \43253_43553 , \43254_43554 , \43255_43555 , \43256_43556 ,
         \43257_43557 , \43258_43558 , \43259_43559 , \43260_43560 , \43261_43561 , \43262_43562 , \43263_43563 , \43264_43564 , \43265_43565 , \43266_43566 ,
         \43267_43567 , \43268_43568 , \43269_43569 , \43270_43570 , \43271_43571 , \43272_43572 , \43273_43573 , \43274_43574 , \43275_43575 , \43276_43576 ,
         \43277_43577 , \43278_43578 , \43279_43579 , \43280_43580 , \43281_43581 , \43282_43582 , \43283_43583 , \43284_43584 , \43285_43585 , \43286_43586 ,
         \43287_43587 , \43288_43588 , \43289_43589 , \43290_43590 , \43291_43591 , \43292_43592 , \43293_43593 , \43294_43594 , \43295_43595 , \43296_43596 ,
         \43297_43597 , \43298_43598 , \43299_43599 , \43300_43600 , \43301_43601 , \43302_43602 , \43303_43603 , \43304_43604 , \43305_43605 , \43306_43606 ,
         \43307_43607 , \43308_43608 , \43309_43609 , \43310_43610 , \43311_43611 , \43312_43612 , \43313_43613 , \43314_43614 , \43315_43615 , \43316_43616 ,
         \43317_43617 , \43318_43618 , \43319_43619 , \43320_43620 , \43321_43621 , \43322_43622 , \43323_43623 , \43324_43624 , \43325_43625 , \43326_43626 ,
         \43327_43627 , \43328_43628 , \43329_43629 , \43330_43630 , \43331_43631 , \43332_43632 , \43333_43633 , \43334_43634 , \43335_43635 , \43336_43636 ,
         \43337_43637 , \43338_43638 , \43339_43639 , \43340_43640 , \43341_43641 , \43342_43642 , \43343_43643 , \43344_43644 , \43345_43645 , \43346_43646 ,
         \43347_43647 , \43348_43648 , \43349_43649 , \43350_43650 , \43351_43651 , \43352_43652 , \43353_43653 , \43354_43654 , \43355_43655 , \43356_43656 ,
         \43357_43657 , \43358_43658 , \43359_43659 , \43360_43660 , \43361_43661 , \43362_43662 , \43363_43663 , \43364_43664 , \43365_43665 , \43366_43666 ,
         \43367_43667 , \43368_43668 , \43369_43669 , \43370_43670 , \43371_43671 , \43372_43672 , \43373_43673 , \43374_43674 , \43375_43675 , \43376_43676 ,
         \43377_43677 , \43378_43678 , \43379_43679 , \43380_43680 , \43381_43681 , \43382_43682 , \43383_43683 , \43384_43684 , \43385_43685 , \43386_43686 ,
         \43387_43687 , \43388_43688 , \43389_43689 , \43390_43690 , \43391_43691 , \43392_43692 , \43393_43693 , \43394_43694 , \43395_43695 , \43396_43696 ,
         \43397_43697 , \43398_43698 , \43399_43699 , \43400_43700 , \43401_43701 , \43402_43702 , \43403_43703 , \43404_43704 , \43405_43705 , \43406_43706 ,
         \43407_43707 , \43408_43708 , \43409_43709 , \43410_43710 , \43411_43711 , \43412_43712 , \43413_43713 , \43414_43714 , \43415_43715 , \43416_43716 ,
         \43417_43717 , \43418_43718 , \43419_43719 , \43420_43720 , \43421_43721 , \43422_43722 , \43423_43723 , \43424_43724 , \43425_43725 , \43426_43726 ,
         \43427_43727 , \43428_43728 , \43429_43729 , \43430_43730 , \43431_43731 , \43432_43732 , \43433_43733 , \43434_43734 , \43435_43735 , \43436_43736 ,
         \43437_43737 , \43438_43738 , \43439_43739 , \43440_43740 , \43441_43741 , \43442_43742 , \43443_43743 , \43444_43744 , \43445_43745 , \43446_43746 ,
         \43447_43747 , \43448_43748 , \43449_43749 , \43450_43750 , \43451_43751 , \43452_43752 , \43453_43753 , \43454_43754 , \43455_43755 , \43456_43756 ,
         \43457_43757 , \43458_43758 , \43459_43759 , \43460_43760 , \43461_43761 , \43462_43762 , \43463_43763 , \43464_43764 , \43465_43765 , \43466_43766 ,
         \43467_43767 , \43468_43768 , \43469_43769 , \43470_43770 , \43471_43771 , \43472_43772 , \43473_43773 , \43474_43774 , \43475_43775 , \43476_43776 ,
         \43477_43777 , \43478_43778 , \43479_43779 , \43480_43780 , \43481_43781 , \43482_43782 , \43483_43783 , \43484_43784 , \43485_43785 , \43486_43786 ,
         \43487_43787 , \43488_43788 , \43489_43789 , \43490_43790 , \43491_43791 , \43492_43792 , \43493_43793 , \43494_43794 , \43495_43795 , \43496_43796 ,
         \43497_43797 , \43498_43798 , \43499_43799 , \43500_43800 , \43501_43801 , \43502_43802 , \43503_43803 , \43504_43804 , \43505_43805 , \43506_43806 ,
         \43507_43807 , \43508_43808 , \43509_43809 , \43510_43810 , \43511_43811 , \43512_43812 , \43513_43813 , \43514_43814 , \43515_43815 , \43516_43816 ,
         \43517_43817 , \43518_43818 , \43519_43819 , \43520_43820 , \43521_43821 , \43522_43822 , \43523_43823 , \43524_43824 , \43525_43825 , \43526_43826 ,
         \43527_43827 , \43528_43828 , \43529_43829 , \43530_43830 , \43531_43831 , \43532_43832 , \43533_43833 , \43534_43834 , \43535_43835 , \43536_43836 ,
         \43537_43837 , \43538_43838 , \43539_43839 , \43540_43840 , \43541_43841 , \43542_43842 , \43543_43843 , \43544_43844 , \43545_43845 , \43546_43846 ,
         \43547_43847 , \43548_43848 , \43549_43849 , \43550_43850 , \43551_43851 , \43552_43852 , \43553_43853 , \43554_43854 , \43555_43855 , \43556_43856 ,
         \43557_43857 , \43558_43858 , \43559_43859 , \43560_43860 , \43561_43861 , \43562_43862 , \43563_43863 , \43564_43864 , \43565_43865 , \43566_43866 ,
         \43567_43867 , \43568_43868 , \43569_43869 , \43570_43870 , \43571_43871 , \43572_43872 , \43573_43873 , \43574_43874 , \43575_43875 , \43576_43876 ,
         \43577_43877 , \43578_43878 , \43579_43879 , \43580_43880 , \43581_43881 , \43582_43882 , \43583_43883 , \43584_43884 , \43585_43885 , \43586_43886 ,
         \43587_43887 , \43588_43888 , \43589_43889 , \43590_43890 , \43591_43891 , \43592_43892 , \43593_43893 , \43594_43894 , \43595_43895 , \43596_43896 ,
         \43597_43897 , \43598_43898 , \43599_43899 , \43600_43900 , \43601_43901 , \43602_43902 , \43603_43903 , \43604_43904 , \43605_43905 , \43606_43906 ,
         \43607_43907 , \43608_43908 , \43609_43909 , \43610_43910 , \43611_43911 , \43612_43912 , \43613_43913 , \43614_43914 , \43615_43915 , \43616_43916 ,
         \43617_43917 , \43618_43918 , \43619_43919 , \43620_43920 , \43621_43921 , \43622_43922 , \43623_43923 , \43624_43924 , \43625_43925 , \43626_43926 ,
         \43627_43927 , \43628_43928 , \43629_43929 , \43630_43930 , \43631_43931 , \43632_43932 , \43633_43933 , \43634_43934 , \43635_43935 , \43636_43936 ,
         \43637_43937 , \43638_43938 , \43639_43939 , \43640_43940 , \43641_43941 , \43642_43942 , \43643_43943 , \43644_43944 , \43645_43945 , \43646_43946 ,
         \43647_43947 , \43648_43948 , \43649_43949 , \43650_43950 , \43651_43951 , \43652_43952 , \43653_43953 , \43654_43954 , \43655_43955 , \43656_43956 ,
         \43657_43957 , \43658_43958 , \43659_43959 , \43660_43960 , \43661_43961 , \43662_43962 , \43663_43963 , \43664_43964 , \43665_43965 , \43666_43966 ,
         \43667_43967 , \43668_43968 , \43669_43969 , \43670_43970 , \43671_43971 , \43672_43972 , \43673_43973 , \43674_43974 , \43675_43975 , \43676_43976 ,
         \43677_43977 , \43678_43978 , \43679_43979 , \43680_43980 , \43681_43981 , \43682_43982 , \43683_43983 , \43684_43984 , \43685_43985 , \43686_43986 ,
         \43687_43987 , \43688_43988 , \43689_43989 , \43690_43990 , \43691_43991 , \43692_43992 , \43693_43993 , \43694_43994 , \43695_43995 , \43696_43996 ,
         \43697_43997 , \43698_43998 , \43699_43999 , \43700_44000 , \43701_44001 , \43702_44002 , \43703_44003 , \43704_44004 , \43705_44005 , \43706_44006 ,
         \43707_44007 , \43708_44008 , \43709_44009 , \43710_44010 , \43711_44011 , \43712_44012 , \43713_44013 , \43714_44014 , \43715_44015 , \43716_44016 ,
         \43717_44017 , \43718_44018 , \43719_44019 , \43720_44020 , \43721_44021 , \43722_44022 , \43723_44023 , \43724_44024 , \43725_44025 , \43726_44026 ,
         \43727_44027 , \43728_44028 , \43729_44029 , \43730_44030 , \43731_44031 , \43732_44032 , \43733_44033 , \43734_44034 , \43735_44035 , \43736_44036 ,
         \43737_44037 , \43738_44038 , \43739_44039 , \43740_44040 , \43741_44041 , \43742_44042 , \43743_44043 , \43744_44044 , \43745_44045 , \43746_44046 ,
         \43747_44047 , \43748_44048 , \43749_44049 , \43750_44050 , \43751_44051 , \43752_44052 , \43753_44053 , \43754_44054 , \43755_44055 , \43756_44056 ,
         \43757_44057 , \43758_44058 , \43759_44059 , \43760_44060 , \43761_44061 , \43762_44062 , \43763_44063 , \43764_44064 , \43765_44065 , \43766_44066 ,
         \43767_44067 , \43768_44068 , \43769_44069 , \43770_44070 , \43771_44071 , \43772_44072 , \43773_44073 , \43774_44074 , \43775_44075 , \43776_44076 ,
         \43777_44077 , \43778_44078 , \43779_44079 , \43780_44080 , \43781_44081 , \43782_44082 , \43783_44083 , \43784_44084 , \43785_44085 , \43786_44086 ,
         \43787_44087 , \43788_44088 , \43789_44089 , \43790_44090 , \43791_44091 , \43792_44092 , \43793_44093 , \43794_44094 , \43795_44095 , \43796_44096 ,
         \43797_44097 , \43798_44098 , \43799_44099 , \43800_44100 , \43801_44101 , \43802_44102 , \43803_44103 , \43804_44104 , \43805_44105 , \43806_44106 ,
         \43807_44107 , \43808_44108 , \43809_44109 , \43810_44110 , \43811_44111 , \43812_44112 , \43813_44113 , \43814_44114 , \43815_44115 , \43816_44116 ,
         \43817_44117 , \43818_44118 , \43819_44119 , \43820_44120 , \43821_44121 , \43822_44122 , \43823_44123 , \43824_44124 , \43825_44125 , \43826_44126 ,
         \43827_44127 , \43828_44128 , \43829_44129 , \43830_44130 , \43831_44131 , \43832_44132 , \43833_44133 , \43834_44134 , \43835_44135 , \43836_44136 ,
         \43837_44137 , \43838_44138 , \43839_44139 , \43840_44140 , \43841_44141 , \43842_44142 , \43843_44143 , \43844_44144 , \43845_44145 , \43846_44146 ,
         \43847_44147 , \43848_44148 , \43849_44149 , \43850_44150 , \43851_44151 , \43852_44152 , \43853_44153 , \43854_44154 , \43855_44155 , \43856_44156 ,
         \43857_44157 , \43858_44158 , \43859_44159 , \43860_44160 , \43861_44161 , \43862_44162 , \43863_44163 , \43864_44164 , \43865_44165 , \43866_44166 ,
         \43867_44167 , \43868_44168 , \43869_44169 , \43870_44170 , \43871_44171 , \43872_44172 , \43873_44173 , \43874_44174 , \43875_44175 , \43876_44176 ,
         \43877_44177 , \43878_44178 , \43879_44179 , \43880_44180 , \43881_44181 , \43882_44182 , \43883_44183 , \43884_44184 , \43885_44185 , \43886_44186 ,
         \43887_44187 , \43888_44188 , \43889_44189 , \43890_44190 , \43891_44191 , \43892_44192 , \43893_44193 , \43894_44194 , \43895_44195 , \43896_44196 ,
         \43897_44197 , \43898_44198 , \43899_44199 , \43900_44200 , \43901_44201 , \43902_44202 , \43903_44203 , \43904_44204 , \43905_44205 , \43906_44206 ,
         \43907_44207 , \43908_44208 , \43909_44209 , \43910_44210 , \43911_44211 , \43912_44212 , \43913_44213 , \43914_44214 , \43915_44215 , \43916_44216 ,
         \43917_44217 , \43918_44218 , \43919_44219 , \43920_44220 , \43921_44221 , \43922_44222 , \43923_44223 , \43924_44224 , \43925_44225 , \43926_44226 ,
         \43927_44227 , \43928_44228 , \43929_44229 , \43930_44230 , \43931_44231 , \43932_44232 , \43933_44233 , \43934_44234 , \43935_44235 , \43936_44236 ,
         \43937_44237 , \43938_44238 , \43939_44239 , \43940_44240 , \43941_44241 , \43942_44242 , \43943_44243 , \43944_44244 , \43945_44245 , \43946_44246 ,
         \43947_44247 , \43948_44248 , \43949_44249 , \43950_44250 , \43951_44251 , \43952_44252 , \43953_44253 , \43954_44254 , \43955_44255 , \43956_44256 ,
         \43957_44257 , \43958_44258 , \43959_44259 , \43960_44260 , \43961_44261 , \43962_44262 , \43963_44263 , \43964_44264 , \43965_44265 , \43966_44266 ,
         \43967_44267 , \43968_44268 , \43969_44269 , \43970_44270 , \43971_44271 , \43972_44272 , \43973_44273 , \43974_44274 , \43975_44275 , \43976_44276 ,
         \43977_44277 , \43978_44278 , \43979_44279 , \43980_44280 , \43981_44281 , \43982_44282 , \43983_44283 , \43984_44284 , \43985_44285 , \43986_44286 ,
         \43987_44287 , \43988_44288 , \43989_44289 , \43990_44290 , \43991_44291 , \43992_44292 , \43993_44293 , \43994_44294 , \43995_44295 , \43996_44296 ,
         \43997_44297 , \43998_44298 , \43999_44299 , \44000_44300 , \44001_44301 , \44002_44302 , \44003_44303 , \44004_44304 , \44005_44305 , \44006_44306 ,
         \44007_44307 , \44008_44308 , \44009_44309 , \44010_44310 , \44011_44311 , \44012_44312 , \44013_44313 , \44014_44314 , \44015_44315 , \44016_44316 ,
         \44017_44317 , \44018_44318 , \44019_44319 , \44020_44320 , \44021_44321 , \44022_44322 , \44023_44323 , \44024_44324 , \44025_44325 , \44026_44326 ,
         \44027_44327 , \44028_44328 , \44029_44329 , \44030_44330 , \44031_44331 , \44032_44332 , \44033_44333 , \44034_44334 , \44035_44335 , \44036_44336 ,
         \44037_44337 , \44038_44338 , \44039_44339 , \44040_44340 , \44041_44341 , \44042_44342 , \44043_44343 , \44044_44344 , \44045_44345 , \44046_44346 ,
         \44047_44347 , \44048_44348 , \44049_44349 , \44050_44350 , \44051_44351 , \44052_44352 , \44053_44353 , \44054_44354 , \44055_44355 , \44056_44356 ,
         \44057_44357 , \44058_44358 , \44059_44359 , \44060_44360 , \44061_44361 , \44062_44362 , \44063_44363 , \44064_44364 , \44065_44365 , \44066_44366 ,
         \44067_44367 , \44068_44368 , \44069_44369 , \44070_44370 , \44071_44371 , \44072_44372 , \44073_44373 , \44074_44374 , \44075_44375 , \44076_44376 ,
         \44077_44377 , \44078_44378 , \44079_44379 , \44080_44380 , \44081_44381 , \44082_44382 , \44083_44383 , \44084_44384 , \44085_44385 , \44086_44386 ,
         \44087_44387 , \44088_44388 , \44089_44389 , \44090_44390 , \44091_44391 , \44092_44392 , \44093_44393 , \44094_44394 , \44095_44395 , \44096_44396 ,
         \44097_44397 , \44098_44398 , \44099_44399 , \44100_44400 , \44101_44401 , \44102_44402 , \44103_44403 , \44104_44404 , \44105_44405 , \44106_44406 ,
         \44107_44407 , \44108_44408 , \44109_44409 , \44110_44410 , \44111_44411 , \44112_44412 , \44113_44413 , \44114_44414 , \44115_44415 , \44116_44416 ,
         \44117_44417 , \44118_44418 , \44119_44419 , \44120_44420 , \44121_44421 , \44122_44422 , \44123_44423 , \44124_44424 , \44125_44425 , \44126_44426 ,
         \44127_44427 , \44128_44428 , \44129_44429 , \44130_44430 , \44131_44431 , \44132_44432 , \44133_44433 , \44134_44434 , \44135_44435 , \44136_44436 ,
         \44137_44437 , \44138_44438 , \44139_44439 , \44140_44440 , \44141_44441 , \44142_44442 , \44143_44443 , \44144_44444 , \44145_44445 , \44146_44446 ,
         \44147_44447 , \44148_44448 , \44149_44449 , \44150_44450 , \44151_44451 , \44152_44452 , \44153_44453 , \44154_44454 , \44155_44455 , \44156_44456 ,
         \44157_44457 , \44158_44458 , \44159_44459 , \44160_44460 , \44161_44461 , \44162_44462 , \44163_44463 , \44164_44464 , \44165_44465 , \44166_44466 ,
         \44167_44467 , \44168_44468 , \44169_44469 , \44170_44470 , \44171_44471 , \44172_44472 , \44173_44473 , \44174_44474 , \44175_44475 , \44176_44476 ,
         \44177_44477 , \44178_44478 , \44179_44479 , \44180_44480 , \44181_44481 , \44182_44482 , \44183_44483 , \44184_44484 , \44185_44485 , \44186_44486 ,
         \44187_44487 , \44188_44488 , \44189_44489 , \44190_44490 , \44191_44491 , \44192_44492 , \44193_44493 , \44194_44494 , \44195_44495 , \44196_44496 ,
         \44197_44497 , \44198_44498 , \44199_44499 , \44200_44500 , \44201_44501 , \44202_44502 , \44203_44503 , \44204_44504 , \44205_44505 , \44206_44506 ,
         \44207_44507 , \44208_44508 , \44209_44509 , \44210_44510 , \44211_44511 , \44212_44512 , \44213_44513 , \44214_44514 , \44215_44515 , \44216_44516 ,
         \44217_44517 , \44218_44518 , \44219_44519 , \44220_44520 , \44221_44521 , \44222_44522 , \44223_44523 , \44224_44524 , \44225_44525 , \44226_44526 ,
         \44227_44527 , \44228_44528 , \44229_44529 , \44230_44530 , \44231_44531 , \44232_44532 , \44233_44533 , \44234_44534 , \44235_44535 , \44236_44536 ,
         \44237_44537 , \44238_44538 , \44239_44539 , \44240_44540 , \44241_44541 , \44242_44542 , \44243_44543 , \44244_44544 , \44245_44545 , \44246_44546 ,
         \44247_44547 , \44248_44548 , \44249_44549 , \44250_44550 , \44251_44551 , \44252_44552 , \44253_44553 , \44254_44554 , \44255_44555 , \44256_44556 ,
         \44257_44557 , \44258_44558 , \44259_44559 , \44260_44560 , \44261_44561 , \44262_44562 , \44263_44563 , \44264_44564 , \44265_44565 , \44266_44566 ,
         \44267_44567 , \44268_44568 , \44269_44569 , \44270_44570 , \44271_44571 , \44272_44572 , \44273_44573 , \44274_44574 , \44275_44575 , \44276_44576 ,
         \44277_44577 , \44278_44578 , \44279_44579 , \44280_44580 , \44281_44581 , \44282_44582 , \44283_44583 , \44284_44584 , \44285_44585 , \44286_44586 ,
         \44287_44587 , \44288_44588 , \44289_44589 , \44290_44590 , \44291_44591 , \44292_44592 , \44293_44593 , \44294_44594 , \44295_44595 , \44296_44596 ,
         \44297_44597 , \44298_44598 , \44299_44599 , \44300_44600 , \44301_44601 , \44302_44602 , \44303_44603 , \44304_44604 , \44305_44605 , \44306_44606 ,
         \44307_44607 , \44308_44608 , \44309_44609 , \44310_44610 , \44311_44611 , \44312_44612 , \44313_44613 , \44314_44614 , \44315_44615 , \44316_44616 ,
         \44317_44617 , \44318_44618 , \44319_44619 , \44320_44620 , \44321_44621 , \44322_44622 , \44323_44623 , \44324_44624 , \44325_44625 , \44326_44626 ,
         \44327_44627 , \44328_44628 , \44329_44629 , \44330_44630 , \44331_44631 , \44332_44632 , \44333_44633 , \44334_44634 , \44335_44635 , \44336_44636 ,
         \44337_44637 , \44338_44638 , \44339_44639 , \44340_44640 , \44341_44641 , \44342_44642 , \44343_44643 , \44344_44644 , \44345_44645 , \44346_44646 ,
         \44347_44647 , \44348_44648 , \44349_44649 , \44350_44650 , \44351_44651 , \44352_44652 , \44353_44653 , \44354_44654 , \44355_44655 , \44356_44656 ,
         \44357_44657 , \44358_44658 , \44359_44659 , \44360_44660 , \44361_44661 , \44362_44662 , \44363_44663 , \44364_44664 , \44365_44665 , \44366_44666 ,
         \44367_44667 , \44368_44668 , \44369_44669 , \44370_44670 , \44371_44671 , \44372_44672 , \44373_44673 , \44374_44674 , \44375_44675 , \44376_44676 ,
         \44377_44677 , \44378_44678 , \44379_44679 , \44380_44680 , \44381_44681 , \44382_44682 , \44383_44683 , \44384_44684 , \44385_44685 , \44386_44686 ,
         \44387_44687 , \44388_44688 , \44389_44689 , \44390_44690 , \44391_44691 , \44392_44692 , \44393_44693 , \44394_44694 , \44395_44695 , \44396_44696 ,
         \44397_44697 , \44398_44698 , \44399_44699 , \44400_44700 , \44401_44701 , \44402_44702 , \44403_44703 , \44404_44704 , \44405_44705 , \44406_44706 ,
         \44407_44707 , \44408_44708 , \44409_44709 , \44410_44710 , \44411_44711 , \44412_44712 , \44413_44713 , \44414_44714 , \44415_44715 , \44416_44716 ,
         \44417_44717 , \44418_44718 , \44419_44719 , \44420_44720 , \44421_44721 , \44422_44722 , \44423_44723 , \44424_44724 , \44425_44725 , \44426_44726 ,
         \44427_44727 , \44428_44728 , \44429_44729 , \44430_44730 , \44431_44731 , \44432_44732 , \44433_44733 , \44434_44734 , \44435_44735 , \44436_44736 ,
         \44437_44737 , \44438_44738 , \44439_44739 , \44440_44740 , \44441_44741 , \44442_44742 , \44443_44743 , \44444_44744 , \44445_44745 , \44446_44746 ,
         \44447_44747 , \44448_44748 , \44449_44749 , \44450_44750 , \44451_44751 , \44452_44752 , \44453_44753 , \44454_44754 , \44455_44755 , \44456_44756 ,
         \44457_44757 , \44458_44758 , \44459_44759 , \44460_44760 , \44461_44761 , \44462_44762 , \44463_44763 , \44464_44764 , \44465_44765 , \44466_44766 ,
         \44467_44767 , \44468_44768 , \44469_44769 , \44470_44770 , \44471_44771 , \44472_44772 , \44473_44773 , \44474_44774 , \44475_44775 , \44476_44776 ,
         \44477_44777 , \44478_44778 , \44479_44779 , \44480_44780 , \44481_44781 , \44482_44782 , \44483_44783 , \44484_44784 , \44485_44785 , \44486_44786 ,
         \44487_44787 , \44488_44788 , \44489_44789 , \44490_44790 , \44491_44791 , \44492_44792 , \44493_44793 , \44494_44794 , \44495_44795 , \44496_44796 ,
         \44497_44797 , \44498_44798 , \44499_44799 , \44500_44800 , \44501_44801 , \44502_44802 , \44503_44803 , \44504_44804 , \44505_44805 , \44506_44806 ,
         \44507_44807 , \44508_44808 , \44509_44809 , \44510_44810 , \44511_44811 , \44512_44812 , \44513_44813 , \44514_44814 , \44515_44815 , \44516_44816 ,
         \44517_44817 , \44518_44818 , \44519_44819 , \44520_44820 , \44521_44821 , \44522_44822 , \44523_44823 , \44524_44824 , \44525_44825 , \44526_44826 ,
         \44527_44827 , \44528_44828 , \44529_44829 , \44530_44830 , \44531_44831 , \44532_44832 , \44533_44833 , \44534_44834 , \44535_44835 , \44536_44836 ,
         \44537_44837 , \44538_44838 , \44539_44839 , \44540_44840 , \44541_44841 , \44542_44842 , \44543_44843 , \44544_44844 , \44545_44845 , \44546_44846 ,
         \44547_44847 , \44548_44848 , \44549_44849 , \44550_44850 , \44551_44851 , \44552_44852 , \44553_44853 , \44554_44854 , \44555_44855 , \44556_44856 ,
         \44557_44857 , \44558_44858 , \44559_44859 , \44560_44860 , \44561_44861 , \44562_44862 , \44563_44863 , \44564_44864 , \44565_44865 , \44566_44866 ,
         \44567_44867 , \44568_44868 , \44569_44869 , \44570_44870 , \44571_44871 , \44572_44872 , \44573_44873 , \44574_44874 , \44575_44875 , \44576_44876 ,
         \44577_44877 , \44578_44878 , \44579_44879 , \44580_44880 , \44581_44881 , \44582_44882 , \44583_44883 , \44584_44884 , \44585_44885 , \44586_44886 ,
         \44587_44887 , \44588_44888 , \44589_44889 , \44590_44890 , \44591_44891 , \44592_44892 , \44593_44893 , \44594_44894 , \44595_44895 , \44596_44896 ,
         \44597_44897 , \44598_44898 , \44599_44899 , \44600_44900 , \44601_44901 , \44602_44902 , \44603_44903 , \44604_44904 , \44605_44905 , \44606_44906 ,
         \44607_44907 , \44608_44908 , \44609_44909 , \44610_44910 , \44611_44911 , \44612_44912 , \44613_44913 , \44614_44914 , \44615_44915 , \44616_44916 ,
         \44617_44917 , \44618_44918 , \44619_44919 , \44620_44920 , \44621_44921 , \44622_44922 , \44623_44923 , \44624_44924 , \44625_44925 , \44626_44926 ,
         \44627_44927 , \44628_44928 , \44629_44929 , \44630_44930 , \44631_44931 , \44632_44932 , \44633_44933 , \44634_44934 , \44635_44935 , \44636_44936 ,
         \44637_44937 , \44638_44938 , \44639_44939 , \44640_44940 , \44641_44941 , \44642_44942 , \44643_44943 , \44644_44944 , \44645_44945 , \44646_44946 ,
         \44647_44947 , \44648_44948 , \44649_44949 , \44650_44950 , \44651_44951 , \44652_44952 , \44653_44953 , \44654_44954 , \44655_44955 , \44656_44956 ,
         \44657_44957 , \44658_44958 , \44659_44959 , \44660_44960 , \44661_44961 , \44662_44962 , \44663_44963 , \44664_44964 , \44665_44965 , \44666_44966 ,
         \44667_44967 , \44668_44968 , \44669_44969 , \44670_44970 , \44671_44971 , \44672_44972 , \44673_44973 , \44674_44974 , \44675_44975 , \44676_44976 ,
         \44677_44977 , \44678_44978 , \44679_44979 , \44680_44980 , \44681_44981 , \44682_44982 , \44683_44983 , \44684_44984 , \44685_44985 , \44686_44986 ,
         \44687_44987 , \44688_44988 , \44689_44989 , \44690_44990 , \44691_44991 , \44692_44992 , \44693_44993 , \44694_44994 , \44695_44995 , \44696_44996 ,
         \44697_44997 , \44698_44998 , \44699_44999 , \44700_45000 , \44701_45001 , \44702_45002 , \44703_45003 , \44704_45004 , \44705_45005 , \44706_45006 ,
         \44707_45007 , \44708_45008 , \44709_45009 , \44710_45010 , \44711_45011 , \44712_45012 , \44713_45013 , \44714_45014 , \44715_45015 , \44716_45016 ,
         \44717_45017 , \44718_45018 , \44719_45019 , \44720_45020 , \44721_45021 , \44722_45022 , \44723_45023 , \44724_45024 , \44725_45025 , \44726_45026 ,
         \44727_45027 , \44728_45028 , \44729_45029 , \44730_45030 , \44731_45031 , \44732_45032 , \44733_45033 , \44734_45034 , \44735_45035 , \44736_45036 ,
         \44737_45037 , \44738_45038 , \44739_45039 , \44740_45040 , \44741_45041 , \44742_45042 , \44743_45043 , \44744_45044 , \44745_45045 , \44746_45046 ,
         \44747_45047 , \44748_45048 , \44749_45049 , \44750_45050 , \44751_45051 , \44752_45052 , \44753_45053 , \44754_45054 , \44755_45055 , \44756_45056 ,
         \44757_45057 , \44758_45058 , \44759_45059 , \44760_45060 , \44761_45061 , \44762_45062 , \44763_45063 , \44764_45064 , \44765_45065 , \44766_45066 ,
         \44767_45067 , \44768_45068 , \44769_45069 , \44770_45070 , \44771_45071 , \44772_45072 , \44773_45073 , \44774_45074 , \44775_45075 , \44776_45076 ,
         \44777_45077 , \44778_45078 , \44779_45079 , \44780_45080 , \44781_45081 , \44782_45082 , \44783_45083 , \44784_45084 , \44785_45085 , \44786_45086 ,
         \44787_45087 , \44788_45088 , \44789_45089 , \44790_45090 , \44791_45091 , \44792_45092 , \44793_45093 , \44794_45094 , \44795_45095 , \44796_45096 ,
         \44797_45097 , \44798_45098 , \44799_45099 , \44800_45100 , \44801_45101 , \44802_45102 , \44803_45103 , \44804_45104 , \44805_45105 , \44806_45106 ,
         \44807_45107 , \44808_45108 , \44809_45109 , \44810_45110 , \44811_45111 , \44812_45112 , \44813_45113 , \44814_45114 , \44815_45115 , \44816_45116 ,
         \44817_45117 , \44818_45118 , \44819_45119 , \44820_45120 , \44821_45121 , \44822_45122 , \44823_45123 , \44824_45124 , \44825_45125 , \44826_45126 ,
         \44827_45127 , \44828_45128 , \44829_45129 , \44830_45130 , \44831_45131 , \44832_45132 , \44833_45133 , \44834_45134 , \44835_45135 , \44836_45136 ,
         \44837_45137 , \44838_45138 , \44839_45139 , \44840_45140 , \44841_45141 , \44842_45142 , \44843_45143 , \44844_45144 , \44845_45145 , \44846_45146 ,
         \44847_45147 , \44848_45148 , \44849_45149 , \44850_45150 , \44851_45151 , \44852_45152 , \44853_45153 , \44854_45154 , \44855_45155 , \44856_45156 ,
         \44857_45157 , \44858_45158 , \44859_45159 , \44860_45160 , \44861_45161 , \44862_45162 , \44863_45163 , \44864_45164 , \44865_45165 , \44866_45166 ,
         \44867_45167 , \44868_45168 , \44869_45169 , \44870_45170 , \44871_45171 , \44872_45172 , \44873_45173 , \44874_45174 , \44875_45175 , \44876_45176 ,
         \44877_45177 , \44878_45178 , \44879_45179 , \44880_45180 , \44881_45181 , \44882_45182 , \44883_45183 , \44884_45184 , \44885_45185 , \44886_45186 ,
         \44887_45187 , \44888_45188 , \44889_45189 , \44890_45190 , \44891_45191 , \44892_45192 , \44893_45193 , \44894_45194 , \44895_45195 , \44896_45196 ,
         \44897_45197 , \44898_45198 , \44899_45199 , \44900_45200 , \44901_45201 , \44902_45202 , \44903_45203 , \44904_45204 , \44905_45205 , \44906_45206 ,
         \44907_45207 , \44908_45208 , \44909_45209 , \44910_45210 , \44911_45211 , \44912_45212 , \44913_45213 , \44914_45214 , \44915_45215 , \44916_45216 ,
         \44917_45217 , \44918_45218 , \44919_45219 , \44920_45220 , \44921_45221 , \44922_45222 , \44923_45223 , \44924_45224 , \44925_45225 , \44926_45226 ,
         \44927_45227 , \44928_45228 , \44929_45229 , \44930_45230 , \44931_45231 , \44932_45232 , \44933_45233 , \44934_45234 , \44935_45235 , \44936_45236 ,
         \44937_45237 , \44938_45238 , \44939_45239 , \44940_45240 , \44941_45241 , \44942_45242 , \44943_45243 , \44944_45244 , \44945_45245 , \44946_45246 ,
         \44947_45247 , \44948_45248 , \44949_45249 , \44950_45250 , \44951_45251 , \44952_45252 , \44953_45253 , \44954_45254 , \44955_45255 , \44956_45256 ,
         \44957_45257 , \44958_45258 , \44959_45259 , \44960_45260 , \44961_45261 , \44962_45262 , \44963_45263 , \44964_45264 , \44965_45265 , \44966_45266 ,
         \44967_45267 , \44968_45268 , \44969_45269 , \44970_45270 , \44971_45271 , \44972_45272 , \44973_45273 , \44974_45274 , \44975_45275 , \44976_45276 ,
         \44977_45277 , \44978_45278 , \44979_45279 , \44980_45280 , \44981_45281 , \44982_45282 , \44983_45283 , \44984_45284 , \44985_45285 , \44986_45286 ,
         \44987_45287 , \44988_45288 , \44989_45289 , \44990_45290 , \44991_45291 , \44992_45292 , \44993_45293 , \44994_45294 , \44995_45295 , \44996_45296 ,
         \44997_45297 , \44998_45298 , \44999_45299 , \45000_45300 , \45001_45301 , \45002_45302 , \45003_45303 , \45004_45304 , \45005_45305 , \45006_45306 ,
         \45007_45307 , \45008_45308 , \45009_45309 , \45010_45310 , \45011_45311 , \45012_45312 , \45013_45313 , \45014_45314 , \45015_45315 , \45016_45316 ,
         \45017_45317 , \45018_45318 , \45019_45319 , \45020_45320 , \45021_45321 , \45022_45322 , \45023_45323 , \45024_45324 , \45025_45325 , \45026_45326 ,
         \45027_45327 , \45028_45328 , \45029_45329 , \45030_45330 , \45031_45331 , \45032_45332 , \45033_45333 , \45034_45334 , \45035_45335 , \45036_45336 ,
         \45037_45337 , \45038_45338 , \45039_45339 , \45040_45340 , \45041_45341 , \45042_45342 , \45043_45343 , \45044_45344 , \45045_45345 , \45046_45346 ,
         \45047_45347 , \45048_45348 , \45049_45349 , \45050_45350 , \45051_45351 , \45052_45352 , \45053_45353 , \45054_45354 , \45055_45355 , \45056_45356 ,
         \45057_45357 , \45058_45358 , \45059_45359 , \45060_45360 , \45061_45361 , \45062_45362 , \45063_45363 , \45064_45364 , \45065_45365 , \45066_45366 ,
         \45067_45367 , \45068_45368 , \45069_45369 , \45070_45370 , \45071_45371 , \45072_45372 , \45073_45373 , \45074_45374 , \45075_45375 , \45076_45376 ,
         \45077_45377 , \45078_45378 , \45079_45379 , \45080_45380 , \45081_45381 , \45082_45382 , \45083_45383 , \45084_45384 , \45085_45385 , \45086_45386 ,
         \45087_45387 , \45088_45388 , \45089_45389 , \45090_45390 , \45091_45391 , \45092_45392 , \45093_45393 , \45094_45394 , \45095_45395 , \45096_45396 ,
         \45097_45397 , \45098_45398 , \45099_45399 , \45100_45400 , \45101_45401 , \45102_45402 , \45103_45403 , \45104_45404 , \45105_45405 , \45106_45406 ,
         \45107_45407 , \45108_45408 , \45109_45409 , \45110_45410 , \45111_45411 , \45112_45412 , \45113_45413 , \45114_45414 , \45115_45415 , \45116_45416 ,
         \45117_45417 , \45118_45418 , \45119_45419 , \45120_45420 , \45121_45421 , \45122_45422 , \45123_45423 , \45124_45424 , \45125_45425 , \45126_45426 ,
         \45127_45427 , \45128_45428 , \45129_45429 , \45130_45430 , \45131_45431 , \45132_45432 , \45133_45433 , \45134_45434 , \45135_45435 , \45136_45436 ,
         \45137_45437 , \45138_45438 , \45139_45439 , \45140_45440 , \45141_45441 , \45142_45442 , \45143_45443 , \45144_45444 , \45145_45445 , \45146_45446 ,
         \45147_45447 , \45148_45448 , \45149_45449 , \45150_45450 , \45151_45451 , \45152_45452 , \45153_45453 , \45154_45454 , \45155_45455 , \45156_45456 ,
         \45157_45457 , \45158_45458 , \45159_45459 , \45160_45460 , \45161_45461 , \45162_45462 , \45163_45463 , \45164_45464 , \45165_45465 , \45166_45466 ,
         \45167_45467 , \45168_45468 , \45169_45469 , \45170_45470 , \45171_45471 , \45172_45472 , \45173_45473 , \45174_45474 , \45175_45475 , \45176_45476 ,
         \45177_45477 , \45178_45478 , \45179_45479 , \45180_45480 , \45181_45481 , \45182_45482 , \45183_45483 , \45184_45484 , \45185_45485 , \45186_45486 ,
         \45187_45487 , \45188_45488 , \45189_45489 , \45190_45490 , \45191_45491 , \45192_45492 , \45193_45493 , \45194_45494 , \45195_45495 , \45196_45496 ,
         \45197_45497 , \45198_45498 , \45199_45499 , \45200_45500 , \45201_45501 , \45202_45502 , \45203_45503 , \45204_45504 , \45205_45505 , \45206_45506 ,
         \45207_45507 , \45208_45508 , \45209_45509 , \45210_45510 , \45211_45511 , \45212_45512 , \45213_45513 , \45214_45514 , \45215_45515 , \45216_45516 ,
         \45217_45517 , \45218_45518 , \45219_45519 , \45220_45520 , \45221_45521 , \45222_45522 , \45223_45523 , \45224_45524 , \45225_45525 , \45226_45526 ,
         \45227_45527 , \45228_45528 , \45229_45529 , \45230_45530 , \45231_45531 , \45232_45532 , \45233_45533 , \45234_45534 , \45235_45535 , \45236_45536 ,
         \45237_45537 , \45238_45538 , \45239_45539 , \45240_45540 , \45241_45541 , \45242_45542 , \45243_45543 , \45244_45544 , \45245_45545 , \45246_45546 ,
         \45247_45547 , \45248_45548 , \45249_45549 , \45250_45550 , \45251_45551 , \45252_45552 , \45253_45553 , \45254_45554 , \45255_45555 , \45256_45556 ,
         \45257_45557 , \45258_45558 , \45259_45559 , \45260_45560 , \45261_45561 , \45262_45562 , \45263_45563 , \45264_45564 , \45265_45565 , \45266_45566 ,
         \45267_45567 , \45268_45568 , \45269_45569 , \45270_45570 , \45271_45571 , \45272_45572 , \45273_45573 , \45274_45574 , \45275_45575 , \45276_45576 ,
         \45277_45577 , \45278_45578 , \45279_45579 , \45280_45580 , \45281_45581 , \45282_45582 , \45283_45583 , \45284_45584 , \45285_45585 , \45286_45586 ,
         \45287_45587 , \45288_45588 , \45289_45589 , \45290_45590 , \45291_45591 , \45292_45592 , \45293_45593 , \45294_45594 , \45295_45595 , \45296_45596 ,
         \45297_45597 , \45298_45598 , \45299_45599 , \45300_45600 , \45301_45601 , \45302_45602 , \45303_45603 , \45304_45604 , \45305_45605 , \45306_45606 ,
         \45307_45607 , \45308_45608 , \45309_45609 , \45310_45610 , \45311_45611 , \45312_45612 , \45313_45613 , \45314_45614 , \45315_45615 , \45316_45616 ,
         \45317_45617 , \45318_45618 , \45319_45619 , \45320_45620 , \45321_45621 , \45322_45622 , \45323_45623 , \45324_45624 , \45325_45625 , \45326_45626 ,
         \45327_45627 , \45328_45628 , \45329_45629 , \45330_45630 , \45331_45631 , \45332_45632 , \45333_45633 , \45334_45634 , \45335_45635 , \45336_45636 ,
         \45337_45637 , \45338_45638 , \45339_45639 , \45340_45640 , \45341_45641 , \45342_45642 , \45343_45643 , \45344_45644 , \45345_45645 , \45346_45646 ,
         \45347_45647 , \45348_45648 , \45349_45649 , \45350_45650 , \45351_45651 , \45352_45652 , \45353_45653 , \45354_45654 , \45355_45655 , \45356_45656 ,
         \45357_45657 , \45358_45658 , \45359_45659 , \45360_45660 , \45361_45661 , \45362_45662 , \45363_45663 , \45364_45664 , \45365_45665 , \45366_45666 ,
         \45367_45667 , \45368_45668 , \45369_45669 , \45370_45670 , \45371_45671 , \45372_45672 , \45373_45673 , \45374_45674 , \45375_45675 , \45376_45676 ,
         \45377_45677 , \45378_45678 , \45379_45679 , \45380_45680 , \45381_45681 , \45382_45682 , \45383_45683 , \45384_45684 , \45385_45685 , \45386_45686 ,
         \45387_45687 , \45388_45688 , \45389_45689 , \45390_45690 , \45391_45691 , \45392_45692 , \45393_45693 , \45394_45694 , \45395_45695 , \45396_45696 ,
         \45397_45697 , \45398_45698 , \45399_45699 , \45400_45700 , \45401_45701 , \45402_45702 , \45403_45703 , \45404_45704 , \45405_45705 , \45406_45706 ,
         \45407_45707 , \45408_45708 , \45409_45709 , \45410_45710 , \45411_45711 , \45412_45712 , \45413_45713 , \45414_45714 , \45415_45715 , \45416_45716 ,
         \45417_45717 , \45418_45718 , \45419_45719 , \45420_45720 , \45421_45721 , \45422_45722 , \45423_45723 , \45424_45724 , \45425_45725 , \45426_45726 ,
         \45427_45727 , \45428_45728 , \45429_45729 , \45430_45730 , \45431_45731 , \45432_45732 , \45433_45733 , \45434_45734 , \45435_45735 , \45436_45736 ,
         \45437_45737 , \45438_45738 , \45439_45739 , \45440_45740 , \45441_45741 , \45442_45742 , \45443_45743 , \45444_45744 , \45445_45745 , \45446_45746 ,
         \45447_45747 , \45448_45748 , \45449_45749 , \45450_45750 , \45451_45751 , \45452_45752 , \45453_45753 , \45454_45754 , \45455_45755 , \45456_45756 ,
         \45457_45757 , \45458_45758 , \45459_45759 , \45460_45760 , \45461_45761 , \45462_45762 , \45463_45763 , \45464_45764 , \45465_45765 , \45466_45766 ,
         \45467_45767 , \45468_45768 , \45469_45769 , \45470_45770 , \45471_45771 , \45472_45772 , \45473_45773 , \45474_45774 , \45475_45775 , \45476_45776 ,
         \45477_45777 , \45478_45778 , \45479_45779 , \45480_45780 , \45481_45781 , \45482_45782 , \45483_45783 , \45484_45784 , \45485_45785 , \45486_45786 ,
         \45487_45787 , \45488_45788 , \45489_45789 , \45490_45790 , \45491_45791 , \45492_45792 , \45493_45793 , \45494_45794 , \45495_45795 , \45496_45796 ,
         \45497_45797 , \45498_45798 , \45499_45799 , \45500_45800 , \45501_45801 , \45502_45802 , \45503_45803 , \45504_45804 , \45505_45805 , \45506_45806 ,
         \45507_45807 , \45508_45808 , \45509_45809 , \45510_45810 , \45511_45811 , \45512_45812 , \45513_45813 , \45514_45814 , \45515_45815 , \45516_45816 ,
         \45517_45817 , \45518_45818 , \45519_45819 , \45520_45820 , \45521_45821 , \45522_45822 , \45523_45823 , \45524_45824 , \45525_45825 , \45526_45826 ,
         \45527_45827 , \45528_45828 , \45529_45829 , \45530_45830 , \45531_45831 , \45532_45832 , \45533_45833 , \45534_45834 , \45535_45835 , \45536_45836 ,
         \45537_45837 , \45538_45838 , \45539_45839 , \45540_45840 , \45541_45841 , \45542_45842 , \45543_45843 , \45544_45844 , \45545_45845 , \45546_45846 ,
         \45547_45847 , \45548_45848 , \45549_45849 , \45550_45850 , \45551_45851 , \45552_45852 , \45553_45853 , \45554_45854 , \45555_45855 , \45556_45856 ,
         \45557_45857 , \45558_45858 , \45559_45859 , \45560_45860 , \45561_45861 , \45562_45862 , \45563_45863 , \45564_45864 , \45565_45865 , \45566_45866 ,
         \45567_45867 , \45568_45868 , \45569_45869 , \45570_45870 , \45571_45871 , \45572_45872 , \45573_45873 , \45574_45874 , \45575_45875 , \45576_45876 ,
         \45577_45877 , \45578_45878 , \45579_45879 , \45580_45880 , \45581_45881 , \45582_45882 , \45583_45883 , \45584_45884 , \45585_45885 , \45586_45886 ,
         \45587_45887 , \45588_45888 , \45589_45889 , \45590_45890 , \45591_45891 , \45592_45892 , \45593_45893 , \45594_45894 , \45595_45895 , \45596_45896 ,
         \45597_45897 , \45598_45898 , \45599_45899 , \45600_45900 , \45601_45901 , \45602_45902 , \45603_45903 , \45604_45904 , \45605_45905 , \45606_45906 ,
         \45607_45907 , \45608_45908 , \45609_45909 , \45610_45910 , \45611_45911 , \45612_45912 , \45613_45913 , \45614_45914 , \45615_45915 , \45616_45916 ,
         \45617_45917 , \45618_45918 , \45619_45919 , \45620_45920 , \45621_45921 , \45622_45922 , \45623_45923 , \45624_45924 , \45625_45925 , \45626_45926 ,
         \45627_45927 , \45628_45928 , \45629_45929 , \45630_45930 , \45631_45931 , \45632_45932 , \45633_45933 , \45634_45934 , \45635_45935 , \45636_45936 ,
         \45637_45937 , \45638_45938 , \45639_45939 , \45640_45940 , \45641_45941 , \45642_45942 , \45643_45943 , \45644_45944 , \45645_45945 , \45646_45946 ,
         \45647_45947 , \45648_45948 , \45649_45949 , \45650_45950 , \45651_45951 , \45652_45952 , \45653_45953 , \45654_45954 , \45655_45955 , \45656_45956 ,
         \45657_45957 , \45658_45958 , \45659_45959 , \45660_45960 , \45661_45961 , \45662_45962 , \45663_45963 , \45664_45964 , \45665_45965 , \45666_45966 ,
         \45667_45967 , \45668_45968 , \45669_45969 , \45670_45970 , \45671_45971 , \45672_45972 , \45673_45973 , \45674_45974 , \45675_45975 , \45676_45976 ,
         \45677_45977 , \45678_45978 , \45679_45979 , \45680_45980 , \45681_45981 , \45682_45982 , \45683_45983 , \45684_45984 , \45685_45985 , \45686_45986 ,
         \45687_45987 , \45688_45988 , \45689_45989 , \45690_45990 , \45691_45991 , \45692_45992 , \45693_45993 , \45694_45994 , \45695_45995 , \45696_45996 ,
         \45697_45997 , \45698_45998 , \45699_45999 , \45700_46000 , \45701_46001 , \45702_46002 , \45703_46003 , \45704_46004 , \45705_46005 , \45706_46006 ,
         \45707_46007 , \45708_46008 , \45709_46009 , \45710_46010 , \45711_46011 , \45712_46012 , \45713_46013 , \45714_46014 , \45715_46015 , \45716_46016 ,
         \45717_46017 , \45718_46018 , \45719_46019 , \45720_46020 , \45721_46021 , \45722_46022 , \45723_46023 , \45724_46024 , \45725_46025 , \45726_46026 ,
         \45727_46027 , \45728_46028 , \45729_46029 , \45730_46030 , \45731_46031 , \45732_46032 , \45733_46033 , \45734_46034 , \45735_46035 , \45736_46036 ,
         \45737_46037 , \45738_46038 , \45739_46039 , \45740_46040 , \45741_46041 , \45742_46042 , \45743_46043 , \45744_46044 , \45745_46045 , \45746_46046 ,
         \45747_46047 , \45748_46048 , \45749_46049 , \45750_46050 , \45751_46051 , \45752_46052 , \45753_46053 , \45754_46054 , \45755_46055 , \45756_46056 ,
         \45757_46057 , \45758_46058 , \45759_46059 , \45760_46060 , \45761_46061 , \45762_46062 , \45763_46063 , \45764_46064 , \45765_46065 , \45766_46066 ,
         \45767_46067 , \45768_46068 , \45769_46069 , \45770_46070 , \45771_46071 , \45772_46072 , \45773_46073 , \45774_46074 , \45775_46075 , \45776_46076 ,
         \45777_46077 , \45778_46078 , \45779_46079 , \45780_46080 , \45781_46081 , \45782_46082 , \45783_46083 , \45784_46084 , \45785_46085 , \45786_46086 ,
         \45787_46087 , \45788_46088 , \45789_46089 , \45790_46090 , \45791_46091 , \45792_46092 , \45793_46093 , \45794_46094 , \45795_46095 , \45796_46096 ,
         \45797_46097 , \45798_46098 , \45799_46099 , \45800_46100 , \45801_46101 , \45802_46102 , \45803_46103 , \45804_46104 , \45805_46105 , \45806_46106 ,
         \45807_46107 , \45808_46108 , \45809_46109 , \45810_46110 , \45811_46111 , \45812_46112 , \45813_46113 , \45814_46114 , \45815_46115 , \45816_46116 ,
         \45817_46117 , \45818_46118 , \45819_46119 , \45820_46120 , \45821_46121 , \45822_46122 , \45823_46123 , \45824_46124 , \45825_46125 , \45826_46126 ,
         \45827_46127 , \45828_46128 , \45829_46129 , \45830_46130 , \45831_46131 , \45832_46132 , \45833_46133 , \45834_46134 , \45835_46135 , \45836_46136 ,
         \45837_46137 , \45838_46138 , \45839_46139 , \45840_46140 , \45841_46141 , \45842_46142 , \45843_46143 , \45844_46144 , \45845_46145 , \45846_46146 ,
         \45847_46147 , \45848_46148 , \45849_46149 , \45850_46150 , \45851_46151 , \45852_46152 , \45853_46153 , \45854_46154 , \45855_46155 , \45856_46156 ,
         \45857_46157 , \45858_46158 , \45859_46159 , \45860_46160 , \45861_46161 , \45862_46162 , \45863_46163 , \45864_46164 , \45865_46165 , \45866_46166 ,
         \45867_46167 , \45868_46168 , \45869_46169 , \45870_46170 , \45871_46171 , \45872_46172 , \45873_46173 , \45874_46174 , \45875_46175 , \45876_46176 ,
         \45877_46177 , \45878_46178 , \45879_46179 , \45880_46180 , \45881_46181 , \45882_46182 , \45883_46183 , \45884_46184 , \45885_46185 , \45886_46186 ,
         \45887_46187 , \45888_46188 , \45889_46189 , \45890_46190 , \45891_46191 , \45892_46192 , \45893_46193 , \45894_46194 , \45895_46195 , \45896_46196 ,
         \45897_46197 , \45898_46198 , \45899_46199 , \45900_46200 , \45901_46201 , \45902_46202 , \45903_46203 , \45904_46204 , \45905_46205 , \45906_46206 ,
         \45907_46207 , \45908_46208 , \45909_46209 , \45910_46210 , \45911_46211 , \45912_46212 , \45913_46213 , \45914_46214 , \45915_46215 , \45916_46216 ,
         \45917_46217 , \45918_46218 , \45919_46219 , \45920_46220 , \45921_46221 , \45922_46222 , \45923_46223 , \45924_46224 , \45925_46225 , \45926_46226 ,
         \45927_46227 , \45928_46228 , \45929_46229 , \45930_46230 , \45931_46231 , \45932_46232 , \45933_46233 , \45934_46234 , \45935_46235 , \45936_46236 ,
         \45937_46237 , \45938_46238 , \45939_46239 , \45940_46240 , \45941_46241 , \45942_46242 , \45943_46243 , \45944_46244 , \45945_46245 , \45946_46246 ,
         \45947_46247 , \45948_46248 , \45949_46249 , \45950_46250 , \45951_46251 , \45952_46252 , \45953_46253 , \45954_46254 , \45955_46255 , \45956_46256 ,
         \45957_46257 , \45958_46258 , \45959_46259 , \45960_46260 , \45961_46261 , \45962_46262 , \45963_46263 , \45964_46264 , \45965_46265 , \45966_46266 ,
         \45967_46267 , \45968_46268 , \45969_46269 , \45970_46270 , \45971_46271 , \45972_46272 , \45973_46273 , \45974_46274 , \45975_46275 , \45976_46276 ,
         \45977_46277 , \45978_46278 , \45979_46279 , \45980_46280 , \45981_46281 , \45982_46282 , \45983_46283 , \45984_46284 , \45985_46285 , \45986_46286 ,
         \45987_46287 , \45988_46288 , \45989_46289 , \45990_46290 , \45991_46291 , \45992_46292 , \45993_46293 , \45994_46294 , \45995_46295 , \45996_46296 ,
         \45997_46297 , \45998_46298 , \45999_46299 , \46000_46300 , \46001_46301 , \46002_46302 , \46003_46303 , \46004_46304 , \46005_46305 , \46006_46306 ,
         \46007_46307 , \46008_46308 , \46009_46309 , \46010_46310 , \46011_46311 , \46012_46312 , \46013_46313 , \46014_46314 , \46015_46315 , \46016_46316 ,
         \46017_46317 , \46018_46318 , \46019_46319 , \46020_46320 , \46021_46321 , \46022_46322 , \46023_46323 , \46024_46324 , \46025_46325 , \46026_46326 ,
         \46027_46327 , \46028_46328 , \46029_46329 , \46030_46330 , \46031_46331 , \46032_46332 , \46033_46333 , \46034_46334 , \46035_46335 , \46036_46336 ,
         \46037_46337 , \46038_46338 , \46039_46339 , \46040_46340 , \46041_46341 , \46042_46342 , \46043_46343 , \46044_46344 , \46045_46345 , \46046_46346 ,
         \46047_46347 , \46048_46348 , \46049_46349 , \46050_46350 , \46051_46351 , \46052_46352 , \46053_46353 , \46054_46354 , \46055_46355 , \46056_46356 ,
         \46057_46357 , \46058_46358 , \46059_46359 , \46060_46360 , \46061_46361 , \46062_46362 , \46063_46363 , \46064_46364 , \46065_46365 , \46066_46366 ,
         \46067_46367 , \46068_46368 , \46069_46369 , \46070_46370 , \46071_46371 , \46072_46372 , \46073_46373 , \46074_46374 , \46075_46375 , \46076_46376 ,
         \46077_46377 , \46078_46378 , \46079_46379 , \46080_46380 , \46081_46381 , \46082_46382 , \46083_46383 , \46084_46384 , \46085_46385 , \46086_46386 ,
         \46087_46387 , \46088_46388 , \46089_46389 , \46090_46390 , \46091_46391 , \46092_46392 , \46093_46393 , \46094_46394 , \46095_46395 , \46096_46396 ,
         \46097_46397 , \46098_46398 , \46099_46399 , \46100_46400 , \46101_46401 , \46102_46402 , \46103_46403 , \46104_46404 , \46105_46405 , \46106_46406 ,
         \46107_46407 , \46108_46408 , \46109_46409 , \46110_46410 , \46111_46411 , \46112_46412 , \46113_46413 , \46114_46414 , \46115_46415 , \46116_46416 ,
         \46117_46417 , \46118_46418 , \46119_46419 , \46120_46420 , \46121_46421 , \46122_46422 , \46123_46423 , \46124_46424 , \46125_46425 , \46126_46426 ,
         \46127_46427 , \46128_46428 , \46129_46429 , \46130_46430 , \46131_46431 , \46132_46432 , \46133_46433 , \46134_46434 , \46135_46435 , \46136_46436 ,
         \46137_46437 , \46138_46438 , \46139_46439 , \46140_46440 , \46141_46441 , \46142_46442 , \46143_46443 , \46144_46444 , \46145_46445 , \46146_46446 ,
         \46147_46447 , \46148_46448 , \46149_46449 , \46150_46450 , \46151_46451 , \46152_46452 , \46153_46453 , \46154_46454 , \46155_46455 , \46156_46456 ,
         \46157_46457 , \46158_46458 , \46159_46459 , \46160_46460 , \46161_46461 , \46162_46462 , \46163_46463 , \46164_46464 , \46165_46465 , \46166_46466 ,
         \46167_46467 , \46168_46468 , \46169_46469 , \46170_46470 , \46171_46471 , \46172_46472 , \46173_46473 , \46174_46474 , \46175_46475 , \46176_46476 ,
         \46177_46477 , \46178_46478 , \46179_46479 , \46180_46480 , \46181_46481 , \46182_46482 , \46183_46483 , \46184_46484 , \46185_46485 , \46186_46486 ,
         \46187_46487 , \46188_46488 , \46189_46489 , \46190_46490 , \46191_46491 , \46192_46492 , \46193_46493 , \46194_46494 , \46195_46495 , \46196_46496 ,
         \46197_46497 , \46198_46498 , \46199_46499 , \46200_46500 , \46201_46501 , \46202_46502 , \46203_46503 , \46204_46504 , \46205_46505 , \46206_46506 ,
         \46207_46507 , \46208_46508 , \46209_46509 , \46210_46510 , \46211_46511 , \46212_46512 , \46213_46513 , \46214_46514 , \46215_46515 , \46216_46516 ,
         \46217_46517 , \46218_46518 , \46219_46519 , \46220_46520 , \46221_46521 , \46222_46522 , \46223_46523 , \46224_46524 , \46225_46525 , \46226_46526 ,
         \46227_46527 , \46228_46528 , \46229_46529 , \46230_46530 , \46231_46531 , \46232_46532 , \46233_46533 , \46234_46534 , \46235_46535 , \46236_46536 ,
         \46237_46537 , \46238_46538 , \46239_46539 , \46240_46540 , \46241_46541 , \46242_46542 , \46243_46543 , \46244_46544 , \46245_46545 , \46246_46546 ,
         \46247_46547 , \46248_46548 , \46249_46549 , \46250_46550 , \46251_46551 , \46252_46552 , \46253_46553 , \46254_46554 , \46255_46555 , \46256_46556 ,
         \46257_46557 , \46258_46558 , \46259_46559 , \46260_46560 , \46261_46561 , \46262_46562 , \46263_46563 , \46264_46564 , \46265_46565 , \46266_46566 ,
         \46267_46567 , \46268_46568 , \46269_46569 , \46270_46570 , \46271_46571 , \46272_46572 , \46273_46573 , \46274_46574 , \46275_46575 , \46276_46576 ,
         \46277_46577 , \46278_46578 , \46279_46579 , \46280_46580 , \46281_46581 , \46282_46582 , \46283_46583 , \46284_46584 , \46285_46585 , \46286_46586 ,
         \46287_46587 , \46288_46588 , \46289_46589 , \46290_46590 , \46291_46591 , \46292_46592 , \46293_46593 , \46294_46594 , \46295_46595 , \46296_46596 ,
         \46297_46597 , \46298_46598 , \46299_46599 , \46300_46600 , \46301_46601 , \46302_46602 , \46303_46603 , \46304_46604 , \46305_46605 , \46306_46606 ,
         \46307_46607 , \46308_46608 , \46309_46609 , \46310_46610 , \46311_46611 , \46312_46612 , \46313_46613 , \46314_46614 , \46315_46615 , \46316_46616 ,
         \46317_46617 , \46318_46618 , \46319_46619 , \46320_46620 , \46321_46621 , \46322_46622 , \46323_46623 , \46324_46624 , \46325_46625 , \46326_46626 ,
         \46327_46627 , \46328_46628 , \46329_46629 , \46330_46630 , \46331_46631 , \46332_46632 , \46333_46633 , \46334_46634 , \46335_46635 , \46336_46636 ,
         \46337_46637 , \46338_46638 , \46339_46639 , \46340_46640 , \46341_46641 , \46342_46642 , \46343_46643 , \46344_46644 , \46345_46645 , \46346_46646 ,
         \46347_46647 , \46348_46648 , \46349_46649 , \46350_46650 , \46351_46651 , \46352_46652 , \46353_46653 , \46354_46654 , \46355_46655 , \46356_46656 ,
         \46357_46657 , \46358_46658 , \46359_46659 , \46360_46660 , \46361_46661 , \46362_46662 , \46363_46663 , \46364_46664 , \46365_46665 , \46366_46666 ,
         \46367_46667 , \46368_46668 , \46369_46669 , \46370_46670 , \46371_46671 , \46372_46672 , \46373_46673 , \46374_46674 , \46375_46675 , \46376_46676 ,
         \46377_46677 , \46378_46678 , \46379_46679 , \46380_46680 , \46381_46681 , \46382_46682 , \46383_46683 , \46384_46684 , \46385_46685 , \46386_46686 ,
         \46387_46687 , \46388_46688 , \46389_46689 , \46390_46690 , \46391_46691 , \46392_46692 , \46393_46693 , \46394_46694 , \46395_46695 , \46396_46696 ,
         \46397_46697 , \46398_46698 , \46399_46699 , \46400_46700 , \46401_46701 , \46402_46702 , \46403_46703 , \46404_46704 , \46405_46705 , \46406_46706 ,
         \46407_46707 , \46408_46708 , \46409_46709 , \46410_46710 , \46411_46711 , \46412_46712 , \46413_46713 , \46414_46714 , \46415_46715 , \46416_46716 ,
         \46417_46717 , \46418_46718 , \46419_46719 , \46420_46720 , \46421_46721 , \46422_46722 , \46423_46723 , \46424_46724 , \46425_46725 , \46426_46726 ,
         \46427_46727 , \46428_46728 , \46429_46729 , \46430_46730 , \46431_46731 , \46432_46732 , \46433_46733 , \46434_46734 , \46435_46735 , \46436_46736 ,
         \46437_46737 , \46438_46738 , \46439_46739 , \46440_46740 , \46441_46741 , \46442_46742 , \46443_46743 , \46444_46744 , \46445_46745 , \46446_46746 ,
         \46447_46747 , \46448_46748 , \46449_46749 , \46450_46750 , \46451_46751 , \46452_46752 , \46453_46753 , \46454_46754 , \46455_46755 , \46456_46756 ,
         \46457_46757 , \46458_46758 , \46459_46759 , \46460_46760 , \46461_46761 , \46462_46762 , \46463_46763 , \46464_46764 , \46465_46765 , \46466_46766 ,
         \46467_46767 , \46468_46768 , \46469_46769 , \46470_46770 , \46471_46771 , \46472_46772 , \46473_46773 , \46474_46774 , \46475_46775 , \46476_46776 ,
         \46477_46777 , \46478_46778 , \46479_46779 , \46480_46780 , \46481_46781 , \46482_46782 , \46483_46783 , \46484_46784 , \46485_46785 , \46486_46786 ,
         \46487_46787 , \46488_46788 , \46489_46789 , \46490_46790 , \46491_46791 , \46492_46792 , \46493_46793 , \46494_46794 , \46495_46795 , \46496_46796 ,
         \46497_46797 , \46498_46798 , \46499_46799 , \46500_46800 , \46501_46801 , \46502_46802 , \46503_46803 , \46504_46804 , \46505_46805 , \46506_46806 ,
         \46507_46807 , \46508_46808 , \46509_46809 , \46510_46810 , \46511_46811 , \46512_46812 , \46513_46813 , \46514_46814 , \46515_46815 , \46516_46816 ,
         \46517_46817 , \46518_46818 , \46519_46819 , \46520_46820 , \46521_46821 , \46522_46822 , \46523_46823 , \46524_46824 , \46525_46825 , \46526_46826 ,
         \46527_46827 , \46528_46828 , \46529_46829 , \46530_46830 , \46531_46831 , \46532_46832 , \46533_46833 , \46534_46834 , \46535_46835 , \46536_46836 ,
         \46537_46837 , \46538_46838 , \46539_46839 , \46540_46840 , \46541_46841 , \46542_46842 , \46543_46843 , \46544_46844 , \46545_46845 , \46546_46846 ,
         \46547_46847 , \46548_46848 , \46549_46849 , \46550_46850 , \46551_46851 , \46552_46852 , \46553_46853 , \46554_46854 , \46555_46855 , \46556_46856 ,
         \46557_46857 , \46558_46858 , \46559_46859 , \46560_46860 , \46561_46861 , \46562_46862 , \46563_46863 , \46564_46864 , \46565_46865 , \46566_46866 ,
         \46567_46867 , \46568_46868 , \46569_46869 , \46570_46870 , \46571_46871 , \46572_46872 , \46573_46873 , \46574_46874 , \46575_46875 , \46576_46876 ,
         \46577_46877 , \46578_46878 , \46579_46879 , \46580_46880 , \46581_46881 , \46582_46882 , \46583_46883 , \46584_46884 , \46585_46885 , \46586_46886 ,
         \46587_46887 , \46588_46888 , \46589_46889 , \46590_46890 , \46591_46891 , \46592_46892 , \46593_46893 , \46594_46894 , \46595_46895 , \46596_46896 ,
         \46597_46897 , \46598_46898 , \46599_46899 , \46600_46900 , \46601_46901 , \46602_46902 , \46603_46903 , \46604_46904 , \46605_46905 , \46606_46906 ,
         \46607_46907 , \46608_46908 , \46609_46909 , \46610_46910 , \46611_46911 , \46612_46912 , \46613_46913 , \46614_46914 , \46615_46915 , \46616_46916 ,
         \46617_46917 , \46618_46918 , \46619_46919 , \46620_46920 , \46621_46921 , \46622_46922 , \46623_46923 , \46624_46924 , \46625_46925 , \46626_46926 ,
         \46627_46927 , \46628_46928 , \46629_46929 , \46630_46930 , \46631_46931 , \46632_46932 , \46633_46933 , \46634_46934 , \46635_46935 , \46636_46936 ,
         \46637_46937 , \46638_46938 , \46639_46939 , \46640_46940 , \46641_46941 , \46642_46942 , \46643_46943 , \46644_46944 , \46645_46945 , \46646_46946 ,
         \46647_46947 , \46648_46948 , \46649_46949 , \46650_46950 , \46651_46951 , \46652_46952 , \46653_46953 , \46654_46954 , \46655_46955 , \46656_46956 ,
         \46657_46957 , \46658_46958 , \46659_46959 , \46660_46960 , \46661_46961 , \46662_46962 , \46663_46963 , \46664_46964 , \46665_46965 , \46666_46966 ,
         \46667_46967 , \46668_46968 , \46669_46969 , \46670_46970 , \46671_46971 , \46672_46972 , \46673_46973 , \46674_46974 , \46675_46975 , \46676_46976 ,
         \46677_46977 , \46678_46978 , \46679_46979 , \46680_46980 , \46681_46981 , \46682_46982 , \46683_46983 , \46684_46984 , \46685_46985 , \46686_46986 ,
         \46687_46987 , \46688_46988 , \46689_46989 , \46690_46990 , \46691_46991 , \46692_46992 , \46693_46993 , \46694_46994 , \46695_46995 , \46696_46996 ,
         \46697_46997 , \46698_46998 , \46699_46999 , \46700_47000 , \46701_47001 , \46702_47002 , \46703_47003 , \46704_47004 , \46705_47005 , \46706_47006 ,
         \46707_47007 , \46708_47008 , \46709_47009 , \46710_47010 , \46711_47011 , \46712_47012 , \46713_47013 , \46714_47014 , \46715_47015 , \46716_47016 ,
         \46717_47017 , \46718_47018 , \46719_47019 , \46720_47020 , \46721_47021 , \46722_47022 , \46723_47023 , \46724_47024 , \46725_47025 , \46726_47026 ,
         \46727_47027 , \46728_47028 , \46729_47029 , \46730_47030 , \46731_47031 , \46732_47032 , \46733_47033 , \46734_47034 , \46735_47035 , \46736_47036 ,
         \46737_47037 , \46738_47038 , \46739_47039 , \46740_47040 , \46741_47041 , \46742_47042 , \46743_47043 , \46744_47044 , \46745_47045 , \46746_47046 ,
         \46747_47047 , \46748_47048 , \46749_47049 , \46750_47050 , \46751_47051 , \46752_47052 , \46753_47053 , \46754_47054 , \46755_47055 , \46756_47056 ,
         \46757_47057 , \46758_47058 , \46759_47059 , \46760_47060 , \46761_47061 , \46762_47062 , \46763_47063 , \46764_47064 , \46765_47065 , \46766_47066 ,
         \46767_47067 , \46768_47068 , \46769_47069 , \46770_47070 , \46771_47071 , \46772_47072 , \46773_47073 , \46774_47074 , \46775_47075 , \46776_47076 ,
         \46777_47077 , \46778_47078 , \46779_47079 , \46780_47080 , \46781_47081 , \46782_47082 , \46783_47083 , \46784_47084 , \46785_47085 , \46786_47086 ,
         \46787_47087 , \46788_47088 , \46789_47089 , \46790_47090 , \46791_47091 , \46792_47092 , \46793_47093 , \46794_47094 , \46795_47095 , \46796_47096 ,
         \46797_47097 , \46798_47098 , \46799_47099 , \46800_47100 , \46801_47101 , \46802_47102 , \46803_47103 , \46804_47104 , \46805_47105 , \46806_47106 ,
         \46807_47107 , \46808_47108 , \46809_47109 , \46810_47110 , \46811_47111 , \46812_47112 , \46813_47113 , \46814_47114 , \46815_47115 , \46816_47116 ,
         \46817_47117 , \46818_47118 , \46819_47119 , \46820_47120 , \46821_47121 , \46822_47122 , \46823_47123 , \46824_47124 , \46825_47125 , \46826_47126 ,
         \46827_47127 , \46828_47128 , \46829_47129 , \46830_47130 , \46831_47131 , \46832_47132 , \46833_47133 , \46834_47134 , \46835_47135 , \46836_47136 ,
         \46837_47137 , \46838_47138 , \46839_47139 , \46840_47140 , \46841_47141 , \46842_47142 , \46843_47143 , \46844_47144 , \46845_47145 , \46846_47146 ,
         \46847_47147 , \46848_47148 , \46849_47149 , \46850_47150 , \46851_47151 , \46852_47152 , \46853_47153 , \46854_47154 , \46855_47155 , \46856_47156 ,
         \46857_47157 , \46858_47158 , \46859_47159 , \46860_47160 , \46861_47161 , \46862_47162 , \46863_47163 , \46864_47164 , \46865_47165 , \46866_47166 ,
         \46867_47167 , \46868_47168 , \46869_47169 , \46870_47170 , \46871_47171 , \46872_47172 , \46873_47173 , \46874_47174 , \46875_47175 , \46876_47176 ,
         \46877_47177 , \46878_47178 , \46879_47179 , \46880_47180 , \46881_47181 , \46882_47182 , \46883_47183 , \46884_47184 , \46885_47185 , \46886_47186 ,
         \46887_47187 , \46888_47188 , \46889_47189 , \46890_47190 , \46891_47191 , \46892_47192 , \46893_47193 , \46894_47194 , \46895_47195 , \46896_47196 ,
         \46897_47197 , \46898_47198 , \46899_47199 , \46900_47200 , \46901_47201 , \46902_47202 , \46903_47203 , \46904_47204 , \46905_47205 , \46906_47206 ,
         \46907_47207 , \46908_47208 , \46909_47209 , \46910_47210 , \46911_47211 , \46912_47212 , \46913_47213 , \46914_47214 , \46915_47215 , \46916_47216 ,
         \46917_47217 , \46918_47218 , \46919_47219 , \46920_47220 , \46921_47221 , \46922_47222 , \46923_47223 , \46924_47224 , \46925_47225 , \46926_47226 ,
         \46927_47227 , \46928_47228 , \46929_47229 , \46930_47230 , \46931_47231 , \46932_47232 , \46933_47233 , \46934_47234 , \46935_47235 , \46936_47236 ,
         \46937_47237 , \46938_47238 , \46939_47239 , \46940_47240 , \46941_47241 , \46942_47242 , \46943_47243 , \46944_47244 , \46945_47245 , \46946_47246 ,
         \46947_47247 , \46948_47248 , \46949_47249 , \46950_47250 , \46951_47251 , \46952_47252 , \46953_47253 , \46954_47254 , \46955_47255 , \46956_47256 ,
         \46957_47257 , \46958_47258 , \46959_47259 , \46960_47260 , \46961_47261 , \46962_47262 , \46963_47263 , \46964_47264 , \46965_47265 , \46966_47266 ,
         \46967_47267 , \46968_47268 , \46969_47269 , \46970_47270 , \46971_47271 , \46972_47272 , \46973_47273 , \46974_47274 , \46975_47275 , \46976_47276 ,
         \46977_47277 , \46978_47278 , \46979_47279 , \46980_47280 , \46981_47281 , \46982_47282 , \46983_47283 , \46984_47284 , \46985_47285 , \46986_47286 ,
         \46987_47287 , \46988_47288 , \46989_47289 , \46990_47290 , \46991_47291 , \46992_47292 , \46993_47293 , \46994_47294 , \46995_47295 , \46996_47296 ,
         \46997_47297 , \46998_47298 , \46999_47299 , \47000_47300 , \47001_47301 , \47002_47302 , \47003_47303 , \47004_47304 , \47005_47305 , \47006_47306 ,
         \47007_47307 , \47008_47308 , \47009_47309 , \47010_47310 , \47011_47311 , \47012_47312 , \47013_47313 , \47014_47314 , \47015_47315 , \47016_47316 ,
         \47017_47317 , \47018_47318 , \47019_47319 , \47020_47320 , \47021_47321 , \47022_47322 , \47023_47323 , \47024_47324 , \47025_47325 , \47026_47326 ,
         \47027_47327 , \47028_47328 , \47029_47329 , \47030_47330 , \47031_47331 , \47032_47332 , \47033_47333 , \47034_47334 , \47035_47335 , \47036_47336 ,
         \47037_47337 , \47038_47338 , \47039_47339 , \47040_47340 , \47041_47341 , \47042_47342 , \47043_47343 , \47044_47344 , \47045_47345 , \47046_47346 ,
         \47047_47347 , \47048_47348 , \47049_47349 , \47050_47350 , \47051_47351 , \47052_47352 , \47053_47353 , \47054_47354 , \47055_47355 , \47056_47356 ,
         \47057_47357 , \47058_47358 , \47059_47359 , \47060_47360 , \47061_47361 , \47062_47362 , \47063_47363 , \47064_47364 , \47065_47365 , \47066_47366 ,
         \47067_47367 , \47068_47368 , \47069_47369 , \47070_47370 , \47071_47371 , \47072_47372 , \47073_47373 , \47074_47374 , \47075_47375 , \47076_47376 ,
         \47077_47377 , \47078_47378 , \47079_47379 , \47080_47380 , \47081_47381 , \47082_47382 , \47083_47383 , \47084_47384 , \47085_47385 , \47086_47386 ,
         \47087_47387 , \47088_47388 , \47089_47389 , \47090_47390 , \47091_47391 , \47092_47392 , \47093_47393 , \47094_47394 , \47095_47395 , \47096_47396 ,
         \47097_47397 , \47098_47398 , \47099_47399 , \47100_47400 , \47101_47401 , \47102_47402 , \47103_47403 , \47104_47404 , \47105_47405 , \47106_47406 ,
         \47107_47407 , \47108_47408 , \47109_47409 , \47110_47410 , \47111_47411 , \47112_47412 , \47113_47413 , \47114_47414 , \47115_47415 , \47116_47416 ,
         \47117_47417 , \47118_47418 , \47119_47419 , \47120_47420 , \47121_47421 , \47122_47422 , \47123_47423 , \47124_47424 , \47125_47425 , \47126_47426 ,
         \47127_47427 , \47128_47428 , \47129_47429 , \47130_47430 , \47131_47431 , \47132_47432 , \47133_47433 , \47134_47434 , \47135_47435 , \47136_47436 ,
         \47137_47437 , \47138_47438 , \47139_47439 , \47140_47440 , \47141_47441 , \47142_47442 , \47143_47443 , \47144_47444 , \47145_47445 , \47146_47446 ,
         \47147_47447 , \47148_47448 , \47149_47449 , \47150_47450 , \47151_47451 , \47152_47452 , \47153_47453 , \47154_47454 , \47155_47455 , \47156_47456 ,
         \47157_47457 , \47158_47458 , \47159_47459 , \47160_47460 , \47161_47461 , \47162_47462 , \47163_47463 , \47164_47464 , \47165_47465 , \47166_47466 ,
         \47167_47467 , \47168_47468 , \47169_47469 , \47170_47470 , \47171_47471 , \47172_47472 , \47173_47473 , \47174_47474 , \47175_47475 , \47176_47476 ,
         \47177_47477 , \47178_47478 , \47179_47479 , \47180_47480 , \47181_47481 , \47182_47482 , \47183_47483 , \47184_47484 , \47185_47485 , \47186_47486 ,
         \47187_47487 , \47188_47488 , \47189_47489 , \47190_47490 , \47191_47491 , \47192_47492 , \47193_47493 , \47194_47494 , \47195_47495 , \47196_47496 ,
         \47197_47497 , \47198_47498 , \47199_47499 , \47200_47500 , \47201_47501 , \47202_47502 , \47203_47503 , \47204_47504 , \47205_47505 , \47206_47506 ,
         \47207_47507 , \47208_47508 , \47209_47509 , \47210_47510 , \47211_47511 , \47212_47512 , \47213_47513 , \47214_47514 , \47215_47515 , \47216_47516 ,
         \47217_47517 , \47218_47518 , \47219_47519 , \47220_47520 , \47221_47521 , \47222_47522 , \47223_47523 , \47224_47524 , \47225_47525 , \47226_47526 ,
         \47227_47527 , \47228_47528 , \47229_47529 , \47230_47530 , \47231_47531 , \47232_47532 , \47233_47533 , \47234_47534 , \47235_47535 , \47236_47536 ,
         \47237_47537 , \47238_47538 , \47239_47539 , \47240_47540 , \47241_47541 , \47242_47542 , \47243_47543 , \47244_47544 , \47245_47545 , \47246_47546 ,
         \47247_47547 , \47248_47548 , \47249_47549 , \47250_47550 , \47251_47551 , \47252_47552 , \47253_47553 , \47254_47554 , \47255_47555 , \47256_47556 ,
         \47257_47557 , \47258_47558 , \47259_47559 , \47260_47560 , \47261_47561 , \47262_47562 , \47263_47563 , \47264_47564 , \47265_47565 , \47266_47566 ,
         \47267_47567 , \47268_47568 , \47269_47569 , \47270_47570 , \47271_47571 , \47272_47572 , \47273_47573 , \47274_47574 , \47275_47575 , \47276_47576 ,
         \47277_47577 , \47278_47578 , \47279_47579 , \47280_47580 , \47281_47581 , \47282_47582 , \47283_47583 , \47284_47584 , \47285_47585 , \47286_47586 ,
         \47287_47587 , \47288_47588 , \47289_47589 , \47290_47590 , \47291_47591 , \47292_47592 , \47293_47593 , \47294_47594 , \47295_47595 , \47296_47596 ,
         \47297_47597 , \47298_47598 , \47299_47599 , \47300_47600 , \47301_47601 , \47302_47602 , \47303_47603 , \47304_47604 , \47305_47605 , \47306_47606 ,
         \47307_47607 , \47308_47608_nGdf4e , \47309_R_58_102f1b78 , \47310_47610 , \47311_47611 , \47312_47612_nGdf51 , \47313_R_59_be1fc68 , \47314_47614 , \47315_47615_nGdf53 , \47316_R_5a_10279198 ,
         \47317_47617 , \47318_47618_nGdf55 , \47319_R_5b_102299e8 , \47320_47620 , \47321_47621_nGdf57 , \47322_R_5c_101d0448 , \47323_47623 , \47324_47624_nGdf59 , \47325_R_5d_f7f82f0 , \47326_47626 ,
         \47327_47627_nGdf5b , \47328_R_5e_be21600 , \47329_47629 , \47330_47630_nGdf5d , \47331_R_5f_f7fa5b8 , \47332_47632 , \47333_47633_nGdf5f , \47334_R_60_1027d530 , \47335_47635 , \47336_47636_nGdf61 ,
         \47337_R_61_10205ae8 , \47338_47638 , \47339_47639_nGdf63 , \47340_R_62_10283510 , \47341_47641 , \47342_47642_nGdf65 , \47343_R_63_f82b578 , \47344_47644 , \47345_47645_nGdf67 , \47346_R_64_ace4e68 ,
         \47347_47647 , \47348_47648_nGdf69 , \47349_R_65_f8204e0 , \47350_47650 , \47351_47651_nGdf6b , \47352_R_66_1027a0b0 , \47353_47653 , \47354_47654_nGdf6d , \47355_R_67_1022dc30 , \47356_47656 ,
         \47357_47657_nGdf6f , \47358_R_68_102478a8 , \47359_47659 , \47360_47660_nGdf71 , \47361_R_69_10286f78 , \47362_47662 , \47363_47663_nGdf73 , \47364_R_6a_f7edd80 , \47365_47665 , \47366_47666_nGdf75 ,
         \47367_R_6b_101c3628 , \47368_47668 , \47369_47669_nGdf77 , \47370_R_6c_f7fbe00 , \47371_47671 , \47372_47672_nGdf79 , \47373_R_6d_f7ce9f8 , \47374_47674 , \47375_47675_nGdf7b , \47376_R_6e_f7c8830 ,
         \47377_47677 , \47378_47678_nGdf7d , \47379_R_6f_101ffc68 , \47380_47680 , \47381_47681_nGdf7f , \47382_R_70_f7d4000 , \47383_47683 , \47384_47684_nGdf81 , \47385_R_71_acee958 , \47386_47686 ,
         \47387_47687_nGdf83 , \47388_R_72_94046c0 , \47389_47689 , \47390_47690_nGdf85 , \47391_R_73_101ee420 , \47392_47692 , \47393_47693_nGdf87 , \47394_R_74_102eb268 , \47395_47695 , \47396_47696_nGdf89 ,
         \47397_R_75_b320c50 , \47398_47698 , \47399_47699_nGdf8b , \47400_R_76_ad80a90 , \47401_47701 , \47402_47702_nGdf8d , \47403_R_77_1027fd48 , \47404_47704 , \47405_47705_nGdf8f , \47406_R_78_f7ce4b8 ,
         \47407_47707 , \47408_47708_nGdf91 , \47409_R_79_ad77048 , \47410_47710 , \47411_47711_nGdf93 , \47412_R_7a_102a6ae0 , \47413_47713 , \47414_47714_nGdf95 , \47415_R_7b_f7e4c78 , \47416_47716 ,
         \47417_47717_nGdf97 , \47418_R_7c_e2a6ce0 , \47419_47719 , \47420_47720_nGdf99 , \47421_R_7d_101e86e0 , \47422_47722 , \47423_47723_nGdf9b , \47424_R_7e_e2a9cc8 , \47425_47725 , \47426_47726_nGdf9d ,
         \47427_R_7f_10292be0 , \47428_47728 , \47429_47729_nGdf9f , \47430_R_80_b33cde8 , \47431_47731 , \47432_47732_nGdfa1 , \47433_R_81_101e2908 , \47434_47734 , \47435_47735_nGdfa3 , \47436_R_82_102e9780 ,
         \47437_47737 , \47438_47738_nGdfa5 , \47439_R_83_f8157a0 , \47440_47740 , \47441_47741_nGdfa7 , \47442_R_84_f819358 , \47443_47743 , \47444_47744_nGdfa9 , \47445_R_85_ace8b70 , \47446_47746 ,
         \47447_47747_nGdfab , \47448_R_86_be142b0 , \47449_47749 , \47450_47750_nGdfad , \47451_R_87_f81b770 , \47452_47752 , \47453_47753_nGdfaf , \47454_R_88_b330278 , \47455_47755 , \47456_47756_nGdfb1 ,
         \47457_R_89_f7fe9f8 , \47458_47758 , \47459_47759_nGdfb3 , \47460_R_8a_101cf488 , \47461_47761 , \47462_47762_nGdfb5 , \47463_R_8b_f8225c0 , \47464_47764 , \47465_47765_nGdfb7 , \47466_R_8c_101d4738 ,
         \47467_47767 , \47468_47768_nGdfb9 , \47469_R_8d_101c4000 , \47470_47770 , \47471_47771_nGdfbb , \47472_R_8e_101fe960 , \47473_47773 , \47474_47774_nGdfbd , \47475_R_8f_102a0330 , \47476_47776 ,
         \47477_47777_nGdfbf , \47478_R_90_f7f4bd0 , \47479_47779 , \47480_47780_nGdfc1 , \47481_R_91_1023e5a8 , \47482_47782 , \47483_47783_nGdfc3 , \47484_R_92_10248da8 , \47485_47785 , \47486_47786_nGdfc5 ,
         \47487_R_93_be2c938 , \47488_47788 , \47489_47789_nGdfc7 , \47490_R_94_f7f5458 , \47491_47791 , \47492_47792 , \47493_47793_nGdfca , \47494_R_95_f7c6808 , \47495_47795 , \47496_47796 ,
         \47497_47797_nGdfcd , \47498_R_96_be316a8 , \47499_47799 , \47500_47800 , \47501_47801_nGdfd0 , \47502_R_97_e2a0328 , \47503_47803 , \47504_47804_nGdfd2 , \47505_R_98_be2d850 , \47506_47806 ,
         \47507_47807 , \47508_47808_nGdfd5 , \47509_R_99_10217db0 , \47510_47810 , \47511_47811_nGdfd7 , \47512_R_9a_f7ec340 , \47513_47813 , \47514_47814 , \47515_47815_nGdfda , \47516_R_9b_be23ec0 ,
         \47517_47817 , \47518_47818_nGdfdc , \47519_R_9c_101d4540 , \47520_47820 , \47521_47821 , \47522_47822_nGdfdf , \47523_R_9d_f800828 , \47524_47824 , \47525_47825_nGdfe1 , \47526_R_9e_102970c8 ,
         \47527_47827 , \47528_47828 , \47529_47829_nGdfe4 , \47530_R_9f_10221de0 , \47531_47831 , \47532_47832_nGdfe6 , \47533_R_a0_ad8d568 , \47534_47834 , \47535_47835 , \47536_47836_nGdfe9 ,
         \47537_R_a1_be4eb58 , \47538_47838 , \47539_47839_nGdfeb , \47540_R_a2_f7c5500 , \47541_47841 , \47542_47842 , \47543_47843_nGdfee , \47544_R_a3_ad88f30 , \47545_47845 , \47546_47846_nGdff0 ,
         \47547_R_a4_f82f088 , \47548_47848 , \47549_47849 , \47550_47850_nGdff3 , \47551_R_a5_f7dcbc8 , \47552_47852 , \47553_47853_nGdff5 , \47554_R_a6_10292940 , \47555_47855 , \47556_47856 ,
         \47557_47857_nGdff8 , \47558_R_a7_be138d8 , \47559_47859 , \47560_47860_nGdffa , \47561_R_a8_acee418 , \47562_47862 , \47563_47863 , \47564_47864_nGdffd , \47565_R_a9_ad84450 , \47566_47866 ,
         \47567_47867_nGdfff , \47568_R_aa_be10838 , \47569_47869 , \47570_47870 , \47571_47871_nGe002 , \47572_R_ab_be31fd8 , \47573_47873 , \47574_47874_nGe004 , \47575_R_ac_acdaef0 , \47576_47876 ,
         \47577_47877 , \47578_47878_nGe007 , \47579_R_ad_acea908 , \47580_47880 , \47581_47881_nGe009 , \47582_R_ae_101f8830 , \47583_47883 , \47584_47884 , \47585_47885_nGe00c , \47586_R_af_f7dec98 ,
         \47587_47887 , \47588_47888_nGe00e , \47589_R_b0_101e2c50 , \47590_47890 , \47591_47891 , \47592_47892_nGe011 , \47593_R_b1_f801b30 , \47594_47894 , \47595_47895_nGe013 , \47596_R_b2_be16e00 ,
         \47597_47897 , \47598_47898 , \47599_47899_nGe016 , \47600_R_b3_102e3cf0 , \47601_47901 , \47602_47902_nGe018 , \47603_R_b4_10291788 ;
buf \U$labajz5598 ( R_58_102f1b78, \47309_R_58_102f1b78 );
buf \U$labajz5599 ( R_59_be1fc68, \47313_R_59_be1fc68 );
buf \U$labajz5600 ( R_5a_10279198, \47316_R_5a_10279198 );
buf \U$labajz5601 ( R_5b_102299e8, \47319_R_5b_102299e8 );
buf \U$labajz5602 ( R_5c_101d0448, \47322_R_5c_101d0448 );
buf \U$labajz5603 ( R_5d_f7f82f0, \47325_R_5d_f7f82f0 );
buf \U$labajz5604 ( R_5e_be21600, \47328_R_5e_be21600 );
buf \U$labajz5605 ( R_5f_f7fa5b8, \47331_R_5f_f7fa5b8 );
buf \U$labajz5606 ( R_60_1027d530, \47334_R_60_1027d530 );
buf \U$labajz5607 ( R_61_10205ae8, \47337_R_61_10205ae8 );
buf \U$labajz5608 ( R_62_10283510, \47340_R_62_10283510 );
buf \U$labajz5609 ( R_63_f82b578, \47343_R_63_f82b578 );
buf \U$labajz5610 ( R_64_ace4e68, \47346_R_64_ace4e68 );
buf \U$labajz5611 ( R_65_f8204e0, \47349_R_65_f8204e0 );
buf \U$labajz5612 ( R_66_1027a0b0, \47352_R_66_1027a0b0 );
buf \U$labajz5613 ( R_67_1022dc30, \47355_R_67_1022dc30 );
buf \U$labajz5614 ( R_68_102478a8, \47358_R_68_102478a8 );
buf \U$labajz5615 ( R_69_10286f78, \47361_R_69_10286f78 );
buf \U$labajz5616 ( R_6a_f7edd80, \47364_R_6a_f7edd80 );
buf \U$labajz5617 ( R_6b_101c3628, \47367_R_6b_101c3628 );
buf \U$labajz5618 ( R_6c_f7fbe00, \47370_R_6c_f7fbe00 );
buf \U$labajz5619 ( R_6d_f7ce9f8, \47373_R_6d_f7ce9f8 );
buf \U$labajz5620 ( R_6e_f7c8830, \47376_R_6e_f7c8830 );
buf \U$labajz5621 ( R_6f_101ffc68, \47379_R_6f_101ffc68 );
buf \U$labajz5622 ( R_70_f7d4000, \47382_R_70_f7d4000 );
buf \U$labajz5623 ( R_71_acee958, \47385_R_71_acee958 );
buf \U$labajz5624 ( R_72_94046c0, \47388_R_72_94046c0 );
buf \U$labajz5625 ( R_73_101ee420, \47391_R_73_101ee420 );
buf \U$labajz5626 ( R_74_102eb268, \47394_R_74_102eb268 );
buf \U$labajz5627 ( R_75_b320c50, \47397_R_75_b320c50 );
buf \U$labajz5628 ( R_76_ad80a90, \47400_R_76_ad80a90 );
buf \U$labajz5629 ( R_77_1027fd48, \47403_R_77_1027fd48 );
buf \U$labajz5630 ( R_78_f7ce4b8, \47406_R_78_f7ce4b8 );
buf \U$labajz5631 ( R_79_ad77048, \47409_R_79_ad77048 );
buf \U$labajz5632 ( R_7a_102a6ae0, \47412_R_7a_102a6ae0 );
buf \U$labajz5633 ( R_7b_f7e4c78, \47415_R_7b_f7e4c78 );
buf \U$labajz5634 ( R_7c_e2a6ce0, \47418_R_7c_e2a6ce0 );
buf \U$labajz5635 ( R_7d_101e86e0, \47421_R_7d_101e86e0 );
buf \U$labajz5636 ( R_7e_e2a9cc8, \47424_R_7e_e2a9cc8 );
buf \U$labajz5637 ( R_7f_10292be0, \47427_R_7f_10292be0 );
buf \U$labajz5638 ( R_80_b33cde8, \47430_R_80_b33cde8 );
buf \U$labajz5639 ( R_81_101e2908, \47433_R_81_101e2908 );
buf \U$labajz5640 ( R_82_102e9780, \47436_R_82_102e9780 );
buf \U$labajz5641 ( R_83_f8157a0, \47439_R_83_f8157a0 );
buf \U$labajz5642 ( R_84_f819358, \47442_R_84_f819358 );
buf \U$labajz5643 ( R_85_ace8b70, \47445_R_85_ace8b70 );
buf \U$labajz5644 ( R_86_be142b0, \47448_R_86_be142b0 );
buf \U$labajz5645 ( R_87_f81b770, \47451_R_87_f81b770 );
buf \U$labajz5646 ( R_88_b330278, \47454_R_88_b330278 );
buf \U$labajz5647 ( R_89_f7fe9f8, \47457_R_89_f7fe9f8 );
buf \U$labajz5648 ( R_8a_101cf488, \47460_R_8a_101cf488 );
buf \U$labajz5649 ( R_8b_f8225c0, \47463_R_8b_f8225c0 );
buf \U$labajz5650 ( R_8c_101d4738, \47466_R_8c_101d4738 );
buf \U$labajz5651 ( R_8d_101c4000, \47469_R_8d_101c4000 );
buf \U$labajz5652 ( R_8e_101fe960, \47472_R_8e_101fe960 );
buf \U$labajz5653 ( R_8f_102a0330, \47475_R_8f_102a0330 );
buf \U$labajz5654 ( R_90_f7f4bd0, \47478_R_90_f7f4bd0 );
buf \U$labajz5655 ( R_91_1023e5a8, \47481_R_91_1023e5a8 );
buf \U$labajz5656 ( R_92_10248da8, \47484_R_92_10248da8 );
buf \U$labajz5657 ( R_93_be2c938, \47487_R_93_be2c938 );
buf \U$labajz5658 ( R_94_f7f5458, \47490_R_94_f7f5458 );
buf \U$labajz5659 ( R_95_f7c6808, \47494_R_95_f7c6808 );
buf \U$labajz5660 ( R_96_be316a8, \47498_R_96_be316a8 );
buf \U$labajz5661 ( R_97_e2a0328, \47502_R_97_e2a0328 );
buf \U$labajz5662 ( R_98_be2d850, \47505_R_98_be2d850 );
buf \U$labajz5663 ( R_99_10217db0, \47509_R_99_10217db0 );
buf \U$labajz5664 ( R_9a_f7ec340, \47512_R_9a_f7ec340 );
buf \U$labajz5665 ( R_9b_be23ec0, \47516_R_9b_be23ec0 );
buf \U$labajz5666 ( R_9c_101d4540, \47519_R_9c_101d4540 );
buf \U$labajz5667 ( R_9d_f800828, \47523_R_9d_f800828 );
buf \U$labajz5668 ( R_9e_102970c8, \47526_R_9e_102970c8 );
buf \U$labajz5669 ( R_9f_10221de0, \47530_R_9f_10221de0 );
buf \U$labajz5670 ( R_a0_ad8d568, \47533_R_a0_ad8d568 );
buf \U$labajz5671 ( R_a1_be4eb58, \47537_R_a1_be4eb58 );
buf \U$labajz5672 ( R_a2_f7c5500, \47540_R_a2_f7c5500 );
buf \U$labajz5673 ( R_a3_ad88f30, \47544_R_a3_ad88f30 );
buf \U$labajz5674 ( R_a4_f82f088, \47547_R_a4_f82f088 );
buf \U$labajz5675 ( R_a5_f7dcbc8, \47551_R_a5_f7dcbc8 );
buf \U$labajz5676 ( R_a6_10292940, \47554_R_a6_10292940 );
buf \U$labajz5677 ( R_a7_be138d8, \47558_R_a7_be138d8 );
buf \U$labajz5678 ( R_a8_acee418, \47561_R_a8_acee418 );
buf \U$labajz5679 ( R_a9_ad84450, \47565_R_a9_ad84450 );
buf \U$labajz5680 ( R_aa_be10838, \47568_R_aa_be10838 );
buf \U$labajz5681 ( R_ab_be31fd8, \47572_R_ab_be31fd8 );
buf \U$labajz5682 ( R_ac_acdaef0, \47575_R_ac_acdaef0 );
buf \U$labajz5683 ( R_ad_acea908, \47579_R_ad_acea908 );
buf \U$labajz5684 ( R_ae_101f8830, \47582_R_ae_101f8830 );
buf \U$labajz5685 ( R_af_f7dec98, \47586_R_af_f7dec98 );
buf \U$labajz5686 ( R_b0_101e2c50, \47589_R_b0_101e2c50 );
buf \U$labajz5687 ( R_b1_f801b30, \47593_R_b1_f801b30 );
buf \U$labajz5688 ( R_b2_be16e00, \47596_R_b2_be16e00 );
buf \U$labajz5689 ( R_b3_102e3cf0, \47600_R_b3_102e3cf0 );
buf \U$labajz5690 ( R_b4_10291788, \47603_R_b4_10291788 );
not \U$1 ( \8753_9052 , RIbc62af0_23);
not \U$2 ( \8754_9053 , RIbc62a78_22);
not \U$3 ( \8755_9054 , RIbc62a00_21);
not \U$4 ( \8756_9055 , RIbc62988_20);
not \U$5 ( \8757_9056 , RIbc62910_19);
not \U$6 ( \8758_9057 , RIbc62898_18);
not \U$7 ( \8759_9058 , RIbc62820_17);
nor \U$8 ( \8760_9059 , \8753_9052 , \8754_9053 , \8755_9054 , \8756_9055 , \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$9 ( \8761_9060 , RIdec64b8_720, \8760_9059 );
nor \U$10 ( \8762_9061 , RIbc62af0_23, \8754_9053 , \8755_9054 , \8756_9055 , \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$11 ( \8763_9062 , RIdec37b8_688, \8762_9061 );
nor \U$12 ( \8764_9063 , \8753_9052 , RIbc62a78_22, \8755_9054 , \8756_9055 , \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$13 ( \8765_9064 , RIfc8daa0_6634, \8764_9063 );
nor \U$14 ( \8766_9065 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , \8756_9055 , \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$15 ( \8767_9066 , RIdec0ab8_656, \8766_9065 );
nor \U$16 ( \8768_9067 , \8753_9052 , \8754_9053 , RIbc62a00_21, \8756_9055 , \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$17 ( \8769_9068 , RIfc56348_6003, \8768_9067 );
nor \U$18 ( \8770_9069 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, \8756_9055 , \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$19 ( \8771_9070 , RIdebddb8_624, \8770_9069 );
nor \U$20 ( \8772_9071 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, \8756_9055 , \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$21 ( \8773_9072 , RIdebb0b8_592, \8772_9071 );
nor \U$22 ( \8774_9073 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \8756_9055 , \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$23 ( \8775_9074 , RIdeb83b8_560, \8774_9073 );
nor \U$24 ( \8776_9075 , \8753_9052 , \8754_9053 , \8755_9054 , RIbc62988_20, \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$25 ( \8777_9076 , RIfc98798_6757, \8776_9075 );
nor \U$26 ( \8778_9077 , RIbc62af0_23, \8754_9053 , \8755_9054 , RIbc62988_20, \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$27 ( \8779_9078 , RIdeb29b8_496, \8778_9077 );
nor \U$28 ( \8780_9079 , \8753_9052 , RIbc62a78_22, \8755_9054 , RIbc62988_20, \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$29 ( \8781_9080 , RIfcbd098_7173, \8780_9079 );
nor \U$30 ( \8782_9081 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , RIbc62988_20, \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$31 ( \8783_9082 , RIdeafcb8_464, \8782_9081 );
nor \U$32 ( \8784_9083 , \8753_9052 , \8754_9053 , RIbc62a00_21, RIbc62988_20, \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$33 ( \8785_9084 , RIfc8dc08_6635, \8784_9083 );
nor \U$34 ( \8786_9085 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, RIbc62988_20, \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$35 ( \8787_9086 , RIdeacb80_432, \8786_9085 );
nor \U$36 ( \8788_9087 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$37 ( \8789_9088 , RIdea6280_400, \8788_9087 );
nor \U$38 ( \8790_9089 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \8757_9056 , \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$39 ( \8791_9090 , RIde9f980_368, \8790_9089 );
nor \U$40 ( \8792_9091 , \8753_9052 , \8754_9053 , \8755_9054 , \8756_9055 , RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$41 ( \8793_9092 , RIfcd6868_7463, \8792_9091 );
nor \U$42 ( \8794_9093 , RIbc62af0_23, \8754_9053 , \8755_9054 , \8756_9055 , RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$43 ( \8795_9094 , RIfc8ded8_6637, \8794_9093 );
nor \U$44 ( \8796_9095 , \8753_9052 , RIbc62a78_22, \8755_9054 , \8756_9055 , RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$45 ( \8797_9096 , RIfc7dd80_6454, \8796_9095 );
nor \U$46 ( \8798_9097 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , \8756_9055 , RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$47 ( \8799_9098 , RIfc56618_6005, \8798_9097 );
nor \U$48 ( \8800_9099 , \8753_9052 , \8754_9053 , RIbc62a00_21, \8756_9055 , RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$49 ( \8801_9100 , RIde92e10_306, \8800_9099 );
nor \U$50 ( \8802_9101 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, \8756_9055 , RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$51 ( \8803_9102 , RIde8f300_288, \8802_9101 );
nor \U$52 ( \8804_9103 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, \8756_9055 , RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$53 ( \8805_9104 , RIde8b160_268, \8804_9103 );
nor \U$54 ( \8806_9105 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \8756_9055 , RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$55 ( \8807_9106 , RIde86fc0_248, \8806_9105 );
nor \U$56 ( \8808_9107 , \8753_9052 , \8754_9053 , \8755_9054 , RIbc62988_20, RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$57 ( \8809_9108 , RIde82ad8_227, \8808_9107 );
nor \U$58 ( \8810_9109 , RIbc62af0_23, \8754_9053 , \8755_9054 , RIbc62988_20, RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$59 ( \8811_9110 , RIfc8e040_6638, \8810_9109 );
nor \U$60 ( \8812_9111 , \8753_9052 , RIbc62a78_22, \8755_9054 , RIbc62988_20, RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$61 ( \8813_9112 , RIfcd96d0_7496, \8812_9111 );
nor \U$62 ( \8814_9113 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , RIbc62988_20, RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$63 ( \8815_9114 , RIfca1e10_6864, \8814_9113 );
nor \U$64 ( \8816_9115 , \8753_9052 , \8754_9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$65 ( \8817_9116 , RIfcbd200_7174, \8816_9115 );
nor \U$66 ( \8818_9117 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$67 ( \8819_9118 , RIe16c5c0_2610, \8818_9117 );
nor \U$68 ( \8820_9119 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$69 ( \8821_9120 , RIe16a298_2585, \8820_9119 );
nor \U$70 ( \8822_9121 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, \8758_9057 , \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$71 ( \8823_9122 , RIe168ab0_2568, \8822_9121 );
nor \U$72 ( \8824_9123 , \8753_9052 , \8754_9053 , \8755_9054 , \8756_9055 , \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$73 ( \8825_9124 , RIe1664b8_2541, \8824_9123 );
nor \U$74 ( \8826_9125 , RIbc62af0_23, \8754_9053 , \8755_9054 , \8756_9055 , \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$75 ( \8827_9126 , RIe1637b8_2509, \8826_9125 );
nor \U$76 ( \8828_9127 , \8753_9052 , RIbc62a78_22, \8755_9054 , \8756_9055 , \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$77 ( \8829_9128 , RIee37f00_5095, \8828_9127 );
nor \U$78 ( \8830_9129 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , \8756_9055 , \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$79 ( \8831_9130 , RIe160ab8_2477, \8830_9129 );
nor \U$80 ( \8832_9131 , \8753_9052 , \8754_9053 , RIbc62a00_21, \8756_9055 , \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$81 ( \8833_9132 , RIfc8ea18_6645, \8832_9131 );
nor \U$82 ( \8834_9133 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, \8756_9055 , \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$83 ( \8835_9134 , RIe15ddb8_2445, \8834_9133 );
nor \U$84 ( \8836_9135 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, \8756_9055 , \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$85 ( \8837_9136 , RIe1583b8_2381, \8836_9135 );
nor \U$86 ( \8838_9137 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \8756_9055 , \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$87 ( \8839_9138 , RIe1556b8_2349, \8838_9137 );
nor \U$88 ( \8840_9139 , \8753_9052 , \8754_9053 , \8755_9054 , RIbc62988_20, \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$89 ( \8841_9140 , RIfe9f828_8159, \8840_9139 );
nor \U$90 ( \8842_9141 , RIbc62af0_23, \8754_9053 , \8755_9054 , RIbc62988_20, \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$91 ( \8843_9142 , RIe1529b8_2317, \8842_9141 );
nor \U$92 ( \8844_9143 , \8753_9052 , RIbc62a78_22, \8755_9054 , RIbc62988_20, \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$93 ( \8845_9144 , RIfe9f990_8160, \8844_9143 );
nor \U$94 ( \8846_9145 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , RIbc62988_20, \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$95 ( \8847_9146 , RIe14fcb8_2285, \8846_9145 );
nor \U$96 ( \8848_9147 , \8753_9052 , \8754_9053 , RIbc62a00_21, RIbc62988_20, \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$97 ( \8849_9148 , RIfcbd368_7175, \8848_9147 );
nor \U$98 ( \8850_9149 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, RIbc62988_20, \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$99 ( \8851_9150 , RIe14cfb8_2253, \8850_9149 );
nor \U$100 ( \8852_9151 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$101 ( \8853_9152 , RIe14a2b8_2221, \8852_9151 );
nor \U$102 ( \8854_9153 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \8757_9056 , RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$103 ( \8855_9154 , RIe1475b8_2189, \8854_9153 );
nor \U$104 ( \8856_9155 , \8753_9052 , \8754_9053 , \8755_9054 , \8756_9055 , RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$105 ( \8857_9156 , RIfc8ee50_6648, \8856_9155 );
nor \U$106 ( \8858_9157 , RIbc62af0_23, \8754_9053 , \8755_9054 , \8756_9055 , RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$107 ( \8859_9158 , RIfc45278_5809, \8858_9157 );
nor \U$108 ( \8860_9159 , \8753_9052 , RIbc62a78_22, \8755_9054 , \8756_9055 , RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$109 ( \8861_9160 , RIfc98360_6754, \8860_9159 );
nor \U$110 ( \8862_9161 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , \8756_9055 , RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$111 ( \8863_9162 , RIfca2248_6867, \8862_9161 );
nor \U$112 ( \8864_9163 , \8753_9052 , \8754_9053 , RIbc62a00_21, \8756_9055 , RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$113 ( \8865_9164 , RIe141d20_2126, \8864_9163 );
nor \U$114 ( \8866_9165 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, \8756_9055 , RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$115 ( \8867_9166 , RIe13f9f8_2101, \8866_9165 );
nor \U$116 ( \8868_9167 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, \8756_9055 , RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$117 ( \8869_9168 , RIdf3d900_2077, \8868_9167 );
nor \U$118 ( \8870_9169 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \8756_9055 , RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$119 ( \8871_9170 , RIdf3b470_2051, \8870_9169 );
nor \U$120 ( \8872_9171 , \8753_9052 , \8754_9053 , \8755_9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$121 ( \8873_9172 , RIfcd6ca0_7466, \8872_9171 );
nor \U$122 ( \8874_9173 , RIbc62af0_23, \8754_9053 , \8755_9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$123 ( \8875_9174 , RIee2ff08_5004, \8874_9173 );
nor \U$124 ( \8876_9175 , \8753_9052 , RIbc62a78_22, \8755_9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$125 ( \8877_9176 , RIfc8ece8_6647, \8876_9175 );
nor \U$126 ( \8878_9177 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$127 ( \8879_9178 , RIee2dd48_4980, \8878_9177 );
nor \U$128 ( \8880_9179 , \8753_9052 , \8754_9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$129 ( \8881_9180 , RIdf36718_1996, \8880_9179 );
nor \U$130 ( \8882_9181 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$131 ( \8883_9182 , RIdf34120_1969, \8882_9181 );
nor \U$132 ( \8884_9183 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$133 ( \8885_9184 , RIdf31f60_1945, \8884_9183 );
nor \U$134 ( \8886_9185 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, \8759_9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$135 ( \8887_9186 , RIfe9f6c0_8158, \8886_9185 );
or \U$136 ( \8888_9187 , \8761_9060 , \8763_9062 , \8765_9064 , \8767_9066 , \8769_9068 , \8771_9070 , \8773_9072 , \8775_9074 , \8777_9076 , \8779_9078 , \8781_9080 , \8783_9082 , \8785_9084 , \8787_9086 , \8789_9088 , \8791_9090 , \8793_9092 , \8795_9094 , \8797_9096 , \8799_9098 , \8801_9100 , \8803_9102 , \8805_9104 , \8807_9106 , \8809_9108 , \8811_9110 , \8813_9112 , \8815_9114 , \8817_9116 , \8819_9118 , \8821_9120 , \8823_9122 , \8825_9124 , \8827_9126 , \8829_9128 , \8831_9130 , \8833_9132 , \8835_9134 , \8837_9136 , \8839_9138 , \8841_9140 , \8843_9142 , \8845_9144 , \8847_9146 , \8849_9148 , \8851_9150 , \8853_9152 , \8855_9154 , \8857_9156 , \8859_9158 , \8861_9160 , \8863_9162 , \8865_9164 , \8867_9166 , \8869_9168 , \8871_9170 , \8873_9172 , \8875_9174 , \8877_9176 , \8879_9178 , \8881_9180 , \8883_9182 , \8885_9184 , \8887_9186 );
nor \U$137 ( \8889_9188 , \8753_9052 , \8754_9053 , \8755_9054 , \8756_9055 , \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$138 ( \8890_9189 , RIfcb4560_7074, \8889_9188 );
nor \U$139 ( \8891_9190 , RIbc62af0_23, \8754_9053 , \8755_9054 , \8756_9055 , \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$140 ( \8892_9191 , RIfc45db8_5817, \8891_9190 );
nor \U$141 ( \8893_9192 , \8753_9052 , RIbc62a78_22, \8755_9054 , \8756_9055 , \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$142 ( \8894_9193 , RIfc8e1a8_6639, \8893_9192 );
nor \U$143 ( \8895_9194 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , \8756_9055 , \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$144 ( \8896_9195 , RIfc7d678_6449, \8895_9194 );
nor \U$145 ( \8897_9196 , \8753_9052 , \8754_9053 , RIbc62a00_21, \8756_9055 , \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$146 ( \8898_9197 , RIdf2aee0_1865, \8897_9196 );
nor \U$147 ( \8899_9198 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, \8756_9055 , \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$148 ( \8900_9199 , RIdf28ff0_1843, \8899_9198 );
nor \U$149 ( \8901_9200 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, \8756_9055 , \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$150 ( \8902_9201 , RIdf26e30_1819, \8901_9200 );
nor \U$151 ( \8903_9202 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \8756_9055 , \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$152 ( \8904_9203 , RIdf25378_1800, \8903_9202 );
nor \U$153 ( \8905_9204 , \8753_9052 , \8754_9053 , \8755_9054 , RIbc62988_20, \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$154 ( \8906_9205 , RIfcb43f8_7073, \8905_9204 );
nor \U$155 ( \8907_9206 , RIbc62af0_23, \8754_9053 , \8755_9054 , RIbc62988_20, \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$156 ( \8908_9207 , RIfc8e748_6643, \8907_9206 );
nor \U$157 ( \8909_9208 , \8753_9052 , RIbc62a78_22, \8755_9054 , RIbc62988_20, \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$158 ( \8910_9209 , RIdf23488_1778, \8909_9208 );
nor \U$159 ( \8911_9210 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , RIbc62988_20, \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$160 ( \8912_9211 , RIfcc2c00_7238, \8911_9210 );
nor \U$161 ( \8913_9212 , \8753_9052 , \8754_9053 , RIbc62a00_21, RIbc62988_20, \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$162 ( \8914_9213 , RIdf21e08_1762, \8913_9212 );
nor \U$163 ( \8915_9214 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, RIbc62988_20, \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$164 ( \8916_9215 , RIdf20788_1746, \8915_9214 );
nor \U$165 ( \8917_9216 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$166 ( \8918_9217 , RIdf1b760_1689, \8917_9216 );
nor \U$167 ( \8919_9218 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \8757_9056 , \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$168 ( \8920_9219 , RIdf1a248_1674, \8919_9218 );
nor \U$169 ( \8921_9220 , \8753_9052 , \8754_9053 , \8755_9054 , \8756_9055 , RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$170 ( \8922_9221 , RIdf18088_1650, \8921_9220 );
nor \U$171 ( \8923_9222 , RIbc62af0_23, \8754_9053 , \8755_9054 , \8756_9055 , RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$172 ( \8924_9223 , RIdf15388_1618, \8923_9222 );
nor \U$173 ( \8925_9224 , \8753_9052 , RIbc62a78_22, \8755_9054 , \8756_9055 , RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$174 ( \8926_9225 , RIdf12688_1586, \8925_9224 );
nor \U$175 ( \8927_9226 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , \8756_9055 , RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$176 ( \8928_9227 , RIdf0f988_1554, \8927_9226 );
nor \U$177 ( \8929_9228 , \8753_9052 , \8754_9053 , RIbc62a00_21, \8756_9055 , RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$178 ( \8930_9229 , RIdf0cc88_1522, \8929_9228 );
nor \U$179 ( \8931_9230 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, \8756_9055 , RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$180 ( \8932_9231 , RIdf09f88_1490, \8931_9230 );
nor \U$181 ( \8933_9232 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, \8756_9055 , RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$182 ( \8934_9233 , RIdf07288_1458, \8933_9232 );
nor \U$183 ( \8935_9234 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \8756_9055 , RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$184 ( \8936_9235 , RIdf04588_1426, \8935_9234 );
nor \U$185 ( \8937_9236 , \8753_9052 , \8754_9053 , \8755_9054 , RIbc62988_20, RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$186 ( \8938_9237 , RIdefeb88_1362, \8937_9236 );
nor \U$187 ( \8939_9238 , RIbc62af0_23, \8754_9053 , \8755_9054 , RIbc62988_20, RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$188 ( \8940_9239 , RIdefbe88_1330, \8939_9238 );
nor \U$189 ( \8941_9240 , \8753_9052 , RIbc62a78_22, \8755_9054 , RIbc62988_20, RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$190 ( \8942_9241 , RIdef9188_1298, \8941_9240 );
nor \U$191 ( \8943_9242 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , RIbc62988_20, RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$192 ( \8944_9243 , RIdef6488_1266, \8943_9242 );
nor \U$193 ( \8945_9244 , \8753_9052 , \8754_9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$194 ( \8946_9245 , RIdef3788_1234, \8945_9244 );
nor \U$195 ( \8947_9246 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$196 ( \8948_9247 , RIdef0a88_1202, \8947_9246 );
nor \U$197 ( \8949_9248 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$198 ( \8950_9249 , RIdeedd88_1170, \8949_9248 );
nor \U$199 ( \8951_9250 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, \8758_9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$200 ( \8952_9251 , RIdeeb088_1138, \8951_9250 );
nor \U$201 ( \8953_9252 , \8753_9052 , \8754_9053 , \8755_9054 , \8756_9055 , \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$202 ( \8954_9253 , RIfc8efb8_6649, \8953_9252 );
nor \U$203 ( \8955_9254 , RIbc62af0_23, \8754_9053 , \8755_9054 , \8756_9055 , \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$204 ( \8956_9255 , RIfc44e40_5806, \8955_9254 );
nor \U$205 ( \8957_9256 , \8753_9052 , RIbc62a78_22, \8755_9054 , \8756_9055 , \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$206 ( \8958_9257 , RIfc57860_6018, \8957_9256 );
nor \U$207 ( \8959_9258 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , \8756_9055 , \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$208 ( \8960_9259 , RIfca23b0_6868, \8959_9258 );
nor \U$209 ( \8961_9260 , \8753_9052 , \8754_9053 , RIbc62a00_21, \8756_9055 , \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$210 ( \8962_9261 , RIfe9faf8_8161, \8961_9260 );
nor \U$211 ( \8963_9262 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, \8756_9055 , \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$212 ( \8964_9263 , RIdee3900_1053, \8963_9262 );
nor \U$213 ( \8965_9264 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, \8756_9055 , \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$214 ( \8966_9265 , RIdee1740_1029, \8965_9264 );
nor \U$215 ( \8967_9266 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \8756_9055 , \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$216 ( \8968_9267 , RIdedf6e8_1006, \8967_9266 );
nor \U$217 ( \8969_9268 , \8753_9052 , \8754_9053 , \8755_9054 , RIbc62988_20, \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$218 ( \8970_9269 , RIfcbd4d0_7176, \8969_9268 );
nor \U$219 ( \8971_9270 , RIbc62af0_23, \8754_9053 , \8755_9054 , RIbc62988_20, \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$220 ( \8972_9271 , RIee22678_4850, \8971_9270 );
nor \U$221 ( \8973_9272 , \8753_9052 , RIbc62a78_22, \8755_9054 , RIbc62988_20, \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$222 ( \8974_9273 , RIfc98090_6752, \8973_9272 );
nor \U$223 ( \8975_9274 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , RIbc62988_20, \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$224 ( \8976_9275 , RIee21598_4838, \8975_9274 );
nor \U$225 ( \8977_9276 , \8753_9052 , \8754_9053 , RIbc62a00_21, RIbc62988_20, \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$226 ( \8978_9277 , RIfe9fc60_8162, \8977_9276 );
nor \U$227 ( \8979_9278 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, RIbc62988_20, \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$228 ( \8980_9279 , RIded80c8_922, \8979_9278 );
nor \U$229 ( \8981_9280 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$230 ( \8982_9281 , RIfe9fdc8_8163, \8981_9280 );
nor \U$231 ( \8983_9282 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \8757_9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$232 ( \8984_9283 , RIded3be0_873, \8983_9282 );
nor \U$233 ( \8985_9284 , \8753_9052 , \8754_9053 , \8755_9054 , \8756_9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$234 ( \8986_9285 , RIded18b8_848, \8985_9284 );
nor \U$235 ( \8987_9286 , RIbc62af0_23, \8754_9053 , \8755_9054 , \8756_9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$236 ( \8988_9287 , RIdecebb8_816, \8987_9286 );
nor \U$237 ( \8989_9288 , \8753_9052 , RIbc62a78_22, \8755_9054 , \8756_9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$238 ( \8990_9289 , RIdecbeb8_784, \8989_9288 );
nor \U$239 ( \8991_9290 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , \8756_9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$240 ( \8992_9291 , RIdec91b8_752, \8991_9290 );
nor \U$241 ( \8993_9292 , \8753_9052 , \8754_9053 , RIbc62a00_21, \8756_9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$242 ( \8994_9293 , RIdeb56b8_528, \8993_9292 );
nor \U$243 ( \8995_9294 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, \8756_9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$244 ( \8996_9295 , RIde99080_336, \8995_9294 );
nor \U$245 ( \8997_9296 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, \8756_9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$246 ( \8998_9297 , RIe16f2c0_2642, \8997_9296 );
nor \U$247 ( \8999_9298 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \8756_9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$248 ( \9000_9299 , RIe15b0b8_2413, \8999_9298 );
nor \U$249 ( \9001_9300 , \8753_9052 , \8754_9053 , \8755_9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$250 ( \9002_9301 , RIe1448b8_2157, \9001_9300 );
nor \U$251 ( \9003_9302 , RIbc62af0_23, \8754_9053 , \8755_9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$252 ( \9004_9303 , RIdf392b0_2027, \9003_9302 );
nor \U$253 ( \9005_9304 , \8753_9052 , RIbc62a78_22, \8755_9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$254 ( \9006_9305 , RIdf2d910_1895, \9005_9304 );
nor \U$255 ( \9007_9306 , RIbc62af0_23, RIbc62a78_22, \8755_9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$256 ( \9008_9307 , RIdf1e190_1719, \9007_9306 );
nor \U$257 ( \9009_9308 , \8753_9052 , \8754_9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$258 ( \9010_9309 , RIdf01888_1394, \9009_9308 );
nor \U$259 ( \9011_9310 , RIbc62af0_23, \8754_9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$260 ( \9012_9311 , RIdee8388_1106, \9011_9310 );
nor \U$261 ( \9013_9312 , \8753_9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$262 ( \9014_9313 , RIdedd0f0_979, \9013_9312 );
nor \U$263 ( \9015_9314 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$264 ( \9016_9315 , RIde7efc8_209, \9015_9314 );
or \U$265 ( \9017_9316 , \8890_9189 , \8892_9191 , \8894_9193 , \8896_9195 , \8898_9197 , \8900_9199 , \8902_9201 , \8904_9203 , \8906_9205 , \8908_9207 , \8910_9209 , \8912_9211 , \8914_9213 , \8916_9215 , \8918_9217 , \8920_9219 , \8922_9221 , \8924_9223 , \8926_9225 , \8928_9227 , \8930_9229 , \8932_9231 , \8934_9233 , \8936_9235 , \8938_9237 , \8940_9239 , \8942_9241 , \8944_9243 , \8946_9245 , \8948_9247 , \8950_9249 , \8952_9251 , \8954_9253 , \8956_9255 , \8958_9257 , \8960_9259 , \8962_9261 , \8964_9263 , \8966_9265 , \8968_9267 , \8970_9269 , \8972_9271 , \8974_9273 , \8976_9275 , \8978_9277 , \8980_9279 , \8982_9281 , \8984_9283 , \8986_9285 , \8988_9287 , \8990_9289 , \8992_9291 , \8994_9293 , \8996_9295 , \8998_9297 , \9000_9299 , \9002_9301 , \9004_9303 , \9006_9305 , \9008_9307 , \9010_9309 , \9012_9311 , \9014_9313 , \9016_9315 );
or \U$266 ( \9018_9317 , \8888_9187 , \9017_9316 );
buf \U$267 ( \9019_9318 , RIbc627a8_16);
buf \U$268 ( \9020_9319 , RIbc62730_15);
buf \U$269 ( \9021_9320 , RIbc626b8_14);
buf \U$270 ( \9022_9321 , RIbc62640_13);
or \U$271 ( \9023_9322 , \9019_9318 , \9020_9319 , \9021_9320 , \9022_9321 );
buf \U$272 ( \9024_9323 , \9023_9322 );
_DC \g30c1/U$1 ( \9025 , \9018_9317 , \9024_9323 );
buf \U$273 ( \9026_9325 , \9025 );
not \U$274 ( \9027_9326 , RIbc625c8_12);
not \U$275 ( \9028_9327 , RIbc62550_11);
not \U$276 ( \9029_9328 , RIbc624d8_10);
not \U$277 ( \9030_9329 , RIbc62460_9);
not \U$278 ( \9031_9330 , RIbc623e8_8);
not \U$279 ( \9032_9331 , RIbc62370_7);
not \U$280 ( \9033_9332 , RIbc622f8_6);
nor \U$281 ( \9034_9333 , \9027_9326 , \9028_9327 , \9029_9328 , \9030_9329 , \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$282 ( \9035_9334 , RIe19e750_3180, \9034_9333 );
nor \U$283 ( \9036_9335 , RIbc625c8_12, \9028_9327 , \9029_9328 , \9030_9329 , \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$284 ( \9037_9336 , RIe19ba50_3148, \9036_9335 );
nor \U$285 ( \9038_9337 , \9027_9326 , RIbc62550_11, \9029_9328 , \9030_9329 , \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$286 ( \9039_9338 , RIfc479d8_5837, \9038_9337 );
nor \U$287 ( \9040_9339 , RIbc625c8_12, RIbc62550_11, \9029_9328 , \9030_9329 , \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$288 ( \9041_9340 , RIe198d50_3116, \9040_9339 );
nor \U$289 ( \9042_9341 , \9027_9326 , \9028_9327 , RIbc624d8_10, \9030_9329 , \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$290 ( \9043_9342 , RIfe9f558_8157, \9042_9341 );
nor \U$291 ( \9044_9343 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, \9030_9329 , \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$292 ( \9045_9344 , RIe196050_3084, \9044_9343 );
nor \U$293 ( \9046_9345 , \9027_9326 , RIbc62550_11, RIbc624d8_10, \9030_9329 , \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$294 ( \9047_9346 , RIe193350_3052, \9046_9345 );
nor \U$295 ( \9048_9347 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9030_9329 , \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$296 ( \9049_9348 , RIe190650_3020, \9048_9347 );
nor \U$297 ( \9050_9349 , \9027_9326 , \9028_9327 , \9029_9328 , RIbc62460_9, \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$298 ( \9051_9350 , RIe18ac50_2956, \9050_9349 );
nor \U$299 ( \9052_9351 , RIbc625c8_12, \9028_9327 , \9029_9328 , RIbc62460_9, \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$300 ( \9053_9352 , RIe187f50_2924, \9052_9351 );
nor \U$301 ( \9054_9353 , \9027_9326 , RIbc62550_11, \9029_9328 , RIbc62460_9, \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$302 ( \9055_9354 , RIfc47870_5836, \9054_9353 );
nor \U$303 ( \9056_9355 , RIbc625c8_12, RIbc62550_11, \9029_9328 , RIbc62460_9, \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$304 ( \9057_9356 , RIe185250_2892, \9056_9355 );
nor \U$305 ( \9058_9357 , \9027_9326 , \9028_9327 , RIbc624d8_10, RIbc62460_9, \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$306 ( \9059_9358 , RIf142ef8_5221, \9058_9357 );
nor \U$307 ( \9060_9359 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, RIbc62460_9, \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$308 ( \9061_9360 , RIe182550_2860, \9060_9359 );
nor \U$309 ( \9062_9361 , \9027_9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$310 ( \9063_9362 , RIe17f850_2828, \9062_9361 );
nor \U$311 ( \9064_9363 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9031_9330 , \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$312 ( \9065_9364 , RIe17cb50_2796, \9064_9363 );
nor \U$313 ( \9066_9365 , \9027_9326 , \9028_9327 , \9029_9328 , \9030_9329 , RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$314 ( \9067_9366 , RIfcb5208_7083, \9066_9365 );
nor \U$315 ( \9068_9367 , RIbc625c8_12, \9028_9327 , \9029_9328 , \9030_9329 , RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$316 ( \9069_9368 , RIfcbc6c0_7166, \9068_9367 );
nor \U$317 ( \9070_9369 , \9027_9326 , RIbc62550_11, \9029_9328 , \9030_9329 , RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$318 ( \9071_9370 , RIe177588_2735, \9070_9369 );
nor \U$319 ( \9072_9371 , RIbc625c8_12, RIbc62550_11, \9029_9328 , \9030_9329 , RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$320 ( \9073_9372 , RIe176610_2724, \9072_9371 );
nor \U$321 ( \9074_9373 , \9027_9326 , \9028_9327 , RIbc624d8_10, \9030_9329 , RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$322 ( \9075_9374 , RIf13fdc0_5186, \9074_9373 );
nor \U$323 ( \9076_9375 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, \9030_9329 , RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$324 ( \9077_9376 , RIfe9f3f0_8156, \9076_9375 );
nor \U$325 ( \9078_9377 , \9027_9326 , RIbc62550_11, RIbc624d8_10, \9030_9329 , RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$326 ( \9079_9378 , RIfce40f8_7617, \9078_9377 );
nor \U$327 ( \9080_9379 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9030_9329 , RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$328 ( \9081_9380 , RIfc47708_5835, \9080_9379 );
nor \U$329 ( \9082_9381 , \9027_9326 , \9028_9327 , \9029_9328 , RIbc62460_9, RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$330 ( \9083_9382 , RIfc47438_5833, \9082_9381 );
nor \U$331 ( \9084_9383 , RIbc625c8_12, \9028_9327 , \9029_9328 , RIbc62460_9, RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$332 ( \9085_9384 , RIfca15a0_6858, \9084_9383 );
nor \U$333 ( \9086_9385 , \9027_9326 , RIbc62550_11, \9029_9328 , RIbc62460_9, RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$334 ( \9087_9386 , RIfc99170_6764, \9086_9385 );
nor \U$335 ( \9088_9387 , RIbc625c8_12, RIbc62550_11, \9029_9328 , RIbc62460_9, RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$336 ( \9089_9388 , RIe1745b8_2701, \9088_9387 );
nor \U$337 ( \9090_9389 , \9027_9326 , \9028_9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$338 ( \9091_9390 , RIfc8cc90_6624, \9090_9389 );
nor \U$339 ( \9092_9391 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$340 ( \9093_9392 , RIfc556a0_5994, \9092_9391 );
nor \U$341 ( \9094_9393 , \9027_9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$342 ( \9095_9394 , RIfc7ee60_6466, \9094_9393 );
nor \U$343 ( \9096_9395 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9032_9331 , \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$344 ( \9097_9396 , RIfce8e50_7672, \9096_9395 );
nor \U$345 ( \9098_9397 , \9027_9326 , \9028_9327 , \9029_9328 , \9030_9329 , \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$346 ( \9099_9398 , RIfe9f288_8155, \9098_9397 );
nor \U$347 ( \9100_9399 , RIbc625c8_12, \9028_9327 , \9029_9328 , \9030_9329 , \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$348 ( \9101_9400 , RIe224aa8_4707, \9100_9399 );
nor \U$349 ( \9102_9401 , \9027_9326 , RIbc62550_11, \9029_9328 , \9030_9329 , \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$350 ( \9103_9402 , RIfc55808_5995, \9102_9401 );
nor \U$351 ( \9104_9403 , RIbc625c8_12, RIbc62550_11, \9029_9328 , \9030_9329 , \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$352 ( \9105_9404 , RIe221da8_4675, \9104_9403 );
nor \U$353 ( \9106_9405 , \9027_9326 , \9028_9327 , RIbc624d8_10, \9030_9329 , \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$354 ( \9107_9406 , RIfcb50a0_7082, \9106_9405 );
nor \U$355 ( \9108_9407 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, \9030_9329 , \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$356 ( \9109_9408 , RIe21f0a8_4643, \9108_9407 );
nor \U$357 ( \9110_9409 , \9027_9326 , RIbc62550_11, RIbc624d8_10, \9030_9329 , \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$358 ( \9111_9410 , RIe2196a8_4579, \9110_9409 );
nor \U$359 ( \9112_9411 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9030_9329 , \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$360 ( \9113_9412 , RIe2169a8_4547, \9112_9411 );
nor \U$361 ( \9114_9413 , \9027_9326 , \9028_9327 , \9029_9328 , RIbc62460_9, \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$362 ( \9115_9414 , RIfcbc828_7167, \9114_9413 );
nor \U$363 ( \9116_9415 , RIbc625c8_12, \9028_9327 , \9029_9328 , RIbc62460_9, \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$364 ( \9117_9416 , RIe213ca8_4515, \9116_9415 );
nor \U$365 ( \9118_9417 , \9027_9326 , RIbc62550_11, \9029_9328 , RIbc62460_9, \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$366 ( \9119_9418 , RIfc47000_5830, \9118_9417 );
nor \U$367 ( \9120_9419 , RIbc625c8_12, RIbc62550_11, \9029_9328 , RIbc62460_9, \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$368 ( \9121_9420 , RIe210fa8_4483, \9120_9419 );
nor \U$369 ( \9122_9421 , \9027_9326 , \9028_9327 , RIbc624d8_10, RIbc62460_9, \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$370 ( \9123_9422 , RIfcbc990_7168, \9122_9421 );
nor \U$371 ( \9124_9423 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, RIbc62460_9, \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$372 ( \9125_9424 , RIe20e2a8_4451, \9124_9423 );
nor \U$373 ( \9126_9425 , \9027_9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$374 ( \9127_9426 , RIe20b5a8_4419, \9126_9425 );
nor \U$375 ( \9128_9427 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9031_9330 , RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$376 ( \9129_9428 , RIe2088a8_4387, \9128_9427 );
nor \U$377 ( \9130_9429 , \9027_9326 , \9028_9327 , \9029_9328 , \9030_9329 , RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$378 ( \9131_9430 , RIfc46bc8_5827, \9130_9429 );
nor \U$379 ( \9132_9431 , RIbc625c8_12, \9028_9327 , \9029_9328 , \9030_9329 , RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$380 ( \9133_9432 , RIfcd6598_7461, \9132_9431 );
nor \U$381 ( \9134_9433 , \9027_9326 , RIbc62550_11, \9029_9328 , \9030_9329 , RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$382 ( \9135_9434 , RIe2032e0_4326, \9134_9433 );
nor \U$383 ( \9136_9435 , RIbc625c8_12, RIbc62550_11, \9029_9328 , \9030_9329 , RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$384 ( \9137_9436 , RIe2016c0_4306, \9136_9435 );
nor \U$385 ( \9138_9437 , \9027_9326 , \9028_9327 , RIbc624d8_10, \9030_9329 , RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$386 ( \9139_9438 , RIfc98ea0_6762, \9138_9437 );
nor \U$387 ( \9140_9439 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, \9030_9329 , RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$388 ( \9141_9440 , RIfc7eb90_6464, \9140_9439 );
nor \U$389 ( \9142_9441 , \9027_9326 , RIbc62550_11, RIbc624d8_10, \9030_9329 , RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$390 ( \9143_9442 , RIfce0318_7573, \9142_9441 );
nor \U$391 ( \9144_9443 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9030_9329 , RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$392 ( \9145_9444 , RIfcbcaf8_7169, \9144_9443 );
nor \U$393 ( \9146_9445 , \9027_9326 , \9028_9327 , \9029_9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$394 ( \9147_9446 , RIfc8cf60_6626, \9146_9445 );
nor \U$395 ( \9148_9447 , RIbc625c8_12, \9028_9327 , \9029_9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$396 ( \9149_9448 , RIfcb4dd0_7080, \9148_9447 );
nor \U$397 ( \9150_9449 , \9027_9326 , RIbc62550_11, \9029_9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$398 ( \9151_9450 , RIe1fd340_4258, \9150_9449 );
nor \U$399 ( \9152_9451 , RIbc625c8_12, RIbc62550_11, \9029_9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$400 ( \9153_9452 , RIe1fc260_4246, \9152_9451 );
nor \U$401 ( \9154_9453 , \9027_9326 , \9028_9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$402 ( \9155_9454 , RIf15cf38_5517, \9154_9453 );
nor \U$403 ( \9156_9455 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$404 ( \9157_9456 , RIfe9f120_8154, \9156_9455 );
nor \U$405 ( \9158_9457 , \9027_9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$406 ( \9159_9458 , RIfc7ea28_6463, \9158_9457 );
nor \U$407 ( \9160_9459 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9033_9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$408 ( \9161_9460 , RIfc8d0c8_6627, \9160_9459 );
or \U$409 ( \9162_9461 , \9035_9334 , \9037_9336 , \9039_9338 , \9041_9340 , \9043_9342 , \9045_9344 , \9047_9346 , \9049_9348 , \9051_9350 , \9053_9352 , \9055_9354 , \9057_9356 , \9059_9358 , \9061_9360 , \9063_9362 , \9065_9364 , \9067_9366 , \9069_9368 , \9071_9370 , \9073_9372 , \9075_9374 , \9077_9376 , \9079_9378 , \9081_9380 , \9083_9382 , \9085_9384 , \9087_9386 , \9089_9388 , \9091_9390 , \9093_9392 , \9095_9394 , \9097_9396 , \9099_9398 , \9101_9400 , \9103_9402 , \9105_9404 , \9107_9406 , \9109_9408 , \9111_9410 , \9113_9412 , \9115_9414 , \9117_9416 , \9119_9418 , \9121_9420 , \9123_9422 , \9125_9424 , \9127_9426 , \9129_9428 , \9131_9430 , \9133_9432 , \9135_9434 , \9137_9436 , \9139_9438 , \9141_9440 , \9143_9442 , \9145_9444 , \9147_9446 , \9149_9448 , \9151_9450 , \9153_9452 , \9155_9454 , \9157_9456 , \9159_9458 , \9161_9460 );
nor \U$410 ( \9163_9462 , \9027_9326 , \9028_9327 , \9029_9328 , \9030_9329 , \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$411 ( \9164_9463 , RIfcbcc60_7170, \9163_9462 );
nor \U$412 ( \9165_9464 , RIbc625c8_12, \9028_9327 , \9029_9328 , \9030_9329 , \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$413 ( \9166_9465 , RIfc98bd0_6760, \9165_9464 );
nor \U$414 ( \9167_9466 , \9027_9326 , RIbc62550_11, \9029_9328 , \9030_9329 , \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$415 ( \9168_9467 , RIfce2d48_7603, \9167_9466 );
nor \U$416 ( \9169_9468 , RIbc625c8_12, RIbc62550_11, \9029_9328 , \9030_9329 , \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$417 ( \9170_9469 , RIe1fb018_4233, \9169_9468 );
nor \U$418 ( \9171_9470 , \9027_9326 , \9028_9327 , RIbc624d8_10, \9030_9329 , \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$419 ( \9172_9471 , RIfc55f10_6000, \9171_9470 );
nor \U$420 ( \9173_9472 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, \9030_9329 , \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$421 ( \9174_9473 , RIfc7e8c0_6462, \9173_9472 );
nor \U$422 ( \9175_9474 , \9027_9326 , RIbc62550_11, RIbc624d8_10, \9030_9329 , \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$423 ( \9176_9475 , RIfc8d230_6628, \9175_9474 );
nor \U$424 ( \9177_9476 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9030_9329 , \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$425 ( \9178_9477 , RIe1f6590_4180, \9177_9476 );
nor \U$426 ( \9179_9478 , \9027_9326 , \9028_9327 , \9029_9328 , RIbc62460_9, \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$427 ( \9180_9479 , RIfce58e0_7634, \9179_9478 );
nor \U$428 ( \9181_9480 , RIbc625c8_12, \9028_9327 , \9029_9328 , RIbc62460_9, \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$429 ( \9182_9481 , RIfc468f8_5825, \9181_9480 );
nor \U$430 ( \9183_9482 , \9027_9326 , RIbc62550_11, \9029_9328 , RIbc62460_9, \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$431 ( \9184_9483 , RIfcc2ed0_7240, \9183_9482 );
nor \U$432 ( \9185_9484 , RIbc625c8_12, RIbc62550_11, \9029_9328 , RIbc62460_9, \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$433 ( \9186_9485 , RIe1f4100_4154, \9185_9484 );
nor \U$434 ( \9187_9486 , \9027_9326 , \9028_9327 , RIbc624d8_10, RIbc62460_9, \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$435 ( \9188_9487 , RIfceedf0_7740, \9187_9486 );
nor \U$436 ( \9189_9488 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, RIbc62460_9, \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$437 ( \9190_9489 , RIfc8d398_6629, \9189_9488 );
nor \U$438 ( \9191_9490 , \9027_9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$439 ( \9192_9491 , RIfc8d500_6630, \9191_9490 );
nor \U$440 ( \9193_9492 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9031_9330 , \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$441 ( \9194_9493 , RIe1eef70_4096, \9193_9492 );
nor \U$442 ( \9195_9494 , \9027_9326 , \9028_9327 , \9029_9328 , \9030_9329 , RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$443 ( \9196_9495 , RIe1ec810_4068, \9195_9494 );
nor \U$444 ( \9197_9496 , RIbc625c8_12, \9028_9327 , \9029_9328 , \9030_9329 , RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$445 ( \9198_9497 , RIe1e9b10_4036, \9197_9496 );
nor \U$446 ( \9199_9498 , \9027_9326 , RIbc62550_11, \9029_9328 , \9030_9329 , RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$447 ( \9200_9499 , RIe1e6e10_4004, \9199_9498 );
nor \U$448 ( \9201_9500 , RIbc625c8_12, RIbc62550_11, \9029_9328 , \9030_9329 , RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$449 ( \9202_9501 , RIe1e4110_3972, \9201_9500 );
nor \U$450 ( \9203_9502 , \9027_9326 , \9028_9327 , RIbc624d8_10, \9030_9329 , RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$451 ( \9204_9503 , RIe1e1410_3940, \9203_9502 );
nor \U$452 ( \9205_9504 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, \9030_9329 , RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$453 ( \9206_9505 , RIe1de710_3908, \9205_9504 );
nor \U$454 ( \9207_9506 , \9027_9326 , RIbc62550_11, RIbc624d8_10, \9030_9329 , RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$455 ( \9208_9507 , RIe1dba10_3876, \9207_9506 );
nor \U$456 ( \9209_9508 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9030_9329 , RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$457 ( \9210_9509 , RIe1d8d10_3844, \9209_9508 );
nor \U$458 ( \9211_9510 , \9027_9326 , \9028_9327 , \9029_9328 , RIbc62460_9, RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$459 ( \9212_9511 , RIe1d3310_3780, \9211_9510 );
nor \U$460 ( \9213_9512 , RIbc625c8_12, \9028_9327 , \9029_9328 , RIbc62460_9, RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$461 ( \9214_9513 , RIe1d0610_3748, \9213_9512 );
nor \U$462 ( \9215_9514 , \9027_9326 , RIbc62550_11, \9029_9328 , RIbc62460_9, RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$463 ( \9216_9515 , RIe1cd910_3716, \9215_9514 );
nor \U$464 ( \9217_9516 , RIbc625c8_12, RIbc62550_11, \9029_9328 , RIbc62460_9, RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$465 ( \9218_9517 , RIe1cac10_3684, \9217_9516 );
nor \U$466 ( \9219_9518 , \9027_9326 , \9028_9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$467 ( \9220_9519 , RIe1c7f10_3652, \9219_9518 );
nor \U$468 ( \9221_9520 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$469 ( \9222_9521 , RIe1c5210_3620, \9221_9520 );
nor \U$470 ( \9223_9522 , \9027_9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$471 ( \9224_9523 , RIe1c2510_3588, \9223_9522 );
nor \U$472 ( \9225_9524 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9032_9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$473 ( \9226_9525 , RIe1bf810_3556, \9225_9524 );
nor \U$474 ( \9227_9526 , \9027_9326 , \9028_9327 , \9029_9328 , \9030_9329 , \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$475 ( \9228_9527 , RIf14d0b0_5336, \9227_9526 );
nor \U$476 ( \9229_9528 , RIbc625c8_12, \9028_9327 , \9029_9328 , \9030_9329 , \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$477 ( \9230_9529 , RIfe9efb8_8153, \9229_9528 );
nor \U$478 ( \9231_9530 , \9027_9326 , RIbc62550_11, \9029_9328 , \9030_9329 , \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$479 ( \9232_9531 , RIe1ba248_3495, \9231_9530 );
nor \U$480 ( \9233_9532 , RIbc625c8_12, RIbc62550_11, \9029_9328 , \9030_9329 , \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$481 ( \9234_9533 , RIe1b8088_3471, \9233_9532 );
nor \U$482 ( \9235_9534 , \9027_9326 , \9028_9327 , RIbc624d8_10, \9030_9329 , \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$483 ( \9236_9535 , RIfec4dd0_8360, \9235_9534 );
nor \U$484 ( \9237_9536 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, \9030_9329 , \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$485 ( \9238_9537 , RIfec50a0_8362, \9237_9536 );
nor \U$486 ( \9239_9538 , \9027_9326 , RIbc62550_11, RIbc624d8_10, \9030_9329 , \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$487 ( \9240_9539 , RIe1b5ec8_3447, \9239_9538 );
nor \U$488 ( \9241_9540 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9030_9329 , \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$489 ( \9242_9541 , RIe1b46e0_3430, \9241_9540 );
nor \U$490 ( \9243_9542 , \9027_9326 , \9028_9327 , \9029_9328 , RIbc62460_9, \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$491 ( \9244_9543 , RIfcb4998_7077, \9243_9542 );
nor \U$492 ( \9245_9544 , RIbc625c8_12, \9028_9327 , \9029_9328 , RIbc62460_9, \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$493 ( \9246_9545 , RIfcb4c68_7079, \9245_9544 );
nor \U$494 ( \9247_9546 , \9027_9326 , RIbc62550_11, \9029_9328 , RIbc62460_9, \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$495 ( \9248_9547 , RIfec5370_8364, \9247_9546 );
nor \U$496 ( \9249_9548 , RIbc625c8_12, RIbc62550_11, \9029_9328 , RIbc62460_9, \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$497 ( \9250_9549 , RIfe9ee50_8152, \9249_9548 );
nor \U$498 ( \9251_9550 , \9027_9326 , \9028_9327 , RIbc624d8_10, RIbc62460_9, \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$499 ( \9252_9551 , RIfcbcdc8_7171, \9251_9550 );
nor \U$500 ( \9253_9552 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, RIbc62460_9, \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$501 ( \9254_9553 , RIfc46358_5821, \9253_9552 );
nor \U$502 ( \9255_9554 , \9027_9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$503 ( \9256_9555 , RIfec5208_8363, \9255_9554 );
nor \U$504 ( \9257_9556 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9031_9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$505 ( \9258_9557 , RIfec4f38_8361, \9257_9556 );
nor \U$506 ( \9259_9558 , \9027_9326 , \9028_9327 , \9029_9328 , \9030_9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$507 ( \9260_9559 , RIe1a9b50_3308, \9259_9558 );
nor \U$508 ( \9261_9560 , RIbc625c8_12, \9028_9327 , \9029_9328 , \9030_9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$509 ( \9262_9561 , RIe1a6e50_3276, \9261_9560 );
nor \U$510 ( \9263_9562 , \9027_9326 , RIbc62550_11, \9029_9328 , \9030_9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$511 ( \9264_9563 , RIe1a4150_3244, \9263_9562 );
nor \U$512 ( \9265_9564 , RIbc625c8_12, RIbc62550_11, \9029_9328 , \9030_9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$513 ( \9266_9565 , RIe1a1450_3212, \9265_9564 );
nor \U$514 ( \9267_9566 , \9027_9326 , \9028_9327 , RIbc624d8_10, \9030_9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$515 ( \9268_9567 , RIe18d950_2988, \9267_9566 );
nor \U$516 ( \9269_9568 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, \9030_9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$517 ( \9270_9569 , RIe179e50_2764, \9269_9568 );
nor \U$518 ( \9271_9570 , \9027_9326 , RIbc62550_11, RIbc624d8_10, \9030_9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$519 ( \9272_9571 , RIe2277a8_4739, \9271_9570 );
nor \U$520 ( \9273_9572 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9030_9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$521 ( \9274_9573 , RIe21c3a8_4611, \9273_9572 );
nor \U$522 ( \9275_9574 , \9027_9326 , \9028_9327 , \9029_9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$523 ( \9276_9575 , RIe205ba8_4355, \9275_9574 );
nor \U$524 ( \9277_9576 , RIbc625c8_12, \9028_9327 , \9029_9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$525 ( \9278_9577 , RIe1ffc08_4287, \9277_9576 );
nor \U$526 ( \9279_9578 , \9027_9326 , RIbc62550_11, \9029_9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$527 ( \9280_9579 , RIe1f8fc0_4210, \9279_9578 );
nor \U$528 ( \9281_9580 , RIbc625c8_12, RIbc62550_11, \9029_9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$529 ( \9282_9581 , RIe1f1b08_4127, \9281_9580 );
nor \U$530 ( \9283_9582 , \9027_9326 , \9028_9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$531 ( \9284_9583 , RIe1d6010_3812, \9283_9582 );
nor \U$532 ( \9285_9584 , RIbc625c8_12, \9028_9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$533 ( \9286_9585 , RIe1bcb10_3524, \9285_9584 );
nor \U$534 ( \9287_9586 , \9027_9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$535 ( \9288_9587 , RIe1af988_3375, \9287_9586 );
nor \U$536 ( \9289_9588 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$537 ( \9290_9589 , RIe171fc0_2674, \9289_9588 );
or \U$538 ( \9291_9590 , \9164_9463 , \9166_9465 , \9168_9467 , \9170_9469 , \9172_9471 , \9174_9473 , \9176_9475 , \9178_9477 , \9180_9479 , \9182_9481 , \9184_9483 , \9186_9485 , \9188_9487 , \9190_9489 , \9192_9491 , \9194_9493 , \9196_9495 , \9198_9497 , \9200_9499 , \9202_9501 , \9204_9503 , \9206_9505 , \9208_9507 , \9210_9509 , \9212_9511 , \9214_9513 , \9216_9515 , \9218_9517 , \9220_9519 , \9222_9521 , \9224_9523 , \9226_9525 , \9228_9527 , \9230_9529 , \9232_9531 , \9234_9533 , \9236_9535 , \9238_9537 , \9240_9539 , \9242_9541 , \9244_9543 , \9246_9545 , \9248_9547 , \9250_9549 , \9252_9551 , \9254_9553 , \9256_9555 , \9258_9557 , \9260_9559 , \9262_9561 , \9264_9563 , \9266_9565 , \9268_9567 , \9270_9569 , \9272_9571 , \9274_9573 , \9276_9575 , \9278_9577 , \9280_9579 , \9282_9581 , \9284_9583 , \9286_9585 , \9288_9587 , \9290_9589 );
or \U$539 ( \9292_9591 , \9162_9461 , \9291_9590 );
buf \U$540 ( \9293_9592 , RIbc62280_5);
buf \U$541 ( \9294_9593 , RIbc62208_4);
buf \U$542 ( \9295_9594 , RIbc62190_3);
buf \U$543 ( \9296_9595 , RIbc62118_2);
or \U$544 ( \9297_9596 , \9293_9592 , \9294_9593 , \9295_9594 , \9296_9595 );
buf \U$545 ( \9298_9597 , \9297_9596 );
_DC \g41ee/U$1 ( \9299 , \9292_9591 , \9298_9597 );
buf \U$546 ( \9300_9599 , \9299 );
xor \U$547 ( \9301_9600 , \9026_9325 , \9300_9599 );
and \U$548 ( \9302_9601 , RIdec6080_717, \8760_9059 );
and \U$549 ( \9303_9602 , RIdec3380_685, \8762_9061 );
and \U$550 ( \9304_9603 , RIee204b8_4826, \8764_9063 );
and \U$551 ( \9305_9604 , RIdec0680_653, \8766_9065 );
and \U$552 ( \9306_9605 , RIfcd70d8_7469, \8768_9067 );
and \U$553 ( \9307_9606 , RIdebd980_621, \8770_9069 );
and \U$554 ( \9308_9607 , RIdebac80_589, \8772_9071 );
and \U$555 ( \9309_9608 , RIdeb7f80_557, \8774_9073 );
and \U$556 ( \9310_9609 , RIfcbe448_7187, \8776_9075 );
and \U$557 ( \9311_9610 , RIdeb2580_493, \8778_9077 );
and \U$558 ( \9312_9611 , RIfcb3480_7062, \8780_9079 );
and \U$559 ( \9313_9612 , RIdeaf880_461, \8782_9081 );
and \U$560 ( \9314_9613 , RIfc43928_5791, \8784_9083 );
and \U$561 ( \9315_9614 , RIdeac1a8_429, \8786_9085 );
and \U$562 ( \9316_9615 , RIdea58a8_397, \8788_9087 );
and \U$563 ( \9317_9616 , RIde9efa8_365, \8790_9089 );
and \U$564 ( \9318_9617 , RIfcd88c0_7486, \8792_9091 );
and \U$565 ( \9319_9618 , RIee1c408_4780, \8794_9093 );
and \U$566 ( \9320_9619 , RIfcc77f0_7292, \8796_9095 );
and \U$567 ( \9321_9620 , RIfea04d0_8168, \8798_9097 );
and \U$568 ( \9322_9621 , RIde92438_303, \8800_9099 );
and \U$569 ( \9323_9622 , RIde8ec70_286, \8802_9101 );
and \U$570 ( \9324_9623 , RIde8aad0_266, \8804_9103 );
and \U$571 ( \9325_9624 , RIde86930_246, \8806_9105 );
and \U$572 ( \9326_9625 , RIfca31c0_6878, \8808_9107 );
and \U$573 ( \9327_9626 , RIfc59a20_6042, \8810_9109 );
and \U$574 ( \9328_9627 , RIfcd1de0_7410, \8812_9111 );
and \U$575 ( \9329_9628 , RIfc91448_6675, \8814_9113 );
and \U$576 ( \9330_9629 , RIfc97280_6742, \8816_9115 );
and \U$577 ( \9331_9630 , RIe16c188_2607, \8818_9117 );
and \U$578 ( \9332_9631 , RIfc97118_6741, \8820_9119 );
and \U$579 ( \9333_9632 , RIe168948_2567, \8822_9121 );
and \U$580 ( \9334_9633 , RIe166080_2538, \8824_9123 );
and \U$581 ( \9335_9634 , RIe163380_2506, \8826_9125 );
and \U$582 ( \9336_9635 , RIee37ac8_5092, \8828_9127 );
and \U$583 ( \9337_9636 , RIe160680_2474, \8830_9129 );
and \U$584 ( \9338_9637 , RIfcd1c78_7409, \8832_9131 );
and \U$585 ( \9339_9638 , RIe15d980_2442, \8834_9133 );
and \U$586 ( \9340_9639 , RIe157f80_2378, \8836_9135 );
and \U$587 ( \9341_9640 , RIe155280_2346, \8838_9137 );
and \U$588 ( \9342_9641 , RIfc3f530_5746, \8840_9139 );
and \U$589 ( \9343_9642 , RIe152580_2314, \8842_9141 );
and \U$590 ( \9344_9643 , RIee35368_5064, \8844_9143 );
and \U$591 ( \9345_9644 , RIe14f880_2282, \8846_9145 );
and \U$592 ( \9346_9645 , RIfc7a3d8_6413, \8848_9147 );
and \U$593 ( \9347_9646 , RIe14cb80_2250, \8850_9149 );
and \U$594 ( \9348_9647 , RIe149e80_2218, \8852_9151 );
and \U$595 ( \9349_9648 , RIe147180_2186, \8854_9153 );
and \U$596 ( \9350_9649 , RIfc42b18_5781, \8856_9155 );
and \U$597 ( \9351_9650 , RIfc7a270_6412, \8858_9157 );
and \U$598 ( \9352_9651 , RIfc5a560_6050, \8860_9159 );
and \U$599 ( \9353_9652 , RIfc96b78_6737, \8862_9161 );
and \U$600 ( \9354_9653 , RIfea6fb0_8216, \8864_9163 );
and \U$601 ( \9355_9654 , RIe13f5c0_2098, \8866_9165 );
and \U$602 ( \9356_9655 , RIdf3d4c8_2074, \8868_9167 );
and \U$603 ( \9357_9656 , RIdf3b038_2048, \8870_9169 );
and \U$604 ( \9358_9657 , RIfce5bb0_7636, \8872_9171 );
and \U$605 ( \9359_9658 , RIee2fc38_5002, \8874_9173 );
and \U$606 ( \9360_9659 , RIfc91cb8_6681, \8876_9175 );
and \U$607 ( \9361_9660 , RIee2d910_4977, \8878_9177 );
and \U$608 ( \9362_9661 , RIdf362e0_1993, \8880_9179 );
and \U$609 ( \9363_9662 , RIdf33e50_1967, \8882_9181 );
and \U$610 ( \9364_9663 , RIdf31c90_1943, \8884_9183 );
and \U$611 ( \9365_9664 , RIdf2fda0_1921, \8886_9185 );
or \U$612 ( \9366_9665 , \9302_9601 , \9303_9602 , \9304_9603 , \9305_9604 , \9306_9605 , \9307_9606 , \9308_9607 , \9309_9608 , \9310_9609 , \9311_9610 , \9312_9611 , \9313_9612 , \9314_9613 , \9315_9614 , \9316_9615 , \9317_9616 , \9318_9617 , \9319_9618 , \9320_9619 , \9321_9620 , \9322_9621 , \9323_9622 , \9324_9623 , \9325_9624 , \9326_9625 , \9327_9626 , \9328_9627 , \9329_9628 , \9330_9629 , \9331_9630 , \9332_9631 , \9333_9632 , \9334_9633 , \9335_9634 , \9336_9635 , \9337_9636 , \9338_9637 , \9339_9638 , \9340_9639 , \9341_9640 , \9342_9641 , \9343_9642 , \9344_9643 , \9345_9644 , \9346_9645 , \9347_9646 , \9348_9647 , \9349_9648 , \9350_9649 , \9351_9650 , \9352_9651 , \9353_9652 , \9354_9653 , \9355_9654 , \9356_9655 , \9357_9656 , \9358_9657 , \9359_9658 , \9360_9659 , \9361_9660 , \9362_9661 , \9363_9662 , \9364_9663 , \9365_9664 );
and \U$613 ( \9367_9666 , RIfc43658_5789, \8889_9188 );
and \U$614 ( \9368_9667 , RIfc59e58_6045, \8891_9190 );
and \U$615 ( \9369_9668 , RIfc96fb0_6740, \8893_9192 );
and \U$616 ( \9370_9669 , RIfc7ac48_6419, \8895_9194 );
and \U$617 ( \9371_9670 , RIfea0368_8167, \8897_9196 );
and \U$618 ( \9372_9671 , RIdf28bb8_1840, \8899_9198 );
and \U$619 ( \9373_9672 , RIdf26cc8_1818, \8901_9200 );
and \U$620 ( \9374_9673 , RIdf25210_1799, \8903_9202 );
and \U$621 ( \9375_9674 , RIfc91718_6677, \8905_9204 );
and \U$622 ( \9376_9675 , RIfcb3318_7061, \8907_9206 );
and \U$623 ( \9377_9676 , RIfc919e8_6679, \8909_9208 );
and \U$624 ( \9378_9677 , RIfc91880_6678, \8911_9210 );
and \U$625 ( \9379_9678 , RIfc430b8_5785, \8913_9212 );
and \U$626 ( \9380_9679 , RIdf20350_1743, \8915_9214 );
and \U$627 ( \9381_9680 , RIfc7a978_6417, \8917_9216 );
and \U$628 ( \9382_9681 , RIdf19e10_1671, \8919_9218 );
and \U$629 ( \9383_9682 , RIdf17c50_1647, \8921_9220 );
and \U$630 ( \9384_9683 , RIdf14f50_1615, \8923_9222 );
and \U$631 ( \9385_9684 , RIdf12250_1583, \8925_9224 );
and \U$632 ( \9386_9685 , RIdf0f550_1551, \8927_9226 );
and \U$633 ( \9387_9686 , RIdf0c850_1519, \8929_9228 );
and \U$634 ( \9388_9687 , RIdf09b50_1487, \8931_9230 );
and \U$635 ( \9389_9688 , RIdf06e50_1455, \8933_9232 );
and \U$636 ( \9390_9689 , RIdf04150_1423, \8935_9234 );
and \U$637 ( \9391_9690 , RIdefe750_1359, \8937_9236 );
and \U$638 ( \9392_9691 , RIdefba50_1327, \8939_9238 );
and \U$639 ( \9393_9692 , RIdef8d50_1295, \8941_9240 );
and \U$640 ( \9394_9693 , RIdef6050_1263, \8943_9242 );
and \U$641 ( \9395_9694 , RIdef3350_1231, \8945_9244 );
and \U$642 ( \9396_9695 , RIdef0650_1199, \8947_9246 );
and \U$643 ( \9397_9696 , RIdeed950_1167, \8949_9248 );
and \U$644 ( \9398_9697 , RIdeeac50_1135, \8951_9250 );
and \U$645 ( \9399_9698 , RIfcd1b10_7408, \8953_9252 );
and \U$646 ( \9400_9699 , RIfc968a8_6735, \8955_9254 );
and \U$647 ( \9401_9700 , RIfc91f88_6683, \8957_9256 );
and \U$648 ( \9402_9701 , RIfcdfc10_7568, \8959_9258 );
and \U$649 ( \9403_9702 , RIfea99e0_8246, \8961_9260 );
and \U$650 ( \9404_9703 , RIdee3630_1051, \8963_9262 );
and \U$651 ( \9405_9704 , RIdee1308_1026, \8965_9264 );
and \U$652 ( \9406_9705 , RIdedf2b0_1003, \8967_9266 );
and \U$653 ( \9407_9706 , RIfcc7d90_7296, \8969_9268 );
and \U$654 ( \9408_9707 , RIfcd85f0_7484, \8971_9270 );
and \U$655 ( \9409_9708 , RIfce3888_7611, \8973_9272 );
and \U$656 ( \9410_9709 , RIfc5a830_6052, \8975_9274 );
and \U$657 ( \9411_9710 , RIdeda3f0_947, \8977_9276 );
and \U$658 ( \9412_9711 , RIfea9878_8245, \8979_9278 );
and \U$659 ( \9413_9712 , RIded5f08_898, \8981_9280 );
and \U$660 ( \9414_9713 , RIded37a8_870, \8983_9282 );
and \U$661 ( \9415_9714 , RIded1480_845, \8985_9284 );
and \U$662 ( \9416_9715 , RIdece780_813, \8987_9286 );
and \U$663 ( \9417_9716 , RIdecba80_781, \8989_9288 );
and \U$664 ( \9418_9717 , RIdec8d80_749, \8991_9290 );
and \U$665 ( \9419_9718 , RIdeb5280_525, \8993_9292 );
and \U$666 ( \9420_9719 , RIde986a8_333, \8995_9294 );
and \U$667 ( \9421_9720 , RIe16ee88_2639, \8997_9296 );
and \U$668 ( \9422_9721 , RIe15ac80_2410, \8999_9298 );
and \U$669 ( \9423_9722 , RIe144480_2154, \9001_9300 );
and \U$670 ( \9424_9723 , RIdf38e78_2024, \9003_9302 );
and \U$671 ( \9425_9724 , RIdf2d4d8_1892, \9005_9304 );
and \U$672 ( \9426_9725 , RIdf1dd58_1716, \9007_9306 );
and \U$673 ( \9427_9726 , RIdf01450_1391, \9009_9308 );
and \U$674 ( \9428_9727 , RIdee7f50_1103, \9011_9310 );
and \U$675 ( \9429_9728 , RIdedccb8_976, \9013_9312 );
and \U$676 ( \9430_9729 , RIde7e5f0_206, \9015_9314 );
or \U$677 ( \9431_9730 , \9367_9666 , \9368_9667 , \9369_9668 , \9370_9669 , \9371_9670 , \9372_9671 , \9373_9672 , \9374_9673 , \9375_9674 , \9376_9675 , \9377_9676 , \9378_9677 , \9379_9678 , \9380_9679 , \9381_9680 , \9382_9681 , \9383_9682 , \9384_9683 , \9385_9684 , \9386_9685 , \9387_9686 , \9388_9687 , \9389_9688 , \9390_9689 , \9391_9690 , \9392_9691 , \9393_9692 , \9394_9693 , \9395_9694 , \9396_9695 , \9397_9696 , \9398_9697 , \9399_9698 , \9400_9699 , \9401_9700 , \9402_9701 , \9403_9702 , \9404_9703 , \9405_9704 , \9406_9705 , \9407_9706 , \9408_9707 , \9409_9708 , \9410_9709 , \9411_9710 , \9412_9711 , \9413_9712 , \9414_9713 , \9415_9714 , \9416_9715 , \9417_9716 , \9418_9717 , \9419_9718 , \9420_9719 , \9421_9720 , \9422_9721 , \9423_9722 , \9424_9723 , \9425_9724 , \9426_9725 , \9427_9726 , \9428_9727 , \9429_9728 , \9430_9729 );
or \U$678 ( \9432_9731 , \9366_9665 , \9431_9730 );
_DC \g3146/U$1 ( \9433 , \9432_9731 , \9024_9323 );
buf \U$679 ( \9434_9733 , \9433 );
and \U$680 ( \9435_9734 , RIe19e318_3177, \9034_9333 );
and \U$681 ( \9436_9735 , RIe19b618_3145, \9036_9335 );
and \U$682 ( \9437_9736 , RIfc8f3f0_6652, \9038_9337 );
and \U$683 ( \9438_9737 , RIe198918_3113, \9040_9339 );
and \U$684 ( \9439_9738 , RIf144b18_5241, \9042_9341 );
and \U$685 ( \9440_9739 , RIe195c18_3081, \9044_9343 );
and \U$686 ( \9441_9740 , RIe192f18_3049, \9046_9345 );
and \U$687 ( \9442_9741 , RIe190218_3017, \9048_9347 );
and \U$688 ( \9443_9742 , RIe18a818_2953, \9050_9349 );
and \U$689 ( \9444_9743 , RIe187b18_2921, \9052_9351 );
and \U$690 ( \9445_9744 , RIf143d08_5231, \9054_9353 );
and \U$691 ( \9446_9745 , RIe184e18_2889, \9056_9355 );
and \U$692 ( \9447_9746 , RIfcb3cf0_7068, \9058_9357 );
and \U$693 ( \9448_9747 , RIe182118_2857, \9060_9359 );
and \U$694 ( \9449_9748 , RIe17f418_2825, \9062_9361 );
and \U$695 ( \9450_9749 , RIe17c718_2793, \9064_9363 );
and \U$696 ( \9451_9750 , RIfc448a0_5802, \9066_9365 );
and \U$697 ( \9452_9751 , RIf141170_5200, \9068_9367 );
and \U$698 ( \9453_9752 , RIfc7c9d0_6440, \9070_9369 );
and \U$699 ( \9454_9753 , RIfea0098_8165, \9072_9371 );
and \U$700 ( \9455_9754 , RIfc57e00_6022, \9074_9373 );
and \U$701 ( \9456_9755 , RIf13f550_5180, \9076_9375 );
and \U$702 ( \9457_9756 , RIfcd6e08_7467, \9078_9377 );
and \U$703 ( \9458_9757 , RIee3d900_5159, \9080_9379 );
and \U$704 ( \9459_9758 , RIfc8f6c0_6654, \9082_9381 );
and \U$705 ( \9460_9759 , RIfce0048_7571, \9084_9383 );
and \U$706 ( \9461_9760 , RIfca27e8_6871, \9086_9385 );
and \U$707 ( \9462_9761 , RIe1742e8_2699, \9088_9387 );
and \U$708 ( \9463_9762 , RIfc7c700_6438, \9090_9389 );
and \U$709 ( \9464_9763 , RIfc8f990_6656, \9092_9391 );
and \U$710 ( \9465_9764 , RIfce9828_7679, \9094_9393 );
and \U$711 ( \9466_9765 , RIfc583a0_6026, \9096_9395 );
and \U$712 ( \9467_9766 , RIf16cdc0_5698, \9098_9397 );
and \U$713 ( \9468_9767 , RIe224670_4704, \9100_9399 );
and \U$714 ( \9469_9768 , RIf16c118_5689, \9102_9401 );
and \U$715 ( \9470_9769 , RIe221970_4672, \9104_9403 );
and \U$716 ( \9471_9770 , RIfc58508_6027, \9106_9405 );
and \U$717 ( \9472_9771 , RIe21ec70_4640, \9108_9407 );
and \U$718 ( \9473_9772 , RIe219270_4576, \9110_9409 );
and \U$719 ( \9474_9773 , RIe216570_4544, \9112_9411 );
and \U$720 ( \9475_9774 , RIfc3ff08_5753, \9114_9413 );
and \U$721 ( \9476_9775 , RIe213870_4512, \9116_9415 );
and \U$722 ( \9477_9776 , RIf1696e8_5659, \9118_9417 );
and \U$723 ( \9478_9777 , RIe210b70_4480, \9120_9419 );
and \U$724 ( \9479_9778 , RIfc58940_6030, \9122_9421 );
and \U$725 ( \9480_9779 , RIe20de70_4448, \9124_9423 );
and \U$726 ( \9481_9780 , RIe20b170_4416, \9126_9425 );
and \U$727 ( \9482_9781 , RIe208470_4384, \9128_9427 );
and \U$728 ( \9483_9782 , RIfc8fc60_6658, \9130_9429 );
and \U$729 ( \9484_9783 , RIfc97820_6746, \9132_9431 );
and \U$730 ( \9485_9784 , RIe202ea8_4323, \9134_9433 );
and \U$731 ( \9486_9785 , RIe201288_4303, \9136_9435 );
and \U$732 ( \9487_9786 , RIfcc27c8_7235, \9138_9437 );
and \U$733 ( \9488_9787 , RIfcdfee0_7570, \9140_9439 );
and \U$734 ( \9489_9788 , RIfc44198_5797, \9142_9441 );
and \U$735 ( \9490_9789 , RIfc58670_6028, \9144_9443 );
and \U$736 ( \9491_9790 , RIf1608e0_5558, \9146_9445 );
and \U$737 ( \9492_9791 , RIf15e9f0_5536, \9148_9447 );
and \U$738 ( \9493_9792 , RIfe9ff30_8164, \9150_9449 );
and \U$739 ( \9494_9793 , RIe1fc0f8_4245, \9152_9451 );
and \U$740 ( \9495_9794 , RIfc7be90_6432, \9154_9453 );
and \U$741 ( \9496_9795 , RIf15bb88_5503, \9156_9455 );
and \U$742 ( \9497_9796 , RIfcd8cf8_7489, \9158_9457 );
and \U$743 ( \9498_9797 , RIfcd8e60_7490, \9160_9459 );
or \U$744 ( \9499_9798 , \9435_9734 , \9436_9735 , \9437_9736 , \9438_9737 , \9439_9738 , \9440_9739 , \9441_9740 , \9442_9741 , \9443_9742 , \9444_9743 , \9445_9744 , \9446_9745 , \9447_9746 , \9448_9747 , \9449_9748 , \9450_9749 , \9451_9750 , \9452_9751 , \9453_9752 , \9454_9753 , \9455_9754 , \9456_9755 , \9457_9756 , \9458_9757 , \9459_9758 , \9460_9759 , \9461_9760 , \9462_9761 , \9463_9762 , \9464_9763 , \9465_9764 , \9466_9765 , \9467_9766 , \9468_9767 , \9469_9768 , \9470_9769 , \9471_9770 , \9472_9771 , \9473_9772 , \9474_9773 , \9475_9774 , \9476_9775 , \9477_9776 , \9478_9777 , \9479_9778 , \9480_9779 , \9481_9780 , \9482_9781 , \9483_9782 , \9484_9783 , \9485_9784 , \9486_9785 , \9487_9786 , \9488_9787 , \9489_9788 , \9490_9789 , \9491_9790 , \9492_9791 , \9493_9792 , \9494_9793 , \9495_9794 , \9496_9795 , \9497_9796 , \9498_9797 );
and \U$745 ( \9500_9799 , RIfca2d88_6875, \9163_9462 );
and \U$746 ( \9501_9800 , RIfcbdea8_7183, \9165_9464 );
and \U$747 ( \9502_9801 , RIfcb3a20_7066, \9167_9466 );
and \U$748 ( \9503_9802 , RIe1fabe0_4230, \9169_9468 );
and \U$749 ( \9504_9803 , RIfc90098_6661, \9171_9470 );
and \U$750 ( \9505_9804 , RIfc90200_6662, \9173_9472 );
and \U$751 ( \9506_9805 , RIfcd20b0_7412, \9175_9474 );
and \U$752 ( \9507_9806 , RIe1f6158_4177, \9177_9476 );
and \U$753 ( \9508_9807 , RIfc904d0_6664, \9179_9478 );
and \U$754 ( \9509_9808 , RIfca2ef0_6876, \9181_9480 );
and \U$755 ( \9510_9809 , RIfc97550_6744, \9183_9482 );
and \U$756 ( \9511_9810 , RIe1f3e30_4152, \9185_9484 );
and \U$757 ( \9512_9811 , RIfc59048_6035, \9187_9486 );
and \U$758 ( \9513_9812 , RIfc907a0_6666, \9189_9488 );
and \U$759 ( \9514_9813 , RIfc90638_6665, \9191_9490 );
and \U$760 ( \9515_9814 , RIe1eeb38_4093, \9193_9492 );
and \U$761 ( \9516_9815 , RIe1ec3d8_4065, \9195_9494 );
and \U$762 ( \9517_9816 , RIe1e96d8_4033, \9197_9496 );
and \U$763 ( \9518_9817 , RIe1e69d8_4001, \9199_9498 );
and \U$764 ( \9519_9818 , RIe1e3cd8_3969, \9201_9500 );
and \U$765 ( \9520_9819 , RIe1e0fd8_3937, \9203_9502 );
and \U$766 ( \9521_9820 , RIe1de2d8_3905, \9205_9504 );
and \U$767 ( \9522_9821 , RIe1db5d8_3873, \9207_9506 );
and \U$768 ( \9523_9822 , RIe1d88d8_3841, \9209_9508 );
and \U$769 ( \9524_9823 , RIe1d2ed8_3777, \9211_9510 );
and \U$770 ( \9525_9824 , RIe1d01d8_3745, \9213_9512 );
and \U$771 ( \9526_9825 , RIe1cd4d8_3713, \9215_9514 );
and \U$772 ( \9527_9826 , RIe1ca7d8_3681, \9217_9516 );
and \U$773 ( \9528_9827 , RIe1c7ad8_3649, \9219_9518 );
and \U$774 ( \9529_9828 , RIe1c4dd8_3617, \9221_9520 );
and \U$775 ( \9530_9829 , RIe1c20d8_3585, \9223_9522 );
and \U$776 ( \9531_9830 , RIe1bf3d8_3553, \9225_9524 );
and \U$777 ( \9532_9831 , RIfcc73b8_7289, \9227_9526 );
and \U$778 ( \9533_9832 , RIfce3cc0_7614, \9229_9528 );
and \U$779 ( \9534_9833 , RIe1b9e10_3492, \9231_9530 );
and \U$780 ( \9535_9834 , RIe1b7c50_3468, \9233_9532 );
and \U$781 ( \9536_9835 , RIfcd6f70_7468, \9235_9534 );
and \U$782 ( \9537_9836 , RIf149e10_5300, \9237_9536 );
and \U$783 ( \9538_9837 , RIe1b5a90_3444, \9239_9538 );
and \U$784 ( \9539_9838 , RIfea0200_8166, \9241_9540 );
and \U$785 ( \9540_9839 , RIfc90bd8_6669, \9243_9542 );
and \U$786 ( \9541_9840 , RIfcdfd78_7569, \9245_9544 );
and \U$787 ( \9542_9841 , RIe1b2ef8_3413, \9247_9546 );
and \U$788 ( \9543_9842 , RIe1b15a8_3395, \9249_9548 );
and \U$789 ( \9544_9843 , RIfc973e8_6743, \9251_9550 );
and \U$790 ( \9545_9844 , RIfcc7520_7290, \9253_9552 );
and \U$791 ( \9546_9845 , RIe1acdf0_3344, \9255_9554 );
and \U$792 ( \9547_9846 , RIe1ab608_3327, \9257_9556 );
and \U$793 ( \9548_9847 , RIe1a9718_3305, \9259_9558 );
and \U$794 ( \9549_9848 , RIe1a6a18_3273, \9261_9560 );
and \U$795 ( \9550_9849 , RIe1a3d18_3241, \9263_9562 );
and \U$796 ( \9551_9850 , RIe1a1018_3209, \9265_9564 );
and \U$797 ( \9552_9851 , RIe18d518_2985, \9267_9566 );
and \U$798 ( \9553_9852 , RIe179a18_2761, \9269_9568 );
and \U$799 ( \9554_9853 , RIe227370_4736, \9271_9570 );
and \U$800 ( \9555_9854 , RIe21bf70_4608, \9273_9572 );
and \U$801 ( \9556_9855 , RIe205770_4352, \9275_9574 );
and \U$802 ( \9557_9856 , RIe1ff7d0_4284, \9277_9576 );
and \U$803 ( \9558_9857 , RIe1f8b88_4207, \9279_9578 );
and \U$804 ( \9559_9858 , RIe1f16d0_4124, \9281_9580 );
and \U$805 ( \9560_9859 , RIe1d5bd8_3809, \9283_9582 );
and \U$806 ( \9561_9860 , RIe1bc6d8_3521, \9285_9584 );
and \U$807 ( \9562_9861 , RIe1af550_3372, \9287_9586 );
and \U$808 ( \9563_9862 , RIe171b88_2671, \9289_9588 );
or \U$809 ( \9564_9863 , \9500_9799 , \9501_9800 , \9502_9801 , \9503_9802 , \9504_9803 , \9505_9804 , \9506_9805 , \9507_9806 , \9508_9807 , \9509_9808 , \9510_9809 , \9511_9810 , \9512_9811 , \9513_9812 , \9514_9813 , \9515_9814 , \9516_9815 , \9517_9816 , \9518_9817 , \9519_9818 , \9520_9819 , \9521_9820 , \9522_9821 , \9523_9822 , \9524_9823 , \9525_9824 , \9526_9825 , \9527_9826 , \9528_9827 , \9529_9828 , \9530_9829 , \9531_9830 , \9532_9831 , \9533_9832 , \9534_9833 , \9535_9834 , \9536_9835 , \9537_9836 , \9538_9837 , \9539_9838 , \9540_9839 , \9541_9840 , \9542_9841 , \9543_9842 , \9544_9843 , \9545_9844 , \9546_9845 , \9547_9846 , \9548_9847 , \9549_9848 , \9550_9849 , \9551_9850 , \9552_9851 , \9553_9852 , \9554_9853 , \9555_9854 , \9556_9855 , \9557_9856 , \9558_9857 , \9559_9858 , \9560_9859 , \9561_9860 , \9562_9861 , \9563_9862 );
or \U$810 ( \9565_9864 , \9499_9798 , \9564_9863 );
_DC \g4273/U$1 ( \9566 , \9565_9864 , \9298_9597 );
buf \U$811 ( \9567_9866 , \9566 );
and \U$812 ( \9568_9867 , \9434_9733 , \9567_9866 );
and \U$813 ( \9569_9868 , RIdec5108_706, \8760_9059 );
and \U$814 ( \9570_9869 , RIdec2408_674, \8762_9061 );
and \U$815 ( \9571_9870 , RIfc93608_6699, \8764_9063 );
and \U$816 ( \9572_9871 , RIdebf708_642, \8766_9065 );
and \U$817 ( \9573_9872 , RIfc934a0_6698, \8768_9067 );
and \U$818 ( \9574_9873 , RIdebca08_610, \8770_9069 );
and \U$819 ( \9575_9874 , RIdeb9d08_578, \8772_9071 );
and \U$820 ( \9576_9875 , RIdeb7008_546, \8774_9073 );
and \U$821 ( \9577_9876 , RIfcdf7d8_7565, \8776_9075 );
and \U$822 ( \9578_9877 , RIdeb1608_482, \8778_9077 );
and \U$823 ( \9579_9878 , RIfc78218_6389, \8780_9079 );
and \U$824 ( \9580_9879 , RIdeae908_450, \8782_9081 );
and \U$825 ( \9581_9880 , RIfcc8498_7301, \8784_9083 );
and \U$826 ( \9582_9881 , RIdea9d90_418, \8786_9085 );
and \U$827 ( \9583_9882 , RIdea3490_386, \8788_9087 );
and \U$828 ( \9584_9883 , RIde9cb90_354, \8790_9089 );
and \U$829 ( \9585_9884 , RIee1cc78_4786, \8792_9091 );
and \U$830 ( \9586_9885 , RIee1bb98_4774, \8794_9093 );
and \U$831 ( \9587_9886 , RIee1b328_4768, \8796_9095 );
and \U$832 ( \9588_9887 , RIee1aab8_4762, \8798_9097 );
and \U$833 ( \9589_9888 , RIde909f8_295, \8800_9099 );
and \U$834 ( \9590_9889 , RIde8d578_279, \8802_9101 );
and \U$835 ( \9591_9890 , RIfea8ea0_8238, \8804_9103 );
and \U$836 ( \9592_9891 , RIde85238_239, \8806_9105 );
and \U$837 ( \9593_9892 , RIde813e0_220, \8808_9107 );
and \U$838 ( \9594_9893 , RIfc938d8_6701, \8810_9109 );
and \U$839 ( \9595_9894 , RIfce5e80_7638, \8812_9111 );
and \U$840 ( \9596_9895 , RIfcbfd98_7205, \8814_9113 );
and \U$841 ( \9597_9896 , RIfce8ce8_7671, \8816_9115 );
and \U$842 ( \9598_9897 , RIe16b4e0_2598, \8818_9117 );
and \U$843 ( \9599_9898 , RIfea8d38_8237, \8820_9119 );
and \U$844 ( \9600_9899 , RIfea9f80_8250, \8822_9121 );
and \U$845 ( \9601_9900 , RIe165108_2527, \8824_9123 );
and \U$846 ( \9602_9901 , RIe162408_2495, \8826_9125 );
and \U$847 ( \9603_9902 , RIfc779a8_6383, \8828_9127 );
and \U$848 ( \9604_9903 , RIe15f708_2463, \8830_9129 );
and \U$849 ( \9605_9904 , RIfe9dc08_8139, \8832_9131 );
and \U$850 ( \9606_9905 , RIe15ca08_2431, \8834_9133 );
and \U$851 ( \9607_9906 , RIe157008_2367, \8836_9135 );
and \U$852 ( \9608_9907 , RIe154308_2335, \8838_9137 );
and \U$853 ( \9609_9908 , RIfea7550_8220, \8840_9139 );
and \U$854 ( \9610_9909 , RIe151608_2303, \8842_9141 );
and \U$855 ( \9611_9910 , RIfcd6160_7458, \8844_9143 );
and \U$856 ( \9612_9911 , RIe14e908_2271, \8846_9145 );
and \U$857 ( \9613_9912 , RIfcd1408_7403, \8848_9147 );
and \U$858 ( \9614_9913 , RIe14bc08_2239, \8850_9149 );
and \U$859 ( \9615_9914 , RIe148f08_2207, \8852_9151 );
and \U$860 ( \9616_9915 , RIe146208_2175, \8854_9153 );
and \U$861 ( \9617_9916 , RIfceb718_7701, \8856_9155 );
and \U$862 ( \9618_9917 , RIfcb19c8_7043, \8858_9157 );
and \U$863 ( \9619_9918 , RIfc93e78_6705, \8860_9159 );
and \U$864 ( \9620_9919 , RIfce7938_7657, \8862_9161 );
and \U$865 ( \9621_9920 , RIe140da8_2115, \8864_9163 );
and \U$866 ( \9622_9921 , RIdf3ecb0_2091, \8866_9165 );
and \U$867 ( \9623_9922 , RIdf3c988_2066, \8868_9167 );
and \U$868 ( \9624_9923 , RIfe9daa0_8138, \8870_9169 );
and \U$869 ( \9625_9924 , RIfce8478_7665, \8872_9171 );
and \U$870 ( \9626_9925 , RIfcdbf98_7525, \8874_9173 );
and \U$871 ( \9627_9926 , RIfc776d8_6381, \8876_9175 );
and \U$872 ( \9628_9927 , RIfc93fe0_6706, \8878_9177 );
and \U$873 ( \9629_9928 , RIdf354d0_1983, \8880_9179 );
and \U$874 ( \9630_9929 , RIdf33040_1957, \8882_9181 );
and \U$875 ( \9631_9930 , RIdf30fe8_1934, \8884_9183 );
and \U$876 ( \9632_9931 , RIdf2ee28_1910, \8886_9185 );
or \U$877 ( \9633_9932 , \9569_9868 , \9570_9869 , \9571_9870 , \9572_9871 , \9573_9872 , \9574_9873 , \9575_9874 , \9576_9875 , \9577_9876 , \9578_9877 , \9579_9878 , \9580_9879 , \9581_9880 , \9582_9881 , \9583_9882 , \9584_9883 , \9585_9884 , \9586_9885 , \9587_9886 , \9588_9887 , \9589_9888 , \9590_9889 , \9591_9890 , \9592_9891 , \9593_9892 , \9594_9893 , \9595_9894 , \9596_9895 , \9597_9896 , \9598_9897 , \9599_9898 , \9600_9899 , \9601_9900 , \9602_9901 , \9603_9902 , \9604_9903 , \9605_9904 , \9606_9905 , \9607_9906 , \9608_9907 , \9609_9908 , \9610_9909 , \9611_9910 , \9612_9911 , \9613_9912 , \9614_9913 , \9615_9914 , \9616_9915 , \9617_9916 , \9618_9917 , \9619_9918 , \9620_9919 , \9621_9920 , \9622_9921 , \9623_9922 , \9624_9923 , \9625_9924 , \9626_9925 , \9627_9926 , \9628_9927 , \9629_9928 , \9630_9929 , \9631_9930 , \9632_9931 );
and \U$878 ( \9634_9933 , RIee2ba20_4955, \8889_9188 );
and \U$879 ( \9635_9934 , RIfc93ba8_6703, \8891_9190 );
and \U$880 ( \9636_9935 , RIfc77de0_6386, \8893_9192 );
and \U$881 ( \9637_9936 , RIee27ad8_4910, \8895_9194 );
and \U$882 ( \9638_9937 , RIfe9d668_8135, \8897_9196 );
and \U$883 ( \9639_9938 , RIfea8bd0_8236, \8899_9198 );
and \U$884 ( \9640_9939 , RIdf26458_1812, \8901_9200 );
and \U$885 ( \9641_9940 , RIfe9d7d0_8136, \8903_9202 );
and \U$886 ( \9642_9941 , RIfcb1c98_7045, \8905_9204 );
and \U$887 ( \9643_9942 , RIee26cc8_4900, \8907_9206 );
and \U$888 ( \9644_9943 , RIdf22ab0_1771, \8909_9208 );
and \U$889 ( \9645_9944 , RIfcc0068_7207, \8911_9210 );
and \U$890 ( \9646_9945 , RIdf21598_1756, \8913_9212 );
and \U$891 ( \9647_9946 , RIdf1f6a8_1734, \8915_9214 );
and \U$892 ( \9648_9947 , RIdf1aef0_1683, \8917_9216 );
and \U$893 ( \9649_9948 , RIfe9d938_8137, \8919_9218 );
and \U$894 ( \9650_9949 , RIdf16cd8_1636, \8921_9220 );
and \U$895 ( \9651_9950 , RIdf13fd8_1604, \8923_9222 );
and \U$896 ( \9652_9951 , RIdf112d8_1572, \8925_9224 );
and \U$897 ( \9653_9952 , RIdf0e5d8_1540, \8927_9226 );
and \U$898 ( \9654_9953 , RIdf0b8d8_1508, \8929_9228 );
and \U$899 ( \9655_9954 , RIdf08bd8_1476, \8931_9230 );
and \U$900 ( \9656_9955 , RIdf05ed8_1444, \8933_9232 );
and \U$901 ( \9657_9956 , RIdf031d8_1412, \8935_9234 );
and \U$902 ( \9658_9957 , RIdefd7d8_1348, \8937_9236 );
and \U$903 ( \9659_9958 , RIdefaad8_1316, \8939_9238 );
and \U$904 ( \9660_9959 , RIdef7dd8_1284, \8941_9240 );
and \U$905 ( \9661_9960 , RIdef50d8_1252, \8943_9242 );
and \U$906 ( \9662_9961 , RIdef23d8_1220, \8945_9244 );
and \U$907 ( \9663_9962 , RIdeef6d8_1188, \8947_9246 );
and \U$908 ( \9664_9963 , RIdeec9d8_1156, \8949_9248 );
and \U$909 ( \9665_9964 , RIdee9cd8_1124, \8951_9250 );
and \U$910 ( \9666_9965 , RIfc942b0_6708, \8953_9252 );
and \U$911 ( \9667_9966 , RIfcde6f8_7553, \8955_9254 );
and \U$912 ( \9668_9967 , RIfcd1138_7401, \8957_9256 );
and \U$913 ( \9669_9968 , RIfcde860_7554, \8959_9258 );
and \U$914 ( \9670_9969 , RIdee4878_1064, \8961_9260 );
and \U$915 ( \9671_9970 , RIdee2af0_1043, \8963_9262 );
and \U$916 ( \9672_9971 , RIdee0a98_1020, \8965_9264 );
and \U$917 ( \9673_9972 , RIdede8d8_996, \8967_9266 );
and \U$918 ( \9674_9973 , RIfc5c9f0_6076, \8969_9268 );
and \U$919 ( \9675_9974 , RIee22240_4847, \8971_9270 );
and \U$920 ( \9676_9975 , RIfcc8768_7303, \8973_9272 );
and \U$921 ( \9677_9976 , RIee21160_4835, \8975_9274 );
and \U$922 ( \9678_9977 , RIded95e0_937, \8977_9276 );
and \U$923 ( \9679_9978 , RIded7150_911, \8979_9278 );
and \U$924 ( \9680_9979 , RIded5260_889, \8981_9280 );
and \U$925 ( \9681_9980 , RIfea76b8_8221, \8983_9282 );
and \U$926 ( \9682_9981 , RIded0508_834, \8985_9284 );
and \U$927 ( \9683_9982 , RIdecd808_802, \8987_9286 );
and \U$928 ( \9684_9983 , RIdecab08_770, \8989_9288 );
and \U$929 ( \9685_9984 , RIdec7e08_738, \8991_9290 );
and \U$930 ( \9686_9985 , RIdeb4308_514, \8993_9292 );
and \U$931 ( \9687_9986 , RIde96290_322, \8995_9294 );
and \U$932 ( \9688_9987 , RIe16df10_2628, \8997_9296 );
and \U$933 ( \9689_9988 , RIe159d08_2399, \8999_9298 );
and \U$934 ( \9690_9989 , RIe143508_2143, \9001_9300 );
and \U$935 ( \9691_9990 , RIdf37f00_2013, \9003_9302 );
and \U$936 ( \9692_9991 , RIdf2c560_1881, \9005_9304 );
and \U$937 ( \9693_9992 , RIdf1cde0_1705, \9007_9306 );
and \U$938 ( \9694_9993 , RIdf004d8_1380, \9009_9308 );
and \U$939 ( \9695_9994 , RIdee6fd8_1092, \9011_9310 );
and \U$940 ( \9696_9995 , RIdedbd40_965, \9013_9312 );
and \U$941 ( \9697_9996 , RIde7c1d8_195, \9015_9314 );
or \U$942 ( \9698_9997 , \9634_9933 , \9635_9934 , \9636_9935 , \9637_9936 , \9638_9937 , \9639_9938 , \9640_9939 , \9641_9940 , \9642_9941 , \9643_9942 , \9644_9943 , \9645_9944 , \9646_9945 , \9647_9946 , \9648_9947 , \9649_9948 , \9650_9949 , \9651_9950 , \9652_9951 , \9653_9952 , \9654_9953 , \9655_9954 , \9656_9955 , \9657_9956 , \9658_9957 , \9659_9958 , \9660_9959 , \9661_9960 , \9662_9961 , \9663_9962 , \9664_9963 , \9665_9964 , \9666_9965 , \9667_9966 , \9668_9967 , \9669_9968 , \9670_9969 , \9671_9970 , \9672_9971 , \9673_9972 , \9674_9973 , \9675_9974 , \9676_9975 , \9677_9976 , \9678_9977 , \9679_9978 , \9680_9979 , \9681_9980 , \9682_9981 , \9683_9982 , \9684_9983 , \9685_9984 , \9686_9985 , \9687_9986 , \9688_9987 , \9689_9988 , \9690_9989 , \9691_9990 , \9692_9991 , \9693_9992 , \9694_9993 , \9695_9994 , \9696_9995 , \9697_9996 );
or \U$943 ( \9699_9998 , \9633_9932 , \9698_9997 );
_DC \g31cb/U$1 ( \9700 , \9699_9998 , \9024_9323 );
buf \U$944 ( \9701_10000 , \9700 );
and \U$945 ( \9702_10001 , RIe19d3a0_3166, \9034_9333 );
and \U$946 ( \9703_10002 , RIe19a6a0_3134, \9036_9335 );
and \U$947 ( \9704_10003 , RIfcb2c10_7056, \9038_9337 );
and \U$948 ( \9705_10004 , RIe1979a0_3102, \9040_9339 );
and \U$949 ( \9706_10005 , RIfc923c0_6686, \9042_9341 );
and \U$950 ( \9707_10006 , RIe194ca0_3070, \9044_9343 );
and \U$951 ( \9708_10007 , RIe191fa0_3038, \9046_9345 );
and \U$952 ( \9709_10008 , RIe18f2a0_3006, \9048_9347 );
and \U$953 ( \9710_10009 , RIe1898a0_2942, \9050_9349 );
and \U$954 ( \9711_10010 , RIe186ba0_2910, \9052_9351 );
and \U$955 ( \9712_10011 , RIfc422a8_5775, \9054_9353 );
and \U$956 ( \9713_10012 , RIe183ea0_2878, \9056_9355 );
and \U$957 ( \9714_10013 , RIfcbecb8_7193, \9058_9357 );
and \U$958 ( \9715_10014 , RIe1811a0_2846, \9060_9359 );
and \U$959 ( \9716_10015 , RIe17e4a0_2814, \9062_9361 );
and \U$960 ( \9717_10016 , RIe17b7a0_2782, \9064_9363 );
and \U$961 ( \9718_10017 , RIf142250_5212, \9066_9365 );
and \U$962 ( \9719_10018 , RIf140bd0_5196, \9068_9367 );
and \U$963 ( \9720_10019 , RIfec43f8_8353, \9070_9369 );
and \U$964 ( \9721_10020 , RIe175968_2715, \9072_9371 );
and \U$965 ( \9722_10021 , RIfc79b68_6407, \9074_9373 );
and \U$966 ( \9723_10022 , RIf13efb0_5176, \9076_9375 );
and \U$967 ( \9724_10023 , RIfc92528_6687, \9078_9377 );
and \U$968 ( \9725_10024 , RIfcb2aa8_7055, \9080_9379 );
and \U$969 ( \9726_10025 , RIfcd8320_7482, \9082_9381 );
and \U$970 ( \9727_10026 , RIfcea200_7686, \9084_9383 );
and \U$971 ( \9728_10027 , RIfc79898_6405, \9086_9385 );
and \U$972 ( \9729_10028 , RIe1734d8_2689, \9088_9387 );
and \U$973 ( \9730_10029 , RIfcd7948_7475, \9090_9389 );
and \U$974 ( \9731_10030 , RIfcd7678_7473, \9092_9391 );
and \U$975 ( \9732_10031 , RIf16e170_5712, \9094_9393 );
and \U$976 ( \9733_10032 , RIfc927f8_6689, \9096_9395 );
and \U$977 ( \9734_10033 , RIfc92960_6690, \9098_9397 );
and \U$978 ( \9735_10034 , RIe2236f8_4693, \9100_9399 );
and \U$979 ( \9736_10035 , RIfc795c8_6403, \9102_9401 );
and \U$980 ( \9737_10036 , RIe2209f8_4661, \9104_9403 );
and \U$981 ( \9738_10037 , RIf16ad68_5675, \9106_9405 );
and \U$982 ( \9739_10038 , RIe21dcf8_4629, \9108_9407 );
and \U$983 ( \9740_10039 , RIe2182f8_4565, \9110_9409 );
and \U$984 ( \9741_10040 , RIe2155f8_4533, \9112_9411 );
and \U$985 ( \9742_10041 , RIfe9d398_8133, \9114_9413 );
and \U$986 ( \9743_10042 , RIe2128f8_4501, \9116_9415 );
and \U$987 ( \9744_10043 , RIfcdb9f8_7521, \9118_9417 );
and \U$988 ( \9745_10044 , RIe20fbf8_4469, \9120_9419 );
and \U$989 ( \9746_10045 , RIfc41d08_5771, \9122_9421 );
and \U$990 ( \9747_10046 , RIe20cef8_4437, \9124_9423 );
and \U$991 ( \9748_10047 , RIe20a1f8_4405, \9126_9425 );
and \U$992 ( \9749_10048 , RIe2074f8_4373, \9128_9427 );
and \U$993 ( \9750_10049 , RIfcd7510_7472, \9130_9429 );
and \U$994 ( \9751_10050 , RIf166010_5620, \9132_9431 );
and \U$995 ( \9752_10051 , RIfe9d230_8132, \9134_9433 );
and \U$996 ( \9753_10052 , RIe2008b0_4296, \9136_9435 );
and \U$997 ( \9754_10053 , RIf165098_5609, \9138_9437 );
and \U$998 ( \9755_10054 , RIfc41ba0_5770, \9140_9439 );
and \U$999 ( \9756_10055 , RIfc41a38_5769, \9142_9441 );
and \U$1000 ( \9757_10056 , RIfc92c30_6692, \9144_9443 );
and \U$1001 ( \9758_10057 , RIfc418d0_5768, \9146_9445 );
and \U$1002 ( \9759_10058 , RIfc79190_6400, \9148_9447 );
and \U$1003 ( \9760_10059 , RIe1fcad0_4252, \9150_9449 );
and \U$1004 ( \9761_10060 , RIfec4560_8354, \9152_9451 );
and \U$1005 ( \9762_10061 , RIfc79028_6399, \9154_9453 );
and \U$1006 ( \9763_10062 , RIfcbf258_7197, \9156_9455 );
and \U$1007 ( \9764_10063 , RIfcc1df0_7228, \9158_9457 );
and \U$1008 ( \9765_10064 , RIfcd81b8_7481, \9160_9459 );
or \U$1009 ( \9766_10065 , \9702_10001 , \9703_10002 , \9704_10003 , \9705_10004 , \9706_10005 , \9707_10006 , \9708_10007 , \9709_10008 , \9710_10009 , \9711_10010 , \9712_10011 , \9713_10012 , \9714_10013 , \9715_10014 , \9716_10015 , \9717_10016 , \9718_10017 , \9719_10018 , \9720_10019 , \9721_10020 , \9722_10021 , \9723_10022 , \9724_10023 , \9725_10024 , \9726_10025 , \9727_10026 , \9728_10027 , \9729_10028 , \9730_10029 , \9731_10030 , \9732_10031 , \9733_10032 , \9734_10033 , \9735_10034 , \9736_10035 , \9737_10036 , \9738_10037 , \9739_10038 , \9740_10039 , \9741_10040 , \9742_10041 , \9743_10042 , \9744_10043 , \9745_10044 , \9746_10045 , \9747_10046 , \9748_10047 , \9749_10048 , \9750_10049 , \9751_10050 , \9752_10051 , \9753_10052 , \9754_10053 , \9755_10054 , \9756_10055 , \9757_10056 , \9758_10057 , \9759_10058 , \9760_10059 , \9761_10060 , \9762_10061 , \9763_10062 , \9764_10063 , \9765_10064 );
and \U$1010 ( \9767_10066 , RIfc92d98_6693, \9163_9462 );
and \U$1011 ( \9768_10067 , RIfc5b4d8_6061, \9165_9464 );
and \U$1012 ( \9769_10068 , RIfcd77e0_7474, \9167_9466 );
and \U$1013 ( \9770_10069 , RIe1fa0a0_4222, \9169_9468 );
and \U$1014 ( \9771_10070 , RIf156188_5439, \9171_9470 );
and \U$1015 ( \9772_10071 , RIfe9d500_8134, \9173_9472 );
and \U$1016 ( \9773_10072 , RIf1546d0_5420, \9175_9474 );
and \U$1017 ( \9774_10073 , RIe1f5348_4167, \9177_9476 );
and \U$1018 ( \9775_10074 , RIfec4830_8356, \9179_9478 );
and \U$1019 ( \9776_10075 , RIfec46c8_8355, \9181_9480 );
and \U$1020 ( \9777_10076 , RIf1508f0_5376, \9183_9482 );
and \U$1021 ( \9778_10077 , RIe1f3020_4142, \9185_9484 );
and \U$1022 ( \9779_10078 , RIfce3180_7606, \9187_9486 );
and \U$1023 ( \9780_10079 , RIfce8fb8_7673, \9189_9488 );
and \U$1024 ( \9781_10080 , RIfcbf690_7200, \9191_9490 );
and \U$1025 ( \9782_10081 , RIe1edd28_4083, \9193_9492 );
and \U$1026 ( \9783_10082 , RIe1eb460_4054, \9195_9494 );
and \U$1027 ( \9784_10083 , RIe1e8760_4022, \9197_9496 );
and \U$1028 ( \9785_10084 , RIe1e5a60_3990, \9199_9498 );
and \U$1029 ( \9786_10085 , RIe1e2d60_3958, \9201_9500 );
and \U$1030 ( \9787_10086 , RIe1e0060_3926, \9203_9502 );
and \U$1031 ( \9788_10087 , RIe1dd360_3894, \9205_9504 );
and \U$1032 ( \9789_10088 , RIe1da660_3862, \9207_9506 );
and \U$1033 ( \9790_10089 , RIe1d7960_3830, \9209_9508 );
and \U$1034 ( \9791_10090 , RIe1d1f60_3766, \9211_9510 );
and \U$1035 ( \9792_10091 , RIe1cf260_3734, \9213_9512 );
and \U$1036 ( \9793_10092 , RIe1cc560_3702, \9215_9514 );
and \U$1037 ( \9794_10093 , RIe1c9860_3670, \9217_9516 );
and \U$1038 ( \9795_10094 , RIe1c6b60_3638, \9219_9518 );
and \U$1039 ( \9796_10095 , RIe1c3e60_3606, \9221_9520 );
and \U$1040 ( \9797_10096 , RIe1c1160_3574, \9223_9522 );
and \U$1041 ( \9798_10097 , RIe1be460_3542, \9225_9524 );
and \U$1042 ( \9799_10098 , RIfe9d0c8_8131, \9227_9526 );
and \U$1043 ( \9800_10099 , RIfe9cc90_8128, \9229_9528 );
and \U$1044 ( \9801_10100 , RIe1b9168_3483, \9231_9530 );
and \U$1045 ( \9802_10101 , RIe1b7110_3460, \9233_9532 );
and \U$1046 ( \9803_10102 , RIf14a3b0_5304, \9235_9534 );
and \U$1047 ( \9804_10103 , RIfe9cb28_8127, \9237_9536 );
and \U$1048 ( \9805_10104 , RIfe9cf60_8130, \9239_9538 );
and \U$1049 ( \9806_10105 , RIfe9c9c0_8126, \9241_9540 );
and \U$1050 ( \9807_10106 , RIfce2208_7595, \9243_9542 );
and \U$1051 ( \9808_10107 , RIfce9558_7677, \9245_9544 );
and \U$1052 ( \9809_10108 , RIfe9c858_8125, \9247_9546 );
and \U$1053 ( \9810_10109 , RIfe9cdf8_8129, \9249_9548 );
and \U$1054 ( \9811_10110 , RIf147110_5268, \9251_9550 );
and \U$1055 ( \9812_10111 , RIf146468_5259, \9253_9552 );
and \U$1056 ( \9813_10112 , RIe1ac2b0_3336, \9255_9554 );
and \U$1057 ( \9814_10113 , RIe1aaac8_3319, \9257_9556 );
and \U$1058 ( \9815_10114 , RIe1a87a0_3294, \9259_9558 );
and \U$1059 ( \9816_10115 , RIe1a5aa0_3262, \9261_9560 );
and \U$1060 ( \9817_10116 , RIe1a2da0_3230, \9263_9562 );
and \U$1061 ( \9818_10117 , RIe1a00a0_3198, \9265_9564 );
and \U$1062 ( \9819_10118 , RIe18c5a0_2974, \9267_9566 );
and \U$1063 ( \9820_10119 , RIe178aa0_2750, \9269_9568 );
and \U$1064 ( \9821_10120 , RIe2263f8_4725, \9271_9570 );
and \U$1065 ( \9822_10121 , RIe21aff8_4597, \9273_9572 );
and \U$1066 ( \9823_10122 , RIe2047f8_4341, \9275_9574 );
and \U$1067 ( \9824_10123 , RIe1fe858_4273, \9277_9576 );
and \U$1068 ( \9825_10124 , RIe1f7c10_4196, \9279_9578 );
and \U$1069 ( \9826_10125 , RIe1f0758_4113, \9281_9580 );
and \U$1070 ( \9827_10126 , RIe1d4c60_3798, \9283_9582 );
and \U$1071 ( \9828_10127 , RIe1bb760_3510, \9285_9584 );
and \U$1072 ( \9829_10128 , RIe1ae5d8_3361, \9287_9586 );
and \U$1073 ( \9830_10129 , RIe170c10_2660, \9289_9588 );
or \U$1074 ( \9831_10130 , \9767_10066 , \9768_10067 , \9769_10068 , \9770_10069 , \9771_10070 , \9772_10071 , \9773_10072 , \9774_10073 , \9775_10074 , \9776_10075 , \9777_10076 , \9778_10077 , \9779_10078 , \9780_10079 , \9781_10080 , \9782_10081 , \9783_10082 , \9784_10083 , \9785_10084 , \9786_10085 , \9787_10086 , \9788_10087 , \9789_10088 , \9790_10089 , \9791_10090 , \9792_10091 , \9793_10092 , \9794_10093 , \9795_10094 , \9796_10095 , \9797_10096 , \9798_10097 , \9799_10098 , \9800_10099 , \9801_10100 , \9802_10101 , \9803_10102 , \9804_10103 , \9805_10104 , \9806_10105 , \9807_10106 , \9808_10107 , \9809_10108 , \9810_10109 , \9811_10110 , \9812_10111 , \9813_10112 , \9814_10113 , \9815_10114 , \9816_10115 , \9817_10116 , \9818_10117 , \9819_10118 , \9820_10119 , \9821_10120 , \9822_10121 , \9823_10122 , \9824_10123 , \9825_10124 , \9826_10125 , \9827_10126 , \9828_10127 , \9829_10128 , \9830_10129 );
or \U$1075 ( \9832_10131 , \9766_10065 , \9831_10130 );
_DC \g42f8/U$1 ( \9833 , \9832_10131 , \9298_9597 );
buf \U$1076 ( \9834_10133 , \9833 );
and \U$1077 ( \9835_10134 , \9701_10000 , \9834_10133 );
and \U$1078 ( \9836_10135 , RIdec4190_695, \8760_9059 );
and \U$1079 ( \9837_10136 , RIdec1490_663, \8762_9061 );
and \U$1080 ( \9838_10137 , RIfceaa70_7692, \8764_9063 );
and \U$1081 ( \9839_10138 , RIdebe790_631, \8766_9065 );
and \U$1082 ( \9840_10139 , RIfc954f8_6721, \8768_9067 );
and \U$1083 ( \9841_10140 , RIdebba90_599, \8770_9069 );
and \U$1084 ( \9842_10141 , RIdeb8d90_567, \8772_9071 );
and \U$1085 ( \9843_10142 , RIdeb6090_535, \8774_9073 );
and \U$1086 ( \9844_10143 , RIfcebb50_7704, \8776_9075 );
and \U$1087 ( \9845_10144 , RIdeb0690_471, \8778_9077 );
and \U$1088 ( \9846_10145 , RIee1e190_4801, \8780_9079 );
and \U$1089 ( \9847_10146 , RIdead990_439, \8782_9081 );
and \U$1090 ( \9848_10147 , RIfcdf0d0_7560, \8784_9083 );
and \U$1091 ( \9849_10148 , RIdea7978_407, \8786_9085 );
and \U$1092 ( \9850_10149 , RIdea1078_375, \8788_9087 );
and \U$1093 ( \9851_10150 , RIde9a778_343, \8790_9089 );
and \U$1094 ( \9852_10151 , RIee1c840_4783, \8792_9091 );
and \U$1095 ( \9853_10152 , RIfc957c8_6723, \8794_9093 );
and \U$1096 ( \9854_10153 , RIfcc8e70_7308, \8796_9095 );
and \U$1097 ( \9855_10154 , RIfc5e610_6096, \8798_9097 );
and \U$1098 ( \9856_10155 , RIfe9e8b0_8148, \8800_9099 );
and \U$1099 ( \9857_10156 , RIde8c1c8_273, \8802_9101 );
and \U$1100 ( \9858_10157 , RIde88028_253, \8804_9103 );
and \U$1101 ( \9859_10158 , RIde83b40_232, \8806_9105 );
and \U$1102 ( \9860_10159 , RIfcb0bb8_7033, \8808_9107 );
and \U$1103 ( \9861_10160 , RIfca4b10_6896, \8810_9109 );
and \U$1104 ( \9862_10161 , RIfc75d88_6363, \8812_9111 );
and \U$1105 ( \9863_10162 , RIfca4c78_6897, \8814_9113 );
and \U$1106 ( \9864_10163 , RIfc95390_6720, \8816_9115 );
and \U$1107 ( \9865_10164 , RIe16a9a0_2590, \8818_9117 );
and \U$1108 ( \9866_10165 , RIfcc8fd8_7309, \8820_9119 );
and \U$1109 ( \9867_10166 , RIe166e90_2548, \8822_9121 );
and \U$1110 ( \9868_10167 , RIe164190_2516, \8824_9123 );
and \U$1111 ( \9869_10168 , RIe161490_2484, \8826_9125 );
and \U$1112 ( \9870_10169 , RIfe9e748_8147, \8828_9127 );
and \U$1113 ( \9871_10170 , RIe15e790_2452, \8830_9129 );
and \U$1114 ( \9872_10171 , RIfc74f78_6353, \8832_9131 );
and \U$1115 ( \9873_10172 , RIe15ba90_2420, \8834_9133 );
and \U$1116 ( \9874_10173 , RIe156090_2356, \8836_9135 );
and \U$1117 ( \9875_10174 , RIe153390_2324, \8838_9137 );
and \U$1118 ( \9876_10175 , RIfc3ecc0_5740, \8840_9139 );
and \U$1119 ( \9877_10176 , RIe150690_2292, \8842_9141 );
and \U$1120 ( \9878_10177 , RIfce8b80_7670, \8844_9143 );
and \U$1121 ( \9879_10178 , RIe14d990_2260, \8846_9145 );
and \U$1122 ( \9880_10179 , RIfca6730_6916, \8848_9147 );
and \U$1123 ( \9881_10180 , RIe14ac90_2228, \8850_9149 );
and \U$1124 ( \9882_10181 , RIe147f90_2196, \8852_9151 );
and \U$1125 ( \9883_10182 , RIe145290_2164, \8854_9153 );
and \U$1126 ( \9884_10183 , RIfcee2b0_7732, \8856_9155 );
and \U$1127 ( \9885_10184 , RIfc5f2b8_6105, \8858_9157 );
and \U$1128 ( \9886_10185 , RIfc753b0_6356, \8860_9159 );
and \U$1129 ( \9887_10186 , RIfc74b40_6350, \8862_9161 );
and \U$1130 ( \9888_10187 , RIe140268_2107, \8864_9163 );
and \U$1131 ( \9889_10188 , RIdf3e170_2083, \8866_9165 );
and \U$1132 ( \9890_10189 , RIdf3be48_2058, \8868_9167 );
and \U$1133 ( \9891_10190 , RIdf39c88_2034, \8870_9169 );
and \U$1134 ( \9892_10191 , RIfcc1c88_7227, \8872_9171 );
and \U$1135 ( \9893_10192 , RIfcc1850_7224, \8874_9173 );
and \U$1136 ( \9894_10193 , RIfc965d8_6733, \8876_9175 );
and \U$1137 ( \9895_10194 , RIfc96038_6729, \8878_9177 );
and \U$1138 ( \9896_10195 , RIdf34828_1974, \8880_9179 );
and \U$1139 ( \9897_10196 , RIdf327d0_1951, \8882_9181 );
and \U$1140 ( \9898_10197 , RIdf301d8_1924, \8884_9183 );
and \U$1141 ( \9899_10198 , RIdf2e2e8_1902, \8886_9185 );
or \U$1142 ( \9900_10199 , \9836_10135 , \9837_10136 , \9838_10137 , \9839_10138 , \9840_10139 , \9841_10140 , \9842_10141 , \9843_10142 , \9844_10143 , \9845_10144 , \9846_10145 , \9847_10146 , \9848_10147 , \9849_10148 , \9850_10149 , \9851_10150 , \9852_10151 , \9853_10152 , \9854_10153 , \9855_10154 , \9856_10155 , \9857_10156 , \9858_10157 , \9859_10158 , \9860_10159 , \9861_10160 , \9862_10161 , \9863_10162 , \9864_10163 , \9865_10164 , \9866_10165 , \9867_10166 , \9868_10167 , \9869_10168 , \9870_10169 , \9871_10170 , \9872_10171 , \9873_10172 , \9874_10173 , \9875_10174 , \9876_10175 , \9877_10176 , \9878_10177 , \9879_10178 , \9880_10179 , \9881_10180 , \9882_10181 , \9883_10182 , \9884_10183 , \9885_10184 , \9886_10185 , \9887_10186 , \9888_10187 , \9889_10188 , \9890_10189 , \9891_10190 , \9892_10191 , \9893_10192 , \9894_10193 , \9895_10194 , \9896_10195 , \9897_10196 , \9898_10197 , \9899_10198 );
and \U$1143 ( \9901_10200 , RIfc5e778_6097, \8889_9188 );
and \U$1144 ( \9902_10201 , RIfcd0328_7391, \8891_9190 );
and \U$1145 ( \9903_10202 , RIfc757e8_6359, \8893_9192 );
and \U$1146 ( \9904_10203 , RIfcee6e8_7735, \8895_9194 );
and \U$1147 ( \9905_10204 , RIdf296f8_1848, \8897_9196 );
and \U$1148 ( \9906_10205 , RIdf273d0_1823, \8899_9198 );
and \U$1149 ( \9907_10206 , RIdf257b0_1803, \8901_9200 );
and \U$1150 ( \9908_10207 , RIdf23b90_1783, \8903_9202 );
and \U$1151 ( \9909_10208 , RIfc95d68_6727, \8905_9204 );
and \U$1152 ( \9910_10209 , RIfceda40_7726, \8907_9206 );
and \U$1153 ( \9911_10210 , RIfe9eb80_8150, \8909_9208 );
and \U$1154 ( \9912_10211 , RIfc75518_6357, \8911_9210 );
and \U$1155 ( \9913_10212 , RIfcd01c0_7390, \8913_9212 );
and \U$1156 ( \9914_10213 , RIdf1eb68_1726, \8915_9214 );
and \U$1157 ( \9915_10214 , RIfe9ece8_8151, \8917_9216 );
and \U$1158 ( \9916_10215 , RIfe9ea18_8149, \8919_9218 );
and \U$1159 ( \9917_10216 , RIdf15d60_1625, \8921_9220 );
and \U$1160 ( \9918_10217 , RIdf13060_1593, \8923_9222 );
and \U$1161 ( \9919_10218 , RIdf10360_1561, \8925_9224 );
and \U$1162 ( \9920_10219 , RIdf0d660_1529, \8927_9226 );
and \U$1163 ( \9921_10220 , RIdf0a960_1497, \8929_9228 );
and \U$1164 ( \9922_10221 , RIdf07c60_1465, \8931_9230 );
and \U$1165 ( \9923_10222 , RIdf04f60_1433, \8933_9232 );
and \U$1166 ( \9924_10223 , RIdf02260_1401, \8935_9234 );
and \U$1167 ( \9925_10224 , RIdefc860_1337, \8937_9236 );
and \U$1168 ( \9926_10225 , RIdef9b60_1305, \8939_9238 );
and \U$1169 ( \9927_10226 , RIdef6e60_1273, \8941_9240 );
and \U$1170 ( \9928_10227 , RIdef4160_1241, \8943_9242 );
and \U$1171 ( \9929_10228 , RIdef1460_1209, \8945_9244 );
and \U$1172 ( \9930_10229 , RIdeee760_1177, \8947_9246 );
and \U$1173 ( \9931_10230 , RIdeeba60_1145, \8949_9248 );
and \U$1174 ( \9932_10231 , RIdee8d60_1113, \8951_9250 );
and \U$1175 ( \9933_10232 , RIfc961a0_6730, \8953_9252 );
and \U$1176 ( \9934_10233 , RIfc96308_6731, \8955_9254 );
and \U$1177 ( \9935_10234 , RIfc5ee80_6102, \8957_9256 );
and \U$1178 ( \9936_10235 , RIfce6150_7640, \8959_9258 );
and \U$1179 ( \9937_10236 , RIdee42d8_1060, \8961_9260 );
and \U$1180 ( \9938_10237 , RIdee1e48_1034, \8963_9262 );
and \U$1181 ( \9939_10238 , RIdee00c0_1013, \8965_9264 );
and \U$1182 ( \9940_10239 , RIdeddac8_986, \8967_9266 );
and \U$1183 ( \9941_10240 , RIfc96470_6732, \8969_9268 );
and \U$1184 ( \9942_10241 , RIfc75248_6355, \8971_9270 );
and \U$1185 ( \9943_10242 , RIfc74ca8_6351, \8973_9272 );
and \U$1186 ( \9944_10243 , RIfcb0618_7029, \8975_9274 );
and \U$1187 ( \9945_10244 , RIded8938_928, \8977_9276 );
and \U$1188 ( \9946_10245 , RIded6610_903, \8979_9278 );
and \U$1189 ( \9947_10246 , RIded4450_879, \8981_9280 );
and \U$1190 ( \9948_10247 , RIded2290_855, \8983_9282 );
and \U$1191 ( \9949_10248 , RIdecf590_823, \8985_9284 );
and \U$1192 ( \9950_10249 , RIdecc890_791, \8987_9286 );
and \U$1193 ( \9951_10250 , RIdec9b90_759, \8989_9288 );
and \U$1194 ( \9952_10251 , RIdec6e90_727, \8991_9290 );
and \U$1195 ( \9953_10252 , RIdeb3390_503, \8993_9292 );
and \U$1196 ( \9954_10253 , RIde93e78_311, \8995_9294 );
and \U$1197 ( \9955_10254 , RIe16cf98_2617, \8997_9296 );
and \U$1198 ( \9956_10255 , RIe158d90_2388, \8999_9298 );
and \U$1199 ( \9957_10256 , RIe142590_2132, \9001_9300 );
and \U$1200 ( \9958_10257 , RIdf36f88_2002, \9003_9302 );
and \U$1201 ( \9959_10258 , RIdf2b5e8_1870, \9005_9304 );
and \U$1202 ( \9960_10259 , RIdf1be68_1694, \9007_9306 );
and \U$1203 ( \9961_10260 , RIdeff560_1369, \9009_9308 );
and \U$1204 ( \9962_10261 , RIdee6060_1081, \9011_9310 );
and \U$1205 ( \9963_10262 , RIdedadc8_954, \9013_9312 );
and \U$1206 ( \9964_10263 , RIde79dc0_184, \9015_9314 );
or \U$1207 ( \9965_10264 , \9901_10200 , \9902_10201 , \9903_10202 , \9904_10203 , \9905_10204 , \9906_10205 , \9907_10206 , \9908_10207 , \9909_10208 , \9910_10209 , \9911_10210 , \9912_10211 , \9913_10212 , \9914_10213 , \9915_10214 , \9916_10215 , \9917_10216 , \9918_10217 , \9919_10218 , \9920_10219 , \9921_10220 , \9922_10221 , \9923_10222 , \9924_10223 , \9925_10224 , \9926_10225 , \9927_10226 , \9928_10227 , \9929_10228 , \9930_10229 , \9931_10230 , \9932_10231 , \9933_10232 , \9934_10233 , \9935_10234 , \9936_10235 , \9937_10236 , \9938_10237 , \9939_10238 , \9940_10239 , \9941_10240 , \9942_10241 , \9943_10242 , \9944_10243 , \9945_10244 , \9946_10245 , \9947_10246 , \9948_10247 , \9949_10248 , \9950_10249 , \9951_10250 , \9952_10251 , \9953_10252 , \9954_10253 , \9955_10254 , \9956_10255 , \9957_10256 , \9958_10257 , \9959_10258 , \9960_10259 , \9961_10260 , \9962_10261 , \9963_10262 , \9964_10263 );
or \U$1208 ( \9966_10265 , \9900_10199 , \9965_10264 );
_DC \g3250/U$1 ( \9967 , \9966_10265 , \9024_9323 );
buf \U$1209 ( \9968_10267 , \9967 );
and \U$1210 ( \9969_10268 , RIe19c428_3155, \9034_9333 );
and \U$1211 ( \9970_10269 , RIe199728_3123, \9036_9335 );
and \U$1212 ( \9971_10270 , RIfe9e310_8144, \9038_9337 );
and \U$1213 ( \9972_10271 , RIe196a28_3091, \9040_9339 );
and \U$1214 ( \9973_10272 , RIfcc04a0_7210, \9042_9341 );
and \U$1215 ( \9974_10273 , RIe193d28_3059, \9044_9343 );
and \U$1216 ( \9975_10274 , RIe191028_3027, \9046_9345 );
and \U$1217 ( \9976_10275 , RIe18e328_2995, \9048_9347 );
and \U$1218 ( \9977_10276 , RIe188928_2931, \9050_9349 );
and \U$1219 ( \9978_10277 , RIe185c28_2899, \9052_9351 );
and \U$1220 ( \9979_10278 , RIfce1830_7588, \9054_9353 );
and \U$1221 ( \9980_10279 , RIe182f28_2867, \9056_9355 );
and \U$1222 ( \9981_10280 , RIfe9e478_8145, \9058_9357 );
and \U$1223 ( \9982_10281 , RIe180228_2835, \9060_9359 );
and \U$1224 ( \9983_10282 , RIe17d528_2803, \9062_9361 );
and \U$1225 ( \9984_10283 , RIe17a828_2771, \9064_9363 );
and \U$1226 ( \9985_10284 , RIf141878_5205, \9066_9365 );
and \U$1227 ( \9986_10285 , RIfcb12c0_7038, \9068_9367 );
and \U$1228 ( \9987_10286 , RIfc94418_6709, \9070_9369 );
and \U$1229 ( \9988_10287 , RIe174f90_2708, \9072_9371 );
and \U$1230 ( \9989_10288 , RIfc77408_6379, \9074_9373 );
and \U$1231 ( \9990_10289 , RIf13ea10_5172, \9076_9375 );
and \U$1232 ( \9991_10290 , RIfcdc100_7526, \9078_9377 );
and \U$1233 ( \9992_10291 , RIfc94580_6710, \9080_9379 );
and \U$1234 ( \9993_10292 , RIfc946e8_6711, \9082_9381 );
and \U$1235 ( \9994_10293 , RIfced338_7721, \9084_9383 );
and \U$1236 ( \9995_10294 , RIfce5fe8_7639, \9086_9385 );
and \U$1237 ( \9996_10295 , RIe172998_2681, \9088_9387 );
and \U$1238 ( \9997_10296 , RIfcdc268_7527, \9090_9389 );
and \U$1239 ( \9998_10297 , RIfcddff0_7548, \9092_9391 );
and \U$1240 ( \9999_10298 , RIfcc0608_7211, \9094_9393 );
and \U$1241 ( \10000_10299 , RIfce7230_7652, \9096_9395 );
and \U$1242 ( \10001_10300 , RIfc40340_5756, \9098_9397 );
and \U$1243 ( \10002_10301 , RIe222780_4682, \9100_9399 );
and \U$1244 ( \10003_10302 , RIfcdd618_7541, \9102_9401 );
and \U$1245 ( \10004_10303 , RIe21fa80_4650, \9104_9403 );
and \U$1246 ( \10005_10304 , RIfcd0b98_7397, \9106_9405 );
and \U$1247 ( \10006_10305 , RIe21cd80_4618, \9108_9407 );
and \U$1248 ( \10007_10306 , RIe217380_4554, \9110_9409 );
and \U$1249 ( \10008_10307 , RIe214680_4522, \9112_9411 );
and \U$1250 ( \10009_10308 , RIfec4998_8357, \9114_9413 );
and \U$1251 ( \10010_10309 , RIe211980_4490, \9116_9415 );
and \U$1252 ( \10011_10310 , RIf168608_5647, \9118_9417 );
and \U$1253 ( \10012_10311 , RIe20ec80_4458, \9120_9419 );
and \U$1254 ( \10013_10312 , RIfcc0770_7212, \9122_9421 );
and \U$1255 ( \10014_10313 , RIe20bf80_4426, \9124_9423 );
and \U$1256 ( \10015_10314 , RIe209280_4394, \9126_9425 );
and \U$1257 ( \10016_10315 , RIe206580_4362, \9128_9427 );
and \U$1258 ( \10017_10316 , RIfce2370_7596, \9130_9429 );
and \U$1259 ( \10018_10317 , RIfcee580_7734, \9132_9431 );
and \U$1260 ( \10019_10318 , RIfec4c68_8359, \9134_9433 );
and \U$1261 ( \10020_10319 , RIfec4b00_8358, \9136_9435 );
and \U$1262 ( \10021_10320 , RIfc949b8_6713, \9138_9437 );
and \U$1263 ( \10022_10321 , RIfcebcb8_7705, \9140_9439 );
and \U$1264 ( \10023_10322 , RIf162938_5581, \9142_9441 );
and \U$1265 ( \10024_10323 , RIf1612b8_5565, \9144_9443 );
and \U$1266 ( \10025_10324 , RIfccd088_7355, \9146_9445 );
and \U$1267 ( \10026_10325 , RIfcc08d8_7213, \9148_9447 );
and \U$1268 ( \10027_10326 , RIfe9e040_8142, \9150_9449 );
and \U$1269 ( \10028_10327 , RIfe9e1a8_8143, \9152_9451 );
and \U$1270 ( \10029_10328 , RIfcead40_7694, \9154_9453 );
and \U$1271 ( \10030_10329 , RIf15ad78_5493, \9156_9455 );
and \U$1272 ( \10031_10330 , RIfc94c88_6715, \9158_9457 );
and \U$1273 ( \10032_10331 , RIfccc3e0_7346, \9160_9459 );
or \U$1274 ( \10033_10332 , \9969_10268 , \9970_10269 , \9971_10270 , \9972_10271 , \9973_10272 , \9974_10273 , \9975_10274 , \9976_10275 , \9977_10276 , \9978_10277 , \9979_10278 , \9980_10279 , \9981_10280 , \9982_10281 , \9983_10282 , \9984_10283 , \9985_10284 , \9986_10285 , \9987_10286 , \9988_10287 , \9989_10288 , \9990_10289 , \9991_10290 , \9992_10291 , \9993_10292 , \9994_10293 , \9995_10294 , \9996_10295 , \9997_10296 , \9998_10297 , \9999_10298 , \10000_10299 , \10001_10300 , \10002_10301 , \10003_10302 , \10004_10303 , \10005_10304 , \10006_10305 , \10007_10306 , \10008_10307 , \10009_10308 , \10010_10309 , \10011_10310 , \10012_10311 , \10013_10312 , \10014_10313 , \10015_10314 , \10016_10315 , \10017_10316 , \10018_10317 , \10019_10318 , \10020_10319 , \10021_10320 , \10022_10321 , \10023_10322 , \10024_10323 , \10025_10324 , \10026_10325 , \10027_10326 , \10028_10327 , \10029_10328 , \10030_10329 , \10031_10330 , \10032_10331 );
and \U$1275 ( \10034_10333 , RIfc765f8_6369, \9163_9462 );
and \U$1276 ( \10035_10334 , RIfc94df0_6716, \9165_9464 );
and \U$1277 ( \10036_10335 , RIfcc0a40_7214, \9167_9466 );
and \U$1278 ( \10037_10336 , RIe1f9998_4217, \9169_9468 );
and \U$1279 ( \10038_10337 , RIfcc8d08_7307, \9171_9470 );
and \U$1280 ( \10039_10338 , RIfce8748_7667, \9173_9472 );
and \U$1281 ( \10040_10339 , RIfceb2e0_7698, \9175_9474 );
and \U$1282 ( \10041_10340 , RIe1f4970_4160, \9177_9476 );
and \U$1283 ( \10042_10341 , RIf152510_5396, \9179_9478 );
and \U$1284 ( \10043_10342 , RIf1512c8_5383, \9181_9480 );
and \U$1285 ( \10044_10343 , RIfcb0ff0_7036, \9183_9482 );
and \U$1286 ( \10045_10344 , RIe1f24e0_4134, \9185_9484 );
and \U$1287 ( \10046_10345 , RIfc761c0_6366, \9187_9486 );
and \U$1288 ( \10047_10346 , RIfc950c0_6718, \9189_9488 );
and \U$1289 ( \10048_10347 , RIfcc0e78_7217, \9191_9490 );
and \U$1290 ( \10049_10348 , RIe1ed1e8_4075, \9193_9492 );
and \U$1291 ( \10050_10349 , RIe1ea4e8_4043, \9195_9494 );
and \U$1292 ( \10051_10350 , RIe1e77e8_4011, \9197_9496 );
and \U$1293 ( \10052_10351 , RIe1e4ae8_3979, \9199_9498 );
and \U$1294 ( \10053_10352 , RIe1e1de8_3947, \9201_9500 );
and \U$1295 ( \10054_10353 , RIe1df0e8_3915, \9203_9502 );
and \U$1296 ( \10055_10354 , RIe1dc3e8_3883, \9205_9504 );
and \U$1297 ( \10056_10355 , RIe1d96e8_3851, \9207_9506 );
and \U$1298 ( \10057_10356 , RIe1d69e8_3819, \9209_9508 );
and \U$1299 ( \10058_10357 , RIe1d0fe8_3755, \9211_9510 );
and \U$1300 ( \10059_10358 , RIe1ce2e8_3723, \9213_9512 );
and \U$1301 ( \10060_10359 , RIe1cb5e8_3691, \9215_9514 );
and \U$1302 ( \10061_10360 , RIe1c88e8_3659, \9217_9516 );
and \U$1303 ( \10062_10361 , RIe1c5be8_3627, \9219_9518 );
and \U$1304 ( \10063_10362 , RIe1c2ee8_3595, \9221_9520 );
and \U$1305 ( \10064_10363 , RIe1c01e8_3563, \9223_9522 );
and \U$1306 ( \10065_10364 , RIe1bd4e8_3531, \9225_9524 );
and \U$1307 ( \10066_10365 , RIf14bfd0_5324, \9227_9526 );
and \U$1308 ( \10067_10366 , RIf14ac20_5310, \9229_9528 );
and \U$1309 ( \10068_10367 , RIfe9ded8_8141, \9231_9530 );
and \U$1310 ( \10069_10368 , RIe1b65d0_3452, \9233_9532 );
and \U$1311 ( \10070_10369 , RIfcecd98_7717, \9235_9534 );
and \U$1312 ( \10071_10370 , RIfc76490_6368, \9237_9536 );
and \U$1313 ( \10072_10371 , RIe1b4c80_3434, \9239_9538 );
and \U$1314 ( \10073_10372 , RIe1b38d0_3420, \9241_9540 );
and \U$1315 ( \10074_10373 , RIfcc0fe0_7218, \9243_9542 );
and \U$1316 ( \10075_10374 , RIfceaea8_7695, \9245_9544 );
and \U$1317 ( \10076_10375 , RIe1b1f80_3402, \9247_9546 );
and \U$1318 ( \10077_10376 , RIe1b0360_3382, \9249_9548 );
and \U$1319 ( \10078_10377 , RIfcd0760_7394, \9251_9550 );
and \U$1320 ( \10079_10378 , RIf145ec8_5255, \9253_9552 );
and \U$1321 ( \10080_10379 , RIfe9e5e0_8146, \9255_9554 );
and \U$1322 ( \10081_10380 , RIfe9dd70_8140, \9257_9556 );
and \U$1323 ( \10082_10381 , RIe1a7828_3283, \9259_9558 );
and \U$1324 ( \10083_10382 , RIe1a4b28_3251, \9261_9560 );
and \U$1325 ( \10084_10383 , RIe1a1e28_3219, \9263_9562 );
and \U$1326 ( \10085_10384 , RIe19f128_3187, \9265_9564 );
and \U$1327 ( \10086_10385 , RIe18b628_2963, \9267_9566 );
and \U$1328 ( \10087_10386 , RIe177b28_2739, \9269_9568 );
and \U$1329 ( \10088_10387 , RIe225480_4714, \9271_9570 );
and \U$1330 ( \10089_10388 , RIe21a080_4586, \9273_9572 );
and \U$1331 ( \10090_10389 , RIe203880_4330, \9275_9574 );
and \U$1332 ( \10091_10390 , RIe1fd8e0_4262, \9277_9576 );
and \U$1333 ( \10092_10391 , RIe1f6c98_4185, \9279_9578 );
and \U$1334 ( \10093_10392 , RIe1ef7e0_4102, \9281_9580 );
and \U$1335 ( \10094_10393 , RIe1d3ce8_3787, \9283_9582 );
and \U$1336 ( \10095_10394 , RIe1ba7e8_3499, \9285_9584 );
and \U$1337 ( \10096_10395 , RIe1ad660_3350, \9287_9586 );
and \U$1338 ( \10097_10396 , RIe16fc98_2649, \9289_9588 );
or \U$1339 ( \10098_10397 , \10034_10333 , \10035_10334 , \10036_10335 , \10037_10336 , \10038_10337 , \10039_10338 , \10040_10339 , \10041_10340 , \10042_10341 , \10043_10342 , \10044_10343 , \10045_10344 , \10046_10345 , \10047_10346 , \10048_10347 , \10049_10348 , \10050_10349 , \10051_10350 , \10052_10351 , \10053_10352 , \10054_10353 , \10055_10354 , \10056_10355 , \10057_10356 , \10058_10357 , \10059_10358 , \10060_10359 , \10061_10360 , \10062_10361 , \10063_10362 , \10064_10363 , \10065_10364 , \10066_10365 , \10067_10366 , \10068_10367 , \10069_10368 , \10070_10369 , \10071_10370 , \10072_10371 , \10073_10372 , \10074_10373 , \10075_10374 , \10076_10375 , \10077_10376 , \10078_10377 , \10079_10378 , \10080_10379 , \10081_10380 , \10082_10381 , \10083_10382 , \10084_10383 , \10085_10384 , \10086_10385 , \10087_10386 , \10088_10387 , \10089_10388 , \10090_10389 , \10091_10390 , \10092_10391 , \10093_10392 , \10094_10393 , \10095_10394 , \10096_10395 , \10097_10396 );
or \U$1340 ( \10099_10398 , \10033_10332 , \10098_10397 );
_DC \g437d/U$1 ( \10100 , \10099_10398 , \9298_9597 );
buf \U$1341 ( \10101_10400 , \10100 );
and \U$1342 ( \10102_10401 , \9968_10267 , \10101_10400 );
and \U$1343 ( \10103_10402 , \9834_10133 , \10102_10401 );
and \U$1344 ( \10104_10403 , \9701_10000 , \10102_10401 );
or \U$1345 ( \10105_10404 , \9835_10134 , \10103_10402 , \10104_10403 );
and \U$1346 ( \10106_10405 , \9567_9866 , \10105_10404 );
and \U$1347 ( \10107_10406 , \9434_9733 , \10105_10404 );
or \U$1348 ( \10108_10407 , \9568_9867 , \10106_10405 , \10107_10406 );
xor \U$1349 ( \10109_10408 , \9301_9600 , \10108_10407 );
buf g444e_GF_PartitionCandidate( \10110_10409_nG444e , \10109_10408 );
xor \U$1350 ( \10111_10410 , \9434_9733 , \9567_9866 );
xor \U$1351 ( \10112_10411 , \10111_10410 , \10105_10404 );
buf g4451_GF_PartitionCandidate( \10113_10412_nG4451 , \10112_10411 );
xor \U$1352 ( \10114_10413 , \9701_10000 , \9834_10133 );
xor \U$1353 ( \10115_10414 , \10114_10413 , \10102_10401 );
buf g4454_GF_PartitionCandidate( \10116_10415_nG4454 , \10115_10414 );
nand \U$1354 ( \10117_10416 , \10113_10412_nG4451 , \10116_10415_nG4454 );
and \U$1355 ( \10118_10417 , \10110_10409_nG444e , \10117_10416 );
xor \U$1356 ( \10119_10418 , \10113_10412_nG4451 , \10116_10415_nG4454 );
and \U$1362 ( \10120_10422 , RIdec4190_695, \9034_9333 );
and \U$1363 ( \10121_10423 , RIdec1490_663, \9036_9335 );
and \U$1364 ( \10122_10424 , RIfceaa70_7692, \9038_9337 );
and \U$1365 ( \10123_10425 , RIdebe790_631, \9040_9339 );
and \U$1366 ( \10124_10426 , RIfc954f8_6721, \9042_9341 );
and \U$1367 ( \10125_10427 , RIdebba90_599, \9044_9343 );
and \U$1368 ( \10126_10428 , RIdeb8d90_567, \9046_9345 );
and \U$1369 ( \10127_10429 , RIdeb6090_535, \9048_9347 );
and \U$1370 ( \10128_10430 , RIfcebb50_7704, \9050_9349 );
and \U$1371 ( \10129_10431 , RIdeb0690_471, \9052_9351 );
and \U$1372 ( \10130_10432 , RIee1e190_4801, \9054_9353 );
and \U$1373 ( \10131_10433 , RIdead990_439, \9056_9355 );
and \U$1374 ( \10132_10434 , RIfcdf0d0_7560, \9058_9357 );
and \U$1375 ( \10133_10435 , RIdea7978_407, \9060_9359 );
and \U$1376 ( \10134_10436 , RIdea1078_375, \9062_9361 );
and \U$1377 ( \10135_10437 , RIde9a778_343, \9064_9363 );
and \U$1378 ( \10136_10438 , RIee1c840_4783, \9066_9365 );
and \U$1379 ( \10137_10439 , RIfc957c8_6723, \9068_9367 );
and \U$1380 ( \10138_10440 , RIfcc8e70_7308, \9070_9369 );
and \U$1381 ( \10139_10441 , RIfc5e610_6096, \9072_9371 );
and \U$1382 ( \10140_10442 , RIfe9e8b0_8148, \9074_9373 );
and \U$1383 ( \10141_10443 , RIde8c1c8_273, \9076_9375 );
and \U$1384 ( \10142_10444 , RIde88028_253, \9078_9377 );
and \U$1385 ( \10143_10445 , RIde83b40_232, \9080_9379 );
and \U$1386 ( \10144_10446 , RIfcb0bb8_7033, \9082_9381 );
and \U$1387 ( \10145_10447 , RIfca4b10_6896, \9084_9383 );
and \U$1388 ( \10146_10448 , RIfc75d88_6363, \9086_9385 );
and \U$1389 ( \10147_10449 , RIfca4c78_6897, \9088_9387 );
and \U$1390 ( \10148_10450 , RIfc95390_6720, \9090_9389 );
and \U$1391 ( \10149_10451 , RIe16a9a0_2590, \9092_9391 );
and \U$1392 ( \10150_10452 , RIfcc8fd8_7309, \9094_9393 );
and \U$1393 ( \10151_10453 , RIe166e90_2548, \9096_9395 );
and \U$1394 ( \10152_10454 , RIe164190_2516, \9098_9397 );
and \U$1395 ( \10153_10455 , RIe161490_2484, \9100_9399 );
and \U$1396 ( \10154_10456 , RIfe9e748_8147, \9102_9401 );
and \U$1397 ( \10155_10457 , RIe15e790_2452, \9104_9403 );
and \U$1398 ( \10156_10458 , RIfc74f78_6353, \9106_9405 );
and \U$1399 ( \10157_10459 , RIe15ba90_2420, \9108_9407 );
and \U$1400 ( \10158_10460 , RIe156090_2356, \9110_9409 );
and \U$1401 ( \10159_10461 , RIe153390_2324, \9112_9411 );
and \U$1402 ( \10160_10462 , RIfc3ecc0_5740, \9114_9413 );
and \U$1403 ( \10161_10463 , RIe150690_2292, \9116_9415 );
and \U$1404 ( \10162_10464 , RIfce8b80_7670, \9118_9417 );
and \U$1405 ( \10163_10465 , RIe14d990_2260, \9120_9419 );
and \U$1406 ( \10164_10466 , RIfca6730_6916, \9122_9421 );
and \U$1407 ( \10165_10467 , RIe14ac90_2228, \9124_9423 );
and \U$1408 ( \10166_10468 , RIe147f90_2196, \9126_9425 );
and \U$1409 ( \10167_10469 , RIe145290_2164, \9128_9427 );
and \U$1410 ( \10168_10470 , RIfcee2b0_7732, \9130_9429 );
and \U$1411 ( \10169_10471 , RIfc5f2b8_6105, \9132_9431 );
and \U$1412 ( \10170_10472 , RIfc753b0_6356, \9134_9433 );
and \U$1413 ( \10171_10473 , RIfc74b40_6350, \9136_9435 );
and \U$1414 ( \10172_10474 , RIe140268_2107, \9138_9437 );
and \U$1415 ( \10173_10475 , RIdf3e170_2083, \9140_9439 );
and \U$1416 ( \10174_10476 , RIdf3be48_2058, \9142_9441 );
and \U$1417 ( \10175_10477 , RIdf39c88_2034, \9144_9443 );
and \U$1418 ( \10176_10478 , RIfcc1c88_7227, \9146_9445 );
and \U$1419 ( \10177_10479 , RIfcc1850_7224, \9148_9447 );
and \U$1420 ( \10178_10480 , RIfc965d8_6733, \9150_9449 );
and \U$1421 ( \10179_10481 , RIfc96038_6729, \9152_9451 );
and \U$1422 ( \10180_10482 , RIdf34828_1974, \9154_9453 );
and \U$1423 ( \10181_10483 , RIdf327d0_1951, \9156_9455 );
and \U$1424 ( \10182_10484 , RIdf301d8_1924, \9158_9457 );
and \U$1425 ( \10183_10485 , RIdf2e2e8_1902, \9160_9459 );
or \U$1426 ( \10184_10486 , \10120_10422 , \10121_10423 , \10122_10424 , \10123_10425 , \10124_10426 , \10125_10427 , \10126_10428 , \10127_10429 , \10128_10430 , \10129_10431 , \10130_10432 , \10131_10433 , \10132_10434 , \10133_10435 , \10134_10436 , \10135_10437 , \10136_10438 , \10137_10439 , \10138_10440 , \10139_10441 , \10140_10442 , \10141_10443 , \10142_10444 , \10143_10445 , \10144_10446 , \10145_10447 , \10146_10448 , \10147_10449 , \10148_10450 , \10149_10451 , \10150_10452 , \10151_10453 , \10152_10454 , \10153_10455 , \10154_10456 , \10155_10457 , \10156_10458 , \10157_10459 , \10158_10460 , \10159_10461 , \10160_10462 , \10161_10463 , \10162_10464 , \10163_10465 , \10164_10466 , \10165_10467 , \10166_10468 , \10167_10469 , \10168_10470 , \10169_10471 , \10170_10472 , \10171_10473 , \10172_10474 , \10173_10475 , \10174_10476 , \10175_10477 , \10176_10478 , \10177_10479 , \10178_10480 , \10179_10481 , \10180_10482 , \10181_10483 , \10182_10484 , \10183_10485 );
and \U$1427 ( \10185_10487 , RIfc5e778_6097, \9163_9462 );
and \U$1428 ( \10186_10488 , RIfcd0328_7391, \9165_9464 );
and \U$1429 ( \10187_10489 , RIfc757e8_6359, \9167_9466 );
and \U$1430 ( \10188_10490 , RIfcee6e8_7735, \9169_9468 );
and \U$1431 ( \10189_10491 , RIdf296f8_1848, \9171_9470 );
and \U$1432 ( \10190_10492 , RIdf273d0_1823, \9173_9472 );
and \U$1433 ( \10191_10493 , RIdf257b0_1803, \9175_9474 );
and \U$1434 ( \10192_10494 , RIdf23b90_1783, \9177_9476 );
and \U$1435 ( \10193_10495 , RIfc95d68_6727, \9179_9478 );
and \U$1436 ( \10194_10496 , RIfceda40_7726, \9181_9480 );
and \U$1437 ( \10195_10497 , RIfe9eb80_8150, \9183_9482 );
and \U$1438 ( \10196_10498 , RIfc75518_6357, \9185_9484 );
and \U$1439 ( \10197_10499 , RIfcd01c0_7390, \9187_9486 );
and \U$1440 ( \10198_10500 , RIdf1eb68_1726, \9189_9488 );
and \U$1441 ( \10199_10501 , RIfe9ece8_8151, \9191_9490 );
and \U$1442 ( \10200_10502 , RIfe9ea18_8149, \9193_9492 );
and \U$1443 ( \10201_10503 , RIdf15d60_1625, \9195_9494 );
and \U$1444 ( \10202_10504 , RIdf13060_1593, \9197_9496 );
and \U$1445 ( \10203_10505 , RIdf10360_1561, \9199_9498 );
and \U$1446 ( \10204_10506 , RIdf0d660_1529, \9201_9500 );
and \U$1447 ( \10205_10507 , RIdf0a960_1497, \9203_9502 );
and \U$1448 ( \10206_10508 , RIdf07c60_1465, \9205_9504 );
and \U$1449 ( \10207_10509 , RIdf04f60_1433, \9207_9506 );
and \U$1450 ( \10208_10510 , RIdf02260_1401, \9209_9508 );
and \U$1451 ( \10209_10511 , RIdefc860_1337, \9211_9510 );
and \U$1452 ( \10210_10512 , RIdef9b60_1305, \9213_9512 );
and \U$1453 ( \10211_10513 , RIdef6e60_1273, \9215_9514 );
and \U$1454 ( \10212_10514 , RIdef4160_1241, \9217_9516 );
and \U$1455 ( \10213_10515 , RIdef1460_1209, \9219_9518 );
and \U$1456 ( \10214_10516 , RIdeee760_1177, \9221_9520 );
and \U$1457 ( \10215_10517 , RIdeeba60_1145, \9223_9522 );
and \U$1458 ( \10216_10518 , RIdee8d60_1113, \9225_9524 );
and \U$1459 ( \10217_10519 , RIfc961a0_6730, \9227_9526 );
and \U$1460 ( \10218_10520 , RIfc96308_6731, \9229_9528 );
and \U$1461 ( \10219_10521 , RIfc5ee80_6102, \9231_9530 );
and \U$1462 ( \10220_10522 , RIfce6150_7640, \9233_9532 );
and \U$1463 ( \10221_10523 , RIdee42d8_1060, \9235_9534 );
and \U$1464 ( \10222_10524 , RIdee1e48_1034, \9237_9536 );
and \U$1465 ( \10223_10525 , RIdee00c0_1013, \9239_9538 );
and \U$1466 ( \10224_10526 , RIdeddac8_986, \9241_9540 );
and \U$1467 ( \10225_10527 , RIfc96470_6732, \9243_9542 );
and \U$1468 ( \10226_10528 , RIfc75248_6355, \9245_9544 );
and \U$1469 ( \10227_10529 , RIfc74ca8_6351, \9247_9546 );
and \U$1470 ( \10228_10530 , RIfcb0618_7029, \9249_9548 );
and \U$1471 ( \10229_10531 , RIded8938_928, \9251_9550 );
and \U$1472 ( \10230_10532 , RIded6610_903, \9253_9552 );
and \U$1473 ( \10231_10533 , RIded4450_879, \9255_9554 );
and \U$1474 ( \10232_10534 , RIded2290_855, \9257_9556 );
and \U$1475 ( \10233_10535 , RIdecf590_823, \9259_9558 );
and \U$1476 ( \10234_10536 , RIdecc890_791, \9261_9560 );
and \U$1477 ( \10235_10537 , RIdec9b90_759, \9263_9562 );
and \U$1478 ( \10236_10538 , RIdec6e90_727, \9265_9564 );
and \U$1479 ( \10237_10539 , RIdeb3390_503, \9267_9566 );
and \U$1480 ( \10238_10540 , RIde93e78_311, \9269_9568 );
and \U$1481 ( \10239_10541 , RIe16cf98_2617, \9271_9570 );
and \U$1482 ( \10240_10542 , RIe158d90_2388, \9273_9572 );
and \U$1483 ( \10241_10543 , RIe142590_2132, \9275_9574 );
and \U$1484 ( \10242_10544 , RIdf36f88_2002, \9277_9576 );
and \U$1485 ( \10243_10545 , RIdf2b5e8_1870, \9279_9578 );
and \U$1486 ( \10244_10546 , RIdf1be68_1694, \9281_9580 );
and \U$1487 ( \10245_10547 , RIdeff560_1369, \9283_9582 );
and \U$1488 ( \10246_10548 , RIdee6060_1081, \9285_9584 );
and \U$1489 ( \10247_10549 , RIdedadc8_954, \9287_9586 );
and \U$1490 ( \10248_10550 , RIde79dc0_184, \9289_9588 );
or \U$1491 ( \10249_10551 , \10185_10487 , \10186_10488 , \10187_10489 , \10188_10490 , \10189_10491 , \10190_10492 , \10191_10493 , \10192_10494 , \10193_10495 , \10194_10496 , \10195_10497 , \10196_10498 , \10197_10499 , \10198_10500 , \10199_10501 , \10200_10502 , \10201_10503 , \10202_10504 , \10203_10505 , \10204_10506 , \10205_10507 , \10206_10508 , \10207_10509 , \10208_10510 , \10209_10511 , \10210_10512 , \10211_10513 , \10212_10514 , \10213_10515 , \10214_10516 , \10215_10517 , \10216_10518 , \10217_10519 , \10218_10520 , \10219_10521 , \10220_10522 , \10221_10523 , \10222_10524 , \10223_10525 , \10224_10526 , \10225_10527 , \10226_10528 , \10227_10529 , \10228_10530 , \10229_10531 , \10230_10532 , \10231_10533 , \10232_10534 , \10233_10535 , \10234_10536 , \10235_10537 , \10236_10538 , \10237_10539 , \10238_10540 , \10239_10541 , \10240_10542 , \10241_10543 , \10242_10544 , \10243_10545 , \10244_10546 , \10245_10547 , \10246_10548 , \10247_10549 , \10248_10550 );
or \U$1492 ( \10250_10552 , \10184_10486 , \10249_10551 );
_DC \g6577/U$1 ( \10251 , \10250_10552 , \9298_9597 );
and \U$1493 ( \10252_10554 , RIe19c428_3155, \8760_9059 );
and \U$1494 ( \10253_10555 , RIe199728_3123, \8762_9061 );
and \U$1495 ( \10254_10556 , RIfe9e310_8144, \8764_9063 );
and \U$1496 ( \10255_10557 , RIe196a28_3091, \8766_9065 );
and \U$1497 ( \10256_10558 , RIfcc04a0_7210, \8768_9067 );
and \U$1498 ( \10257_10559 , RIe193d28_3059, \8770_9069 );
and \U$1499 ( \10258_10560 , RIe191028_3027, \8772_9071 );
and \U$1500 ( \10259_10561 , RIe18e328_2995, \8774_9073 );
and \U$1501 ( \10260_10562 , RIe188928_2931, \8776_9075 );
and \U$1502 ( \10261_10563 , RIe185c28_2899, \8778_9077 );
and \U$1503 ( \10262_10564 , RIfce1830_7588, \8780_9079 );
and \U$1504 ( \10263_10565 , RIe182f28_2867, \8782_9081 );
and \U$1505 ( \10264_10566 , RIfe9e478_8145, \8784_9083 );
and \U$1506 ( \10265_10567 , RIe180228_2835, \8786_9085 );
and \U$1507 ( \10266_10568 , RIe17d528_2803, \8788_9087 );
and \U$1508 ( \10267_10569 , RIe17a828_2771, \8790_9089 );
and \U$1509 ( \10268_10570 , RIf141878_5205, \8792_9091 );
and \U$1510 ( \10269_10571 , RIfcb12c0_7038, \8794_9093 );
and \U$1511 ( \10270_10572 , RIfc94418_6709, \8796_9095 );
and \U$1512 ( \10271_10573 , RIe174f90_2708, \8798_9097 );
and \U$1513 ( \10272_10574 , RIfc77408_6379, \8800_9099 );
and \U$1514 ( \10273_10575 , RIf13ea10_5172, \8802_9101 );
and \U$1515 ( \10274_10576 , RIfcdc100_7526, \8804_9103 );
and \U$1516 ( \10275_10577 , RIfc94580_6710, \8806_9105 );
and \U$1517 ( \10276_10578 , RIfc946e8_6711, \8808_9107 );
and \U$1518 ( \10277_10579 , RIfced338_7721, \8810_9109 );
and \U$1519 ( \10278_10580 , RIfce5fe8_7639, \8812_9111 );
and \U$1520 ( \10279_10581 , RIe172998_2681, \8814_9113 );
and \U$1521 ( \10280_10582 , RIfcdc268_7527, \8816_9115 );
and \U$1522 ( \10281_10583 , RIfcddff0_7548, \8818_9117 );
and \U$1523 ( \10282_10584 , RIfcc0608_7211, \8820_9119 );
and \U$1524 ( \10283_10585 , RIfce7230_7652, \8822_9121 );
and \U$1525 ( \10284_10586 , RIfc40340_5756, \8824_9123 );
and \U$1526 ( \10285_10587 , RIe222780_4682, \8826_9125 );
and \U$1527 ( \10286_10588 , RIfcdd618_7541, \8828_9127 );
and \U$1528 ( \10287_10589 , RIe21fa80_4650, \8830_9129 );
and \U$1529 ( \10288_10590 , RIfcd0b98_7397, \8832_9131 );
and \U$1530 ( \10289_10591 , RIe21cd80_4618, \8834_9133 );
and \U$1531 ( \10290_10592 , RIe217380_4554, \8836_9135 );
and \U$1532 ( \10291_10593 , RIe214680_4522, \8838_9137 );
and \U$1533 ( \10292_10594 , RIfec4998_8357, \8840_9139 );
and \U$1534 ( \10293_10595 , RIe211980_4490, \8842_9141 );
and \U$1535 ( \10294_10596 , RIf168608_5647, \8844_9143 );
and \U$1536 ( \10295_10597 , RIe20ec80_4458, \8846_9145 );
and \U$1537 ( \10296_10598 , RIfcc0770_7212, \8848_9147 );
and \U$1538 ( \10297_10599 , RIe20bf80_4426, \8850_9149 );
and \U$1539 ( \10298_10600 , RIe209280_4394, \8852_9151 );
and \U$1540 ( \10299_10601 , RIe206580_4362, \8854_9153 );
and \U$1541 ( \10300_10602 , RIfce2370_7596, \8856_9155 );
and \U$1542 ( \10301_10603 , RIfcee580_7734, \8858_9157 );
and \U$1543 ( \10302_10604 , RIfec4c68_8359, \8860_9159 );
and \U$1544 ( \10303_10605 , RIfec4b00_8358, \8862_9161 );
and \U$1545 ( \10304_10606 , RIfc949b8_6713, \8864_9163 );
and \U$1546 ( \10305_10607 , RIfcebcb8_7705, \8866_9165 );
and \U$1547 ( \10306_10608 , RIf162938_5581, \8868_9167 );
and \U$1548 ( \10307_10609 , RIf1612b8_5565, \8870_9169 );
and \U$1549 ( \10308_10610 , RIfccd088_7355, \8872_9171 );
and \U$1550 ( \10309_10611 , RIfcc08d8_7213, \8874_9173 );
and \U$1551 ( \10310_10612 , RIfe9e040_8142, \8876_9175 );
and \U$1552 ( \10311_10613 , RIfe9e1a8_8143, \8878_9177 );
and \U$1553 ( \10312_10614 , RIfcead40_7694, \8880_9179 );
and \U$1554 ( \10313_10615 , RIf15ad78_5493, \8882_9181 );
and \U$1555 ( \10314_10616 , RIfc94c88_6715, \8884_9183 );
and \U$1556 ( \10315_10617 , RIfccc3e0_7346, \8886_9185 );
or \U$1557 ( \10316_10618 , \10252_10554 , \10253_10555 , \10254_10556 , \10255_10557 , \10256_10558 , \10257_10559 , \10258_10560 , \10259_10561 , \10260_10562 , \10261_10563 , \10262_10564 , \10263_10565 , \10264_10566 , \10265_10567 , \10266_10568 , \10267_10569 , \10268_10570 , \10269_10571 , \10270_10572 , \10271_10573 , \10272_10574 , \10273_10575 , \10274_10576 , \10275_10577 , \10276_10578 , \10277_10579 , \10278_10580 , \10279_10581 , \10280_10582 , \10281_10583 , \10282_10584 , \10283_10585 , \10284_10586 , \10285_10587 , \10286_10588 , \10287_10589 , \10288_10590 , \10289_10591 , \10290_10592 , \10291_10593 , \10292_10594 , \10293_10595 , \10294_10596 , \10295_10597 , \10296_10598 , \10297_10599 , \10298_10600 , \10299_10601 , \10300_10602 , \10301_10603 , \10302_10604 , \10303_10605 , \10304_10606 , \10305_10607 , \10306_10608 , \10307_10609 , \10308_10610 , \10309_10611 , \10310_10612 , \10311_10613 , \10312_10614 , \10313_10615 , \10314_10616 , \10315_10617 );
and \U$1558 ( \10317_10619 , RIfc765f8_6369, \8889_9188 );
and \U$1559 ( \10318_10620 , RIfc94df0_6716, \8891_9190 );
and \U$1560 ( \10319_10621 , RIfcc0a40_7214, \8893_9192 );
and \U$1561 ( \10320_10622 , RIe1f9998_4217, \8895_9194 );
and \U$1562 ( \10321_10623 , RIfcc8d08_7307, \8897_9196 );
and \U$1563 ( \10322_10624 , RIfce8748_7667, \8899_9198 );
and \U$1564 ( \10323_10625 , RIfceb2e0_7698, \8901_9200 );
and \U$1565 ( \10324_10626 , RIe1f4970_4160, \8903_9202 );
and \U$1566 ( \10325_10627 , RIf152510_5396, \8905_9204 );
and \U$1567 ( \10326_10628 , RIf1512c8_5383, \8907_9206 );
and \U$1568 ( \10327_10629 , RIfcb0ff0_7036, \8909_9208 );
and \U$1569 ( \10328_10630 , RIe1f24e0_4134, \8911_9210 );
and \U$1570 ( \10329_10631 , RIfc761c0_6366, \8913_9212 );
and \U$1571 ( \10330_10632 , RIfc950c0_6718, \8915_9214 );
and \U$1572 ( \10331_10633 , RIfcc0e78_7217, \8917_9216 );
and \U$1573 ( \10332_10634 , RIe1ed1e8_4075, \8919_9218 );
and \U$1574 ( \10333_10635 , RIe1ea4e8_4043, \8921_9220 );
and \U$1575 ( \10334_10636 , RIe1e77e8_4011, \8923_9222 );
and \U$1576 ( \10335_10637 , RIe1e4ae8_3979, \8925_9224 );
and \U$1577 ( \10336_10638 , RIe1e1de8_3947, \8927_9226 );
and \U$1578 ( \10337_10639 , RIe1df0e8_3915, \8929_9228 );
and \U$1579 ( \10338_10640 , RIe1dc3e8_3883, \8931_9230 );
and \U$1580 ( \10339_10641 , RIe1d96e8_3851, \8933_9232 );
and \U$1581 ( \10340_10642 , RIe1d69e8_3819, \8935_9234 );
and \U$1582 ( \10341_10643 , RIe1d0fe8_3755, \8937_9236 );
and \U$1583 ( \10342_10644 , RIe1ce2e8_3723, \8939_9238 );
and \U$1584 ( \10343_10645 , RIe1cb5e8_3691, \8941_9240 );
and \U$1585 ( \10344_10646 , RIe1c88e8_3659, \8943_9242 );
and \U$1586 ( \10345_10647 , RIe1c5be8_3627, \8945_9244 );
and \U$1587 ( \10346_10648 , RIe1c2ee8_3595, \8947_9246 );
and \U$1588 ( \10347_10649 , RIe1c01e8_3563, \8949_9248 );
and \U$1589 ( \10348_10650 , RIe1bd4e8_3531, \8951_9250 );
and \U$1590 ( \10349_10651 , RIf14bfd0_5324, \8953_9252 );
and \U$1591 ( \10350_10652 , RIf14ac20_5310, \8955_9254 );
and \U$1592 ( \10351_10653 , RIfe9ded8_8141, \8957_9256 );
and \U$1593 ( \10352_10654 , RIe1b65d0_3452, \8959_9258 );
and \U$1594 ( \10353_10655 , RIfcecd98_7717, \8961_9260 );
and \U$1595 ( \10354_10656 , RIfc76490_6368, \8963_9262 );
and \U$1596 ( \10355_10657 , RIe1b4c80_3434, \8965_9264 );
and \U$1597 ( \10356_10658 , RIe1b38d0_3420, \8967_9266 );
and \U$1598 ( \10357_10659 , RIfcc0fe0_7218, \8969_9268 );
and \U$1599 ( \10358_10660 , RIfceaea8_7695, \8971_9270 );
and \U$1600 ( \10359_10661 , RIe1b1f80_3402, \8973_9272 );
and \U$1601 ( \10360_10662 , RIe1b0360_3382, \8975_9274 );
and \U$1602 ( \10361_10663 , RIfcd0760_7394, \8977_9276 );
and \U$1603 ( \10362_10664 , RIf145ec8_5255, \8979_9278 );
and \U$1604 ( \10363_10665 , RIfe9e5e0_8146, \8981_9280 );
and \U$1605 ( \10364_10666 , RIfe9dd70_8140, \8983_9282 );
and \U$1606 ( \10365_10667 , RIe1a7828_3283, \8985_9284 );
and \U$1607 ( \10366_10668 , RIe1a4b28_3251, \8987_9286 );
and \U$1608 ( \10367_10669 , RIe1a1e28_3219, \8989_9288 );
and \U$1609 ( \10368_10670 , RIe19f128_3187, \8991_9290 );
and \U$1610 ( \10369_10671 , RIe18b628_2963, \8993_9292 );
and \U$1611 ( \10370_10672 , RIe177b28_2739, \8995_9294 );
and \U$1612 ( \10371_10673 , RIe225480_4714, \8997_9296 );
and \U$1613 ( \10372_10674 , RIe21a080_4586, \8999_9298 );
and \U$1614 ( \10373_10675 , RIe203880_4330, \9001_9300 );
and \U$1615 ( \10374_10676 , RIe1fd8e0_4262, \9003_9302 );
and \U$1616 ( \10375_10677 , RIe1f6c98_4185, \9005_9304 );
and \U$1617 ( \10376_10678 , RIe1ef7e0_4102, \9007_9306 );
and \U$1618 ( \10377_10679 , RIe1d3ce8_3787, \9009_9308 );
and \U$1619 ( \10378_10680 , RIe1ba7e8_3499, \9011_9310 );
and \U$1620 ( \10379_10681 , RIe1ad660_3350, \9013_9312 );
and \U$1621 ( \10380_10682 , RIe16fc98_2649, \9015_9314 );
or \U$1622 ( \10381_10683 , \10317_10619 , \10318_10620 , \10319_10621 , \10320_10622 , \10321_10623 , \10322_10624 , \10323_10625 , \10324_10626 , \10325_10627 , \10326_10628 , \10327_10629 , \10328_10630 , \10329_10631 , \10330_10632 , \10331_10633 , \10332_10634 , \10333_10635 , \10334_10636 , \10335_10637 , \10336_10638 , \10337_10639 , \10338_10640 , \10339_10641 , \10340_10642 , \10341_10643 , \10342_10644 , \10343_10645 , \10344_10646 , \10345_10647 , \10346_10648 , \10347_10649 , \10348_10650 , \10349_10651 , \10350_10652 , \10351_10653 , \10352_10654 , \10353_10655 , \10354_10656 , \10355_10657 , \10356_10658 , \10357_10659 , \10358_10660 , \10359_10661 , \10360_10662 , \10361_10663 , \10362_10664 , \10363_10665 , \10364_10666 , \10365_10667 , \10366_10668 , \10367_10669 , \10368_10670 , \10369_10671 , \10370_10672 , \10371_10673 , \10372_10674 , \10373_10675 , \10374_10676 , \10375_10677 , \10376_10678 , \10377_10679 , \10378_10680 , \10379_10681 , \10380_10682 );
or \U$1623 ( \10382_10684 , \10316_10618 , \10381_10683 );
_DC \g6578/U$1 ( \10383 , \10382_10684 , \9024_9323 );
and g6579_GF_PartitionCandidate( \10384_10686_nG6579 , \10251 , \10383 );
buf \U$1624 ( \10385_10687 , \10384_10686_nG6579 );
_DC \g44da/U$1 ( \10386 , \10250_10552 , \9298_9597 );
_DC \g455e/U$1 ( \10387 , \10382_10684 , \9024_9323 );
xor g455f_GF_PartitionCandidate( \10388_10690_nG455f , \10386 , \10387 );
buf \U$1625 ( \10389_10691 , \10388_10690_nG455f );
and \U$1626 ( \10390_10692 , \10385_10687 , \10389_10691 );
buf \U$1627 ( \10391_10693 , \10390_10692 );
buf g9c0e_GF_PartitionCandidate( \10392_10694_nG9c0e , \10391_10693 );
and \U$1628 ( \10393_10695 , \10119_10418 , \10392_10694_nG9c0e );
or \U$1629 ( \10394_10696 , 1'b0 , \10393_10695 );
xor \U$1630 ( \10395_10697 , \10118_10417 , \10394_10696 );
xor \U$1631 ( \10396_10698 , \10118_10417 , \10395_10697 );
buf \U$1632 ( \10397_10699 , \10396_10698 );
buf \U$1633 ( \10398_10700 , \10397_10699 );
and \U$1637 ( \10399_10703 , \10116_10415_nG4454 , 1'b1 );
xor \U$1634 ( \10400_10701 , \9968_10267 , \10101_10400 );
buf g4456_GF_PartitionCandidate( \10401_10702_nG4456 , \10400_10701 );
xor \U$1638 ( \10402_10704 , \10401_10702_nG4456 , 1'b0 );
and \U$1643 ( \10403_10708 , \10402_10704 , \10392_10694_nG9c0e );
or \U$1644 ( \10404_10709 , 1'b0 , \10403_10708 );
xor \U$1645 ( \10405_10710 , \10399_10703 , \10404_10709 );
and \U$1646 ( \10406_10711 , \10399_10703 , \10405_10710 );
buf \U$1647 ( \10407_10712 , \10406_10711 );
buf \U$1649 ( \10408_10713 , \10407_10712 );
not \U$1639 ( \10409_10705 , \10402_10704 );
xor \U$1640 ( \10410_10706 , \10116_10415_nG4454 , \10401_10702_nG4456 );
and \U$1641 ( \10411_10707 , \10409_10705 , \10410_10706 );
and \U$1650 ( \10412_10714 , \10411_10707 , \10392_10694_nG9c0e );
and \U$1651 ( \10413_10715 , RIdec5108_706, \9034_9333 );
and \U$1652 ( \10414_10716 , RIdec2408_674, \9036_9335 );
and \U$1653 ( \10415_10717 , RIfc93608_6699, \9038_9337 );
and \U$1654 ( \10416_10718 , RIdebf708_642, \9040_9339 );
and \U$1655 ( \10417_10719 , RIfc934a0_6698, \9042_9341 );
and \U$1656 ( \10418_10720 , RIdebca08_610, \9044_9343 );
and \U$1657 ( \10419_10721 , RIdeb9d08_578, \9046_9345 );
and \U$1658 ( \10420_10722 , RIdeb7008_546, \9048_9347 );
and \U$1659 ( \10421_10723 , RIfcdf7d8_7565, \9050_9349 );
and \U$1660 ( \10422_10724 , RIdeb1608_482, \9052_9351 );
and \U$1661 ( \10423_10725 , RIfc78218_6389, \9054_9353 );
and \U$1662 ( \10424_10726 , RIdeae908_450, \9056_9355 );
and \U$1663 ( \10425_10727 , RIfcc8498_7301, \9058_9357 );
and \U$1664 ( \10426_10728 , RIdea9d90_418, \9060_9359 );
and \U$1665 ( \10427_10729 , RIdea3490_386, \9062_9361 );
and \U$1666 ( \10428_10730 , RIde9cb90_354, \9064_9363 );
and \U$1667 ( \10429_10731 , RIee1cc78_4786, \9066_9365 );
and \U$1668 ( \10430_10732 , RIee1bb98_4774, \9068_9367 );
and \U$1669 ( \10431_10733 , RIee1b328_4768, \9070_9369 );
and \U$1670 ( \10432_10734 , RIee1aab8_4762, \9072_9371 );
and \U$1671 ( \10433_10735 , RIde909f8_295, \9074_9373 );
and \U$1672 ( \10434_10736 , RIde8d578_279, \9076_9375 );
and \U$1673 ( \10435_10737 , RIfea8ea0_8238, \9078_9377 );
and \U$1674 ( \10436_10738 , RIde85238_239, \9080_9379 );
and \U$1675 ( \10437_10739 , RIde813e0_220, \9082_9381 );
and \U$1676 ( \10438_10740 , RIfc938d8_6701, \9084_9383 );
and \U$1677 ( \10439_10741 , RIfce5e80_7638, \9086_9385 );
and \U$1678 ( \10440_10742 , RIfcbfd98_7205, \9088_9387 );
and \U$1679 ( \10441_10743 , RIfce8ce8_7671, \9090_9389 );
and \U$1680 ( \10442_10744 , RIe16b4e0_2598, \9092_9391 );
and \U$1681 ( \10443_10745 , RIfea8d38_8237, \9094_9393 );
and \U$1682 ( \10444_10746 , RIfea9f80_8250, \9096_9395 );
and \U$1683 ( \10445_10747 , RIe165108_2527, \9098_9397 );
and \U$1684 ( \10446_10748 , RIe162408_2495, \9100_9399 );
and \U$1685 ( \10447_10749 , RIfc779a8_6383, \9102_9401 );
and \U$1686 ( \10448_10750 , RIe15f708_2463, \9104_9403 );
and \U$1687 ( \10449_10751 , RIfe9dc08_8139, \9106_9405 );
and \U$1688 ( \10450_10752 , RIe15ca08_2431, \9108_9407 );
and \U$1689 ( \10451_10753 , RIe157008_2367, \9110_9409 );
and \U$1690 ( \10452_10754 , RIe154308_2335, \9112_9411 );
and \U$1691 ( \10453_10755 , RIfea7550_8220, \9114_9413 );
and \U$1692 ( \10454_10756 , RIe151608_2303, \9116_9415 );
and \U$1693 ( \10455_10757 , RIfcd6160_7458, \9118_9417 );
and \U$1694 ( \10456_10758 , RIe14e908_2271, \9120_9419 );
and \U$1695 ( \10457_10759 , RIfcd1408_7403, \9122_9421 );
and \U$1696 ( \10458_10760 , RIe14bc08_2239, \9124_9423 );
and \U$1697 ( \10459_10761 , RIe148f08_2207, \9126_9425 );
and \U$1698 ( \10460_10762 , RIe146208_2175, \9128_9427 );
and \U$1699 ( \10461_10763 , RIfceb718_7701, \9130_9429 );
and \U$1700 ( \10462_10764 , RIfcb19c8_7043, \9132_9431 );
and \U$1701 ( \10463_10765 , RIfc93e78_6705, \9134_9433 );
and \U$1702 ( \10464_10766 , RIfce7938_7657, \9136_9435 );
and \U$1703 ( \10465_10767 , RIe140da8_2115, \9138_9437 );
and \U$1704 ( \10466_10768 , RIdf3ecb0_2091, \9140_9439 );
and \U$1705 ( \10467_10769 , RIdf3c988_2066, \9142_9441 );
and \U$1706 ( \10468_10770 , RIfe9daa0_8138, \9144_9443 );
and \U$1707 ( \10469_10771 , RIfce8478_7665, \9146_9445 );
and \U$1708 ( \10470_10772 , RIfcdbf98_7525, \9148_9447 );
and \U$1709 ( \10471_10773 , RIfc776d8_6381, \9150_9449 );
and \U$1710 ( \10472_10774 , RIfc93fe0_6706, \9152_9451 );
and \U$1711 ( \10473_10775 , RIdf354d0_1983, \9154_9453 );
and \U$1712 ( \10474_10776 , RIdf33040_1957, \9156_9455 );
and \U$1713 ( \10475_10777 , RIdf30fe8_1934, \9158_9457 );
and \U$1714 ( \10476_10778 , RIdf2ee28_1910, \9160_9459 );
or \U$1715 ( \10477_10779 , \10413_10715 , \10414_10716 , \10415_10717 , \10416_10718 , \10417_10719 , \10418_10720 , \10419_10721 , \10420_10722 , \10421_10723 , \10422_10724 , \10423_10725 , \10424_10726 , \10425_10727 , \10426_10728 , \10427_10729 , \10428_10730 , \10429_10731 , \10430_10732 , \10431_10733 , \10432_10734 , \10433_10735 , \10434_10736 , \10435_10737 , \10436_10738 , \10437_10739 , \10438_10740 , \10439_10741 , \10440_10742 , \10441_10743 , \10442_10744 , \10443_10745 , \10444_10746 , \10445_10747 , \10446_10748 , \10447_10749 , \10448_10750 , \10449_10751 , \10450_10752 , \10451_10753 , \10452_10754 , \10453_10755 , \10454_10756 , \10455_10757 , \10456_10758 , \10457_10759 , \10458_10760 , \10459_10761 , \10460_10762 , \10461_10763 , \10462_10764 , \10463_10765 , \10464_10766 , \10465_10767 , \10466_10768 , \10467_10769 , \10468_10770 , \10469_10771 , \10470_10772 , \10471_10773 , \10472_10774 , \10473_10775 , \10474_10776 , \10475_10777 , \10476_10778 );
and \U$1716 ( \10478_10780 , RIee2ba20_4955, \9163_9462 );
and \U$1717 ( \10479_10781 , RIfc93ba8_6703, \9165_9464 );
and \U$1718 ( \10480_10782 , RIfc77de0_6386, \9167_9466 );
and \U$1719 ( \10481_10783 , RIee27ad8_4910, \9169_9468 );
and \U$1720 ( \10482_10784 , RIfe9d668_8135, \9171_9470 );
and \U$1721 ( \10483_10785 , RIfea8bd0_8236, \9173_9472 );
and \U$1722 ( \10484_10786 , RIdf26458_1812, \9175_9474 );
and \U$1723 ( \10485_10787 , RIfe9d7d0_8136, \9177_9476 );
and \U$1724 ( \10486_10788 , RIfcb1c98_7045, \9179_9478 );
and \U$1725 ( \10487_10789 , RIee26cc8_4900, \9181_9480 );
and \U$1726 ( \10488_10790 , RIdf22ab0_1771, \9183_9482 );
and \U$1727 ( \10489_10791 , RIfcc0068_7207, \9185_9484 );
and \U$1728 ( \10490_10792 , RIdf21598_1756, \9187_9486 );
and \U$1729 ( \10491_10793 , RIdf1f6a8_1734, \9189_9488 );
and \U$1730 ( \10492_10794 , RIdf1aef0_1683, \9191_9490 );
and \U$1731 ( \10493_10795 , RIfe9d938_8137, \9193_9492 );
and \U$1732 ( \10494_10796 , RIdf16cd8_1636, \9195_9494 );
and \U$1733 ( \10495_10797 , RIdf13fd8_1604, \9197_9496 );
and \U$1734 ( \10496_10798 , RIdf112d8_1572, \9199_9498 );
and \U$1735 ( \10497_10799 , RIdf0e5d8_1540, \9201_9500 );
and \U$1736 ( \10498_10800 , RIdf0b8d8_1508, \9203_9502 );
and \U$1737 ( \10499_10801 , RIdf08bd8_1476, \9205_9504 );
and \U$1738 ( \10500_10802 , RIdf05ed8_1444, \9207_9506 );
and \U$1739 ( \10501_10803 , RIdf031d8_1412, \9209_9508 );
and \U$1740 ( \10502_10804 , RIdefd7d8_1348, \9211_9510 );
and \U$1741 ( \10503_10805 , RIdefaad8_1316, \9213_9512 );
and \U$1742 ( \10504_10806 , RIdef7dd8_1284, \9215_9514 );
and \U$1743 ( \10505_10807 , RIdef50d8_1252, \9217_9516 );
and \U$1744 ( \10506_10808 , RIdef23d8_1220, \9219_9518 );
and \U$1745 ( \10507_10809 , RIdeef6d8_1188, \9221_9520 );
and \U$1746 ( \10508_10810 , RIdeec9d8_1156, \9223_9522 );
and \U$1747 ( \10509_10811 , RIdee9cd8_1124, \9225_9524 );
and \U$1748 ( \10510_10812 , RIfc942b0_6708, \9227_9526 );
and \U$1749 ( \10511_10813 , RIfcde6f8_7553, \9229_9528 );
and \U$1750 ( \10512_10814 , RIfcd1138_7401, \9231_9530 );
and \U$1751 ( \10513_10815 , RIfcde860_7554, \9233_9532 );
and \U$1752 ( \10514_10816 , RIdee4878_1064, \9235_9534 );
and \U$1753 ( \10515_10817 , RIdee2af0_1043, \9237_9536 );
and \U$1754 ( \10516_10818 , RIdee0a98_1020, \9239_9538 );
and \U$1755 ( \10517_10819 , RIdede8d8_996, \9241_9540 );
and \U$1756 ( \10518_10820 , RIfc5c9f0_6076, \9243_9542 );
and \U$1757 ( \10519_10821 , RIee22240_4847, \9245_9544 );
and \U$1758 ( \10520_10822 , RIfcc8768_7303, \9247_9546 );
and \U$1759 ( \10521_10823 , RIee21160_4835, \9249_9548 );
and \U$1760 ( \10522_10824 , RIded95e0_937, \9251_9550 );
and \U$1761 ( \10523_10825 , RIded7150_911, \9253_9552 );
and \U$1762 ( \10524_10826 , RIded5260_889, \9255_9554 );
and \U$1763 ( \10525_10827 , RIfea76b8_8221, \9257_9556 );
and \U$1764 ( \10526_10828 , RIded0508_834, \9259_9558 );
and \U$1765 ( \10527_10829 , RIdecd808_802, \9261_9560 );
and \U$1766 ( \10528_10830 , RIdecab08_770, \9263_9562 );
and \U$1767 ( \10529_10831 , RIdec7e08_738, \9265_9564 );
and \U$1768 ( \10530_10832 , RIdeb4308_514, \9267_9566 );
and \U$1769 ( \10531_10833 , RIde96290_322, \9269_9568 );
and \U$1770 ( \10532_10834 , RIe16df10_2628, \9271_9570 );
and \U$1771 ( \10533_10835 , RIe159d08_2399, \9273_9572 );
and \U$1772 ( \10534_10836 , RIe143508_2143, \9275_9574 );
and \U$1773 ( \10535_10837 , RIdf37f00_2013, \9277_9576 );
and \U$1774 ( \10536_10838 , RIdf2c560_1881, \9279_9578 );
and \U$1775 ( \10537_10839 , RIdf1cde0_1705, \9281_9580 );
and \U$1776 ( \10538_10840 , RIdf004d8_1380, \9283_9582 );
and \U$1777 ( \10539_10841 , RIdee6fd8_1092, \9285_9584 );
and \U$1778 ( \10540_10842 , RIdedbd40_965, \9287_9586 );
and \U$1779 ( \10541_10843 , RIde7c1d8_195, \9289_9588 );
or \U$1780 ( \10542_10844 , \10478_10780 , \10479_10781 , \10480_10782 , \10481_10783 , \10482_10784 , \10483_10785 , \10484_10786 , \10485_10787 , \10486_10788 , \10487_10789 , \10488_10790 , \10489_10791 , \10490_10792 , \10491_10793 , \10492_10794 , \10493_10795 , \10494_10796 , \10495_10797 , \10496_10798 , \10497_10799 , \10498_10800 , \10499_10801 , \10500_10802 , \10501_10803 , \10502_10804 , \10503_10805 , \10504_10806 , \10505_10807 , \10506_10808 , \10507_10809 , \10508_10810 , \10509_10811 , \10510_10812 , \10511_10813 , \10512_10814 , \10513_10815 , \10514_10816 , \10515_10817 , \10516_10818 , \10517_10819 , \10518_10820 , \10519_10821 , \10520_10822 , \10521_10823 , \10522_10824 , \10523_10825 , \10524_10826 , \10525_10827 , \10526_10828 , \10527_10829 , \10528_10830 , \10529_10831 , \10530_10832 , \10531_10833 , \10532_10834 , \10533_10835 , \10534_10836 , \10535_10837 , \10536_10838 , \10537_10839 , \10538_10840 , \10539_10841 , \10540_10842 , \10541_10843 );
or \U$1781 ( \10543_10845 , \10477_10779 , \10542_10844 );
_DC \g45e3/U$1 ( \10544 , \10543_10845 , \9298_9597 );
and \U$1782 ( \10545_10847 , RIe19d3a0_3166, \8760_9059 );
and \U$1783 ( \10546_10848 , RIe19a6a0_3134, \8762_9061 );
and \U$1784 ( \10547_10849 , RIfcb2c10_7056, \8764_9063 );
and \U$1785 ( \10548_10850 , RIe1979a0_3102, \8766_9065 );
and \U$1786 ( \10549_10851 , RIfc923c0_6686, \8768_9067 );
and \U$1787 ( \10550_10852 , RIe194ca0_3070, \8770_9069 );
and \U$1788 ( \10551_10853 , RIe191fa0_3038, \8772_9071 );
and \U$1789 ( \10552_10854 , RIe18f2a0_3006, \8774_9073 );
and \U$1790 ( \10553_10855 , RIe1898a0_2942, \8776_9075 );
and \U$1791 ( \10554_10856 , RIe186ba0_2910, \8778_9077 );
and \U$1792 ( \10555_10857 , RIfc422a8_5775, \8780_9079 );
and \U$1793 ( \10556_10858 , RIe183ea0_2878, \8782_9081 );
and \U$1794 ( \10557_10859 , RIfcbecb8_7193, \8784_9083 );
and \U$1795 ( \10558_10860 , RIe1811a0_2846, \8786_9085 );
and \U$1796 ( \10559_10861 , RIe17e4a0_2814, \8788_9087 );
and \U$1797 ( \10560_10862 , RIe17b7a0_2782, \8790_9089 );
and \U$1798 ( \10561_10863 , RIf142250_5212, \8792_9091 );
and \U$1799 ( \10562_10864 , RIf140bd0_5196, \8794_9093 );
and \U$1800 ( \10563_10865 , RIfec43f8_8353, \8796_9095 );
and \U$1801 ( \10564_10866 , RIe175968_2715, \8798_9097 );
and \U$1802 ( \10565_10867 , RIfc79b68_6407, \8800_9099 );
and \U$1803 ( \10566_10868 , RIf13efb0_5176, \8802_9101 );
and \U$1804 ( \10567_10869 , RIfc92528_6687, \8804_9103 );
and \U$1805 ( \10568_10870 , RIfcb2aa8_7055, \8806_9105 );
and \U$1806 ( \10569_10871 , RIfcd8320_7482, \8808_9107 );
and \U$1807 ( \10570_10872 , RIfcea200_7686, \8810_9109 );
and \U$1808 ( \10571_10873 , RIfc79898_6405, \8812_9111 );
and \U$1809 ( \10572_10874 , RIe1734d8_2689, \8814_9113 );
and \U$1810 ( \10573_10875 , RIfcd7948_7475, \8816_9115 );
and \U$1811 ( \10574_10876 , RIfcd7678_7473, \8818_9117 );
and \U$1812 ( \10575_10877 , RIf16e170_5712, \8820_9119 );
and \U$1813 ( \10576_10878 , RIfc927f8_6689, \8822_9121 );
and \U$1814 ( \10577_10879 , RIfc92960_6690, \8824_9123 );
and \U$1815 ( \10578_10880 , RIe2236f8_4693, \8826_9125 );
and \U$1816 ( \10579_10881 , RIfc795c8_6403, \8828_9127 );
and \U$1817 ( \10580_10882 , RIe2209f8_4661, \8830_9129 );
and \U$1818 ( \10581_10883 , RIf16ad68_5675, \8832_9131 );
and \U$1819 ( \10582_10884 , RIe21dcf8_4629, \8834_9133 );
and \U$1820 ( \10583_10885 , RIe2182f8_4565, \8836_9135 );
and \U$1821 ( \10584_10886 , RIe2155f8_4533, \8838_9137 );
and \U$1822 ( \10585_10887 , RIfe9d398_8133, \8840_9139 );
and \U$1823 ( \10586_10888 , RIe2128f8_4501, \8842_9141 );
and \U$1824 ( \10587_10889 , RIfcdb9f8_7521, \8844_9143 );
and \U$1825 ( \10588_10890 , RIe20fbf8_4469, \8846_9145 );
and \U$1826 ( \10589_10891 , RIfc41d08_5771, \8848_9147 );
and \U$1827 ( \10590_10892 , RIe20cef8_4437, \8850_9149 );
and \U$1828 ( \10591_10893 , RIe20a1f8_4405, \8852_9151 );
and \U$1829 ( \10592_10894 , RIe2074f8_4373, \8854_9153 );
and \U$1830 ( \10593_10895 , RIfcd7510_7472, \8856_9155 );
and \U$1831 ( \10594_10896 , RIf166010_5620, \8858_9157 );
and \U$1832 ( \10595_10897 , RIfe9d230_8132, \8860_9159 );
and \U$1833 ( \10596_10898 , RIe2008b0_4296, \8862_9161 );
and \U$1834 ( \10597_10899 , RIf165098_5609, \8864_9163 );
and \U$1835 ( \10598_10900 , RIfc41ba0_5770, \8866_9165 );
and \U$1836 ( \10599_10901 , RIfc41a38_5769, \8868_9167 );
and \U$1837 ( \10600_10902 , RIfc92c30_6692, \8870_9169 );
and \U$1838 ( \10601_10903 , RIfc418d0_5768, \8872_9171 );
and \U$1839 ( \10602_10904 , RIfc79190_6400, \8874_9173 );
and \U$1840 ( \10603_10905 , RIe1fcad0_4252, \8876_9175 );
and \U$1841 ( \10604_10906 , RIfec4560_8354, \8878_9177 );
and \U$1842 ( \10605_10907 , RIfc79028_6399, \8880_9179 );
and \U$1843 ( \10606_10908 , RIfcbf258_7197, \8882_9181 );
and \U$1844 ( \10607_10909 , RIfcc1df0_7228, \8884_9183 );
and \U$1845 ( \10608_10910 , RIfcd81b8_7481, \8886_9185 );
or \U$1846 ( \10609_10911 , \10545_10847 , \10546_10848 , \10547_10849 , \10548_10850 , \10549_10851 , \10550_10852 , \10551_10853 , \10552_10854 , \10553_10855 , \10554_10856 , \10555_10857 , \10556_10858 , \10557_10859 , \10558_10860 , \10559_10861 , \10560_10862 , \10561_10863 , \10562_10864 , \10563_10865 , \10564_10866 , \10565_10867 , \10566_10868 , \10567_10869 , \10568_10870 , \10569_10871 , \10570_10872 , \10571_10873 , \10572_10874 , \10573_10875 , \10574_10876 , \10575_10877 , \10576_10878 , \10577_10879 , \10578_10880 , \10579_10881 , \10580_10882 , \10581_10883 , \10582_10884 , \10583_10885 , \10584_10886 , \10585_10887 , \10586_10888 , \10587_10889 , \10588_10890 , \10589_10891 , \10590_10892 , \10591_10893 , \10592_10894 , \10593_10895 , \10594_10896 , \10595_10897 , \10596_10898 , \10597_10899 , \10598_10900 , \10599_10901 , \10600_10902 , \10601_10903 , \10602_10904 , \10603_10905 , \10604_10906 , \10605_10907 , \10606_10908 , \10607_10909 , \10608_10910 );
and \U$1847 ( \10610_10912 , RIfc92d98_6693, \8889_9188 );
and \U$1848 ( \10611_10913 , RIfc5b4d8_6061, \8891_9190 );
and \U$1849 ( \10612_10914 , RIfcd77e0_7474, \8893_9192 );
and \U$1850 ( \10613_10915 , RIe1fa0a0_4222, \8895_9194 );
and \U$1851 ( \10614_10916 , RIf156188_5439, \8897_9196 );
and \U$1852 ( \10615_10917 , RIfe9d500_8134, \8899_9198 );
and \U$1853 ( \10616_10918 , RIf1546d0_5420, \8901_9200 );
and \U$1854 ( \10617_10919 , RIe1f5348_4167, \8903_9202 );
and \U$1855 ( \10618_10920 , RIfec4830_8356, \8905_9204 );
and \U$1856 ( \10619_10921 , RIfec46c8_8355, \8907_9206 );
and \U$1857 ( \10620_10922 , RIf1508f0_5376, \8909_9208 );
and \U$1858 ( \10621_10923 , RIe1f3020_4142, \8911_9210 );
and \U$1859 ( \10622_10924 , RIfce3180_7606, \8913_9212 );
and \U$1860 ( \10623_10925 , RIfce8fb8_7673, \8915_9214 );
and \U$1861 ( \10624_10926 , RIfcbf690_7200, \8917_9216 );
and \U$1862 ( \10625_10927 , RIe1edd28_4083, \8919_9218 );
and \U$1863 ( \10626_10928 , RIe1eb460_4054, \8921_9220 );
and \U$1864 ( \10627_10929 , RIe1e8760_4022, \8923_9222 );
and \U$1865 ( \10628_10930 , RIe1e5a60_3990, \8925_9224 );
and \U$1866 ( \10629_10931 , RIe1e2d60_3958, \8927_9226 );
and \U$1867 ( \10630_10932 , RIe1e0060_3926, \8929_9228 );
and \U$1868 ( \10631_10933 , RIe1dd360_3894, \8931_9230 );
and \U$1869 ( \10632_10934 , RIe1da660_3862, \8933_9232 );
and \U$1870 ( \10633_10935 , RIe1d7960_3830, \8935_9234 );
and \U$1871 ( \10634_10936 , RIe1d1f60_3766, \8937_9236 );
and \U$1872 ( \10635_10937 , RIe1cf260_3734, \8939_9238 );
and \U$1873 ( \10636_10938 , RIe1cc560_3702, \8941_9240 );
and \U$1874 ( \10637_10939 , RIe1c9860_3670, \8943_9242 );
and \U$1875 ( \10638_10940 , RIe1c6b60_3638, \8945_9244 );
and \U$1876 ( \10639_10941 , RIe1c3e60_3606, \8947_9246 );
and \U$1877 ( \10640_10942 , RIe1c1160_3574, \8949_9248 );
and \U$1878 ( \10641_10943 , RIe1be460_3542, \8951_9250 );
and \U$1879 ( \10642_10944 , RIfe9d0c8_8131, \8953_9252 );
and \U$1880 ( \10643_10945 , RIfe9cc90_8128, \8955_9254 );
and \U$1881 ( \10644_10946 , RIe1b9168_3483, \8957_9256 );
and \U$1882 ( \10645_10947 , RIe1b7110_3460, \8959_9258 );
and \U$1883 ( \10646_10948 , RIf14a3b0_5304, \8961_9260 );
and \U$1884 ( \10647_10949 , RIfe9cb28_8127, \8963_9262 );
and \U$1885 ( \10648_10950 , RIfe9cf60_8130, \8965_9264 );
and \U$1886 ( \10649_10951 , RIfe9c9c0_8126, \8967_9266 );
and \U$1887 ( \10650_10952 , RIfce2208_7595, \8969_9268 );
and \U$1888 ( \10651_10953 , RIfce9558_7677, \8971_9270 );
and \U$1889 ( \10652_10954 , RIfe9c858_8125, \8973_9272 );
and \U$1890 ( \10653_10955 , RIfe9cdf8_8129, \8975_9274 );
and \U$1891 ( \10654_10956 , RIf147110_5268, \8977_9276 );
and \U$1892 ( \10655_10957 , RIf146468_5259, \8979_9278 );
and \U$1893 ( \10656_10958 , RIe1ac2b0_3336, \8981_9280 );
and \U$1894 ( \10657_10959 , RIe1aaac8_3319, \8983_9282 );
and \U$1895 ( \10658_10960 , RIe1a87a0_3294, \8985_9284 );
and \U$1896 ( \10659_10961 , RIe1a5aa0_3262, \8987_9286 );
and \U$1897 ( \10660_10962 , RIe1a2da0_3230, \8989_9288 );
and \U$1898 ( \10661_10963 , RIe1a00a0_3198, \8991_9290 );
and \U$1899 ( \10662_10964 , RIe18c5a0_2974, \8993_9292 );
and \U$1900 ( \10663_10965 , RIe178aa0_2750, \8995_9294 );
and \U$1901 ( \10664_10966 , RIe2263f8_4725, \8997_9296 );
and \U$1902 ( \10665_10967 , RIe21aff8_4597, \8999_9298 );
and \U$1903 ( \10666_10968 , RIe2047f8_4341, \9001_9300 );
and \U$1904 ( \10667_10969 , RIe1fe858_4273, \9003_9302 );
and \U$1905 ( \10668_10970 , RIe1f7c10_4196, \9005_9304 );
and \U$1906 ( \10669_10971 , RIe1f0758_4113, \9007_9306 );
and \U$1907 ( \10670_10972 , RIe1d4c60_3798, \9009_9308 );
and \U$1908 ( \10671_10973 , RIe1bb760_3510, \9011_9310 );
and \U$1909 ( \10672_10974 , RIe1ae5d8_3361, \9013_9312 );
and \U$1910 ( \10673_10975 , RIe170c10_2660, \9015_9314 );
or \U$1911 ( \10674_10976 , \10610_10912 , \10611_10913 , \10612_10914 , \10613_10915 , \10614_10916 , \10615_10917 , \10616_10918 , \10617_10919 , \10618_10920 , \10619_10921 , \10620_10922 , \10621_10923 , \10622_10924 , \10623_10925 , \10624_10926 , \10625_10927 , \10626_10928 , \10627_10929 , \10628_10930 , \10629_10931 , \10630_10932 , \10631_10933 , \10632_10934 , \10633_10935 , \10634_10936 , \10635_10937 , \10636_10938 , \10637_10939 , \10638_10940 , \10639_10941 , \10640_10942 , \10641_10943 , \10642_10944 , \10643_10945 , \10644_10946 , \10645_10947 , \10646_10948 , \10647_10949 , \10648_10950 , \10649_10951 , \10650_10952 , \10651_10953 , \10652_10954 , \10653_10955 , \10654_10956 , \10655_10957 , \10656_10958 , \10657_10959 , \10658_10960 , \10659_10961 , \10660_10962 , \10661_10963 , \10662_10964 , \10663_10965 , \10664_10966 , \10665_10967 , \10666_10968 , \10667_10969 , \10668_10970 , \10669_10971 , \10670_10972 , \10671_10973 , \10672_10974 , \10673_10975 );
or \U$1912 ( \10675_10977 , \10609_10911 , \10674_10976 );
_DC \g4667/U$1 ( \10676 , \10675_10977 , \9024_9323 );
xor g4668_GF_PartitionCandidate( \10677_10979_nG4668 , \10544 , \10676 );
buf \U$1913 ( \10678_10980 , \10677_10979_nG4668 );
xor \U$1914 ( \10679_10981 , \10678_10980 , \10389_10691 );
not \U$1915 ( \10680_10982 , \10389_10691 );
and \U$1916 ( \10681_10983 , \10679_10981 , \10680_10982 );
and \U$1917 ( \10682_10984 , \10385_10687 , \10681_10983 );
_DC \g657a/U$1 ( \10683 , \10543_10845 , \9298_9597 );
_DC \g657b/U$1 ( \10684 , \10675_10977 , \9024_9323 );
and g657c_GF_PartitionCandidate( \10685_10987_nG657c , \10683 , \10684 );
buf \U$1918 ( \10686_10988 , \10685_10987_nG657c );
and \U$1919 ( \10687_10989 , \10686_10988 , \10389_10691 );
nor \U$1920 ( \10688_10990 , \10682_10984 , \10687_10989 );
xnor \U$1921 ( \10689_10991 , \10688_10990 , \10678_10980 );
not \U$1922 ( \10690_10992 , \10390_10692 );
and \U$1923 ( \10691_10993 , \10690_10992 , \10678_10980 );
xor \U$1924 ( \10692_10994 , \10689_10991 , \10691_10993 );
buf g9c0b_GF_PartitionCandidate( \10693_10995_nG9c0b , \10692_10994 );
and \U$1925 ( \10694_10996 , \10402_10704 , \10693_10995_nG9c0b );
or \U$1926 ( \10695_10997 , \10412_10714 , \10694_10996 );
xor \U$1927 ( \10696_10998 , \10399_10703 , \10695_10997 );
buf \U$1928 ( \10697_10999 , \10696_10998 );
buf \U$1930 ( \10698_11000 , \10697_10999 );
and \U$1931 ( \10699_11001 , \10408_10713 , \10698_11000 );
buf \U$1932 ( \10700_11002 , \10699_11001 );
and \U$1933 ( \10701_11003 , \10411_10707 , \10693_10995_nG9c0b );
and \U$1934 ( \10702_11004 , \10686_10988 , \10681_10983 );
and \U$1935 ( \10703_11005 , RIdec6080_717, \9034_9333 );
and \U$1936 ( \10704_11006 , RIdec3380_685, \9036_9335 );
and \U$1937 ( \10705_11007 , RIee204b8_4826, \9038_9337 );
and \U$1938 ( \10706_11008 , RIdec0680_653, \9040_9339 );
and \U$1939 ( \10707_11009 , RIfcd70d8_7469, \9042_9341 );
and \U$1940 ( \10708_11010 , RIdebd980_621, \9044_9343 );
and \U$1941 ( \10709_11011 , RIdebac80_589, \9046_9345 );
and \U$1942 ( \10710_11012 , RIdeb7f80_557, \9048_9347 );
and \U$1943 ( \10711_11013 , RIfcbe448_7187, \9050_9349 );
and \U$1944 ( \10712_11014 , RIdeb2580_493, \9052_9351 );
and \U$1945 ( \10713_11015 , RIfcb3480_7062, \9054_9353 );
and \U$1946 ( \10714_11016 , RIdeaf880_461, \9056_9355 );
and \U$1947 ( \10715_11017 , RIfc43928_5791, \9058_9357 );
and \U$1948 ( \10716_11018 , RIdeac1a8_429, \9060_9359 );
and \U$1949 ( \10717_11019 , RIdea58a8_397, \9062_9361 );
and \U$1950 ( \10718_11020 , RIde9efa8_365, \9064_9363 );
and \U$1951 ( \10719_11021 , RIfcd88c0_7486, \9066_9365 );
and \U$1952 ( \10720_11022 , RIee1c408_4780, \9068_9367 );
and \U$1953 ( \10721_11023 , RIfcc77f0_7292, \9070_9369 );
and \U$1954 ( \10722_11024 , RIfea04d0_8168, \9072_9371 );
and \U$1955 ( \10723_11025 , RIde92438_303, \9074_9373 );
and \U$1956 ( \10724_11026 , RIde8ec70_286, \9076_9375 );
and \U$1957 ( \10725_11027 , RIde8aad0_266, \9078_9377 );
and \U$1958 ( \10726_11028 , RIde86930_246, \9080_9379 );
and \U$1959 ( \10727_11029 , RIfca31c0_6878, \9082_9381 );
and \U$1960 ( \10728_11030 , RIfc59a20_6042, \9084_9383 );
and \U$1961 ( \10729_11031 , RIfcd1de0_7410, \9086_9385 );
and \U$1962 ( \10730_11032 , RIfc91448_6675, \9088_9387 );
and \U$1963 ( \10731_11033 , RIfc97280_6742, \9090_9389 );
and \U$1964 ( \10732_11034 , RIe16c188_2607, \9092_9391 );
and \U$1965 ( \10733_11035 , RIfc97118_6741, \9094_9393 );
and \U$1966 ( \10734_11036 , RIe168948_2567, \9096_9395 );
and \U$1967 ( \10735_11037 , RIe166080_2538, \9098_9397 );
and \U$1968 ( \10736_11038 , RIe163380_2506, \9100_9399 );
and \U$1969 ( \10737_11039 , RIee37ac8_5092, \9102_9401 );
and \U$1970 ( \10738_11040 , RIe160680_2474, \9104_9403 );
and \U$1971 ( \10739_11041 , RIfcd1c78_7409, \9106_9405 );
and \U$1972 ( \10740_11042 , RIe15d980_2442, \9108_9407 );
and \U$1973 ( \10741_11043 , RIe157f80_2378, \9110_9409 );
and \U$1974 ( \10742_11044 , RIe155280_2346, \9112_9411 );
and \U$1975 ( \10743_11045 , RIfc3f530_5746, \9114_9413 );
and \U$1976 ( \10744_11046 , RIe152580_2314, \9116_9415 );
and \U$1977 ( \10745_11047 , RIee35368_5064, \9118_9417 );
and \U$1978 ( \10746_11048 , RIe14f880_2282, \9120_9419 );
and \U$1979 ( \10747_11049 , RIfc7a3d8_6413, \9122_9421 );
and \U$1980 ( \10748_11050 , RIe14cb80_2250, \9124_9423 );
and \U$1981 ( \10749_11051 , RIe149e80_2218, \9126_9425 );
and \U$1982 ( \10750_11052 , RIe147180_2186, \9128_9427 );
and \U$1983 ( \10751_11053 , RIfc42b18_5781, \9130_9429 );
and \U$1984 ( \10752_11054 , RIfc7a270_6412, \9132_9431 );
and \U$1985 ( \10753_11055 , RIfc5a560_6050, \9134_9433 );
and \U$1986 ( \10754_11056 , RIfc96b78_6737, \9136_9435 );
and \U$1987 ( \10755_11057 , RIfea6fb0_8216, \9138_9437 );
and \U$1988 ( \10756_11058 , RIe13f5c0_2098, \9140_9439 );
and \U$1989 ( \10757_11059 , RIdf3d4c8_2074, \9142_9441 );
and \U$1990 ( \10758_11060 , RIdf3b038_2048, \9144_9443 );
and \U$1991 ( \10759_11061 , RIfce5bb0_7636, \9146_9445 );
and \U$1992 ( \10760_11062 , RIee2fc38_5002, \9148_9447 );
and \U$1993 ( \10761_11063 , RIfc91cb8_6681, \9150_9449 );
and \U$1994 ( \10762_11064 , RIee2d910_4977, \9152_9451 );
and \U$1995 ( \10763_11065 , RIdf362e0_1993, \9154_9453 );
and \U$1996 ( \10764_11066 , RIdf33e50_1967, \9156_9455 );
and \U$1997 ( \10765_11067 , RIdf31c90_1943, \9158_9457 );
and \U$1998 ( \10766_11068 , RIdf2fda0_1921, \9160_9459 );
or \U$1999 ( \10767_11069 , \10703_11005 , \10704_11006 , \10705_11007 , \10706_11008 , \10707_11009 , \10708_11010 , \10709_11011 , \10710_11012 , \10711_11013 , \10712_11014 , \10713_11015 , \10714_11016 , \10715_11017 , \10716_11018 , \10717_11019 , \10718_11020 , \10719_11021 , \10720_11022 , \10721_11023 , \10722_11024 , \10723_11025 , \10724_11026 , \10725_11027 , \10726_11028 , \10727_11029 , \10728_11030 , \10729_11031 , \10730_11032 , \10731_11033 , \10732_11034 , \10733_11035 , \10734_11036 , \10735_11037 , \10736_11038 , \10737_11039 , \10738_11040 , \10739_11041 , \10740_11042 , \10741_11043 , \10742_11044 , \10743_11045 , \10744_11046 , \10745_11047 , \10746_11048 , \10747_11049 , \10748_11050 , \10749_11051 , \10750_11052 , \10751_11053 , \10752_11054 , \10753_11055 , \10754_11056 , \10755_11057 , \10756_11058 , \10757_11059 , \10758_11060 , \10759_11061 , \10760_11062 , \10761_11063 , \10762_11064 , \10763_11065 , \10764_11066 , \10765_11067 , \10766_11068 );
and \U$2000 ( \10768_11070 , RIfc43658_5789, \9163_9462 );
and \U$2001 ( \10769_11071 , RIfc59e58_6045, \9165_9464 );
and \U$2002 ( \10770_11072 , RIfc96fb0_6740, \9167_9466 );
and \U$2003 ( \10771_11073 , RIfc7ac48_6419, \9169_9468 );
and \U$2004 ( \10772_11074 , RIfea0368_8167, \9171_9470 );
and \U$2005 ( \10773_11075 , RIdf28bb8_1840, \9173_9472 );
and \U$2006 ( \10774_11076 , RIdf26cc8_1818, \9175_9474 );
and \U$2007 ( \10775_11077 , RIdf25210_1799, \9177_9476 );
and \U$2008 ( \10776_11078 , RIfc91718_6677, \9179_9478 );
and \U$2009 ( \10777_11079 , RIfcb3318_7061, \9181_9480 );
and \U$2010 ( \10778_11080 , RIfc919e8_6679, \9183_9482 );
and \U$2011 ( \10779_11081 , RIfc91880_6678, \9185_9484 );
and \U$2012 ( \10780_11082 , RIfc430b8_5785, \9187_9486 );
and \U$2013 ( \10781_11083 , RIdf20350_1743, \9189_9488 );
and \U$2014 ( \10782_11084 , RIfc7a978_6417, \9191_9490 );
and \U$2015 ( \10783_11085 , RIdf19e10_1671, \9193_9492 );
and \U$2016 ( \10784_11086 , RIdf17c50_1647, \9195_9494 );
and \U$2017 ( \10785_11087 , RIdf14f50_1615, \9197_9496 );
and \U$2018 ( \10786_11088 , RIdf12250_1583, \9199_9498 );
and \U$2019 ( \10787_11089 , RIdf0f550_1551, \9201_9500 );
and \U$2020 ( \10788_11090 , RIdf0c850_1519, \9203_9502 );
and \U$2021 ( \10789_11091 , RIdf09b50_1487, \9205_9504 );
and \U$2022 ( \10790_11092 , RIdf06e50_1455, \9207_9506 );
and \U$2023 ( \10791_11093 , RIdf04150_1423, \9209_9508 );
and \U$2024 ( \10792_11094 , RIdefe750_1359, \9211_9510 );
and \U$2025 ( \10793_11095 , RIdefba50_1327, \9213_9512 );
and \U$2026 ( \10794_11096 , RIdef8d50_1295, \9215_9514 );
and \U$2027 ( \10795_11097 , RIdef6050_1263, \9217_9516 );
and \U$2028 ( \10796_11098 , RIdef3350_1231, \9219_9518 );
and \U$2029 ( \10797_11099 , RIdef0650_1199, \9221_9520 );
and \U$2030 ( \10798_11100 , RIdeed950_1167, \9223_9522 );
and \U$2031 ( \10799_11101 , RIdeeac50_1135, \9225_9524 );
and \U$2032 ( \10800_11102 , RIfcd1b10_7408, \9227_9526 );
and \U$2033 ( \10801_11103 , RIfc968a8_6735, \9229_9528 );
and \U$2034 ( \10802_11104 , RIfc91f88_6683, \9231_9530 );
and \U$2035 ( \10803_11105 , RIfcdfc10_7568, \9233_9532 );
and \U$2036 ( \10804_11106 , RIfea99e0_8246, \9235_9534 );
and \U$2037 ( \10805_11107 , RIdee3630_1051, \9237_9536 );
and \U$2038 ( \10806_11108 , RIdee1308_1026, \9239_9538 );
and \U$2039 ( \10807_11109 , RIdedf2b0_1003, \9241_9540 );
and \U$2040 ( \10808_11110 , RIfcc7d90_7296, \9243_9542 );
and \U$2041 ( \10809_11111 , RIfcd85f0_7484, \9245_9544 );
and \U$2042 ( \10810_11112 , RIfce3888_7611, \9247_9546 );
and \U$2043 ( \10811_11113 , RIfc5a830_6052, \9249_9548 );
and \U$2044 ( \10812_11114 , RIdeda3f0_947, \9251_9550 );
and \U$2045 ( \10813_11115 , RIfea9878_8245, \9253_9552 );
and \U$2046 ( \10814_11116 , RIded5f08_898, \9255_9554 );
and \U$2047 ( \10815_11117 , RIded37a8_870, \9257_9556 );
and \U$2048 ( \10816_11118 , RIded1480_845, \9259_9558 );
and \U$2049 ( \10817_11119 , RIdece780_813, \9261_9560 );
and \U$2050 ( \10818_11120 , RIdecba80_781, \9263_9562 );
and \U$2051 ( \10819_11121 , RIdec8d80_749, \9265_9564 );
and \U$2052 ( \10820_11122 , RIdeb5280_525, \9267_9566 );
and \U$2053 ( \10821_11123 , RIde986a8_333, \9269_9568 );
and \U$2054 ( \10822_11124 , RIe16ee88_2639, \9271_9570 );
and \U$2055 ( \10823_11125 , RIe15ac80_2410, \9273_9572 );
and \U$2056 ( \10824_11126 , RIe144480_2154, \9275_9574 );
and \U$2057 ( \10825_11127 , RIdf38e78_2024, \9277_9576 );
and \U$2058 ( \10826_11128 , RIdf2d4d8_1892, \9279_9578 );
and \U$2059 ( \10827_11129 , RIdf1dd58_1716, \9281_9580 );
and \U$2060 ( \10828_11130 , RIdf01450_1391, \9283_9582 );
and \U$2061 ( \10829_11131 , RIdee7f50_1103, \9285_9584 );
and \U$2062 ( \10830_11132 , RIdedccb8_976, \9287_9586 );
and \U$2063 ( \10831_11133 , RIde7e5f0_206, \9289_9588 );
or \U$2064 ( \10832_11134 , \10768_11070 , \10769_11071 , \10770_11072 , \10771_11073 , \10772_11074 , \10773_11075 , \10774_11076 , \10775_11077 , \10776_11078 , \10777_11079 , \10778_11080 , \10779_11081 , \10780_11082 , \10781_11083 , \10782_11084 , \10783_11085 , \10784_11086 , \10785_11087 , \10786_11088 , \10787_11089 , \10788_11090 , \10789_11091 , \10790_11092 , \10791_11093 , \10792_11094 , \10793_11095 , \10794_11096 , \10795_11097 , \10796_11098 , \10797_11099 , \10798_11100 , \10799_11101 , \10800_11102 , \10801_11103 , \10802_11104 , \10803_11105 , \10804_11106 , \10805_11107 , \10806_11108 , \10807_11109 , \10808_11110 , \10809_11111 , \10810_11112 , \10811_11113 , \10812_11114 , \10813_11115 , \10814_11116 , \10815_11117 , \10816_11118 , \10817_11119 , \10818_11120 , \10819_11121 , \10820_11122 , \10821_11123 , \10822_11124 , \10823_11125 , \10824_11126 , \10825_11127 , \10826_11128 , \10827_11129 , \10828_11130 , \10829_11131 , \10830_11132 , \10831_11133 );
or \U$2065 ( \10833_11135 , \10767_11069 , \10832_11134 );
_DC \g657d/U$1 ( \10834 , \10833_11135 , \9298_9597 );
and \U$2066 ( \10835_11137 , RIe19e318_3177, \8760_9059 );
and \U$2067 ( \10836_11138 , RIe19b618_3145, \8762_9061 );
and \U$2068 ( \10837_11139 , RIfc8f3f0_6652, \8764_9063 );
and \U$2069 ( \10838_11140 , RIe198918_3113, \8766_9065 );
and \U$2070 ( \10839_11141 , RIf144b18_5241, \8768_9067 );
and \U$2071 ( \10840_11142 , RIe195c18_3081, \8770_9069 );
and \U$2072 ( \10841_11143 , RIe192f18_3049, \8772_9071 );
and \U$2073 ( \10842_11144 , RIe190218_3017, \8774_9073 );
and \U$2074 ( \10843_11145 , RIe18a818_2953, \8776_9075 );
and \U$2075 ( \10844_11146 , RIe187b18_2921, \8778_9077 );
and \U$2076 ( \10845_11147 , RIf143d08_5231, \8780_9079 );
and \U$2077 ( \10846_11148 , RIe184e18_2889, \8782_9081 );
and \U$2078 ( \10847_11149 , RIfcb3cf0_7068, \8784_9083 );
and \U$2079 ( \10848_11150 , RIe182118_2857, \8786_9085 );
and \U$2080 ( \10849_11151 , RIe17f418_2825, \8788_9087 );
and \U$2081 ( \10850_11152 , RIe17c718_2793, \8790_9089 );
and \U$2082 ( \10851_11153 , RIfc448a0_5802, \8792_9091 );
and \U$2083 ( \10852_11154 , RIf141170_5200, \8794_9093 );
and \U$2084 ( \10853_11155 , RIfc7c9d0_6440, \8796_9095 );
and \U$2085 ( \10854_11156 , RIfea0098_8165, \8798_9097 );
and \U$2086 ( \10855_11157 , RIfc57e00_6022, \8800_9099 );
and \U$2087 ( \10856_11158 , RIf13f550_5180, \8802_9101 );
and \U$2088 ( \10857_11159 , RIfcd6e08_7467, \8804_9103 );
and \U$2089 ( \10858_11160 , RIee3d900_5159, \8806_9105 );
and \U$2090 ( \10859_11161 , RIfc8f6c0_6654, \8808_9107 );
and \U$2091 ( \10860_11162 , RIfce0048_7571, \8810_9109 );
and \U$2092 ( \10861_11163 , RIfca27e8_6871, \8812_9111 );
and \U$2093 ( \10862_11164 , RIe1742e8_2699, \8814_9113 );
and \U$2094 ( \10863_11165 , RIfc7c700_6438, \8816_9115 );
and \U$2095 ( \10864_11166 , RIfc8f990_6656, \8818_9117 );
and \U$2096 ( \10865_11167 , RIfce9828_7679, \8820_9119 );
and \U$2097 ( \10866_11168 , RIfc583a0_6026, \8822_9121 );
and \U$2098 ( \10867_11169 , RIf16cdc0_5698, \8824_9123 );
and \U$2099 ( \10868_11170 , RIe224670_4704, \8826_9125 );
and \U$2100 ( \10869_11171 , RIf16c118_5689, \8828_9127 );
and \U$2101 ( \10870_11172 , RIe221970_4672, \8830_9129 );
and \U$2102 ( \10871_11173 , RIfc58508_6027, \8832_9131 );
and \U$2103 ( \10872_11174 , RIe21ec70_4640, \8834_9133 );
and \U$2104 ( \10873_11175 , RIe219270_4576, \8836_9135 );
and \U$2105 ( \10874_11176 , RIe216570_4544, \8838_9137 );
and \U$2106 ( \10875_11177 , RIfc3ff08_5753, \8840_9139 );
and \U$2107 ( \10876_11178 , RIe213870_4512, \8842_9141 );
and \U$2108 ( \10877_11179 , RIf1696e8_5659, \8844_9143 );
and \U$2109 ( \10878_11180 , RIe210b70_4480, \8846_9145 );
and \U$2110 ( \10879_11181 , RIfc58940_6030, \8848_9147 );
and \U$2111 ( \10880_11182 , RIe20de70_4448, \8850_9149 );
and \U$2112 ( \10881_11183 , RIe20b170_4416, \8852_9151 );
and \U$2113 ( \10882_11184 , RIe208470_4384, \8854_9153 );
and \U$2114 ( \10883_11185 , RIfc8fc60_6658, \8856_9155 );
and \U$2115 ( \10884_11186 , RIfc97820_6746, \8858_9157 );
and \U$2116 ( \10885_11187 , RIe202ea8_4323, \8860_9159 );
and \U$2117 ( \10886_11188 , RIe201288_4303, \8862_9161 );
and \U$2118 ( \10887_11189 , RIfcc27c8_7235, \8864_9163 );
and \U$2119 ( \10888_11190 , RIfcdfee0_7570, \8866_9165 );
and \U$2120 ( \10889_11191 , RIfc44198_5797, \8868_9167 );
and \U$2121 ( \10890_11192 , RIfc58670_6028, \8870_9169 );
and \U$2122 ( \10891_11193 , RIf1608e0_5558, \8872_9171 );
and \U$2123 ( \10892_11194 , RIf15e9f0_5536, \8874_9173 );
and \U$2124 ( \10893_11195 , RIfe9ff30_8164, \8876_9175 );
and \U$2125 ( \10894_11196 , RIe1fc0f8_4245, \8878_9177 );
and \U$2126 ( \10895_11197 , RIfc7be90_6432, \8880_9179 );
and \U$2127 ( \10896_11198 , RIf15bb88_5503, \8882_9181 );
and \U$2128 ( \10897_11199 , RIfcd8cf8_7489, \8884_9183 );
and \U$2129 ( \10898_11200 , RIfcd8e60_7490, \8886_9185 );
or \U$2130 ( \10899_11201 , \10835_11137 , \10836_11138 , \10837_11139 , \10838_11140 , \10839_11141 , \10840_11142 , \10841_11143 , \10842_11144 , \10843_11145 , \10844_11146 , \10845_11147 , \10846_11148 , \10847_11149 , \10848_11150 , \10849_11151 , \10850_11152 , \10851_11153 , \10852_11154 , \10853_11155 , \10854_11156 , \10855_11157 , \10856_11158 , \10857_11159 , \10858_11160 , \10859_11161 , \10860_11162 , \10861_11163 , \10862_11164 , \10863_11165 , \10864_11166 , \10865_11167 , \10866_11168 , \10867_11169 , \10868_11170 , \10869_11171 , \10870_11172 , \10871_11173 , \10872_11174 , \10873_11175 , \10874_11176 , \10875_11177 , \10876_11178 , \10877_11179 , \10878_11180 , \10879_11181 , \10880_11182 , \10881_11183 , \10882_11184 , \10883_11185 , \10884_11186 , \10885_11187 , \10886_11188 , \10887_11189 , \10888_11190 , \10889_11191 , \10890_11192 , \10891_11193 , \10892_11194 , \10893_11195 , \10894_11196 , \10895_11197 , \10896_11198 , \10897_11199 , \10898_11200 );
and \U$2131 ( \10900_11202 , RIfca2d88_6875, \8889_9188 );
and \U$2132 ( \10901_11203 , RIfcbdea8_7183, \8891_9190 );
and \U$2133 ( \10902_11204 , RIfcb3a20_7066, \8893_9192 );
and \U$2134 ( \10903_11205 , RIe1fabe0_4230, \8895_9194 );
and \U$2135 ( \10904_11206 , RIfc90098_6661, \8897_9196 );
and \U$2136 ( \10905_11207 , RIfc90200_6662, \8899_9198 );
and \U$2137 ( \10906_11208 , RIfcd20b0_7412, \8901_9200 );
and \U$2138 ( \10907_11209 , RIe1f6158_4177, \8903_9202 );
and \U$2139 ( \10908_11210 , RIfc904d0_6664, \8905_9204 );
and \U$2140 ( \10909_11211 , RIfca2ef0_6876, \8907_9206 );
and \U$2141 ( \10910_11212 , RIfc97550_6744, \8909_9208 );
and \U$2142 ( \10911_11213 , RIe1f3e30_4152, \8911_9210 );
and \U$2143 ( \10912_11214 , RIfc59048_6035, \8913_9212 );
and \U$2144 ( \10913_11215 , RIfc907a0_6666, \8915_9214 );
and \U$2145 ( \10914_11216 , RIfc90638_6665, \8917_9216 );
and \U$2146 ( \10915_11217 , RIe1eeb38_4093, \8919_9218 );
and \U$2147 ( \10916_11218 , RIe1ec3d8_4065, \8921_9220 );
and \U$2148 ( \10917_11219 , RIe1e96d8_4033, \8923_9222 );
and \U$2149 ( \10918_11220 , RIe1e69d8_4001, \8925_9224 );
and \U$2150 ( \10919_11221 , RIe1e3cd8_3969, \8927_9226 );
and \U$2151 ( \10920_11222 , RIe1e0fd8_3937, \8929_9228 );
and \U$2152 ( \10921_11223 , RIe1de2d8_3905, \8931_9230 );
and \U$2153 ( \10922_11224 , RIe1db5d8_3873, \8933_9232 );
and \U$2154 ( \10923_11225 , RIe1d88d8_3841, \8935_9234 );
and \U$2155 ( \10924_11226 , RIe1d2ed8_3777, \8937_9236 );
and \U$2156 ( \10925_11227 , RIe1d01d8_3745, \8939_9238 );
and \U$2157 ( \10926_11228 , RIe1cd4d8_3713, \8941_9240 );
and \U$2158 ( \10927_11229 , RIe1ca7d8_3681, \8943_9242 );
and \U$2159 ( \10928_11230 , RIe1c7ad8_3649, \8945_9244 );
and \U$2160 ( \10929_11231 , RIe1c4dd8_3617, \8947_9246 );
and \U$2161 ( \10930_11232 , RIe1c20d8_3585, \8949_9248 );
and \U$2162 ( \10931_11233 , RIe1bf3d8_3553, \8951_9250 );
and \U$2163 ( \10932_11234 , RIfcc73b8_7289, \8953_9252 );
and \U$2164 ( \10933_11235 , RIfce3cc0_7614, \8955_9254 );
and \U$2165 ( \10934_11236 , RIe1b9e10_3492, \8957_9256 );
and \U$2166 ( \10935_11237 , RIe1b7c50_3468, \8959_9258 );
and \U$2167 ( \10936_11238 , RIfcd6f70_7468, \8961_9260 );
and \U$2168 ( \10937_11239 , RIf149e10_5300, \8963_9262 );
and \U$2169 ( \10938_11240 , RIe1b5a90_3444, \8965_9264 );
and \U$2170 ( \10939_11241 , RIfea0200_8166, \8967_9266 );
and \U$2171 ( \10940_11242 , RIfc90bd8_6669, \8969_9268 );
and \U$2172 ( \10941_11243 , RIfcdfd78_7569, \8971_9270 );
and \U$2173 ( \10942_11244 , RIe1b2ef8_3413, \8973_9272 );
and \U$2174 ( \10943_11245 , RIe1b15a8_3395, \8975_9274 );
and \U$2175 ( \10944_11246 , RIfc973e8_6743, \8977_9276 );
and \U$2176 ( \10945_11247 , RIfcc7520_7290, \8979_9278 );
and \U$2177 ( \10946_11248 , RIe1acdf0_3344, \8981_9280 );
and \U$2178 ( \10947_11249 , RIe1ab608_3327, \8983_9282 );
and \U$2179 ( \10948_11250 , RIe1a9718_3305, \8985_9284 );
and \U$2180 ( \10949_11251 , RIe1a6a18_3273, \8987_9286 );
and \U$2181 ( \10950_11252 , RIe1a3d18_3241, \8989_9288 );
and \U$2182 ( \10951_11253 , RIe1a1018_3209, \8991_9290 );
and \U$2183 ( \10952_11254 , RIe18d518_2985, \8993_9292 );
and \U$2184 ( \10953_11255 , RIe179a18_2761, \8995_9294 );
and \U$2185 ( \10954_11256 , RIe227370_4736, \8997_9296 );
and \U$2186 ( \10955_11257 , RIe21bf70_4608, \8999_9298 );
and \U$2187 ( \10956_11258 , RIe205770_4352, \9001_9300 );
and \U$2188 ( \10957_11259 , RIe1ff7d0_4284, \9003_9302 );
and \U$2189 ( \10958_11260 , RIe1f8b88_4207, \9005_9304 );
and \U$2190 ( \10959_11261 , RIe1f16d0_4124, \9007_9306 );
and \U$2191 ( \10960_11262 , RIe1d5bd8_3809, \9009_9308 );
and \U$2192 ( \10961_11263 , RIe1bc6d8_3521, \9011_9310 );
and \U$2193 ( \10962_11264 , RIe1af550_3372, \9013_9312 );
and \U$2194 ( \10963_11265 , RIe171b88_2671, \9015_9314 );
or \U$2195 ( \10964_11266 , \10900_11202 , \10901_11203 , \10902_11204 , \10903_11205 , \10904_11206 , \10905_11207 , \10906_11208 , \10907_11209 , \10908_11210 , \10909_11211 , \10910_11212 , \10911_11213 , \10912_11214 , \10913_11215 , \10914_11216 , \10915_11217 , \10916_11218 , \10917_11219 , \10918_11220 , \10919_11221 , \10920_11222 , \10921_11223 , \10922_11224 , \10923_11225 , \10924_11226 , \10925_11227 , \10926_11228 , \10927_11229 , \10928_11230 , \10929_11231 , \10930_11232 , \10931_11233 , \10932_11234 , \10933_11235 , \10934_11236 , \10935_11237 , \10936_11238 , \10937_11239 , \10938_11240 , \10939_11241 , \10940_11242 , \10941_11243 , \10942_11244 , \10943_11245 , \10944_11246 , \10945_11247 , \10946_11248 , \10947_11249 , \10948_11250 , \10949_11251 , \10950_11252 , \10951_11253 , \10952_11254 , \10953_11255 , \10954_11256 , \10955_11257 , \10956_11258 , \10957_11259 , \10958_11260 , \10959_11261 , \10960_11262 , \10961_11263 , \10962_11264 , \10963_11265 );
or \U$2196 ( \10965_11267 , \10899_11201 , \10964_11266 );
_DC \g657e/U$1 ( \10966 , \10965_11267 , \9024_9323 );
and g657f_GF_PartitionCandidate( \10967_11269_nG657f , \10834 , \10966 );
buf \U$2197 ( \10968_11270 , \10967_11269_nG657f );
and \U$2198 ( \10969_11271 , \10968_11270 , \10389_10691 );
nor \U$2199 ( \10970_11272 , \10702_11004 , \10969_11271 );
xnor \U$2200 ( \10971_11273 , \10970_11272 , \10678_10980 );
_DC \g46ec/U$1 ( \10972 , \10833_11135 , \9298_9597 );
_DC \g4770/U$1 ( \10973 , \10965_11267 , \9024_9323 );
xor g4771_GF_PartitionCandidate( \10974_11276_nG4771 , \10972 , \10973 );
buf \U$2201 ( \10975_11277 , \10974_11276_nG4771 );
xor \U$2202 ( \10976_11278 , \10975_11277 , \10678_10980 );
and \U$2203 ( \10977_11279 , \10385_10687 , \10976_11278 );
xor \U$2204 ( \10978_11280 , \10971_11273 , \10977_11279 );
and \U$2205 ( \10979_11281 , \10689_10991 , \10691_10993 );
xor \U$2206 ( \10980_11282 , \10978_11280 , \10979_11281 );
buf g9c08_GF_PartitionCandidate( \10981_11283_nG9c08 , \10980_11282 );
and \U$2207 ( \10982_11284 , \10402_10704 , \10981_11283_nG9c08 );
or \U$2208 ( \10983_11285 , \10701_11003 , \10982_11284 );
xor \U$2209 ( \10984_11286 , \10399_10703 , \10983_11285 );
buf \U$2210 ( \10985_11287 , \10984_11286 );
buf \U$2212 ( \10986_11288 , \10985_11287 );
xor \U$2213 ( \10987_11289 , \10700_11002 , \10986_11288 );
and \U$2214 ( \10988_11290 , \10398_10700 , \10987_11289 );
and \U$2215 ( \10989_11291 , \10700_11002 , \10986_11288 );
buf \U$2216 ( \10990_11292 , \10989_11291 );
and \U$2217 ( \10991_11293 , \10118_10417 , \10395_10697 );
buf \U$2218 ( \10992_11294 , \10991_11293 );
buf \U$2220 ( \10993_11295 , \10992_11294 );
not \U$1357 ( \10994_10419 , \10119_10418 );
xor \U$1358 ( \10995_10420 , \10110_10409_nG444e , \10113_10412_nG4451 );
and \U$1359 ( \10996_10421 , \10994_10419 , \10995_10420 );
and \U$2221 ( \10997_11296 , \10996_10421 , \10392_10694_nG9c0e );
and \U$2222 ( \10998_11297 , \10119_10418 , \10693_10995_nG9c0b );
or \U$2223 ( \10999_11298 , \10997_11296 , \10998_11297 );
xor \U$2224 ( \11000_11299 , \10118_10417 , \10999_11298 );
buf \U$2225 ( \11001_11300 , \11000_11299 );
buf \U$2227 ( \11002_11301 , \11001_11300 );
xor \U$2228 ( \11003_11302 , \10993_11295 , \11002_11301 );
buf \U$2229 ( \11004_11303 , \11003_11302 );
xor \U$2230 ( \11005_11304 , \10990_11292 , \11004_11303 );
and \U$2231 ( \11006_11305 , \10411_10707 , \10981_11283_nG9c08 );
and \U$2232 ( \11007_11306 , RIdec64b8_720, \9034_9333 );
and \U$2233 ( \11008_11307 , RIdec37b8_688, \9036_9335 );
and \U$2234 ( \11009_11308 , RIfc8daa0_6634, \9038_9337 );
and \U$2235 ( \11010_11309 , RIdec0ab8_656, \9040_9339 );
and \U$2236 ( \11011_11310 , RIfc56348_6003, \9042_9341 );
and \U$2237 ( \11012_11311 , RIdebddb8_624, \9044_9343 );
and \U$2238 ( \11013_11312 , RIdebb0b8_592, \9046_9345 );
and \U$2239 ( \11014_11313 , RIdeb83b8_560, \9048_9347 );
and \U$2240 ( \11015_11314 , RIfc98798_6757, \9050_9349 );
and \U$2241 ( \11016_11315 , RIdeb29b8_496, \9052_9351 );
and \U$2242 ( \11017_11316 , RIfcbd098_7173, \9054_9353 );
and \U$2243 ( \11018_11317 , RIdeafcb8_464, \9056_9355 );
and \U$2244 ( \11019_11318 , RIfc8dc08_6635, \9058_9357 );
and \U$2245 ( \11020_11319 , RIdeacb80_432, \9060_9359 );
and \U$2246 ( \11021_11320 , RIdea6280_400, \9062_9361 );
and \U$2247 ( \11022_11321 , RIde9f980_368, \9064_9363 );
and \U$2248 ( \11023_11322 , RIfcd6868_7463, \9066_9365 );
and \U$2249 ( \11024_11323 , RIfc8ded8_6637, \9068_9367 );
and \U$2250 ( \11025_11324 , RIfc7dd80_6454, \9070_9369 );
and \U$2251 ( \11026_11325 , RIfc56618_6005, \9072_9371 );
and \U$2252 ( \11027_11326 , RIde92e10_306, \9074_9373 );
and \U$2253 ( \11028_11327 , RIde8f300_288, \9076_9375 );
and \U$2254 ( \11029_11328 , RIde8b160_268, \9078_9377 );
and \U$2255 ( \11030_11329 , RIde86fc0_248, \9080_9379 );
and \U$2256 ( \11031_11330 , RIde82ad8_227, \9082_9381 );
and \U$2257 ( \11032_11331 , RIfc8e040_6638, \9084_9383 );
and \U$2258 ( \11033_11332 , RIfcd96d0_7496, \9086_9385 );
and \U$2259 ( \11034_11333 , RIfca1e10_6864, \9088_9387 );
and \U$2260 ( \11035_11334 , RIfcbd200_7174, \9090_9389 );
and \U$2261 ( \11036_11335 , RIe16c5c0_2610, \9092_9391 );
and \U$2262 ( \11037_11336 , RIe16a298_2585, \9094_9393 );
and \U$2263 ( \11038_11337 , RIe168ab0_2568, \9096_9395 );
and \U$2264 ( \11039_11338 , RIe1664b8_2541, \9098_9397 );
and \U$2265 ( \11040_11339 , RIe1637b8_2509, \9100_9399 );
and \U$2266 ( \11041_11340 , RIee37f00_5095, \9102_9401 );
and \U$2267 ( \11042_11341 , RIe160ab8_2477, \9104_9403 );
and \U$2268 ( \11043_11342 , RIfc8ea18_6645, \9106_9405 );
and \U$2269 ( \11044_11343 , RIe15ddb8_2445, \9108_9407 );
and \U$2270 ( \11045_11344 , RIe1583b8_2381, \9110_9409 );
and \U$2271 ( \11046_11345 , RIe1556b8_2349, \9112_9411 );
and \U$2272 ( \11047_11346 , RIfe9f828_8159, \9114_9413 );
and \U$2273 ( \11048_11347 , RIe1529b8_2317, \9116_9415 );
and \U$2274 ( \11049_11348 , RIfe9f990_8160, \9118_9417 );
and \U$2275 ( \11050_11349 , RIe14fcb8_2285, \9120_9419 );
and \U$2276 ( \11051_11350 , RIfcbd368_7175, \9122_9421 );
and \U$2277 ( \11052_11351 , RIe14cfb8_2253, \9124_9423 );
and \U$2278 ( \11053_11352 , RIe14a2b8_2221, \9126_9425 );
and \U$2279 ( \11054_11353 , RIe1475b8_2189, \9128_9427 );
and \U$2280 ( \11055_11354 , RIfc8ee50_6648, \9130_9429 );
and \U$2281 ( \11056_11355 , RIfc45278_5809, \9132_9431 );
and \U$2282 ( \11057_11356 , RIfc98360_6754, \9134_9433 );
and \U$2283 ( \11058_11357 , RIfca2248_6867, \9136_9435 );
and \U$2284 ( \11059_11358 , RIe141d20_2126, \9138_9437 );
and \U$2285 ( \11060_11359 , RIe13f9f8_2101, \9140_9439 );
and \U$2286 ( \11061_11360 , RIdf3d900_2077, \9142_9441 );
and \U$2287 ( \11062_11361 , RIdf3b470_2051, \9144_9443 );
and \U$2288 ( \11063_11362 , RIfcd6ca0_7466, \9146_9445 );
and \U$2289 ( \11064_11363 , RIee2ff08_5004, \9148_9447 );
and \U$2290 ( \11065_11364 , RIfc8ece8_6647, \9150_9449 );
and \U$2291 ( \11066_11365 , RIee2dd48_4980, \9152_9451 );
and \U$2292 ( \11067_11366 , RIdf36718_1996, \9154_9453 );
and \U$2293 ( \11068_11367 , RIdf34120_1969, \9156_9455 );
and \U$2294 ( \11069_11368 , RIdf31f60_1945, \9158_9457 );
and \U$2295 ( \11070_11369 , RIfe9f6c0_8158, \9160_9459 );
or \U$2296 ( \11071_11370 , \11007_11306 , \11008_11307 , \11009_11308 , \11010_11309 , \11011_11310 , \11012_11311 , \11013_11312 , \11014_11313 , \11015_11314 , \11016_11315 , \11017_11316 , \11018_11317 , \11019_11318 , \11020_11319 , \11021_11320 , \11022_11321 , \11023_11322 , \11024_11323 , \11025_11324 , \11026_11325 , \11027_11326 , \11028_11327 , \11029_11328 , \11030_11329 , \11031_11330 , \11032_11331 , \11033_11332 , \11034_11333 , \11035_11334 , \11036_11335 , \11037_11336 , \11038_11337 , \11039_11338 , \11040_11339 , \11041_11340 , \11042_11341 , \11043_11342 , \11044_11343 , \11045_11344 , \11046_11345 , \11047_11346 , \11048_11347 , \11049_11348 , \11050_11349 , \11051_11350 , \11052_11351 , \11053_11352 , \11054_11353 , \11055_11354 , \11056_11355 , \11057_11356 , \11058_11357 , \11059_11358 , \11060_11359 , \11061_11360 , \11062_11361 , \11063_11362 , \11064_11363 , \11065_11364 , \11066_11365 , \11067_11366 , \11068_11367 , \11069_11368 , \11070_11369 );
and \U$2297 ( \11072_11371 , RIfcb4560_7074, \9163_9462 );
and \U$2298 ( \11073_11372 , RIfc45db8_5817, \9165_9464 );
and \U$2299 ( \11074_11373 , RIfc8e1a8_6639, \9167_9466 );
and \U$2300 ( \11075_11374 , RIfc7d678_6449, \9169_9468 );
and \U$2301 ( \11076_11375 , RIdf2aee0_1865, \9171_9470 );
and \U$2302 ( \11077_11376 , RIdf28ff0_1843, \9173_9472 );
and \U$2303 ( \11078_11377 , RIdf26e30_1819, \9175_9474 );
and \U$2304 ( \11079_11378 , RIdf25378_1800, \9177_9476 );
and \U$2305 ( \11080_11379 , RIfcb43f8_7073, \9179_9478 );
and \U$2306 ( \11081_11380 , RIfc8e748_6643, \9181_9480 );
and \U$2307 ( \11082_11381 , RIdf23488_1778, \9183_9482 );
and \U$2308 ( \11083_11382 , RIfcc2c00_7238, \9185_9484 );
and \U$2309 ( \11084_11383 , RIdf21e08_1762, \9187_9486 );
and \U$2310 ( \11085_11384 , RIdf20788_1746, \9189_9488 );
and \U$2311 ( \11086_11385 , RIdf1b760_1689, \9191_9490 );
and \U$2312 ( \11087_11386 , RIdf1a248_1674, \9193_9492 );
and \U$2313 ( \11088_11387 , RIdf18088_1650, \9195_9494 );
and \U$2314 ( \11089_11388 , RIdf15388_1618, \9197_9496 );
and \U$2315 ( \11090_11389 , RIdf12688_1586, \9199_9498 );
and \U$2316 ( \11091_11390 , RIdf0f988_1554, \9201_9500 );
and \U$2317 ( \11092_11391 , RIdf0cc88_1522, \9203_9502 );
and \U$2318 ( \11093_11392 , RIdf09f88_1490, \9205_9504 );
and \U$2319 ( \11094_11393 , RIdf07288_1458, \9207_9506 );
and \U$2320 ( \11095_11394 , RIdf04588_1426, \9209_9508 );
and \U$2321 ( \11096_11395 , RIdefeb88_1362, \9211_9510 );
and \U$2322 ( \11097_11396 , RIdefbe88_1330, \9213_9512 );
and \U$2323 ( \11098_11397 , RIdef9188_1298, \9215_9514 );
and \U$2324 ( \11099_11398 , RIdef6488_1266, \9217_9516 );
and \U$2325 ( \11100_11399 , RIdef3788_1234, \9219_9518 );
and \U$2326 ( \11101_11400 , RIdef0a88_1202, \9221_9520 );
and \U$2327 ( \11102_11401 , RIdeedd88_1170, \9223_9522 );
and \U$2328 ( \11103_11402 , RIdeeb088_1138, \9225_9524 );
and \U$2329 ( \11104_11403 , RIfc8efb8_6649, \9227_9526 );
and \U$2330 ( \11105_11404 , RIfc44e40_5806, \9229_9528 );
and \U$2331 ( \11106_11405 , RIfc57860_6018, \9231_9530 );
and \U$2332 ( \11107_11406 , RIfca23b0_6868, \9233_9532 );
and \U$2333 ( \11108_11407 , RIfe9faf8_8161, \9235_9534 );
and \U$2334 ( \11109_11408 , RIdee3900_1053, \9237_9536 );
and \U$2335 ( \11110_11409 , RIdee1740_1029, \9239_9538 );
and \U$2336 ( \11111_11410 , RIdedf6e8_1006, \9241_9540 );
and \U$2337 ( \11112_11411 , RIfcbd4d0_7176, \9243_9542 );
and \U$2338 ( \11113_11412 , RIee22678_4850, \9245_9544 );
and \U$2339 ( \11114_11413 , RIfc98090_6752, \9247_9546 );
and \U$2340 ( \11115_11414 , RIee21598_4838, \9249_9548 );
and \U$2341 ( \11116_11415 , RIfe9fc60_8162, \9251_9550 );
and \U$2342 ( \11117_11416 , RIded80c8_922, \9253_9552 );
and \U$2343 ( \11118_11417 , RIfe9fdc8_8163, \9255_9554 );
and \U$2344 ( \11119_11418 , RIded3be0_873, \9257_9556 );
and \U$2345 ( \11120_11419 , RIded18b8_848, \9259_9558 );
and \U$2346 ( \11121_11420 , RIdecebb8_816, \9261_9560 );
and \U$2347 ( \11122_11421 , RIdecbeb8_784, \9263_9562 );
and \U$2348 ( \11123_11422 , RIdec91b8_752, \9265_9564 );
and \U$2349 ( \11124_11423 , RIdeb56b8_528, \9267_9566 );
and \U$2350 ( \11125_11424 , RIde99080_336, \9269_9568 );
and \U$2351 ( \11126_11425 , RIe16f2c0_2642, \9271_9570 );
and \U$2352 ( \11127_11426 , RIe15b0b8_2413, \9273_9572 );
and \U$2353 ( \11128_11427 , RIe1448b8_2157, \9275_9574 );
and \U$2354 ( \11129_11428 , RIdf392b0_2027, \9277_9576 );
and \U$2355 ( \11130_11429 , RIdf2d910_1895, \9279_9578 );
and \U$2356 ( \11131_11430 , RIdf1e190_1719, \9281_9580 );
and \U$2357 ( \11132_11431 , RIdf01888_1394, \9283_9582 );
and \U$2358 ( \11133_11432 , RIdee8388_1106, \9285_9584 );
and \U$2359 ( \11134_11433 , RIdedd0f0_979, \9287_9586 );
and \U$2360 ( \11135_11434 , RIde7efc8_209, \9289_9588 );
or \U$2361 ( \11136_11435 , \11072_11371 , \11073_11372 , \11074_11373 , \11075_11374 , \11076_11375 , \11077_11376 , \11078_11377 , \11079_11378 , \11080_11379 , \11081_11380 , \11082_11381 , \11083_11382 , \11084_11383 , \11085_11384 , \11086_11385 , \11087_11386 , \11088_11387 , \11089_11388 , \11090_11389 , \11091_11390 , \11092_11391 , \11093_11392 , \11094_11393 , \11095_11394 , \11096_11395 , \11097_11396 , \11098_11397 , \11099_11398 , \11100_11399 , \11101_11400 , \11102_11401 , \11103_11402 , \11104_11403 , \11105_11404 , \11106_11405 , \11107_11406 , \11108_11407 , \11109_11408 , \11110_11409 , \11111_11410 , \11112_11411 , \11113_11412 , \11114_11413 , \11115_11414 , \11116_11415 , \11117_11416 , \11118_11417 , \11119_11418 , \11120_11419 , \11121_11420 , \11122_11421 , \11123_11422 , \11124_11423 , \11125_11424 , \11126_11425 , \11127_11426 , \11128_11427 , \11129_11428 , \11130_11429 , \11131_11430 , \11132_11431 , \11133_11432 , \11134_11433 , \11135_11434 );
or \U$2362 ( \11137_11436 , \11071_11370 , \11136_11435 );
_DC \g47f5/U$1 ( \11138 , \11137_11436 , \9298_9597 );
and \U$2363 ( \11139_11438 , RIe19e750_3180, \8760_9059 );
and \U$2364 ( \11140_11439 , RIe19ba50_3148, \8762_9061 );
and \U$2365 ( \11141_11440 , RIfc479d8_5837, \8764_9063 );
and \U$2366 ( \11142_11441 , RIe198d50_3116, \8766_9065 );
and \U$2367 ( \11143_11442 , RIfe9f558_8157, \8768_9067 );
and \U$2368 ( \11144_11443 , RIe196050_3084, \8770_9069 );
and \U$2369 ( \11145_11444 , RIe193350_3052, \8772_9071 );
and \U$2370 ( \11146_11445 , RIe190650_3020, \8774_9073 );
and \U$2371 ( \11147_11446 , RIe18ac50_2956, \8776_9075 );
and \U$2372 ( \11148_11447 , RIe187f50_2924, \8778_9077 );
and \U$2373 ( \11149_11448 , RIfc47870_5836, \8780_9079 );
and \U$2374 ( \11150_11449 , RIe185250_2892, \8782_9081 );
and \U$2375 ( \11151_11450 , RIf142ef8_5221, \8784_9083 );
and \U$2376 ( \11152_11451 , RIe182550_2860, \8786_9085 );
and \U$2377 ( \11153_11452 , RIe17f850_2828, \8788_9087 );
and \U$2378 ( \11154_11453 , RIe17cb50_2796, \8790_9089 );
and \U$2379 ( \11155_11454 , RIfcb5208_7083, \8792_9091 );
and \U$2380 ( \11156_11455 , RIfcbc6c0_7166, \8794_9093 );
and \U$2381 ( \11157_11456 , RIe177588_2735, \8796_9095 );
and \U$2382 ( \11158_11457 , RIe176610_2724, \8798_9097 );
and \U$2383 ( \11159_11458 , RIf13fdc0_5186, \8800_9099 );
and \U$2384 ( \11160_11459 , RIfe9f3f0_8156, \8802_9101 );
and \U$2385 ( \11161_11460 , RIfce40f8_7617, \8804_9103 );
and \U$2386 ( \11162_11461 , RIfc47708_5835, \8806_9105 );
and \U$2387 ( \11163_11462 , RIfc47438_5833, \8808_9107 );
and \U$2388 ( \11164_11463 , RIfca15a0_6858, \8810_9109 );
and \U$2389 ( \11165_11464 , RIfc99170_6764, \8812_9111 );
and \U$2390 ( \11166_11465 , RIe1745b8_2701, \8814_9113 );
and \U$2391 ( \11167_11466 , RIfc8cc90_6624, \8816_9115 );
and \U$2392 ( \11168_11467 , RIfc556a0_5994, \8818_9117 );
and \U$2393 ( \11169_11468 , RIfc7ee60_6466, \8820_9119 );
and \U$2394 ( \11170_11469 , RIfce8e50_7672, \8822_9121 );
and \U$2395 ( \11171_11470 , RIfe9f288_8155, \8824_9123 );
and \U$2396 ( \11172_11471 , RIe224aa8_4707, \8826_9125 );
and \U$2397 ( \11173_11472 , RIfc55808_5995, \8828_9127 );
and \U$2398 ( \11174_11473 , RIe221da8_4675, \8830_9129 );
and \U$2399 ( \11175_11474 , RIfcb50a0_7082, \8832_9131 );
and \U$2400 ( \11176_11475 , RIe21f0a8_4643, \8834_9133 );
and \U$2401 ( \11177_11476 , RIe2196a8_4579, \8836_9135 );
and \U$2402 ( \11178_11477 , RIe2169a8_4547, \8838_9137 );
and \U$2403 ( \11179_11478 , RIfcbc828_7167, \8840_9139 );
and \U$2404 ( \11180_11479 , RIe213ca8_4515, \8842_9141 );
and \U$2405 ( \11181_11480 , RIfc47000_5830, \8844_9143 );
and \U$2406 ( \11182_11481 , RIe210fa8_4483, \8846_9145 );
and \U$2407 ( \11183_11482 , RIfcbc990_7168, \8848_9147 );
and \U$2408 ( \11184_11483 , RIe20e2a8_4451, \8850_9149 );
and \U$2409 ( \11185_11484 , RIe20b5a8_4419, \8852_9151 );
and \U$2410 ( \11186_11485 , RIe2088a8_4387, \8854_9153 );
and \U$2411 ( \11187_11486 , RIfc46bc8_5827, \8856_9155 );
and \U$2412 ( \11188_11487 , RIfcd6598_7461, \8858_9157 );
and \U$2413 ( \11189_11488 , RIe2032e0_4326, \8860_9159 );
and \U$2414 ( \11190_11489 , RIe2016c0_4306, \8862_9161 );
and \U$2415 ( \11191_11490 , RIfc98ea0_6762, \8864_9163 );
and \U$2416 ( \11192_11491 , RIfc7eb90_6464, \8866_9165 );
and \U$2417 ( \11193_11492 , RIfce0318_7573, \8868_9167 );
and \U$2418 ( \11194_11493 , RIfcbcaf8_7169, \8870_9169 );
and \U$2419 ( \11195_11494 , RIfc8cf60_6626, \8872_9171 );
and \U$2420 ( \11196_11495 , RIfcb4dd0_7080, \8874_9173 );
and \U$2421 ( \11197_11496 , RIe1fd340_4258, \8876_9175 );
and \U$2422 ( \11198_11497 , RIe1fc260_4246, \8878_9177 );
and \U$2423 ( \11199_11498 , RIf15cf38_5517, \8880_9179 );
and \U$2424 ( \11200_11499 , RIfe9f120_8154, \8882_9181 );
and \U$2425 ( \11201_11500 , RIfc7ea28_6463, \8884_9183 );
and \U$2426 ( \11202_11501 , RIfc8d0c8_6627, \8886_9185 );
or \U$2427 ( \11203_11502 , \11139_11438 , \11140_11439 , \11141_11440 , \11142_11441 , \11143_11442 , \11144_11443 , \11145_11444 , \11146_11445 , \11147_11446 , \11148_11447 , \11149_11448 , \11150_11449 , \11151_11450 , \11152_11451 , \11153_11452 , \11154_11453 , \11155_11454 , \11156_11455 , \11157_11456 , \11158_11457 , \11159_11458 , \11160_11459 , \11161_11460 , \11162_11461 , \11163_11462 , \11164_11463 , \11165_11464 , \11166_11465 , \11167_11466 , \11168_11467 , \11169_11468 , \11170_11469 , \11171_11470 , \11172_11471 , \11173_11472 , \11174_11473 , \11175_11474 , \11176_11475 , \11177_11476 , \11178_11477 , \11179_11478 , \11180_11479 , \11181_11480 , \11182_11481 , \11183_11482 , \11184_11483 , \11185_11484 , \11186_11485 , \11187_11486 , \11188_11487 , \11189_11488 , \11190_11489 , \11191_11490 , \11192_11491 , \11193_11492 , \11194_11493 , \11195_11494 , \11196_11495 , \11197_11496 , \11198_11497 , \11199_11498 , \11200_11499 , \11201_11500 , \11202_11501 );
and \U$2428 ( \11204_11503 , RIfcbcc60_7170, \8889_9188 );
and \U$2429 ( \11205_11504 , RIfc98bd0_6760, \8891_9190 );
and \U$2430 ( \11206_11505 , RIfce2d48_7603, \8893_9192 );
and \U$2431 ( \11207_11506 , RIe1fb018_4233, \8895_9194 );
and \U$2432 ( \11208_11507 , RIfc55f10_6000, \8897_9196 );
and \U$2433 ( \11209_11508 , RIfc7e8c0_6462, \8899_9198 );
and \U$2434 ( \11210_11509 , RIfc8d230_6628, \8901_9200 );
and \U$2435 ( \11211_11510 , RIe1f6590_4180, \8903_9202 );
and \U$2436 ( \11212_11511 , RIfce58e0_7634, \8905_9204 );
and \U$2437 ( \11213_11512 , RIfc468f8_5825, \8907_9206 );
and \U$2438 ( \11214_11513 , RIfcc2ed0_7240, \8909_9208 );
and \U$2439 ( \11215_11514 , RIe1f4100_4154, \8911_9210 );
and \U$2440 ( \11216_11515 , RIfceedf0_7740, \8913_9212 );
and \U$2441 ( \11217_11516 , RIfc8d398_6629, \8915_9214 );
and \U$2442 ( \11218_11517 , RIfc8d500_6630, \8917_9216 );
and \U$2443 ( \11219_11518 , RIe1eef70_4096, \8919_9218 );
and \U$2444 ( \11220_11519 , RIe1ec810_4068, \8921_9220 );
and \U$2445 ( \11221_11520 , RIe1e9b10_4036, \8923_9222 );
and \U$2446 ( \11222_11521 , RIe1e6e10_4004, \8925_9224 );
and \U$2447 ( \11223_11522 , RIe1e4110_3972, \8927_9226 );
and \U$2448 ( \11224_11523 , RIe1e1410_3940, \8929_9228 );
and \U$2449 ( \11225_11524 , RIe1de710_3908, \8931_9230 );
and \U$2450 ( \11226_11525 , RIe1dba10_3876, \8933_9232 );
and \U$2451 ( \11227_11526 , RIe1d8d10_3844, \8935_9234 );
and \U$2452 ( \11228_11527 , RIe1d3310_3780, \8937_9236 );
and \U$2453 ( \11229_11528 , RIe1d0610_3748, \8939_9238 );
and \U$2454 ( \11230_11529 , RIe1cd910_3716, \8941_9240 );
and \U$2455 ( \11231_11530 , RIe1cac10_3684, \8943_9242 );
and \U$2456 ( \11232_11531 , RIe1c7f10_3652, \8945_9244 );
and \U$2457 ( \11233_11532 , RIe1c5210_3620, \8947_9246 );
and \U$2458 ( \11234_11533 , RIe1c2510_3588, \8949_9248 );
and \U$2459 ( \11235_11534 , RIe1bf810_3556, \8951_9250 );
and \U$2460 ( \11236_11535 , RIf14d0b0_5336, \8953_9252 );
and \U$2461 ( \11237_11536 , RIfe9efb8_8153, \8955_9254 );
and \U$2462 ( \11238_11537 , RIe1ba248_3495, \8957_9256 );
and \U$2463 ( \11239_11538 , RIe1b8088_3471, \8959_9258 );
and \U$2464 ( \11240_11539 , RIfec4dd0_8360, \8961_9260 );
and \U$2465 ( \11241_11540 , RIfec50a0_8362, \8963_9262 );
and \U$2466 ( \11242_11541 , RIe1b5ec8_3447, \8965_9264 );
and \U$2467 ( \11243_11542 , RIe1b46e0_3430, \8967_9266 );
and \U$2468 ( \11244_11543 , RIfcb4998_7077, \8969_9268 );
and \U$2469 ( \11245_11544 , RIfcb4c68_7079, \8971_9270 );
and \U$2470 ( \11246_11545 , RIfec5370_8364, \8973_9272 );
and \U$2471 ( \11247_11546 , RIfe9ee50_8152, \8975_9274 );
and \U$2472 ( \11248_11547 , RIfcbcdc8_7171, \8977_9276 );
and \U$2473 ( \11249_11548 , RIfc46358_5821, \8979_9278 );
and \U$2474 ( \11250_11549 , RIfec5208_8363, \8981_9280 );
and \U$2475 ( \11251_11550 , RIfec4f38_8361, \8983_9282 );
and \U$2476 ( \11252_11551 , RIe1a9b50_3308, \8985_9284 );
and \U$2477 ( \11253_11552 , RIe1a6e50_3276, \8987_9286 );
and \U$2478 ( \11254_11553 , RIe1a4150_3244, \8989_9288 );
and \U$2479 ( \11255_11554 , RIe1a1450_3212, \8991_9290 );
and \U$2480 ( \11256_11555 , RIe18d950_2988, \8993_9292 );
and \U$2481 ( \11257_11556 , RIe179e50_2764, \8995_9294 );
and \U$2482 ( \11258_11557 , RIe2277a8_4739, \8997_9296 );
and \U$2483 ( \11259_11558 , RIe21c3a8_4611, \8999_9298 );
and \U$2484 ( \11260_11559 , RIe205ba8_4355, \9001_9300 );
and \U$2485 ( \11261_11560 , RIe1ffc08_4287, \9003_9302 );
and \U$2486 ( \11262_11561 , RIe1f8fc0_4210, \9005_9304 );
and \U$2487 ( \11263_11562 , RIe1f1b08_4127, \9007_9306 );
and \U$2488 ( \11264_11563 , RIe1d6010_3812, \9009_9308 );
and \U$2489 ( \11265_11564 , RIe1bcb10_3524, \9011_9310 );
and \U$2490 ( \11266_11565 , RIe1af988_3375, \9013_9312 );
and \U$2491 ( \11267_11566 , RIe171fc0_2674, \9015_9314 );
or \U$2492 ( \11268_11567 , \11204_11503 , \11205_11504 , \11206_11505 , \11207_11506 , \11208_11507 , \11209_11508 , \11210_11509 , \11211_11510 , \11212_11511 , \11213_11512 , \11214_11513 , \11215_11514 , \11216_11515 , \11217_11516 , \11218_11517 , \11219_11518 , \11220_11519 , \11221_11520 , \11222_11521 , \11223_11522 , \11224_11523 , \11225_11524 , \11226_11525 , \11227_11526 , \11228_11527 , \11229_11528 , \11230_11529 , \11231_11530 , \11232_11531 , \11233_11532 , \11234_11533 , \11235_11534 , \11236_11535 , \11237_11536 , \11238_11537 , \11239_11538 , \11240_11539 , \11241_11540 , \11242_11541 , \11243_11542 , \11244_11543 , \11245_11544 , \11246_11545 , \11247_11546 , \11248_11547 , \11249_11548 , \11250_11549 , \11251_11550 , \11252_11551 , \11253_11552 , \11254_11553 , \11255_11554 , \11256_11555 , \11257_11556 , \11258_11557 , \11259_11558 , \11260_11559 , \11261_11560 , \11262_11561 , \11263_11562 , \11264_11563 , \11265_11564 , \11266_11565 , \11267_11566 );
or \U$2493 ( \11269_11568 , \11203_11502 , \11268_11567 );
_DC \g4879/U$1 ( \11270 , \11269_11568 , \9024_9323 );
xor g487a_GF_PartitionCandidate( \11271_11570_nG487a , \11138 , \11270 );
buf \U$2494 ( \11272_11571 , \11271_11570_nG487a );
xor \U$2495 ( \11273_11572 , \11272_11571 , \10975_11277 );
not \U$2496 ( \11274_11573 , \10976_11278 );
and \U$2497 ( \11275_11574 , \11273_11572 , \11274_11573 );
and \U$2498 ( \11276_11575 , \10385_10687 , \11275_11574 );
and \U$2499 ( \11277_11576 , \10686_10988 , \10976_11278 );
nor \U$2500 ( \11278_11577 , \11276_11575 , \11277_11576 );
and \U$2501 ( \11279_11578 , \10975_11277 , \10678_10980 );
not \U$2502 ( \11280_11579 , \11279_11578 );
and \U$2503 ( \11281_11580 , \11272_11571 , \11280_11579 );
xnor \U$2504 ( \11282_11581 , \11278_11577 , \11281_11580 );
and \U$2505 ( \11283_11582 , \10968_11270 , \10681_10983 );
_DC \g6580/U$1 ( \11284 , \11137_11436 , \9298_9597 );
_DC \g6581/U$1 ( \11285 , \11269_11568 , \9024_9323 );
and g6582_GF_PartitionCandidate( \11286_11585_nG6582 , \11284 , \11285 );
buf \U$2506 ( \11287_11586 , \11286_11585_nG6582 );
and \U$2507 ( \11288_11587 , \11287_11586 , \10389_10691 );
nor \U$2508 ( \11289_11588 , \11283_11582 , \11288_11587 );
xnor \U$2509 ( \11290_11589 , \11289_11588 , \10678_10980 );
not \U$2510 ( \11291_11590 , \10977_11279 );
and \U$2511 ( \11292_11591 , \11291_11590 , \11281_11580 );
xor \U$2512 ( \11293_11592 , \11290_11589 , \11292_11591 );
xor \U$2513 ( \11294_11593 , \11282_11581 , \11293_11592 );
and \U$2514 ( \11295_11594 , \10971_11273 , \10977_11279 );
and \U$2515 ( \11296_11595 , \10978_11280 , \10979_11281 );
or \U$2516 ( \11297_11596 , \11295_11594 , \11296_11595 );
xor \U$2517 ( \11298_11597 , \11294_11593 , \11297_11596 );
buf g9c05_GF_PartitionCandidate( \11299_11598_nG9c05 , \11298_11597 );
and \U$2518 ( \11300_11599 , \10402_10704 , \11299_11598_nG9c05 );
or \U$2519 ( \11301_11600 , \11006_11305 , \11300_11599 );
xor \U$2520 ( \11302_11601 , \10399_10703 , \11301_11600 );
buf \U$2521 ( \11303_11602 , \11302_11601 );
buf \U$2523 ( \11304_11603 , \11303_11602 );
xor \U$2524 ( \11305_11604 , \11005_11304 , \11304_11603 );
and \U$2525 ( \11306_11605 , \10988_11290 , \11305_11604 );
and \U$2526 ( \11307_11606 , RIdec6788_722, \8760_9059 );
and \U$2527 ( \11308_11607 , RIdec3a88_690, \8762_9061 );
and \U$2528 ( \11309_11608 , RIee20788_4828, \8764_9063 );
and \U$2529 ( \11310_11609 , RIdec0d88_658, \8766_9065 );
and \U$2530 ( \11311_11610 , RIee1f810_4817, \8768_9067 );
and \U$2531 ( \11312_11611 , RIdebe088_626, \8770_9069 );
and \U$2532 ( \11313_11612 , RIdebb388_594, \8772_9071 );
and \U$2533 ( \11314_11613 , RIdeb8688_562, \8774_9073 );
and \U$2534 ( \11315_11614 , RIfc9b1c8_6787, \8776_9075 );
and \U$2535 ( \11316_11615 , RIdeb2c88_498, \8778_9077 );
and \U$2536 ( \11317_11616 , RIfce1f38_7593, \8780_9079 );
and \U$2537 ( \11318_11617 , RIdeaff88_466, \8782_9081 );
and \U$2538 ( \11319_11618 , RIfc892e8_6583, \8784_9083 );
and \U$2539 ( \11320_11619 , RIdead210_434, \8786_9085 );
and \U$2540 ( \11321_11620 , RIdea6910_402, \8788_9087 );
and \U$2541 ( \11322_11621 , RIdea0010_370, \8790_9089 );
and \U$2542 ( \11323_11622 , RIee1d650_4793, \8792_9091 );
and \U$2543 ( \11324_11623 , RIee1c570_4781, \8794_9093 );
and \U$2544 ( \11325_11624 , RIee1b5f8_4770, \8796_9095 );
and \U$2545 ( \11326_11625 , RIee1aef0_4765, \8798_9097 );
and \U$2546 ( \11327_11626 , RIfe99888_8091, \8800_9099 );
and \U$2547 ( \11328_11627 , RIfe99450_8088, \8802_9101 );
and \U$2548 ( \11329_11628 , RIfe99720_8090, \8804_9103 );
and \U$2549 ( \11330_11629 , RIfe995b8_8089, \8806_9105 );
and \U$2550 ( \11331_11630 , RIde83168_229, \8808_9107 );
and \U$2551 ( \11332_11631 , RIfcc43e8_7255, \8810_9109 );
and \U$2552 ( \11333_11632 , RIfcd5a58_7453, \8812_9111 );
and \U$2553 ( \11334_11633 , RIfc89450_6584, \8814_9113 );
and \U$2554 ( \11335_11634 , RIfcc5798_7269, \8816_9115 );
and \U$2555 ( \11336_11635 , RIe16c890_2612, \8818_9117 );
and \U$2556 ( \11337_11636 , RIe16a568_2587, \8820_9119 );
and \U$2557 ( \11338_11637 , RIe168d80_2570, \8822_9121 );
and \U$2558 ( \11339_11638 , RIe166788_2543, \8824_9123 );
and \U$2559 ( \11340_11639 , RIe163a88_2511, \8826_9125 );
and \U$2560 ( \11341_11640 , RIfc83618_6517, \8828_9127 );
and \U$2561 ( \11342_11641 , RIe160d88_2479, \8830_9129 );
and \U$2562 ( \11343_11642 , RIee36718_5078, \8832_9131 );
and \U$2563 ( \11344_11643 , RIe15e088_2447, \8834_9133 );
and \U$2564 ( \11345_11644 , RIe158688_2383, \8836_9135 );
and \U$2565 ( \11346_11645 , RIe155988_2351, \8838_9137 );
and \U$2566 ( \11347_11646 , RIfc3f800_5748, \8840_9139 );
and \U$2567 ( \11348_11647 , RIe152c88_2319, \8842_9141 );
and \U$2568 ( \11349_11648 , RIfc895b8_6585, \8844_9143 );
and \U$2569 ( \11350_11649 , RIe14ff88_2287, \8846_9145 );
and \U$2570 ( \11351_11650 , RIfc51cf8_5953, \8848_9147 );
and \U$2571 ( \11352_11651 , RIe14d288_2255, \8850_9149 );
and \U$2572 ( \11353_11652 , RIe14a588_2223, \8852_9151 );
and \U$2573 ( \11354_11653 , RIe147888_2191, \8854_9153 );
and \U$2574 ( \11355_11654 , RIee34990_5057, \8856_9155 );
and \U$2575 ( \11356_11655 , RIee338b0_5045, \8858_9157 );
and \U$2576 ( \11357_11656 , RIfc831e0_6514, \8860_9159 );
and \U$2577 ( \11358_11657 , RIfcd3b68_7431, \8862_9161 );
and \U$2578 ( \11359_11658 , RIe141ff0_2128, \8864_9163 );
and \U$2579 ( \11360_11659 , RIe13fcc8_2103, \8866_9165 );
and \U$2580 ( \11361_11660 , RIdf3dbd0_2079, \8868_9167 );
and \U$2581 ( \11362_11661 , RIdf3b740_2053, \8870_9169 );
and \U$2582 ( \11363_11662 , RIfcb6f90_7104, \8872_9171 );
and \U$2583 ( \11364_11663 , RIee301d8_5006, \8874_9173 );
and \U$2584 ( \11365_11664 , RIfcba938_7145, \8876_9175 );
and \U$2585 ( \11366_11665 , RIee2e018_4982, \8878_9177 );
and \U$2586 ( \11367_11666 , RIdf369e8_1998, \8880_9179 );
and \U$2587 ( \11368_11667 , RIdf343f0_1971, \8882_9181 );
and \U$2588 ( \11369_11668 , RIdf32230_1947, \8884_9183 );
and \U$2589 ( \11370_11669 , RIfe99e28_8095, \8886_9185 );
or \U$2590 ( \11371_11670 , \11307_11606 , \11308_11607 , \11309_11608 , \11310_11609 , \11311_11610 , \11312_11611 , \11313_11612 , \11314_11613 , \11315_11614 , \11316_11615 , \11317_11616 , \11318_11617 , \11319_11618 , \11320_11619 , \11321_11620 , \11322_11621 , \11323_11622 , \11324_11623 , \11325_11624 , \11326_11625 , \11327_11626 , \11328_11627 , \11329_11628 , \11330_11629 , \11331_11630 , \11332_11631 , \11333_11632 , \11334_11633 , \11335_11634 , \11336_11635 , \11337_11636 , \11338_11637 , \11339_11638 , \11340_11639 , \11341_11640 , \11342_11641 , \11343_11642 , \11344_11643 , \11345_11644 , \11346_11645 , \11347_11646 , \11348_11647 , \11349_11648 , \11350_11649 , \11351_11650 , \11352_11651 , \11353_11652 , \11354_11653 , \11355_11654 , \11356_11655 , \11357_11656 , \11358_11657 , \11359_11658 , \11360_11659 , \11361_11660 , \11362_11661 , \11363_11662 , \11364_11663 , \11365_11664 , \11366_11665 , \11367_11666 , \11368_11667 , \11369_11668 , \11370_11669 );
and \U$2591 ( \11372_11671 , RIfc83078_6513, \8889_9188 );
and \U$2592 ( \11373_11672 , RIfcb6e28_7103, \8891_9190 );
and \U$2593 ( \11374_11673 , RIfc9ad90_6784, \8893_9192 );
and \U$2594 ( \11375_11674 , RIfcbad70_7148, \8895_9194 );
and \U$2595 ( \11376_11675 , RIdf2b1b0_1867, \8897_9196 );
and \U$2596 ( \11377_11676 , RIdf292c0_1845, \8899_9198 );
and \U$2597 ( \11378_11677 , RIfe99b58_8093, \8901_9200 );
and \U$2598 ( \11379_11678 , RIfe999f0_8092, \8903_9202 );
and \U$2599 ( \11380_11679 , RIfc9ac28_6783, \8905_9204 );
and \U$2600 ( \11381_11680 , RIfc4a9a8_5871, \8907_9206 );
and \U$2601 ( \11382_11681 , RIdf23758_1780, \8909_9208 );
and \U$2602 ( \11383_11682 , RIfc82da8_6511, \8911_9210 );
and \U$2603 ( \11384_11683 , RIdf220d8_1764, \8913_9212 );
and \U$2604 ( \11385_11684 , RIdf20a58_1748, \8915_9214 );
and \U$2605 ( \11386_11685 , RIdf1ba30_1691, \8917_9216 );
and \U$2606 ( \11387_11686 , RIfe99cc0_8094, \8919_9218 );
and \U$2607 ( \11388_11687 , RIdf18358_1652, \8921_9220 );
and \U$2608 ( \11389_11688 , RIdf15658_1620, \8923_9222 );
and \U$2609 ( \11390_11689 , RIdf12958_1588, \8925_9224 );
and \U$2610 ( \11391_11690 , RIdf0fc58_1556, \8927_9226 );
and \U$2611 ( \11392_11691 , RIdf0cf58_1524, \8929_9228 );
and \U$2612 ( \11393_11692 , RIdf0a258_1492, \8931_9230 );
and \U$2613 ( \11394_11693 , RIdf07558_1460, \8933_9232 );
and \U$2614 ( \11395_11694 , RIdf04858_1428, \8935_9234 );
and \U$2615 ( \11396_11695 , RIdefee58_1364, \8937_9236 );
and \U$2616 ( \11397_11696 , RIdefc158_1332, \8939_9238 );
and \U$2617 ( \11398_11697 , RIdef9458_1300, \8941_9240 );
and \U$2618 ( \11399_11698 , RIdef6758_1268, \8943_9242 );
and \U$2619 ( \11400_11699 , RIdef3a58_1236, \8945_9244 );
and \U$2620 ( \11401_11700 , RIdef0d58_1204, \8947_9246 );
and \U$2621 ( \11402_11701 , RIdeee058_1172, \8949_9248 );
and \U$2622 ( \11403_11702 , RIdeeb358_1140, \8951_9250 );
and \U$2623 ( \11404_11703 , RIee25918_4886, \8953_9252 );
and \U$2624 ( \11405_11704 , RIee24b08_4876, \8955_9254 );
and \U$2625 ( \11406_11705 , RIfc52568_5959, \8957_9256 );
and \U$2626 ( \11407_11706 , RIfc826a0_6506, \8959_9258 );
and \U$2627 ( \11408_11707 , RIdee5958_1076, \8961_9260 );
and \U$2628 ( \11409_11708 , RIdee3bd0_1055, \8963_9262 );
and \U$2629 ( \11410_11709 , RIfe99f90_8096, \8965_9264 );
and \U$2630 ( \11411_11710 , RIdedf9b8_1008, \8967_9266 );
and \U$2631 ( \11412_11711 , RIfce4800_7622, \8969_9268 );
and \U$2632 ( \11413_11712 , RIfc89b58_6589, \8971_9270 );
and \U$2633 ( \11414_11713 , RIfc9f3e0_6834, \8973_9272 );
and \U$2634 ( \11415_11714 , RIfc82538_6505, \8975_9274 );
and \U$2635 ( \11416_11715 , RIdeda828_950, \8977_9276 );
and \U$2636 ( \11417_11716 , RIded8398_924, \8979_9278 );
and \U$2637 ( \11418_11717 , RIfeabe70_8272, \8981_9280 );
and \U$2638 ( \11419_11718 , RIded3eb0_875, \8983_9282 );
and \U$2639 ( \11420_11719 , RIded1b88_850, \8985_9284 );
and \U$2640 ( \11421_11720 , RIdecee88_818, \8987_9286 );
and \U$2641 ( \11422_11721 , RIdecc188_786, \8989_9288 );
and \U$2642 ( \11423_11722 , RIdec9488_754, \8991_9290 );
and \U$2643 ( \11424_11723 , RIdeb5988_530, \8993_9292 );
and \U$2644 ( \11425_11724 , RIde99710_338, \8995_9294 );
and \U$2645 ( \11426_11725 , RIe16f590_2644, \8997_9296 );
and \U$2646 ( \11427_11726 , RIe15b388_2415, \8999_9298 );
and \U$2647 ( \11428_11727 , RIe144b88_2159, \9001_9300 );
and \U$2648 ( \11429_11728 , RIdf39580_2029, \9003_9302 );
and \U$2649 ( \11430_11729 , RIdf2dbe0_1897, \9005_9304 );
and \U$2650 ( \11431_11730 , RIdf1e460_1721, \9007_9306 );
and \U$2651 ( \11432_11731 , RIdf01b58_1396, \9009_9308 );
and \U$2652 ( \11433_11732 , RIdee8658_1108, \9011_9310 );
and \U$2653 ( \11434_11733 , RIdedd3c0_981, \9013_9312 );
and \U$2654 ( \11435_11734 , RIde7f658_211, \9015_9314 );
or \U$2655 ( \11436_11735 , \11372_11671 , \11373_11672 , \11374_11673 , \11375_11674 , \11376_11675 , \11377_11676 , \11378_11677 , \11379_11678 , \11380_11679 , \11381_11680 , \11382_11681 , \11383_11682 , \11384_11683 , \11385_11684 , \11386_11685 , \11387_11686 , \11388_11687 , \11389_11688 , \11390_11689 , \11391_11690 , \11392_11691 , \11393_11692 , \11394_11693 , \11395_11694 , \11396_11695 , \11397_11696 , \11398_11697 , \11399_11698 , \11400_11699 , \11401_11700 , \11402_11701 , \11403_11702 , \11404_11703 , \11405_11704 , \11406_11705 , \11407_11706 , \11408_11707 , \11409_11708 , \11410_11709 , \11411_11710 , \11412_11711 , \11413_11712 , \11414_11713 , \11415_11714 , \11416_11715 , \11417_11716 , \11418_11717 , \11419_11718 , \11420_11719 , \11421_11720 , \11422_11721 , \11423_11722 , \11424_11723 , \11425_11724 , \11426_11725 , \11427_11726 , \11428_11727 , \11429_11728 , \11430_11729 , \11431_11730 , \11432_11731 , \11433_11732 , \11434_11733 , \11435_11734 );
or \U$2656 ( \11437_11736 , \11371_11670 , \11436_11735 );
_DC \g2fb7/U$1 ( \11438 , \11437_11736 , \9024_9323 );
buf \U$2657 ( \11439_11738 , \11438 );
and \U$2658 ( \11440_11739 , RIe19ea20_3182, \9034_9333 );
and \U$2659 ( \11441_11740 , RIe19bd20_3150, \9036_9335 );
and \U$2660 ( \11442_11741 , RIf145928_5251, \9038_9337 );
and \U$2661 ( \11443_11742 , RIe199020_3118, \9040_9339 );
and \U$2662 ( \11444_11743 , RIfe98910_8080, \9042_9341 );
and \U$2663 ( \11445_11744 , RIe196320_3086, \9044_9343 );
and \U$2664 ( \11446_11745 , RIe193620_3054, \9046_9345 );
and \U$2665 ( \11447_11746 , RIe190920_3022, \9048_9347 );
and \U$2666 ( \11448_11747 , RIe18af20_2958, \9050_9349 );
and \U$2667 ( \11449_11748 , RIe188220_2926, \9052_9351 );
and \U$2668 ( \11450_11749 , RIf143e70_5232, \9054_9353 );
and \U$2669 ( \11451_11750 , RIe185520_2894, \9056_9355 );
and \U$2670 ( \11452_11751 , RIfc95c00_6726, \9058_9357 );
and \U$2671 ( \11453_11752 , RIe182820_2862, \9060_9359 );
and \U$2672 ( \11454_11753 , RIe17fb20_2830, \9062_9361 );
and \U$2673 ( \11455_11754 , RIe17ce20_2798, \9064_9363 );
and \U$2674 ( \11456_11755 , RIf142520_5214, \9066_9365 );
and \U$2675 ( \11457_11756 , RIf141440_5202, \9068_9367 );
and \U$2676 ( \11458_11757 , RIe1776f0_2736, \9070_9369 );
and \U$2677 ( \11459_11758 , RIfeab8d0_8268, \9072_9371 );
and \U$2678 ( \11460_11759 , RIfcc5bd0_7272, \9074_9373 );
and \U$2679 ( \11461_11760 , RIfc62dc8_6147, \9076_9375 );
and \U$2680 ( \11462_11761 , RIee3e710_5169, \9078_9377 );
and \U$2681 ( \11463_11762 , RIfc9cb18_6805, \9080_9379 );
and \U$2682 ( \11464_11763 , RIee3c820_5147, \9082_9381 );
and \U$2683 ( \11465_11764 , RIee3b470_5133, \9084_9383 );
and \U$2684 ( \11466_11765 , RIee3a390_5121, \9086_9385 );
and \U$2685 ( \11467_11766 , RIe174888_2703, \9088_9387 );
and \U$2686 ( \11468_11767 , RIf170498_5737, \9090_9389 );
and \U$2687 ( \11469_11768 , RIfc68660_6210, \9092_9391 );
and \U$2688 ( \11470_11769 , RIf16e878_5717, \9094_9393 );
and \U$2689 ( \11471_11770 , RIfc6ea38_6281, \9096_9395 );
and \U$2690 ( \11472_11771 , RIfe98d48_8083, \9098_9397 );
and \U$2691 ( \11473_11772 , RIe224d78_4709, \9100_9399 );
and \U$2692 ( \11474_11773 , RIf16c280_5690, \9102_9401 );
and \U$2693 ( \11475_11774 , RIe222078_4677, \9104_9403 );
and \U$2694 ( \11476_11775 , RIf16b308_5679, \9106_9405 );
and \U$2695 ( \11477_11776 , RIe21f378_4645, \9108_9407 );
and \U$2696 ( \11478_11777 , RIe219978_4581, \9110_9409 );
and \U$2697 ( \11479_11778 , RIe216c78_4549, \9112_9411 );
and \U$2698 ( \11480_11779 , RIf16a390_5668, \9114_9413 );
and \U$2699 ( \11481_11780 , RIe213f78_4517, \9116_9415 );
and \U$2700 ( \11482_11781 , RIf169b20_5662, \9118_9417 );
and \U$2701 ( \11483_11782 , RIe211278_4485, \9120_9419 );
and \U$2702 ( \11484_11783 , RIf1681d0_5644, \9122_9421 );
and \U$2703 ( \11485_11784 , RIe20e578_4453, \9124_9423 );
and \U$2704 ( \11486_11785 , RIe20b878_4421, \9126_9425 );
and \U$2705 ( \11487_11786 , RIe208b78_4389, \9128_9427 );
and \U$2706 ( \11488_11787 , RIfcd4ae0_7442, \9130_9429 );
and \U$2707 ( \11489_11788 , RIfc61478_6129, \9132_9431 );
and \U$2708 ( \11490_11789 , RIfeab060_8262, \9134_9433 );
and \U$2709 ( \11491_11790 , RIe201990_4308, \9136_9435 );
and \U$2710 ( \11492_11791 , RIfc70ec8_6307, \9138_9437 );
and \U$2711 ( \11493_11792 , RIfc70928_6303, \9140_9439 );
and \U$2712 ( \11494_11793 , RIfcec528_7711, \9142_9441 );
and \U$2713 ( \11495_11794 , RIfcbe880_7190, \9144_9443 );
and \U$2714 ( \11496_11795 , RIf160d18_5561, \9146_9445 );
and \U$2715 ( \11497_11796 , RIf15ee28_5539, \9148_9447 );
and \U$2716 ( \11498_11797 , RIfe98be0_8082, \9150_9449 );
and \U$2717 ( \11499_11798 , RIfe98eb0_8084, \9152_9451 );
and \U$2718 ( \11500_11799 , RIf15d0a0_5518, \9154_9453 );
and \U$2719 ( \11501_11800 , RIf15bcf0_5504, \9156_9455 );
and \U$2720 ( \11502_11801 , RIfcd4540_7438, \9158_9457 );
and \U$2721 ( \11503_11802 , RIf159e00_5482, \9160_9459 );
or \U$2722 ( \11504_11803 , \11440_11739 , \11441_11740 , \11442_11741 , \11443_11742 , \11444_11743 , \11445_11744 , \11446_11745 , \11447_11746 , \11448_11747 , \11449_11748 , \11450_11749 , \11451_11750 , \11452_11751 , \11453_11752 , \11454_11753 , \11455_11754 , \11456_11755 , \11457_11756 , \11458_11757 , \11459_11758 , \11460_11759 , \11461_11760 , \11462_11761 , \11463_11762 , \11464_11763 , \11465_11764 , \11466_11765 , \11467_11766 , \11468_11767 , \11469_11768 , \11470_11769 , \11471_11770 , \11472_11771 , \11473_11772 , \11474_11773 , \11475_11774 , \11476_11775 , \11477_11776 , \11478_11777 , \11479_11778 , \11480_11779 , \11481_11780 , \11482_11781 , \11483_11782 , \11484_11783 , \11485_11784 , \11486_11785 , \11487_11786 , \11488_11787 , \11489_11788 , \11490_11789 , \11491_11790 , \11492_11791 , \11493_11792 , \11494_11793 , \11495_11794 , \11496_11795 , \11497_11796 , \11498_11797 , \11499_11798 , \11500_11799 , \11501_11800 , \11502_11801 , \11503_11802 );
and \U$2723 ( \11505_11804 , RIf1592c0_5474, \9163_9462 );
and \U$2724 ( \11506_11805 , RIf158078_5461, \9165_9464 );
and \U$2725 ( \11507_11806 , RIfca3a30_6884, \9167_9466 );
and \U$2726 ( \11508_11807 , RIfea7988_8223, \9169_9468 );
and \U$2727 ( \11509_11808 , RIf156728_5443, \9171_9470 );
and \U$2728 ( \11510_11809 , RIf155be8_5435, \9173_9472 );
and \U$2729 ( \11511_11810 , RIf154b08_5423, \9175_9474 );
and \U$2730 ( \11512_11811 , RIfe98a78_8081, \9177_9476 );
and \U$2731 ( \11513_11812 , RIf1538c0_5410, \9179_9478 );
and \U$2732 ( \11514_11813 , RIf1520d8_5393, \9181_9480 );
and \U$2733 ( \11515_11814 , RIf150e90_5380, \9183_9482 );
and \U$2734 ( \11516_11815 , RIe1f43d0_4156, \9185_9484 );
and \U$2735 ( \11517_11816 , RIf14fdb0_5368, \9187_9486 );
and \U$2736 ( \11518_11817 , RIfcd2380_7414, \9189_9488 );
and \U$2737 ( \11519_11818 , RIf14e2f8_5349, \9191_9490 );
and \U$2738 ( \11520_11819 , RIe1ef240_4098, \9193_9492 );
and \U$2739 ( \11521_11820 , RIe1ecae0_4070, \9195_9494 );
and \U$2740 ( \11522_11821 , RIe1e9de0_4038, \9197_9496 );
and \U$2741 ( \11523_11822 , RIe1e70e0_4006, \9199_9498 );
and \U$2742 ( \11524_11823 , RIe1e43e0_3974, \9201_9500 );
and \U$2743 ( \11525_11824 , RIe1e16e0_3942, \9203_9502 );
and \U$2744 ( \11526_11825 , RIe1de9e0_3910, \9205_9504 );
and \U$2745 ( \11527_11826 , RIe1dbce0_3878, \9207_9506 );
and \U$2746 ( \11528_11827 , RIe1d8fe0_3846, \9209_9508 );
and \U$2747 ( \11529_11828 , RIe1d35e0_3782, \9211_9510 );
and \U$2748 ( \11530_11829 , RIe1d08e0_3750, \9213_9512 );
and \U$2749 ( \11531_11830 , RIe1cdbe0_3718, \9215_9514 );
and \U$2750 ( \11532_11831 , RIe1caee0_3686, \9217_9516 );
and \U$2751 ( \11533_11832 , RIe1c81e0_3654, \9219_9518 );
and \U$2752 ( \11534_11833 , RIe1c54e0_3622, \9221_9520 );
and \U$2753 ( \11535_11834 , RIe1c27e0_3590, \9223_9522 );
and \U$2754 ( \11536_11835 , RIe1bfae0_3558, \9225_9524 );
and \U$2755 ( \11537_11836 , RIfc44b70_5804, \9227_9526 );
and \U$2756 ( \11538_11837 , RIf14bd00_5322, \9229_9528 );
and \U$2757 ( \11539_11838 , RIfe992e8_8087, \9231_9530 );
and \U$2758 ( \11540_11839 , RIfe987a8_8079, \9233_9532 );
and \U$2759 ( \11541_11840 , RIf14a950_5308, \9235_9534 );
and \U$2760 ( \11542_11841 , RIf149f78_5301, \9237_9536 );
and \U$2761 ( \11543_11842 , RIfe99180_8086, \9239_9538 );
and \U$2762 ( \11544_11843 , RIfe98640_8078, \9241_9540 );
and \U$2763 ( \11545_11844 , RIf149438_5293, \9243_9542 );
and \U$2764 ( \11546_11845 , RIfcec7f8_7713, \9245_9544 );
and \U$2765 ( \11547_11846 , RIfe984d8_8077, \9247_9546 );
and \U$2766 ( \11548_11847 , RIe1b1b48_3399, \9249_9548 );
and \U$2767 ( \11549_11848 , RIfc4b650_5880, \9251_9550 );
and \U$2768 ( \11550_11849 , RIfcda918_7509, \9253_9552 );
and \U$2769 ( \11551_11850 , RIfe98370_8076, \9255_9554 );
and \U$2770 ( \11552_11851 , RIfe99018_8085, \9257_9556 );
and \U$2771 ( \11553_11852 , RIe1a9e20_3310, \9259_9558 );
and \U$2772 ( \11554_11853 , RIe1a7120_3278, \9261_9560 );
and \U$2773 ( \11555_11854 , RIe1a4420_3246, \9263_9562 );
and \U$2774 ( \11556_11855 , RIe1a1720_3214, \9265_9564 );
and \U$2775 ( \11557_11856 , RIe18dc20_2990, \9267_9566 );
and \U$2776 ( \11558_11857 , RIe17a120_2766, \9269_9568 );
and \U$2777 ( \11559_11858 , RIe227a78_4741, \9271_9570 );
and \U$2778 ( \11560_11859 , RIe21c678_4613, \9273_9572 );
and \U$2779 ( \11561_11860 , RIe205e78_4357, \9275_9574 );
and \U$2780 ( \11562_11861 , RIe1ffed8_4289, \9277_9576 );
and \U$2781 ( \11563_11862 , RIe1f9290_4212, \9279_9578 );
and \U$2782 ( \11564_11863 , RIe1f1dd8_4129, \9281_9580 );
and \U$2783 ( \11565_11864 , RIe1d62e0_3814, \9283_9582 );
and \U$2784 ( \11566_11865 , RIe1bcde0_3526, \9285_9584 );
and \U$2785 ( \11567_11866 , RIe1afc58_3377, \9287_9586 );
and \U$2786 ( \11568_11867 , RIe172290_2676, \9289_9588 );
or \U$2787 ( \11569_11868 , \11505_11804 , \11506_11805 , \11507_11806 , \11508_11807 , \11509_11808 , \11510_11809 , \11511_11810 , \11512_11811 , \11513_11812 , \11514_11813 , \11515_11814 , \11516_11815 , \11517_11816 , \11518_11817 , \11519_11818 , \11520_11819 , \11521_11820 , \11522_11821 , \11523_11822 , \11524_11823 , \11525_11824 , \11526_11825 , \11527_11826 , \11528_11827 , \11529_11828 , \11530_11829 , \11531_11830 , \11532_11831 , \11533_11832 , \11534_11833 , \11535_11834 , \11536_11835 , \11537_11836 , \11538_11837 , \11539_11838 , \11540_11839 , \11541_11840 , \11542_11841 , \11543_11842 , \11544_11843 , \11545_11844 , \11546_11845 , \11547_11846 , \11548_11847 , \11549_11848 , \11550_11849 , \11551_11850 , \11552_11851 , \11553_11852 , \11554_11853 , \11555_11854 , \11556_11855 , \11557_11856 , \11558_11857 , \11559_11858 , \11560_11859 , \11561_11860 , \11562_11861 , \11563_11862 , \11564_11863 , \11565_11864 , \11566_11865 , \11567_11866 , \11568_11867 );
or \U$2788 ( \11570_11869 , \11504_11803 , \11569_11868 );
_DC \g40e4/U$1 ( \11571 , \11570_11869 , \9298_9597 );
buf \U$2789 ( \11572_11871 , \11571 );
xor \U$2790 ( \11573_11872 , \11439_11738 , \11572_11871 );
and \U$2791 ( \11574_11873 , RIdec6620_721, \8760_9059 );
and \U$2792 ( \11575_11874 , RIdec3920_689, \8762_9061 );
and \U$2793 ( \11576_11875 , RIfc49328_5855, \8764_9063 );
and \U$2794 ( \11577_11876 , RIdec0c20_657, \8766_9065 );
and \U$2795 ( \11578_11877 , RIfc80eb8_6489, \8768_9067 );
and \U$2796 ( \11579_11878 , RIdebdf20_625, \8770_9069 );
and \U$2797 ( \11580_11879 , RIdebb220_593, \8772_9071 );
and \U$2798 ( \11581_11880 , RIdeb8520_561, \8774_9073 );
and \U$2799 ( \11582_11881 , RIfc80648_6483, \8776_9075 );
and \U$2800 ( \11583_11882 , RIdeb2b20_497, \8778_9077 );
and \U$2801 ( \11584_11883 , RIfc8b340_6606, \8780_9079 );
and \U$2802 ( \11585_11884 , RIdeafe20_465, \8782_9081 );
and \U$2803 ( \11586_11885 , RIfc491c0_5854, \8784_9083 );
and \U$2804 ( \11587_11886 , RIdeacec8_433, \8786_9085 );
and \U$2805 ( \11588_11887 , RIdea65c8_401, \8788_9087 );
and \U$2806 ( \11589_11888 , RIde9fcc8_369, \8790_9089 );
and \U$2807 ( \11590_11889 , RIfcd9c70_7500, \8792_9091 );
and \U$2808 ( \11591_11890 , RIfe98208_8075, \8794_9093 );
and \U$2809 ( \11592_11891 , RIfce4698_7621, \8796_9095 );
and \U$2810 ( \11593_11892 , RIfe980a0_8074, \8798_9097 );
and \U$2811 ( \11594_11893 , RIde93158_307, \8800_9099 );
and \U$2812 ( \11595_11894 , RIde8f648_289, \8802_9101 );
and \U$2813 ( \11596_11895 , RIde8b4a8_269, \8804_9103 );
and \U$2814 ( \11597_11896 , RIde87308_249, \8806_9105 );
and \U$2815 ( \11598_11897 , RIde82e20_228, \8808_9107 );
and \U$2816 ( \11599_11898 , RIfcbba18_7157, \8810_9109 );
and \U$2817 ( \11600_11899 , RIfc48d88_5851, \8812_9111 );
and \U$2818 ( \11601_11900 , RIfc99f80_6774, \8814_9113 );
and \U$2819 ( \11602_11901 , RIfc8b4a8_6607, \8816_9115 );
and \U$2820 ( \11603_11902 , RIe16c728_2611, \8818_9117 );
and \U$2821 ( \11604_11903 , RIe16a400_2586, \8820_9119 );
and \U$2822 ( \11605_11904 , RIe168c18_2569, \8822_9121 );
and \U$2823 ( \11606_11905 , RIe166620_2542, \8824_9123 );
and \U$2824 ( \11607_11906 , RIe163920_2510, \8826_9125 );
and \U$2825 ( \11608_11907 , RIee38068_5096, \8828_9127 );
and \U$2826 ( \11609_11908 , RIe160c20_2478, \8830_9129 );
and \U$2827 ( \11610_11909 , RIfc48248_5843, \8832_9131 );
and \U$2828 ( \11611_11910 , RIe15df20_2446, \8834_9133 );
and \U$2829 ( \11612_11911 , RIe158520_2382, \8836_9135 );
and \U$2830 ( \11613_11912 , RIe155820_2350, \8838_9137 );
and \U$2831 ( \11614_11913 , RIfcbbe50_7160, \8840_9139 );
and \U$2832 ( \11615_11914 , RIe152b20_2318, \8842_9141 );
and \U$2833 ( \11616_11915 , RIfc47e10_5840, \8844_9143 );
and \U$2834 ( \11617_11916 , RIe14fe20_2286, \8846_9145 );
and \U$2835 ( \11618_11917 , RIfca0e98_6853, \8848_9147 );
and \U$2836 ( \11619_11918 , RIe14d120_2254, \8850_9149 );
and \U$2837 ( \11620_11919 , RIe14a420_2222, \8852_9151 );
and \U$2838 ( \11621_11920 , RIe147720_2190, \8854_9153 );
and \U$2839 ( \11622_11921 , RIfc8be80_6614, \8856_9155 );
and \U$2840 ( \11623_11922 , RIfc7fb08_6475, \8858_9157 );
and \U$2841 ( \11624_11923 , RIfc480e0_5842, \8860_9159 );
and \U$2842 ( \11625_11924 , RIfc99878_6769, \8862_9161 );
and \U$2843 ( \11626_11925 , RIe141e88_2127, \8864_9163 );
and \U$2844 ( \11627_11926 , RIe13fb60_2102, \8866_9165 );
and \U$2845 ( \11628_11927 , RIdf3da68_2078, \8868_9167 );
and \U$2846 ( \11629_11928 , RIdf3b5d8_2052, \8870_9169 );
and \U$2847 ( \11630_11929 , RIfe97f38_8073, \8872_9171 );
and \U$2848 ( \11631_11930 , RIee30070_5005, \8874_9173 );
and \U$2849 ( \11632_11931 , RIee2eb58_4990, \8876_9175 );
and \U$2850 ( \11633_11932 , RIee2deb0_4981, \8878_9177 );
and \U$2851 ( \11634_11933 , RIdf36880_1997, \8880_9179 );
and \U$2852 ( \11635_11934 , RIdf34288_1970, \8882_9181 );
and \U$2853 ( \11636_11935 , RIdf320c8_1946, \8884_9183 );
and \U$2854 ( \11637_11936 , RIfe97dd0_8072, \8886_9185 );
or \U$2855 ( \11638_11937 , \11574_11873 , \11575_11874 , \11576_11875 , \11577_11876 , \11578_11877 , \11579_11878 , \11580_11879 , \11581_11880 , \11582_11881 , \11583_11882 , \11584_11883 , \11585_11884 , \11586_11885 , \11587_11886 , \11588_11887 , \11589_11888 , \11590_11889 , \11591_11890 , \11592_11891 , \11593_11892 , \11594_11893 , \11595_11894 , \11596_11895 , \11597_11896 , \11598_11897 , \11599_11898 , \11600_11899 , \11601_11900 , \11602_11901 , \11603_11902 , \11604_11903 , \11605_11904 , \11606_11905 , \11607_11906 , \11608_11907 , \11609_11908 , \11610_11909 , \11611_11910 , \11612_11911 , \11613_11912 , \11614_11913 , \11615_11914 , \11616_11915 , \11617_11916 , \11618_11917 , \11619_11918 , \11620_11919 , \11621_11920 , \11622_11921 , \11623_11922 , \11624_11923 , \11625_11924 , \11626_11925 , \11627_11926 , \11628_11927 , \11629_11928 , \11630_11929 , \11631_11930 , \11632_11931 , \11633_11932 , \11634_11933 , \11635_11934 , \11636_11935 , \11637_11936 );
and \U$2856 ( \11639_11938 , RIfcc3740_7246, \8889_9188 );
and \U$2857 ( \11640_11939 , RIfc48ab8_5849, \8891_9190 );
and \U$2858 ( \11641_11940 , RIfce05e8_7575, \8893_9192 );
and \U$2859 ( \11642_11941 , RIfc80210_6480, \8895_9194 );
and \U$2860 ( \11643_11942 , RIdf2b048_1866, \8897_9196 );
and \U$2861 ( \11644_11943 , RIdf29158_1844, \8899_9198 );
and \U$2862 ( \11645_11944 , RIdf26f98_1820, \8901_9200 );
and \U$2863 ( \11646_11945 , RIdf254e0_1801, \8903_9202 );
and \U$2864 ( \11647_11946 , RIfc8bbb0_6612, \8905_9204 );
and \U$2865 ( \11648_11947 , RIfc48950_5848, \8907_9206 );
and \U$2866 ( \11649_11948 , RIdf235f0_1779, \8909_9208 );
and \U$2867 ( \11650_11949 , RIfc8bd18_6613, \8911_9210 );
and \U$2868 ( \11651_11950 , RIdf21f70_1763, \8913_9212 );
and \U$2869 ( \11652_11951 , RIdf208f0_1747, \8915_9214 );
and \U$2870 ( \11653_11952 , RIdf1b8c8_1690, \8917_9216 );
and \U$2871 ( \11654_11953 , RIdf1a3b0_1675, \8919_9218 );
and \U$2872 ( \11655_11954 , RIdf181f0_1651, \8921_9220 );
and \U$2873 ( \11656_11955 , RIdf154f0_1619, \8923_9222 );
and \U$2874 ( \11657_11956 , RIdf127f0_1587, \8925_9224 );
and \U$2875 ( \11658_11957 , RIdf0faf0_1555, \8927_9226 );
and \U$2876 ( \11659_11958 , RIdf0cdf0_1523, \8929_9228 );
and \U$2877 ( \11660_11959 , RIdf0a0f0_1491, \8931_9230 );
and \U$2878 ( \11661_11960 , RIdf073f0_1459, \8933_9232 );
and \U$2879 ( \11662_11961 , RIdf046f0_1427, \8935_9234 );
and \U$2880 ( \11663_11962 , RIdefecf0_1363, \8937_9236 );
and \U$2881 ( \11664_11963 , RIdefbff0_1331, \8939_9238 );
and \U$2882 ( \11665_11964 , RIdef92f0_1299, \8941_9240 );
and \U$2883 ( \11666_11965 , RIdef65f0_1267, \8943_9242 );
and \U$2884 ( \11667_11966 , RIdef38f0_1235, \8945_9244 );
and \U$2885 ( \11668_11967 , RIdef0bf0_1203, \8947_9246 );
and \U$2886 ( \11669_11968 , RIdeedef0_1171, \8949_9248 );
and \U$2887 ( \11670_11969 , RIdeeb1f0_1139, \8951_9250 );
and \U$2888 ( \11671_11970 , RIfcbc120_7162, \8953_9252 );
and \U$2889 ( \11672_11971 , RIfcd9838_7497, \8955_9254 );
and \U$2890 ( \11673_11972 , RIfc99710_6768, \8957_9256 );
and \U$2891 ( \11674_11973 , RIfca1168_6855, \8959_9258 );
and \U$2892 ( \11675_11974 , RIdee57f0_1075, \8961_9260 );
and \U$2893 ( \11676_11975 , RIdee3a68_1054, \8963_9262 );
and \U$2894 ( \11677_11976 , RIdee18a8_1030, \8965_9264 );
and \U$2895 ( \11678_11977 , RIdedf850_1007, \8967_9266 );
and \U$2896 ( \11679_11978 , RIfc549f8_5985, \8969_9268 );
and \U$2897 ( \11680_11979 , RIfcb5370_7084, \8971_9270 );
and \U$2898 ( \11681_11980 , RIfce43c8_7619, \8973_9272 );
and \U$2899 ( \11682_11981 , RIfce0480_7574, \8975_9274 );
and \U$2900 ( \11683_11982 , RIdeda6c0_949, \8977_9276 );
and \U$2901 ( \11684_11983 , RIded8230_923, \8979_9278 );
and \U$2902 ( \11685_11984 , RIded6070_899, \8981_9280 );
and \U$2903 ( \11686_11985 , RIded3d48_874, \8983_9282 );
and \U$2904 ( \11687_11986 , RIded1a20_849, \8985_9284 );
and \U$2905 ( \11688_11987 , RIdeced20_817, \8987_9286 );
and \U$2906 ( \11689_11988 , RIdecc020_785, \8989_9288 );
and \U$2907 ( \11690_11989 , RIdec9320_753, \8991_9290 );
and \U$2908 ( \11691_11990 , RIdeb5820_529, \8993_9292 );
and \U$2909 ( \11692_11991 , RIde993c8_337, \8995_9294 );
and \U$2910 ( \11693_11992 , RIe16f428_2643, \8997_9296 );
and \U$2911 ( \11694_11993 , RIe15b220_2414, \8999_9298 );
and \U$2912 ( \11695_11994 , RIe144a20_2158, \9001_9300 );
and \U$2913 ( \11696_11995 , RIdf39418_2028, \9003_9302 );
and \U$2914 ( \11697_11996 , RIdf2da78_1896, \9005_9304 );
and \U$2915 ( \11698_11997 , RIdf1e2f8_1720, \9007_9306 );
and \U$2916 ( \11699_11998 , RIdf019f0_1395, \9009_9308 );
and \U$2917 ( \11700_11999 , RIdee84f0_1107, \9011_9310 );
and \U$2918 ( \11701_12000 , RIdedd258_980, \9013_9312 );
and \U$2919 ( \11702_12001 , RIde7f310_210, \9015_9314 );
or \U$2920 ( \11703_12002 , \11639_11938 , \11640_11939 , \11641_11940 , \11642_11941 , \11643_11942 , \11644_11943 , \11645_11944 , \11646_11945 , \11647_11946 , \11648_11947 , \11649_11948 , \11650_11949 , \11651_11950 , \11652_11951 , \11653_11952 , \11654_11953 , \11655_11954 , \11656_11955 , \11657_11956 , \11658_11957 , \11659_11958 , \11660_11959 , \11661_11960 , \11662_11961 , \11663_11962 , \11664_11963 , \11665_11964 , \11666_11965 , \11667_11966 , \11668_11967 , \11669_11968 , \11670_11969 , \11671_11970 , \11672_11971 , \11673_11972 , \11674_11973 , \11675_11974 , \11676_11975 , \11677_11976 , \11678_11977 , \11679_11978 , \11680_11979 , \11681_11980 , \11682_11981 , \11683_11982 , \11684_11983 , \11685_11984 , \11686_11985 , \11687_11986 , \11688_11987 , \11689_11988 , \11690_11989 , \11691_11990 , \11692_11991 , \11693_11992 , \11694_11993 , \11695_11994 , \11696_11995 , \11697_11996 , \11698_11997 , \11699_11998 , \11700_11999 , \11701_12000 , \11702_12001 );
or \U$2921 ( \11704_12003 , \11638_11937 , \11703_12002 );
_DC \g303c/U$1 ( \11705 , \11704_12003 , \9024_9323 );
buf \U$2922 ( \11706_12005 , \11705 );
and \U$2923 ( \11707_12006 , RIe19e8b8_3181, \9034_9333 );
and \U$2924 ( \11708_12007 , RIe19bbb8_3149, \9036_9335 );
and \U$2925 ( \11709_12008 , RIfe976c8_8067, \9038_9337 );
and \U$2926 ( \11710_12009 , RIe198eb8_3117, \9040_9339 );
and \U$2927 ( \11711_12010 , RIf144c80_5242, \9042_9341 );
and \U$2928 ( \11712_12011 , RIe1961b8_3085, \9044_9343 );
and \U$2929 ( \11713_12012 , RIe1934b8_3053, \9046_9345 );
and \U$2930 ( \11714_12013 , RIe1907b8_3021, \9048_9347 );
and \U$2931 ( \11715_12014 , RIe18adb8_2957, \9050_9349 );
and \U$2932 ( \11716_12015 , RIe1880b8_2925, \9052_9351 );
and \U$2933 ( \11717_12016 , RIfe97560_8066, \9054_9353 );
and \U$2934 ( \11718_12017 , RIe1853b8_2893, \9056_9355 );
and \U$2935 ( \11719_12018 , RIfcc3fb0_7252, \9058_9357 );
and \U$2936 ( \11720_12019 , RIe1826b8_2861, \9060_9359 );
and \U$2937 ( \11721_12020 , RIe17f9b8_2829, \9062_9361 );
and \U$2938 ( \11722_12021 , RIe17ccb8_2797, \9064_9363 );
and \U$2939 ( \11723_12022 , RIfcd3730_7428, \9066_9365 );
and \U$2940 ( \11724_12023 , RIf1412d8_5201, \9068_9367 );
and \U$2941 ( \11725_12024 , RIfcc4118_7253, \9070_9369 );
and \U$2942 ( \11726_12025 , RIfe97830_8068, \9072_9371 );
and \U$2943 ( \11727_12026 , RIfc4a6d8_5869, \9074_9373 );
and \U$2944 ( \11728_12027 , RIf13f6b8_5181, \9076_9375 );
and \U$2945 ( \11729_12028 , RIfc9f980_6838, \9078_9377 );
and \U$2946 ( \11730_12029 , RIfc9fae8_6839, \9080_9379 );
and \U$2947 ( \11731_12030 , RIfcc3e48_7251, \9082_9381 );
and \U$2948 ( \11732_12031 , RIfc89e28_6591, \9084_9383 );
and \U$2949 ( \11733_12032 , RIfc89cc0_6590, \9086_9385 );
and \U$2950 ( \11734_12033 , RIe174720_2702, \9088_9387 );
and \U$2951 ( \11735_12034 , RIfc4a408_5867, \9090_9389 );
and \U$2952 ( \11736_12035 , RIfce27a8_7599, \9092_9391 );
and \U$2953 ( \11737_12036 , RIfc530a8_5967, \9094_9393 );
and \U$2954 ( \11738_12037 , RIfcd5d28_7455, \9096_9395 );
and \U$2955 ( \11739_12038 , RIf16cf28_5699, \9098_9397 );
and \U$2956 ( \11740_12039 , RIe224c10_4708, \9100_9399 );
and \U$2957 ( \11741_12040 , RIfc53210_5968, \9102_9401 );
and \U$2958 ( \11742_12041 , RIe221f10_4676, \9104_9403 );
and \U$2959 ( \11743_12042 , RIf16b1a0_5678, \9106_9405 );
and \U$2960 ( \11744_12043 , RIe21f210_4644, \9108_9407 );
and \U$2961 ( \11745_12044 , RIe219810_4580, \9110_9409 );
and \U$2962 ( \11746_12045 , RIe216b10_4548, \9112_9411 );
and \U$2963 ( \11747_12046 , RIfc401d8_5755, \9114_9413 );
and \U$2964 ( \11748_12047 , RIe213e10_4516, \9116_9415 );
and \U$2965 ( \11749_12048 , RIf1699b8_5661, \9118_9417 );
and \U$2966 ( \11750_12049 , RIe211110_4484, \9120_9419 );
and \U$2967 ( \11751_12050 , RIfc81cc8_6499, \9122_9421 );
and \U$2968 ( \11752_12051 , RIe20e410_4452, \9124_9423 );
and \U$2969 ( \11753_12052 , RIe20b710_4420, \9126_9425 );
and \U$2970 ( \11754_12053 , RIe208a10_4388, \9128_9427 );
and \U$2971 ( \11755_12054 , RIfc8a0f8_6593, \9130_9429 );
and \U$2972 ( \11756_12055 , RIfcb6720_7098, \9132_9431 );
and \U$2973 ( \11757_12056 , RIe203448_4327, \9134_9433 );
and \U$2974 ( \11758_12057 , RIe201828_4307, \9136_9435 );
and \U$2975 ( \11759_12058 , RIfc53378_5969, \9138_9437 );
and \U$2976 ( \11760_12059 , RIfc8a3c8_6595, \9140_9439 );
and \U$2977 ( \11761_12060 , RIfcb65b8_7097, \9142_9441 );
and \U$2978 ( \11762_12061 , RIfc49fd0_5864, \9144_9443 );
and \U$2979 ( \11763_12062 , RIf160bb0_5560, \9146_9445 );
and \U$2980 ( \11764_12063 , RIf15ecc0_5538, \9148_9447 );
and \U$2981 ( \11765_12064 , RIe1fd4a8_4259, \9150_9449 );
and \U$2982 ( \11766_12065 , RIfe97b00_8070, \9152_9451 );
and \U$2983 ( \11767_12066 , RIfc8a530_6596, \9154_9453 );
and \U$2984 ( \11768_12067 , RIfe97c68_8071, \9156_9455 );
and \U$2985 ( \11769_12068 , RIfc8a800_6598, \9158_9457 );
and \U$2986 ( \11770_12069 , RIfc8a698_6597, \9160_9459 );
or \U$2987 ( \11771_12070 , \11707_12006 , \11708_12007 , \11709_12008 , \11710_12009 , \11711_12010 , \11712_12011 , \11713_12012 , \11714_12013 , \11715_12014 , \11716_12015 , \11717_12016 , \11718_12017 , \11719_12018 , \11720_12019 , \11721_12020 , \11722_12021 , \11723_12022 , \11724_12023 , \11725_12024 , \11726_12025 , \11727_12026 , \11728_12027 , \11729_12028 , \11730_12029 , \11731_12030 , \11732_12031 , \11733_12032 , \11734_12033 , \11735_12034 , \11736_12035 , \11737_12036 , \11738_12037 , \11739_12038 , \11740_12039 , \11741_12040 , \11742_12041 , \11743_12042 , \11744_12043 , \11745_12044 , \11746_12045 , \11747_12046 , \11748_12047 , \11749_12048 , \11750_12049 , \11751_12050 , \11752_12051 , \11753_12052 , \11754_12053 , \11755_12054 , \11756_12055 , \11757_12056 , \11758_12057 , \11759_12058 , \11760_12059 , \11761_12060 , \11762_12061 , \11763_12062 , \11764_12063 , \11765_12064 , \11766_12065 , \11767_12066 , \11768_12067 , \11769_12068 , \11770_12069 );
and \U$2988 ( \11772_12071 , RIfc9a7f0_6780, \9163_9462 );
and \U$2989 ( \11773_12072 , RIfc81890_6496, \9165_9464 );
and \U$2990 ( \11774_12073 , RIfcd5e90_7456, \9167_9466 );
and \U$2991 ( \11775_12074 , RIe1fb180_4234, \9169_9468 );
and \U$2992 ( \11776_12075 , RIfc49e68_5863, \9171_9470 );
and \U$2993 ( \11777_12076 , RIfc81728_6495, \9173_9472 );
and \U$2994 ( \11778_12077 , RIfcbb1a8_7151, \9175_9474 );
and \U$2995 ( \11779_12078 , RIe1f66f8_4181, \9177_9476 );
and \U$2996 ( \11780_12079 , RIfcd3460_7426, \9179_9478 );
and \U$2997 ( \11781_12080 , RIfcb62e8_7095, \9181_9480 );
and \U$2998 ( \11782_12081 , RIfc9a520_6778, \9183_9482 );
and \U$2999 ( \11783_12082 , RIe1f4268_4155, \9185_9484 );
and \U$3000 ( \11784_12083 , RIfc49d00_5862, \9187_9486 );
and \U$3001 ( \11785_12084 , RIfcd9dd8_7501, \9189_9488 );
and \U$3002 ( \11786_12085 , RIfcbb310_7152, \9191_9490 );
and \U$3003 ( \11787_12086 , RIe1ef0d8_4097, \9193_9492 );
and \U$3004 ( \11788_12087 , RIe1ec978_4069, \9195_9494 );
and \U$3005 ( \11789_12088 , RIe1e9c78_4037, \9197_9496 );
and \U$3006 ( \11790_12089 , RIe1e6f78_4005, \9199_9498 );
and \U$3007 ( \11791_12090 , RIe1e4278_3973, \9201_9500 );
and \U$3008 ( \11792_12091 , RIe1e1578_3941, \9203_9502 );
and \U$3009 ( \11793_12092 , RIe1de878_3909, \9205_9504 );
and \U$3010 ( \11794_12093 , RIe1dbb78_3877, \9207_9506 );
and \U$3011 ( \11795_12094 , RIe1d8e78_3845, \9209_9508 );
and \U$3012 ( \11796_12095 , RIe1d3478_3781, \9211_9510 );
and \U$3013 ( \11797_12096 , RIe1d0778_3749, \9213_9512 );
and \U$3014 ( \11798_12097 , RIe1cda78_3717, \9215_9514 );
and \U$3015 ( \11799_12098 , RIe1cad78_3685, \9217_9516 );
and \U$3016 ( \11800_12099 , RIe1c8078_3653, \9219_9518 );
and \U$3017 ( \11801_12100 , RIe1c5378_3621, \9221_9520 );
and \U$3018 ( \11802_12101 , RIe1c2678_3589, \9223_9522 );
and \U$3019 ( \11803_12102 , RIe1bf978_3557, \9225_9524 );
and \U$3020 ( \11804_12103 , RIfc49a30_5860, \9227_9526 );
and \U$3021 ( \11805_12104 , RIfcb6018_7093, \9229_9528 );
and \U$3022 ( \11806_12105 , RIe1ba3b0_3496, \9231_9530 );
and \U$3023 ( \11807_12106 , RIe1b81f0_3472, \9233_9532 );
and \U$3024 ( \11808_12107 , RIfce0a20_7578, \9235_9534 );
and \U$3025 ( \11809_12108 , RIfcbb5e0_7154, \9237_9536 );
and \U$3026 ( \11810_12109 , RIe1b6030_3448, \9239_9538 );
and \U$3027 ( \11811_12110 , RIfe97998_8069, \9241_9540 );
and \U$3028 ( \11812_12111 , RIfce5610_7632, \9243_9542 );
and \U$3029 ( \11813_12112 , RIfcc3a10_7248, \9245_9544 );
and \U$3030 ( \11814_12113 , RIe1b3330_3416, \9247_9546 );
and \U$3031 ( \11815_12114 , RIe1b19e0_3398, \9249_9548 );
and \U$3032 ( \11816_12115 , RIfc495f8_5857, \9251_9550 );
and \U$3033 ( \11817_12116 , RIfc81188_6491, \9253_9552 );
and \U$3034 ( \11818_12117 , RIe1ad228_3347, \9255_9554 );
and \U$3035 ( \11819_12118 , RIe1aba40_3330, \9257_9556 );
and \U$3036 ( \11820_12119 , RIe1a9cb8_3309, \9259_9558 );
and \U$3037 ( \11821_12120 , RIe1a6fb8_3277, \9261_9560 );
and \U$3038 ( \11822_12121 , RIe1a42b8_3245, \9263_9562 );
and \U$3039 ( \11823_12122 , RIe1a15b8_3213, \9265_9564 );
and \U$3040 ( \11824_12123 , RIe18dab8_2989, \9267_9566 );
and \U$3041 ( \11825_12124 , RIe179fb8_2765, \9269_9568 );
and \U$3042 ( \11826_12125 , RIe227910_4740, \9271_9570 );
and \U$3043 ( \11827_12126 , RIe21c510_4612, \9273_9572 );
and \U$3044 ( \11828_12127 , RIe205d10_4356, \9275_9574 );
and \U$3045 ( \11829_12128 , RIe1ffd70_4288, \9277_9576 );
and \U$3046 ( \11830_12129 , RIe1f9128_4211, \9279_9578 );
and \U$3047 ( \11831_12130 , RIe1f1c70_4128, \9281_9580 );
and \U$3048 ( \11832_12131 , RIe1d6178_3813, \9283_9582 );
and \U$3049 ( \11833_12132 , RIe1bcc78_3525, \9285_9584 );
and \U$3050 ( \11834_12133 , RIe1afaf0_3376, \9287_9586 );
and \U$3051 ( \11835_12134 , RIe172128_2675, \9289_9588 );
or \U$3052 ( \11836_12135 , \11772_12071 , \11773_12072 , \11774_12073 , \11775_12074 , \11776_12075 , \11777_12076 , \11778_12077 , \11779_12078 , \11780_12079 , \11781_12080 , \11782_12081 , \11783_12082 , \11784_12083 , \11785_12084 , \11786_12085 , \11787_12086 , \11788_12087 , \11789_12088 , \11790_12089 , \11791_12090 , \11792_12091 , \11793_12092 , \11794_12093 , \11795_12094 , \11796_12095 , \11797_12096 , \11798_12097 , \11799_12098 , \11800_12099 , \11801_12100 , \11802_12101 , \11803_12102 , \11804_12103 , \11805_12104 , \11806_12105 , \11807_12106 , \11808_12107 , \11809_12108 , \11810_12109 , \11811_12110 , \11812_12111 , \11813_12112 , \11814_12113 , \11815_12114 , \11816_12115 , \11817_12116 , \11818_12117 , \11819_12118 , \11820_12119 , \11821_12120 , \11822_12121 , \11823_12122 , \11824_12123 , \11825_12124 , \11826_12125 , \11827_12126 , \11828_12127 , \11829_12128 , \11830_12129 , \11831_12130 , \11832_12131 , \11833_12132 , \11834_12133 , \11835_12134 );
or \U$3053 ( \11837_12136 , \11771_12070 , \11836_12135 );
_DC \g4169/U$1 ( \11838 , \11837_12136 , \9298_9597 );
buf \U$3054 ( \11839_12138 , \11838 );
and \U$3055 ( \11840_12139 , \11706_12005 , \11839_12138 );
and \U$3056 ( \11841_12140 , \9026_9325 , \9300_9599 );
and \U$3057 ( \11842_12141 , \9300_9599 , \10108_10407 );
and \U$3058 ( \11843_12142 , \9026_9325 , \10108_10407 );
or \U$3059 ( \11844_12143 , \11841_12140 , \11842_12141 , \11843_12142 );
and \U$3060 ( \11845_12144 , \11839_12138 , \11844_12143 );
and \U$3061 ( \11846_12145 , \11706_12005 , \11844_12143 );
or \U$3062 ( \11847_12146 , \11840_12139 , \11845_12144 , \11846_12145 );
xor \U$3063 ( \11848_12147 , \11573_11872 , \11847_12146 );
buf g4448_GF_PartitionCandidate( \11849_12148_nG4448 , \11848_12147 );
xor \U$3064 ( \11850_12149 , \11706_12005 , \11839_12138 );
xor \U$3065 ( \11851_12150 , \11850_12149 , \11844_12143 );
buf g444b_GF_PartitionCandidate( \11852_12151_nG444b , \11851_12150 );
nand \U$3066 ( \11853_12152 , \11852_12151_nG444b , \10110_10409_nG444e );
and \U$3067 ( \11854_12153 , \11849_12148_nG4448 , \11853_12152 );
xor \U$3068 ( \11855_12154 , \11852_12151_nG444b , \10110_10409_nG444e );
and \U$3073 ( \11856_12158 , \11855_12154 , \10392_10694_nG9c0e );
or \U$3074 ( \11857_12159 , 1'b0 , \11856_12158 );
xor \U$3075 ( \11858_12160 , \11854_12153 , \11857_12159 );
xor \U$3076 ( \11859_12161 , \11854_12153 , \11858_12160 );
buf \U$3077 ( \11860_12162 , \11859_12161 );
buf \U$3078 ( \11861_12163 , \11860_12162 );
and \U$3079 ( \11862_12164 , \11306_11605 , \11861_12163 );
and \U$3080 ( \11863_12165 , \10993_11295 , \11002_11301 );
buf \U$3081 ( \11864_12166 , \11863_12165 );
and \U$3082 ( \11865_12167 , \10996_10421 , \10693_10995_nG9c0b );
and \U$3083 ( \11866_12168 , \10119_10418 , \10981_11283_nG9c08 );
or \U$3084 ( \11867_12169 , \11865_12167 , \11866_12168 );
xor \U$3085 ( \11868_12170 , \10118_10417 , \11867_12169 );
buf \U$3086 ( \11869_12171 , \11868_12170 );
buf \U$3088 ( \11870_12172 , \11869_12171 );
xor \U$3089 ( \11871_12173 , \11864_12166 , \11870_12172 );
buf \U$3090 ( \11872_12174 , \11871_12173 );
and \U$3091 ( \11873_12175 , \10990_11292 , \11004_11303 );
and \U$3092 ( \11874_12176 , \10990_11292 , \11304_11603 );
and \U$3093 ( \11875_12177 , \11004_11303 , \11304_11603 );
or \U$3094 ( \11876_12178 , \11873_12175 , \11874_12176 , \11875_12177 );
buf \U$3095 ( \11877_12179 , \11876_12178 );
xor \U$3096 ( \11878_12180 , \11872_12174 , \11877_12179 );
and \U$3097 ( \11879_12181 , \10411_10707 , \11299_11598_nG9c05 );
and \U$3098 ( \11880_12182 , \11287_11586 , \10681_10983 );
and \U$3099 ( \11881_12183 , RIdec6620_721, \9034_9333 );
and \U$3100 ( \11882_12184 , RIdec3920_689, \9036_9335 );
and \U$3101 ( \11883_12185 , RIfc49328_5855, \9038_9337 );
and \U$3102 ( \11884_12186 , RIdec0c20_657, \9040_9339 );
and \U$3103 ( \11885_12187 , RIfc80eb8_6489, \9042_9341 );
and \U$3104 ( \11886_12188 , RIdebdf20_625, \9044_9343 );
and \U$3105 ( \11887_12189 , RIdebb220_593, \9046_9345 );
and \U$3106 ( \11888_12190 , RIdeb8520_561, \9048_9347 );
and \U$3107 ( \11889_12191 , RIfc80648_6483, \9050_9349 );
and \U$3108 ( \11890_12192 , RIdeb2b20_497, \9052_9351 );
and \U$3109 ( \11891_12193 , RIfc8b340_6606, \9054_9353 );
and \U$3110 ( \11892_12194 , RIdeafe20_465, \9056_9355 );
and \U$3111 ( \11893_12195 , RIfc491c0_5854, \9058_9357 );
and \U$3112 ( \11894_12196 , RIdeacec8_433, \9060_9359 );
and \U$3113 ( \11895_12197 , RIdea65c8_401, \9062_9361 );
and \U$3114 ( \11896_12198 , RIde9fcc8_369, \9064_9363 );
and \U$3115 ( \11897_12199 , RIfcd9c70_7500, \9066_9365 );
and \U$3116 ( \11898_12200 , RIfe98208_8075, \9068_9367 );
and \U$3117 ( \11899_12201 , RIfce4698_7621, \9070_9369 );
and \U$3118 ( \11900_12202 , RIfe980a0_8074, \9072_9371 );
and \U$3119 ( \11901_12203 , RIde93158_307, \9074_9373 );
and \U$3120 ( \11902_12204 , RIde8f648_289, \9076_9375 );
and \U$3121 ( \11903_12205 , RIde8b4a8_269, \9078_9377 );
and \U$3122 ( \11904_12206 , RIde87308_249, \9080_9379 );
and \U$3123 ( \11905_12207 , RIde82e20_228, \9082_9381 );
and \U$3124 ( \11906_12208 , RIfcbba18_7157, \9084_9383 );
and \U$3125 ( \11907_12209 , RIfc48d88_5851, \9086_9385 );
and \U$3126 ( \11908_12210 , RIfc99f80_6774, \9088_9387 );
and \U$3127 ( \11909_12211 , RIfc8b4a8_6607, \9090_9389 );
and \U$3128 ( \11910_12212 , RIe16c728_2611, \9092_9391 );
and \U$3129 ( \11911_12213 , RIe16a400_2586, \9094_9393 );
and \U$3130 ( \11912_12214 , RIe168c18_2569, \9096_9395 );
and \U$3131 ( \11913_12215 , RIe166620_2542, \9098_9397 );
and \U$3132 ( \11914_12216 , RIe163920_2510, \9100_9399 );
and \U$3133 ( \11915_12217 , RIee38068_5096, \9102_9401 );
and \U$3134 ( \11916_12218 , RIe160c20_2478, \9104_9403 );
and \U$3135 ( \11917_12219 , RIfc48248_5843, \9106_9405 );
and \U$3136 ( \11918_12220 , RIe15df20_2446, \9108_9407 );
and \U$3137 ( \11919_12221 , RIe158520_2382, \9110_9409 );
and \U$3138 ( \11920_12222 , RIe155820_2350, \9112_9411 );
and \U$3139 ( \11921_12223 , RIfcbbe50_7160, \9114_9413 );
and \U$3140 ( \11922_12224 , RIe152b20_2318, \9116_9415 );
and \U$3141 ( \11923_12225 , RIfc47e10_5840, \9118_9417 );
and \U$3142 ( \11924_12226 , RIe14fe20_2286, \9120_9419 );
and \U$3143 ( \11925_12227 , RIfca0e98_6853, \9122_9421 );
and \U$3144 ( \11926_12228 , RIe14d120_2254, \9124_9423 );
and \U$3145 ( \11927_12229 , RIe14a420_2222, \9126_9425 );
and \U$3146 ( \11928_12230 , RIe147720_2190, \9128_9427 );
and \U$3147 ( \11929_12231 , RIfc8be80_6614, \9130_9429 );
and \U$3148 ( \11930_12232 , RIfc7fb08_6475, \9132_9431 );
and \U$3149 ( \11931_12233 , RIfc480e0_5842, \9134_9433 );
and \U$3150 ( \11932_12234 , RIfc99878_6769, \9136_9435 );
and \U$3151 ( \11933_12235 , RIe141e88_2127, \9138_9437 );
and \U$3152 ( \11934_12236 , RIe13fb60_2102, \9140_9439 );
and \U$3153 ( \11935_12237 , RIdf3da68_2078, \9142_9441 );
and \U$3154 ( \11936_12238 , RIdf3b5d8_2052, \9144_9443 );
and \U$3155 ( \11937_12239 , RIfe97f38_8073, \9146_9445 );
and \U$3156 ( \11938_12240 , RIee30070_5005, \9148_9447 );
and \U$3157 ( \11939_12241 , RIee2eb58_4990, \9150_9449 );
and \U$3158 ( \11940_12242 , RIee2deb0_4981, \9152_9451 );
and \U$3159 ( \11941_12243 , RIdf36880_1997, \9154_9453 );
and \U$3160 ( \11942_12244 , RIdf34288_1970, \9156_9455 );
and \U$3161 ( \11943_12245 , RIdf320c8_1946, \9158_9457 );
and \U$3162 ( \11944_12246 , RIfe97dd0_8072, \9160_9459 );
or \U$3163 ( \11945_12247 , \11881_12183 , \11882_12184 , \11883_12185 , \11884_12186 , \11885_12187 , \11886_12188 , \11887_12189 , \11888_12190 , \11889_12191 , \11890_12192 , \11891_12193 , \11892_12194 , \11893_12195 , \11894_12196 , \11895_12197 , \11896_12198 , \11897_12199 , \11898_12200 , \11899_12201 , \11900_12202 , \11901_12203 , \11902_12204 , \11903_12205 , \11904_12206 , \11905_12207 , \11906_12208 , \11907_12209 , \11908_12210 , \11909_12211 , \11910_12212 , \11911_12213 , \11912_12214 , \11913_12215 , \11914_12216 , \11915_12217 , \11916_12218 , \11917_12219 , \11918_12220 , \11919_12221 , \11920_12222 , \11921_12223 , \11922_12224 , \11923_12225 , \11924_12226 , \11925_12227 , \11926_12228 , \11927_12229 , \11928_12230 , \11929_12231 , \11930_12232 , \11931_12233 , \11932_12234 , \11933_12235 , \11934_12236 , \11935_12237 , \11936_12238 , \11937_12239 , \11938_12240 , \11939_12241 , \11940_12242 , \11941_12243 , \11942_12244 , \11943_12245 , \11944_12246 );
and \U$3164 ( \11946_12248 , RIfcc3740_7246, \9163_9462 );
and \U$3165 ( \11947_12249 , RIfc48ab8_5849, \9165_9464 );
and \U$3166 ( \11948_12250 , RIfce05e8_7575, \9167_9466 );
and \U$3167 ( \11949_12251 , RIfc80210_6480, \9169_9468 );
and \U$3168 ( \11950_12252 , RIdf2b048_1866, \9171_9470 );
and \U$3169 ( \11951_12253 , RIdf29158_1844, \9173_9472 );
and \U$3170 ( \11952_12254 , RIdf26f98_1820, \9175_9474 );
and \U$3171 ( \11953_12255 , RIdf254e0_1801, \9177_9476 );
and \U$3172 ( \11954_12256 , RIfc8bbb0_6612, \9179_9478 );
and \U$3173 ( \11955_12257 , RIfc48950_5848, \9181_9480 );
and \U$3174 ( \11956_12258 , RIdf235f0_1779, \9183_9482 );
and \U$3175 ( \11957_12259 , RIfc8bd18_6613, \9185_9484 );
and \U$3176 ( \11958_12260 , RIdf21f70_1763, \9187_9486 );
and \U$3177 ( \11959_12261 , RIdf208f0_1747, \9189_9488 );
and \U$3178 ( \11960_12262 , RIdf1b8c8_1690, \9191_9490 );
and \U$3179 ( \11961_12263 , RIdf1a3b0_1675, \9193_9492 );
and \U$3180 ( \11962_12264 , RIdf181f0_1651, \9195_9494 );
and \U$3181 ( \11963_12265 , RIdf154f0_1619, \9197_9496 );
and \U$3182 ( \11964_12266 , RIdf127f0_1587, \9199_9498 );
and \U$3183 ( \11965_12267 , RIdf0faf0_1555, \9201_9500 );
and \U$3184 ( \11966_12268 , RIdf0cdf0_1523, \9203_9502 );
and \U$3185 ( \11967_12269 , RIdf0a0f0_1491, \9205_9504 );
and \U$3186 ( \11968_12270 , RIdf073f0_1459, \9207_9506 );
and \U$3187 ( \11969_12271 , RIdf046f0_1427, \9209_9508 );
and \U$3188 ( \11970_12272 , RIdefecf0_1363, \9211_9510 );
and \U$3189 ( \11971_12273 , RIdefbff0_1331, \9213_9512 );
and \U$3190 ( \11972_12274 , RIdef92f0_1299, \9215_9514 );
and \U$3191 ( \11973_12275 , RIdef65f0_1267, \9217_9516 );
and \U$3192 ( \11974_12276 , RIdef38f0_1235, \9219_9518 );
and \U$3193 ( \11975_12277 , RIdef0bf0_1203, \9221_9520 );
and \U$3194 ( \11976_12278 , RIdeedef0_1171, \9223_9522 );
and \U$3195 ( \11977_12279 , RIdeeb1f0_1139, \9225_9524 );
and \U$3196 ( \11978_12280 , RIfcbc120_7162, \9227_9526 );
and \U$3197 ( \11979_12281 , RIfcd9838_7497, \9229_9528 );
and \U$3198 ( \11980_12282 , RIfc99710_6768, \9231_9530 );
and \U$3199 ( \11981_12283 , RIfca1168_6855, \9233_9532 );
and \U$3200 ( \11982_12284 , RIdee57f0_1075, \9235_9534 );
and \U$3201 ( \11983_12285 , RIdee3a68_1054, \9237_9536 );
and \U$3202 ( \11984_12286 , RIdee18a8_1030, \9239_9538 );
and \U$3203 ( \11985_12287 , RIdedf850_1007, \9241_9540 );
and \U$3204 ( \11986_12288 , RIfc549f8_5985, \9243_9542 );
and \U$3205 ( \11987_12289 , RIfcb5370_7084, \9245_9544 );
and \U$3206 ( \11988_12290 , RIfce43c8_7619, \9247_9546 );
and \U$3207 ( \11989_12291 , RIfce0480_7574, \9249_9548 );
and \U$3208 ( \11990_12292 , RIdeda6c0_949, \9251_9550 );
and \U$3209 ( \11991_12293 , RIded8230_923, \9253_9552 );
and \U$3210 ( \11992_12294 , RIded6070_899, \9255_9554 );
and \U$3211 ( \11993_12295 , RIded3d48_874, \9257_9556 );
and \U$3212 ( \11994_12296 , RIded1a20_849, \9259_9558 );
and \U$3213 ( \11995_12297 , RIdeced20_817, \9261_9560 );
and \U$3214 ( \11996_12298 , RIdecc020_785, \9263_9562 );
and \U$3215 ( \11997_12299 , RIdec9320_753, \9265_9564 );
and \U$3216 ( \11998_12300 , RIdeb5820_529, \9267_9566 );
and \U$3217 ( \11999_12301 , RIde993c8_337, \9269_9568 );
and \U$3218 ( \12000_12302 , RIe16f428_2643, \9271_9570 );
and \U$3219 ( \12001_12303 , RIe15b220_2414, \9273_9572 );
and \U$3220 ( \12002_12304 , RIe144a20_2158, \9275_9574 );
and \U$3221 ( \12003_12305 , RIdf39418_2028, \9277_9576 );
and \U$3222 ( \12004_12306 , RIdf2da78_1896, \9279_9578 );
and \U$3223 ( \12005_12307 , RIdf1e2f8_1720, \9281_9580 );
and \U$3224 ( \12006_12308 , RIdf019f0_1395, \9283_9582 );
and \U$3225 ( \12007_12309 , RIdee84f0_1107, \9285_9584 );
and \U$3226 ( \12008_12310 , RIdedd258_980, \9287_9586 );
and \U$3227 ( \12009_12311 , RIde7f310_210, \9289_9588 );
or \U$3228 ( \12010_12312 , \11946_12248 , \11947_12249 , \11948_12250 , \11949_12251 , \11950_12252 , \11951_12253 , \11952_12254 , \11953_12255 , \11954_12256 , \11955_12257 , \11956_12258 , \11957_12259 , \11958_12260 , \11959_12261 , \11960_12262 , \11961_12263 , \11962_12264 , \11963_12265 , \11964_12266 , \11965_12267 , \11966_12268 , \11967_12269 , \11968_12270 , \11969_12271 , \11970_12272 , \11971_12273 , \11972_12274 , \11973_12275 , \11974_12276 , \11975_12277 , \11976_12278 , \11977_12279 , \11978_12280 , \11979_12281 , \11980_12282 , \11981_12283 , \11982_12284 , \11983_12285 , \11984_12286 , \11985_12287 , \11986_12288 , \11987_12289 , \11988_12290 , \11989_12291 , \11990_12292 , \11991_12293 , \11992_12294 , \11993_12295 , \11994_12296 , \11995_12297 , \11996_12298 , \11997_12299 , \11998_12300 , \11999_12301 , \12000_12302 , \12001_12303 , \12002_12304 , \12003_12305 , \12004_12306 , \12005_12307 , \12006_12308 , \12007_12309 , \12008_12310 , \12009_12311 );
or \U$3229 ( \12011_12313 , \11945_12247 , \12010_12312 );
_DC \g6583/U$1 ( \12012 , \12011_12313 , \9298_9597 );
and \U$3230 ( \12013_12315 , RIe19e8b8_3181, \8760_9059 );
and \U$3231 ( \12014_12316 , RIe19bbb8_3149, \8762_9061 );
and \U$3232 ( \12015_12317 , RIfe976c8_8067, \8764_9063 );
and \U$3233 ( \12016_12318 , RIe198eb8_3117, \8766_9065 );
and \U$3234 ( \12017_12319 , RIf144c80_5242, \8768_9067 );
and \U$3235 ( \12018_12320 , RIe1961b8_3085, \8770_9069 );
and \U$3236 ( \12019_12321 , RIe1934b8_3053, \8772_9071 );
and \U$3237 ( \12020_12322 , RIe1907b8_3021, \8774_9073 );
and \U$3238 ( \12021_12323 , RIe18adb8_2957, \8776_9075 );
and \U$3239 ( \12022_12324 , RIe1880b8_2925, \8778_9077 );
and \U$3240 ( \12023_12325 , RIfe97560_8066, \8780_9079 );
and \U$3241 ( \12024_12326 , RIe1853b8_2893, \8782_9081 );
and \U$3242 ( \12025_12327 , RIfcc3fb0_7252, \8784_9083 );
and \U$3243 ( \12026_12328 , RIe1826b8_2861, \8786_9085 );
and \U$3244 ( \12027_12329 , RIe17f9b8_2829, \8788_9087 );
and \U$3245 ( \12028_12330 , RIe17ccb8_2797, \8790_9089 );
and \U$3246 ( \12029_12331 , RIfcd3730_7428, \8792_9091 );
and \U$3247 ( \12030_12332 , RIf1412d8_5201, \8794_9093 );
and \U$3248 ( \12031_12333 , RIfcc4118_7253, \8796_9095 );
and \U$3249 ( \12032_12334 , RIfe97830_8068, \8798_9097 );
and \U$3250 ( \12033_12335 , RIfc4a6d8_5869, \8800_9099 );
and \U$3251 ( \12034_12336 , RIf13f6b8_5181, \8802_9101 );
and \U$3252 ( \12035_12337 , RIfc9f980_6838, \8804_9103 );
and \U$3253 ( \12036_12338 , RIfc9fae8_6839, \8806_9105 );
and \U$3254 ( \12037_12339 , RIfcc3e48_7251, \8808_9107 );
and \U$3255 ( \12038_12340 , RIfc89e28_6591, \8810_9109 );
and \U$3256 ( \12039_12341 , RIfc89cc0_6590, \8812_9111 );
and \U$3257 ( \12040_12342 , RIe174720_2702, \8814_9113 );
and \U$3258 ( \12041_12343 , RIfc4a408_5867, \8816_9115 );
and \U$3259 ( \12042_12344 , RIfce27a8_7599, \8818_9117 );
and \U$3260 ( \12043_12345 , RIfc530a8_5967, \8820_9119 );
and \U$3261 ( \12044_12346 , RIfcd5d28_7455, \8822_9121 );
and \U$3262 ( \12045_12347 , RIf16cf28_5699, \8824_9123 );
and \U$3263 ( \12046_12348 , RIe224c10_4708, \8826_9125 );
and \U$3264 ( \12047_12349 , RIfc53210_5968, \8828_9127 );
and \U$3265 ( \12048_12350 , RIe221f10_4676, \8830_9129 );
and \U$3266 ( \12049_12351 , RIf16b1a0_5678, \8832_9131 );
and \U$3267 ( \12050_12352 , RIe21f210_4644, \8834_9133 );
and \U$3268 ( \12051_12353 , RIe219810_4580, \8836_9135 );
and \U$3269 ( \12052_12354 , RIe216b10_4548, \8838_9137 );
and \U$3270 ( \12053_12355 , RIfc401d8_5755, \8840_9139 );
and \U$3271 ( \12054_12356 , RIe213e10_4516, \8842_9141 );
and \U$3272 ( \12055_12357 , RIf1699b8_5661, \8844_9143 );
and \U$3273 ( \12056_12358 , RIe211110_4484, \8846_9145 );
and \U$3274 ( \12057_12359 , RIfc81cc8_6499, \8848_9147 );
and \U$3275 ( \12058_12360 , RIe20e410_4452, \8850_9149 );
and \U$3276 ( \12059_12361 , RIe20b710_4420, \8852_9151 );
and \U$3277 ( \12060_12362 , RIe208a10_4388, \8854_9153 );
and \U$3278 ( \12061_12363 , RIfc8a0f8_6593, \8856_9155 );
and \U$3279 ( \12062_12364 , RIfcb6720_7098, \8858_9157 );
and \U$3280 ( \12063_12365 , RIe203448_4327, \8860_9159 );
and \U$3281 ( \12064_12366 , RIe201828_4307, \8862_9161 );
and \U$3282 ( \12065_12367 , RIfc53378_5969, \8864_9163 );
and \U$3283 ( \12066_12368 , RIfc8a3c8_6595, \8866_9165 );
and \U$3284 ( \12067_12369 , RIfcb65b8_7097, \8868_9167 );
and \U$3285 ( \12068_12370 , RIfc49fd0_5864, \8870_9169 );
and \U$3286 ( \12069_12371 , RIf160bb0_5560, \8872_9171 );
and \U$3287 ( \12070_12372 , RIf15ecc0_5538, \8874_9173 );
and \U$3288 ( \12071_12373 , RIe1fd4a8_4259, \8876_9175 );
and \U$3289 ( \12072_12374 , RIfe97b00_8070, \8878_9177 );
and \U$3290 ( \12073_12375 , RIfc8a530_6596, \8880_9179 );
and \U$3291 ( \12074_12376 , RIfe97c68_8071, \8882_9181 );
and \U$3292 ( \12075_12377 , RIfc8a800_6598, \8884_9183 );
and \U$3293 ( \12076_12378 , RIfc8a698_6597, \8886_9185 );
or \U$3294 ( \12077_12379 , \12013_12315 , \12014_12316 , \12015_12317 , \12016_12318 , \12017_12319 , \12018_12320 , \12019_12321 , \12020_12322 , \12021_12323 , \12022_12324 , \12023_12325 , \12024_12326 , \12025_12327 , \12026_12328 , \12027_12329 , \12028_12330 , \12029_12331 , \12030_12332 , \12031_12333 , \12032_12334 , \12033_12335 , \12034_12336 , \12035_12337 , \12036_12338 , \12037_12339 , \12038_12340 , \12039_12341 , \12040_12342 , \12041_12343 , \12042_12344 , \12043_12345 , \12044_12346 , \12045_12347 , \12046_12348 , \12047_12349 , \12048_12350 , \12049_12351 , \12050_12352 , \12051_12353 , \12052_12354 , \12053_12355 , \12054_12356 , \12055_12357 , \12056_12358 , \12057_12359 , \12058_12360 , \12059_12361 , \12060_12362 , \12061_12363 , \12062_12364 , \12063_12365 , \12064_12366 , \12065_12367 , \12066_12368 , \12067_12369 , \12068_12370 , \12069_12371 , \12070_12372 , \12071_12373 , \12072_12374 , \12073_12375 , \12074_12376 , \12075_12377 , \12076_12378 );
and \U$3295 ( \12078_12380 , RIfc9a7f0_6780, \8889_9188 );
and \U$3296 ( \12079_12381 , RIfc81890_6496, \8891_9190 );
and \U$3297 ( \12080_12382 , RIfcd5e90_7456, \8893_9192 );
and \U$3298 ( \12081_12383 , RIe1fb180_4234, \8895_9194 );
and \U$3299 ( \12082_12384 , RIfc49e68_5863, \8897_9196 );
and \U$3300 ( \12083_12385 , RIfc81728_6495, \8899_9198 );
and \U$3301 ( \12084_12386 , RIfcbb1a8_7151, \8901_9200 );
and \U$3302 ( \12085_12387 , RIe1f66f8_4181, \8903_9202 );
and \U$3303 ( \12086_12388 , RIfcd3460_7426, \8905_9204 );
and \U$3304 ( \12087_12389 , RIfcb62e8_7095, \8907_9206 );
and \U$3305 ( \12088_12390 , RIfc9a520_6778, \8909_9208 );
and \U$3306 ( \12089_12391 , RIe1f4268_4155, \8911_9210 );
and \U$3307 ( \12090_12392 , RIfc49d00_5862, \8913_9212 );
and \U$3308 ( \12091_12393 , RIfcd9dd8_7501, \8915_9214 );
and \U$3309 ( \12092_12394 , RIfcbb310_7152, \8917_9216 );
and \U$3310 ( \12093_12395 , RIe1ef0d8_4097, \8919_9218 );
and \U$3311 ( \12094_12396 , RIe1ec978_4069, \8921_9220 );
and \U$3312 ( \12095_12397 , RIe1e9c78_4037, \8923_9222 );
and \U$3313 ( \12096_12398 , RIe1e6f78_4005, \8925_9224 );
and \U$3314 ( \12097_12399 , RIe1e4278_3973, \8927_9226 );
and \U$3315 ( \12098_12400 , RIe1e1578_3941, \8929_9228 );
and \U$3316 ( \12099_12401 , RIe1de878_3909, \8931_9230 );
and \U$3317 ( \12100_12402 , RIe1dbb78_3877, \8933_9232 );
and \U$3318 ( \12101_12403 , RIe1d8e78_3845, \8935_9234 );
and \U$3319 ( \12102_12404 , RIe1d3478_3781, \8937_9236 );
and \U$3320 ( \12103_12405 , RIe1d0778_3749, \8939_9238 );
and \U$3321 ( \12104_12406 , RIe1cda78_3717, \8941_9240 );
and \U$3322 ( \12105_12407 , RIe1cad78_3685, \8943_9242 );
and \U$3323 ( \12106_12408 , RIe1c8078_3653, \8945_9244 );
and \U$3324 ( \12107_12409 , RIe1c5378_3621, \8947_9246 );
and \U$3325 ( \12108_12410 , RIe1c2678_3589, \8949_9248 );
and \U$3326 ( \12109_12411 , RIe1bf978_3557, \8951_9250 );
and \U$3327 ( \12110_12412 , RIfc49a30_5860, \8953_9252 );
and \U$3328 ( \12111_12413 , RIfcb6018_7093, \8955_9254 );
and \U$3329 ( \12112_12414 , RIe1ba3b0_3496, \8957_9256 );
and \U$3330 ( \12113_12415 , RIe1b81f0_3472, \8959_9258 );
and \U$3331 ( \12114_12416 , RIfce0a20_7578, \8961_9260 );
and \U$3332 ( \12115_12417 , RIfcbb5e0_7154, \8963_9262 );
and \U$3333 ( \12116_12418 , RIe1b6030_3448, \8965_9264 );
and \U$3334 ( \12117_12419 , RIfe97998_8069, \8967_9266 );
and \U$3335 ( \12118_12420 , RIfce5610_7632, \8969_9268 );
and \U$3336 ( \12119_12421 , RIfcc3a10_7248, \8971_9270 );
and \U$3337 ( \12120_12422 , RIe1b3330_3416, \8973_9272 );
and \U$3338 ( \12121_12423 , RIe1b19e0_3398, \8975_9274 );
and \U$3339 ( \12122_12424 , RIfc495f8_5857, \8977_9276 );
and \U$3340 ( \12123_12425 , RIfc81188_6491, \8979_9278 );
and \U$3341 ( \12124_12426 , RIe1ad228_3347, \8981_9280 );
and \U$3342 ( \12125_12427 , RIe1aba40_3330, \8983_9282 );
and \U$3343 ( \12126_12428 , RIe1a9cb8_3309, \8985_9284 );
and \U$3344 ( \12127_12429 , RIe1a6fb8_3277, \8987_9286 );
and \U$3345 ( \12128_12430 , RIe1a42b8_3245, \8989_9288 );
and \U$3346 ( \12129_12431 , RIe1a15b8_3213, \8991_9290 );
and \U$3347 ( \12130_12432 , RIe18dab8_2989, \8993_9292 );
and \U$3348 ( \12131_12433 , RIe179fb8_2765, \8995_9294 );
and \U$3349 ( \12132_12434 , RIe227910_4740, \8997_9296 );
and \U$3350 ( \12133_12435 , RIe21c510_4612, \8999_9298 );
and \U$3351 ( \12134_12436 , RIe205d10_4356, \9001_9300 );
and \U$3352 ( \12135_12437 , RIe1ffd70_4288, \9003_9302 );
and \U$3353 ( \12136_12438 , RIe1f9128_4211, \9005_9304 );
and \U$3354 ( \12137_12439 , RIe1f1c70_4128, \9007_9306 );
and \U$3355 ( \12138_12440 , RIe1d6178_3813, \9009_9308 );
and \U$3356 ( \12139_12441 , RIe1bcc78_3525, \9011_9310 );
and \U$3357 ( \12140_12442 , RIe1afaf0_3376, \9013_9312 );
and \U$3358 ( \12141_12443 , RIe172128_2675, \9015_9314 );
or \U$3359 ( \12142_12444 , \12078_12380 , \12079_12381 , \12080_12382 , \12081_12383 , \12082_12384 , \12083_12385 , \12084_12386 , \12085_12387 , \12086_12388 , \12087_12389 , \12088_12390 , \12089_12391 , \12090_12392 , \12091_12393 , \12092_12394 , \12093_12395 , \12094_12396 , \12095_12397 , \12096_12398 , \12097_12399 , \12098_12400 , \12099_12401 , \12100_12402 , \12101_12403 , \12102_12404 , \12103_12405 , \12104_12406 , \12105_12407 , \12106_12408 , \12107_12409 , \12108_12410 , \12109_12411 , \12110_12412 , \12111_12413 , \12112_12414 , \12113_12415 , \12114_12416 , \12115_12417 , \12116_12418 , \12117_12419 , \12118_12420 , \12119_12421 , \12120_12422 , \12121_12423 , \12122_12424 , \12123_12425 , \12124_12426 , \12125_12427 , \12126_12428 , \12127_12429 , \12128_12430 , \12129_12431 , \12130_12432 , \12131_12433 , \12132_12434 , \12133_12435 , \12134_12436 , \12135_12437 , \12136_12438 , \12137_12439 , \12138_12440 , \12139_12441 , \12140_12442 , \12141_12443 );
or \U$3360 ( \12143_12445 , \12077_12379 , \12142_12444 );
_DC \g6584/U$1 ( \12144 , \12143_12445 , \9024_9323 );
and g6585_GF_PartitionCandidate( \12145_12447_nG6585 , \12012 , \12144 );
buf \U$3361 ( \12146_12448 , \12145_12447_nG6585 );
and \U$3362 ( \12147_12449 , \12146_12448 , \10389_10691 );
nor \U$3363 ( \12148_12450 , \11880_12182 , \12147_12449 );
xnor \U$3364 ( \12149_12451 , \12148_12450 , \10678_10980 );
and \U$3365 ( \12150_12452 , \10686_10988 , \11275_11574 );
and \U$3366 ( \12151_12453 , \10968_11270 , \10976_11278 );
nor \U$3367 ( \12152_12454 , \12150_12452 , \12151_12453 );
xnor \U$3368 ( \12153_12455 , \12152_12454 , \11281_11580 );
xor \U$3369 ( \12154_12456 , \12149_12451 , \12153_12455 );
_DC \g48fe/U$1 ( \12155 , \12011_12313 , \9298_9597 );
_DC \g4982/U$1 ( \12156 , \12143_12445 , \9024_9323 );
xor g4983_GF_PartitionCandidate( \12157_12459_nG4983 , \12155 , \12156 );
buf \U$3370 ( \12158_12460 , \12157_12459_nG4983 );
xor \U$3371 ( \12159_12461 , \12158_12460 , \11272_11571 );
and \U$3372 ( \12160_12462 , \10385_10687 , \12159_12461 );
xor \U$3373 ( \12161_12463 , \12154_12456 , \12160_12462 );
and \U$3374 ( \12162_12464 , \11290_11589 , \11292_11591 );
xor \U$3375 ( \12163_12465 , \12161_12463 , \12162_12464 );
and \U$3376 ( \12164_12466 , \11282_11581 , \11293_11592 );
and \U$3377 ( \12165_12467 , \11294_11593 , \11297_11596 );
or \U$3378 ( \12166_12468 , \12164_12466 , \12165_12467 );
xor \U$3379 ( \12167_12469 , \12163_12465 , \12166_12468 );
buf g9c02_GF_PartitionCandidate( \12168_12470_nG9c02 , \12167_12469 );
and \U$3380 ( \12169_12471 , \10402_10704 , \12168_12470_nG9c02 );
or \U$3381 ( \12170_12472 , \11879_12181 , \12169_12471 );
xor \U$3382 ( \12171_12473 , \10399_10703 , \12170_12472 );
buf \U$3383 ( \12172_12474 , \12171_12473 );
buf \U$3385 ( \12173_12475 , \12172_12474 );
xor \U$3386 ( \12174_12476 , \11878_12180 , \12173_12475 );
and \U$3387 ( \12175_12477 , \11306_11605 , \12174_12476 );
and \U$3388 ( \12176_12478 , \11861_12163 , \12174_12476 );
or \U$3389 ( \12177_12479 , \11862_12164 , \12175_12477 , \12176_12478 );
and \U$3390 ( \12178_12480 , \11854_12153 , \11858_12160 );
buf \U$3391 ( \12179_12481 , \12178_12480 );
buf \U$3393 ( \12180_12482 , \12179_12481 );
not \U$3069 ( \12181_12155 , \11855_12154 );
xor \U$3070 ( \12182_12156 , \11849_12148_nG4448 , \11852_12151_nG444b );
and \U$3071 ( \12183_12157 , \12181_12155 , \12182_12156 );
and \U$3394 ( \12184_12483 , \12183_12157 , \10392_10694_nG9c0e );
and \U$3395 ( \12185_12484 , \11855_12154 , \10693_10995_nG9c0b );
or \U$3396 ( \12186_12485 , \12184_12483 , \12185_12484 );
xor \U$3397 ( \12187_12486 , \11854_12153 , \12186_12485 );
buf \U$3398 ( \12188_12487 , \12187_12486 );
buf \U$3400 ( \12189_12488 , \12188_12487 );
xor \U$3401 ( \12190_12489 , \12180_12482 , \12189_12488 );
buf \U$3402 ( \12191_12490 , \12190_12489 );
and \U$3403 ( \12192_12491 , \10996_10421 , \10981_11283_nG9c08 );
and \U$3404 ( \12193_12492 , \10119_10418 , \11299_11598_nG9c05 );
or \U$3405 ( \12194_12493 , \12192_12491 , \12193_12492 );
xor \U$3406 ( \12195_12494 , \10118_10417 , \12194_12493 );
buf \U$3407 ( \12196_12495 , \12195_12494 );
buf \U$3409 ( \12197_12496 , \12196_12495 );
xor \U$3410 ( \12198_12497 , \12191_12490 , \12197_12496 );
and \U$3411 ( \12199_12498 , \10411_10707 , \12168_12470_nG9c02 );
and \U$3412 ( \12200_12499 , \12149_12451 , \12153_12455 );
and \U$3413 ( \12201_12500 , \12153_12455 , \12160_12462 );
and \U$3414 ( \12202_12501 , \12149_12451 , \12160_12462 );
or \U$3415 ( \12203_12502 , \12200_12499 , \12201_12500 , \12202_12501 );
and \U$3416 ( \12204_12503 , \12146_12448 , \10681_10983 );
and \U$3417 ( \12205_12504 , RIdec6788_722, \9034_9333 );
and \U$3418 ( \12206_12505 , RIdec3a88_690, \9036_9335 );
and \U$3419 ( \12207_12506 , RIee20788_4828, \9038_9337 );
and \U$3420 ( \12208_12507 , RIdec0d88_658, \9040_9339 );
and \U$3421 ( \12209_12508 , RIee1f810_4817, \9042_9341 );
and \U$3422 ( \12210_12509 , RIdebe088_626, \9044_9343 );
and \U$3423 ( \12211_12510 , RIdebb388_594, \9046_9345 );
and \U$3424 ( \12212_12511 , RIdeb8688_562, \9048_9347 );
and \U$3425 ( \12213_12512 , RIfc9b1c8_6787, \9050_9349 );
and \U$3426 ( \12214_12513 , RIdeb2c88_498, \9052_9351 );
and \U$3427 ( \12215_12514 , RIfce1f38_7593, \9054_9353 );
and \U$3428 ( \12216_12515 , RIdeaff88_466, \9056_9355 );
and \U$3429 ( \12217_12516 , RIfc892e8_6583, \9058_9357 );
and \U$3430 ( \12218_12517 , RIdead210_434, \9060_9359 );
and \U$3431 ( \12219_12518 , RIdea6910_402, \9062_9361 );
and \U$3432 ( \12220_12519 , RIdea0010_370, \9064_9363 );
and \U$3433 ( \12221_12520 , RIee1d650_4793, \9066_9365 );
and \U$3434 ( \12222_12521 , RIee1c570_4781, \9068_9367 );
and \U$3435 ( \12223_12522 , RIee1b5f8_4770, \9070_9369 );
and \U$3436 ( \12224_12523 , RIee1aef0_4765, \9072_9371 );
and \U$3437 ( \12225_12524 , RIfe99888_8091, \9074_9373 );
and \U$3438 ( \12226_12525 , RIfe99450_8088, \9076_9375 );
and \U$3439 ( \12227_12526 , RIfe99720_8090, \9078_9377 );
and \U$3440 ( \12228_12527 , RIfe995b8_8089, \9080_9379 );
and \U$3441 ( \12229_12528 , RIde83168_229, \9082_9381 );
and \U$3442 ( \12230_12529 , RIfcc43e8_7255, \9084_9383 );
and \U$3443 ( \12231_12530 , RIfcd5a58_7453, \9086_9385 );
and \U$3444 ( \12232_12531 , RIfc89450_6584, \9088_9387 );
and \U$3445 ( \12233_12532 , RIfcc5798_7269, \9090_9389 );
and \U$3446 ( \12234_12533 , RIe16c890_2612, \9092_9391 );
and \U$3447 ( \12235_12534 , RIe16a568_2587, \9094_9393 );
and \U$3448 ( \12236_12535 , RIe168d80_2570, \9096_9395 );
and \U$3449 ( \12237_12536 , RIe166788_2543, \9098_9397 );
and \U$3450 ( \12238_12537 , RIe163a88_2511, \9100_9399 );
and \U$3451 ( \12239_12538 , RIfc83618_6517, \9102_9401 );
and \U$3452 ( \12240_12539 , RIe160d88_2479, \9104_9403 );
and \U$3453 ( \12241_12540 , RIee36718_5078, \9106_9405 );
and \U$3454 ( \12242_12541 , RIe15e088_2447, \9108_9407 );
and \U$3455 ( \12243_12542 , RIe158688_2383, \9110_9409 );
and \U$3456 ( \12244_12543 , RIe155988_2351, \9112_9411 );
and \U$3457 ( \12245_12544 , RIfc3f800_5748, \9114_9413 );
and \U$3458 ( \12246_12545 , RIe152c88_2319, \9116_9415 );
and \U$3459 ( \12247_12546 , RIfc895b8_6585, \9118_9417 );
and \U$3460 ( \12248_12547 , RIe14ff88_2287, \9120_9419 );
and \U$3461 ( \12249_12548 , RIfc51cf8_5953, \9122_9421 );
and \U$3462 ( \12250_12549 , RIe14d288_2255, \9124_9423 );
and \U$3463 ( \12251_12550 , RIe14a588_2223, \9126_9425 );
and \U$3464 ( \12252_12551 , RIe147888_2191, \9128_9427 );
and \U$3465 ( \12253_12552 , RIee34990_5057, \9130_9429 );
and \U$3466 ( \12254_12553 , RIee338b0_5045, \9132_9431 );
and \U$3467 ( \12255_12554 , RIfc831e0_6514, \9134_9433 );
and \U$3468 ( \12256_12555 , RIfcd3b68_7431, \9136_9435 );
and \U$3469 ( \12257_12556 , RIe141ff0_2128, \9138_9437 );
and \U$3470 ( \12258_12557 , RIe13fcc8_2103, \9140_9439 );
and \U$3471 ( \12259_12558 , RIdf3dbd0_2079, \9142_9441 );
and \U$3472 ( \12260_12559 , RIdf3b740_2053, \9144_9443 );
and \U$3473 ( \12261_12560 , RIfcb6f90_7104, \9146_9445 );
and \U$3474 ( \12262_12561 , RIee301d8_5006, \9148_9447 );
and \U$3475 ( \12263_12562 , RIfcba938_7145, \9150_9449 );
and \U$3476 ( \12264_12563 , RIee2e018_4982, \9152_9451 );
and \U$3477 ( \12265_12564 , RIdf369e8_1998, \9154_9453 );
and \U$3478 ( \12266_12565 , RIdf343f0_1971, \9156_9455 );
and \U$3479 ( \12267_12566 , RIdf32230_1947, \9158_9457 );
and \U$3480 ( \12268_12567 , RIfe99e28_8095, \9160_9459 );
or \U$3481 ( \12269_12568 , \12205_12504 , \12206_12505 , \12207_12506 , \12208_12507 , \12209_12508 , \12210_12509 , \12211_12510 , \12212_12511 , \12213_12512 , \12214_12513 , \12215_12514 , \12216_12515 , \12217_12516 , \12218_12517 , \12219_12518 , \12220_12519 , \12221_12520 , \12222_12521 , \12223_12522 , \12224_12523 , \12225_12524 , \12226_12525 , \12227_12526 , \12228_12527 , \12229_12528 , \12230_12529 , \12231_12530 , \12232_12531 , \12233_12532 , \12234_12533 , \12235_12534 , \12236_12535 , \12237_12536 , \12238_12537 , \12239_12538 , \12240_12539 , \12241_12540 , \12242_12541 , \12243_12542 , \12244_12543 , \12245_12544 , \12246_12545 , \12247_12546 , \12248_12547 , \12249_12548 , \12250_12549 , \12251_12550 , \12252_12551 , \12253_12552 , \12254_12553 , \12255_12554 , \12256_12555 , \12257_12556 , \12258_12557 , \12259_12558 , \12260_12559 , \12261_12560 , \12262_12561 , \12263_12562 , \12264_12563 , \12265_12564 , \12266_12565 , \12267_12566 , \12268_12567 );
and \U$3482 ( \12270_12569 , RIfc83078_6513, \9163_9462 );
and \U$3483 ( \12271_12570 , RIfcb6e28_7103, \9165_9464 );
and \U$3484 ( \12272_12571 , RIfc9ad90_6784, \9167_9466 );
and \U$3485 ( \12273_12572 , RIfcbad70_7148, \9169_9468 );
and \U$3486 ( \12274_12573 , RIdf2b1b0_1867, \9171_9470 );
and \U$3487 ( \12275_12574 , RIdf292c0_1845, \9173_9472 );
and \U$3488 ( \12276_12575 , RIfe99b58_8093, \9175_9474 );
and \U$3489 ( \12277_12576 , RIfe999f0_8092, \9177_9476 );
and \U$3490 ( \12278_12577 , RIfc9ac28_6783, \9179_9478 );
and \U$3491 ( \12279_12578 , RIfc4a9a8_5871, \9181_9480 );
and \U$3492 ( \12280_12579 , RIdf23758_1780, \9183_9482 );
and \U$3493 ( \12281_12580 , RIfc82da8_6511, \9185_9484 );
and \U$3494 ( \12282_12581 , RIdf220d8_1764, \9187_9486 );
and \U$3495 ( \12283_12582 , RIdf20a58_1748, \9189_9488 );
and \U$3496 ( \12284_12583 , RIdf1ba30_1691, \9191_9490 );
and \U$3497 ( \12285_12584 , RIfe99cc0_8094, \9193_9492 );
and \U$3498 ( \12286_12585 , RIdf18358_1652, \9195_9494 );
and \U$3499 ( \12287_12586 , RIdf15658_1620, \9197_9496 );
and \U$3500 ( \12288_12587 , RIdf12958_1588, \9199_9498 );
and \U$3501 ( \12289_12588 , RIdf0fc58_1556, \9201_9500 );
and \U$3502 ( \12290_12589 , RIdf0cf58_1524, \9203_9502 );
and \U$3503 ( \12291_12590 , RIdf0a258_1492, \9205_9504 );
and \U$3504 ( \12292_12591 , RIdf07558_1460, \9207_9506 );
and \U$3505 ( \12293_12592 , RIdf04858_1428, \9209_9508 );
and \U$3506 ( \12294_12593 , RIdefee58_1364, \9211_9510 );
and \U$3507 ( \12295_12594 , RIdefc158_1332, \9213_9512 );
and \U$3508 ( \12296_12595 , RIdef9458_1300, \9215_9514 );
and \U$3509 ( \12297_12596 , RIdef6758_1268, \9217_9516 );
and \U$3510 ( \12298_12597 , RIdef3a58_1236, \9219_9518 );
and \U$3511 ( \12299_12598 , RIdef0d58_1204, \9221_9520 );
and \U$3512 ( \12300_12599 , RIdeee058_1172, \9223_9522 );
and \U$3513 ( \12301_12600 , RIdeeb358_1140, \9225_9524 );
and \U$3514 ( \12302_12601 , RIee25918_4886, \9227_9526 );
and \U$3515 ( \12303_12602 , RIee24b08_4876, \9229_9528 );
and \U$3516 ( \12304_12603 , RIfc52568_5959, \9231_9530 );
and \U$3517 ( \12305_12604 , RIfc826a0_6506, \9233_9532 );
and \U$3518 ( \12306_12605 , RIdee5958_1076, \9235_9534 );
and \U$3519 ( \12307_12606 , RIdee3bd0_1055, \9237_9536 );
and \U$3520 ( \12308_12607 , RIfe99f90_8096, \9239_9538 );
and \U$3521 ( \12309_12608 , RIdedf9b8_1008, \9241_9540 );
and \U$3522 ( \12310_12609 , RIfce4800_7622, \9243_9542 );
and \U$3523 ( \12311_12610 , RIfc89b58_6589, \9245_9544 );
and \U$3524 ( \12312_12611 , RIfc9f3e0_6834, \9247_9546 );
and \U$3525 ( \12313_12612 , RIfc82538_6505, \9249_9548 );
and \U$3526 ( \12314_12613 , RIdeda828_950, \9251_9550 );
and \U$3527 ( \12315_12614 , RIded8398_924, \9253_9552 );
and \U$3528 ( \12316_12615 , RIfeabe70_8272, \9255_9554 );
and \U$3529 ( \12317_12616 , RIded3eb0_875, \9257_9556 );
and \U$3530 ( \12318_12617 , RIded1b88_850, \9259_9558 );
and \U$3531 ( \12319_12618 , RIdecee88_818, \9261_9560 );
and \U$3532 ( \12320_12619 , RIdecc188_786, \9263_9562 );
and \U$3533 ( \12321_12620 , RIdec9488_754, \9265_9564 );
and \U$3534 ( \12322_12621 , RIdeb5988_530, \9267_9566 );
and \U$3535 ( \12323_12622 , RIde99710_338, \9269_9568 );
and \U$3536 ( \12324_12623 , RIe16f590_2644, \9271_9570 );
and \U$3537 ( \12325_12624 , RIe15b388_2415, \9273_9572 );
and \U$3538 ( \12326_12625 , RIe144b88_2159, \9275_9574 );
and \U$3539 ( \12327_12626 , RIdf39580_2029, \9277_9576 );
and \U$3540 ( \12328_12627 , RIdf2dbe0_1897, \9279_9578 );
and \U$3541 ( \12329_12628 , RIdf1e460_1721, \9281_9580 );
and \U$3542 ( \12330_12629 , RIdf01b58_1396, \9283_9582 );
and \U$3543 ( \12331_12630 , RIdee8658_1108, \9285_9584 );
and \U$3544 ( \12332_12631 , RIdedd3c0_981, \9287_9586 );
and \U$3545 ( \12333_12632 , RIde7f658_211, \9289_9588 );
or \U$3546 ( \12334_12633 , \12270_12569 , \12271_12570 , \12272_12571 , \12273_12572 , \12274_12573 , \12275_12574 , \12276_12575 , \12277_12576 , \12278_12577 , \12279_12578 , \12280_12579 , \12281_12580 , \12282_12581 , \12283_12582 , \12284_12583 , \12285_12584 , \12286_12585 , \12287_12586 , \12288_12587 , \12289_12588 , \12290_12589 , \12291_12590 , \12292_12591 , \12293_12592 , \12294_12593 , \12295_12594 , \12296_12595 , \12297_12596 , \12298_12597 , \12299_12598 , \12300_12599 , \12301_12600 , \12302_12601 , \12303_12602 , \12304_12603 , \12305_12604 , \12306_12605 , \12307_12606 , \12308_12607 , \12309_12608 , \12310_12609 , \12311_12610 , \12312_12611 , \12313_12612 , \12314_12613 , \12315_12614 , \12316_12615 , \12317_12616 , \12318_12617 , \12319_12618 , \12320_12619 , \12321_12620 , \12322_12621 , \12323_12622 , \12324_12623 , \12325_12624 , \12326_12625 , \12327_12626 , \12328_12627 , \12329_12628 , \12330_12629 , \12331_12630 , \12332_12631 , \12333_12632 );
or \U$3547 ( \12335_12634 , \12269_12568 , \12334_12633 );
_DC \g6586/U$1 ( \12336 , \12335_12634 , \9298_9597 );
and \U$3548 ( \12337_12636 , RIe19ea20_3182, \8760_9059 );
and \U$3549 ( \12338_12637 , RIe19bd20_3150, \8762_9061 );
and \U$3550 ( \12339_12638 , RIf145928_5251, \8764_9063 );
and \U$3551 ( \12340_12639 , RIe199020_3118, \8766_9065 );
and \U$3552 ( \12341_12640 , RIfe98910_8080, \8768_9067 );
and \U$3553 ( \12342_12641 , RIe196320_3086, \8770_9069 );
and \U$3554 ( \12343_12642 , RIe193620_3054, \8772_9071 );
and \U$3555 ( \12344_12643 , RIe190920_3022, \8774_9073 );
and \U$3556 ( \12345_12644 , RIe18af20_2958, \8776_9075 );
and \U$3557 ( \12346_12645 , RIe188220_2926, \8778_9077 );
and \U$3558 ( \12347_12646 , RIf143e70_5232, \8780_9079 );
and \U$3559 ( \12348_12647 , RIe185520_2894, \8782_9081 );
and \U$3560 ( \12349_12648 , RIfc95c00_6726, \8784_9083 );
and \U$3561 ( \12350_12649 , RIe182820_2862, \8786_9085 );
and \U$3562 ( \12351_12650 , RIe17fb20_2830, \8788_9087 );
and \U$3563 ( \12352_12651 , RIe17ce20_2798, \8790_9089 );
and \U$3564 ( \12353_12652 , RIf142520_5214, \8792_9091 );
and \U$3565 ( \12354_12653 , RIf141440_5202, \8794_9093 );
and \U$3566 ( \12355_12654 , RIe1776f0_2736, \8796_9095 );
and \U$3567 ( \12356_12655 , RIfeab8d0_8268, \8798_9097 );
and \U$3568 ( \12357_12656 , RIfcc5bd0_7272, \8800_9099 );
and \U$3569 ( \12358_12657 , RIfc62dc8_6147, \8802_9101 );
and \U$3570 ( \12359_12658 , RIee3e710_5169, \8804_9103 );
and \U$3571 ( \12360_12659 , RIfc9cb18_6805, \8806_9105 );
and \U$3572 ( \12361_12660 , RIee3c820_5147, \8808_9107 );
and \U$3573 ( \12362_12661 , RIee3b470_5133, \8810_9109 );
and \U$3574 ( \12363_12662 , RIee3a390_5121, \8812_9111 );
and \U$3575 ( \12364_12663 , RIe174888_2703, \8814_9113 );
and \U$3576 ( \12365_12664 , RIf170498_5737, \8816_9115 );
and \U$3577 ( \12366_12665 , RIfc68660_6210, \8818_9117 );
and \U$3578 ( \12367_12666 , RIf16e878_5717, \8820_9119 );
and \U$3579 ( \12368_12667 , RIfc6ea38_6281, \8822_9121 );
and \U$3580 ( \12369_12668 , RIfe98d48_8083, \8824_9123 );
and \U$3581 ( \12370_12669 , RIe224d78_4709, \8826_9125 );
and \U$3582 ( \12371_12670 , RIf16c280_5690, \8828_9127 );
and \U$3583 ( \12372_12671 , RIe222078_4677, \8830_9129 );
and \U$3584 ( \12373_12672 , RIf16b308_5679, \8832_9131 );
and \U$3585 ( \12374_12673 , RIe21f378_4645, \8834_9133 );
and \U$3586 ( \12375_12674 , RIe219978_4581, \8836_9135 );
and \U$3587 ( \12376_12675 , RIe216c78_4549, \8838_9137 );
and \U$3588 ( \12377_12676 , RIf16a390_5668, \8840_9139 );
and \U$3589 ( \12378_12677 , RIe213f78_4517, \8842_9141 );
and \U$3590 ( \12379_12678 , RIf169b20_5662, \8844_9143 );
and \U$3591 ( \12380_12679 , RIe211278_4485, \8846_9145 );
and \U$3592 ( \12381_12680 , RIf1681d0_5644, \8848_9147 );
and \U$3593 ( \12382_12681 , RIe20e578_4453, \8850_9149 );
and \U$3594 ( \12383_12682 , RIe20b878_4421, \8852_9151 );
and \U$3595 ( \12384_12683 , RIe208b78_4389, \8854_9153 );
and \U$3596 ( \12385_12684 , RIfcd4ae0_7442, \8856_9155 );
and \U$3597 ( \12386_12685 , RIfc61478_6129, \8858_9157 );
and \U$3598 ( \12387_12686 , RIfeab060_8262, \8860_9159 );
and \U$3599 ( \12388_12687 , RIe201990_4308, \8862_9161 );
and \U$3600 ( \12389_12688 , RIfc70ec8_6307, \8864_9163 );
and \U$3601 ( \12390_12689 , RIfc70928_6303, \8866_9165 );
and \U$3602 ( \12391_12690 , RIfcec528_7711, \8868_9167 );
and \U$3603 ( \12392_12691 , RIfcbe880_7190, \8870_9169 );
and \U$3604 ( \12393_12692 , RIf160d18_5561, \8872_9171 );
and \U$3605 ( \12394_12693 , RIf15ee28_5539, \8874_9173 );
and \U$3606 ( \12395_12694 , RIfe98be0_8082, \8876_9175 );
and \U$3607 ( \12396_12695 , RIfe98eb0_8084, \8878_9177 );
and \U$3608 ( \12397_12696 , RIf15d0a0_5518, \8880_9179 );
and \U$3609 ( \12398_12697 , RIf15bcf0_5504, \8882_9181 );
and \U$3610 ( \12399_12698 , RIfcd4540_7438, \8884_9183 );
and \U$3611 ( \12400_12699 , RIf159e00_5482, \8886_9185 );
or \U$3612 ( \12401_12700 , \12337_12636 , \12338_12637 , \12339_12638 , \12340_12639 , \12341_12640 , \12342_12641 , \12343_12642 , \12344_12643 , \12345_12644 , \12346_12645 , \12347_12646 , \12348_12647 , \12349_12648 , \12350_12649 , \12351_12650 , \12352_12651 , \12353_12652 , \12354_12653 , \12355_12654 , \12356_12655 , \12357_12656 , \12358_12657 , \12359_12658 , \12360_12659 , \12361_12660 , \12362_12661 , \12363_12662 , \12364_12663 , \12365_12664 , \12366_12665 , \12367_12666 , \12368_12667 , \12369_12668 , \12370_12669 , \12371_12670 , \12372_12671 , \12373_12672 , \12374_12673 , \12375_12674 , \12376_12675 , \12377_12676 , \12378_12677 , \12379_12678 , \12380_12679 , \12381_12680 , \12382_12681 , \12383_12682 , \12384_12683 , \12385_12684 , \12386_12685 , \12387_12686 , \12388_12687 , \12389_12688 , \12390_12689 , \12391_12690 , \12392_12691 , \12393_12692 , \12394_12693 , \12395_12694 , \12396_12695 , \12397_12696 , \12398_12697 , \12399_12698 , \12400_12699 );
and \U$3613 ( \12402_12701 , RIf1592c0_5474, \8889_9188 );
and \U$3614 ( \12403_12702 , RIf158078_5461, \8891_9190 );
and \U$3615 ( \12404_12703 , RIfca3a30_6884, \8893_9192 );
and \U$3616 ( \12405_12704 , RIfea7988_8223, \8895_9194 );
and \U$3617 ( \12406_12705 , RIf156728_5443, \8897_9196 );
and \U$3618 ( \12407_12706 , RIf155be8_5435, \8899_9198 );
and \U$3619 ( \12408_12707 , RIf154b08_5423, \8901_9200 );
and \U$3620 ( \12409_12708 , RIfe98a78_8081, \8903_9202 );
and \U$3621 ( \12410_12709 , RIf1538c0_5410, \8905_9204 );
and \U$3622 ( \12411_12710 , RIf1520d8_5393, \8907_9206 );
and \U$3623 ( \12412_12711 , RIf150e90_5380, \8909_9208 );
and \U$3624 ( \12413_12712 , RIe1f43d0_4156, \8911_9210 );
and \U$3625 ( \12414_12713 , RIf14fdb0_5368, \8913_9212 );
and \U$3626 ( \12415_12714 , RIfcd2380_7414, \8915_9214 );
and \U$3627 ( \12416_12715 , RIf14e2f8_5349, \8917_9216 );
and \U$3628 ( \12417_12716 , RIe1ef240_4098, \8919_9218 );
and \U$3629 ( \12418_12717 , RIe1ecae0_4070, \8921_9220 );
and \U$3630 ( \12419_12718 , RIe1e9de0_4038, \8923_9222 );
and \U$3631 ( \12420_12719 , RIe1e70e0_4006, \8925_9224 );
and \U$3632 ( \12421_12720 , RIe1e43e0_3974, \8927_9226 );
and \U$3633 ( \12422_12721 , RIe1e16e0_3942, \8929_9228 );
and \U$3634 ( \12423_12722 , RIe1de9e0_3910, \8931_9230 );
and \U$3635 ( \12424_12723 , RIe1dbce0_3878, \8933_9232 );
and \U$3636 ( \12425_12724 , RIe1d8fe0_3846, \8935_9234 );
and \U$3637 ( \12426_12725 , RIe1d35e0_3782, \8937_9236 );
and \U$3638 ( \12427_12726 , RIe1d08e0_3750, \8939_9238 );
and \U$3639 ( \12428_12727 , RIe1cdbe0_3718, \8941_9240 );
and \U$3640 ( \12429_12728 , RIe1caee0_3686, \8943_9242 );
and \U$3641 ( \12430_12729 , RIe1c81e0_3654, \8945_9244 );
and \U$3642 ( \12431_12730 , RIe1c54e0_3622, \8947_9246 );
and \U$3643 ( \12432_12731 , RIe1c27e0_3590, \8949_9248 );
and \U$3644 ( \12433_12732 , RIe1bfae0_3558, \8951_9250 );
and \U$3645 ( \12434_12733 , RIfc44b70_5804, \8953_9252 );
and \U$3646 ( \12435_12734 , RIf14bd00_5322, \8955_9254 );
and \U$3647 ( \12436_12735 , RIfe992e8_8087, \8957_9256 );
and \U$3648 ( \12437_12736 , RIfe987a8_8079, \8959_9258 );
and \U$3649 ( \12438_12737 , RIf14a950_5308, \8961_9260 );
and \U$3650 ( \12439_12738 , RIf149f78_5301, \8963_9262 );
and \U$3651 ( \12440_12739 , RIfe99180_8086, \8965_9264 );
and \U$3652 ( \12441_12740 , RIfe98640_8078, \8967_9266 );
and \U$3653 ( \12442_12741 , RIf149438_5293, \8969_9268 );
and \U$3654 ( \12443_12742 , RIfcec7f8_7713, \8971_9270 );
and \U$3655 ( \12444_12743 , RIfe984d8_8077, \8973_9272 );
and \U$3656 ( \12445_12744 , RIe1b1b48_3399, \8975_9274 );
and \U$3657 ( \12446_12745 , RIfc4b650_5880, \8977_9276 );
and \U$3658 ( \12447_12746 , RIfcda918_7509, \8979_9278 );
and \U$3659 ( \12448_12747 , RIfe98370_8076, \8981_9280 );
and \U$3660 ( \12449_12748 , RIfe99018_8085, \8983_9282 );
and \U$3661 ( \12450_12749 , RIe1a9e20_3310, \8985_9284 );
and \U$3662 ( \12451_12750 , RIe1a7120_3278, \8987_9286 );
and \U$3663 ( \12452_12751 , RIe1a4420_3246, \8989_9288 );
and \U$3664 ( \12453_12752 , RIe1a1720_3214, \8991_9290 );
and \U$3665 ( \12454_12753 , RIe18dc20_2990, \8993_9292 );
and \U$3666 ( \12455_12754 , RIe17a120_2766, \8995_9294 );
and \U$3667 ( \12456_12755 , RIe227a78_4741, \8997_9296 );
and \U$3668 ( \12457_12756 , RIe21c678_4613, \8999_9298 );
and \U$3669 ( \12458_12757 , RIe205e78_4357, \9001_9300 );
and \U$3670 ( \12459_12758 , RIe1ffed8_4289, \9003_9302 );
and \U$3671 ( \12460_12759 , RIe1f9290_4212, \9005_9304 );
and \U$3672 ( \12461_12760 , RIe1f1dd8_4129, \9007_9306 );
and \U$3673 ( \12462_12761 , RIe1d62e0_3814, \9009_9308 );
and \U$3674 ( \12463_12762 , RIe1bcde0_3526, \9011_9310 );
and \U$3675 ( \12464_12763 , RIe1afc58_3377, \9013_9312 );
and \U$3676 ( \12465_12764 , RIe172290_2676, \9015_9314 );
or \U$3677 ( \12466_12765 , \12402_12701 , \12403_12702 , \12404_12703 , \12405_12704 , \12406_12705 , \12407_12706 , \12408_12707 , \12409_12708 , \12410_12709 , \12411_12710 , \12412_12711 , \12413_12712 , \12414_12713 , \12415_12714 , \12416_12715 , \12417_12716 , \12418_12717 , \12419_12718 , \12420_12719 , \12421_12720 , \12422_12721 , \12423_12722 , \12424_12723 , \12425_12724 , \12426_12725 , \12427_12726 , \12428_12727 , \12429_12728 , \12430_12729 , \12431_12730 , \12432_12731 , \12433_12732 , \12434_12733 , \12435_12734 , \12436_12735 , \12437_12736 , \12438_12737 , \12439_12738 , \12440_12739 , \12441_12740 , \12442_12741 , \12443_12742 , \12444_12743 , \12445_12744 , \12446_12745 , \12447_12746 , \12448_12747 , \12449_12748 , \12450_12749 , \12451_12750 , \12452_12751 , \12453_12752 , \12454_12753 , \12455_12754 , \12456_12755 , \12457_12756 , \12458_12757 , \12459_12758 , \12460_12759 , \12461_12760 , \12462_12761 , \12463_12762 , \12464_12763 , \12465_12764 );
or \U$3678 ( \12467_12766 , \12401_12700 , \12466_12765 );
_DC \g6587/U$1 ( \12468 , \12467_12766 , \9024_9323 );
and g6588_GF_PartitionCandidate( \12469_12768_nG6588 , \12336 , \12468 );
buf \U$3679 ( \12470_12769 , \12469_12768_nG6588 );
and \U$3680 ( \12471_12770 , \12470_12769 , \10389_10691 );
nor \U$3681 ( \12472_12771 , \12204_12503 , \12471_12770 );
xnor \U$3682 ( \12473_12772 , \12472_12771 , \10678_10980 );
not \U$3683 ( \12474_12773 , \12160_12462 );
_DC \g4a07/U$1 ( \12475 , \12335_12634 , \9298_9597 );
_DC \g4a8b/U$1 ( \12476 , \12467_12766 , \9024_9323 );
xor g4a8c_GF_PartitionCandidate( \12477_12776_nG4a8c , \12475 , \12476 );
buf \U$3684 ( \12478_12777 , \12477_12776_nG4a8c );
and \U$3685 ( \12479_12778 , \12158_12460 , \11272_11571 );
not \U$3686 ( \12480_12779 , \12479_12778 );
and \U$3687 ( \12481_12780 , \12478_12777 , \12480_12779 );
and \U$3688 ( \12482_12781 , \12474_12773 , \12481_12780 );
xor \U$3689 ( \12483_12782 , \12473_12772 , \12482_12781 );
and \U$3690 ( \12484_12783 , \10968_11270 , \11275_11574 );
and \U$3691 ( \12485_12784 , \11287_11586 , \10976_11278 );
nor \U$3692 ( \12486_12785 , \12484_12783 , \12485_12784 );
xnor \U$3693 ( \12487_12786 , \12486_12785 , \11281_11580 );
xor \U$3694 ( \12488_12787 , \12483_12782 , \12487_12786 );
xor \U$3695 ( \12489_12788 , \12478_12777 , \12158_12460 );
not \U$3696 ( \12490_12789 , \12159_12461 );
and \U$3697 ( \12491_12790 , \12489_12788 , \12490_12789 );
and \U$3698 ( \12492_12791 , \10385_10687 , \12491_12790 );
and \U$3699 ( \12493_12792 , \10686_10988 , \12159_12461 );
nor \U$3700 ( \12494_12793 , \12492_12791 , \12493_12792 );
xnor \U$3701 ( \12495_12794 , \12494_12793 , \12481_12780 );
xor \U$3702 ( \12496_12795 , \12488_12787 , \12495_12794 );
xor \U$3703 ( \12497_12796 , \12203_12502 , \12496_12795 );
and \U$3704 ( \12498_12797 , \12161_12463 , \12162_12464 );
and \U$3705 ( \12499_12798 , \12163_12465 , \12166_12468 );
or \U$3706 ( \12500_12799 , \12498_12797 , \12499_12798 );
xor \U$3707 ( \12501_12800 , \12497_12796 , \12500_12799 );
buf g9bff_GF_PartitionCandidate( \12502_12801_nG9bff , \12501_12800 );
and \U$3708 ( \12503_12802 , \10402_10704 , \12502_12801_nG9bff );
or \U$3709 ( \12504_12803 , \12199_12498 , \12503_12802 );
xor \U$3710 ( \12505_12804 , \10399_10703 , \12504_12803 );
buf \U$3711 ( \12506_12805 , \12505_12804 );
buf \U$3713 ( \12507_12806 , \12506_12805 );
xor \U$3714 ( \12508_12807 , \12198_12497 , \12507_12806 );
buf \U$3715 ( \12509_12808 , \12508_12807 );
and \U$3716 ( \12510_12809 , \11872_12174 , \11877_12179 );
and \U$3717 ( \12511_12810 , \11872_12174 , \12173_12475 );
and \U$3718 ( \12512_12811 , \11877_12179 , \12173_12475 );
or \U$3719 ( \12513_12812 , \12510_12809 , \12511_12810 , \12512_12811 );
buf \U$3720 ( \12514_12813 , \12513_12812 );
xor \U$3721 ( \12515_12814 , \12509_12808 , \12514_12813 );
and \U$3722 ( \12516_12815 , \11864_12166 , \11870_12172 );
buf \U$3723 ( \12517_12816 , \12516_12815 );
xor \U$3724 ( \12518_12817 , \12515_12814 , \12517_12816 );
and \U$3725 ( \12519_12818 , \12177_12479 , \12518_12817 );
and \U$3726 ( \12520_12819 , RIdec6a58_724, \8760_9059 );
and \U$3727 ( \12521_12820 , RIdec3d58_692, \8762_9061 );
and \U$3728 ( \12522_12821 , RIfc723e0_6322, \8764_9063 );
and \U$3729 ( \12523_12822 , RIdec1058_660, \8766_9065 );
and \U$3730 ( \12524_12823 , RIfc59fc0_6046, \8768_9067 );
and \U$3731 ( \12525_12824 , RIdebe358_628, \8770_9069 );
and \U$3732 ( \12526_12825 , RIdebb658_596, \8772_9071 );
and \U$3733 ( \12527_12826 , RIdeb8958_564, \8774_9073 );
and \U$3734 ( \12528_12827 , RIfcb96f0_7132, \8776_9075 );
and \U$3735 ( \12529_12828 , RIdeb2f58_500, \8778_9077 );
and \U$3736 ( \12530_12829 , RIfce1c68_7591, \8780_9079 );
and \U$3737 ( \12531_12830 , RIdeb0258_468, \8782_9081 );
and \U$3738 ( \12532_12831 , RIfc9b498_6789, \8784_9083 );
and \U$3739 ( \12533_12832 , RIdead558_436, \8786_9085 );
and \U$3740 ( \12534_12833 , RIdea6fa0_404, \8788_9087 );
and \U$3741 ( \12535_12834 , RIdea06a0_372, \8790_9089 );
and \U$3742 ( \12536_12835 , RIfc81458_6493, \8792_9091 );
and \U$3743 ( \12537_12836 , RIfc83780_6518, \8794_9093 );
and \U$3744 ( \12538_12837 , RIfc4e620_5914, \8796_9095 );
and \U$3745 ( \12539_12838 , RIfcd3e38_7433, \8798_9097 );
and \U$3746 ( \12540_12839 , RIde937e8_309, \8800_9099 );
and \U$3747 ( \12541_12840 , RIde8f990_290, \8802_9101 );
and \U$3748 ( \12542_12841 , RIde8bb38_271, \8804_9103 );
and \U$3749 ( \12543_12842 , RIde87650_250, \8806_9105 );
and \U$3750 ( \12544_12843 , RIde834b0_230, \8808_9107 );
and \U$3751 ( \12545_12844 , RIfc42c80_5782, \8810_9109 );
and \U$3752 ( \12546_12845 , RIfc65960_6178, \8812_9111 );
and \U$3753 ( \12547_12846 , RIfc6c710_6256, \8814_9113 );
and \U$3754 ( \12548_12847 , RIee392b0_5109, \8816_9115 );
and \U$3755 ( \12549_12848 , RIe16cb60_2614, \8818_9117 );
and \U$3756 ( \12550_12849 , RIe16a6d0_2588, \8820_9119 );
and \U$3757 ( \12551_12850 , RIe169050_2572, \8822_9121 );
and \U$3758 ( \12552_12851 , RIe166a58_2545, \8824_9123 );
and \U$3759 ( \12553_12852 , RIe163d58_2513, \8826_9125 );
and \U$3760 ( \12554_12853 , RIfec3cf0_8348, \8828_9127 );
and \U$3761 ( \12555_12854 , RIe161058_2481, \8830_9129 );
and \U$3762 ( \12556_12855 , RIfcd54b8_7449, \8832_9131 );
and \U$3763 ( \12557_12856 , RIe15e358_2449, \8834_9133 );
and \U$3764 ( \12558_12857 , RIe158958_2385, \8836_9135 );
and \U$3765 ( \12559_12858 , RIe155c58_2353, \8838_9137 );
and \U$3766 ( \12560_12859 , RIfe9ba48_8115, \8840_9139 );
and \U$3767 ( \12561_12860 , RIe152f58_2321, \8842_9141 );
and \U$3768 ( \12562_12861 , RIfec4128_8351, \8844_9143 );
and \U$3769 ( \12563_12862 , RIe150258_2289, \8846_9145 );
and \U$3770 ( \12564_12863 , RIfcb9b28_7135, \8848_9147 );
and \U$3771 ( \12565_12864 , RIe14d558_2257, \8850_9149 );
and \U$3772 ( \12566_12865 , RIe14a858_2225, \8852_9151 );
and \U$3773 ( \12567_12866 , RIe147b58_2193, \8854_9153 );
and \U$3774 ( \12568_12867 , RIfcdb2f0_7516, \8856_9155 );
and \U$3775 ( \12569_12868 , RIfc553d0_5992, \8858_9157 );
and \U$3776 ( \12570_12869 , RIfc9a0e8_6775, \8860_9159 );
and \U$3777 ( \12571_12870 , RIfcbd908_7179, \8862_9161 );
and \U$3778 ( \12572_12871 , RIe1422c0_2130, \8864_9163 );
and \U$3779 ( \12573_12872 , RIe13ff98_2105, \8866_9165 );
and \U$3780 ( \12574_12873 , RIdf3dea0_2081, \8868_9167 );
and \U$3781 ( \12575_12874 , RIdf3ba10_2055, \8870_9169 );
and \U$3782 ( \12576_12875 , RIfc87128_6559, \8872_9171 );
and \U$3783 ( \12577_12876 , RIee304a8_5008, \8874_9173 );
and \U$3784 ( \12578_12877 , RIfcc51f8_7265, \8876_9175 );
and \U$3785 ( \12579_12878 , RIee2e2e8_4984, \8878_9177 );
and \U$3786 ( \12580_12879 , RIdf36cb8_2000, \8880_9179 );
and \U$3787 ( \12581_12880 , RIfec3fc0_8350, \8882_9181 );
and \U$3788 ( \12582_12881 , RIdf32500_1949, \8884_9183 );
and \U$3789 ( \12583_12882 , RIfec3e58_8349, \8886_9185 );
or \U$3790 ( \12584_12883 , \12520_12819 , \12521_12820 , \12522_12821 , \12523_12822 , \12524_12823 , \12525_12824 , \12526_12825 , \12527_12826 , \12528_12827 , \12529_12828 , \12530_12829 , \12531_12830 , \12532_12831 , \12533_12832 , \12534_12833 , \12535_12834 , \12536_12835 , \12537_12836 , \12538_12837 , \12539_12838 , \12540_12839 , \12541_12840 , \12542_12841 , \12543_12842 , \12544_12843 , \12545_12844 , \12546_12845 , \12547_12846 , \12548_12847 , \12549_12848 , \12550_12849 , \12551_12850 , \12552_12851 , \12553_12852 , \12554_12853 , \12555_12854 , \12556_12855 , \12557_12856 , \12558_12857 , \12559_12858 , \12560_12859 , \12561_12860 , \12562_12861 , \12563_12862 , \12564_12863 , \12565_12864 , \12566_12865 , \12567_12866 , \12568_12867 , \12569_12868 , \12570_12869 , \12571_12870 , \12572_12871 , \12573_12872 , \12574_12873 , \12575_12874 , \12576_12875 , \12577_12876 , \12578_12877 , \12579_12878 , \12580_12879 , \12581_12880 , \12582_12881 , \12583_12882 );
and \U$3791 ( \12585_12884 , RIee2c830_4965, \8889_9188 );
and \U$3792 ( \12586_12885 , RIee2ad78_4946, \8891_9190 );
and \U$3793 ( \12587_12886 , RIee296f8_4930, \8893_9192 );
and \U$3794 ( \12588_12887 , RIee284b0_4917, \8895_9194 );
and \U$3795 ( \12589_12888 , RIfe9b8e0_8114, \8897_9196 );
and \U$3796 ( \12590_12889 , RIfe9b610_8112, \8899_9198 );
and \U$3797 ( \12591_12890 , RIfe9b778_8113, \8901_9200 );
and \U$3798 ( \12592_12891 , RIfe9b4a8_8111, \8903_9202 );
and \U$3799 ( \12593_12892 , RIfcb7c38_7113, \8905_9204 );
and \U$3800 ( \12594_12893 , RIfc86b88_6555, \8907_9206 );
and \U$3801 ( \12595_12894 , RIdf238c0_1781, \8909_9208 );
and \U$3802 ( \12596_12895 , RIfc75ab8_6361, \8911_9210 );
and \U$3803 ( \12597_12896 , RIdf22240_1765, \8913_9212 );
and \U$3804 ( \12598_12897 , RIfeaa3b8_8253, \8915_9214 );
and \U$3805 ( \12599_12898 , RIdf1bb98_1692, \8917_9216 );
and \U$3806 ( \12600_12899 , RIdf1a680_1677, \8919_9218 );
and \U$3807 ( \12601_12900 , RIdf18628_1654, \8921_9220 );
and \U$3808 ( \12602_12901 , RIdf15928_1622, \8923_9222 );
and \U$3809 ( \12603_12902 , RIdf12c28_1590, \8925_9224 );
and \U$3810 ( \12604_12903 , RIdf0ff28_1558, \8927_9226 );
and \U$3811 ( \12605_12904 , RIdf0d228_1526, \8929_9228 );
and \U$3812 ( \12606_12905 , RIdf0a528_1494, \8931_9230 );
and \U$3813 ( \12607_12906 , RIdf07828_1462, \8933_9232 );
and \U$3814 ( \12608_12907 , RIdf04b28_1430, \8935_9234 );
and \U$3815 ( \12609_12908 , RIdeff128_1366, \8937_9236 );
and \U$3816 ( \12610_12909 , RIdefc428_1334, \8939_9238 );
and \U$3817 ( \12611_12910 , RIdef9728_1302, \8941_9240 );
and \U$3818 ( \12612_12911 , RIdef6a28_1270, \8943_9242 );
and \U$3819 ( \12613_12912 , RIdef3d28_1238, \8945_9244 );
and \U$3820 ( \12614_12913 , RIdef1028_1206, \8947_9246 );
and \U$3821 ( \12615_12914 , RIdeee328_1174, \8949_9248 );
and \U$3822 ( \12616_12915 , RIdeeb628_1142, \8951_9250 );
and \U$3823 ( \12617_12916 , RIee25a80_4887, \8953_9252 );
and \U$3824 ( \12618_12917 , RIee24c70_4877, \8955_9254 );
and \U$3825 ( \12619_12918 , RIfcddd20_7546, \8957_9256 );
and \U$3826 ( \12620_12919 , RIfccc110_7344, \8959_9258 );
and \U$3827 ( \12621_12920 , RIdee5c28_1078, \8961_9260 );
and \U$3828 ( \12622_12921 , RIdee3ea0_1057, \8963_9262 );
and \U$3829 ( \12623_12922 , RIdee1b78_1032, \8965_9264 );
and \U$3830 ( \12624_12923 , RIdedfc88_1010, \8967_9266 );
and \U$3831 ( \12625_12924 , RIfc6a6b8_6233, \8969_9268 );
and \U$3832 ( \12626_12925 , RIee227e0_4851, \8971_9270 );
and \U$3833 ( \12627_12926 , RIfc88be0_6578, \8973_9272 );
and \U$3834 ( \12628_12927 , RIee21868_4840, \8975_9274 );
and \U$3835 ( \12629_12928 , RIdedaaf8_952, \8977_9276 );
and \U$3836 ( \12630_12929 , RIded8668_926, \8979_9278 );
and \U$3837 ( \12631_12930 , RIded6340_901, \8981_9280 );
and \U$3838 ( \12632_12931 , RIded4180_877, \8983_9282 );
and \U$3839 ( \12633_12932 , RIded1e58_852, \8985_9284 );
and \U$3840 ( \12634_12933 , RIdecf158_820, \8987_9286 );
and \U$3841 ( \12635_12934 , RIdecc458_788, \8989_9288 );
and \U$3842 ( \12636_12935 , RIdec9758_756, \8991_9290 );
and \U$3843 ( \12637_12936 , RIdeb5c58_532, \8993_9292 );
and \U$3844 ( \12638_12937 , RIde99da0_340, \8995_9294 );
and \U$3845 ( \12639_12938 , RIe16f860_2646, \8997_9296 );
and \U$3846 ( \12640_12939 , RIe15b658_2417, \8999_9298 );
and \U$3847 ( \12641_12940 , RIe144e58_2161, \9001_9300 );
and \U$3848 ( \12642_12941 , RIdf39850_2031, \9003_9302 );
and \U$3849 ( \12643_12942 , RIdf2deb0_1899, \9005_9304 );
and \U$3850 ( \12644_12943 , RIdf1e730_1723, \9007_9306 );
and \U$3851 ( \12645_12944 , RIdf01e28_1398, \9009_9308 );
and \U$3852 ( \12646_12945 , RIdee8928_1110, \9011_9310 );
and \U$3853 ( \12647_12946 , RIdedd690_983, \9013_9312 );
and \U$3854 ( \12648_12947 , RIde7fce8_213, \9015_9314 );
or \U$3855 ( \12649_12948 , \12585_12884 , \12586_12885 , \12587_12886 , \12588_12887 , \12589_12888 , \12590_12889 , \12591_12890 , \12592_12891 , \12593_12892 , \12594_12893 , \12595_12894 , \12596_12895 , \12597_12896 , \12598_12897 , \12599_12898 , \12600_12899 , \12601_12900 , \12602_12901 , \12603_12902 , \12604_12903 , \12605_12904 , \12606_12905 , \12607_12906 , \12608_12907 , \12609_12908 , \12610_12909 , \12611_12910 , \12612_12911 , \12613_12912 , \12614_12913 , \12615_12914 , \12616_12915 , \12617_12916 , \12618_12917 , \12619_12918 , \12620_12919 , \12621_12920 , \12622_12921 , \12623_12922 , \12624_12923 , \12625_12924 , \12626_12925 , \12627_12926 , \12628_12927 , \12629_12928 , \12630_12929 , \12631_12930 , \12632_12931 , \12633_12932 , \12634_12933 , \12635_12934 , \12636_12935 , \12637_12936 , \12638_12937 , \12639_12938 , \12640_12939 , \12641_12940 , \12642_12941 , \12643_12942 , \12644_12943 , \12645_12944 , \12646_12945 , \12647_12946 , \12648_12947 );
or \U$3856 ( \12650_12949 , \12584_12883 , \12649_12948 );
_DC \g2ead/U$1 ( \12651 , \12650_12949 , \9024_9323 );
buf \U$3857 ( \12652_12951 , \12651 );
and \U$3858 ( \12653_12952 , RIe19ecf0_3184, \9034_9333 );
and \U$3859 ( \12654_12953 , RIe19bff0_3152, \9036_9335 );
and \U$3860 ( \12655_12954 , RIf145a90_5252, \9038_9337 );
and \U$3861 ( \12656_12955 , RIe1992f0_3120, \9040_9339 );
and \U$3862 ( \12657_12956 , RIf144de8_5243, \9042_9341 );
and \U$3863 ( \12658_12957 , RIe1965f0_3088, \9044_9343 );
and \U$3864 ( \12659_12958 , RIe1938f0_3056, \9046_9345 );
and \U$3865 ( \12660_12959 , RIe190bf0_3024, \9048_9347 );
and \U$3866 ( \12661_12960 , RIe18b1f0_2960, \9050_9349 );
and \U$3867 ( \12662_12961 , RIe1884f0_2928, \9052_9351 );
and \U$3868 ( \12663_12962 , RIfc72980_6326, \9054_9353 );
and \U$3869 ( \12664_12963 , RIe1857f0_2896, \9056_9355 );
and \U$3870 ( \12665_12964 , RIf143060_5222, \9058_9357 );
and \U$3871 ( \12666_12965 , RIe182af0_2864, \9060_9359 );
and \U$3872 ( \12667_12966 , RIe17fdf0_2832, \9062_9361 );
and \U$3873 ( \12668_12967 , RIe17d0f0_2800, \9064_9363 );
and \U$3874 ( \12669_12968 , RIf142688_5215, \9066_9365 );
and \U$3875 ( \12670_12969 , RIf141710_5204, \9068_9367 );
and \U$3876 ( \12671_12970 , RIe177858_2737, \9070_9369 );
and \U$3877 ( \12672_12971 , RIe176778_2725, \9072_9371 );
and \U$3878 ( \12673_12972 , RIfcea638_7689, \9074_9373 );
and \U$3879 ( \12674_12973 , RIfca54e8_6903, \9076_9375 );
and \U$3880 ( \12675_12974 , RIee3e878_5170, \9078_9377 );
and \U$3881 ( \12676_12975 , RIee3dbd0_5161, \9080_9379 );
and \U$3882 ( \12677_12976 , RIee3c988_5148, \9082_9381 );
and \U$3883 ( \12678_12977 , RIee3b5d8_5134, \9084_9383 );
and \U$3884 ( \12679_12978 , RIee3a4f8_5122, \9086_9385 );
and \U$3885 ( \12680_12979 , RIe174b58_2705, \9088_9387 );
and \U$3886 ( \12681_12980 , RIf170600_5738, \9090_9389 );
and \U$3887 ( \12682_12981 , RIfc76fd0_6376, \9092_9391 );
and \U$3888 ( \12683_12982 , RIf16e9e0_5718, \9094_9393 );
and \U$3889 ( \12684_12983 , RIfced608_7723, \9096_9395 );
and \U$3890 ( \12685_12984 , RIf16d090_5700, \9098_9397 );
and \U$3891 ( \12686_12985 , RIe225048_4711, \9100_9399 );
and \U$3892 ( \12687_12986 , RIf16c550_5692, \9102_9401 );
and \U$3893 ( \12688_12987 , RIe222348_4679, \9104_9403 );
and \U$3894 ( \12689_12988 , RIf16b470_5680, \9106_9405 );
and \U$3895 ( \12690_12989 , RIe21f648_4647, \9108_9407 );
and \U$3896 ( \12691_12990 , RIe219c48_4583, \9110_9409 );
and \U$3897 ( \12692_12991 , RIe216f48_4551, \9112_9411 );
and \U$3898 ( \12693_12992 , RIf16a4f8_5669, \9114_9413 );
and \U$3899 ( \12694_12993 , RIe214248_4519, \9116_9415 );
and \U$3900 ( \12695_12994 , RIf169df0_5664, \9118_9417 );
and \U$3901 ( \12696_12995 , RIe211548_4487, \9120_9419 );
and \U$3902 ( \12697_12996 , RIf1684a0_5646, \9122_9421 );
and \U$3903 ( \12698_12997 , RIe20e848_4455, \9124_9423 );
and \U$3904 ( \12699_12998 , RIe20bb48_4423, \9126_9425 );
and \U$3905 ( \12700_12999 , RIe208e48_4391, \9128_9427 );
and \U$3906 ( \12701_13000 , RIf1673c0_5634, \9130_9429 );
and \U$3907 ( \12702_13001 , RIf166448_5623, \9132_9431 );
and \U$3908 ( \12703_13002 , RIfe9c6f0_8124, \9134_9433 );
and \U$3909 ( \12704_13003 , RIfe9c150_8120, \9136_9435 );
and \U$3910 ( \12705_13004 , RIf1654d0_5612, \9138_9437 );
and \U$3911 ( \12706_13005 , RIfcc4550_7256, \9140_9439 );
and \U$3912 ( \12707_13006 , RIf1635e0_5590, \9142_9441 );
and \U$3913 ( \12708_13007 , RIf162500_5578, \9144_9443 );
and \U$3914 ( \12709_13008 , RIf160fe8_5563, \9146_9445 );
and \U$3915 ( \12710_13009 , RIf15f0f8_5541, \9148_9447 );
and \U$3916 ( \12711_13010 , RIfe9bfe8_8119, \9150_9449 );
and \U$3917 ( \12712_13011 , RIfe9c588_8123, \9152_9451 );
and \U$3918 ( \12713_13012 , RIf15d208_5519, \9154_9453 );
and \U$3919 ( \12714_13013 , RIf15bfc0_5506, \9156_9455 );
and \U$3920 ( \12715_13014 , RIfc4d540_5902, \9158_9457 );
and \U$3921 ( \12716_13015 , RIfc9c848_6803, \9160_9459 );
or \U$3922 ( \12717_13016 , \12653_12952 , \12654_12953 , \12655_12954 , \12656_12955 , \12657_12956 , \12658_12957 , \12659_12958 , \12660_12959 , \12661_12960 , \12662_12961 , \12663_12962 , \12664_12963 , \12665_12964 , \12666_12965 , \12667_12966 , \12668_12967 , \12669_12968 , \12670_12969 , \12671_12970 , \12672_12971 , \12673_12972 , \12674_12973 , \12675_12974 , \12676_12975 , \12677_12976 , \12678_12977 , \12679_12978 , \12680_12979 , \12681_12980 , \12682_12981 , \12683_12982 , \12684_12983 , \12685_12984 , \12686_12985 , \12687_12986 , \12688_12987 , \12689_12988 , \12690_12989 , \12691_12990 , \12692_12991 , \12693_12992 , \12694_12993 , \12695_12994 , \12696_12995 , \12697_12996 , \12698_12997 , \12699_12998 , \12700_12999 , \12701_13000 , \12702_13001 , \12703_13002 , \12704_13003 , \12705_13004 , \12706_13005 , \12707_13006 , \12708_13007 , \12709_13008 , \12710_13009 , \12711_13010 , \12712_13011 , \12713_13012 , \12714_13013 , \12715_13014 , \12716_13015 );
and \U$3923 ( \12718_13017 , RIfec4290_8352, \9163_9462 );
and \U$3924 ( \12719_13018 , RIfe9c2b8_8121, \9165_9464 );
and \U$3925 ( \12720_13019 , RIfcc01d0_7208, \9167_9466 );
and \U$3926 ( \12721_13020 , RIe1fb2e8_4235, \9169_9468 );
and \U$3927 ( \12722_13021 , RIfe9c420_8122, \9171_9470 );
and \U$3928 ( \12723_13022 , RIfca3e68_6887, \9173_9472 );
and \U$3929 ( \12724_13023 , RIf154c70_5424, \9175_9474 );
and \U$3930 ( \12725_13024 , RIe1f69c8_4183, \9177_9476 );
and \U$3931 ( \12726_13025 , RIf153a28_5411, \9179_9478 );
and \U$3932 ( \12727_13026 , RIf152240_5394, \9181_9480 );
and \U$3933 ( \12728_13027 , RIf150ff8_5381, \9183_9482 );
and \U$3934 ( \12729_13028 , RIe1f46a0_4158, \9185_9484 );
and \U$3935 ( \12730_13029 , RIfca6028_6911, \9187_9486 );
and \U$3936 ( \12731_13030 , RIfc43bf8_5793, \9189_9488 );
and \U$3937 ( \12732_13031 , RIf14e460_5350, \9191_9490 );
and \U$3938 ( \12733_13032 , RIe1ef3a8_4099, \9193_9492 );
and \U$3939 ( \12734_13033 , RIe1ecdb0_4072, \9195_9494 );
and \U$3940 ( \12735_13034 , RIe1ea0b0_4040, \9197_9496 );
and \U$3941 ( \12736_13035 , RIe1e73b0_4008, \9199_9498 );
and \U$3942 ( \12737_13036 , RIe1e46b0_3976, \9201_9500 );
and \U$3943 ( \12738_13037 , RIe1e19b0_3944, \9203_9502 );
and \U$3944 ( \12739_13038 , RIe1decb0_3912, \9205_9504 );
and \U$3945 ( \12740_13039 , RIe1dbfb0_3880, \9207_9506 );
and \U$3946 ( \12741_13040 , RIe1d92b0_3848, \9209_9508 );
and \U$3947 ( \12742_13041 , RIe1d38b0_3784, \9211_9510 );
and \U$3948 ( \12743_13042 , RIe1d0bb0_3752, \9213_9512 );
and \U$3949 ( \12744_13043 , RIe1cdeb0_3720, \9215_9514 );
and \U$3950 ( \12745_13044 , RIe1cb1b0_3688, \9217_9516 );
and \U$3951 ( \12746_13045 , RIe1c84b0_3656, \9219_9518 );
and \U$3952 ( \12747_13046 , RIe1c57b0_3624, \9221_9520 );
and \U$3953 ( \12748_13047 , RIe1c2ab0_3592, \9223_9522 );
and \U$3954 ( \12749_13048 , RIe1bfdb0_3560, \9225_9524 );
and \U$3955 ( \12750_13049 , RIfc4d6a8_5903, \9227_9526 );
and \U$3956 ( \12751_13050 , RIf14be68_5323, \9229_9528 );
and \U$3957 ( \12752_13051 , RIe1ba680_3498, \9231_9530 );
and \U$3958 ( \12753_13052 , RIfe9be80_8118, \9233_9532 );
and \U$3959 ( \12754_13053 , RIfc86e58_6557, \9235_9534 );
and \U$3960 ( \12755_13054 , RIfcd46a8_7439, \9237_9536 );
and \U$3961 ( \12756_13055 , RIe1b6300_3450, \9239_9538 );
and \U$3962 ( \12757_13056 , RIfe9bd18_8117, \9241_9540 );
and \U$3963 ( \12758_13057 , RIf1495a0_5294, \9243_9542 );
and \U$3964 ( \12759_13058 , RIf1481f0_5280, \9245_9544 );
and \U$3965 ( \12760_13059 , RIe1b3600_3418, \9247_9546 );
and \U$3966 ( \12761_13060 , RIe1b1e18_3401, \9249_9548 );
and \U$3967 ( \12762_13061 , RIfc69470_6220, \9251_9550 );
and \U$3968 ( \12763_13062 , RIfcbfac8_7203, \9253_9552 );
and \U$3969 ( \12764_13063 , RIfe9bbb0_8116, \9255_9554 );
and \U$3970 ( \12765_13064 , RIe1abd10_3332, \9257_9556 );
and \U$3971 ( \12766_13065 , RIe1aa0f0_3312, \9259_9558 );
and \U$3972 ( \12767_13066 , RIe1a73f0_3280, \9261_9560 );
and \U$3973 ( \12768_13067 , RIe1a46f0_3248, \9263_9562 );
and \U$3974 ( \12769_13068 , RIe1a19f0_3216, \9265_9564 );
and \U$3975 ( \12770_13069 , RIe18def0_2992, \9267_9566 );
and \U$3976 ( \12771_13070 , RIe17a3f0_2768, \9269_9568 );
and \U$3977 ( \12772_13071 , RIe227d48_4743, \9271_9570 );
and \U$3978 ( \12773_13072 , RIe21c948_4615, \9273_9572 );
and \U$3979 ( \12774_13073 , RIe206148_4359, \9275_9574 );
and \U$3980 ( \12775_13074 , RIe2001a8_4291, \9277_9576 );
and \U$3981 ( \12776_13075 , RIe1f9560_4214, \9279_9578 );
and \U$3982 ( \12777_13076 , RIe1f20a8_4131, \9281_9580 );
and \U$3983 ( \12778_13077 , RIe1d65b0_3816, \9283_9582 );
and \U$3984 ( \12779_13078 , RIe1bd0b0_3528, \9285_9584 );
and \U$3985 ( \12780_13079 , RIe1aff28_3379, \9287_9586 );
and \U$3986 ( \12781_13080 , RIe172560_2678, \9289_9588 );
or \U$3987 ( \12782_13081 , \12718_13017 , \12719_13018 , \12720_13019 , \12721_13020 , \12722_13021 , \12723_13022 , \12724_13023 , \12725_13024 , \12726_13025 , \12727_13026 , \12728_13027 , \12729_13028 , \12730_13029 , \12731_13030 , \12732_13031 , \12733_13032 , \12734_13033 , \12735_13034 , \12736_13035 , \12737_13036 , \12738_13037 , \12739_13038 , \12740_13039 , \12741_13040 , \12742_13041 , \12743_13042 , \12744_13043 , \12745_13044 , \12746_13045 , \12747_13046 , \12748_13047 , \12749_13048 , \12750_13049 , \12751_13050 , \12752_13051 , \12753_13052 , \12754_13053 , \12755_13054 , \12756_13055 , \12757_13056 , \12758_13057 , \12759_13058 , \12760_13059 , \12761_13060 , \12762_13061 , \12763_13062 , \12764_13063 , \12765_13064 , \12766_13065 , \12767_13066 , \12768_13067 , \12769_13068 , \12770_13069 , \12771_13070 , \12772_13071 , \12773_13072 , \12774_13073 , \12775_13074 , \12776_13075 , \12777_13076 , \12778_13077 , \12779_13078 , \12780_13079 , \12781_13080 );
or \U$3988 ( \12783_13082 , \12717_13016 , \12782_13081 );
_DC \g3fda/U$1 ( \12784 , \12783_13082 , \9298_9597 );
buf \U$3989 ( \12785_13084 , \12784 );
xor \U$3990 ( \12786_13085 , \12652_12951 , \12785_13084 );
and \U$3991 ( \12787_13086 , RIdec68f0_723, \8760_9059 );
and \U$3992 ( \12788_13087 , RIdec3bf0_691, \8762_9061 );
and \U$3993 ( \12789_13088 , RIee208f0_4829, \8764_9063 );
and \U$3994 ( \12790_13089 , RIdec0ef0_659, \8766_9065 );
and \U$3995 ( \12791_13090 , RIfc7ce08_6443, \8768_9067 );
and \U$3996 ( \12792_13091 , RIdebe1f0_627, \8770_9069 );
and \U$3997 ( \12793_13092 , RIdebb4f0_595, \8772_9071 );
and \U$3998 ( \12794_13093 , RIdeb87f0_563, \8774_9073 );
and \U$3999 ( \12795_13094 , RIfc9b8d0_6792, \8776_9075 );
and \U$4000 ( \12796_13095 , RIdeb2df0_499, \8778_9077 );
and \U$4001 ( \12797_13096 , RIfcc6710_7280, \8780_9079 );
and \U$4002 ( \12798_13097 , RIdeb00f0_467, \8782_9081 );
and \U$4003 ( \12799_13098 , RIfc5ff60_6114, \8784_9083 );
and \U$4004 ( \12800_13099 , RIdead3f0_435, \8786_9085 );
and \U$4005 ( \12801_13100 , RIdea6c58_403, \8788_9087 );
and \U$4006 ( \12802_13101 , RIdea0358_371, \8790_9089 );
and \U$4007 ( \12803_13102 , RIfce5070_7628, \8792_9091 );
and \U$4008 ( \12804_13103 , RIee1c6d8_4782, \8794_9093 );
and \U$4009 ( \12805_13104 , RIfce70c8_7651, \8796_9095 );
and \U$4010 ( \12806_13105 , RIee1b058_4766, \8798_9097 );
and \U$4011 ( \12807_13106 , RIde934a0_308, \8800_9099 );
and \U$4012 ( \12808_13107 , RIfe9b1d8_8109, \8802_9101 );
and \U$4013 ( \12809_13108 , RIde8b7f0_270, \8804_9103 );
and \U$4014 ( \12810_13109 , RIfe9b340_8110, \8806_9105 );
and \U$4015 ( \12811_13110 , RIfc6b798_6245, \8808_9107 );
and \U$4016 ( \12812_13111 , RIfcb2238_7049, \8810_9109 );
and \U$4017 ( \12813_13112 , RIfcd3a00_7430, \8812_9111 );
and \U$4018 ( \12814_13113 , RIfcdb020_7514, \8814_9113 );
and \U$4019 ( \12815_13114 , RIfc511b8_5945, \8816_9115 );
and \U$4020 ( \12816_13115 , RIe16c9f8_2613, \8818_9117 );
and \U$4021 ( \12817_13116 , RIfcb27d8_7053, \8820_9119 );
and \U$4022 ( \12818_13117 , RIe168ee8_2571, \8822_9121 );
and \U$4023 ( \12819_13118 , RIe1668f0_2544, \8824_9123 );
and \U$4024 ( \12820_13119 , RIe163bf0_2512, \8826_9125 );
and \U$4025 ( \12821_13120 , RIee381d0_5097, \8828_9127 );
and \U$4026 ( \12822_13121 , RIe160ef0_2480, \8830_9129 );
and \U$4027 ( \12823_13122 , RIfcdfaa8_7567, \8832_9131 );
and \U$4028 ( \12824_13123 , RIe15e1f0_2448, \8834_9133 );
and \U$4029 ( \12825_13124 , RIe1587f0_2384, \8836_9135 );
and \U$4030 ( \12826_13125 , RIe155af0_2352, \8838_9137 );
and \U$4031 ( \12827_13126 , RIfc3f968_5749, \8840_9139 );
and \U$4032 ( \12828_13127 , RIe152df0_2320, \8842_9141 );
and \U$4033 ( \12829_13128 , RIfcd5080_7446, \8844_9143 );
and \U$4034 ( \12830_13129 , RIe1500f0_2288, \8846_9145 );
and \U$4035 ( \12831_13130 , RIfc84b30_6532, \8848_9147 );
and \U$4036 ( \12832_13131 , RIe14d3f0_2256, \8850_9149 );
and \U$4037 ( \12833_13132 , RIe14a6f0_2224, \8852_9151 );
and \U$4038 ( \12834_13133 , RIe1479f0_2192, \8854_9153 );
and \U$4039 ( \12835_13134 , RIfcea098_7685, \8856_9155 );
and \U$4040 ( \12836_13135 , RIfc92f00_6694, \8858_9157 );
and \U$4041 ( \12837_13136 , RIfc54890_5984, \8860_9159 );
and \U$4042 ( \12838_13137 , RIfcdcc40_7534, \8862_9161 );
and \U$4043 ( \12839_13138 , RIe142158_2129, \8864_9163 );
and \U$4044 ( \12840_13139 , RIe13fe30_2104, \8866_9165 );
and \U$4045 ( \12841_13140 , RIdf3dd38_2080, \8868_9167 );
and \U$4046 ( \12842_13141 , RIdf3b8a8_2054, \8870_9169 );
and \U$4047 ( \12843_13142 , RIfc57590_6016, \8872_9171 );
and \U$4048 ( \12844_13143 , RIee30340_5007, \8874_9173 );
and \U$4049 ( \12845_13144 , RIfcd0490_7392, \8876_9175 );
and \U$4050 ( \12846_13145 , RIee2e180_4983, \8878_9177 );
and \U$4051 ( \12847_13146 , RIdf36b50_1999, \8880_9179 );
and \U$4052 ( \12848_13147 , RIdf34558_1972, \8882_9181 );
and \U$4053 ( \12849_13148 , RIdf32398_1948, \8884_9183 );
and \U$4054 ( \12850_13149 , RIfe9b070_8108, \8886_9185 );
or \U$4055 ( \12851_13150 , \12787_13086 , \12788_13087 , \12789_13088 , \12790_13089 , \12791_13090 , \12792_13091 , \12793_13092 , \12794_13093 , \12795_13094 , \12796_13095 , \12797_13096 , \12798_13097 , \12799_13098 , \12800_13099 , \12801_13100 , \12802_13101 , \12803_13102 , \12804_13103 , \12805_13104 , \12806_13105 , \12807_13106 , \12808_13107 , \12809_13108 , \12810_13109 , \12811_13110 , \12812_13111 , \12813_13112 , \12814_13113 , \12815_13114 , \12816_13115 , \12817_13116 , \12818_13117 , \12819_13118 , \12820_13119 , \12821_13120 , \12822_13121 , \12823_13122 , \12824_13123 , \12825_13124 , \12826_13125 , \12827_13126 , \12828_13127 , \12829_13128 , \12830_13129 , \12831_13130 , \12832_13131 , \12833_13132 , \12834_13133 , \12835_13134 , \12836_13135 , \12837_13136 , \12838_13137 , \12839_13138 , \12840_13139 , \12841_13140 , \12842_13141 , \12843_13142 , \12844_13143 , \12845_13144 , \12846_13145 , \12847_13146 , \12848_13147 , \12849_13148 , \12850_13149 );
and \U$4056 ( \12852_13151 , RIfcb1860_7042, \8889_9188 );
and \U$4057 ( \12853_13152 , RIfca1b40_6862, \8891_9190 );
and \U$4058 ( \12854_13153 , RIfc5c018_6069, \8893_9192 );
and \U$4059 ( \12855_13154 , RIfe9ada0_8106, \8895_9194 );
and \U$4060 ( \12856_13155 , RIdf2b318_1868, \8897_9196 );
and \U$4061 ( \12857_13156 , RIdf29428_1846, \8899_9198 );
and \U$4062 ( \12858_13157 , RIdf27100_1821, \8901_9200 );
and \U$4063 ( \12859_13158 , RIfe9af08_8107, \8903_9202 );
and \U$4064 ( \12860_13159 , RIfc5e1d8_6093, \8905_9204 );
and \U$4065 ( \12861_13160 , RIfcdcda8_7535, \8907_9206 );
and \U$4066 ( \12862_13161 , RIfcac400_6982, \8909_9208 );
and \U$4067 ( \12863_13162 , RIfc691a0_6218, \8911_9210 );
and \U$4068 ( \12864_13163 , RIfcaad80_6966, \8913_9212 );
and \U$4069 ( \12865_13164 , RIdf20bc0_1749, \8915_9214 );
and \U$4070 ( \12866_13165 , RIfc61b80_6134, \8917_9216 );
and \U$4071 ( \12867_13166 , RIdf1a518_1676, \8919_9218 );
and \U$4072 ( \12868_13167 , RIdf184c0_1653, \8921_9220 );
and \U$4073 ( \12869_13168 , RIdf157c0_1621, \8923_9222 );
and \U$4074 ( \12870_13169 , RIdf12ac0_1589, \8925_9224 );
and \U$4075 ( \12871_13170 , RIdf0fdc0_1557, \8927_9226 );
and \U$4076 ( \12872_13171 , RIdf0d0c0_1525, \8929_9228 );
and \U$4077 ( \12873_13172 , RIdf0a3c0_1493, \8931_9230 );
and \U$4078 ( \12874_13173 , RIdf076c0_1461, \8933_9232 );
and \U$4079 ( \12875_13174 , RIdf049c0_1429, \8935_9234 );
and \U$4080 ( \12876_13175 , RIdefefc0_1365, \8937_9236 );
and \U$4081 ( \12877_13176 , RIdefc2c0_1333, \8939_9238 );
and \U$4082 ( \12878_13177 , RIdef95c0_1301, \8941_9240 );
and \U$4083 ( \12879_13178 , RIdef68c0_1269, \8943_9242 );
and \U$4084 ( \12880_13179 , RIdef3bc0_1237, \8945_9244 );
and \U$4085 ( \12881_13180 , RIdef0ec0_1205, \8947_9246 );
and \U$4086 ( \12882_13181 , RIdeee1c0_1173, \8949_9248 );
and \U$4087 ( \12883_13182 , RIdeeb4c0_1141, \8951_9250 );
and \U$4088 ( \12884_13183 , RIfc69b78_6225, \8953_9252 );
and \U$4089 ( \12885_13184 , RIfc6b900_6246, \8955_9254 );
and \U$4090 ( \12886_13185 , RIfc4d270_5900, \8957_9256 );
and \U$4091 ( \12887_13186 , RIfced770_7724, \8959_9258 );
and \U$4092 ( \12888_13187 , RIdee5ac0_1077, \8961_9260 );
and \U$4093 ( \12889_13188 , RIdee3d38_1056, \8963_9262 );
and \U$4094 ( \12890_13189 , RIdee1a10_1031, \8965_9264 );
and \U$4095 ( \12891_13190 , RIdedfb20_1009, \8967_9266 );
and \U$4096 ( \12892_13191 , RIfc7ff40_6478, \8969_9268 );
and \U$4097 ( \12893_13192 , RIfca4408_6891, \8971_9270 );
and \U$4098 ( \12894_13193 , RIfcb5640_7086, \8973_9272 );
and \U$4099 ( \12895_13194 , RIee21700_4839, \8975_9274 );
and \U$4100 ( \12896_13195 , RIdeda990_951, \8977_9276 );
and \U$4101 ( \12897_13196 , RIded8500_925, \8979_9278 );
and \U$4102 ( \12898_13197 , RIded61d8_900, \8981_9280 );
and \U$4103 ( \12899_13198 , RIded4018_876, \8983_9282 );
and \U$4104 ( \12900_13199 , RIded1cf0_851, \8985_9284 );
and \U$4105 ( \12901_13200 , RIdeceff0_819, \8987_9286 );
and \U$4106 ( \12902_13201 , RIdecc2f0_787, \8989_9288 );
and \U$4107 ( \12903_13202 , RIdec95f0_755, \8991_9290 );
and \U$4108 ( \12904_13203 , RIdeb5af0_531, \8993_9292 );
and \U$4109 ( \12905_13204 , RIde99a58_339, \8995_9294 );
and \U$4110 ( \12906_13205 , RIe16f6f8_2645, \8997_9296 );
and \U$4111 ( \12907_13206 , RIe15b4f0_2416, \8999_9298 );
and \U$4112 ( \12908_13207 , RIe144cf0_2160, \9001_9300 );
and \U$4113 ( \12909_13208 , RIdf396e8_2030, \9003_9302 );
and \U$4114 ( \12910_13209 , RIdf2dd48_1898, \9005_9304 );
and \U$4115 ( \12911_13210 , RIdf1e5c8_1722, \9007_9306 );
and \U$4116 ( \12912_13211 , RIdf01cc0_1397, \9009_9308 );
and \U$4117 ( \12913_13212 , RIdee87c0_1109, \9011_9310 );
and \U$4118 ( \12914_13213 , RIdedd528_982, \9013_9312 );
and \U$4119 ( \12915_13214 , RIde7f9a0_212, \9015_9314 );
or \U$4120 ( \12916_13215 , \12852_13151 , \12853_13152 , \12854_13153 , \12855_13154 , \12856_13155 , \12857_13156 , \12858_13157 , \12859_13158 , \12860_13159 , \12861_13160 , \12862_13161 , \12863_13162 , \12864_13163 , \12865_13164 , \12866_13165 , \12867_13166 , \12868_13167 , \12869_13168 , \12870_13169 , \12871_13170 , \12872_13171 , \12873_13172 , \12874_13173 , \12875_13174 , \12876_13175 , \12877_13176 , \12878_13177 , \12879_13178 , \12880_13179 , \12881_13180 , \12882_13181 , \12883_13182 , \12884_13183 , \12885_13184 , \12886_13185 , \12887_13186 , \12888_13187 , \12889_13188 , \12890_13189 , \12891_13190 , \12892_13191 , \12893_13192 , \12894_13193 , \12895_13194 , \12896_13195 , \12897_13196 , \12898_13197 , \12899_13198 , \12900_13199 , \12901_13200 , \12902_13201 , \12903_13202 , \12904_13203 , \12905_13204 , \12906_13205 , \12907_13206 , \12908_13207 , \12909_13208 , \12910_13209 , \12911_13210 , \12912_13211 , \12913_13212 , \12914_13213 , \12915_13214 );
or \U$4121 ( \12917_13216 , \12851_13150 , \12916_13215 );
_DC \g2f32/U$1 ( \12918 , \12917_13216 , \9024_9323 );
buf \U$4122 ( \12919_13218 , \12918 );
and \U$4123 ( \12920_13219 , RIe19eb88_3183, \9034_9333 );
and \U$4124 ( \12921_13220 , RIe19be88_3151, \9036_9335 );
and \U$4125 ( \12922_13221 , RIfe9a698_8101, \9038_9337 );
and \U$4126 ( \12923_13222 , RIe199188_3119, \9040_9339 );
and \U$4127 ( \12924_13223 , RIfe9a530_8100, \9042_9341 );
and \U$4128 ( \12925_13224 , RIe196488_3087, \9044_9343 );
and \U$4129 ( \12926_13225 , RIe193788_3055, \9046_9345 );
and \U$4130 ( \12927_13226 , RIe190a88_3023, \9048_9347 );
and \U$4131 ( \12928_13227 , RIe18b088_2959, \9050_9349 );
and \U$4132 ( \12929_13228 , RIe188388_2927, \9052_9351 );
and \U$4133 ( \12930_13229 , RIfe9a800_8102, \9054_9353 );
and \U$4134 ( \12931_13230 , RIe185688_2895, \9056_9355 );
and \U$4135 ( \12932_13231 , RIfc8d938_6633, \9058_9357 );
and \U$4136 ( \12933_13232 , RIe182988_2863, \9060_9359 );
and \U$4137 ( \12934_13233 , RIe17fc88_2831, \9062_9361 );
and \U$4138 ( \12935_13234 , RIe17cf88_2799, \9064_9363 );
and \U$4139 ( \12936_13235 , RIfe9a3c8_8099, \9066_9365 );
and \U$4140 ( \12937_13236 , RIf1415a8_5203, \9068_9367 );
and \U$4141 ( \12938_13237 , RIfe9a260_8098, \9070_9369 );
and \U$4142 ( \12939_13238 , RIfe9a0f8_8097, \9072_9371 );
and \U$4143 ( \12940_13239 , RIfcb9150_7128, \9074_9373 );
and \U$4144 ( \12941_13240 , RIf13f820_5182, \9076_9375 );
and \U$4145 ( \12942_13241 , RIfc9fc50_6840, \9078_9377 );
and \U$4146 ( \12943_13242 , RIfce5340_7630, \9080_9379 );
and \U$4147 ( \12944_13243 , RIfc5cb58_6077, \9082_9381 );
and \U$4148 ( \12945_13244 , RIfc576f8_6017, \9084_9383 );
and \U$4149 ( \12946_13245 , RIfc780b0_6388, \9086_9385 );
and \U$4150 ( \12947_13246 , RIe1749f0_2704, \9088_9387 );
and \U$4151 ( \12948_13247 , RIfc7adb0_6420, \9090_9389 );
and \U$4152 ( \12949_13248 , RIfc7c2c8_6435, \9092_9391 );
and \U$4153 ( \12950_13249 , RIfcb2d78_7057, \9094_9393 );
and \U$4154 ( \12951_13250 , RIfc7e758_6461, \9096_9395 );
and \U$4155 ( \12952_13251 , RIfe9aad0_8104, \9098_9397 );
and \U$4156 ( \12953_13252 , RIe224ee0_4710, \9100_9399 );
and \U$4157 ( \12954_13253 , RIf16c3e8_5691, \9102_9401 );
and \U$4158 ( \12955_13254 , RIe2221e0_4678, \9104_9403 );
and \U$4159 ( \12956_13255 , RIfcd3898_7429, \9106_9405 );
and \U$4160 ( \12957_13256 , RIe21f4e0_4646, \9108_9407 );
and \U$4161 ( \12958_13257 , RIe219ae0_4582, \9110_9409 );
and \U$4162 ( \12959_13258 , RIe216de0_4550, \9112_9411 );
and \U$4163 ( \12960_13259 , RIfc880a0_6570, \9114_9413 );
and \U$4164 ( \12961_13260 , RIe2140e0_4518, \9116_9415 );
and \U$4165 ( \12962_13261 , RIf169c88_5663, \9118_9417 );
and \U$4166 ( \12963_13262 , RIe2113e0_4486, \9120_9419 );
and \U$4167 ( \12964_13263 , RIf168338_5645, \9122_9421 );
and \U$4168 ( \12965_13264 , RIe20e6e0_4454, \9124_9423 );
and \U$4169 ( \12966_13265 , RIe20b9e0_4422, \9126_9425 );
and \U$4170 ( \12967_13266 , RIe208ce0_4390, \9128_9427 );
and \U$4171 ( \12968_13267 , RIfce4c38_7625, \9130_9429 );
and \U$4172 ( \12969_13268 , RIfc9c6e0_6802, \9132_9431 );
and \U$4173 ( \12970_13269 , RIe2035b0_4328, \9134_9433 );
and \U$4174 ( \12971_13270 , RIe201af8_4309, \9136_9435 );
and \U$4175 ( \12972_13271 , RIfc500d8_5933, \9138_9437 );
and \U$4176 ( \12973_13272 , RIfc85c10_6544, \9140_9439 );
and \U$4177 ( \12974_13273 , RIfce81a8_7663, \9142_9441 );
and \U$4178 ( \12975_13274 , RIfce9c60_7682, \9144_9443 );
and \U$4179 ( \12976_13275 , RIf160e80_5562, \9146_9445 );
and \U$4180 ( \12977_13276 , RIf15ef90_5540, \9148_9447 );
and \U$4181 ( \12978_13277 , RIfe9a968_8103, \9150_9449 );
and \U$4182 ( \12979_13278 , RIfe9ac38_8105, \9152_9451 );
and \U$4183 ( \12980_13279 , RIfca8d28_6943, \9154_9453 );
and \U$4184 ( \12981_13280 , RIf15be58_5505, \9156_9455 );
and \U$4185 ( \12982_13281 , RIfcedba8_7727, \9158_9457 );
and \U$4186 ( \12983_13282 , RIfc6a988_6235, \9160_9459 );
or \U$4187 ( \12984_13283 , \12920_13219 , \12921_13220 , \12922_13221 , \12923_13222 , \12924_13223 , \12925_13224 , \12926_13225 , \12927_13226 , \12928_13227 , \12929_13228 , \12930_13229 , \12931_13230 , \12932_13231 , \12933_13232 , \12934_13233 , \12935_13234 , \12936_13235 , \12937_13236 , \12938_13237 , \12939_13238 , \12940_13239 , \12941_13240 , \12942_13241 , \12943_13242 , \12944_13243 , \12945_13244 , \12946_13245 , \12947_13246 , \12948_13247 , \12949_13248 , \12950_13249 , \12951_13250 , \12952_13251 , \12953_13252 , \12954_13253 , \12955_13254 , \12956_13255 , \12957_13256 , \12958_13257 , \12959_13258 , \12960_13259 , \12961_13260 , \12962_13261 , \12963_13262 , \12964_13263 , \12965_13264 , \12966_13265 , \12967_13266 , \12968_13267 , \12969_13268 , \12970_13269 , \12971_13270 , \12972_13271 , \12973_13272 , \12974_13273 , \12975_13274 , \12976_13275 , \12977_13276 , \12978_13277 , \12979_13278 , \12980_13279 , \12981_13280 , \12982_13281 , \12983_13282 );
and \U$4188 ( \12985_13284 , RIfc71cd8_6317, \9163_9462 );
and \U$4189 ( \12986_13285 , RIfccb198_7333, \9165_9464 );
and \U$4190 ( \12987_13286 , RIfcaa3a8_6959, \9167_9466 );
and \U$4191 ( \12988_13287 , RIfec3b88_8347, \9169_9468 );
and \U$4192 ( \12989_13288 , RIfc4c730_5892, \9171_9470 );
and \U$4193 ( \12990_13289 , RIfc6d688_6267, \9173_9472 );
and \U$4194 ( \12991_13290 , RIfca8e90_6944, \9175_9474 );
and \U$4195 ( \12992_13291 , RIe1f6860_4182, \9177_9476 );
and \U$4196 ( \12993_13292 , RIfc64e20_6170, \9179_9478 );
and \U$4197 ( \12994_13293 , RIfcaee30_7012, \9181_9480 );
and \U$4198 ( \12995_13294 , RIfccee10_7376, \9183_9482 );
and \U$4199 ( \12996_13295 , RIe1f4538_4157, \9185_9484 );
and \U$4200 ( \12997_13296 , RIfc63ea8_6159, \9187_9486 );
and \U$4201 ( \12998_13297 , RIfcaecc8_7011, \9189_9488 );
and \U$4202 ( \12999_13298 , RIfcae458_7005, \9191_9490 );
and \U$4203 ( \13000_13299 , RIfeab1c8_8263, \9193_9492 );
and \U$4204 ( \13001_13300 , RIe1ecc48_4071, \9195_9494 );
and \U$4205 ( \13002_13301 , RIe1e9f48_4039, \9197_9496 );
and \U$4206 ( \13003_13302 , RIe1e7248_4007, \9199_9498 );
and \U$4207 ( \13004_13303 , RIe1e4548_3975, \9201_9500 );
and \U$4208 ( \13005_13304 , RIe1e1848_3943, \9203_9502 );
and \U$4209 ( \13006_13305 , RIe1deb48_3911, \9205_9504 );
and \U$4210 ( \13007_13306 , RIe1dbe48_3879, \9207_9506 );
and \U$4211 ( \13008_13307 , RIe1d9148_3847, \9209_9508 );
and \U$4212 ( \13009_13308 , RIe1d3748_3783, \9211_9510 );
and \U$4213 ( \13010_13309 , RIe1d0a48_3751, \9213_9512 );
and \U$4214 ( \13011_13310 , RIe1cdd48_3719, \9215_9514 );
and \U$4215 ( \13012_13311 , RIe1cb048_3687, \9217_9516 );
and \U$4216 ( \13013_13312 , RIe1c8348_3655, \9219_9518 );
and \U$4217 ( \13014_13313 , RIe1c5648_3623, \9221_9520 );
and \U$4218 ( \13015_13314 , RIe1c2948_3591, \9223_9522 );
and \U$4219 ( \13016_13315 , RIe1bfc48_3559, \9225_9524 );
and \U$4220 ( \13017_13316 , RIfcc70e8_7287, \9227_9526 );
and \U$4221 ( \13018_13317 , RIfca7ae0_6930, \9229_9528 );
and \U$4222 ( \13019_13318 , RIe1ba518_3497, \9231_9530 );
and \U$4223 ( \13020_13319 , RIe1b8358_3473, \9233_9532 );
and \U$4224 ( \13021_13320 , RIfc598b8_6041, \9235_9534 );
and \U$4225 ( \13022_13321 , RIfcc2228_7231, \9237_9536 );
and \U$4226 ( \13023_13322 , RIe1b6198_3449, \9239_9538 );
and \U$4227 ( \13024_13323 , RIe1b4848_3431, \9241_9540 );
and \U$4228 ( \13025_13324 , RIfc82f10_6512, \9243_9542 );
and \U$4229 ( \13026_13325 , RIfc55970_5996, \9245_9544 );
and \U$4230 ( \13027_13326 , RIe1b3498_3417, \9247_9546 );
and \U$4231 ( \13028_13327 , RIe1b1cb0_3400, \9249_9548 );
and \U$4232 ( \13029_13328 , RIfcb7698_7109, \9251_9550 );
and \U$4233 ( \13030_13329 , RIfc4b4e8_5879, \9253_9552 );
and \U$4234 ( \13031_13330 , RIe1ad390_3348, \9255_9554 );
and \U$4235 ( \13032_13331 , RIe1abba8_3331, \9257_9556 );
and \U$4236 ( \13033_13332 , RIe1a9f88_3311, \9259_9558 );
and \U$4237 ( \13034_13333 , RIe1a7288_3279, \9261_9560 );
and \U$4238 ( \13035_13334 , RIe1a4588_3247, \9263_9562 );
and \U$4239 ( \13036_13335 , RIe1a1888_3215, \9265_9564 );
and \U$4240 ( \13037_13336 , RIe18dd88_2991, \9267_9566 );
and \U$4241 ( \13038_13337 , RIe17a288_2767, \9269_9568 );
and \U$4242 ( \13039_13338 , RIe227be0_4742, \9271_9570 );
and \U$4243 ( \13040_13339 , RIe21c7e0_4614, \9273_9572 );
and \U$4244 ( \13041_13340 , RIe205fe0_4358, \9275_9574 );
and \U$4245 ( \13042_13341 , RIe200040_4290, \9277_9576 );
and \U$4246 ( \13043_13342 , RIe1f93f8_4213, \9279_9578 );
and \U$4247 ( \13044_13343 , RIe1f1f40_4130, \9281_9580 );
and \U$4248 ( \13045_13344 , RIe1d6448_3815, \9283_9582 );
and \U$4249 ( \13046_13345 , RIe1bcf48_3527, \9285_9584 );
and \U$4250 ( \13047_13346 , RIe1afdc0_3378, \9287_9586 );
and \U$4251 ( \13048_13347 , RIe1723f8_2677, \9289_9588 );
or \U$4252 ( \13049_13348 , \12985_13284 , \12986_13285 , \12987_13286 , \12988_13287 , \12989_13288 , \12990_13289 , \12991_13290 , \12992_13291 , \12993_13292 , \12994_13293 , \12995_13294 , \12996_13295 , \12997_13296 , \12998_13297 , \12999_13298 , \13000_13299 , \13001_13300 , \13002_13301 , \13003_13302 , \13004_13303 , \13005_13304 , \13006_13305 , \13007_13306 , \13008_13307 , \13009_13308 , \13010_13309 , \13011_13310 , \13012_13311 , \13013_13312 , \13014_13313 , \13015_13314 , \13016_13315 , \13017_13316 , \13018_13317 , \13019_13318 , \13020_13319 , \13021_13320 , \13022_13321 , \13023_13322 , \13024_13323 , \13025_13324 , \13026_13325 , \13027_13326 , \13028_13327 , \13029_13328 , \13030_13329 , \13031_13330 , \13032_13331 , \13033_13332 , \13034_13333 , \13035_13334 , \13036_13335 , \13037_13336 , \13038_13337 , \13039_13338 , \13040_13339 , \13041_13340 , \13042_13341 , \13043_13342 , \13044_13343 , \13045_13344 , \13046_13345 , \13047_13346 , \13048_13347 );
or \U$4253 ( \13050_13349 , \12984_13283 , \13049_13348 );
_DC \g405f/U$1 ( \13051 , \13050_13349 , \9298_9597 );
buf \U$4254 ( \13052_13351 , \13051 );
and \U$4255 ( \13053_13352 , \12919_13218 , \13052_13351 );
and \U$4256 ( \13054_13353 , \11439_11738 , \11572_11871 );
and \U$4257 ( \13055_13354 , \11572_11871 , \11847_12146 );
and \U$4258 ( \13056_13355 , \11439_11738 , \11847_12146 );
or \U$4259 ( \13057_13356 , \13054_13353 , \13055_13354 , \13056_13355 );
and \U$4260 ( \13058_13357 , \13052_13351 , \13057_13356 );
and \U$4261 ( \13059_13358 , \12919_13218 , \13057_13356 );
or \U$4262 ( \13060_13359 , \13053_13352 , \13058_13357 , \13059_13358 );
xor \U$4263 ( \13061_13360 , \12786_13085 , \13060_13359 );
buf g4442_GF_PartitionCandidate( \13062_13361_nG4442 , \13061_13360 );
xor \U$4264 ( \13063_13362 , \12919_13218 , \13052_13351 );
xor \U$4265 ( \13064_13363 , \13063_13362 , \13057_13356 );
buf g4445_GF_PartitionCandidate( \13065_13364_nG4445 , \13064_13363 );
nand \U$4266 ( \13066_13365 , \13065_13364_nG4445 , \11849_12148_nG4448 );
and \U$4267 ( \13067_13366 , \13062_13361_nG4442 , \13066_13365 );
xor \U$4268 ( \13068_13367 , \13065_13364_nG4445 , \11849_12148_nG4448 );
and \U$4273 ( \13069_13371 , \13068_13367 , \10392_10694_nG9c0e );
or \U$4274 ( \13070_13372 , 1'b0 , \13069_13371 );
xor \U$4275 ( \13071_13373 , \13067_13366 , \13070_13372 );
xor \U$4276 ( \13072_13374 , \13067_13366 , \13071_13373 );
buf \U$4277 ( \13073_13375 , \13072_13374 );
buf \U$4278 ( \13074_13376 , \13073_13375 );
and \U$4279 ( \13075_13377 , \12519_12818 , \13074_13376 );
and \U$4280 ( \13076_13378 , \12509_12808 , \12514_12813 );
and \U$4281 ( \13077_13379 , \12509_12808 , \12517_12816 );
and \U$4282 ( \13078_13380 , \12514_12813 , \12517_12816 );
or \U$4283 ( \13079_13381 , \13076_13378 , \13077_13379 , \13078_13380 );
buf \U$4284 ( \13080_13382 , \13079_13381 );
and \U$4285 ( \13081_13383 , \12191_12490 , \12197_12496 );
and \U$4286 ( \13082_13384 , \12191_12490 , \12507_12806 );
and \U$4287 ( \13083_13385 , \12197_12496 , \12507_12806 );
or \U$4288 ( \13084_13386 , \13081_13383 , \13082_13384 , \13083_13385 );
buf \U$4289 ( \13085_13387 , \13084_13386 );
xor \U$4290 ( \13086_13388 , \13080_13382 , \13085_13387 );
and \U$4291 ( \13087_13389 , \12180_12482 , \12189_12488 );
buf \U$4292 ( \13088_13390 , \13087_13389 );
and \U$4293 ( \13089_13391 , \12183_12157 , \10693_10995_nG9c0b );
and \U$4294 ( \13090_13392 , \11855_12154 , \10981_11283_nG9c08 );
or \U$4295 ( \13091_13393 , \13089_13391 , \13090_13392 );
xor \U$4296 ( \13092_13394 , \11854_12153 , \13091_13393 );
buf \U$4297 ( \13093_13395 , \13092_13394 );
buf \U$4299 ( \13094_13396 , \13093_13395 );
xor \U$4300 ( \13095_13397 , \13088_13390 , \13094_13396 );
buf \U$4301 ( \13096_13398 , \13095_13397 );
and \U$4302 ( \13097_13399 , \10996_10421 , \11299_11598_nG9c05 );
and \U$4303 ( \13098_13400 , \10119_10418 , \12168_12470_nG9c02 );
or \U$4304 ( \13099_13401 , \13097_13399 , \13098_13400 );
xor \U$4305 ( \13100_13402 , \10118_10417 , \13099_13401 );
buf \U$4306 ( \13101_13403 , \13100_13402 );
buf \U$4308 ( \13102_13404 , \13101_13403 );
xor \U$4309 ( \13103_13405 , \13096_13398 , \13102_13404 );
and \U$4310 ( \13104_13406 , \10411_10707 , \12502_12801_nG9bff );
and \U$4311 ( \13105_13407 , \12473_12772 , \12482_12781 );
and \U$4312 ( \13106_13408 , \10686_10988 , \12491_12790 );
and \U$4313 ( \13107_13409 , \10968_11270 , \12159_12461 );
nor \U$4314 ( \13108_13410 , \13106_13408 , \13107_13409 );
xnor \U$4315 ( \13109_13411 , \13108_13410 , \12481_12780 );
xor \U$4316 ( \13110_13412 , \13105_13407 , \13109_13411 );
and \U$4317 ( \13111_13413 , \12470_12769 , \10681_10983 );
and \U$4318 ( \13112_13414 , RIdec68f0_723, \9034_9333 );
and \U$4319 ( \13113_13415 , RIdec3bf0_691, \9036_9335 );
and \U$4320 ( \13114_13416 , RIee208f0_4829, \9038_9337 );
and \U$4321 ( \13115_13417 , RIdec0ef0_659, \9040_9339 );
and \U$4322 ( \13116_13418 , RIfc7ce08_6443, \9042_9341 );
and \U$4323 ( \13117_13419 , RIdebe1f0_627, \9044_9343 );
and \U$4324 ( \13118_13420 , RIdebb4f0_595, \9046_9345 );
and \U$4325 ( \13119_13421 , RIdeb87f0_563, \9048_9347 );
and \U$4326 ( \13120_13422 , RIfc9b8d0_6792, \9050_9349 );
and \U$4327 ( \13121_13423 , RIdeb2df0_499, \9052_9351 );
and \U$4328 ( \13122_13424 , RIfcc6710_7280, \9054_9353 );
and \U$4329 ( \13123_13425 , RIdeb00f0_467, \9056_9355 );
and \U$4330 ( \13124_13426 , RIfc5ff60_6114, \9058_9357 );
and \U$4331 ( \13125_13427 , RIdead3f0_435, \9060_9359 );
and \U$4332 ( \13126_13428 , RIdea6c58_403, \9062_9361 );
and \U$4333 ( \13127_13429 , RIdea0358_371, \9064_9363 );
and \U$4334 ( \13128_13430 , RIfce5070_7628, \9066_9365 );
and \U$4335 ( \13129_13431 , RIee1c6d8_4782, \9068_9367 );
and \U$4336 ( \13130_13432 , RIfce70c8_7651, \9070_9369 );
and \U$4337 ( \13131_13433 , RIee1b058_4766, \9072_9371 );
and \U$4338 ( \13132_13434 , RIde934a0_308, \9074_9373 );
and \U$4339 ( \13133_13435 , RIfe9b1d8_8109, \9076_9375 );
and \U$4340 ( \13134_13436 , RIde8b7f0_270, \9078_9377 );
and \U$4341 ( \13135_13437 , RIfe9b340_8110, \9080_9379 );
and \U$4342 ( \13136_13438 , RIfc6b798_6245, \9082_9381 );
and \U$4343 ( \13137_13439 , RIfcb2238_7049, \9084_9383 );
and \U$4344 ( \13138_13440 , RIfcd3a00_7430, \9086_9385 );
and \U$4345 ( \13139_13441 , RIfcdb020_7514, \9088_9387 );
and \U$4346 ( \13140_13442 , RIfc511b8_5945, \9090_9389 );
and \U$4347 ( \13141_13443 , RIe16c9f8_2613, \9092_9391 );
and \U$4348 ( \13142_13444 , RIfcb27d8_7053, \9094_9393 );
and \U$4349 ( \13143_13445 , RIe168ee8_2571, \9096_9395 );
and \U$4350 ( \13144_13446 , RIe1668f0_2544, \9098_9397 );
and \U$4351 ( \13145_13447 , RIe163bf0_2512, \9100_9399 );
and \U$4352 ( \13146_13448 , RIee381d0_5097, \9102_9401 );
and \U$4353 ( \13147_13449 , RIe160ef0_2480, \9104_9403 );
and \U$4354 ( \13148_13450 , RIfcdfaa8_7567, \9106_9405 );
and \U$4355 ( \13149_13451 , RIe15e1f0_2448, \9108_9407 );
and \U$4356 ( \13150_13452 , RIe1587f0_2384, \9110_9409 );
and \U$4357 ( \13151_13453 , RIe155af0_2352, \9112_9411 );
and \U$4358 ( \13152_13454 , RIfc3f968_5749, \9114_9413 );
and \U$4359 ( \13153_13455 , RIe152df0_2320, \9116_9415 );
and \U$4360 ( \13154_13456 , RIfcd5080_7446, \9118_9417 );
and \U$4361 ( \13155_13457 , RIe1500f0_2288, \9120_9419 );
and \U$4362 ( \13156_13458 , RIfc84b30_6532, \9122_9421 );
and \U$4363 ( \13157_13459 , RIe14d3f0_2256, \9124_9423 );
and \U$4364 ( \13158_13460 , RIe14a6f0_2224, \9126_9425 );
and \U$4365 ( \13159_13461 , RIe1479f0_2192, \9128_9427 );
and \U$4366 ( \13160_13462 , RIfcea098_7685, \9130_9429 );
and \U$4367 ( \13161_13463 , RIfc92f00_6694, \9132_9431 );
and \U$4368 ( \13162_13464 , RIfc54890_5984, \9134_9433 );
and \U$4369 ( \13163_13465 , RIfcdcc40_7534, \9136_9435 );
and \U$4370 ( \13164_13466 , RIe142158_2129, \9138_9437 );
and \U$4371 ( \13165_13467 , RIe13fe30_2104, \9140_9439 );
and \U$4372 ( \13166_13468 , RIdf3dd38_2080, \9142_9441 );
and \U$4373 ( \13167_13469 , RIdf3b8a8_2054, \9144_9443 );
and \U$4374 ( \13168_13470 , RIfc57590_6016, \9146_9445 );
and \U$4375 ( \13169_13471 , RIee30340_5007, \9148_9447 );
and \U$4376 ( \13170_13472 , RIfcd0490_7392, \9150_9449 );
and \U$4377 ( \13171_13473 , RIee2e180_4983, \9152_9451 );
and \U$4378 ( \13172_13474 , RIdf36b50_1999, \9154_9453 );
and \U$4379 ( \13173_13475 , RIdf34558_1972, \9156_9455 );
and \U$4380 ( \13174_13476 , RIdf32398_1948, \9158_9457 );
and \U$4381 ( \13175_13477 , RIfe9b070_8108, \9160_9459 );
or \U$4382 ( \13176_13478 , \13112_13414 , \13113_13415 , \13114_13416 , \13115_13417 , \13116_13418 , \13117_13419 , \13118_13420 , \13119_13421 , \13120_13422 , \13121_13423 , \13122_13424 , \13123_13425 , \13124_13426 , \13125_13427 , \13126_13428 , \13127_13429 , \13128_13430 , \13129_13431 , \13130_13432 , \13131_13433 , \13132_13434 , \13133_13435 , \13134_13436 , \13135_13437 , \13136_13438 , \13137_13439 , \13138_13440 , \13139_13441 , \13140_13442 , \13141_13443 , \13142_13444 , \13143_13445 , \13144_13446 , \13145_13447 , \13146_13448 , \13147_13449 , \13148_13450 , \13149_13451 , \13150_13452 , \13151_13453 , \13152_13454 , \13153_13455 , \13154_13456 , \13155_13457 , \13156_13458 , \13157_13459 , \13158_13460 , \13159_13461 , \13160_13462 , \13161_13463 , \13162_13464 , \13163_13465 , \13164_13466 , \13165_13467 , \13166_13468 , \13167_13469 , \13168_13470 , \13169_13471 , \13170_13472 , \13171_13473 , \13172_13474 , \13173_13475 , \13174_13476 , \13175_13477 );
and \U$4383 ( \13177_13479 , RIfcb1860_7042, \9163_9462 );
and \U$4384 ( \13178_13480 , RIfca1b40_6862, \9165_9464 );
and \U$4385 ( \13179_13481 , RIfc5c018_6069, \9167_9466 );
and \U$4386 ( \13180_13482 , RIfe9ada0_8106, \9169_9468 );
and \U$4387 ( \13181_13483 , RIdf2b318_1868, \9171_9470 );
and \U$4388 ( \13182_13484 , RIdf29428_1846, \9173_9472 );
and \U$4389 ( \13183_13485 , RIdf27100_1821, \9175_9474 );
and \U$4390 ( \13184_13486 , RIfe9af08_8107, \9177_9476 );
and \U$4391 ( \13185_13487 , RIfc5e1d8_6093, \9179_9478 );
and \U$4392 ( \13186_13488 , RIfcdcda8_7535, \9181_9480 );
and \U$4393 ( \13187_13489 , RIfcac400_6982, \9183_9482 );
and \U$4394 ( \13188_13490 , RIfc691a0_6218, \9185_9484 );
and \U$4395 ( \13189_13491 , RIfcaad80_6966, \9187_9486 );
and \U$4396 ( \13190_13492 , RIdf20bc0_1749, \9189_9488 );
and \U$4397 ( \13191_13493 , RIfc61b80_6134, \9191_9490 );
and \U$4398 ( \13192_13494 , RIdf1a518_1676, \9193_9492 );
and \U$4399 ( \13193_13495 , RIdf184c0_1653, \9195_9494 );
and \U$4400 ( \13194_13496 , RIdf157c0_1621, \9197_9496 );
and \U$4401 ( \13195_13497 , RIdf12ac0_1589, \9199_9498 );
and \U$4402 ( \13196_13498 , RIdf0fdc0_1557, \9201_9500 );
and \U$4403 ( \13197_13499 , RIdf0d0c0_1525, \9203_9502 );
and \U$4404 ( \13198_13500 , RIdf0a3c0_1493, \9205_9504 );
and \U$4405 ( \13199_13501 , RIdf076c0_1461, \9207_9506 );
and \U$4406 ( \13200_13502 , RIdf049c0_1429, \9209_9508 );
and \U$4407 ( \13201_13503 , RIdefefc0_1365, \9211_9510 );
and \U$4408 ( \13202_13504 , RIdefc2c0_1333, \9213_9512 );
and \U$4409 ( \13203_13505 , RIdef95c0_1301, \9215_9514 );
and \U$4410 ( \13204_13506 , RIdef68c0_1269, \9217_9516 );
and \U$4411 ( \13205_13507 , RIdef3bc0_1237, \9219_9518 );
and \U$4412 ( \13206_13508 , RIdef0ec0_1205, \9221_9520 );
and \U$4413 ( \13207_13509 , RIdeee1c0_1173, \9223_9522 );
and \U$4414 ( \13208_13510 , RIdeeb4c0_1141, \9225_9524 );
and \U$4415 ( \13209_13511 , RIfc69b78_6225, \9227_9526 );
and \U$4416 ( \13210_13512 , RIfc6b900_6246, \9229_9528 );
and \U$4417 ( \13211_13513 , RIfc4d270_5900, \9231_9530 );
and \U$4418 ( \13212_13514 , RIfced770_7724, \9233_9532 );
and \U$4419 ( \13213_13515 , RIdee5ac0_1077, \9235_9534 );
and \U$4420 ( \13214_13516 , RIdee3d38_1056, \9237_9536 );
and \U$4421 ( \13215_13517 , RIdee1a10_1031, \9239_9538 );
and \U$4422 ( \13216_13518 , RIdedfb20_1009, \9241_9540 );
and \U$4423 ( \13217_13519 , RIfc7ff40_6478, \9243_9542 );
and \U$4424 ( \13218_13520 , RIfca4408_6891, \9245_9544 );
and \U$4425 ( \13219_13521 , RIfcb5640_7086, \9247_9546 );
and \U$4426 ( \13220_13522 , RIee21700_4839, \9249_9548 );
and \U$4427 ( \13221_13523 , RIdeda990_951, \9251_9550 );
and \U$4428 ( \13222_13524 , RIded8500_925, \9253_9552 );
and \U$4429 ( \13223_13525 , RIded61d8_900, \9255_9554 );
and \U$4430 ( \13224_13526 , RIded4018_876, \9257_9556 );
and \U$4431 ( \13225_13527 , RIded1cf0_851, \9259_9558 );
and \U$4432 ( \13226_13528 , RIdeceff0_819, \9261_9560 );
and \U$4433 ( \13227_13529 , RIdecc2f0_787, \9263_9562 );
and \U$4434 ( \13228_13530 , RIdec95f0_755, \9265_9564 );
and \U$4435 ( \13229_13531 , RIdeb5af0_531, \9267_9566 );
and \U$4436 ( \13230_13532 , RIde99a58_339, \9269_9568 );
and \U$4437 ( \13231_13533 , RIe16f6f8_2645, \9271_9570 );
and \U$4438 ( \13232_13534 , RIe15b4f0_2416, \9273_9572 );
and \U$4439 ( \13233_13535 , RIe144cf0_2160, \9275_9574 );
and \U$4440 ( \13234_13536 , RIdf396e8_2030, \9277_9576 );
and \U$4441 ( \13235_13537 , RIdf2dd48_1898, \9279_9578 );
and \U$4442 ( \13236_13538 , RIdf1e5c8_1722, \9281_9580 );
and \U$4443 ( \13237_13539 , RIdf01cc0_1397, \9283_9582 );
and \U$4444 ( \13238_13540 , RIdee87c0_1109, \9285_9584 );
and \U$4445 ( \13239_13541 , RIdedd528_982, \9287_9586 );
and \U$4446 ( \13240_13542 , RIde7f9a0_212, \9289_9588 );
or \U$4447 ( \13241_13543 , \13177_13479 , \13178_13480 , \13179_13481 , \13180_13482 , \13181_13483 , \13182_13484 , \13183_13485 , \13184_13486 , \13185_13487 , \13186_13488 , \13187_13489 , \13188_13490 , \13189_13491 , \13190_13492 , \13191_13493 , \13192_13494 , \13193_13495 , \13194_13496 , \13195_13497 , \13196_13498 , \13197_13499 , \13198_13500 , \13199_13501 , \13200_13502 , \13201_13503 , \13202_13504 , \13203_13505 , \13204_13506 , \13205_13507 , \13206_13508 , \13207_13509 , \13208_13510 , \13209_13511 , \13210_13512 , \13211_13513 , \13212_13514 , \13213_13515 , \13214_13516 , \13215_13517 , \13216_13518 , \13217_13519 , \13218_13520 , \13219_13521 , \13220_13522 , \13221_13523 , \13222_13524 , \13223_13525 , \13224_13526 , \13225_13527 , \13226_13528 , \13227_13529 , \13228_13530 , \13229_13531 , \13230_13532 , \13231_13533 , \13232_13534 , \13233_13535 , \13234_13536 , \13235_13537 , \13236_13538 , \13237_13539 , \13238_13540 , \13239_13541 , \13240_13542 );
or \U$4448 ( \13242_13544 , \13176_13478 , \13241_13543 );
_DC \g6589/U$1 ( \13243 , \13242_13544 , \9298_9597 );
and \U$4449 ( \13244_13546 , RIe19eb88_3183, \8760_9059 );
and \U$4450 ( \13245_13547 , RIe19be88_3151, \8762_9061 );
and \U$4451 ( \13246_13548 , RIfe9a698_8101, \8764_9063 );
and \U$4452 ( \13247_13549 , RIe199188_3119, \8766_9065 );
and \U$4453 ( \13248_13550 , RIfe9a530_8100, \8768_9067 );
and \U$4454 ( \13249_13551 , RIe196488_3087, \8770_9069 );
and \U$4455 ( \13250_13552 , RIe193788_3055, \8772_9071 );
and \U$4456 ( \13251_13553 , RIe190a88_3023, \8774_9073 );
and \U$4457 ( \13252_13554 , RIe18b088_2959, \8776_9075 );
and \U$4458 ( \13253_13555 , RIe188388_2927, \8778_9077 );
and \U$4459 ( \13254_13556 , RIfe9a800_8102, \8780_9079 );
and \U$4460 ( \13255_13557 , RIe185688_2895, \8782_9081 );
and \U$4461 ( \13256_13558 , RIfc8d938_6633, \8784_9083 );
and \U$4462 ( \13257_13559 , RIe182988_2863, \8786_9085 );
and \U$4463 ( \13258_13560 , RIe17fc88_2831, \8788_9087 );
and \U$4464 ( \13259_13561 , RIe17cf88_2799, \8790_9089 );
and \U$4465 ( \13260_13562 , RIfe9a3c8_8099, \8792_9091 );
and \U$4466 ( \13261_13563 , RIf1415a8_5203, \8794_9093 );
and \U$4467 ( \13262_13564 , RIfe9a260_8098, \8796_9095 );
and \U$4468 ( \13263_13565 , RIfe9a0f8_8097, \8798_9097 );
and \U$4469 ( \13264_13566 , RIfcb9150_7128, \8800_9099 );
and \U$4470 ( \13265_13567 , RIf13f820_5182, \8802_9101 );
and \U$4471 ( \13266_13568 , RIfc9fc50_6840, \8804_9103 );
and \U$4472 ( \13267_13569 , RIfce5340_7630, \8806_9105 );
and \U$4473 ( \13268_13570 , RIfc5cb58_6077, \8808_9107 );
and \U$4474 ( \13269_13571 , RIfc576f8_6017, \8810_9109 );
and \U$4475 ( \13270_13572 , RIfc780b0_6388, \8812_9111 );
and \U$4476 ( \13271_13573 , RIe1749f0_2704, \8814_9113 );
and \U$4477 ( \13272_13574 , RIfc7adb0_6420, \8816_9115 );
and \U$4478 ( \13273_13575 , RIfc7c2c8_6435, \8818_9117 );
and \U$4479 ( \13274_13576 , RIfcb2d78_7057, \8820_9119 );
and \U$4480 ( \13275_13577 , RIfc7e758_6461, \8822_9121 );
and \U$4481 ( \13276_13578 , RIfe9aad0_8104, \8824_9123 );
and \U$4482 ( \13277_13579 , RIe224ee0_4710, \8826_9125 );
and \U$4483 ( \13278_13580 , RIf16c3e8_5691, \8828_9127 );
and \U$4484 ( \13279_13581 , RIe2221e0_4678, \8830_9129 );
and \U$4485 ( \13280_13582 , RIfcd3898_7429, \8832_9131 );
and \U$4486 ( \13281_13583 , RIe21f4e0_4646, \8834_9133 );
and \U$4487 ( \13282_13584 , RIe219ae0_4582, \8836_9135 );
and \U$4488 ( \13283_13585 , RIe216de0_4550, \8838_9137 );
and \U$4489 ( \13284_13586 , RIfc880a0_6570, \8840_9139 );
and \U$4490 ( \13285_13587 , RIe2140e0_4518, \8842_9141 );
and \U$4491 ( \13286_13588 , RIf169c88_5663, \8844_9143 );
and \U$4492 ( \13287_13589 , RIe2113e0_4486, \8846_9145 );
and \U$4493 ( \13288_13590 , RIf168338_5645, \8848_9147 );
and \U$4494 ( \13289_13591 , RIe20e6e0_4454, \8850_9149 );
and \U$4495 ( \13290_13592 , RIe20b9e0_4422, \8852_9151 );
and \U$4496 ( \13291_13593 , RIe208ce0_4390, \8854_9153 );
and \U$4497 ( \13292_13594 , RIfce4c38_7625, \8856_9155 );
and \U$4498 ( \13293_13595 , RIfc9c6e0_6802, \8858_9157 );
and \U$4499 ( \13294_13596 , RIe2035b0_4328, \8860_9159 );
and \U$4500 ( \13295_13597 , RIe201af8_4309, \8862_9161 );
and \U$4501 ( \13296_13598 , RIfc500d8_5933, \8864_9163 );
and \U$4502 ( \13297_13599 , RIfc85c10_6544, \8866_9165 );
and \U$4503 ( \13298_13600 , RIfce81a8_7663, \8868_9167 );
and \U$4504 ( \13299_13601 , RIfce9c60_7682, \8870_9169 );
and \U$4505 ( \13300_13602 , RIf160e80_5562, \8872_9171 );
and \U$4506 ( \13301_13603 , RIf15ef90_5540, \8874_9173 );
and \U$4507 ( \13302_13604 , RIfe9a968_8103, \8876_9175 );
and \U$4508 ( \13303_13605 , RIfe9ac38_8105, \8878_9177 );
and \U$4509 ( \13304_13606 , RIfca8d28_6943, \8880_9179 );
and \U$4510 ( \13305_13607 , RIf15be58_5505, \8882_9181 );
and \U$4511 ( \13306_13608 , RIfcedba8_7727, \8884_9183 );
and \U$4512 ( \13307_13609 , RIfc6a988_6235, \8886_9185 );
or \U$4513 ( \13308_13610 , \13244_13546 , \13245_13547 , \13246_13548 , \13247_13549 , \13248_13550 , \13249_13551 , \13250_13552 , \13251_13553 , \13252_13554 , \13253_13555 , \13254_13556 , \13255_13557 , \13256_13558 , \13257_13559 , \13258_13560 , \13259_13561 , \13260_13562 , \13261_13563 , \13262_13564 , \13263_13565 , \13264_13566 , \13265_13567 , \13266_13568 , \13267_13569 , \13268_13570 , \13269_13571 , \13270_13572 , \13271_13573 , \13272_13574 , \13273_13575 , \13274_13576 , \13275_13577 , \13276_13578 , \13277_13579 , \13278_13580 , \13279_13581 , \13280_13582 , \13281_13583 , \13282_13584 , \13283_13585 , \13284_13586 , \13285_13587 , \13286_13588 , \13287_13589 , \13288_13590 , \13289_13591 , \13290_13592 , \13291_13593 , \13292_13594 , \13293_13595 , \13294_13596 , \13295_13597 , \13296_13598 , \13297_13599 , \13298_13600 , \13299_13601 , \13300_13602 , \13301_13603 , \13302_13604 , \13303_13605 , \13304_13606 , \13305_13607 , \13306_13608 , \13307_13609 );
and \U$4514 ( \13309_13611 , RIfc71cd8_6317, \8889_9188 );
and \U$4515 ( \13310_13612 , RIfccb198_7333, \8891_9190 );
and \U$4516 ( \13311_13613 , RIfcaa3a8_6959, \8893_9192 );
and \U$4517 ( \13312_13614 , RIfec3b88_8347, \8895_9194 );
and \U$4518 ( \13313_13615 , RIfc4c730_5892, \8897_9196 );
and \U$4519 ( \13314_13616 , RIfc6d688_6267, \8899_9198 );
and \U$4520 ( \13315_13617 , RIfca8e90_6944, \8901_9200 );
and \U$4521 ( \13316_13618 , RIe1f6860_4182, \8903_9202 );
and \U$4522 ( \13317_13619 , RIfc64e20_6170, \8905_9204 );
and \U$4523 ( \13318_13620 , RIfcaee30_7012, \8907_9206 );
and \U$4524 ( \13319_13621 , RIfccee10_7376, \8909_9208 );
and \U$4525 ( \13320_13622 , RIe1f4538_4157, \8911_9210 );
and \U$4526 ( \13321_13623 , RIfc63ea8_6159, \8913_9212 );
and \U$4527 ( \13322_13624 , RIfcaecc8_7011, \8915_9214 );
and \U$4528 ( \13323_13625 , RIfcae458_7005, \8917_9216 );
and \U$4529 ( \13324_13626 , RIfeab1c8_8263, \8919_9218 );
and \U$4530 ( \13325_13627 , RIe1ecc48_4071, \8921_9220 );
and \U$4531 ( \13326_13628 , RIe1e9f48_4039, \8923_9222 );
and \U$4532 ( \13327_13629 , RIe1e7248_4007, \8925_9224 );
and \U$4533 ( \13328_13630 , RIe1e4548_3975, \8927_9226 );
and \U$4534 ( \13329_13631 , RIe1e1848_3943, \8929_9228 );
and \U$4535 ( \13330_13632 , RIe1deb48_3911, \8931_9230 );
and \U$4536 ( \13331_13633 , RIe1dbe48_3879, \8933_9232 );
and \U$4537 ( \13332_13634 , RIe1d9148_3847, \8935_9234 );
and \U$4538 ( \13333_13635 , RIe1d3748_3783, \8937_9236 );
and \U$4539 ( \13334_13636 , RIe1d0a48_3751, \8939_9238 );
and \U$4540 ( \13335_13637 , RIe1cdd48_3719, \8941_9240 );
and \U$4541 ( \13336_13638 , RIe1cb048_3687, \8943_9242 );
and \U$4542 ( \13337_13639 , RIe1c8348_3655, \8945_9244 );
and \U$4543 ( \13338_13640 , RIe1c5648_3623, \8947_9246 );
and \U$4544 ( \13339_13641 , RIe1c2948_3591, \8949_9248 );
and \U$4545 ( \13340_13642 , RIe1bfc48_3559, \8951_9250 );
and \U$4546 ( \13341_13643 , RIfcc70e8_7287, \8953_9252 );
and \U$4547 ( \13342_13644 , RIfca7ae0_6930, \8955_9254 );
and \U$4548 ( \13343_13645 , RIe1ba518_3497, \8957_9256 );
and \U$4549 ( \13344_13646 , RIe1b8358_3473, \8959_9258 );
and \U$4550 ( \13345_13647 , RIfc598b8_6041, \8961_9260 );
and \U$4551 ( \13346_13648 , RIfcc2228_7231, \8963_9262 );
and \U$4552 ( \13347_13649 , RIe1b6198_3449, \8965_9264 );
and \U$4553 ( \13348_13650 , RIe1b4848_3431, \8967_9266 );
and \U$4554 ( \13349_13651 , RIfc82f10_6512, \8969_9268 );
and \U$4555 ( \13350_13652 , RIfc55970_5996, \8971_9270 );
and \U$4556 ( \13351_13653 , RIe1b3498_3417, \8973_9272 );
and \U$4557 ( \13352_13654 , RIe1b1cb0_3400, \8975_9274 );
and \U$4558 ( \13353_13655 , RIfcb7698_7109, \8977_9276 );
and \U$4559 ( \13354_13656 , RIfc4b4e8_5879, \8979_9278 );
and \U$4560 ( \13355_13657 , RIe1ad390_3348, \8981_9280 );
and \U$4561 ( \13356_13658 , RIe1abba8_3331, \8983_9282 );
and \U$4562 ( \13357_13659 , RIe1a9f88_3311, \8985_9284 );
and \U$4563 ( \13358_13660 , RIe1a7288_3279, \8987_9286 );
and \U$4564 ( \13359_13661 , RIe1a4588_3247, \8989_9288 );
and \U$4565 ( \13360_13662 , RIe1a1888_3215, \8991_9290 );
and \U$4566 ( \13361_13663 , RIe18dd88_2991, \8993_9292 );
and \U$4567 ( \13362_13664 , RIe17a288_2767, \8995_9294 );
and \U$4568 ( \13363_13665 , RIe227be0_4742, \8997_9296 );
and \U$4569 ( \13364_13666 , RIe21c7e0_4614, \8999_9298 );
and \U$4570 ( \13365_13667 , RIe205fe0_4358, \9001_9300 );
and \U$4571 ( \13366_13668 , RIe200040_4290, \9003_9302 );
and \U$4572 ( \13367_13669 , RIe1f93f8_4213, \9005_9304 );
and \U$4573 ( \13368_13670 , RIe1f1f40_4130, \9007_9306 );
and \U$4574 ( \13369_13671 , RIe1d6448_3815, \9009_9308 );
and \U$4575 ( \13370_13672 , RIe1bcf48_3527, \9011_9310 );
and \U$4576 ( \13371_13673 , RIe1afdc0_3378, \9013_9312 );
and \U$4577 ( \13372_13674 , RIe1723f8_2677, \9015_9314 );
or \U$4578 ( \13373_13675 , \13309_13611 , \13310_13612 , \13311_13613 , \13312_13614 , \13313_13615 , \13314_13616 , \13315_13617 , \13316_13618 , \13317_13619 , \13318_13620 , \13319_13621 , \13320_13622 , \13321_13623 , \13322_13624 , \13323_13625 , \13324_13626 , \13325_13627 , \13326_13628 , \13327_13629 , \13328_13630 , \13329_13631 , \13330_13632 , \13331_13633 , \13332_13634 , \13333_13635 , \13334_13636 , \13335_13637 , \13336_13638 , \13337_13639 , \13338_13640 , \13339_13641 , \13340_13642 , \13341_13643 , \13342_13644 , \13343_13645 , \13344_13646 , \13345_13647 , \13346_13648 , \13347_13649 , \13348_13650 , \13349_13651 , \13350_13652 , \13351_13653 , \13352_13654 , \13353_13655 , \13354_13656 , \13355_13657 , \13356_13658 , \13357_13659 , \13358_13660 , \13359_13661 , \13360_13662 , \13361_13663 , \13362_13664 , \13363_13665 , \13364_13666 , \13365_13667 , \13366_13668 , \13367_13669 , \13368_13670 , \13369_13671 , \13370_13672 , \13371_13673 , \13372_13674 );
or \U$4579 ( \13374_13676 , \13308_13610 , \13373_13675 );
_DC \g658a/U$1 ( \13375 , \13374_13676 , \9024_9323 );
and g658b_GF_PartitionCandidate( \13376_13678_nG658b , \13243 , \13375 );
buf \U$4580 ( \13377_13679 , \13376_13678_nG658b );
and \U$4581 ( \13378_13680 , \13377_13679 , \10389_10691 );
nor \U$4582 ( \13379_13681 , \13111_13413 , \13378_13680 );
xnor \U$4583 ( \13380_13682 , \13379_13681 , \10678_10980 );
and \U$4584 ( \13381_13683 , \11287_11586 , \11275_11574 );
and \U$4585 ( \13382_13684 , \12146_12448 , \10976_11278 );
nor \U$4586 ( \13383_13685 , \13381_13683 , \13382_13684 );
xnor \U$4587 ( \13384_13686 , \13383_13685 , \11281_11580 );
xor \U$4588 ( \13385_13687 , \13380_13682 , \13384_13686 );
_DC \g4b10/U$1 ( \13386 , \13242_13544 , \9298_9597 );
_DC \g4b94/U$1 ( \13387 , \13374_13676 , \9024_9323 );
xor g4b95_GF_PartitionCandidate( \13388_13690_nG4b95 , \13386 , \13387 );
buf \U$4589 ( \13389_13691 , \13388_13690_nG4b95 );
xor \U$4590 ( \13390_13692 , \13389_13691 , \12478_12777 );
and \U$4591 ( \13391_13693 , \10385_10687 , \13390_13692 );
xor \U$4592 ( \13392_13694 , \13385_13687 , \13391_13693 );
xor \U$4593 ( \13393_13695 , \13110_13412 , \13392_13694 );
and \U$4594 ( \13394_13696 , \12483_12782 , \12487_12786 );
and \U$4595 ( \13395_13697 , \12487_12786 , \12495_12794 );
and \U$4596 ( \13396_13698 , \12483_12782 , \12495_12794 );
or \U$4597 ( \13397_13699 , \13394_13696 , \13395_13697 , \13396_13698 );
xor \U$4598 ( \13398_13700 , \13393_13695 , \13397_13699 );
and \U$4599 ( \13399_13701 , \12203_12502 , \12496_12795 );
and \U$4600 ( \13400_13702 , \12497_12796 , \12500_12799 );
or \U$4601 ( \13401_13703 , \13399_13701 , \13400_13702 );
xor \U$4602 ( \13402_13704 , \13398_13700 , \13401_13703 );
buf g9bfc_GF_PartitionCandidate( \13403_13705_nG9bfc , \13402_13704 );
and \U$4603 ( \13404_13706 , \10402_10704 , \13403_13705_nG9bfc );
or \U$4604 ( \13405_13707 , \13104_13406 , \13404_13706 );
xor \U$4605 ( \13406_13708 , \10399_10703 , \13405_13707 );
buf \U$4606 ( \13407_13709 , \13406_13708 );
buf \U$4608 ( \13408_13710 , \13407_13709 );
xor \U$4609 ( \13409_13711 , \13103_13405 , \13408_13710 );
buf \U$4610 ( \13410_13712 , \13409_13711 );
xor \U$4611 ( \13411_13713 , \13086_13388 , \13410_13712 );
and \U$4612 ( \13412_13714 , \12519_12818 , \13411_13713 );
and \U$4613 ( \13413_13715 , \13074_13376 , \13411_13713 );
or \U$4614 ( \13414_13716 , \13075_13377 , \13412_13714 , \13413_13715 );
and \U$4615 ( \13415_13717 , \13080_13382 , \13085_13387 );
and \U$4616 ( \13416_13718 , \13080_13382 , \13410_13712 );
and \U$4617 ( \13417_13719 , \13085_13387 , \13410_13712 );
or \U$4618 ( \13418_13720 , \13415_13717 , \13416_13718 , \13417_13719 );
buf \U$4619 ( \13419_13721 , \13418_13720 );
and \U$4620 ( \13420_13722 , \13096_13398 , \13102_13404 );
and \U$4621 ( \13421_13723 , \13096_13398 , \13408_13710 );
and \U$4622 ( \13422_13724 , \13102_13404 , \13408_13710 );
or \U$4623 ( \13423_13725 , \13420_13722 , \13421_13723 , \13422_13724 );
buf \U$4624 ( \13424_13726 , \13423_13725 );
xor \U$4625 ( \13425_13727 , \13419_13721 , \13424_13726 );
and \U$4626 ( \13426_13728 , \13067_13366 , \13071_13373 );
buf \U$4627 ( \13427_13729 , \13426_13728 );
buf \U$4629 ( \13428_13730 , \13427_13729 );
not \U$4269 ( \13429_13368 , \13068_13367 );
xor \U$4270 ( \13430_13369 , \13062_13361_nG4442 , \13065_13364_nG4445 );
and \U$4271 ( \13431_13370 , \13429_13368 , \13430_13369 );
and \U$4630 ( \13432_13731 , \13431_13370 , \10392_10694_nG9c0e );
and \U$4631 ( \13433_13732 , \13068_13367 , \10693_10995_nG9c0b );
or \U$4632 ( \13434_13733 , \13432_13731 , \13433_13732 );
xor \U$4633 ( \13435_13734 , \13067_13366 , \13434_13733 );
buf \U$4634 ( \13436_13735 , \13435_13734 );
buf \U$4636 ( \13437_13736 , \13436_13735 );
xor \U$4637 ( \13438_13737 , \13428_13730 , \13437_13736 );
buf \U$4638 ( \13439_13738 , \13438_13737 );
and \U$4639 ( \13440_13739 , \12183_12157 , \10981_11283_nG9c08 );
and \U$4640 ( \13441_13740 , \11855_12154 , \11299_11598_nG9c05 );
or \U$4641 ( \13442_13741 , \13440_13739 , \13441_13740 );
xor \U$4642 ( \13443_13742 , \11854_12153 , \13442_13741 );
buf \U$4643 ( \13444_13743 , \13443_13742 );
buf \U$4645 ( \13445_13744 , \13444_13743 );
xor \U$4646 ( \13446_13745 , \13439_13738 , \13445_13744 );
and \U$4647 ( \13447_13746 , \10996_10421 , \12168_12470_nG9c02 );
and \U$4648 ( \13448_13747 , \10119_10418 , \12502_12801_nG9bff );
or \U$4649 ( \13449_13748 , \13447_13746 , \13448_13747 );
xor \U$4650 ( \13450_13749 , \10118_10417 , \13449_13748 );
buf \U$4651 ( \13451_13750 , \13450_13749 );
buf \U$4653 ( \13452_13751 , \13451_13750 );
xor \U$4654 ( \13453_13752 , \13446_13745 , \13452_13751 );
buf \U$4655 ( \13454_13753 , \13453_13752 );
and \U$4656 ( \13455_13754 , \13088_13390 , \13094_13396 );
buf \U$4657 ( \13456_13755 , \13455_13754 );
xor \U$4658 ( \13457_13756 , \13454_13753 , \13456_13755 );
and \U$4659 ( \13458_13757 , \10411_10707 , \13403_13705_nG9bfc );
and \U$4660 ( \13459_13758 , \13377_13679 , \10681_10983 );
and \U$4661 ( \13460_13759 , RIdec6a58_724, \9034_9333 );
and \U$4662 ( \13461_13760 , RIdec3d58_692, \9036_9335 );
and \U$4663 ( \13462_13761 , RIfc723e0_6322, \9038_9337 );
and \U$4664 ( \13463_13762 , RIdec1058_660, \9040_9339 );
and \U$4665 ( \13464_13763 , RIfc59fc0_6046, \9042_9341 );
and \U$4666 ( \13465_13764 , RIdebe358_628, \9044_9343 );
and \U$4667 ( \13466_13765 , RIdebb658_596, \9046_9345 );
and \U$4668 ( \13467_13766 , RIdeb8958_564, \9048_9347 );
and \U$4669 ( \13468_13767 , RIfcb96f0_7132, \9050_9349 );
and \U$4670 ( \13469_13768 , RIdeb2f58_500, \9052_9351 );
and \U$4671 ( \13470_13769 , RIfce1c68_7591, \9054_9353 );
and \U$4672 ( \13471_13770 , RIdeb0258_468, \9056_9355 );
and \U$4673 ( \13472_13771 , RIfc9b498_6789, \9058_9357 );
and \U$4674 ( \13473_13772 , RIdead558_436, \9060_9359 );
and \U$4675 ( \13474_13773 , RIdea6fa0_404, \9062_9361 );
and \U$4676 ( \13475_13774 , RIdea06a0_372, \9064_9363 );
and \U$4677 ( \13476_13775 , RIfc81458_6493, \9066_9365 );
and \U$4678 ( \13477_13776 , RIfc83780_6518, \9068_9367 );
and \U$4679 ( \13478_13777 , RIfc4e620_5914, \9070_9369 );
and \U$4680 ( \13479_13778 , RIfcd3e38_7433, \9072_9371 );
and \U$4681 ( \13480_13779 , RIde937e8_309, \9074_9373 );
and \U$4682 ( \13481_13780 , RIde8f990_290, \9076_9375 );
and \U$4683 ( \13482_13781 , RIde8bb38_271, \9078_9377 );
and \U$4684 ( \13483_13782 , RIde87650_250, \9080_9379 );
and \U$4685 ( \13484_13783 , RIde834b0_230, \9082_9381 );
and \U$4686 ( \13485_13784 , RIfc42c80_5782, \9084_9383 );
and \U$4687 ( \13486_13785 , RIfc65960_6178, \9086_9385 );
and \U$4688 ( \13487_13786 , RIfc6c710_6256, \9088_9387 );
and \U$4689 ( \13488_13787 , RIee392b0_5109, \9090_9389 );
and \U$4690 ( \13489_13788 , RIe16cb60_2614, \9092_9391 );
and \U$4691 ( \13490_13789 , RIe16a6d0_2588, \9094_9393 );
and \U$4692 ( \13491_13790 , RIe169050_2572, \9096_9395 );
and \U$4693 ( \13492_13791 , RIe166a58_2545, \9098_9397 );
and \U$4694 ( \13493_13792 , RIe163d58_2513, \9100_9399 );
and \U$4695 ( \13494_13793 , RIfec3cf0_8348, \9102_9401 );
and \U$4696 ( \13495_13794 , RIe161058_2481, \9104_9403 );
and \U$4697 ( \13496_13795 , RIfcd54b8_7449, \9106_9405 );
and \U$4698 ( \13497_13796 , RIe15e358_2449, \9108_9407 );
and \U$4699 ( \13498_13797 , RIe158958_2385, \9110_9409 );
and \U$4700 ( \13499_13798 , RIe155c58_2353, \9112_9411 );
and \U$4701 ( \13500_13799 , RIfe9ba48_8115, \9114_9413 );
and \U$4702 ( \13501_13800 , RIe152f58_2321, \9116_9415 );
and \U$4703 ( \13502_13801 , RIfec4128_8351, \9118_9417 );
and \U$4704 ( \13503_13802 , RIe150258_2289, \9120_9419 );
and \U$4705 ( \13504_13803 , RIfcb9b28_7135, \9122_9421 );
and \U$4706 ( \13505_13804 , RIe14d558_2257, \9124_9423 );
and \U$4707 ( \13506_13805 , RIe14a858_2225, \9126_9425 );
and \U$4708 ( \13507_13806 , RIe147b58_2193, \9128_9427 );
and \U$4709 ( \13508_13807 , RIfcdb2f0_7516, \9130_9429 );
and \U$4710 ( \13509_13808 , RIfc553d0_5992, \9132_9431 );
and \U$4711 ( \13510_13809 , RIfc9a0e8_6775, \9134_9433 );
and \U$4712 ( \13511_13810 , RIfcbd908_7179, \9136_9435 );
and \U$4713 ( \13512_13811 , RIe1422c0_2130, \9138_9437 );
and \U$4714 ( \13513_13812 , RIe13ff98_2105, \9140_9439 );
and \U$4715 ( \13514_13813 , RIdf3dea0_2081, \9142_9441 );
and \U$4716 ( \13515_13814 , RIdf3ba10_2055, \9144_9443 );
and \U$4717 ( \13516_13815 , RIfc87128_6559, \9146_9445 );
and \U$4718 ( \13517_13816 , RIee304a8_5008, \9148_9447 );
and \U$4719 ( \13518_13817 , RIfcc51f8_7265, \9150_9449 );
and \U$4720 ( \13519_13818 , RIee2e2e8_4984, \9152_9451 );
and \U$4721 ( \13520_13819 , RIdf36cb8_2000, \9154_9453 );
and \U$4722 ( \13521_13820 , RIfec3fc0_8350, \9156_9455 );
and \U$4723 ( \13522_13821 , RIdf32500_1949, \9158_9457 );
and \U$4724 ( \13523_13822 , RIfec3e58_8349, \9160_9459 );
or \U$4725 ( \13524_13823 , \13460_13759 , \13461_13760 , \13462_13761 , \13463_13762 , \13464_13763 , \13465_13764 , \13466_13765 , \13467_13766 , \13468_13767 , \13469_13768 , \13470_13769 , \13471_13770 , \13472_13771 , \13473_13772 , \13474_13773 , \13475_13774 , \13476_13775 , \13477_13776 , \13478_13777 , \13479_13778 , \13480_13779 , \13481_13780 , \13482_13781 , \13483_13782 , \13484_13783 , \13485_13784 , \13486_13785 , \13487_13786 , \13488_13787 , \13489_13788 , \13490_13789 , \13491_13790 , \13492_13791 , \13493_13792 , \13494_13793 , \13495_13794 , \13496_13795 , \13497_13796 , \13498_13797 , \13499_13798 , \13500_13799 , \13501_13800 , \13502_13801 , \13503_13802 , \13504_13803 , \13505_13804 , \13506_13805 , \13507_13806 , \13508_13807 , \13509_13808 , \13510_13809 , \13511_13810 , \13512_13811 , \13513_13812 , \13514_13813 , \13515_13814 , \13516_13815 , \13517_13816 , \13518_13817 , \13519_13818 , \13520_13819 , \13521_13820 , \13522_13821 , \13523_13822 );
and \U$4726 ( \13525_13824 , RIee2c830_4965, \9163_9462 );
and \U$4727 ( \13526_13825 , RIee2ad78_4946, \9165_9464 );
and \U$4728 ( \13527_13826 , RIee296f8_4930, \9167_9466 );
and \U$4729 ( \13528_13827 , RIee284b0_4917, \9169_9468 );
and \U$4730 ( \13529_13828 , RIfe9b8e0_8114, \9171_9470 );
and \U$4731 ( \13530_13829 , RIfe9b610_8112, \9173_9472 );
and \U$4732 ( \13531_13830 , RIfe9b778_8113, \9175_9474 );
and \U$4733 ( \13532_13831 , RIfe9b4a8_8111, \9177_9476 );
and \U$4734 ( \13533_13832 , RIfcb7c38_7113, \9179_9478 );
and \U$4735 ( \13534_13833 , RIfc86b88_6555, \9181_9480 );
and \U$4736 ( \13535_13834 , RIdf238c0_1781, \9183_9482 );
and \U$4737 ( \13536_13835 , RIfc75ab8_6361, \9185_9484 );
and \U$4738 ( \13537_13836 , RIdf22240_1765, \9187_9486 );
and \U$4739 ( \13538_13837 , RIfeaa3b8_8253, \9189_9488 );
and \U$4740 ( \13539_13838 , RIdf1bb98_1692, \9191_9490 );
and \U$4741 ( \13540_13839 , RIdf1a680_1677, \9193_9492 );
and \U$4742 ( \13541_13840 , RIdf18628_1654, \9195_9494 );
and \U$4743 ( \13542_13841 , RIdf15928_1622, \9197_9496 );
and \U$4744 ( \13543_13842 , RIdf12c28_1590, \9199_9498 );
and \U$4745 ( \13544_13843 , RIdf0ff28_1558, \9201_9500 );
and \U$4746 ( \13545_13844 , RIdf0d228_1526, \9203_9502 );
and \U$4747 ( \13546_13845 , RIdf0a528_1494, \9205_9504 );
and \U$4748 ( \13547_13846 , RIdf07828_1462, \9207_9506 );
and \U$4749 ( \13548_13847 , RIdf04b28_1430, \9209_9508 );
and \U$4750 ( \13549_13848 , RIdeff128_1366, \9211_9510 );
and \U$4751 ( \13550_13849 , RIdefc428_1334, \9213_9512 );
and \U$4752 ( \13551_13850 , RIdef9728_1302, \9215_9514 );
and \U$4753 ( \13552_13851 , RIdef6a28_1270, \9217_9516 );
and \U$4754 ( \13553_13852 , RIdef3d28_1238, \9219_9518 );
and \U$4755 ( \13554_13853 , RIdef1028_1206, \9221_9520 );
and \U$4756 ( \13555_13854 , RIdeee328_1174, \9223_9522 );
and \U$4757 ( \13556_13855 , RIdeeb628_1142, \9225_9524 );
and \U$4758 ( \13557_13856 , RIee25a80_4887, \9227_9526 );
and \U$4759 ( \13558_13857 , RIee24c70_4877, \9229_9528 );
and \U$4760 ( \13559_13858 , RIfcddd20_7546, \9231_9530 );
and \U$4761 ( \13560_13859 , RIfccc110_7344, \9233_9532 );
and \U$4762 ( \13561_13860 , RIdee5c28_1078, \9235_9534 );
and \U$4763 ( \13562_13861 , RIdee3ea0_1057, \9237_9536 );
and \U$4764 ( \13563_13862 , RIdee1b78_1032, \9239_9538 );
and \U$4765 ( \13564_13863 , RIdedfc88_1010, \9241_9540 );
and \U$4766 ( \13565_13864 , RIfc6a6b8_6233, \9243_9542 );
and \U$4767 ( \13566_13865 , RIee227e0_4851, \9245_9544 );
and \U$4768 ( \13567_13866 , RIfc88be0_6578, \9247_9546 );
and \U$4769 ( \13568_13867 , RIee21868_4840, \9249_9548 );
and \U$4770 ( \13569_13868 , RIdedaaf8_952, \9251_9550 );
and \U$4771 ( \13570_13869 , RIded8668_926, \9253_9552 );
and \U$4772 ( \13571_13870 , RIded6340_901, \9255_9554 );
and \U$4773 ( \13572_13871 , RIded4180_877, \9257_9556 );
and \U$4774 ( \13573_13872 , RIded1e58_852, \9259_9558 );
and \U$4775 ( \13574_13873 , RIdecf158_820, \9261_9560 );
and \U$4776 ( \13575_13874 , RIdecc458_788, \9263_9562 );
and \U$4777 ( \13576_13875 , RIdec9758_756, \9265_9564 );
and \U$4778 ( \13577_13876 , RIdeb5c58_532, \9267_9566 );
and \U$4779 ( \13578_13877 , RIde99da0_340, \9269_9568 );
and \U$4780 ( \13579_13878 , RIe16f860_2646, \9271_9570 );
and \U$4781 ( \13580_13879 , RIe15b658_2417, \9273_9572 );
and \U$4782 ( \13581_13880 , RIe144e58_2161, \9275_9574 );
and \U$4783 ( \13582_13881 , RIdf39850_2031, \9277_9576 );
and \U$4784 ( \13583_13882 , RIdf2deb0_1899, \9279_9578 );
and \U$4785 ( \13584_13883 , RIdf1e730_1723, \9281_9580 );
and \U$4786 ( \13585_13884 , RIdf01e28_1398, \9283_9582 );
and \U$4787 ( \13586_13885 , RIdee8928_1110, \9285_9584 );
and \U$4788 ( \13587_13886 , RIdedd690_983, \9287_9586 );
and \U$4789 ( \13588_13887 , RIde7fce8_213, \9289_9588 );
or \U$4790 ( \13589_13888 , \13525_13824 , \13526_13825 , \13527_13826 , \13528_13827 , \13529_13828 , \13530_13829 , \13531_13830 , \13532_13831 , \13533_13832 , \13534_13833 , \13535_13834 , \13536_13835 , \13537_13836 , \13538_13837 , \13539_13838 , \13540_13839 , \13541_13840 , \13542_13841 , \13543_13842 , \13544_13843 , \13545_13844 , \13546_13845 , \13547_13846 , \13548_13847 , \13549_13848 , \13550_13849 , \13551_13850 , \13552_13851 , \13553_13852 , \13554_13853 , \13555_13854 , \13556_13855 , \13557_13856 , \13558_13857 , \13559_13858 , \13560_13859 , \13561_13860 , \13562_13861 , \13563_13862 , \13564_13863 , \13565_13864 , \13566_13865 , \13567_13866 , \13568_13867 , \13569_13868 , \13570_13869 , \13571_13870 , \13572_13871 , \13573_13872 , \13574_13873 , \13575_13874 , \13576_13875 , \13577_13876 , \13578_13877 , \13579_13878 , \13580_13879 , \13581_13880 , \13582_13881 , \13583_13882 , \13584_13883 , \13585_13884 , \13586_13885 , \13587_13886 , \13588_13887 );
or \U$4791 ( \13590_13889 , \13524_13823 , \13589_13888 );
_DC \g658c/U$1 ( \13591 , \13590_13889 , \9298_9597 );
and \U$4792 ( \13592_13891 , RIe19ecf0_3184, \8760_9059 );
and \U$4793 ( \13593_13892 , RIe19bff0_3152, \8762_9061 );
and \U$4794 ( \13594_13893 , RIf145a90_5252, \8764_9063 );
and \U$4795 ( \13595_13894 , RIe1992f0_3120, \8766_9065 );
and \U$4796 ( \13596_13895 , RIf144de8_5243, \8768_9067 );
and \U$4797 ( \13597_13896 , RIe1965f0_3088, \8770_9069 );
and \U$4798 ( \13598_13897 , RIe1938f0_3056, \8772_9071 );
and \U$4799 ( \13599_13898 , RIe190bf0_3024, \8774_9073 );
and \U$4800 ( \13600_13899 , RIe18b1f0_2960, \8776_9075 );
and \U$4801 ( \13601_13900 , RIe1884f0_2928, \8778_9077 );
and \U$4802 ( \13602_13901 , RIfc72980_6326, \8780_9079 );
and \U$4803 ( \13603_13902 , RIe1857f0_2896, \8782_9081 );
and \U$4804 ( \13604_13903 , RIf143060_5222, \8784_9083 );
and \U$4805 ( \13605_13904 , RIe182af0_2864, \8786_9085 );
and \U$4806 ( \13606_13905 , RIe17fdf0_2832, \8788_9087 );
and \U$4807 ( \13607_13906 , RIe17d0f0_2800, \8790_9089 );
and \U$4808 ( \13608_13907 , RIf142688_5215, \8792_9091 );
and \U$4809 ( \13609_13908 , RIf141710_5204, \8794_9093 );
and \U$4810 ( \13610_13909 , RIe177858_2737, \8796_9095 );
and \U$4811 ( \13611_13910 , RIe176778_2725, \8798_9097 );
and \U$4812 ( \13612_13911 , RIfcea638_7689, \8800_9099 );
and \U$4813 ( \13613_13912 , RIfca54e8_6903, \8802_9101 );
and \U$4814 ( \13614_13913 , RIee3e878_5170, \8804_9103 );
and \U$4815 ( \13615_13914 , RIee3dbd0_5161, \8806_9105 );
and \U$4816 ( \13616_13915 , RIee3c988_5148, \8808_9107 );
and \U$4817 ( \13617_13916 , RIee3b5d8_5134, \8810_9109 );
and \U$4818 ( \13618_13917 , RIee3a4f8_5122, \8812_9111 );
and \U$4819 ( \13619_13918 , RIe174b58_2705, \8814_9113 );
and \U$4820 ( \13620_13919 , RIf170600_5738, \8816_9115 );
and \U$4821 ( \13621_13920 , RIfc76fd0_6376, \8818_9117 );
and \U$4822 ( \13622_13921 , RIf16e9e0_5718, \8820_9119 );
and \U$4823 ( \13623_13922 , RIfced608_7723, \8822_9121 );
and \U$4824 ( \13624_13923 , RIf16d090_5700, \8824_9123 );
and \U$4825 ( \13625_13924 , RIe225048_4711, \8826_9125 );
and \U$4826 ( \13626_13925 , RIf16c550_5692, \8828_9127 );
and \U$4827 ( \13627_13926 , RIe222348_4679, \8830_9129 );
and \U$4828 ( \13628_13927 , RIf16b470_5680, \8832_9131 );
and \U$4829 ( \13629_13928 , RIe21f648_4647, \8834_9133 );
and \U$4830 ( \13630_13929 , RIe219c48_4583, \8836_9135 );
and \U$4831 ( \13631_13930 , RIe216f48_4551, \8838_9137 );
and \U$4832 ( \13632_13931 , RIf16a4f8_5669, \8840_9139 );
and \U$4833 ( \13633_13932 , RIe214248_4519, \8842_9141 );
and \U$4834 ( \13634_13933 , RIf169df0_5664, \8844_9143 );
and \U$4835 ( \13635_13934 , RIe211548_4487, \8846_9145 );
and \U$4836 ( \13636_13935 , RIf1684a0_5646, \8848_9147 );
and \U$4837 ( \13637_13936 , RIe20e848_4455, \8850_9149 );
and \U$4838 ( \13638_13937 , RIe20bb48_4423, \8852_9151 );
and \U$4839 ( \13639_13938 , RIe208e48_4391, \8854_9153 );
and \U$4840 ( \13640_13939 , RIf1673c0_5634, \8856_9155 );
and \U$4841 ( \13641_13940 , RIf166448_5623, \8858_9157 );
and \U$4842 ( \13642_13941 , RIfe9c6f0_8124, \8860_9159 );
and \U$4843 ( \13643_13942 , RIfe9c150_8120, \8862_9161 );
and \U$4844 ( \13644_13943 , RIf1654d0_5612, \8864_9163 );
and \U$4845 ( \13645_13944 , RIfcc4550_7256, \8866_9165 );
and \U$4846 ( \13646_13945 , RIf1635e0_5590, \8868_9167 );
and \U$4847 ( \13647_13946 , RIf162500_5578, \8870_9169 );
and \U$4848 ( \13648_13947 , RIf160fe8_5563, \8872_9171 );
and \U$4849 ( \13649_13948 , RIf15f0f8_5541, \8874_9173 );
and \U$4850 ( \13650_13949 , RIfe9bfe8_8119, \8876_9175 );
and \U$4851 ( \13651_13950 , RIfe9c588_8123, \8878_9177 );
and \U$4852 ( \13652_13951 , RIf15d208_5519, \8880_9179 );
and \U$4853 ( \13653_13952 , RIf15bfc0_5506, \8882_9181 );
and \U$4854 ( \13654_13953 , RIfc4d540_5902, \8884_9183 );
and \U$4855 ( \13655_13954 , RIfc9c848_6803, \8886_9185 );
or \U$4856 ( \13656_13955 , \13592_13891 , \13593_13892 , \13594_13893 , \13595_13894 , \13596_13895 , \13597_13896 , \13598_13897 , \13599_13898 , \13600_13899 , \13601_13900 , \13602_13901 , \13603_13902 , \13604_13903 , \13605_13904 , \13606_13905 , \13607_13906 , \13608_13907 , \13609_13908 , \13610_13909 , \13611_13910 , \13612_13911 , \13613_13912 , \13614_13913 , \13615_13914 , \13616_13915 , \13617_13916 , \13618_13917 , \13619_13918 , \13620_13919 , \13621_13920 , \13622_13921 , \13623_13922 , \13624_13923 , \13625_13924 , \13626_13925 , \13627_13926 , \13628_13927 , \13629_13928 , \13630_13929 , \13631_13930 , \13632_13931 , \13633_13932 , \13634_13933 , \13635_13934 , \13636_13935 , \13637_13936 , \13638_13937 , \13639_13938 , \13640_13939 , \13641_13940 , \13642_13941 , \13643_13942 , \13644_13943 , \13645_13944 , \13646_13945 , \13647_13946 , \13648_13947 , \13649_13948 , \13650_13949 , \13651_13950 , \13652_13951 , \13653_13952 , \13654_13953 , \13655_13954 );
and \U$4857 ( \13657_13956 , RIfec4290_8352, \8889_9188 );
and \U$4858 ( \13658_13957 , RIfe9c2b8_8121, \8891_9190 );
and \U$4859 ( \13659_13958 , RIfcc01d0_7208, \8893_9192 );
and \U$4860 ( \13660_13959 , RIe1fb2e8_4235, \8895_9194 );
and \U$4861 ( \13661_13960 , RIfe9c420_8122, \8897_9196 );
and \U$4862 ( \13662_13961 , RIfca3e68_6887, \8899_9198 );
and \U$4863 ( \13663_13962 , RIf154c70_5424, \8901_9200 );
and \U$4864 ( \13664_13963 , RIe1f69c8_4183, \8903_9202 );
and \U$4865 ( \13665_13964 , RIf153a28_5411, \8905_9204 );
and \U$4866 ( \13666_13965 , RIf152240_5394, \8907_9206 );
and \U$4867 ( \13667_13966 , RIf150ff8_5381, \8909_9208 );
and \U$4868 ( \13668_13967 , RIe1f46a0_4158, \8911_9210 );
and \U$4869 ( \13669_13968 , RIfca6028_6911, \8913_9212 );
and \U$4870 ( \13670_13969 , RIfc43bf8_5793, \8915_9214 );
and \U$4871 ( \13671_13970 , RIf14e460_5350, \8917_9216 );
and \U$4872 ( \13672_13971 , RIe1ef3a8_4099, \8919_9218 );
and \U$4873 ( \13673_13972 , RIe1ecdb0_4072, \8921_9220 );
and \U$4874 ( \13674_13973 , RIe1ea0b0_4040, \8923_9222 );
and \U$4875 ( \13675_13974 , RIe1e73b0_4008, \8925_9224 );
and \U$4876 ( \13676_13975 , RIe1e46b0_3976, \8927_9226 );
and \U$4877 ( \13677_13976 , RIe1e19b0_3944, \8929_9228 );
and \U$4878 ( \13678_13977 , RIe1decb0_3912, \8931_9230 );
and \U$4879 ( \13679_13978 , RIe1dbfb0_3880, \8933_9232 );
and \U$4880 ( \13680_13979 , RIe1d92b0_3848, \8935_9234 );
and \U$4881 ( \13681_13980 , RIe1d38b0_3784, \8937_9236 );
and \U$4882 ( \13682_13981 , RIe1d0bb0_3752, \8939_9238 );
and \U$4883 ( \13683_13982 , RIe1cdeb0_3720, \8941_9240 );
and \U$4884 ( \13684_13983 , RIe1cb1b0_3688, \8943_9242 );
and \U$4885 ( \13685_13984 , RIe1c84b0_3656, \8945_9244 );
and \U$4886 ( \13686_13985 , RIe1c57b0_3624, \8947_9246 );
and \U$4887 ( \13687_13986 , RIe1c2ab0_3592, \8949_9248 );
and \U$4888 ( \13688_13987 , RIe1bfdb0_3560, \8951_9250 );
and \U$4889 ( \13689_13988 , RIfc4d6a8_5903, \8953_9252 );
and \U$4890 ( \13690_13989 , RIf14be68_5323, \8955_9254 );
and \U$4891 ( \13691_13990 , RIe1ba680_3498, \8957_9256 );
and \U$4892 ( \13692_13991 , RIfe9be80_8118, \8959_9258 );
and \U$4893 ( \13693_13992 , RIfc86e58_6557, \8961_9260 );
and \U$4894 ( \13694_13993 , RIfcd46a8_7439, \8963_9262 );
and \U$4895 ( \13695_13994 , RIe1b6300_3450, \8965_9264 );
and \U$4896 ( \13696_13995 , RIfe9bd18_8117, \8967_9266 );
and \U$4897 ( \13697_13996 , RIf1495a0_5294, \8969_9268 );
and \U$4898 ( \13698_13997 , RIf1481f0_5280, \8971_9270 );
and \U$4899 ( \13699_13998 , RIe1b3600_3418, \8973_9272 );
and \U$4900 ( \13700_13999 , RIe1b1e18_3401, \8975_9274 );
and \U$4901 ( \13701_14000 , RIfc69470_6220, \8977_9276 );
and \U$4902 ( \13702_14001 , RIfcbfac8_7203, \8979_9278 );
and \U$4903 ( \13703_14002 , RIfe9bbb0_8116, \8981_9280 );
and \U$4904 ( \13704_14003 , RIe1abd10_3332, \8983_9282 );
and \U$4905 ( \13705_14004 , RIe1aa0f0_3312, \8985_9284 );
and \U$4906 ( \13706_14005 , RIe1a73f0_3280, \8987_9286 );
and \U$4907 ( \13707_14006 , RIe1a46f0_3248, \8989_9288 );
and \U$4908 ( \13708_14007 , RIe1a19f0_3216, \8991_9290 );
and \U$4909 ( \13709_14008 , RIe18def0_2992, \8993_9292 );
and \U$4910 ( \13710_14009 , RIe17a3f0_2768, \8995_9294 );
and \U$4911 ( \13711_14010 , RIe227d48_4743, \8997_9296 );
and \U$4912 ( \13712_14011 , RIe21c948_4615, \8999_9298 );
and \U$4913 ( \13713_14012 , RIe206148_4359, \9001_9300 );
and \U$4914 ( \13714_14013 , RIe2001a8_4291, \9003_9302 );
and \U$4915 ( \13715_14014 , RIe1f9560_4214, \9005_9304 );
and \U$4916 ( \13716_14015 , RIe1f20a8_4131, \9007_9306 );
and \U$4917 ( \13717_14016 , RIe1d65b0_3816, \9009_9308 );
and \U$4918 ( \13718_14017 , RIe1bd0b0_3528, \9011_9310 );
and \U$4919 ( \13719_14018 , RIe1aff28_3379, \9013_9312 );
and \U$4920 ( \13720_14019 , RIe172560_2678, \9015_9314 );
or \U$4921 ( \13721_14020 , \13657_13956 , \13658_13957 , \13659_13958 , \13660_13959 , \13661_13960 , \13662_13961 , \13663_13962 , \13664_13963 , \13665_13964 , \13666_13965 , \13667_13966 , \13668_13967 , \13669_13968 , \13670_13969 , \13671_13970 , \13672_13971 , \13673_13972 , \13674_13973 , \13675_13974 , \13676_13975 , \13677_13976 , \13678_13977 , \13679_13978 , \13680_13979 , \13681_13980 , \13682_13981 , \13683_13982 , \13684_13983 , \13685_13984 , \13686_13985 , \13687_13986 , \13688_13987 , \13689_13988 , \13690_13989 , \13691_13990 , \13692_13991 , \13693_13992 , \13694_13993 , \13695_13994 , \13696_13995 , \13697_13996 , \13698_13997 , \13699_13998 , \13700_13999 , \13701_14000 , \13702_14001 , \13703_14002 , \13704_14003 , \13705_14004 , \13706_14005 , \13707_14006 , \13708_14007 , \13709_14008 , \13710_14009 , \13711_14010 , \13712_14011 , \13713_14012 , \13714_14013 , \13715_14014 , \13716_14015 , \13717_14016 , \13718_14017 , \13719_14018 , \13720_14019 );
or \U$4922 ( \13722_14021 , \13656_13955 , \13721_14020 );
_DC \g658d/U$1 ( \13723 , \13722_14021 , \9024_9323 );
and g658e_GF_PartitionCandidate( \13724_14023_nG658e , \13591 , \13723 );
buf \U$4923 ( \13725_14024 , \13724_14023_nG658e );
and \U$4924 ( \13726_14025 , \13725_14024 , \10389_10691 );
nor \U$4925 ( \13727_14026 , \13459_13758 , \13726_14025 );
xnor \U$4926 ( \13728_14027 , \13727_14026 , \10678_10980 );
not \U$4927 ( \13729_14028 , \13391_13693 );
_DC \g4c19/U$1 ( \13730 , \13590_13889 , \9298_9597 );
_DC \g4c9d/U$1 ( \13731 , \13722_14021 , \9024_9323 );
xor g4c9e_GF_PartitionCandidate( \13732_14031_nG4c9e , \13730 , \13731 );
buf \U$4928 ( \13733_14032 , \13732_14031_nG4c9e );
and \U$4929 ( \13734_14033 , \13389_13691 , \12478_12777 );
not \U$4930 ( \13735_14034 , \13734_14033 );
and \U$4931 ( \13736_14035 , \13733_14032 , \13735_14034 );
and \U$4932 ( \13737_14036 , \13729_14028 , \13736_14035 );
xor \U$4933 ( \13738_14037 , \13728_14027 , \13737_14036 );
and \U$4934 ( \13739_14038 , \13380_13682 , \13384_13686 );
and \U$4935 ( \13740_14039 , \13384_13686 , \13391_13693 );
and \U$4936 ( \13741_14040 , \13380_13682 , \13391_13693 );
or \U$4937 ( \13742_14041 , \13739_14038 , \13740_14039 , \13741_14040 );
xor \U$4938 ( \13743_14042 , \13738_14037 , \13742_14041 );
and \U$4939 ( \13744_14043 , \12146_12448 , \11275_11574 );
and \U$4940 ( \13745_14044 , \12470_12769 , \10976_11278 );
nor \U$4941 ( \13746_14045 , \13744_14043 , \13745_14044 );
xnor \U$4942 ( \13747_14046 , \13746_14045 , \11281_11580 );
and \U$4943 ( \13748_14047 , \10968_11270 , \12491_12790 );
and \U$4944 ( \13749_14048 , \11287_11586 , \12159_12461 );
nor \U$4945 ( \13750_14049 , \13748_14047 , \13749_14048 );
xnor \U$4946 ( \13751_14050 , \13750_14049 , \12481_12780 );
xor \U$4947 ( \13752_14051 , \13747_14046 , \13751_14050 );
xor \U$4948 ( \13753_14052 , \13733_14032 , \13389_13691 );
not \U$4949 ( \13754_14053 , \13390_13692 );
and \U$4950 ( \13755_14054 , \13753_14052 , \13754_14053 );
and \U$4951 ( \13756_14055 , \10385_10687 , \13755_14054 );
and \U$4952 ( \13757_14056 , \10686_10988 , \13390_13692 );
nor \U$4953 ( \13758_14057 , \13756_14055 , \13757_14056 );
xnor \U$4954 ( \13759_14058 , \13758_14057 , \13736_14035 );
xor \U$4955 ( \13760_14059 , \13752_14051 , \13759_14058 );
xor \U$4956 ( \13761_14060 , \13743_14042 , \13760_14059 );
and \U$4957 ( \13762_14061 , \13105_13407 , \13109_13411 );
and \U$4958 ( \13763_14062 , \13109_13411 , \13392_13694 );
and \U$4959 ( \13764_14063 , \13105_13407 , \13392_13694 );
or \U$4960 ( \13765_14064 , \13762_14061 , \13763_14062 , \13764_14063 );
xor \U$4961 ( \13766_14065 , \13761_14060 , \13765_14064 );
and \U$4962 ( \13767_14066 , \13393_13695 , \13397_13699 );
and \U$4963 ( \13768_14067 , \13398_13700 , \13401_13703 );
or \U$4964 ( \13769_14068 , \13767_14066 , \13768_14067 );
xor \U$4965 ( \13770_14069 , \13766_14065 , \13769_14068 );
buf g9bf9_GF_PartitionCandidate( \13771_14070_nG9bf9 , \13770_14069 );
and \U$4966 ( \13772_14071 , \10402_10704 , \13771_14070_nG9bf9 );
or \U$4967 ( \13773_14072 , \13458_13757 , \13772_14071 );
xor \U$4968 ( \13774_14073 , \10399_10703 , \13773_14072 );
buf \U$4969 ( \13775_14074 , \13774_14073 );
buf \U$4971 ( \13776_14075 , \13775_14074 );
xor \U$4972 ( \13777_14076 , \13457_13756 , \13776_14075 );
buf \U$4973 ( \13778_14077 , \13777_14076 );
xor \U$4974 ( \13779_14078 , \13425_13727 , \13778_14077 );
and \U$4975 ( \13780_14079 , \13414_13716 , \13779_14078 );
and \U$4976 ( \13781_14080 , RIdec6d28_726, \8760_9059 );
and \U$4977 ( \13782_14081 , RIdec4028_694, \8762_9061 );
and \U$4978 ( \13783_14082 , RIee20bc0_4831, \8764_9063 );
and \U$4979 ( \13784_14083 , RIdec1328_662, \8766_9065 );
and \U$4980 ( \13785_14084 , RIfcbaed8_7149, \8768_9067 );
and \U$4981 ( \13786_14085 , RIdebe628_630, \8770_9069 );
and \U$4982 ( \13787_14086 , RIdebb928_598, \8772_9071 );
and \U$4983 ( \13788_14087 , RIdeb8c28_566, \8774_9073 );
and \U$4984 ( \13789_14088 , RIfc412b8_5767, \8776_9075 );
and \U$4985 ( \13790_14089 , RIdeb3228_502, \8778_9077 );
and \U$4986 ( \13791_14090 , RIfc9ea08_6827, \8780_9079 );
and \U$4987 ( \13792_14091 , RIdeb0528_470, \8782_9081 );
and \U$4988 ( \13793_14092 , RIee1e028_4800, \8784_9083 );
and \U$4989 ( \13794_14093 , RIdead828_438, \8786_9085 );
and \U$4990 ( \13795_14094 , RIdea7630_406, \8788_9087 );
and \U$4991 ( \13796_14095 , RIdea0d30_374, \8790_9089 );
and \U$4992 ( \13797_14096 , RIfcbac08_7147, \8792_9091 );
and \U$4993 ( \13798_14097 , RIfc55538_5993, \8794_9093 );
and \U$4994 ( \13799_14098 , RIfcba668_7143, \8796_9095 );
and \U$4995 ( \13800_14099 , RIfc4af48_5875, \8798_9097 );
and \U$4996 ( \13801_14100 , RIfe912f0_7996, \8800_9099 );
and \U$4997 ( \13802_14101 , RIfe91458_7997, \8802_9101 );
and \U$4998 ( \13803_14102 , RIde8be80_272, \8804_9103 );
and \U$4999 ( \13804_14103 , RIde87ce0_252, \8806_9105 );
and \U$5000 ( \13805_14104 , RIfc85238_6537, \8808_9107 );
and \U$5001 ( \13806_14105 , RIfc88640_6574, \8810_9109 );
and \U$5002 ( \13807_14106 , RIfcda210_7504, \8812_9111 );
and \U$5003 ( \13808_14107 , RIfcd5788_7451, \8814_9113 );
and \U$5004 ( \13809_14108 , RIee39418_5110, \8816_9115 );
and \U$5005 ( \13810_14109 , RIe16ce30_2616, \8818_9117 );
and \U$5006 ( \13811_14110 , RIfc884d8_6573, \8820_9119 );
and \U$5007 ( \13812_14111 , RIe169320_2574, \8822_9121 );
and \U$5008 ( \13813_14112 , RIe166d28_2547, \8824_9123 );
and \U$5009 ( \13814_14113 , RIe164028_2515, \8826_9125 );
and \U$5010 ( \13815_14114 , RIfe90918_7989, \8828_9127 );
and \U$5011 ( \13816_14115 , RIe161328_2483, \8830_9129 );
and \U$5012 ( \13817_14116 , RIee36880_5079, \8832_9131 );
and \U$5013 ( \13818_14117 , RIe15e628_2451, \8834_9133 );
and \U$5014 ( \13819_14118 , RIe158c28_2387, \8836_9135 );
and \U$5015 ( \13820_14119 , RIe155f28_2355, \8838_9137 );
and \U$5016 ( \13821_14120 , RIfe91188_7995, \8840_9139 );
and \U$5017 ( \13822_14121 , RIe153228_2323, \8842_9141 );
and \U$5018 ( \13823_14122 , RIfe91020_7994, \8844_9143 );
and \U$5019 ( \13824_14123 , RIe150528_2291, \8846_9145 );
and \U$5020 ( \13825_14124 , RIfcda378_7505, \8848_9147 );
and \U$5021 ( \13826_14125 , RIe14d828_2259, \8850_9149 );
and \U$5022 ( \13827_14126 , RIe14ab28_2227, \8852_9151 );
and \U$5023 ( \13828_14127 , RIe147e28_2195, \8854_9153 );
and \U$5024 ( \13829_14128 , RIfe90eb8_7993, \8856_9155 );
and \U$5025 ( \13830_14129 , RIfe90d50_7992, \8858_9157 );
and \U$5026 ( \13831_14130 , RIfcb99c0_7134, \8860_9159 );
and \U$5027 ( \13832_14131 , RIfc9c2a8_6799, \8862_9161 );
and \U$5028 ( \13833_14132 , RIfe90be8_7991, \8864_9163 );
and \U$5029 ( \13834_14133 , RIfe90a80_7990, \8866_9165 );
and \U$5030 ( \13835_14134 , RIdf3e008_2082, \8868_9167 );
and \U$5031 ( \13836_14135 , RIdf3bce0_2057, \8870_9169 );
and \U$5032 ( \13837_14136 , RIfcec690_7712, \8872_9171 );
and \U$5033 ( \13838_14137 , RIee30778_5010, \8874_9173 );
and \U$5034 ( \13839_14138 , RIfc87dd0_6568, \8876_9175 );
and \U$5035 ( \13840_14139 , RIee2e5b8_4986, \8878_9177 );
and \U$5036 ( \13841_14140 , RIdf36e20_2001, \8880_9179 );
and \U$5037 ( \13842_14141 , RIdf346c0_1973, \8882_9181 );
and \U$5038 ( \13843_14142 , RIdf32668_1950, \8884_9183 );
and \U$5039 ( \13844_14143 , RIdf30070_1923, \8886_9185 );
or \U$5040 ( \13845_14144 , \13781_14080 , \13782_14081 , \13783_14082 , \13784_14083 , \13785_14084 , \13786_14085 , \13787_14086 , \13788_14087 , \13789_14088 , \13790_14089 , \13791_14090 , \13792_14091 , \13793_14092 , \13794_14093 , \13795_14094 , \13796_14095 , \13797_14096 , \13798_14097 , \13799_14098 , \13800_14099 , \13801_14100 , \13802_14101 , \13803_14102 , \13804_14103 , \13805_14104 , \13806_14105 , \13807_14106 , \13808_14107 , \13809_14108 , \13810_14109 , \13811_14110 , \13812_14111 , \13813_14112 , \13814_14113 , \13815_14114 , \13816_14115 , \13817_14116 , \13818_14117 , \13819_14118 , \13820_14119 , \13821_14120 , \13822_14121 , \13823_14122 , \13824_14123 , \13825_14124 , \13826_14125 , \13827_14126 , \13828_14127 , \13829_14128 , \13830_14129 , \13831_14130 , \13832_14131 , \13833_14132 , \13834_14133 , \13835_14134 , \13836_14135 , \13837_14136 , \13838_14137 , \13839_14138 , \13840_14139 , \13841_14140 , \13842_14141 , \13843_14142 , \13844_14143 );
and \U$5041 ( \13846_14145 , RIee2c998_4966, \8889_9188 );
and \U$5042 ( \13847_14146 , RIee2aee0_4947, \8891_9190 );
and \U$5043 ( \13848_14147 , RIee299c8_4932, \8893_9192 );
and \U$5044 ( \13849_14148 , RIee28618_4918, \8895_9194 );
and \U$5045 ( \13850_14149 , RIfe90378_7985, \8897_9196 );
and \U$5046 ( \13851_14150 , RIfe907b0_7988, \8899_9198 );
and \U$5047 ( \13852_14151 , RIfe904e0_7986, \8901_9200 );
and \U$5048 ( \13853_14152 , RIfe90648_7987, \8903_9202 );
and \U$5049 ( \13854_14153 , RIfc9d928_6815, \8905_9204 );
and \U$5050 ( \13855_14154 , RIfc86048_6547, \8907_9206 );
and \U$5051 ( \13856_14155 , RIfcb92b8_7129, \8909_9208 );
and \U$5052 ( \13857_14156 , RIfc4ee90_5920, \8911_9210 );
and \U$5053 ( \13858_14157 , RIfc86a20_6554, \8913_9212 );
and \U$5054 ( \13859_14158 , RIdf20e90_1751, \8915_9214 );
and \U$5055 ( \13860_14159 , RIfcb8fe8_7127, \8917_9216 );
and \U$5056 ( \13861_14160 , RIdf1a950_1679, \8919_9218 );
and \U$5057 ( \13862_14161 , RIdf188f8_1656, \8921_9220 );
and \U$5058 ( \13863_14162 , RIdf15bf8_1624, \8923_9222 );
and \U$5059 ( \13864_14163 , RIdf12ef8_1592, \8925_9224 );
and \U$5060 ( \13865_14164 , RIdf101f8_1560, \8927_9226 );
and \U$5061 ( \13866_14165 , RIdf0d4f8_1528, \8929_9228 );
and \U$5062 ( \13867_14166 , RIdf0a7f8_1496, \8931_9230 );
and \U$5063 ( \13868_14167 , RIdf07af8_1464, \8933_9232 );
and \U$5064 ( \13869_14168 , RIdf04df8_1432, \8935_9234 );
and \U$5065 ( \13870_14169 , RIdeff3f8_1368, \8937_9236 );
and \U$5066 ( \13871_14170 , RIdefc6f8_1336, \8939_9238 );
and \U$5067 ( \13872_14171 , RIdef99f8_1304, \8941_9240 );
and \U$5068 ( \13873_14172 , RIdef6cf8_1272, \8943_9242 );
and \U$5069 ( \13874_14173 , RIdef3ff8_1240, \8945_9244 );
and \U$5070 ( \13875_14174 , RIdef12f8_1208, \8947_9246 );
and \U$5071 ( \13876_14175 , RIdeee5f8_1176, \8949_9248 );
and \U$5072 ( \13877_14176 , RIdeeb8f8_1144, \8951_9250 );
and \U$5073 ( \13878_14177 , RIfc857d8_6541, \8953_9252 );
and \U$5074 ( \13879_14178 , RIee24dd8_4878, \8955_9254 );
and \U$5075 ( \13880_14179 , RIfc4ff70_5932, \8957_9256 );
and \U$5076 ( \13881_14180 , RIfc50240_5934, \8959_9258 );
and \U$5077 ( \13882_14181 , RIdee5ef8_1080, \8961_9260 );
and \U$5078 ( \13883_14182 , RIdee4170_1059, \8963_9262 );
and \U$5079 ( \13884_14183 , RIfe915c0_7998, \8965_9264 );
and \U$5080 ( \13885_14184 , RIdedff58_1012, \8967_9266 );
and \U$5081 ( \13886_14185 , RIfcd4810_7440, \8969_9268 );
and \U$5082 ( \13887_14186 , RIee22948_4852, \8971_9270 );
and \U$5083 ( \13888_14187 , RIfce1560_7586, \8973_9272 );
and \U$5084 ( \13889_14188 , RIee219d0_4841, \8975_9274 );
and \U$5085 ( \13890_14189 , RIdedac60_953, \8977_9276 );
and \U$5086 ( \13891_14190 , RIfe91728_7999, \8979_9278 );
and \U$5087 ( \13892_14191 , RIded64a8_902, \8981_9280 );
and \U$5088 ( \13893_14192 , RIfe91890_8000, \8983_9282 );
and \U$5089 ( \13894_14193 , RIded2128_854, \8985_9284 );
and \U$5090 ( \13895_14194 , RIdecf428_822, \8987_9286 );
and \U$5091 ( \13896_14195 , RIdecc728_790, \8989_9288 );
and \U$5092 ( \13897_14196 , RIdec9a28_758, \8991_9290 );
and \U$5093 ( \13898_14197 , RIdeb5f28_534, \8993_9292 );
and \U$5094 ( \13899_14198 , RIde9a430_342, \8995_9294 );
and \U$5095 ( \13900_14199 , RIe16fb30_2648, \8997_9296 );
and \U$5096 ( \13901_14200 , RIe15b928_2419, \8999_9298 );
and \U$5097 ( \13902_14201 , RIe145128_2163, \9001_9300 );
and \U$5098 ( \13903_14202 , RIdf39b20_2033, \9003_9302 );
and \U$5099 ( \13904_14203 , RIdf2e180_1901, \9005_9304 );
and \U$5100 ( \13905_14204 , RIdf1ea00_1725, \9007_9306 );
and \U$5101 ( \13906_14205 , RIdf020f8_1400, \9009_9308 );
and \U$5102 ( \13907_14206 , RIdee8bf8_1112, \9011_9310 );
and \U$5103 ( \13908_14207 , RIdedd960_985, \9013_9312 );
and \U$5104 ( \13909_14208 , RIde80378_215, \9015_9314 );
or \U$5105 ( \13910_14209 , \13846_14145 , \13847_14146 , \13848_14147 , \13849_14148 , \13850_14149 , \13851_14150 , \13852_14151 , \13853_14152 , \13854_14153 , \13855_14154 , \13856_14155 , \13857_14156 , \13858_14157 , \13859_14158 , \13860_14159 , \13861_14160 , \13862_14161 , \13863_14162 , \13864_14163 , \13865_14164 , \13866_14165 , \13867_14166 , \13868_14167 , \13869_14168 , \13870_14169 , \13871_14170 , \13872_14171 , \13873_14172 , \13874_14173 , \13875_14174 , \13876_14175 , \13877_14176 , \13878_14177 , \13879_14178 , \13880_14179 , \13881_14180 , \13882_14181 , \13883_14182 , \13884_14183 , \13885_14184 , \13886_14185 , \13887_14186 , \13888_14187 , \13889_14188 , \13890_14189 , \13891_14190 , \13892_14191 , \13893_14192 , \13894_14193 , \13895_14194 , \13896_14195 , \13897_14196 , \13898_14197 , \13899_14198 , \13900_14199 , \13901_14200 , \13902_14201 , \13903_14202 , \13904_14203 , \13905_14204 , \13906_14205 , \13907_14206 , \13908_14207 , \13909_14208 );
or \U$5106 ( \13911_14210 , \13845_14144 , \13910_14209 );
_DC \g2da3/U$1 ( \13912 , \13911_14210 , \9024_9323 );
buf \U$5107 ( \13913_14212 , \13912 );
and \U$5108 ( \13914_14213 , RIe19efc0_3186, \9034_9333 );
and \U$5109 ( \13915_14214 , RIe19c2c0_3154, \9036_9335 );
and \U$5110 ( \13916_14215 , RIf145d60_5254, \9038_9337 );
and \U$5111 ( \13917_14216 , RIe1995c0_3122, \9040_9339 );
and \U$5112 ( \13918_14217 , RIfc637a0_6154, \9042_9341 );
and \U$5113 ( \13919_14218 , RIe1968c0_3090, \9044_9343 );
and \U$5114 ( \13920_14219 , RIe193bc0_3058, \9046_9345 );
and \U$5115 ( \13921_14220 , RIe190ec0_3026, \9048_9347 );
and \U$5116 ( \13922_14221 , RIe18b4c0_2962, \9050_9349 );
and \U$5117 ( \13923_14222 , RIe1887c0_2930, \9052_9351 );
and \U$5118 ( \13924_14223 , RIfc62af8_6145, \9054_9353 );
and \U$5119 ( \13925_14224 , RIe185ac0_2898, \9056_9355 );
and \U$5120 ( \13926_14225 , RIfe8fc70_7980, \9058_9357 );
and \U$5121 ( \13927_14226 , RIe182dc0_2866, \9060_9359 );
and \U$5122 ( \13928_14227 , RIe1800c0_2834, \9062_9361 );
and \U$5123 ( \13929_14228 , RIe17d3c0_2802, \9064_9363 );
and \U$5124 ( \13930_14229 , RIfe90210_7984, \9066_9365 );
and \U$5125 ( \13931_14230 , RIfe8ff40_7982, \9068_9367 );
and \U$5126 ( \13932_14231 , RIfc72f20_6330, \9070_9369 );
and \U$5127 ( \13933_14232 , RIe176a48_2727, \9072_9371 );
and \U$5128 ( \13934_14233 , RIfcaf6a0_7018, \9074_9373 );
and \U$5129 ( \13935_14234 , RIfc61040_6126, \9076_9375 );
and \U$5130 ( \13936_14235 , RIf13e8a8_5171, \9078_9377 );
and \U$5131 ( \13937_14236 , RIfe900a8_7983, \9080_9379 );
and \U$5132 ( \13938_14237 , RIee3caf0_5149, \9082_9381 );
and \U$5133 ( \13939_14238 , RIee3b740_5135, \9084_9383 );
and \U$5134 ( \13940_14239 , RIee3a660_5123, \9086_9385 );
and \U$5135 ( \13941_14240 , RIe174e28_2707, \9088_9387 );
and \U$5136 ( \13942_14241 , RIf170768_5739, \9090_9389 );
and \U$5137 ( \13943_14242 , RIfc5fdf8_6113, \9092_9391 );
and \U$5138 ( \13944_14243 , RIf16eb48_5719, \9094_9393 );
and \U$5139 ( \13945_14244 , RIfcaaab0_6964, \9096_9395 );
and \U$5140 ( \13946_14245 , RIf16d1f8_5701, \9098_9397 );
and \U$5141 ( \13947_14246 , RIe225318_4713, \9100_9399 );
and \U$5142 ( \13948_14247 , RIf16c6b8_5693, \9102_9401 );
and \U$5143 ( \13949_14248 , RIe222618_4681, \9104_9403 );
and \U$5144 ( \13950_14249 , RIf16b5d8_5681, \9106_9405 );
and \U$5145 ( \13951_14250 , RIe21f918_4649, \9108_9407 );
and \U$5146 ( \13952_14251 , RIe219f18_4585, \9110_9409 );
and \U$5147 ( \13953_14252 , RIe217218_4553, \9112_9411 );
and \U$5148 ( \13954_14253 , RIfca62f8_6913, \9114_9413 );
and \U$5149 ( \13955_14254 , RIe214518_4521, \9116_9415 );
and \U$5150 ( \13956_14255 , RIfcc9578_7313, \9118_9417 );
and \U$5151 ( \13957_14256 , RIe211818_4489, \9120_9419 );
and \U$5152 ( \13958_14257 , RIfca5a88_6907, \9122_9421 );
and \U$5153 ( \13959_14258 , RIe20eb18_4457, \9124_9423 );
and \U$5154 ( \13960_14259 , RIe20be18_4425, \9126_9425 );
and \U$5155 ( \13961_14260 , RIe209118_4393, \9128_9427 );
and \U$5156 ( \13962_14261 , RIf167690_5636, \9130_9429 );
and \U$5157 ( \13963_14262 , RIf166718_5625, \9132_9431 );
and \U$5158 ( \13964_14263 , RIfe8f9a0_7978, \9134_9433 );
and \U$5159 ( \13965_14264 , RIfe8f838_7977, \9136_9435 );
and \U$5160 ( \13966_14265 , RIf165638_5613, \9138_9437 );
and \U$5161 ( \13967_14266 , RIf164990_5604, \9140_9439 );
and \U$5162 ( \13968_14267 , RIf1638b0_5592, \9142_9441 );
and \U$5163 ( \13969_14268 , RIf1627d0_5580, \9144_9443 );
and \U$5164 ( \13970_14269 , RIf161150_5564, \9146_9445 );
and \U$5165 ( \13971_14270 , RIf15f260_5542, \9148_9447 );
and \U$5166 ( \13972_14271 , RIe1fd778_4261, \9150_9449 );
and \U$5167 ( \13973_14272 , RIe1fc530_4248, \9152_9451 );
and \U$5168 ( \13974_14273 , RIf15d4d8_5521, \9154_9453 );
and \U$5169 ( \13975_14274 , RIf15c290_5508, \9156_9455 );
and \U$5170 ( \13976_14275 , RIfca20e0_6866, \9158_9457 );
and \U$5171 ( \13977_14276 , RIf159f68_5483, \9160_9459 );
or \U$5172 ( \13978_14277 , \13914_14213 , \13915_14214 , \13916_14215 , \13917_14216 , \13918_14217 , \13919_14218 , \13920_14219 , \13921_14220 , \13922_14221 , \13923_14222 , \13924_14223 , \13925_14224 , \13926_14225 , \13927_14226 , \13928_14227 , \13929_14228 , \13930_14229 , \13931_14230 , \13932_14231 , \13933_14232 , \13934_14233 , \13935_14234 , \13936_14235 , \13937_14236 , \13938_14237 , \13939_14238 , \13940_14239 , \13941_14240 , \13942_14241 , \13943_14242 , \13944_14243 , \13945_14244 , \13946_14245 , \13947_14246 , \13948_14247 , \13949_14248 , \13950_14249 , \13951_14250 , \13952_14251 , \13953_14252 , \13954_14253 , \13955_14254 , \13956_14255 , \13957_14256 , \13958_14257 , \13959_14258 , \13960_14259 , \13961_14260 , \13962_14261 , \13963_14262 , \13964_14263 , \13965_14264 , \13966_14265 , \13967_14266 , \13968_14267 , \13969_14268 , \13970_14269 , \13971_14270 , \13972_14271 , \13973_14272 , \13974_14273 , \13975_14274 , \13976_14275 , \13977_14276 );
and \U$5173 ( \13979_14278 , RIf159428_5475, \9163_9462 );
and \U$5174 ( \13980_14279 , RIf1581e0_5462, \9165_9464 );
and \U$5175 ( \13981_14280 , RIfc5ebb0_6100, \9167_9466 );
and \U$5176 ( \13982_14281 , RIfe8fdd8_7981, \9169_9468 );
and \U$5177 ( \13983_14282 , RIfc69e48_6227, \9171_9470 );
and \U$5178 ( \13984_14283 , RIfc5e8e0_6098, \9173_9472 );
and \U$5179 ( \13985_14284 , RIf154f40_5426, \9175_9474 );
and \U$5180 ( \13986_14285 , RIe1f6b30_4184, \9177_9476 );
and \U$5181 ( \13987_14286 , RIf153b90_5412, \9179_9478 );
and \U$5182 ( \13988_14287 , RIf1523a8_5395, \9181_9480 );
and \U$5183 ( \13989_14288 , RIfce88b0_7668, \9183_9482 );
and \U$5184 ( \13990_14289 , RIfe8fb08_7979, \9185_9484 );
and \U$5185 ( \13991_14290 , RIfcebe20_7706, \9187_9486 );
and \U$5186 ( \13992_14291 , RIfcb1158_7037, \9189_9488 );
and \U$5187 ( \13993_14292 , RIf14e730_5352, \9191_9490 );
and \U$5188 ( \13994_14293 , RIe1ef678_4101, \9193_9492 );
and \U$5189 ( \13995_14294 , RIe1ed080_4074, \9195_9494 );
and \U$5190 ( \13996_14295 , RIe1ea380_4042, \9197_9496 );
and \U$5191 ( \13997_14296 , RIe1e7680_4010, \9199_9498 );
and \U$5192 ( \13998_14297 , RIe1e4980_3978, \9201_9500 );
and \U$5193 ( \13999_14298 , RIe1e1c80_3946, \9203_9502 );
and \U$5194 ( \14000_14299 , RIe1def80_3914, \9205_9504 );
and \U$5195 ( \14001_14300 , RIe1dc280_3882, \9207_9506 );
and \U$5196 ( \14002_14301 , RIe1d9580_3850, \9209_9508 );
and \U$5197 ( \14003_14302 , RIe1d3b80_3786, \9211_9510 );
and \U$5198 ( \14004_14303 , RIe1d0e80_3754, \9213_9512 );
and \U$5199 ( \14005_14304 , RIe1ce180_3722, \9215_9514 );
and \U$5200 ( \14006_14305 , RIe1cb480_3690, \9217_9516 );
and \U$5201 ( \14007_14306 , RIe1c8780_3658, \9219_9518 );
and \U$5202 ( \14008_14307 , RIe1c5a80_3626, \9221_9520 );
and \U$5203 ( \14009_14308 , RIe1c2d80_3594, \9223_9522 );
and \U$5204 ( \14010_14309 , RIe1c0080_3562, \9225_9524 );
and \U$5205 ( \14011_14310 , RIfcc8ba0_7306, \9227_9526 );
and \U$5206 ( \14012_14311 , RIfc5d698_6085, \9229_9528 );
and \U$5207 ( \14013_14312 , RIfec35e8_8343, \9231_9530 );
and \U$5208 ( \14014_14313 , RIfeabd08_8271, \9233_9532 );
and \U$5209 ( \14015_14314 , RIfc5cf90_6080, \9235_9534 );
and \U$5210 ( \14016_14315 , RIfc5ce28_6079, \9237_9536 );
and \U$5211 ( \14017_14316 , RIfec31b0_8340, \9239_9538 );
and \U$5212 ( \14018_14317 , RIe1b4b18_3433, \9241_9540 );
and \U$5213 ( \14019_14318 , RIf149708_5295, \9243_9542 );
and \U$5214 ( \14020_14319 , RIf148358_5281, \9245_9544 );
and \U$5215 ( \14021_14320 , RIe1b3768_3419, \9247_9546 );
and \U$5216 ( \14022_14321 , RIfec3480_8342, \9249_9548 );
and \U$5217 ( \14023_14322 , RIfc483b0_5844, \9251_9550 );
and \U$5218 ( \14024_14323 , RIfc80be8_6487, \9253_9552 );
and \U$5219 ( \14025_14324 , RIe1ad4f8_3349, \9255_9554 );
and \U$5220 ( \14026_14325 , RIfec3318_8341, \9257_9556 );
and \U$5221 ( \14027_14326 , RIe1aa3c0_3314, \9259_9558 );
and \U$5222 ( \14028_14327 , RIe1a76c0_3282, \9261_9560 );
and \U$5223 ( \14029_14328 , RIe1a49c0_3250, \9263_9562 );
and \U$5224 ( \14030_14329 , RIe1a1cc0_3218, \9265_9564 );
and \U$5225 ( \14031_14330 , RIe18e1c0_2994, \9267_9566 );
and \U$5226 ( \14032_14331 , RIe17a6c0_2770, \9269_9568 );
and \U$5227 ( \14033_14332 , RIe228018_4745, \9271_9570 );
and \U$5228 ( \14034_14333 , RIe21cc18_4617, \9273_9572 );
and \U$5229 ( \14035_14334 , RIe206418_4361, \9275_9574 );
and \U$5230 ( \14036_14335 , RIe200478_4293, \9277_9576 );
and \U$5231 ( \14037_14336 , RIe1f9830_4216, \9279_9578 );
and \U$5232 ( \14038_14337 , RIe1f2378_4133, \9281_9580 );
and \U$5233 ( \14039_14338 , RIe1d6880_3818, \9283_9582 );
and \U$5234 ( \14040_14339 , RIe1bd380_3530, \9285_9584 );
and \U$5235 ( \14041_14340 , RIe1b01f8_3381, \9287_9586 );
and \U$5236 ( \14042_14341 , RIe172830_2680, \9289_9588 );
or \U$5237 ( \14043_14342 , \13979_14278 , \13980_14279 , \13981_14280 , \13982_14281 , \13983_14282 , \13984_14283 , \13985_14284 , \13986_14285 , \13987_14286 , \13988_14287 , \13989_14288 , \13990_14289 , \13991_14290 , \13992_14291 , \13993_14292 , \13994_14293 , \13995_14294 , \13996_14295 , \13997_14296 , \13998_14297 , \13999_14298 , \14000_14299 , \14001_14300 , \14002_14301 , \14003_14302 , \14004_14303 , \14005_14304 , \14006_14305 , \14007_14306 , \14008_14307 , \14009_14308 , \14010_14309 , \14011_14310 , \14012_14311 , \14013_14312 , \14014_14313 , \14015_14314 , \14016_14315 , \14017_14316 , \14018_14317 , \14019_14318 , \14020_14319 , \14021_14320 , \14022_14321 , \14023_14322 , \14024_14323 , \14025_14324 , \14026_14325 , \14027_14326 , \14028_14327 , \14029_14328 , \14030_14329 , \14031_14330 , \14032_14331 , \14033_14332 , \14034_14333 , \14035_14334 , \14036_14335 , \14037_14336 , \14038_14337 , \14039_14338 , \14040_14339 , \14041_14340 , \14042_14341 );
or \U$5238 ( \14044_14343 , \13978_14277 , \14043_14342 );
_DC \g3ed0/U$1 ( \14045 , \14044_14343 , \9298_9597 );
buf \U$5239 ( \14046_14345 , \14045 );
xor \U$5240 ( \14047_14346 , \13913_14212 , \14046_14345 );
and \U$5241 ( \14048_14347 , RIdec6bc0_725, \8760_9059 );
and \U$5242 ( \14049_14348 , RIdec3ec0_693, \8762_9061 );
and \U$5243 ( \14050_14349 , RIee20a58_4830, \8764_9063 );
and \U$5244 ( \14051_14350 , RIdec11c0_661, \8766_9065 );
and \U$5245 ( \14052_14351 , RIee1f978_4818, \8768_9067 );
and \U$5246 ( \14053_14352 , RIdebe4c0_629, \8770_9069 );
and \U$5247 ( \14054_14353 , RIdebb7c0_597, \8772_9071 );
and \U$5248 ( \14055_14354 , RIdeb8ac0_565, \8774_9073 );
and \U$5249 ( \14056_14355 , RIee1efa0_4811, \8776_9075 );
and \U$5250 ( \14057_14356 , RIdeb30c0_501, \8778_9077 );
and \U$5251 ( \14058_14357 , RIfcb04b0_7028, \8780_9079 );
and \U$5252 ( \14059_14358 , RIdeb03c0_469, \8782_9081 );
and \U$5253 ( \14060_14359 , RIfc5e4a8_6095, \8784_9083 );
and \U$5254 ( \14061_14360 , RIdead6c0_437, \8786_9085 );
and \U$5255 ( \14062_14361 , RIdea72e8_405, \8788_9087 );
and \U$5256 ( \14063_14362 , RIdea09e8_373, \8790_9089 );
and \U$5257 ( \14064_14363 , RIfcb2508_7051, \8792_9091 );
and \U$5258 ( \14065_14364 , RIfcd16d8_7405, \8794_9093 );
and \U$5259 ( \14066_14365 , RIfc5d800_6086, \8796_9095 );
and \U$5260 ( \14067_14366 , RIfc63d40_6158, \8798_9097 );
and \U$5261 ( \14068_14367 , RIde93b30_310, \8800_9099 );
and \U$5262 ( \14069_14368 , RIfea7820_8222, \8802_9101 );
and \U$5263 ( \14070_14369 , RIfea73e8_8219, \8804_9103 );
and \U$5264 ( \14071_14370 , RIde87998_251, \8806_9105 );
and \U$5265 ( \14072_14371 , RIde837f8_231, \8808_9107 );
and \U$5266 ( \14073_14372 , RIfc7bd28_6431, \8810_9109 );
and \U$5267 ( \14074_14373 , RIfcc7ef8_7297, \8812_9111 );
and \U$5268 ( \14075_14374 , RIfc7a108_6411, \8814_9113 );
and \U$5269 ( \14076_14375 , RIfc7a6a8_6415, \8816_9115 );
and \U$5270 ( \14077_14376 , RIe16ccc8_2615, \8818_9117 );
and \U$5271 ( \14078_14377 , RIe16a838_2589, \8820_9119 );
and \U$5272 ( \14079_14378 , RIe1691b8_2573, \8822_9121 );
and \U$5273 ( \14080_14379 , RIe166bc0_2546, \8824_9123 );
and \U$5274 ( \14081_14380 , RIe163ec0_2514, \8826_9125 );
and \U$5275 ( \14082_14381 , RIee38338_5098, \8828_9127 );
and \U$5276 ( \14083_14382 , RIe1611c0_2482, \8830_9129 );
and \U$5277 ( \14084_14383 , RIfc54b60_5986, \8832_9131 );
and \U$5278 ( \14085_14384 , RIe15e4c0_2450, \8834_9133 );
and \U$5279 ( \14086_14385 , RIe158ac0_2386, \8836_9135 );
and \U$5280 ( \14087_14386 , RIe155dc0_2354, \8838_9137 );
and \U$5281 ( \14088_14387 , RIee35a70_5069, \8840_9139 );
and \U$5282 ( \14089_14388 , RIe1530c0_2322, \8842_9141 );
and \U$5283 ( \14090_14389 , RIee357a0_5067, \8844_9143 );
and \U$5284 ( \14091_14390 , RIe1503c0_2290, \8846_9145 );
and \U$5285 ( \14092_14391 , RIfc9fdb8_6841, \8848_9147 );
and \U$5286 ( \14093_14392 , RIe14d6c0_2258, \8850_9149 );
and \U$5287 ( \14094_14393 , RIe14a9c0_2226, \8852_9151 );
and \U$5288 ( \14095_14394 , RIe147cc0_2194, \8854_9153 );
and \U$5289 ( \14096_14395 , RIee34af8_5058, \8856_9155 );
and \U$5290 ( \14097_14396 , RIee33a18_5046, \8858_9157 );
and \U$5291 ( \14098_14397 , RIee327d0_5033, \8860_9159 );
and \U$5292 ( \14099_14398 , RIfcbcf30_7172, \8862_9161 );
and \U$5293 ( \14100_14399 , RIe142428_2131, \8864_9163 );
and \U$5294 ( \14101_14400 , RIe140100_2106, \8866_9165 );
and \U$5295 ( \14102_14401 , RIfea7280_8218, \8868_9167 );
and \U$5296 ( \14103_14402 , RIdf3bb78_2056, \8870_9169 );
and \U$5297 ( \14104_14403 , RIfc731f0_6332, \8872_9171 );
and \U$5298 ( \14105_14404 , RIee30610_5009, \8874_9173 );
and \U$5299 ( \14106_14405 , RIfcbe010_7184, \8876_9175 );
and \U$5300 ( \14107_14406 , RIee2e450_4985, \8878_9177 );
and \U$5301 ( \14108_14407 , RIfec2ee0_8338, \8880_9179 );
and \U$5302 ( \14109_14408 , RIfec3048_8339, \8882_9181 );
and \U$5303 ( \14110_14409 , RIfec2c10_8336, \8884_9183 );
and \U$5304 ( \14111_14410 , RIfec2d78_8337, \8886_9185 );
or \U$5305 ( \14112_14411 , \14048_14347 , \14049_14348 , \14050_14349 , \14051_14350 , \14052_14351 , \14053_14352 , \14054_14353 , \14055_14354 , \14056_14355 , \14057_14356 , \14058_14357 , \14059_14358 , \14060_14359 , \14061_14360 , \14062_14361 , \14063_14362 , \14064_14363 , \14065_14364 , \14066_14365 , \14067_14366 , \14068_14367 , \14069_14368 , \14070_14369 , \14071_14370 , \14072_14371 , \14073_14372 , \14074_14373 , \14075_14374 , \14076_14375 , \14077_14376 , \14078_14377 , \14079_14378 , \14080_14379 , \14081_14380 , \14082_14381 , \14083_14382 , \14084_14383 , \14085_14384 , \14086_14385 , \14087_14386 , \14088_14387 , \14089_14388 , \14090_14389 , \14091_14390 , \14092_14391 , \14093_14392 , \14094_14393 , \14095_14394 , \14096_14395 , \14097_14396 , \14098_14397 , \14099_14398 , \14100_14399 , \14101_14400 , \14102_14401 , \14103_14402 , \14104_14403 , \14105_14404 , \14106_14405 , \14107_14406 , \14108_14407 , \14109_14408 , \14110_14409 , \14111_14410 );
and \U$5306 ( \14113_14412 , RIfcb46c8_7075, \8889_9188 );
and \U$5307 ( \14114_14413 , RIfcb4830_7076, \8891_9190 );
and \U$5308 ( \14115_14414 , RIee29860_4931, \8893_9192 );
and \U$5309 ( \14116_14415 , RIfcb88e0_7122, \8895_9194 );
and \U$5310 ( \14117_14416 , RIdf2b480_1869, \8897_9196 );
and \U$5311 ( \14118_14417 , RIdf29590_1847, \8899_9198 );
and \U$5312 ( \14119_14418 , RIdf27268_1822, \8901_9200 );
and \U$5313 ( \14120_14419 , RIdf25648_1802, \8903_9202 );
and \U$5314 ( \14121_14420 , RIfcc9de8_7319, \8905_9204 );
and \U$5315 ( \14122_14421 , RIfc53648_5971, \8907_9206 );
and \U$5316 ( \14123_14422 , RIdf23a28_1782, \8909_9208 );
and \U$5317 ( \14124_14423 , RIfc823d0_6504, \8911_9210 );
and \U$5318 ( \14125_14424 , RIdf223a8_1766, \8913_9212 );
and \U$5319 ( \14126_14425 , RIdf20d28_1750, \8915_9214 );
and \U$5320 ( \14127_14426 , RIdf1bd00_1693, \8917_9216 );
and \U$5321 ( \14128_14427 , RIdf1a7e8_1678, \8919_9218 );
and \U$5322 ( \14129_14428 , RIdf18790_1655, \8921_9220 );
and \U$5323 ( \14130_14429 , RIdf15a90_1623, \8923_9222 );
and \U$5324 ( \14131_14430 , RIdf12d90_1591, \8925_9224 );
and \U$5325 ( \14132_14431 , RIdf10090_1559, \8927_9226 );
and \U$5326 ( \14133_14432 , RIdf0d390_1527, \8929_9228 );
and \U$5327 ( \14134_14433 , RIdf0a690_1495, \8931_9230 );
and \U$5328 ( \14135_14434 , RIdf07990_1463, \8933_9232 );
and \U$5329 ( \14136_14435 , RIdf04c90_1431, \8935_9234 );
and \U$5330 ( \14137_14436 , RIdeff290_1367, \8937_9236 );
and \U$5331 ( \14138_14437 , RIdefc590_1335, \8939_9238 );
and \U$5332 ( \14139_14438 , RIdef9890_1303, \8941_9240 );
and \U$5333 ( \14140_14439 , RIdef6b90_1271, \8943_9242 );
and \U$5334 ( \14141_14440 , RIdef3e90_1239, \8945_9244 );
and \U$5335 ( \14142_14441 , RIdef1190_1207, \8947_9246 );
and \U$5336 ( \14143_14442 , RIdeee490_1175, \8949_9248 );
and \U$5337 ( \14144_14443 , RIdeeb790_1143, \8951_9250 );
and \U$5338 ( \14145_14444 , RIee25be8_4888, \8953_9252 );
and \U$5339 ( \14146_14445 , RIfc6af28_6239, \8955_9254 );
and \U$5340 ( \14147_14446 , RIee23fc8_4868, \8957_9256 );
and \U$5341 ( \14148_14447 , RIfccf680_7382, \8959_9258 );
and \U$5342 ( \14149_14448 , RIdee5d90_1079, \8961_9260 );
and \U$5343 ( \14150_14449 , RIdee4008_1058, \8963_9262 );
and \U$5344 ( \14151_14450 , RIdee1ce0_1033, \8965_9264 );
and \U$5345 ( \14152_14451 , RIdedfdf0_1011, \8967_9266 );
and \U$5346 ( \14153_14452 , RIfc6b090_6240, \8969_9268 );
and \U$5347 ( \14154_14453 , RIfc534e0_5970, \8971_9270 );
and \U$5348 ( \14155_14454 , RIfca5920_6906, \8973_9272 );
and \U$5349 ( \14156_14455 , RIfc66770_6188, \8975_9274 );
and \U$5350 ( \14157_14456 , RIfe8f6d0_7976, \8977_9276 );
and \U$5351 ( \14158_14457 , RIded87d0_927, \8979_9278 );
and \U$5352 ( \14159_14458 , RIfe8f568_7975, \8981_9280 );
and \U$5353 ( \14160_14459 , RIded42e8_878, \8983_9282 );
and \U$5354 ( \14161_14460 , RIded1fc0_853, \8985_9284 );
and \U$5355 ( \14162_14461 , RIdecf2c0_821, \8987_9286 );
and \U$5356 ( \14163_14462 , RIdecc5c0_789, \8989_9288 );
and \U$5357 ( \14164_14463 , RIdec98c0_757, \8991_9290 );
and \U$5358 ( \14165_14464 , RIdeb5dc0_533, \8993_9292 );
and \U$5359 ( \14166_14465 , RIde9a0e8_341, \8995_9294 );
and \U$5360 ( \14167_14466 , RIe16f9c8_2647, \8997_9296 );
and \U$5361 ( \14168_14467 , RIe15b7c0_2418, \8999_9298 );
and \U$5362 ( \14169_14468 , RIe144fc0_2162, \9001_9300 );
and \U$5363 ( \14170_14469 , RIdf399b8_2032, \9003_9302 );
and \U$5364 ( \14171_14470 , RIdf2e018_1900, \9005_9304 );
and \U$5365 ( \14172_14471 , RIdf1e898_1724, \9007_9306 );
and \U$5366 ( \14173_14472 , RIdf01f90_1399, \9009_9308 );
and \U$5367 ( \14174_14473 , RIdee8a90_1111, \9011_9310 );
and \U$5368 ( \14175_14474 , RIdedd7f8_984, \9013_9312 );
and \U$5369 ( \14176_14475 , RIde80030_214, \9015_9314 );
or \U$5370 ( \14177_14476 , \14113_14412 , \14114_14413 , \14115_14414 , \14116_14415 , \14117_14416 , \14118_14417 , \14119_14418 , \14120_14419 , \14121_14420 , \14122_14421 , \14123_14422 , \14124_14423 , \14125_14424 , \14126_14425 , \14127_14426 , \14128_14427 , \14129_14428 , \14130_14429 , \14131_14430 , \14132_14431 , \14133_14432 , \14134_14433 , \14135_14434 , \14136_14435 , \14137_14436 , \14138_14437 , \14139_14438 , \14140_14439 , \14141_14440 , \14142_14441 , \14143_14442 , \14144_14443 , \14145_14444 , \14146_14445 , \14147_14446 , \14148_14447 , \14149_14448 , \14150_14449 , \14151_14450 , \14152_14451 , \14153_14452 , \14154_14453 , \14155_14454 , \14156_14455 , \14157_14456 , \14158_14457 , \14159_14458 , \14160_14459 , \14161_14460 , \14162_14461 , \14163_14462 , \14164_14463 , \14165_14464 , \14166_14465 , \14167_14466 , \14168_14467 , \14169_14468 , \14170_14469 , \14171_14470 , \14172_14471 , \14173_14472 , \14174_14473 , \14175_14474 , \14176_14475 );
or \U$5371 ( \14178_14477 , \14112_14411 , \14177_14476 );
_DC \g2e28/U$1 ( \14179 , \14178_14477 , \9024_9323 );
buf \U$5372 ( \14180_14479 , \14179 );
and \U$5373 ( \14181_14480 , RIe19ee58_3185, \9034_9333 );
and \U$5374 ( \14182_14481 , RIe19c158_3153, \9036_9335 );
and \U$5375 ( \14183_14482 , RIf145bf8_5253, \9038_9337 );
and \U$5376 ( \14184_14483 , RIe199458_3121, \9040_9339 );
and \U$5377 ( \14185_14484 , RIfe8f298_7973, \9042_9341 );
and \U$5378 ( \14186_14485 , RIe196758_3089, \9044_9343 );
and \U$5379 ( \14187_14486 , RIe193a58_3057, \9046_9345 );
and \U$5380 ( \14188_14487 , RIe190d58_3025, \9048_9347 );
and \U$5381 ( \14189_14488 , RIe18b358_2961, \9050_9349 );
and \U$5382 ( \14190_14489 , RIe188658_2929, \9052_9351 );
and \U$5383 ( \14191_14490 , RIfe8f130_7972, \9054_9353 );
and \U$5384 ( \14192_14491 , RIe185958_2897, \9056_9355 );
and \U$5385 ( \14193_14492 , RIfc9f278_6833, \9058_9357 );
and \U$5386 ( \14194_14493 , RIe182c58_2865, \9060_9359 );
and \U$5387 ( \14195_14494 , RIe17ff58_2833, \9062_9361 );
and \U$5388 ( \14196_14495 , RIe17d258_2801, \9064_9363 );
and \U$5389 ( \14197_14496 , RIf1427f0_5216, \9066_9365 );
and \U$5390 ( \14198_14497 , RIfe8efc8_7971, \9068_9367 );
and \U$5391 ( \14199_14498 , RIe1779c0_2738, \9070_9369 );
and \U$5392 ( \14200_14499 , RIe1768e0_2726, \9072_9371 );
and \U$5393 ( \14201_14500 , RIfc81e30_6500, \9074_9373 );
and \U$5394 ( \14202_14501 , RIfc9ff20_6842, \9076_9375 );
and \U$5395 ( \14203_14502 , RIfca0088_6843, \9078_9377 );
and \U$5396 ( \14204_14503 , RIfc81b60_6498, \9080_9379 );
and \U$5397 ( \14205_14504 , RIfce5778_7633, \9082_9381 );
and \U$5398 ( \14206_14505 , RIfce08b8_7577, \9084_9383 );
and \U$5399 ( \14207_14506 , RIfc815c0_6494, \9086_9385 );
and \U$5400 ( \14208_14507 , RIe174cc0_2706, \9088_9387 );
and \U$5401 ( \14209_14508 , RIfca04c0_6846, \9090_9389 );
and \U$5402 ( \14210_14509 , RIfc53eb8_5977, \9092_9391 );
and \U$5403 ( \14211_14510 , RIfcc65a8_7279, \9094_9393 );
and \U$5404 ( \14212_14511 , RIfc80d50_6488, \9096_9395 );
and \U$5405 ( \14213_14512 , RIfc804e0_6482, \9098_9397 );
and \U$5406 ( \14214_14513 , RIe2251b0_4712, \9100_9399 );
and \U$5407 ( \14215_14514 , RIfc80378_6481, \9102_9401 );
and \U$5408 ( \14216_14515 , RIe2224b0_4680, \9104_9403 );
and \U$5409 ( \14217_14516 , RIfcb5910_7088, \9106_9405 );
and \U$5410 ( \14218_14517 , RIe21f7b0_4648, \9108_9407 );
and \U$5411 ( \14219_14518 , RIe219db0_4584, \9110_9409 );
and \U$5412 ( \14220_14519 , RIe2170b0_4552, \9112_9411 );
and \U$5413 ( \14221_14520 , RIfca01f0_6844, \9114_9413 );
and \U$5414 ( \14222_14521 , RIe2143b0_4520, \9116_9415 );
and \U$5415 ( \14223_14522 , RIfc82c40_6510, \9118_9417 );
and \U$5416 ( \14224_14523 , RIe2116b0_4488, \9120_9419 );
and \U$5417 ( \14225_14524 , RIfc7f6d0_6472, \9122_9421 );
and \U$5418 ( \14226_14525 , RIe20e9b0_4456, \9124_9423 );
and \U$5419 ( \14227_14526 , RIe20bcb0_4424, \9126_9425 );
and \U$5420 ( \14228_14527 , RIe208fb0_4392, \9128_9427 );
and \U$5421 ( \14229_14528 , RIf167528_5635, \9130_9429 );
and \U$5422 ( \14230_14529 , RIf1665b0_5624, \9132_9431 );
and \U$5423 ( \14231_14530 , RIe203718_4329, \9134_9433 );
and \U$5424 ( \14232_14531 , RIe201c60_4310, \9136_9435 );
and \U$5425 ( \14233_14532 , RIfc9da90_6816, \9138_9437 );
and \U$5426 ( \14234_14533 , RIfcc5360_7266, \9140_9439 );
and \U$5427 ( \14235_14534 , RIf163748_5591, \9142_9441 );
and \U$5428 ( \14236_14535 , RIf162668_5579, \9144_9443 );
and \U$5429 ( \14237_14536 , RIfc7e320_6458, \9146_9445 );
and \U$5430 ( \14238_14537 , RIfc87998_6565, \9148_9447 );
and \U$5431 ( \14239_14538 , RIe1fd610_4260, \9150_9449 );
and \U$5432 ( \14240_14539 , RIe1fc3c8_4247, \9152_9451 );
and \U$5433 ( \14241_14540 , RIf15d370_5520, \9154_9453 );
and \U$5434 ( \14242_14541 , RIf15c128_5507, \9156_9455 );
and \U$5435 ( \14243_14542 , RIfcc5d38_7273, \9158_9457 );
and \U$5436 ( \14244_14543 , RIfce7d70_7660, \9160_9459 );
or \U$5437 ( \14245_14544 , \14181_14480 , \14182_14481 , \14183_14482 , \14184_14483 , \14185_14484 , \14186_14485 , \14187_14486 , \14188_14487 , \14189_14488 , \14190_14489 , \14191_14490 , \14192_14491 , \14193_14492 , \14194_14493 , \14195_14494 , \14196_14495 , \14197_14496 , \14198_14497 , \14199_14498 , \14200_14499 , \14201_14500 , \14202_14501 , \14203_14502 , \14204_14503 , \14205_14504 , \14206_14505 , \14207_14506 , \14208_14507 , \14209_14508 , \14210_14509 , \14211_14510 , \14212_14511 , \14213_14512 , \14214_14513 , \14215_14514 , \14216_14515 , \14217_14516 , \14218_14517 , \14219_14518 , \14220_14519 , \14221_14520 , \14222_14521 , \14223_14522 , \14224_14523 , \14225_14524 , \14226_14525 , \14227_14526 , \14228_14527 , \14229_14528 , \14230_14529 , \14231_14530 , \14232_14531 , \14233_14532 , \14234_14533 , \14235_14534 , \14236_14535 , \14237_14536 , \14238_14537 , \14239_14538 , \14240_14539 , \14241_14540 , \14242_14541 , \14243_14542 , \14244_14543 );
and \U$5438 ( \14246_14545 , RIfc4bd58_5885, \9163_9462 );
and \U$5439 ( \14247_14546 , RIfc55c40_5998, \9165_9464 );
and \U$5440 ( \14248_14547 , RIfca2ab8_6873, \9167_9466 );
and \U$5441 ( \14249_14548 , RIe1fb450_4236, \9169_9468 );
and \U$5442 ( \14250_14549 , RIf156890_5444, \9171_9470 );
and \U$5443 ( \14251_14550 , RIfcd5ff8_7457, \9173_9472 );
and \U$5444 ( \14252_14551 , RIf154dd8_5425, \9175_9474 );
and \U$5445 ( \14253_14552 , RIfec2aa8_8335, \9177_9476 );
and \U$5446 ( \14254_14553 , RIfcb4b00_7078, \9179_9478 );
and \U$5447 ( \14255_14554 , RIfcd9400_7494, \9181_9480 );
and \U$5448 ( \14256_14555 , RIf151160_5382, \9183_9482 );
and \U$5449 ( \14257_14556 , RIe1f4808_4159, \9185_9484 );
and \U$5450 ( \14258_14557 , RIfc44738_5801, \9187_9486 );
and \U$5451 ( \14259_14558 , RIfc90908_6667, \9189_9488 );
and \U$5452 ( \14260_14559 , RIf14e5c8_5351, \9191_9490 );
and \U$5453 ( \14261_14560 , RIe1ef510_4100, \9193_9492 );
and \U$5454 ( \14262_14561 , RIe1ecf18_4073, \9195_9494 );
and \U$5455 ( \14263_14562 , RIe1ea218_4041, \9197_9496 );
and \U$5456 ( \14264_14563 , RIe1e7518_4009, \9199_9498 );
and \U$5457 ( \14265_14564 , RIe1e4818_3977, \9201_9500 );
and \U$5458 ( \14266_14565 , RIe1e1b18_3945, \9203_9502 );
and \U$5459 ( \14267_14566 , RIe1dee18_3913, \9205_9504 );
and \U$5460 ( \14268_14567 , RIe1dc118_3881, \9207_9506 );
and \U$5461 ( \14269_14568 , RIe1d9418_3849, \9209_9508 );
and \U$5462 ( \14270_14569 , RIe1d3a18_3785, \9211_9510 );
and \U$5463 ( \14271_14570 , RIe1d0d18_3753, \9213_9512 );
and \U$5464 ( \14272_14571 , RIe1ce018_3721, \9215_9514 );
and \U$5465 ( \14273_14572 , RIe1cb318_3689, \9217_9516 );
and \U$5466 ( \14274_14573 , RIe1c8618_3657, \9219_9518 );
and \U$5467 ( \14275_14574 , RIe1c5918_3625, \9221_9520 );
and \U$5468 ( \14276_14575 , RIe1c2c18_3593, \9223_9522 );
and \U$5469 ( \14277_14576 , RIe1bff18_3561, \9225_9524 );
and \U$5470 ( \14278_14577 , RIf14d218_5337, \9227_9526 );
and \U$5471 ( \14279_14578 , RIfe8ee60_7970, \9229_9528 );
and \U$5472 ( \14280_14579 , RIfea8090_8228, \9231_9530 );
and \U$5473 ( \14281_14580 , RIe1b84c0_3474, \9233_9532 );
and \U$5474 ( \14282_14581 , RIf14aab8_5309, \9235_9534 );
and \U$5475 ( \14283_14582 , RIfc6c170_6252, \9237_9536 );
and \U$5476 ( \14284_14583 , RIe1b6468_3451, \9239_9538 );
and \U$5477 ( \14285_14584 , RIe1b49b0_3432, \9241_9540 );
and \U$5478 ( \14286_14585 , RIfcafad8_7021, \9243_9542 );
and \U$5479 ( \14287_14586 , RIfcaa948_6963, \9245_9544 );
and \U$5480 ( \14288_14587 , RIfe8ecf8_7969, \9247_9546 );
and \U$5481 ( \14289_14588 , RIfe8f400_7974, \9249_9548 );
and \U$5482 ( \14290_14589 , RIfc67f58_6205, \9251_9550 );
and \U$5483 ( \14291_14590 , RIfca8ff8_6945, \9253_9552 );
and \U$5484 ( \14292_14591 , RIfe8eb90_7968, \9255_9554 );
and \U$5485 ( \14293_14592 , RIe1abe78_3333, \9257_9556 );
and \U$5486 ( \14294_14593 , RIe1aa258_3313, \9259_9558 );
and \U$5487 ( \14295_14594 , RIe1a7558_3281, \9261_9560 );
and \U$5488 ( \14296_14595 , RIe1a4858_3249, \9263_9562 );
and \U$5489 ( \14297_14596 , RIe1a1b58_3217, \9265_9564 );
and \U$5490 ( \14298_14597 , RIe18e058_2993, \9267_9566 );
and \U$5491 ( \14299_14598 , RIe17a558_2769, \9269_9568 );
and \U$5492 ( \14300_14599 , RIe227eb0_4744, \9271_9570 );
and \U$5493 ( \14301_14600 , RIe21cab0_4616, \9273_9572 );
and \U$5494 ( \14302_14601 , RIe2062b0_4360, \9275_9574 );
and \U$5495 ( \14303_14602 , RIe200310_4292, \9277_9576 );
and \U$5496 ( \14304_14603 , RIe1f96c8_4215, \9279_9578 );
and \U$5497 ( \14305_14604 , RIe1f2210_4132, \9281_9580 );
and \U$5498 ( \14306_14605 , RIe1d6718_3817, \9283_9582 );
and \U$5499 ( \14307_14606 , RIe1bd218_3529, \9285_9584 );
and \U$5500 ( \14308_14607 , RIe1b0090_3380, \9287_9586 );
and \U$5501 ( \14309_14608 , RIe1726c8_2679, \9289_9588 );
or \U$5502 ( \14310_14609 , \14246_14545 , \14247_14546 , \14248_14547 , \14249_14548 , \14250_14549 , \14251_14550 , \14252_14551 , \14253_14552 , \14254_14553 , \14255_14554 , \14256_14555 , \14257_14556 , \14258_14557 , \14259_14558 , \14260_14559 , \14261_14560 , \14262_14561 , \14263_14562 , \14264_14563 , \14265_14564 , \14266_14565 , \14267_14566 , \14268_14567 , \14269_14568 , \14270_14569 , \14271_14570 , \14272_14571 , \14273_14572 , \14274_14573 , \14275_14574 , \14276_14575 , \14277_14576 , \14278_14577 , \14279_14578 , \14280_14579 , \14281_14580 , \14282_14581 , \14283_14582 , \14284_14583 , \14285_14584 , \14286_14585 , \14287_14586 , \14288_14587 , \14289_14588 , \14290_14589 , \14291_14590 , \14292_14591 , \14293_14592 , \14294_14593 , \14295_14594 , \14296_14595 , \14297_14596 , \14298_14597 , \14299_14598 , \14300_14599 , \14301_14600 , \14302_14601 , \14303_14602 , \14304_14603 , \14305_14604 , \14306_14605 , \14307_14606 , \14308_14607 , \14309_14608 );
or \U$5503 ( \14311_14610 , \14245_14544 , \14310_14609 );
_DC \g3f55/U$1 ( \14312 , \14311_14610 , \9298_9597 );
buf \U$5504 ( \14313_14612 , \14312 );
and \U$5505 ( \14314_14613 , \14180_14479 , \14313_14612 );
and \U$5506 ( \14315_14614 , \12652_12951 , \12785_13084 );
and \U$5507 ( \14316_14615 , \12785_13084 , \13060_13359 );
and \U$5508 ( \14317_14616 , \12652_12951 , \13060_13359 );
or \U$5509 ( \14318_14617 , \14315_14614 , \14316_14615 , \14317_14616 );
and \U$5510 ( \14319_14618 , \14313_14612 , \14318_14617 );
and \U$5511 ( \14320_14619 , \14180_14479 , \14318_14617 );
or \U$5512 ( \14321_14620 , \14314_14613 , \14319_14618 , \14320_14619 );
xor \U$5513 ( \14322_14621 , \14047_14346 , \14321_14620 );
buf g443c_GF_PartitionCandidate( \14323_14622_nG443c , \14322_14621 );
xor \U$5514 ( \14324_14623 , \14180_14479 , \14313_14612 );
xor \U$5515 ( \14325_14624 , \14324_14623 , \14318_14617 );
buf g443f_GF_PartitionCandidate( \14326_14625_nG443f , \14325_14624 );
nand \U$5516 ( \14327_14626 , \14326_14625_nG443f , \13062_13361_nG4442 );
and \U$5517 ( \14328_14627 , \14323_14622_nG443c , \14327_14626 );
xor \U$5518 ( \14329_14628 , \14326_14625_nG443f , \13062_13361_nG4442 );
and \U$5523 ( \14330_14632 , \14329_14628 , \10392_10694_nG9c0e );
or \U$5524 ( \14331_14633 , 1'b0 , \14330_14632 );
xor \U$5525 ( \14332_14634 , \14328_14627 , \14331_14633 );
xor \U$5526 ( \14333_14635 , \14328_14627 , \14332_14634 );
buf \U$5527 ( \14334_14636 , \14333_14635 );
buf \U$5528 ( \14335_14637 , \14334_14636 );
and \U$5529 ( \14336_14638 , \13780_14079 , \14335_14637 );
and \U$5530 ( \14337_14639 , \13419_13721 , \13424_13726 );
and \U$5531 ( \14338_14640 , \13419_13721 , \13778_14077 );
and \U$5532 ( \14339_14641 , \13424_13726 , \13778_14077 );
or \U$5533 ( \14340_14642 , \14337_14639 , \14338_14640 , \14339_14641 );
buf \U$5534 ( \14341_14643 , \14340_14642 );
and \U$5535 ( \14342_14644 , \13428_13730 , \13437_13736 );
buf \U$5536 ( \14343_14645 , \14342_14644 );
and \U$5537 ( \14344_14646 , \13431_13370 , \10693_10995_nG9c0b );
and \U$5538 ( \14345_14647 , \13068_13367 , \10981_11283_nG9c08 );
or \U$5539 ( \14346_14648 , \14344_14646 , \14345_14647 );
xor \U$5540 ( \14347_14649 , \13067_13366 , \14346_14648 );
buf \U$5541 ( \14348_14650 , \14347_14649 );
buf \U$5543 ( \14349_14651 , \14348_14650 );
xor \U$5544 ( \14350_14652 , \14343_14645 , \14349_14651 );
buf \U$5545 ( \14351_14653 , \14350_14652 );
and \U$5546 ( \14352_14654 , \12183_12157 , \11299_11598_nG9c05 );
and \U$5547 ( \14353_14655 , \11855_12154 , \12168_12470_nG9c02 );
or \U$5548 ( \14354_14656 , \14352_14654 , \14353_14655 );
xor \U$5549 ( \14355_14657 , \11854_12153 , \14354_14656 );
buf \U$5550 ( \14356_14658 , \14355_14657 );
buf \U$5552 ( \14357_14659 , \14356_14658 );
xor \U$5553 ( \14358_14660 , \14351_14653 , \14357_14659 );
and \U$5554 ( \14359_14661 , \10996_10421 , \12502_12801_nG9bff );
and \U$5555 ( \14360_14662 , \10119_10418 , \13403_13705_nG9bfc );
or \U$5556 ( \14361_14663 , \14359_14661 , \14360_14662 );
xor \U$5557 ( \14362_14664 , \10118_10417 , \14361_14663 );
buf \U$5558 ( \14363_14665 , \14362_14664 );
buf \U$5560 ( \14364_14666 , \14363_14665 );
xor \U$5561 ( \14365_14667 , \14358_14660 , \14364_14666 );
buf \U$5562 ( \14366_14668 , \14365_14667 );
and \U$5563 ( \14367_14669 , \13439_13738 , \13445_13744 );
and \U$5564 ( \14368_14670 , \13439_13738 , \13452_13751 );
and \U$5565 ( \14369_14671 , \13445_13744 , \13452_13751 );
or \U$5566 ( \14370_14672 , \14367_14669 , \14368_14670 , \14369_14671 );
buf \U$5567 ( \14371_14673 , \14370_14672 );
xor \U$5568 ( \14372_14674 , \14366_14668 , \14371_14673 );
and \U$5569 ( \14373_14675 , \10411_10707 , \13771_14070_nG9bf9 );
and \U$5570 ( \14374_14676 , \13738_14037 , \13742_14041 );
and \U$5571 ( \14375_14677 , \13742_14041 , \13760_14059 );
and \U$5572 ( \14376_14678 , \13738_14037 , \13760_14059 );
or \U$5573 ( \14377_14679 , \14374_14676 , \14375_14677 , \14376_14678 );
and \U$5574 ( \14378_14680 , \13747_14046 , \13751_14050 );
and \U$5575 ( \14379_14681 , \13751_14050 , \13759_14058 );
and \U$5576 ( \14380_14682 , \13747_14046 , \13759_14058 );
or \U$5577 ( \14381_14683 , \14378_14680 , \14379_14681 , \14380_14682 );
and \U$5578 ( \14382_14684 , \13725_14024 , \10681_10983 );
and \U$5579 ( \14383_14685 , RIdec6bc0_725, \9034_9333 );
and \U$5580 ( \14384_14686 , RIdec3ec0_693, \9036_9335 );
and \U$5581 ( \14385_14687 , RIee20a58_4830, \9038_9337 );
and \U$5582 ( \14386_14688 , RIdec11c0_661, \9040_9339 );
and \U$5583 ( \14387_14689 , RIee1f978_4818, \9042_9341 );
and \U$5584 ( \14388_14690 , RIdebe4c0_629, \9044_9343 );
and \U$5585 ( \14389_14691 , RIdebb7c0_597, \9046_9345 );
and \U$5586 ( \14390_14692 , RIdeb8ac0_565, \9048_9347 );
and \U$5587 ( \14391_14693 , RIee1efa0_4811, \9050_9349 );
and \U$5588 ( \14392_14694 , RIdeb30c0_501, \9052_9351 );
and \U$5589 ( \14393_14695 , RIfcb04b0_7028, \9054_9353 );
and \U$5590 ( \14394_14696 , RIdeb03c0_469, \9056_9355 );
and \U$5591 ( \14395_14697 , RIfc5e4a8_6095, \9058_9357 );
and \U$5592 ( \14396_14698 , RIdead6c0_437, \9060_9359 );
and \U$5593 ( \14397_14699 , RIdea72e8_405, \9062_9361 );
and \U$5594 ( \14398_14700 , RIdea09e8_373, \9064_9363 );
and \U$5595 ( \14399_14701 , RIfcb2508_7051, \9066_9365 );
and \U$5596 ( \14400_14702 , RIfcd16d8_7405, \9068_9367 );
and \U$5597 ( \14401_14703 , RIfc5d800_6086, \9070_9369 );
and \U$5598 ( \14402_14704 , RIfc63d40_6158, \9072_9371 );
and \U$5599 ( \14403_14705 , RIde93b30_310, \9074_9373 );
and \U$5600 ( \14404_14706 , RIfea7820_8222, \9076_9375 );
and \U$5601 ( \14405_14707 , RIfea73e8_8219, \9078_9377 );
and \U$5602 ( \14406_14708 , RIde87998_251, \9080_9379 );
and \U$5603 ( \14407_14709 , RIde837f8_231, \9082_9381 );
and \U$5604 ( \14408_14710 , RIfc7bd28_6431, \9084_9383 );
and \U$5605 ( \14409_14711 , RIfcc7ef8_7297, \9086_9385 );
and \U$5606 ( \14410_14712 , RIfc7a108_6411, \9088_9387 );
and \U$5607 ( \14411_14713 , RIfc7a6a8_6415, \9090_9389 );
and \U$5608 ( \14412_14714 , RIe16ccc8_2615, \9092_9391 );
and \U$5609 ( \14413_14715 , RIe16a838_2589, \9094_9393 );
and \U$5610 ( \14414_14716 , RIe1691b8_2573, \9096_9395 );
and \U$5611 ( \14415_14717 , RIe166bc0_2546, \9098_9397 );
and \U$5612 ( \14416_14718 , RIe163ec0_2514, \9100_9399 );
and \U$5613 ( \14417_14719 , RIee38338_5098, \9102_9401 );
and \U$5614 ( \14418_14720 , RIe1611c0_2482, \9104_9403 );
and \U$5615 ( \14419_14721 , RIfc54b60_5986, \9106_9405 );
and \U$5616 ( \14420_14722 , RIe15e4c0_2450, \9108_9407 );
and \U$5617 ( \14421_14723 , RIe158ac0_2386, \9110_9409 );
and \U$5618 ( \14422_14724 , RIe155dc0_2354, \9112_9411 );
and \U$5619 ( \14423_14725 , RIee35a70_5069, \9114_9413 );
and \U$5620 ( \14424_14726 , RIe1530c0_2322, \9116_9415 );
and \U$5621 ( \14425_14727 , RIee357a0_5067, \9118_9417 );
and \U$5622 ( \14426_14728 , RIe1503c0_2290, \9120_9419 );
and \U$5623 ( \14427_14729 , RIfc9fdb8_6841, \9122_9421 );
and \U$5624 ( \14428_14730 , RIe14d6c0_2258, \9124_9423 );
and \U$5625 ( \14429_14731 , RIe14a9c0_2226, \9126_9425 );
and \U$5626 ( \14430_14732 , RIe147cc0_2194, \9128_9427 );
and \U$5627 ( \14431_14733 , RIee34af8_5058, \9130_9429 );
and \U$5628 ( \14432_14734 , RIee33a18_5046, \9132_9431 );
and \U$5629 ( \14433_14735 , RIee327d0_5033, \9134_9433 );
and \U$5630 ( \14434_14736 , RIfcbcf30_7172, \9136_9435 );
and \U$5631 ( \14435_14737 , RIe142428_2131, \9138_9437 );
and \U$5632 ( \14436_14738 , RIe140100_2106, \9140_9439 );
and \U$5633 ( \14437_14739 , RIfea7280_8218, \9142_9441 );
and \U$5634 ( \14438_14740 , RIdf3bb78_2056, \9144_9443 );
and \U$5635 ( \14439_14741 , RIfc731f0_6332, \9146_9445 );
and \U$5636 ( \14440_14742 , RIee30610_5009, \9148_9447 );
and \U$5637 ( \14441_14743 , RIfcbe010_7184, \9150_9449 );
and \U$5638 ( \14442_14744 , RIee2e450_4985, \9152_9451 );
and \U$5639 ( \14443_14745 , RIfec2ee0_8338, \9154_9453 );
and \U$5640 ( \14444_14746 , RIfec3048_8339, \9156_9455 );
and \U$5641 ( \14445_14747 , RIfec2c10_8336, \9158_9457 );
and \U$5642 ( \14446_14748 , RIfec2d78_8337, \9160_9459 );
or \U$5643 ( \14447_14749 , \14383_14685 , \14384_14686 , \14385_14687 , \14386_14688 , \14387_14689 , \14388_14690 , \14389_14691 , \14390_14692 , \14391_14693 , \14392_14694 , \14393_14695 , \14394_14696 , \14395_14697 , \14396_14698 , \14397_14699 , \14398_14700 , \14399_14701 , \14400_14702 , \14401_14703 , \14402_14704 , \14403_14705 , \14404_14706 , \14405_14707 , \14406_14708 , \14407_14709 , \14408_14710 , \14409_14711 , \14410_14712 , \14411_14713 , \14412_14714 , \14413_14715 , \14414_14716 , \14415_14717 , \14416_14718 , \14417_14719 , \14418_14720 , \14419_14721 , \14420_14722 , \14421_14723 , \14422_14724 , \14423_14725 , \14424_14726 , \14425_14727 , \14426_14728 , \14427_14729 , \14428_14730 , \14429_14731 , \14430_14732 , \14431_14733 , \14432_14734 , \14433_14735 , \14434_14736 , \14435_14737 , \14436_14738 , \14437_14739 , \14438_14740 , \14439_14741 , \14440_14742 , \14441_14743 , \14442_14744 , \14443_14745 , \14444_14746 , \14445_14747 , \14446_14748 );
and \U$5644 ( \14448_14750 , RIfcb46c8_7075, \9163_9462 );
and \U$5645 ( \14449_14751 , RIfcb4830_7076, \9165_9464 );
and \U$5646 ( \14450_14752 , RIee29860_4931, \9167_9466 );
and \U$5647 ( \14451_14753 , RIfcb88e0_7122, \9169_9468 );
and \U$5648 ( \14452_14754 , RIdf2b480_1869, \9171_9470 );
and \U$5649 ( \14453_14755 , RIdf29590_1847, \9173_9472 );
and \U$5650 ( \14454_14756 , RIdf27268_1822, \9175_9474 );
and \U$5651 ( \14455_14757 , RIdf25648_1802, \9177_9476 );
and \U$5652 ( \14456_14758 , RIfcc9de8_7319, \9179_9478 );
and \U$5653 ( \14457_14759 , RIfc53648_5971, \9181_9480 );
and \U$5654 ( \14458_14760 , RIdf23a28_1782, \9183_9482 );
and \U$5655 ( \14459_14761 , RIfc823d0_6504, \9185_9484 );
and \U$5656 ( \14460_14762 , RIdf223a8_1766, \9187_9486 );
and \U$5657 ( \14461_14763 , RIdf20d28_1750, \9189_9488 );
and \U$5658 ( \14462_14764 , RIdf1bd00_1693, \9191_9490 );
and \U$5659 ( \14463_14765 , RIdf1a7e8_1678, \9193_9492 );
and \U$5660 ( \14464_14766 , RIdf18790_1655, \9195_9494 );
and \U$5661 ( \14465_14767 , RIdf15a90_1623, \9197_9496 );
and \U$5662 ( \14466_14768 , RIdf12d90_1591, \9199_9498 );
and \U$5663 ( \14467_14769 , RIdf10090_1559, \9201_9500 );
and \U$5664 ( \14468_14770 , RIdf0d390_1527, \9203_9502 );
and \U$5665 ( \14469_14771 , RIdf0a690_1495, \9205_9504 );
and \U$5666 ( \14470_14772 , RIdf07990_1463, \9207_9506 );
and \U$5667 ( \14471_14773 , RIdf04c90_1431, \9209_9508 );
and \U$5668 ( \14472_14774 , RIdeff290_1367, \9211_9510 );
and \U$5669 ( \14473_14775 , RIdefc590_1335, \9213_9512 );
and \U$5670 ( \14474_14776 , RIdef9890_1303, \9215_9514 );
and \U$5671 ( \14475_14777 , RIdef6b90_1271, \9217_9516 );
and \U$5672 ( \14476_14778 , RIdef3e90_1239, \9219_9518 );
and \U$5673 ( \14477_14779 , RIdef1190_1207, \9221_9520 );
and \U$5674 ( \14478_14780 , RIdeee490_1175, \9223_9522 );
and \U$5675 ( \14479_14781 , RIdeeb790_1143, \9225_9524 );
and \U$5676 ( \14480_14782 , RIee25be8_4888, \9227_9526 );
and \U$5677 ( \14481_14783 , RIfc6af28_6239, \9229_9528 );
and \U$5678 ( \14482_14784 , RIee23fc8_4868, \9231_9530 );
and \U$5679 ( \14483_14785 , RIfccf680_7382, \9233_9532 );
and \U$5680 ( \14484_14786 , RIdee5d90_1079, \9235_9534 );
and \U$5681 ( \14485_14787 , RIdee4008_1058, \9237_9536 );
and \U$5682 ( \14486_14788 , RIdee1ce0_1033, \9239_9538 );
and \U$5683 ( \14487_14789 , RIdedfdf0_1011, \9241_9540 );
and \U$5684 ( \14488_14790 , RIfc6b090_6240, \9243_9542 );
and \U$5685 ( \14489_14791 , RIfc534e0_5970, \9245_9544 );
and \U$5686 ( \14490_14792 , RIfca5920_6906, \9247_9546 );
and \U$5687 ( \14491_14793 , RIfc66770_6188, \9249_9548 );
and \U$5688 ( \14492_14794 , RIfe8f6d0_7976, \9251_9550 );
and \U$5689 ( \14493_14795 , RIded87d0_927, \9253_9552 );
and \U$5690 ( \14494_14796 , RIfe8f568_7975, \9255_9554 );
and \U$5691 ( \14495_14797 , RIded42e8_878, \9257_9556 );
and \U$5692 ( \14496_14798 , RIded1fc0_853, \9259_9558 );
and \U$5693 ( \14497_14799 , RIdecf2c0_821, \9261_9560 );
and \U$5694 ( \14498_14800 , RIdecc5c0_789, \9263_9562 );
and \U$5695 ( \14499_14801 , RIdec98c0_757, \9265_9564 );
and \U$5696 ( \14500_14802 , RIdeb5dc0_533, \9267_9566 );
and \U$5697 ( \14501_14803 , RIde9a0e8_341, \9269_9568 );
and \U$5698 ( \14502_14804 , RIe16f9c8_2647, \9271_9570 );
and \U$5699 ( \14503_14805 , RIe15b7c0_2418, \9273_9572 );
and \U$5700 ( \14504_14806 , RIe144fc0_2162, \9275_9574 );
and \U$5701 ( \14505_14807 , RIdf399b8_2032, \9277_9576 );
and \U$5702 ( \14506_14808 , RIdf2e018_1900, \9279_9578 );
and \U$5703 ( \14507_14809 , RIdf1e898_1724, \9281_9580 );
and \U$5704 ( \14508_14810 , RIdf01f90_1399, \9283_9582 );
and \U$5705 ( \14509_14811 , RIdee8a90_1111, \9285_9584 );
and \U$5706 ( \14510_14812 , RIdedd7f8_984, \9287_9586 );
and \U$5707 ( \14511_14813 , RIde80030_214, \9289_9588 );
or \U$5708 ( \14512_14814 , \14448_14750 , \14449_14751 , \14450_14752 , \14451_14753 , \14452_14754 , \14453_14755 , \14454_14756 , \14455_14757 , \14456_14758 , \14457_14759 , \14458_14760 , \14459_14761 , \14460_14762 , \14461_14763 , \14462_14764 , \14463_14765 , \14464_14766 , \14465_14767 , \14466_14768 , \14467_14769 , \14468_14770 , \14469_14771 , \14470_14772 , \14471_14773 , \14472_14774 , \14473_14775 , \14474_14776 , \14475_14777 , \14476_14778 , \14477_14779 , \14478_14780 , \14479_14781 , \14480_14782 , \14481_14783 , \14482_14784 , \14483_14785 , \14484_14786 , \14485_14787 , \14486_14788 , \14487_14789 , \14488_14790 , \14489_14791 , \14490_14792 , \14491_14793 , \14492_14794 , \14493_14795 , \14494_14796 , \14495_14797 , \14496_14798 , \14497_14799 , \14498_14800 , \14499_14801 , \14500_14802 , \14501_14803 , \14502_14804 , \14503_14805 , \14504_14806 , \14505_14807 , \14506_14808 , \14507_14809 , \14508_14810 , \14509_14811 , \14510_14812 , \14511_14813 );
or \U$5709 ( \14513_14815 , \14447_14749 , \14512_14814 );
_DC \g658f/U$1 ( \14514 , \14513_14815 , \9298_9597 );
and \U$5710 ( \14515_14817 , RIe19ee58_3185, \8760_9059 );
and \U$5711 ( \14516_14818 , RIe19c158_3153, \8762_9061 );
and \U$5712 ( \14517_14819 , RIf145bf8_5253, \8764_9063 );
and \U$5713 ( \14518_14820 , RIe199458_3121, \8766_9065 );
and \U$5714 ( \14519_14821 , RIfe8f298_7973, \8768_9067 );
and \U$5715 ( \14520_14822 , RIe196758_3089, \8770_9069 );
and \U$5716 ( \14521_14823 , RIe193a58_3057, \8772_9071 );
and \U$5717 ( \14522_14824 , RIe190d58_3025, \8774_9073 );
and \U$5718 ( \14523_14825 , RIe18b358_2961, \8776_9075 );
and \U$5719 ( \14524_14826 , RIe188658_2929, \8778_9077 );
and \U$5720 ( \14525_14827 , RIfe8f130_7972, \8780_9079 );
and \U$5721 ( \14526_14828 , RIe185958_2897, \8782_9081 );
and \U$5722 ( \14527_14829 , RIfc9f278_6833, \8784_9083 );
and \U$5723 ( \14528_14830 , RIe182c58_2865, \8786_9085 );
and \U$5724 ( \14529_14831 , RIe17ff58_2833, \8788_9087 );
and \U$5725 ( \14530_14832 , RIe17d258_2801, \8790_9089 );
and \U$5726 ( \14531_14833 , RIf1427f0_5216, \8792_9091 );
and \U$5727 ( \14532_14834 , RIfe8efc8_7971, \8794_9093 );
and \U$5728 ( \14533_14835 , RIe1779c0_2738, \8796_9095 );
and \U$5729 ( \14534_14836 , RIe1768e0_2726, \8798_9097 );
and \U$5730 ( \14535_14837 , RIfc81e30_6500, \8800_9099 );
and \U$5731 ( \14536_14838 , RIfc9ff20_6842, \8802_9101 );
and \U$5732 ( \14537_14839 , RIfca0088_6843, \8804_9103 );
and \U$5733 ( \14538_14840 , RIfc81b60_6498, \8806_9105 );
and \U$5734 ( \14539_14841 , RIfce5778_7633, \8808_9107 );
and \U$5735 ( \14540_14842 , RIfce08b8_7577, \8810_9109 );
and \U$5736 ( \14541_14843 , RIfc815c0_6494, \8812_9111 );
and \U$5737 ( \14542_14844 , RIe174cc0_2706, \8814_9113 );
and \U$5738 ( \14543_14845 , RIfca04c0_6846, \8816_9115 );
and \U$5739 ( \14544_14846 , RIfc53eb8_5977, \8818_9117 );
and \U$5740 ( \14545_14847 , RIfcc65a8_7279, \8820_9119 );
and \U$5741 ( \14546_14848 , RIfc80d50_6488, \8822_9121 );
and \U$5742 ( \14547_14849 , RIfc804e0_6482, \8824_9123 );
and \U$5743 ( \14548_14850 , RIe2251b0_4712, \8826_9125 );
and \U$5744 ( \14549_14851 , RIfc80378_6481, \8828_9127 );
and \U$5745 ( \14550_14852 , RIe2224b0_4680, \8830_9129 );
and \U$5746 ( \14551_14853 , RIfcb5910_7088, \8832_9131 );
and \U$5747 ( \14552_14854 , RIe21f7b0_4648, \8834_9133 );
and \U$5748 ( \14553_14855 , RIe219db0_4584, \8836_9135 );
and \U$5749 ( \14554_14856 , RIe2170b0_4552, \8838_9137 );
and \U$5750 ( \14555_14857 , RIfca01f0_6844, \8840_9139 );
and \U$5751 ( \14556_14858 , RIe2143b0_4520, \8842_9141 );
and \U$5752 ( \14557_14859 , RIfc82c40_6510, \8844_9143 );
and \U$5753 ( \14558_14860 , RIe2116b0_4488, \8846_9145 );
and \U$5754 ( \14559_14861 , RIfc7f6d0_6472, \8848_9147 );
and \U$5755 ( \14560_14862 , RIe20e9b0_4456, \8850_9149 );
and \U$5756 ( \14561_14863 , RIe20bcb0_4424, \8852_9151 );
and \U$5757 ( \14562_14864 , RIe208fb0_4392, \8854_9153 );
and \U$5758 ( \14563_14865 , RIf167528_5635, \8856_9155 );
and \U$5759 ( \14564_14866 , RIf1665b0_5624, \8858_9157 );
and \U$5760 ( \14565_14867 , RIe203718_4329, \8860_9159 );
and \U$5761 ( \14566_14868 , RIe201c60_4310, \8862_9161 );
and \U$5762 ( \14567_14869 , RIfc9da90_6816, \8864_9163 );
and \U$5763 ( \14568_14870 , RIfcc5360_7266, \8866_9165 );
and \U$5764 ( \14569_14871 , RIf163748_5591, \8868_9167 );
and \U$5765 ( \14570_14872 , RIf162668_5579, \8870_9169 );
and \U$5766 ( \14571_14873 , RIfc7e320_6458, \8872_9171 );
and \U$5767 ( \14572_14874 , RIfc87998_6565, \8874_9173 );
and \U$5768 ( \14573_14875 , RIe1fd610_4260, \8876_9175 );
and \U$5769 ( \14574_14876 , RIe1fc3c8_4247, \8878_9177 );
and \U$5770 ( \14575_14877 , RIf15d370_5520, \8880_9179 );
and \U$5771 ( \14576_14878 , RIf15c128_5507, \8882_9181 );
and \U$5772 ( \14577_14879 , RIfcc5d38_7273, \8884_9183 );
and \U$5773 ( \14578_14880 , RIfce7d70_7660, \8886_9185 );
or \U$5774 ( \14579_14881 , \14515_14817 , \14516_14818 , \14517_14819 , \14518_14820 , \14519_14821 , \14520_14822 , \14521_14823 , \14522_14824 , \14523_14825 , \14524_14826 , \14525_14827 , \14526_14828 , \14527_14829 , \14528_14830 , \14529_14831 , \14530_14832 , \14531_14833 , \14532_14834 , \14533_14835 , \14534_14836 , \14535_14837 , \14536_14838 , \14537_14839 , \14538_14840 , \14539_14841 , \14540_14842 , \14541_14843 , \14542_14844 , \14543_14845 , \14544_14846 , \14545_14847 , \14546_14848 , \14547_14849 , \14548_14850 , \14549_14851 , \14550_14852 , \14551_14853 , \14552_14854 , \14553_14855 , \14554_14856 , \14555_14857 , \14556_14858 , \14557_14859 , \14558_14860 , \14559_14861 , \14560_14862 , \14561_14863 , \14562_14864 , \14563_14865 , \14564_14866 , \14565_14867 , \14566_14868 , \14567_14869 , \14568_14870 , \14569_14871 , \14570_14872 , \14571_14873 , \14572_14874 , \14573_14875 , \14574_14876 , \14575_14877 , \14576_14878 , \14577_14879 , \14578_14880 );
and \U$5775 ( \14580_14882 , RIfc4bd58_5885, \8889_9188 );
and \U$5776 ( \14581_14883 , RIfc55c40_5998, \8891_9190 );
and \U$5777 ( \14582_14884 , RIfca2ab8_6873, \8893_9192 );
and \U$5778 ( \14583_14885 , RIe1fb450_4236, \8895_9194 );
and \U$5779 ( \14584_14886 , RIf156890_5444, \8897_9196 );
and \U$5780 ( \14585_14887 , RIfcd5ff8_7457, \8899_9198 );
and \U$5781 ( \14586_14888 , RIf154dd8_5425, \8901_9200 );
and \U$5782 ( \14587_14889 , RIfec2aa8_8335, \8903_9202 );
and \U$5783 ( \14588_14890 , RIfcb4b00_7078, \8905_9204 );
and \U$5784 ( \14589_14891 , RIfcd9400_7494, \8907_9206 );
and \U$5785 ( \14590_14892 , RIf151160_5382, \8909_9208 );
and \U$5786 ( \14591_14893 , RIe1f4808_4159, \8911_9210 );
and \U$5787 ( \14592_14894 , RIfc44738_5801, \8913_9212 );
and \U$5788 ( \14593_14895 , RIfc90908_6667, \8915_9214 );
and \U$5789 ( \14594_14896 , RIf14e5c8_5351, \8917_9216 );
and \U$5790 ( \14595_14897 , RIe1ef510_4100, \8919_9218 );
and \U$5791 ( \14596_14898 , RIe1ecf18_4073, \8921_9220 );
and \U$5792 ( \14597_14899 , RIe1ea218_4041, \8923_9222 );
and \U$5793 ( \14598_14900 , RIe1e7518_4009, \8925_9224 );
and \U$5794 ( \14599_14901 , RIe1e4818_3977, \8927_9226 );
and \U$5795 ( \14600_14902 , RIe1e1b18_3945, \8929_9228 );
and \U$5796 ( \14601_14903 , RIe1dee18_3913, \8931_9230 );
and \U$5797 ( \14602_14904 , RIe1dc118_3881, \8933_9232 );
and \U$5798 ( \14603_14905 , RIe1d9418_3849, \8935_9234 );
and \U$5799 ( \14604_14906 , RIe1d3a18_3785, \8937_9236 );
and \U$5800 ( \14605_14907 , RIe1d0d18_3753, \8939_9238 );
and \U$5801 ( \14606_14908 , RIe1ce018_3721, \8941_9240 );
and \U$5802 ( \14607_14909 , RIe1cb318_3689, \8943_9242 );
and \U$5803 ( \14608_14910 , RIe1c8618_3657, \8945_9244 );
and \U$5804 ( \14609_14911 , RIe1c5918_3625, \8947_9246 );
and \U$5805 ( \14610_14912 , RIe1c2c18_3593, \8949_9248 );
and \U$5806 ( \14611_14913 , RIe1bff18_3561, \8951_9250 );
and \U$5807 ( \14612_14914 , RIf14d218_5337, \8953_9252 );
and \U$5808 ( \14613_14915 , RIfe8ee60_7970, \8955_9254 );
and \U$5809 ( \14614_14916 , RIfea8090_8228, \8957_9256 );
and \U$5810 ( \14615_14917 , RIe1b84c0_3474, \8959_9258 );
and \U$5811 ( \14616_14918 , RIf14aab8_5309, \8961_9260 );
and \U$5812 ( \14617_14919 , RIfc6c170_6252, \8963_9262 );
and \U$5813 ( \14618_14920 , RIe1b6468_3451, \8965_9264 );
and \U$5814 ( \14619_14921 , RIe1b49b0_3432, \8967_9266 );
and \U$5815 ( \14620_14922 , RIfcafad8_7021, \8969_9268 );
and \U$5816 ( \14621_14923 , RIfcaa948_6963, \8971_9270 );
and \U$5817 ( \14622_14924 , RIfe8ecf8_7969, \8973_9272 );
and \U$5818 ( \14623_14925 , RIfe8f400_7974, \8975_9274 );
and \U$5819 ( \14624_14926 , RIfc67f58_6205, \8977_9276 );
and \U$5820 ( \14625_14927 , RIfca8ff8_6945, \8979_9278 );
and \U$5821 ( \14626_14928 , RIfe8eb90_7968, \8981_9280 );
and \U$5822 ( \14627_14929 , RIe1abe78_3333, \8983_9282 );
and \U$5823 ( \14628_14930 , RIe1aa258_3313, \8985_9284 );
and \U$5824 ( \14629_14931 , RIe1a7558_3281, \8987_9286 );
and \U$5825 ( \14630_14932 , RIe1a4858_3249, \8989_9288 );
and \U$5826 ( \14631_14933 , RIe1a1b58_3217, \8991_9290 );
and \U$5827 ( \14632_14934 , RIe18e058_2993, \8993_9292 );
and \U$5828 ( \14633_14935 , RIe17a558_2769, \8995_9294 );
and \U$5829 ( \14634_14936 , RIe227eb0_4744, \8997_9296 );
and \U$5830 ( \14635_14937 , RIe21cab0_4616, \8999_9298 );
and \U$5831 ( \14636_14938 , RIe2062b0_4360, \9001_9300 );
and \U$5832 ( \14637_14939 , RIe200310_4292, \9003_9302 );
and \U$5833 ( \14638_14940 , RIe1f96c8_4215, \9005_9304 );
and \U$5834 ( \14639_14941 , RIe1f2210_4132, \9007_9306 );
and \U$5835 ( \14640_14942 , RIe1d6718_3817, \9009_9308 );
and \U$5836 ( \14641_14943 , RIe1bd218_3529, \9011_9310 );
and \U$5837 ( \14642_14944 , RIe1b0090_3380, \9013_9312 );
and \U$5838 ( \14643_14945 , RIe1726c8_2679, \9015_9314 );
or \U$5839 ( \14644_14946 , \14580_14882 , \14581_14883 , \14582_14884 , \14583_14885 , \14584_14886 , \14585_14887 , \14586_14888 , \14587_14889 , \14588_14890 , \14589_14891 , \14590_14892 , \14591_14893 , \14592_14894 , \14593_14895 , \14594_14896 , \14595_14897 , \14596_14898 , \14597_14899 , \14598_14900 , \14599_14901 , \14600_14902 , \14601_14903 , \14602_14904 , \14603_14905 , \14604_14906 , \14605_14907 , \14606_14908 , \14607_14909 , \14608_14910 , \14609_14911 , \14610_14912 , \14611_14913 , \14612_14914 , \14613_14915 , \14614_14916 , \14615_14917 , \14616_14918 , \14617_14919 , \14618_14920 , \14619_14921 , \14620_14922 , \14621_14923 , \14622_14924 , \14623_14925 , \14624_14926 , \14625_14927 , \14626_14928 , \14627_14929 , \14628_14930 , \14629_14931 , \14630_14932 , \14631_14933 , \14632_14934 , \14633_14935 , \14634_14936 , \14635_14937 , \14636_14938 , \14637_14939 , \14638_14940 , \14639_14941 , \14640_14942 , \14641_14943 , \14642_14944 , \14643_14945 );
or \U$5840 ( \14645_14947 , \14579_14881 , \14644_14946 );
_DC \g6590/U$1 ( \14646 , \14645_14947 , \9024_9323 );
and g6591_GF_PartitionCandidate( \14647_14949_nG6591 , \14514 , \14646 );
buf \U$5841 ( \14648_14950 , \14647_14949_nG6591 );
and \U$5842 ( \14649_14951 , \14648_14950 , \10389_10691 );
nor \U$5843 ( \14650_14952 , \14382_14684 , \14649_14951 );
xnor \U$5844 ( \14651_14953 , \14650_14952 , \10678_10980 );
and \U$5845 ( \14652_14954 , \10686_10988 , \13755_14054 );
and \U$5846 ( \14653_14955 , \10968_11270 , \13390_13692 );
nor \U$5847 ( \14654_14956 , \14652_14954 , \14653_14955 );
xnor \U$5848 ( \14655_14957 , \14654_14956 , \13736_14035 );
xor \U$5849 ( \14656_14958 , \14651_14953 , \14655_14957 );
_DC \g4d22/U$1 ( \14657 , \14513_14815 , \9298_9597 );
_DC \g4da6/U$1 ( \14658 , \14645_14947 , \9024_9323 );
xor g4da7_GF_PartitionCandidate( \14659_14961_nG4da7 , \14657 , \14658 );
buf \U$5850 ( \14660_14962 , \14659_14961_nG4da7 );
xor \U$5851 ( \14661_14963 , \14660_14962 , \13733_14032 );
and \U$5852 ( \14662_14964 , \10385_10687 , \14661_14963 );
xor \U$5853 ( \14663_14965 , \14656_14958 , \14662_14964 );
xor \U$5854 ( \14664_14966 , \14381_14683 , \14663_14965 );
and \U$5855 ( \14665_14967 , \13728_14027 , \13737_14036 );
and \U$5856 ( \14666_14968 , \12470_12769 , \11275_11574 );
and \U$5857 ( \14667_14969 , \13377_13679 , \10976_11278 );
nor \U$5858 ( \14668_14970 , \14666_14968 , \14667_14969 );
xnor \U$5859 ( \14669_14971 , \14668_14970 , \11281_11580 );
xor \U$5860 ( \14670_14972 , \14665_14967 , \14669_14971 );
and \U$5861 ( \14671_14973 , \11287_11586 , \12491_12790 );
and \U$5862 ( \14672_14974 , \12146_12448 , \12159_12461 );
nor \U$5863 ( \14673_14975 , \14671_14973 , \14672_14974 );
xnor \U$5864 ( \14674_14976 , \14673_14975 , \12481_12780 );
xor \U$5865 ( \14675_14977 , \14670_14972 , \14674_14976 );
xor \U$5866 ( \14676_14978 , \14664_14966 , \14675_14977 );
xor \U$5867 ( \14677_14979 , \14377_14679 , \14676_14978 );
and \U$5868 ( \14678_14980 , \13761_14060 , \13765_14064 );
and \U$5869 ( \14679_14981 , \13766_14065 , \13769_14068 );
or \U$5870 ( \14680_14982 , \14678_14980 , \14679_14981 );
xor \U$5871 ( \14681_14983 , \14677_14979 , \14680_14982 );
buf g9bf6_GF_PartitionCandidate( \14682_14984_nG9bf6 , \14681_14983 );
and \U$5872 ( \14683_14985 , \10402_10704 , \14682_14984_nG9bf6 );
or \U$5873 ( \14684_14986 , \14373_14675 , \14683_14985 );
xor \U$5874 ( \14685_14987 , \10399_10703 , \14684_14986 );
buf \U$5875 ( \14686_14988 , \14685_14987 );
buf \U$5877 ( \14687_14989 , \14686_14988 );
xor \U$5878 ( \14688_14990 , \14372_14674 , \14687_14989 );
buf \U$5879 ( \14689_14991 , \14688_14990 );
xor \U$5880 ( \14690_14992 , \14341_14643 , \14689_14991 );
and \U$5881 ( \14691_14993 , \13454_13753 , \13456_13755 );
and \U$5882 ( \14692_14994 , \13454_13753 , \13776_14075 );
and \U$5883 ( \14693_14995 , \13456_13755 , \13776_14075 );
or \U$5884 ( \14694_14996 , \14691_14993 , \14692_14994 , \14693_14995 );
buf \U$5885 ( \14695_14997 , \14694_14996 );
xor \U$5886 ( \14696_14998 , \14690_14992 , \14695_14997 );
and \U$5887 ( \14697_14999 , \13780_14079 , \14696_14998 );
and \U$5888 ( \14698_15000 , \14335_14637 , \14696_14998 );
or \U$5889 ( \14699_15001 , \14336_14638 , \14697_14999 , \14698_15000 );
and \U$5890 ( \14700_15002 , \14366_14668 , \14371_14673 );
and \U$5891 ( \14701_15003 , \14366_14668 , \14687_14989 );
and \U$5892 ( \14702_15004 , \14371_14673 , \14687_14989 );
or \U$5893 ( \14703_15005 , \14700_15002 , \14701_15003 , \14702_15004 );
buf \U$5894 ( \14704_15006 , \14703_15005 );
and \U$5895 ( \14705_15007 , \14328_14627 , \14332_14634 );
buf \U$5896 ( \14706_15008 , \14705_15007 );
buf \U$5898 ( \14707_15009 , \14706_15008 );
not \U$5519 ( \14708_14629 , \14329_14628 );
xor \U$5520 ( \14709_14630 , \14323_14622_nG443c , \14326_14625_nG443f );
and \U$5521 ( \14710_14631 , \14708_14629 , \14709_14630 );
and \U$5899 ( \14711_15010 , \14710_14631 , \10392_10694_nG9c0e );
and \U$5900 ( \14712_15011 , \14329_14628 , \10693_10995_nG9c0b );
or \U$5901 ( \14713_15012 , \14711_15010 , \14712_15011 );
xor \U$5902 ( \14714_15013 , \14328_14627 , \14713_15012 );
buf \U$5903 ( \14715_15014 , \14714_15013 );
buf \U$5905 ( \14716_15015 , \14715_15014 );
xor \U$5906 ( \14717_15016 , \14707_15009 , \14716_15015 );
buf \U$5907 ( \14718_15017 , \14717_15016 );
and \U$5908 ( \14719_15018 , \13431_13370 , \10981_11283_nG9c08 );
and \U$5909 ( \14720_15019 , \13068_13367 , \11299_11598_nG9c05 );
or \U$5910 ( \14721_15020 , \14719_15018 , \14720_15019 );
xor \U$5911 ( \14722_15021 , \13067_13366 , \14721_15020 );
buf \U$5912 ( \14723_15022 , \14722_15021 );
buf \U$5914 ( \14724_15023 , \14723_15022 );
xor \U$5915 ( \14725_15024 , \14718_15017 , \14724_15023 );
and \U$5916 ( \14726_15025 , \12183_12157 , \12168_12470_nG9c02 );
and \U$5917 ( \14727_15026 , \11855_12154 , \12502_12801_nG9bff );
or \U$5918 ( \14728_15027 , \14726_15025 , \14727_15026 );
xor \U$5919 ( \14729_15028 , \11854_12153 , \14728_15027 );
buf \U$5920 ( \14730_15029 , \14729_15028 );
buf \U$5922 ( \14731_15030 , \14730_15029 );
xor \U$5923 ( \14732_15031 , \14725_15024 , \14731_15030 );
buf \U$5924 ( \14733_15032 , \14732_15031 );
and \U$5925 ( \14734_15033 , \14351_14653 , \14357_14659 );
and \U$5926 ( \14735_15034 , \14351_14653 , \14364_14666 );
and \U$5927 ( \14736_15035 , \14357_14659 , \14364_14666 );
or \U$5928 ( \14737_15036 , \14734_15033 , \14735_15034 , \14736_15035 );
buf \U$5929 ( \14738_15037 , \14737_15036 );
and \U$5930 ( \14739_15038 , \14343_14645 , \14349_14651 );
buf \U$5931 ( \14740_15039 , \14739_15038 );
xor \U$5932 ( \14741_15040 , \14738_15037 , \14740_15039 );
and \U$5933 ( \14742_15041 , \10996_10421 , \13403_13705_nG9bfc );
and \U$5934 ( \14743_15042 , \10119_10418 , \13771_14070_nG9bf9 );
or \U$5935 ( \14744_15043 , \14742_15041 , \14743_15042 );
xor \U$5936 ( \14745_15044 , \10118_10417 , \14744_15043 );
buf \U$5937 ( \14746_15045 , \14745_15044 );
buf \U$5939 ( \14747_15046 , \14746_15045 );
xor \U$5940 ( \14748_15047 , \14741_15040 , \14747_15046 );
buf \U$5941 ( \14749_15048 , \14748_15047 );
xor \U$5942 ( \14750_15049 , \14733_15032 , \14749_15048 );
and \U$5943 ( \14751_15050 , \10411_10707 , \14682_14984_nG9bf6 );
and \U$5944 ( \14752_15051 , \14665_14967 , \14669_14971 );
and \U$5945 ( \14753_15052 , \14669_14971 , \14674_14976 );
and \U$5946 ( \14754_15053 , \14665_14967 , \14674_14976 );
or \U$5947 ( \14755_15054 , \14752_15051 , \14753_15052 , \14754_15053 );
and \U$5948 ( \14756_15055 , \14648_14950 , \10681_10983 );
and \U$5949 ( \14757_15056 , RIdec6d28_726, \9034_9333 );
and \U$5950 ( \14758_15057 , RIdec4028_694, \9036_9335 );
and \U$5951 ( \14759_15058 , RIee20bc0_4831, \9038_9337 );
and \U$5952 ( \14760_15059 , RIdec1328_662, \9040_9339 );
and \U$5953 ( \14761_15060 , RIfcbaed8_7149, \9042_9341 );
and \U$5954 ( \14762_15061 , RIdebe628_630, \9044_9343 );
and \U$5955 ( \14763_15062 , RIdebb928_598, \9046_9345 );
and \U$5956 ( \14764_15063 , RIdeb8c28_566, \9048_9347 );
and \U$5957 ( \14765_15064 , RIfc412b8_5767, \9050_9349 );
and \U$5958 ( \14766_15065 , RIdeb3228_502, \9052_9351 );
and \U$5959 ( \14767_15066 , RIfc9ea08_6827, \9054_9353 );
and \U$5960 ( \14768_15067 , RIdeb0528_470, \9056_9355 );
and \U$5961 ( \14769_15068 , RIee1e028_4800, \9058_9357 );
and \U$5962 ( \14770_15069 , RIdead828_438, \9060_9359 );
and \U$5963 ( \14771_15070 , RIdea7630_406, \9062_9361 );
and \U$5964 ( \14772_15071 , RIdea0d30_374, \9064_9363 );
and \U$5965 ( \14773_15072 , RIfcbac08_7147, \9066_9365 );
and \U$5966 ( \14774_15073 , RIfc55538_5993, \9068_9367 );
and \U$5967 ( \14775_15074 , RIfcba668_7143, \9070_9369 );
and \U$5968 ( \14776_15075 , RIfc4af48_5875, \9072_9371 );
and \U$5969 ( \14777_15076 , RIfe912f0_7996, \9074_9373 );
and \U$5970 ( \14778_15077 , RIfe91458_7997, \9076_9375 );
and \U$5971 ( \14779_15078 , RIde8be80_272, \9078_9377 );
and \U$5972 ( \14780_15079 , RIde87ce0_252, \9080_9379 );
and \U$5973 ( \14781_15080 , RIfc85238_6537, \9082_9381 );
and \U$5974 ( \14782_15081 , RIfc88640_6574, \9084_9383 );
and \U$5975 ( \14783_15082 , RIfcda210_7504, \9086_9385 );
and \U$5976 ( \14784_15083 , RIfcd5788_7451, \9088_9387 );
and \U$5977 ( \14785_15084 , RIee39418_5110, \9090_9389 );
and \U$5978 ( \14786_15085 , RIe16ce30_2616, \9092_9391 );
and \U$5979 ( \14787_15086 , RIfc884d8_6573, \9094_9393 );
and \U$5980 ( \14788_15087 , RIe169320_2574, \9096_9395 );
and \U$5981 ( \14789_15088 , RIe166d28_2547, \9098_9397 );
and \U$5982 ( \14790_15089 , RIe164028_2515, \9100_9399 );
and \U$5983 ( \14791_15090 , RIfe90918_7989, \9102_9401 );
and \U$5984 ( \14792_15091 , RIe161328_2483, \9104_9403 );
and \U$5985 ( \14793_15092 , RIee36880_5079, \9106_9405 );
and \U$5986 ( \14794_15093 , RIe15e628_2451, \9108_9407 );
and \U$5987 ( \14795_15094 , RIe158c28_2387, \9110_9409 );
and \U$5988 ( \14796_15095 , RIe155f28_2355, \9112_9411 );
and \U$5989 ( \14797_15096 , RIfe91188_7995, \9114_9413 );
and \U$5990 ( \14798_15097 , RIe153228_2323, \9116_9415 );
and \U$5991 ( \14799_15098 , RIfe91020_7994, \9118_9417 );
and \U$5992 ( \14800_15099 , RIe150528_2291, \9120_9419 );
and \U$5993 ( \14801_15100 , RIfcda378_7505, \9122_9421 );
and \U$5994 ( \14802_15101 , RIe14d828_2259, \9124_9423 );
and \U$5995 ( \14803_15102 , RIe14ab28_2227, \9126_9425 );
and \U$5996 ( \14804_15103 , RIe147e28_2195, \9128_9427 );
and \U$5997 ( \14805_15104 , RIfe90eb8_7993, \9130_9429 );
and \U$5998 ( \14806_15105 , RIfe90d50_7992, \9132_9431 );
and \U$5999 ( \14807_15106 , RIfcb99c0_7134, \9134_9433 );
and \U$6000 ( \14808_15107 , RIfc9c2a8_6799, \9136_9435 );
and \U$6001 ( \14809_15108 , RIfe90be8_7991, \9138_9437 );
and \U$6002 ( \14810_15109 , RIfe90a80_7990, \9140_9439 );
and \U$6003 ( \14811_15110 , RIdf3e008_2082, \9142_9441 );
and \U$6004 ( \14812_15111 , RIdf3bce0_2057, \9144_9443 );
and \U$6005 ( \14813_15112 , RIfcec690_7712, \9146_9445 );
and \U$6006 ( \14814_15113 , RIee30778_5010, \9148_9447 );
and \U$6007 ( \14815_15114 , RIfc87dd0_6568, \9150_9449 );
and \U$6008 ( \14816_15115 , RIee2e5b8_4986, \9152_9451 );
and \U$6009 ( \14817_15116 , RIdf36e20_2001, \9154_9453 );
and \U$6010 ( \14818_15117 , RIdf346c0_1973, \9156_9455 );
and \U$6011 ( \14819_15118 , RIdf32668_1950, \9158_9457 );
and \U$6012 ( \14820_15119 , RIdf30070_1923, \9160_9459 );
or \U$6013 ( \14821_15120 , \14757_15056 , \14758_15057 , \14759_15058 , \14760_15059 , \14761_15060 , \14762_15061 , \14763_15062 , \14764_15063 , \14765_15064 , \14766_15065 , \14767_15066 , \14768_15067 , \14769_15068 , \14770_15069 , \14771_15070 , \14772_15071 , \14773_15072 , \14774_15073 , \14775_15074 , \14776_15075 , \14777_15076 , \14778_15077 , \14779_15078 , \14780_15079 , \14781_15080 , \14782_15081 , \14783_15082 , \14784_15083 , \14785_15084 , \14786_15085 , \14787_15086 , \14788_15087 , \14789_15088 , \14790_15089 , \14791_15090 , \14792_15091 , \14793_15092 , \14794_15093 , \14795_15094 , \14796_15095 , \14797_15096 , \14798_15097 , \14799_15098 , \14800_15099 , \14801_15100 , \14802_15101 , \14803_15102 , \14804_15103 , \14805_15104 , \14806_15105 , \14807_15106 , \14808_15107 , \14809_15108 , \14810_15109 , \14811_15110 , \14812_15111 , \14813_15112 , \14814_15113 , \14815_15114 , \14816_15115 , \14817_15116 , \14818_15117 , \14819_15118 , \14820_15119 );
and \U$6014 ( \14822_15121 , RIee2c998_4966, \9163_9462 );
and \U$6015 ( \14823_15122 , RIee2aee0_4947, \9165_9464 );
and \U$6016 ( \14824_15123 , RIee299c8_4932, \9167_9466 );
and \U$6017 ( \14825_15124 , RIee28618_4918, \9169_9468 );
and \U$6018 ( \14826_15125 , RIfe90378_7985, \9171_9470 );
and \U$6019 ( \14827_15126 , RIfe907b0_7988, \9173_9472 );
and \U$6020 ( \14828_15127 , RIfe904e0_7986, \9175_9474 );
and \U$6021 ( \14829_15128 , RIfe90648_7987, \9177_9476 );
and \U$6022 ( \14830_15129 , RIfc9d928_6815, \9179_9478 );
and \U$6023 ( \14831_15130 , RIfc86048_6547, \9181_9480 );
and \U$6024 ( \14832_15131 , RIfcb92b8_7129, \9183_9482 );
and \U$6025 ( \14833_15132 , RIfc4ee90_5920, \9185_9484 );
and \U$6026 ( \14834_15133 , RIfc86a20_6554, \9187_9486 );
and \U$6027 ( \14835_15134 , RIdf20e90_1751, \9189_9488 );
and \U$6028 ( \14836_15135 , RIfcb8fe8_7127, \9191_9490 );
and \U$6029 ( \14837_15136 , RIdf1a950_1679, \9193_9492 );
and \U$6030 ( \14838_15137 , RIdf188f8_1656, \9195_9494 );
and \U$6031 ( \14839_15138 , RIdf15bf8_1624, \9197_9496 );
and \U$6032 ( \14840_15139 , RIdf12ef8_1592, \9199_9498 );
and \U$6033 ( \14841_15140 , RIdf101f8_1560, \9201_9500 );
and \U$6034 ( \14842_15141 , RIdf0d4f8_1528, \9203_9502 );
and \U$6035 ( \14843_15142 , RIdf0a7f8_1496, \9205_9504 );
and \U$6036 ( \14844_15143 , RIdf07af8_1464, \9207_9506 );
and \U$6037 ( \14845_15144 , RIdf04df8_1432, \9209_9508 );
and \U$6038 ( \14846_15145 , RIdeff3f8_1368, \9211_9510 );
and \U$6039 ( \14847_15146 , RIdefc6f8_1336, \9213_9512 );
and \U$6040 ( \14848_15147 , RIdef99f8_1304, \9215_9514 );
and \U$6041 ( \14849_15148 , RIdef6cf8_1272, \9217_9516 );
and \U$6042 ( \14850_15149 , RIdef3ff8_1240, \9219_9518 );
and \U$6043 ( \14851_15150 , RIdef12f8_1208, \9221_9520 );
and \U$6044 ( \14852_15151 , RIdeee5f8_1176, \9223_9522 );
and \U$6045 ( \14853_15152 , RIdeeb8f8_1144, \9225_9524 );
and \U$6046 ( \14854_15153 , RIfc857d8_6541, \9227_9526 );
and \U$6047 ( \14855_15154 , RIee24dd8_4878, \9229_9528 );
and \U$6048 ( \14856_15155 , RIfc4ff70_5932, \9231_9530 );
and \U$6049 ( \14857_15156 , RIfc50240_5934, \9233_9532 );
and \U$6050 ( \14858_15157 , RIdee5ef8_1080, \9235_9534 );
and \U$6051 ( \14859_15158 , RIdee4170_1059, \9237_9536 );
and \U$6052 ( \14860_15159 , RIfe915c0_7998, \9239_9538 );
and \U$6053 ( \14861_15160 , RIdedff58_1012, \9241_9540 );
and \U$6054 ( \14862_15161 , RIfcd4810_7440, \9243_9542 );
and \U$6055 ( \14863_15162 , RIee22948_4852, \9245_9544 );
and \U$6056 ( \14864_15163 , RIfce1560_7586, \9247_9546 );
and \U$6057 ( \14865_15164 , RIee219d0_4841, \9249_9548 );
and \U$6058 ( \14866_15165 , RIdedac60_953, \9251_9550 );
and \U$6059 ( \14867_15166 , RIfe91728_7999, \9253_9552 );
and \U$6060 ( \14868_15167 , RIded64a8_902, \9255_9554 );
and \U$6061 ( \14869_15168 , RIfe91890_8000, \9257_9556 );
and \U$6062 ( \14870_15169 , RIded2128_854, \9259_9558 );
and \U$6063 ( \14871_15170 , RIdecf428_822, \9261_9560 );
and \U$6064 ( \14872_15171 , RIdecc728_790, \9263_9562 );
and \U$6065 ( \14873_15172 , RIdec9a28_758, \9265_9564 );
and \U$6066 ( \14874_15173 , RIdeb5f28_534, \9267_9566 );
and \U$6067 ( \14875_15174 , RIde9a430_342, \9269_9568 );
and \U$6068 ( \14876_15175 , RIe16fb30_2648, \9271_9570 );
and \U$6069 ( \14877_15176 , RIe15b928_2419, \9273_9572 );
and \U$6070 ( \14878_15177 , RIe145128_2163, \9275_9574 );
and \U$6071 ( \14879_15178 , RIdf39b20_2033, \9277_9576 );
and \U$6072 ( \14880_15179 , RIdf2e180_1901, \9279_9578 );
and \U$6073 ( \14881_15180 , RIdf1ea00_1725, \9281_9580 );
and \U$6074 ( \14882_15181 , RIdf020f8_1400, \9283_9582 );
and \U$6075 ( \14883_15182 , RIdee8bf8_1112, \9285_9584 );
and \U$6076 ( \14884_15183 , RIdedd960_985, \9287_9586 );
and \U$6077 ( \14885_15184 , RIde80378_215, \9289_9588 );
or \U$6078 ( \14886_15185 , \14822_15121 , \14823_15122 , \14824_15123 , \14825_15124 , \14826_15125 , \14827_15126 , \14828_15127 , \14829_15128 , \14830_15129 , \14831_15130 , \14832_15131 , \14833_15132 , \14834_15133 , \14835_15134 , \14836_15135 , \14837_15136 , \14838_15137 , \14839_15138 , \14840_15139 , \14841_15140 , \14842_15141 , \14843_15142 , \14844_15143 , \14845_15144 , \14846_15145 , \14847_15146 , \14848_15147 , \14849_15148 , \14850_15149 , \14851_15150 , \14852_15151 , \14853_15152 , \14854_15153 , \14855_15154 , \14856_15155 , \14857_15156 , \14858_15157 , \14859_15158 , \14860_15159 , \14861_15160 , \14862_15161 , \14863_15162 , \14864_15163 , \14865_15164 , \14866_15165 , \14867_15166 , \14868_15167 , \14869_15168 , \14870_15169 , \14871_15170 , \14872_15171 , \14873_15172 , \14874_15173 , \14875_15174 , \14876_15175 , \14877_15176 , \14878_15177 , \14879_15178 , \14880_15179 , \14881_15180 , \14882_15181 , \14883_15182 , \14884_15183 , \14885_15184 );
or \U$6079 ( \14887_15186 , \14821_15120 , \14886_15185 );
_DC \g6592/U$1 ( \14888 , \14887_15186 , \9298_9597 );
and \U$6080 ( \14889_15188 , RIe19efc0_3186, \8760_9059 );
and \U$6081 ( \14890_15189 , RIe19c2c0_3154, \8762_9061 );
and \U$6082 ( \14891_15190 , RIf145d60_5254, \8764_9063 );
and \U$6083 ( \14892_15191 , RIe1995c0_3122, \8766_9065 );
and \U$6084 ( \14893_15192 , RIfc637a0_6154, \8768_9067 );
and \U$6085 ( \14894_15193 , RIe1968c0_3090, \8770_9069 );
and \U$6086 ( \14895_15194 , RIe193bc0_3058, \8772_9071 );
and \U$6087 ( \14896_15195 , RIe190ec0_3026, \8774_9073 );
and \U$6088 ( \14897_15196 , RIe18b4c0_2962, \8776_9075 );
and \U$6089 ( \14898_15197 , RIe1887c0_2930, \8778_9077 );
and \U$6090 ( \14899_15198 , RIfc62af8_6145, \8780_9079 );
and \U$6091 ( \14900_15199 , RIe185ac0_2898, \8782_9081 );
and \U$6092 ( \14901_15200 , RIfe8fc70_7980, \8784_9083 );
and \U$6093 ( \14902_15201 , RIe182dc0_2866, \8786_9085 );
and \U$6094 ( \14903_15202 , RIe1800c0_2834, \8788_9087 );
and \U$6095 ( \14904_15203 , RIe17d3c0_2802, \8790_9089 );
and \U$6096 ( \14905_15204 , RIfe90210_7984, \8792_9091 );
and \U$6097 ( \14906_15205 , RIfe8ff40_7982, \8794_9093 );
and \U$6098 ( \14907_15206 , RIfc72f20_6330, \8796_9095 );
and \U$6099 ( \14908_15207 , RIe176a48_2727, \8798_9097 );
and \U$6100 ( \14909_15208 , RIfcaf6a0_7018, \8800_9099 );
and \U$6101 ( \14910_15209 , RIfc61040_6126, \8802_9101 );
and \U$6102 ( \14911_15210 , RIf13e8a8_5171, \8804_9103 );
and \U$6103 ( \14912_15211 , RIfe900a8_7983, \8806_9105 );
and \U$6104 ( \14913_15212 , RIee3caf0_5149, \8808_9107 );
and \U$6105 ( \14914_15213 , RIee3b740_5135, \8810_9109 );
and \U$6106 ( \14915_15214 , RIee3a660_5123, \8812_9111 );
and \U$6107 ( \14916_15215 , RIe174e28_2707, \8814_9113 );
and \U$6108 ( \14917_15216 , RIf170768_5739, \8816_9115 );
and \U$6109 ( \14918_15217 , RIfc5fdf8_6113, \8818_9117 );
and \U$6110 ( \14919_15218 , RIf16eb48_5719, \8820_9119 );
and \U$6111 ( \14920_15219 , RIfcaaab0_6964, \8822_9121 );
and \U$6112 ( \14921_15220 , RIf16d1f8_5701, \8824_9123 );
and \U$6113 ( \14922_15221 , RIe225318_4713, \8826_9125 );
and \U$6114 ( \14923_15222 , RIf16c6b8_5693, \8828_9127 );
and \U$6115 ( \14924_15223 , RIe222618_4681, \8830_9129 );
and \U$6116 ( \14925_15224 , RIf16b5d8_5681, \8832_9131 );
and \U$6117 ( \14926_15225 , RIe21f918_4649, \8834_9133 );
and \U$6118 ( \14927_15226 , RIe219f18_4585, \8836_9135 );
and \U$6119 ( \14928_15227 , RIe217218_4553, \8838_9137 );
and \U$6120 ( \14929_15228 , RIfca62f8_6913, \8840_9139 );
and \U$6121 ( \14930_15229 , RIe214518_4521, \8842_9141 );
and \U$6122 ( \14931_15230 , RIfcc9578_7313, \8844_9143 );
and \U$6123 ( \14932_15231 , RIe211818_4489, \8846_9145 );
and \U$6124 ( \14933_15232 , RIfca5a88_6907, \8848_9147 );
and \U$6125 ( \14934_15233 , RIe20eb18_4457, \8850_9149 );
and \U$6126 ( \14935_15234 , RIe20be18_4425, \8852_9151 );
and \U$6127 ( \14936_15235 , RIe209118_4393, \8854_9153 );
and \U$6128 ( \14937_15236 , RIf167690_5636, \8856_9155 );
and \U$6129 ( \14938_15237 , RIf166718_5625, \8858_9157 );
and \U$6130 ( \14939_15238 , RIfe8f9a0_7978, \8860_9159 );
and \U$6131 ( \14940_15239 , RIfe8f838_7977, \8862_9161 );
and \U$6132 ( \14941_15240 , RIf165638_5613, \8864_9163 );
and \U$6133 ( \14942_15241 , RIf164990_5604, \8866_9165 );
and \U$6134 ( \14943_15242 , RIf1638b0_5592, \8868_9167 );
and \U$6135 ( \14944_15243 , RIf1627d0_5580, \8870_9169 );
and \U$6136 ( \14945_15244 , RIf161150_5564, \8872_9171 );
and \U$6137 ( \14946_15245 , RIf15f260_5542, \8874_9173 );
and \U$6138 ( \14947_15246 , RIe1fd778_4261, \8876_9175 );
and \U$6139 ( \14948_15247 , RIe1fc530_4248, \8878_9177 );
and \U$6140 ( \14949_15248 , RIf15d4d8_5521, \8880_9179 );
and \U$6141 ( \14950_15249 , RIf15c290_5508, \8882_9181 );
and \U$6142 ( \14951_15250 , RIfca20e0_6866, \8884_9183 );
and \U$6143 ( \14952_15251 , RIf159f68_5483, \8886_9185 );
or \U$6144 ( \14953_15252 , \14889_15188 , \14890_15189 , \14891_15190 , \14892_15191 , \14893_15192 , \14894_15193 , \14895_15194 , \14896_15195 , \14897_15196 , \14898_15197 , \14899_15198 , \14900_15199 , \14901_15200 , \14902_15201 , \14903_15202 , \14904_15203 , \14905_15204 , \14906_15205 , \14907_15206 , \14908_15207 , \14909_15208 , \14910_15209 , \14911_15210 , \14912_15211 , \14913_15212 , \14914_15213 , \14915_15214 , \14916_15215 , \14917_15216 , \14918_15217 , \14919_15218 , \14920_15219 , \14921_15220 , \14922_15221 , \14923_15222 , \14924_15223 , \14925_15224 , \14926_15225 , \14927_15226 , \14928_15227 , \14929_15228 , \14930_15229 , \14931_15230 , \14932_15231 , \14933_15232 , \14934_15233 , \14935_15234 , \14936_15235 , \14937_15236 , \14938_15237 , \14939_15238 , \14940_15239 , \14941_15240 , \14942_15241 , \14943_15242 , \14944_15243 , \14945_15244 , \14946_15245 , \14947_15246 , \14948_15247 , \14949_15248 , \14950_15249 , \14951_15250 , \14952_15251 );
and \U$6145 ( \14954_15253 , RIf159428_5475, \8889_9188 );
and \U$6146 ( \14955_15254 , RIf1581e0_5462, \8891_9190 );
and \U$6147 ( \14956_15255 , RIfc5ebb0_6100, \8893_9192 );
and \U$6148 ( \14957_15256 , RIfe8fdd8_7981, \8895_9194 );
and \U$6149 ( \14958_15257 , RIfc69e48_6227, \8897_9196 );
and \U$6150 ( \14959_15258 , RIfc5e8e0_6098, \8899_9198 );
and \U$6151 ( \14960_15259 , RIf154f40_5426, \8901_9200 );
and \U$6152 ( \14961_15260 , RIe1f6b30_4184, \8903_9202 );
and \U$6153 ( \14962_15261 , RIf153b90_5412, \8905_9204 );
and \U$6154 ( \14963_15262 , RIf1523a8_5395, \8907_9206 );
and \U$6155 ( \14964_15263 , RIfce88b0_7668, \8909_9208 );
and \U$6156 ( \14965_15264 , RIfe8fb08_7979, \8911_9210 );
and \U$6157 ( \14966_15265 , RIfcebe20_7706, \8913_9212 );
and \U$6158 ( \14967_15266 , RIfcb1158_7037, \8915_9214 );
and \U$6159 ( \14968_15267 , RIf14e730_5352, \8917_9216 );
and \U$6160 ( \14969_15268 , RIe1ef678_4101, \8919_9218 );
and \U$6161 ( \14970_15269 , RIe1ed080_4074, \8921_9220 );
and \U$6162 ( \14971_15270 , RIe1ea380_4042, \8923_9222 );
and \U$6163 ( \14972_15271 , RIe1e7680_4010, \8925_9224 );
and \U$6164 ( \14973_15272 , RIe1e4980_3978, \8927_9226 );
and \U$6165 ( \14974_15273 , RIe1e1c80_3946, \8929_9228 );
and \U$6166 ( \14975_15274 , RIe1def80_3914, \8931_9230 );
and \U$6167 ( \14976_15275 , RIe1dc280_3882, \8933_9232 );
and \U$6168 ( \14977_15276 , RIe1d9580_3850, \8935_9234 );
and \U$6169 ( \14978_15277 , RIe1d3b80_3786, \8937_9236 );
and \U$6170 ( \14979_15278 , RIe1d0e80_3754, \8939_9238 );
and \U$6171 ( \14980_15279 , RIe1ce180_3722, \8941_9240 );
and \U$6172 ( \14981_15280 , RIe1cb480_3690, \8943_9242 );
and \U$6173 ( \14982_15281 , RIe1c8780_3658, \8945_9244 );
and \U$6174 ( \14983_15282 , RIe1c5a80_3626, \8947_9246 );
and \U$6175 ( \14984_15283 , RIe1c2d80_3594, \8949_9248 );
and \U$6176 ( \14985_15284 , RIe1c0080_3562, \8951_9250 );
and \U$6177 ( \14986_15285 , RIfcc8ba0_7306, \8953_9252 );
and \U$6178 ( \14987_15286 , RIfc5d698_6085, \8955_9254 );
and \U$6179 ( \14988_15287 , RIfec35e8_8343, \8957_9256 );
and \U$6180 ( \14989_15288 , RIfeabd08_8271, \8959_9258 );
and \U$6181 ( \14990_15289 , RIfc5cf90_6080, \8961_9260 );
and \U$6182 ( \14991_15290 , RIfc5ce28_6079, \8963_9262 );
and \U$6183 ( \14992_15291 , RIfec31b0_8340, \8965_9264 );
and \U$6184 ( \14993_15292 , RIe1b4b18_3433, \8967_9266 );
and \U$6185 ( \14994_15293 , RIf149708_5295, \8969_9268 );
and \U$6186 ( \14995_15294 , RIf148358_5281, \8971_9270 );
and \U$6187 ( \14996_15295 , RIe1b3768_3419, \8973_9272 );
and \U$6188 ( \14997_15296 , RIfec3480_8342, \8975_9274 );
and \U$6189 ( \14998_15297 , RIfc483b0_5844, \8977_9276 );
and \U$6190 ( \14999_15298 , RIfc80be8_6487, \8979_9278 );
and \U$6191 ( \15000_15299 , RIe1ad4f8_3349, \8981_9280 );
and \U$6192 ( \15001_15300 , RIfec3318_8341, \8983_9282 );
and \U$6193 ( \15002_15301 , RIe1aa3c0_3314, \8985_9284 );
and \U$6194 ( \15003_15302 , RIe1a76c0_3282, \8987_9286 );
and \U$6195 ( \15004_15303 , RIe1a49c0_3250, \8989_9288 );
and \U$6196 ( \15005_15304 , RIe1a1cc0_3218, \8991_9290 );
and \U$6197 ( \15006_15305 , RIe18e1c0_2994, \8993_9292 );
and \U$6198 ( \15007_15306 , RIe17a6c0_2770, \8995_9294 );
and \U$6199 ( \15008_15307 , RIe228018_4745, \8997_9296 );
and \U$6200 ( \15009_15308 , RIe21cc18_4617, \8999_9298 );
and \U$6201 ( \15010_15309 , RIe206418_4361, \9001_9300 );
and \U$6202 ( \15011_15310 , RIe200478_4293, \9003_9302 );
and \U$6203 ( \15012_15311 , RIe1f9830_4216, \9005_9304 );
and \U$6204 ( \15013_15312 , RIe1f2378_4133, \9007_9306 );
and \U$6205 ( \15014_15313 , RIe1d6880_3818, \9009_9308 );
and \U$6206 ( \15015_15314 , RIe1bd380_3530, \9011_9310 );
and \U$6207 ( \15016_15315 , RIe1b01f8_3381, \9013_9312 );
and \U$6208 ( \15017_15316 , RIe172830_2680, \9015_9314 );
or \U$6209 ( \15018_15317 , \14954_15253 , \14955_15254 , \14956_15255 , \14957_15256 , \14958_15257 , \14959_15258 , \14960_15259 , \14961_15260 , \14962_15261 , \14963_15262 , \14964_15263 , \14965_15264 , \14966_15265 , \14967_15266 , \14968_15267 , \14969_15268 , \14970_15269 , \14971_15270 , \14972_15271 , \14973_15272 , \14974_15273 , \14975_15274 , \14976_15275 , \14977_15276 , \14978_15277 , \14979_15278 , \14980_15279 , \14981_15280 , \14982_15281 , \14983_15282 , \14984_15283 , \14985_15284 , \14986_15285 , \14987_15286 , \14988_15287 , \14989_15288 , \14990_15289 , \14991_15290 , \14992_15291 , \14993_15292 , \14994_15293 , \14995_15294 , \14996_15295 , \14997_15296 , \14998_15297 , \14999_15298 , \15000_15299 , \15001_15300 , \15002_15301 , \15003_15302 , \15004_15303 , \15005_15304 , \15006_15305 , \15007_15306 , \15008_15307 , \15009_15308 , \15010_15309 , \15011_15310 , \15012_15311 , \15013_15312 , \15014_15313 , \15015_15314 , \15016_15315 , \15017_15316 );
or \U$6210 ( \15019_15318 , \14953_15252 , \15018_15317 );
_DC \g6593/U$1 ( \15020 , \15019_15318 , \9024_9323 );
and g6594_GF_PartitionCandidate( \15021_15320_nG6594 , \14888 , \15020 );
buf \U$6211 ( \15022_15321 , \15021_15320_nG6594 );
and \U$6212 ( \15023_15322 , \15022_15321 , \10389_10691 );
nor \U$6213 ( \15024_15323 , \14756_15055 , \15023_15322 );
xnor \U$6214 ( \15025_15324 , \15024_15323 , \10678_10980 );
and \U$6215 ( \15026_15325 , \10968_11270 , \13755_14054 );
and \U$6216 ( \15027_15326 , \11287_11586 , \13390_13692 );
nor \U$6217 ( \15028_15327 , \15026_15325 , \15027_15326 );
xnor \U$6218 ( \15029_15328 , \15028_15327 , \13736_14035 );
xor \U$6219 ( \15030_15329 , \15025_15324 , \15029_15328 );
_DC \g4e2b/U$1 ( \15031 , \14887_15186 , \9298_9597 );
_DC \g4eaf/U$1 ( \15032 , \15019_15318 , \9024_9323 );
xor g4eb0_GF_PartitionCandidate( \15033_15332_nG4eb0 , \15031 , \15032 );
buf \U$6220 ( \15034_15333 , \15033_15332_nG4eb0 );
xor \U$6221 ( \15035_15334 , \15034_15333 , \14660_14962 );
not \U$6222 ( \15036_15335 , \14661_14963 );
and \U$6223 ( \15037_15336 , \15035_15334 , \15036_15335 );
and \U$6224 ( \15038_15337 , \10385_10687 , \15037_15336 );
and \U$6225 ( \15039_15338 , \10686_10988 , \14661_14963 );
nor \U$6226 ( \15040_15339 , \15038_15337 , \15039_15338 );
and \U$6227 ( \15041_15340 , \14660_14962 , \13733_14032 );
not \U$6228 ( \15042_15341 , \15041_15340 );
and \U$6229 ( \15043_15342 , \15034_15333 , \15042_15341 );
xnor \U$6230 ( \15044_15343 , \15040_15339 , \15043_15342 );
xor \U$6231 ( \15045_15344 , \15030_15329 , \15044_15343 );
xor \U$6232 ( \15046_15345 , \14755_15054 , \15045_15344 );
and \U$6233 ( \15047_15346 , \13377_13679 , \11275_11574 );
and \U$6234 ( \15048_15347 , \13725_14024 , \10976_11278 );
nor \U$6235 ( \15049_15348 , \15047_15346 , \15048_15347 );
xnor \U$6236 ( \15050_15349 , \15049_15348 , \11281_11580 );
not \U$6237 ( \15051_15350 , \14662_14964 );
and \U$6238 ( \15052_15351 , \15051_15350 , \15043_15342 );
xor \U$6239 ( \15053_15352 , \15050_15349 , \15052_15351 );
and \U$6240 ( \15054_15353 , \14651_14953 , \14655_14957 );
and \U$6241 ( \15055_15354 , \14655_14957 , \14662_14964 );
and \U$6242 ( \15056_15355 , \14651_14953 , \14662_14964 );
or \U$6243 ( \15057_15356 , \15054_15353 , \15055_15354 , \15056_15355 );
xor \U$6244 ( \15058_15357 , \15053_15352 , \15057_15356 );
and \U$6245 ( \15059_15358 , \12146_12448 , \12491_12790 );
and \U$6246 ( \15060_15359 , \12470_12769 , \12159_12461 );
nor \U$6247 ( \15061_15360 , \15059_15358 , \15060_15359 );
xnor \U$6248 ( \15062_15361 , \15061_15360 , \12481_12780 );
xor \U$6249 ( \15063_15362 , \15058_15357 , \15062_15361 );
xor \U$6250 ( \15064_15363 , \15046_15345 , \15063_15362 );
and \U$6251 ( \15065_15364 , \14381_14683 , \14663_14965 );
and \U$6252 ( \15066_15365 , \14663_14965 , \14675_14977 );
and \U$6253 ( \15067_15366 , \14381_14683 , \14675_14977 );
or \U$6254 ( \15068_15367 , \15065_15364 , \15066_15365 , \15067_15366 );
xor \U$6255 ( \15069_15368 , \15064_15363 , \15068_15367 );
and \U$6256 ( \15070_15369 , \14377_14679 , \14676_14978 );
and \U$6257 ( \15071_15370 , \14677_14979 , \14680_14982 );
or \U$6258 ( \15072_15371 , \15070_15369 , \15071_15370 );
xor \U$6259 ( \15073_15372 , \15069_15368 , \15072_15371 );
buf g9bf3_GF_PartitionCandidate( \15074_15373_nG9bf3 , \15073_15372 );
and \U$6260 ( \15075_15374 , \10402_10704 , \15074_15373_nG9bf3 );
or \U$6261 ( \15076_15375 , \14751_15050 , \15075_15374 );
xor \U$6262 ( \15077_15376 , \10399_10703 , \15076_15375 );
buf \U$6263 ( \15078_15377 , \15077_15376 );
buf \U$6265 ( \15079_15378 , \15078_15377 );
xor \U$6266 ( \15080_15379 , \14750_15049 , \15079_15378 );
buf \U$6267 ( \15081_15380 , \15080_15379 );
xor \U$6268 ( \15082_15381 , \14704_15006 , \15081_15380 );
and \U$6269 ( \15083_15382 , \14341_14643 , \14689_14991 );
and \U$6270 ( \15084_15383 , \14341_14643 , \14695_14997 );
and \U$6271 ( \15085_15384 , \14689_14991 , \14695_14997 );
or \U$6272 ( \15086_15385 , \15083_15382 , \15084_15383 , \15085_15384 );
buf \U$6273 ( \15087_15386 , \15086_15385 );
xor \U$6274 ( \15088_15387 , \15082_15381 , \15087_15386 );
and \U$6275 ( \15089_15388 , \14699_15001 , \15088_15387 );
and \U$6276 ( \15090_15389 , RIdec4460_697, \8760_9059 );
and \U$6277 ( \15091_15390 , RIdec1760_665, \8762_9061 );
and \U$6278 ( \15092_15391 , RIee1fae0_4819, \8764_9063 );
and \U$6279 ( \15093_15392 , RIdebea60_633, \8766_9065 );
and \U$6280 ( \15094_15393 , RIee1f108_4812, \8768_9067 );
and \U$6281 ( \15095_15394 , RIdebbd60_601, \8770_9069 );
and \U$6282 ( \15096_15395 , RIdeb9060_569, \8772_9071 );
and \U$6283 ( \15097_15396 , RIdeb6360_537, \8774_9073 );
and \U$6284 ( \15098_15397 , RIee1eb68_4808, \8776_9075 );
and \U$6285 ( \15099_15398 , RIdeb0960_473, \8778_9077 );
and \U$6286 ( \15100_15399 , RIee1e460_4803, \8780_9079 );
and \U$6287 ( \15101_15400 , RIdeadc60_441, \8782_9081 );
and \U$6288 ( \15102_15401 , RIee1d7b8_4794, \8784_9083 );
and \U$6289 ( \15103_15402 , RIdea8008_409, \8786_9085 );
and \U$6290 ( \15104_15403 , RIdea1708_377, \8788_9087 );
and \U$6291 ( \15105_15404 , RIde9ae08_345, \8790_9089 );
and \U$6292 ( \15106_15405 , RIfe957d8_8045, \8792_9091 );
and \U$6293 ( \15107_15406 , RIfe95508_8043, \8794_9093 );
and \U$6294 ( \15108_15407 , RIfe95670_8044, \8796_9095 );
and \U$6295 ( \15109_15408 , RIee1a7e8_4760, \8798_9097 );
and \U$6296 ( \15110_15409 , RIfe95aa8_8047, \8800_9099 );
and \U$6297 ( \15111_15410 , RIfe95238_8041, \8802_9101 );
and \U$6298 ( \15112_15411 , RIfe95940_8046, \8804_9103 );
and \U$6299 ( \15113_15412 , RIfe953a0_8042, \8806_9105 );
and \U$6300 ( \15114_15413 , RIee1a0e0_4755, \8808_9107 );
and \U$6301 ( \15115_15414 , RIee19ca8_4752, \8810_9109 );
and \U$6302 ( \15116_15415 , RIee19870_4749, \8812_9111 );
and \U$6303 ( \15117_15416 , RIee19438_4746, \8814_9113 );
and \U$6304 ( \15118_15417 , RIee38ba8_5104, \8816_9115 );
and \U$6305 ( \15119_15418 , RIfe95c10_8048, \8818_9117 );
and \U$6306 ( \15120_15419 , RIee384a0_5099, \8820_9119 );
and \U$6307 ( \15121_15420 , RIfea9440_8242, \8822_9121 );
and \U$6308 ( \15122_15421 , RIe164460_2518, \8824_9123 );
and \U$6309 ( \15123_15422 , RIe161760_2486, \8826_9125 );
and \U$6310 ( \15124_15423 , RIfe942c0_8030, \8828_9127 );
and \U$6311 ( \15125_15424 , RIe15ea60_2454, \8830_9129 );
and \U$6312 ( \15126_15425 , RIfe94158_8029, \8832_9131 );
and \U$6313 ( \15127_15426 , RIe15bd60_2422, \8834_9133 );
and \U$6314 ( \15128_15427 , RIe156360_2358, \8836_9135 );
and \U$6315 ( \15129_15428 , RIe153660_2326, \8838_9137 );
and \U$6316 ( \15130_15429 , RIfe94428_8031, \8840_9139 );
and \U$6317 ( \15131_15430 , RIe150960_2294, \8842_9141 );
and \U$6318 ( \15132_15431 , RIfe94590_8032, \8844_9143 );
and \U$6319 ( \15133_15432 , RIe14dc60_2262, \8846_9145 );
and \U$6320 ( \15134_15433 , RIfc5c2e8_6071, \8848_9147 );
and \U$6321 ( \15135_15434 , RIe14af60_2230, \8850_9149 );
and \U$6322 ( \15136_15435 , RIe148260_2198, \8852_9151 );
and \U$6323 ( \15137_15436 , RIe145560_2166, \8854_9153 );
and \U$6324 ( \15138_15437 , RIee33ce8_5048, \8856_9155 );
and \U$6325 ( \15139_15438 , RIee32aa0_5035, \8858_9157 );
and \U$6326 ( \15140_15439 , RIee31858_5022, \8860_9159 );
and \U$6327 ( \15141_15440 , RIfc5d530_6084, \8862_9161 );
and \U$6328 ( \15142_15441 , RIe140538_2109, \8864_9163 );
and \U$6329 ( \15143_15442 , RIdf3e2d8_2084, \8866_9165 );
and \U$6330 ( \15144_15443 , RIdf3c118_2060, \8868_9167 );
and \U$6331 ( \15145_15444 , RIdf39df0_2035, \8870_9169 );
and \U$6332 ( \15146_15445 , RIfcdd780_7542, \8872_9171 );
and \U$6333 ( \15147_15446 , RIee2ee28_4992, \8874_9173 );
and \U$6334 ( \15148_15447 , RIfcc88d0_7304, \8876_9175 );
and \U$6335 ( \15149_15448 , RIee2cc68_4968, \8878_9177 );
and \U$6336 ( \15150_15449 , RIdf34990_1975, \8880_9179 );
and \U$6337 ( \15151_15450 , RIdf32aa0_1953, \8882_9181 );
and \U$6338 ( \15152_15451 , RIdf304a8_1926, \8884_9183 );
and \U$6339 ( \15153_15452 , RIdf2e5b8_1904, \8886_9185 );
or \U$6340 ( \15154_15453 , \15090_15389 , \15091_15390 , \15092_15391 , \15093_15392 , \15094_15393 , \15095_15394 , \15096_15395 , \15097_15396 , \15098_15397 , \15099_15398 , \15100_15399 , \15101_15400 , \15102_15401 , \15103_15402 , \15104_15403 , \15105_15404 , \15106_15405 , \15107_15406 , \15108_15407 , \15109_15408 , \15110_15409 , \15111_15410 , \15112_15411 , \15113_15412 , \15114_15413 , \15115_15414 , \15116_15415 , \15117_15416 , \15118_15417 , \15119_15418 , \15120_15419 , \15121_15420 , \15122_15421 , \15123_15422 , \15124_15423 , \15125_15424 , \15126_15425 , \15127_15426 , \15128_15427 , \15129_15428 , \15130_15429 , \15131_15430 , \15132_15431 , \15133_15432 , \15134_15433 , \15135_15434 , \15136_15435 , \15137_15436 , \15138_15437 , \15139_15438 , \15140_15439 , \15141_15440 , \15142_15441 , \15143_15442 , \15144_15443 , \15145_15444 , \15146_15445 , \15147_15446 , \15148_15447 , \15149_15448 , \15150_15449 , \15151_15450 , \15152_15451 , \15153_15452 );
and \U$6341 ( \15155_15454 , RIee2b1b0_4949, \8889_9188 );
and \U$6342 ( \15156_15455 , RIfe946f8_8033, \8891_9190 );
and \U$6343 ( \15157_15456 , RIfcb2940_7054, \8893_9192 );
and \U$6344 ( \15158_15457 , RIee273d0_4905, \8895_9194 );
and \U$6345 ( \15159_15458 , RIfe949c8_8035, \8897_9196 );
and \U$6346 ( \15160_15459 , RIdf27538_1824, \8899_9198 );
and \U$6347 ( \15161_15460 , RIfe94b30_8036, \8901_9200 );
and \U$6348 ( \15162_15461 , RIfe94860_8034, \8903_9202 );
and \U$6349 ( \15163_15462 , RIee26f98_4902, \8905_9204 );
and \U$6350 ( \15164_15463 , RIee269f8_4898, \8907_9206 );
and \U$6351 ( \15165_15464 , RIee26728_4896, \8909_9208 );
and \U$6352 ( \15166_15465 , RIee26458_4894, \8911_9210 );
and \U$6353 ( \15167_15466 , RIee26188_4892, \8913_9212 );
and \U$6354 ( \15168_15467 , RIfe94c98_8037, \8915_9214 );
and \U$6355 ( \15169_15468 , RIee25d50_4889, \8917_9216 );
and \U$6356 ( \15170_15469 , RIfea9170_8240, \8919_9218 );
and \U$6357 ( \15171_15470 , RIdf16030_1627, \8921_9220 );
and \U$6358 ( \15172_15471 , RIdf13330_1595, \8923_9222 );
and \U$6359 ( \15173_15472 , RIdf10630_1563, \8925_9224 );
and \U$6360 ( \15174_15473 , RIdf0d930_1531, \8927_9226 );
and \U$6361 ( \15175_15474 , RIdf0ac30_1499, \8929_9228 );
and \U$6362 ( \15176_15475 , RIdf07f30_1467, \8931_9230 );
and \U$6363 ( \15177_15476 , RIdf05230_1435, \8933_9232 );
and \U$6364 ( \15178_15477 , RIdf02530_1403, \8935_9234 );
and \U$6365 ( \15179_15478 , RIdefcb30_1339, \8937_9236 );
and \U$6366 ( \15180_15479 , RIdef9e30_1307, \8939_9238 );
and \U$6367 ( \15181_15480 , RIdef7130_1275, \8941_9240 );
and \U$6368 ( \15182_15481 , RIdef4430_1243, \8943_9242 );
and \U$6369 ( \15183_15482 , RIdef1730_1211, \8945_9244 );
and \U$6370 ( \15184_15483 , RIdeeea30_1179, \8947_9246 );
and \U$6371 ( \15185_15484 , RIdeebd30_1147, \8949_9248 );
and \U$6372 ( \15186_15485 , RIdee9030_1115, \8951_9250 );
and \U$6373 ( \15187_15486 , RIee250a8_4880, \8953_9252 );
and \U$6374 ( \15188_15487 , RIee24298_4870, \8955_9254 );
and \U$6375 ( \15189_15488 , RIee23758_4862, \8957_9256 );
and \U$6376 ( \15190_15489 , RIee22d80_4855, \8959_9258 );
and \U$6377 ( \15191_15490 , RIfe950d0_8040, \8961_9260 );
and \U$6378 ( \15192_15491 , RIfe94f68_8039, \8963_9262 );
and \U$6379 ( \15193_15492 , RIfe94e00_8038, \8965_9264 );
and \U$6380 ( \15194_15493 , RIdeddd98_988, \8967_9266 );
and \U$6381 ( \15195_15494 , RIee22ab0_4853, \8969_9268 );
and \U$6382 ( \15196_15495 , RIee21e08_4844, \8971_9270 );
and \U$6383 ( \15197_15496 , RIfca46d8_6893, \8973_9272 );
and \U$6384 ( \15198_15497 , RIfc5dad0_6088, \8975_9274 );
and \U$6385 ( \15199_15498 , RIfeaa250_8252, \8977_9276 );
and \U$6386 ( \15200_15499 , RIfe96048_8051, \8979_9278 );
and \U$6387 ( \15201_15500 , RIfe95d78_8049, \8981_9280 );
and \U$6388 ( \15202_15501 , RIfe95ee0_8050, \8983_9282 );
and \U$6389 ( \15203_15502 , RIdecf860_825, \8985_9284 );
and \U$6390 ( \15204_15503 , RIdeccb60_793, \8987_9286 );
and \U$6391 ( \15205_15504 , RIdec9e60_761, \8989_9288 );
and \U$6392 ( \15206_15505 , RIdec7160_729, \8991_9290 );
and \U$6393 ( \15207_15506 , RIdeb3660_505, \8993_9292 );
and \U$6394 ( \15208_15507 , RIde94508_313, \8995_9294 );
and \U$6395 ( \15209_15508 , RIe16d268_2619, \8997_9296 );
and \U$6396 ( \15210_15509 , RIe159060_2390, \8999_9298 );
and \U$6397 ( \15211_15510 , RIe142860_2134, \9001_9300 );
and \U$6398 ( \15212_15511 , RIdf37258_2004, \9003_9302 );
and \U$6399 ( \15213_15512 , RIdf2b8b8_1872, \9005_9304 );
and \U$6400 ( \15214_15513 , RIdf1c138_1696, \9007_9306 );
and \U$6401 ( \15215_15514 , RIdeff830_1371, \9009_9308 );
and \U$6402 ( \15216_15515 , RIdee6330_1083, \9011_9310 );
and \U$6403 ( \15217_15516 , RIdedb098_956, \9013_9312 );
and \U$6404 ( \15218_15517 , RIde7a450_186, \9015_9314 );
or \U$6405 ( \15219_15518 , \15155_15454 , \15156_15455 , \15157_15456 , \15158_15457 , \15159_15458 , \15160_15459 , \15161_15460 , \15162_15461 , \15163_15462 , \15164_15463 , \15165_15464 , \15166_15465 , \15167_15466 , \15168_15467 , \15169_15468 , \15170_15469 , \15171_15470 , \15172_15471 , \15173_15472 , \15174_15473 , \15175_15474 , \15176_15475 , \15177_15476 , \15178_15477 , \15179_15478 , \15180_15479 , \15181_15480 , \15182_15481 , \15183_15482 , \15184_15483 , \15185_15484 , \15186_15485 , \15187_15486 , \15188_15487 , \15189_15488 , \15190_15489 , \15191_15490 , \15192_15491 , \15193_15492 , \15194_15493 , \15195_15494 , \15196_15495 , \15197_15496 , \15198_15497 , \15199_15498 , \15200_15499 , \15201_15500 , \15202_15501 , \15203_15502 , \15204_15503 , \15205_15504 , \15206_15505 , \15207_15506 , \15208_15507 , \15209_15508 , \15210_15509 , \15211_15510 , \15212_15511 , \15213_15512 , \15214_15513 , \15215_15514 , \15216_15515 , \15217_15516 , \15218_15517 );
or \U$6406 ( \15220_15519 , \15154_15453 , \15219_15518 );
_DC \g2c99/U$1 ( \15221 , \15220_15519 , \9024_9323 );
buf \U$6407 ( \15222_15521 , \15221 );
and \U$6408 ( \15223_15522 , RIe19c6f8_3157, \9034_9333 );
and \U$6409 ( \15224_15523 , RIe1999f8_3125, \9036_9335 );
and \U$6410 ( \15225_15524 , RIf1450b8_5245, \9038_9337 );
and \U$6411 ( \15226_15525 , RIe196cf8_3093, \9040_9339 );
and \U$6412 ( \15227_15526 , RIf143fd8_5233, \9042_9341 );
and \U$6413 ( \15228_15527 , RIe193ff8_3061, \9044_9343 );
and \U$6414 ( \15229_15528 , RIe1912f8_3029, \9046_9345 );
and \U$6415 ( \15230_15529 , RIe18e5f8_2997, \9048_9347 );
and \U$6416 ( \15231_15530 , RIe188bf8_2933, \9050_9349 );
and \U$6417 ( \15232_15531 , RIe185ef8_2901, \9052_9351 );
and \U$6418 ( \15233_15532 , RIfe973f8_8065, \9054_9353 );
and \U$6419 ( \15234_15533 , RIe1831f8_2869, \9056_9355 );
and \U$6420 ( \15235_15534 , RIf142958_5217, \9058_9357 );
and \U$6421 ( \15236_15535 , RIe1804f8_2837, \9060_9359 );
and \U$6422 ( \15237_15536 , RIe17d7f8_2805, \9062_9361 );
and \U$6423 ( \15238_15537 , RIe17aaf8_2773, \9064_9363 );
and \U$6424 ( \15239_15538 , RIf141b48_5207, \9066_9365 );
and \U$6425 ( \15240_15539 , RIfc542f0_5980, \9068_9367 );
and \U$6426 ( \15241_15540 , RIfc800a8_6479, \9070_9369 );
and \U$6427 ( \15242_15541 , RIe175260_2710, \9072_9371 );
and \U$6428 ( \15243_15542 , RIfca0bc8_6851, \9074_9373 );
and \U$6429 ( \15244_15543 , RIfc48680_5846, \9076_9375 );
and \U$6430 ( \15245_15544 , RIee3dea0_5163, \9078_9377 );
and \U$6431 ( \15246_15545 , RIfcc6878_7281, \9080_9379 );
and \U$6432 ( \15247_15546 , RIee3ba10_5137, \9082_9381 );
and \U$6433 ( \15248_15547 , RIee3a930_5125, \9084_9383 );
and \U$6434 ( \15249_15548 , RIfe97290_8064, \9086_9385 );
and \U$6435 ( \15250_15549 , RIe172b00_2682, \9088_9387 );
and \U$6436 ( \15251_15550 , RIf16f958_5729, \9090_9389 );
and \U$6437 ( \15252_15551 , RIf16ee18_5721, \9092_9391 );
and \U$6438 ( \15253_15552 , RIf16da68_5707, \9094_9393 );
and \U$6439 ( \15254_15553 , RIf16d360_5702, \9096_9395 );
and \U$6440 ( \15255_15554 , RIfe96e58_8061, \9098_9397 );
and \U$6441 ( \15256_15555 , RIe222a50_4684, \9100_9399 );
and \U$6442 ( \15257_15556 , RIfe96cf0_8060, \9102_9401 );
and \U$6443 ( \15258_15557 , RIe21fd50_4652, \9104_9403 );
and \U$6444 ( \15259_15558 , RIf16a660_5670, \9106_9405 );
and \U$6445 ( \15260_15559 , RIe21d050_4620, \9108_9407 );
and \U$6446 ( \15261_15560 , RIe217650_4556, \9110_9409 );
and \U$6447 ( \15262_15561 , RIe214950_4524, \9112_9411 );
and \U$6448 ( \15263_15562 , RIf169f58_5665, \9114_9413 );
and \U$6449 ( \15264_15563 , RIe211c50_4492, \9116_9415 );
and \U$6450 ( \15265_15564 , RIf168770_5648, \9118_9417 );
and \U$6451 ( \15266_15565 , RIe20ef50_4460, \9120_9419 );
and \U$6452 ( \15267_15566 , RIf1677f8_5637, \9122_9421 );
and \U$6453 ( \15268_15567 , RIe20c250_4428, \9124_9423 );
and \U$6454 ( \15269_15568 , RIe209550_4396, \9126_9425 );
and \U$6455 ( \15270_15569 , RIe206850_4364, \9128_9427 );
and \U$6456 ( \15271_15570 , RIf166880_5626, \9130_9429 );
and \U$6457 ( \15272_15571 , RIf1657a0_5614, \9132_9431 );
and \U$6458 ( \15273_15572 , RIe201dc8_4311, \9134_9433 );
and \U$6459 ( \15274_15573 , RIe2005e0_4294, \9136_9435 );
and \U$6460 ( \15275_15574 , RIfe96b88_8059, \9138_9437 );
and \U$6461 ( \15276_15575 , RIf163b80_5594, \9140_9439 );
and \U$6462 ( \15277_15576 , RIf162c08_5583, \9142_9441 );
and \U$6463 ( \15278_15577 , RIf161420_5566, \9144_9443 );
and \U$6464 ( \15279_15578 , RIf15f530_5544, \9146_9445 );
and \U$6465 ( \15280_15579 , RIf15d7a8_5523, \9148_9447 );
and \U$6466 ( \15281_15580 , RIfe968b8_8057, \9150_9449 );
and \U$6467 ( \15282_15581 , RIfe96a20_8058, \9152_9451 );
and \U$6468 ( \15283_15582 , RIfcb3fc0_7070, \9154_9453 );
and \U$6469 ( \15284_15583 , RIfc7cf70_6444, \9156_9455 );
and \U$6470 ( \15285_15584 , RIfc579c8_6019, \9158_9457 );
and \U$6471 ( \15286_15585 , RIf159590_5476, \9160_9459 );
or \U$6472 ( \15287_15586 , \15223_15522 , \15224_15523 , \15225_15524 , \15226_15525 , \15227_15526 , \15228_15527 , \15229_15528 , \15230_15529 , \15231_15530 , \15232_15531 , \15233_15532 , \15234_15533 , \15235_15534 , \15236_15535 , \15237_15536 , \15238_15537 , \15239_15538 , \15240_15539 , \15241_15540 , \15242_15541 , \15243_15542 , \15244_15543 , \15245_15544 , \15246_15545 , \15247_15546 , \15248_15547 , \15249_15548 , \15250_15549 , \15251_15550 , \15252_15551 , \15253_15552 , \15254_15553 , \15255_15554 , \15256_15555 , \15257_15556 , \15258_15557 , \15259_15558 , \15260_15559 , \15261_15560 , \15262_15561 , \15263_15562 , \15264_15563 , \15265_15564 , \15266_15565 , \15267_15566 , \15268_15567 , \15269_15568 , \15270_15569 , \15271_15570 , \15272_15571 , \15273_15572 , \15274_15573 , \15275_15574 , \15276_15575 , \15277_15576 , \15278_15577 , \15279_15578 , \15280_15579 , \15281_15580 , \15282_15581 , \15283_15582 , \15284_15583 , \15285_15584 , \15286_15585 );
and \U$6473 ( \15288_15587 , RIf1584b0_5464, \9163_9462 );
and \U$6474 ( \15289_15588 , RIf157268_5451, \9165_9464 );
and \U$6475 ( \15290_15589 , RIf1569f8_5445, \9167_9466 );
and \U$6476 ( \15291_15590 , RIfe965e8_8055, \9169_9468 );
and \U$6477 ( \15292_15591 , RIf155d50_5436, \9171_9470 );
and \U$6478 ( \15293_15592 , RIf155210_5428, \9173_9472 );
and \U$6479 ( \15294_15593 , RIf153e60_5414, \9175_9474 );
and \U$6480 ( \15295_15594 , RIfe96750_8056, \9177_9476 );
and \U$6481 ( \15296_15595 , RIf1527e0_5398, \9179_9478 );
and \U$6482 ( \15297_15596 , RIf151430_5384, \9181_9480 );
and \U$6483 ( \15298_15597 , RIfcd2650_7416, \9183_9482 );
and \U$6484 ( \15299_15598 , RIe1f2648_4135, \9185_9484 );
and \U$6485 ( \15300_15599 , RIf14f108_5359, \9187_9486 );
and \U$6486 ( \15301_15600 , RIfc7f298_6469, \9189_9488 );
and \U$6487 ( \15302_15601 , RIf14d4e8_5339, \9191_9490 );
and \U$6488 ( \15303_15602 , RIe1ed350_4076, \9193_9492 );
and \U$6489 ( \15304_15603 , RIe1ea7b8_4045, \9195_9494 );
and \U$6490 ( \15305_15604 , RIe1e7ab8_4013, \9197_9496 );
and \U$6491 ( \15306_15605 , RIe1e4db8_3981, \9199_9498 );
and \U$6492 ( \15307_15606 , RIe1e20b8_3949, \9201_9500 );
and \U$6493 ( \15308_15607 , RIe1df3b8_3917, \9203_9502 );
and \U$6494 ( \15309_15608 , RIe1dc6b8_3885, \9205_9504 );
and \U$6495 ( \15310_15609 , RIe1d99b8_3853, \9207_9506 );
and \U$6496 ( \15311_15610 , RIe1d6cb8_3821, \9209_9508 );
and \U$6497 ( \15312_15611 , RIe1d12b8_3757, \9211_9510 );
and \U$6498 ( \15313_15612 , RIe1ce5b8_3725, \9213_9512 );
and \U$6499 ( \15314_15613 , RIe1cb8b8_3693, \9215_9514 );
and \U$6500 ( \15315_15614 , RIe1c8bb8_3661, \9217_9516 );
and \U$6501 ( \15316_15615 , RIe1c5eb8_3629, \9219_9518 );
and \U$6502 ( \15317_15616 , RIe1c31b8_3597, \9221_9520 );
and \U$6503 ( \15318_15617 , RIe1c04b8_3565, \9223_9522 );
and \U$6504 ( \15319_15618 , RIe1bd7b8_3533, \9225_9524 );
and \U$6505 ( \15320_15619 , RIf14c138_5325, \9227_9526 );
and \U$6506 ( \15321_15620 , RIf14ad88_5311, \9229_9528 );
and \U$6507 ( \15322_15621 , RIe1b8790_3476, \9231_9530 );
and \U$6508 ( \15323_15622 , RIfe96480_8054, \9233_9532 );
and \U$6509 ( \15324_15623 , RIf14a0e0_5302, \9235_9534 );
and \U$6510 ( \15325_15624 , RIf149870_5296, \9237_9536 );
and \U$6511 ( \15326_15625 , RIfe97128_8063, \9239_9538 );
and \U$6512 ( \15327_15626 , RIfe96318_8053, \9241_9540 );
and \U$6513 ( \15328_15627 , RIf148628_5283, \9243_9542 );
and \U$6514 ( \15329_15628 , RIfc58d78_6033, \9245_9544 );
and \U$6515 ( \15330_15629 , RIe1b20e8_3403, \9247_9546 );
and \U$6516 ( \15331_15630 , RIe1b04c8_3383, \9249_9548 );
and \U$6517 ( \15332_15631 , RIf146cd8_5265, \9251_9550 );
and \U$6518 ( \15333_15632 , RIfc591b0_6036, \9253_9552 );
and \U$6519 ( \15334_15633 , RIfe961b0_8052, \9255_9554 );
and \U$6520 ( \15335_15634 , RIfe96fc0_8062, \9257_9556 );
and \U$6521 ( \15336_15635 , RIe1a7af8_3285, \9259_9558 );
and \U$6522 ( \15337_15636 , RIe1a4df8_3253, \9261_9560 );
and \U$6523 ( \15338_15637 , RIe1a20f8_3221, \9263_9562 );
and \U$6524 ( \15339_15638 , RIe19f3f8_3189, \9265_9564 );
and \U$6525 ( \15340_15639 , RIe18b8f8_2965, \9267_9566 );
and \U$6526 ( \15341_15640 , RIe177df8_2741, \9269_9568 );
and \U$6527 ( \15342_15641 , RIe225750_4716, \9271_9570 );
and \U$6528 ( \15343_15642 , RIe21a350_4588, \9273_9572 );
and \U$6529 ( \15344_15643 , RIe203b50_4332, \9275_9574 );
and \U$6530 ( \15345_15644 , RIe1fdbb0_4264, \9277_9576 );
and \U$6531 ( \15346_15645 , RIe1f6f68_4187, \9279_9578 );
and \U$6532 ( \15347_15646 , RIe1efab0_4104, \9281_9580 );
and \U$6533 ( \15348_15647 , RIe1d3fb8_3789, \9283_9582 );
and \U$6534 ( \15349_15648 , RIe1baab8_3501, \9285_9584 );
and \U$6535 ( \15350_15649 , RIe1ad930_3352, \9287_9586 );
and \U$6536 ( \15351_15650 , RIe16ff68_2651, \9289_9588 );
or \U$6537 ( \15352_15651 , \15288_15587 , \15289_15588 , \15290_15589 , \15291_15590 , \15292_15591 , \15293_15592 , \15294_15593 , \15295_15594 , \15296_15595 , \15297_15596 , \15298_15597 , \15299_15598 , \15300_15599 , \15301_15600 , \15302_15601 , \15303_15602 , \15304_15603 , \15305_15604 , \15306_15605 , \15307_15606 , \15308_15607 , \15309_15608 , \15310_15609 , \15311_15610 , \15312_15611 , \15313_15612 , \15314_15613 , \15315_15614 , \15316_15615 , \15317_15616 , \15318_15617 , \15319_15618 , \15320_15619 , \15321_15620 , \15322_15621 , \15323_15622 , \15324_15623 , \15325_15624 , \15326_15625 , \15327_15626 , \15328_15627 , \15329_15628 , \15330_15629 , \15331_15630 , \15332_15631 , \15333_15632 , \15334_15633 , \15335_15634 , \15336_15635 , \15337_15636 , \15338_15637 , \15339_15638 , \15340_15639 , \15341_15640 , \15342_15641 , \15343_15642 , \15344_15643 , \15345_15644 , \15346_15645 , \15347_15646 , \15348_15647 , \15349_15648 , \15350_15649 , \15351_15650 );
or \U$6538 ( \15353_15652 , \15287_15586 , \15352_15651 );
_DC \g3dc6/U$1 ( \15354 , \15353_15652 , \9298_9597 );
buf \U$6539 ( \15355_15654 , \15354 );
xor \U$6540 ( \15356_15655 , \15222_15521 , \15355_15654 );
and \U$6541 ( \15357_15656 , RIdec42f8_696, \8760_9059 );
and \U$6542 ( \15358_15657 , RIdec15f8_664, \8762_9061 );
and \U$6543 ( \15359_15658 , RIfcc6cb0_7284, \8764_9063 );
and \U$6544 ( \15360_15659 , RIdebe8f8_632, \8766_9065 );
and \U$6545 ( \15361_15660 , RIfe93780_8022, \8768_9067 );
and \U$6546 ( \15362_15661 , RIdebbbf8_600, \8770_9069 );
and \U$6547 ( \15363_15662 , RIdeb8ef8_568, \8772_9071 );
and \U$6548 ( \15364_15663 , RIdeb61f8_536, \8774_9073 );
and \U$6549 ( \15365_15664 , RIee1ea00_4807, \8776_9075 );
and \U$6550 ( \15366_15665 , RIdeb07f8_472, \8778_9077 );
and \U$6551 ( \15367_15666 , RIee1e2f8_4802, \8780_9079 );
and \U$6552 ( \15368_15667 , RIdeadaf8_440, \8782_9081 );
and \U$6553 ( \15369_15668 , RIfc5d3c8_6083, \8784_9083 );
and \U$6554 ( \15370_15669 , RIdea7cc0_408, \8786_9085 );
and \U$6555 ( \15371_15670 , RIdea13c0_376, \8788_9087 );
and \U$6556 ( \15372_15671 , RIde9aac0_344, \8790_9089 );
and \U$6557 ( \15373_15672 , RIfc58238_6025, \8792_9091 );
and \U$6558 ( \15374_15673 , RIfcc3b78_7249, \8794_9093 );
and \U$6559 ( \15375_15674 , RIfc7d0d8_6445, \8796_9095 );
and \U$6560 ( \15376_15675 , RIfc59750_6040, \8798_9097 );
and \U$6561 ( \15377_15676 , RIfe93a50_8024, \8800_9099 );
and \U$6562 ( \15378_15677 , RIfe938e8_8023, \8802_9101 );
and \U$6563 ( \15379_15678 , RIde88370_254, \8804_9103 );
and \U$6564 ( \15380_15679 , RIde83e88_233, \8806_9105 );
and \U$6565 ( \15381_15680 , RIfc5f420_6106, \8808_9107 );
and \U$6566 ( \15382_15681 , RIfc976b8_6745, \8810_9109 );
and \U$6567 ( \15383_15682 , RIfc90a70_6668, \8812_9111 );
and \U$6568 ( \15384_15683 , RIfc60500_6118, \8814_9113 );
and \U$6569 ( \15385_15684 , RIee38a40_5103, \8816_9115 );
and \U$6570 ( \15386_15685 , RIe16ab08_2591, \8818_9117 );
and \U$6571 ( \15387_15686 , RIe169488_2575, \8820_9119 );
and \U$6572 ( \15388_15687 , RIe166ff8_2549, \8822_9121 );
and \U$6573 ( \15389_15688 , RIe1642f8_2517, \8824_9123 );
and \U$6574 ( \15390_15689 , RIe1615f8_2485, \8826_9125 );
and \U$6575 ( \15391_15690 , RIee369e8_5080, \8828_9127 );
and \U$6576 ( \15392_15691 , RIe15e8f8_2453, \8830_9129 );
and \U$6577 ( \15393_15692 , RIee35bd8_5070, \8832_9131 );
and \U$6578 ( \15394_15693 , RIe15bbf8_2421, \8834_9133 );
and \U$6579 ( \15395_15694 , RIe1561f8_2357, \8836_9135 );
and \U$6580 ( \15396_15695 , RIe1534f8_2325, \8838_9137 );
and \U$6581 ( \15397_15696 , RIfc3ee28_5741, \8840_9139 );
and \U$6582 ( \15398_15697 , RIe1507f8_2293, \8842_9141 );
and \U$6583 ( \15399_15698 , RIfce6c90_7648, \8844_9143 );
and \U$6584 ( \15400_15699 , RIe14daf8_2261, \8846_9145 );
and \U$6585 ( \15401_15700 , RIfcca7c0_7326, \8848_9147 );
and \U$6586 ( \15402_15701 , RIe14adf8_2229, \8850_9149 );
and \U$6587 ( \15403_15702 , RIe1480f8_2197, \8852_9151 );
and \U$6588 ( \15404_15703 , RIe1453f8_2165, \8854_9153 );
and \U$6589 ( \15405_15704 , RIee33b80_5047, \8856_9155 );
and \U$6590 ( \15406_15705 , RIee32938_5034, \8858_9157 );
and \U$6591 ( \15407_15706 , RIee316f0_5021, \8860_9159 );
and \U$6592 ( \15408_15707 , RIee30bb0_5013, \8862_9161 );
and \U$6593 ( \15409_15708 , RIe1403d0_2108, \8864_9163 );
and \U$6594 ( \15410_15709 , RIfe93618_8021, \8866_9165 );
and \U$6595 ( \15411_15710 , RIdf3bfb0_2059, \8868_9167 );
and \U$6596 ( \15412_15711 , RIfe934b0_8020, \8870_9169 );
and \U$6597 ( \15413_15712 , RIfcd0d00_7398, \8872_9171 );
and \U$6598 ( \15414_15713 , RIee2ecc0_4991, \8874_9173 );
and \U$6599 ( \15415_15714 , RIee2e720_4987, \8876_9175 );
and \U$6600 ( \15416_15715 , RIee2cb00_4967, \8878_9177 );
and \U$6601 ( \15417_15716 , RIfe93bb8_8025, \8880_9179 );
and \U$6602 ( \15418_15717 , RIdf32938_1952, \8882_9181 );
and \U$6603 ( \15419_15718 , RIdf30340_1925, \8884_9183 );
and \U$6604 ( \15420_15719 , RIdf2e450_1903, \8886_9185 );
or \U$6605 ( \15421_15720 , \15357_15656 , \15358_15657 , \15359_15658 , \15360_15659 , \15361_15660 , \15362_15661 , \15363_15662 , \15364_15663 , \15365_15664 , \15366_15665 , \15367_15666 , \15368_15667 , \15369_15668 , \15370_15669 , \15371_15670 , \15372_15671 , \15373_15672 , \15374_15673 , \15375_15674 , \15376_15675 , \15377_15676 , \15378_15677 , \15379_15678 , \15380_15679 , \15381_15680 , \15382_15681 , \15383_15682 , \15384_15683 , \15385_15684 , \15386_15685 , \15387_15686 , \15388_15687 , \15389_15688 , \15390_15689 , \15391_15690 , \15392_15691 , \15393_15692 , \15394_15693 , \15395_15694 , \15396_15695 , \15397_15696 , \15398_15697 , \15399_15698 , \15400_15699 , \15401_15700 , \15402_15701 , \15403_15702 , \15404_15703 , \15405_15704 , \15406_15705 , \15407_15706 , \15408_15707 , \15409_15708 , \15410_15709 , \15411_15710 , \15412_15711 , \15413_15712 , \15414_15713 , \15415_15714 , \15416_15715 , \15417_15716 , \15418_15717 , \15419_15718 , \15420_15719 );
and \U$6606 ( \15422_15721 , RIee2b048_4948, \8889_9188 );
and \U$6607 ( \15423_15722 , RIee29b30_4933, \8891_9190 );
and \U$6608 ( \15424_15723 , RIfc67148_6195, \8893_9192 );
and \U$6609 ( \15425_15724 , RIfc6fb18_6293, \8895_9194 );
and \U$6610 ( \15426_15725 , RIdf29860_1849, \8897_9196 );
and \U$6611 ( \15427_15726 , RIfe931e0_8018, \8899_9198 );
and \U$6612 ( \15428_15727 , RIfe93348_8019, \8901_9200 );
and \U$6613 ( \15429_15728 , RIfe93078_8017, \8903_9202 );
and \U$6614 ( \15430_15729 , RIfc672b0_6196, \8905_9204 );
and \U$6615 ( \15431_15730 , RIfca8788_6939, \8907_9206 );
and \U$6616 ( \15432_15731 , RIdf22510_1767, \8909_9208 );
and \U$6617 ( \15433_15732 , RIfcea7a0_7690, \8911_9210 );
and \U$6618 ( \15434_15733 , RIdf20ff8_1752, \8913_9212 );
and \U$6619 ( \15435_15734 , RIdf1ecd0_1727, \8915_9214 );
and \U$6620 ( \15436_15735 , RIdf1aab8_1680, \8917_9216 );
and \U$6621 ( \15437_15736 , RIfea7c58_8225, \8919_9218 );
and \U$6622 ( \15438_15737 , RIdf15ec8_1626, \8921_9220 );
and \U$6623 ( \15439_15738 , RIdf131c8_1594, \8923_9222 );
and \U$6624 ( \15440_15739 , RIdf104c8_1562, \8925_9224 );
and \U$6625 ( \15441_15740 , RIdf0d7c8_1530, \8927_9226 );
and \U$6626 ( \15442_15741 , RIdf0aac8_1498, \8929_9228 );
and \U$6627 ( \15443_15742 , RIdf07dc8_1466, \8931_9230 );
and \U$6628 ( \15444_15743 , RIdf050c8_1434, \8933_9232 );
and \U$6629 ( \15445_15744 , RIdf023c8_1402, \8935_9234 );
and \U$6630 ( \15446_15745 , RIdefc9c8_1338, \8937_9236 );
and \U$6631 ( \15447_15746 , RIdef9cc8_1306, \8939_9238 );
and \U$6632 ( \15448_15747 , RIdef6fc8_1274, \8941_9240 );
and \U$6633 ( \15449_15748 , RIdef42c8_1242, \8943_9242 );
and \U$6634 ( \15450_15749 , RIdef15c8_1210, \8945_9244 );
and \U$6635 ( \15451_15750 , RIdeee8c8_1178, \8947_9246 );
and \U$6636 ( \15452_15751 , RIdeebbc8_1146, \8949_9248 );
and \U$6637 ( \15453_15752 , RIdee8ec8_1114, \8951_9250 );
and \U$6638 ( \15454_15753 , RIee24f40_4879, \8953_9252 );
and \U$6639 ( \15455_15754 , RIee24130_4869, \8955_9254 );
and \U$6640 ( \15456_15755 , RIee235f0_4861, \8957_9256 );
and \U$6641 ( \15457_15756 , RIee22c18_4854, \8959_9258 );
and \U$6642 ( \15458_15757 , RIfe93d20_8026, \8961_9260 );
and \U$6643 ( \15459_15758 , RIdee1fb0_1035, \8963_9262 );
and \U$6644 ( \15460_15759 , RIdee0228_1014, \8965_9264 );
and \U$6645 ( \15461_15760 , RIdeddc30_987, \8967_9266 );
and \U$6646 ( \15462_15761 , RIfc684f8_6209, \8969_9268 );
and \U$6647 ( \15463_15762 , RIee21ca0_4843, \8971_9270 );
and \U$6648 ( \15464_15763 , RIfc68390_6208, \8973_9272 );
and \U$6649 ( \15465_15764 , RIee20d28_4832, \8975_9274 );
and \U$6650 ( \15466_15765 , RIded8aa0_929, \8977_9276 );
and \U$6651 ( \15467_15766 , RIfe93ff0_8028, \8979_9278 );
and \U$6652 ( \15468_15767 , RIded45b8_880, \8981_9280 );
and \U$6653 ( \15469_15768 , RIfe93e88_8027, \8983_9282 );
and \U$6654 ( \15470_15769 , RIdecf6f8_824, \8985_9284 );
and \U$6655 ( \15471_15770 , RIdecc9f8_792, \8987_9286 );
and \U$6656 ( \15472_15771 , RIdec9cf8_760, \8989_9288 );
and \U$6657 ( \15473_15772 , RIdec6ff8_728, \8991_9290 );
and \U$6658 ( \15474_15773 , RIdeb34f8_504, \8993_9292 );
and \U$6659 ( \15475_15774 , RIde941c0_312, \8995_9294 );
and \U$6660 ( \15476_15775 , RIe16d100_2618, \8997_9296 );
and \U$6661 ( \15477_15776 , RIe158ef8_2389, \8999_9298 );
and \U$6662 ( \15478_15777 , RIe1426f8_2133, \9001_9300 );
and \U$6663 ( \15479_15778 , RIdf370f0_2003, \9003_9302 );
and \U$6664 ( \15480_15779 , RIdf2b750_1871, \9005_9304 );
and \U$6665 ( \15481_15780 , RIdf1bfd0_1695, \9007_9306 );
and \U$6666 ( \15482_15781 , RIdeff6c8_1370, \9009_9308 );
and \U$6667 ( \15483_15782 , RIdee61c8_1082, \9011_9310 );
and \U$6668 ( \15484_15783 , RIdedaf30_955, \9013_9312 );
and \U$6669 ( \15485_15784 , RIde7a108_185, \9015_9314 );
or \U$6670 ( \15486_15785 , \15422_15721 , \15423_15722 , \15424_15723 , \15425_15724 , \15426_15725 , \15427_15726 , \15428_15727 , \15429_15728 , \15430_15729 , \15431_15730 , \15432_15731 , \15433_15732 , \15434_15733 , \15435_15734 , \15436_15735 , \15437_15736 , \15438_15737 , \15439_15738 , \15440_15739 , \15441_15740 , \15442_15741 , \15443_15742 , \15444_15743 , \15445_15744 , \15446_15745 , \15447_15746 , \15448_15747 , \15449_15748 , \15450_15749 , \15451_15750 , \15452_15751 , \15453_15752 , \15454_15753 , \15455_15754 , \15456_15755 , \15457_15756 , \15458_15757 , \15459_15758 , \15460_15759 , \15461_15760 , \15462_15761 , \15463_15762 , \15464_15763 , \15465_15764 , \15466_15765 , \15467_15766 , \15468_15767 , \15469_15768 , \15470_15769 , \15471_15770 , \15472_15771 , \15473_15772 , \15474_15773 , \15475_15774 , \15476_15775 , \15477_15776 , \15478_15777 , \15479_15778 , \15480_15779 , \15481_15780 , \15482_15781 , \15483_15782 , \15484_15783 , \15485_15784 );
or \U$6671 ( \15487_15786 , \15421_15720 , \15486_15785 );
_DC \g2d1e/U$1 ( \15488 , \15487_15786 , \9024_9323 );
buf \U$6672 ( \15489_15788 , \15488 );
and \U$6673 ( \15490_15789 , RIe19c590_3156, \9034_9333 );
and \U$6674 ( \15491_15790 , RIe199890_3124, \9036_9335 );
and \U$6675 ( \15492_15791 , RIf144f50_5244, \9038_9337 );
and \U$6676 ( \15493_15792 , RIe196b90_3092, \9040_9339 );
and \U$6677 ( \15494_15793 , RIfc76058_6365, \9042_9341 );
and \U$6678 ( \15495_15794 , RIe193e90_3060, \9044_9343 );
and \U$6679 ( \15496_15795 , RIe191190_3028, \9046_9345 );
and \U$6680 ( \15497_15796 , RIe18e490_2996, \9048_9347 );
and \U$6681 ( \15498_15797 , RIe188a90_2932, \9050_9349 );
and \U$6682 ( \15499_15798 , RIe185d90_2900, \9052_9351 );
and \U$6683 ( \15500_15799 , RIfccd8f8_7361, \9054_9353 );
and \U$6684 ( \15501_15800 , RIe183090_2868, \9056_9355 );
and \U$6685 ( \15502_15801 , RIfc76e68_6375, \9058_9357 );
and \U$6686 ( \15503_15802 , RIe180390_2836, \9060_9359 );
and \U$6687 ( \15504_15803 , RIe17d690_2804, \9062_9361 );
and \U$6688 ( \15505_15804 , RIe17a990_2772, \9064_9363 );
and \U$6689 ( \15506_15805 , RIf1419e0_5206, \9066_9365 );
and \U$6690 ( \15507_15806 , RIf140630_5192, \9068_9367 );
and \U$6691 ( \15508_15807 , RIe176bb0_2728, \9070_9369 );
and \U$6692 ( \15509_15808 , RIe1750f8_2709, \9072_9371 );
and \U$6693 ( \15510_15809 , RIfcd1840_7406, \9074_9373 );
and \U$6694 ( \15511_15810 , RIfc5f6f0_6108, \9076_9375 );
and \U$6695 ( \15512_15811 , RIee3dd38_5162, \9078_9377 );
and \U$6696 ( \15513_15812 , RIee3cc58_5150, \9080_9379 );
and \U$6697 ( \15514_15813 , RIee3b8a8_5136, \9082_9381 );
and \U$6698 ( \15515_15814 , RIee3a7c8_5124, \9084_9383 );
and \U$6699 ( \15516_15815 , RIee39580_5111, \9086_9385 );
and \U$6700 ( \15517_15816 , RIfea9008_8239, \9088_9387 );
and \U$6701 ( \15518_15817 , RIf16f7f0_5728, \9090_9389 );
and \U$6702 ( \15519_15818 , RIf16ecb0_5720, \9092_9391 );
and \U$6703 ( \15520_15819 , RIf16d900_5706, \9094_9393 );
and \U$6704 ( \15521_15820 , RIfc78ec0_6398, \9096_9395 );
and \U$6705 ( \15522_15821 , RIfcc8060_7298, \9098_9397 );
and \U$6706 ( \15523_15822 , RIe2228e8_4683, \9100_9399 );
and \U$6707 ( \15524_15823 , RIfc5a3f8_6049, \9102_9401 );
and \U$6708 ( \15525_15824 , RIe21fbe8_4651, \9104_9403 );
and \U$6709 ( \15526_15825 , RIfc74000_6342, \9106_9405 );
and \U$6710 ( \15527_15826 , RIe21cee8_4619, \9108_9407 );
and \U$6711 ( \15528_15827 , RIe2174e8_4555, \9110_9409 );
and \U$6712 ( \15529_15828 , RIe2147e8_4523, \9112_9411 );
and \U$6713 ( \15530_15829 , RIfca2c20_6874, \9114_9413 );
and \U$6714 ( \15531_15830 , RIe211ae8_4491, \9116_9415 );
and \U$6715 ( \15532_15831 , RIfca2950_6872, \9118_9417 );
and \U$6716 ( \15533_15832 , RIe20ede8_4459, \9120_9419 );
and \U$6717 ( \15534_15833 , RIfcc24f8_7233, \9122_9421 );
and \U$6718 ( \15535_15834 , RIe20c0e8_4427, \9124_9423 );
and \U$6719 ( \15536_15835 , RIe2093e8_4395, \9126_9425 );
and \U$6720 ( \15537_15836 , RIe2066e8_4363, \9128_9427 );
and \U$6721 ( \15538_15837 , RIfc45110_5808, \9130_9429 );
and \U$6722 ( \15539_15838 , RIfcc6f80_7286, \9132_9431 );
and \U$6723 ( \15540_15839 , RIfe92f10_8016, \9134_9433 );
and \U$6724 ( \15541_15840 , RIfe92970_8012, \9136_9435 );
and \U$6725 ( \15542_15841 , RIf164af8_5605, \9138_9437 );
and \U$6726 ( \15543_15842 , RIf163a18_5593, \9140_9439 );
and \U$6727 ( \15544_15843 , RIf162aa0_5582, \9142_9441 );
and \U$6728 ( \15545_15844 , RIfe92ad8_8013, \9144_9443 );
and \U$6729 ( \15546_15845 , RIf15f3c8_5543, \9146_9445 );
and \U$6730 ( \15547_15846 , RIf15d640_5522, \9148_9447 );
and \U$6731 ( \15548_15847 , RIfe92808_8011, \9150_9449 );
and \U$6732 ( \15549_15848 , RIfe92c40_8014, \9152_9451 );
and \U$6733 ( \15550_15849 , RIfe926a0_8010, \9154_9453 );
and \U$6734 ( \15551_15850 , RIfe92da8_8015, \9156_9455 );
and \U$6735 ( \15552_15851 , RIfe92538_8009, \9158_9457 );
and \U$6736 ( \15553_15852 , RIfcb5a78_7089, \9160_9459 );
or \U$6737 ( \15554_15853 , \15490_15789 , \15491_15790 , \15492_15791 , \15493_15792 , \15494_15793 , \15495_15794 , \15496_15795 , \15497_15796 , \15498_15797 , \15499_15798 , \15500_15799 , \15501_15800 , \15502_15801 , \15503_15802 , \15504_15803 , \15505_15804 , \15506_15805 , \15507_15806 , \15508_15807 , \15509_15808 , \15510_15809 , \15511_15810 , \15512_15811 , \15513_15812 , \15514_15813 , \15515_15814 , \15516_15815 , \15517_15816 , \15518_15817 , \15519_15818 , \15520_15819 , \15521_15820 , \15522_15821 , \15523_15822 , \15524_15823 , \15525_15824 , \15526_15825 , \15527_15826 , \15528_15827 , \15529_15828 , \15530_15829 , \15531_15830 , \15532_15831 , \15533_15832 , \15534_15833 , \15535_15834 , \15536_15835 , \15537_15836 , \15538_15837 , \15539_15838 , \15540_15839 , \15541_15840 , \15542_15841 , \15543_15842 , \15544_15843 , \15545_15844 , \15546_15845 , \15547_15846 , \15548_15847 , \15549_15848 , \15550_15849 , \15551_15850 , \15552_15851 , \15553_15852 );
and \U$6738 ( \15555_15854 , RIf158348_5463, \9163_9462 );
and \U$6739 ( \15556_15855 , RIf157100_5450, \9165_9464 );
and \U$6740 ( \15557_15856 , RIfc53be8_5975, \9167_9466 );
and \U$6741 ( \15558_15857 , RIfec38b8_8345, \9169_9468 );
and \U$6742 ( \15559_15858 , RIfcc5ea0_7274, \9171_9470 );
and \U$6743 ( \15560_15859 , RIf1550a8_5427, \9173_9472 );
and \U$6744 ( \15561_15860 , RIf153cf8_5413, \9175_9474 );
and \U$6745 ( \15562_15861 , RIfec3a20_8346, \9177_9476 );
and \U$6746 ( \15563_15862 , RIf152678_5397, \9179_9478 );
and \U$6747 ( \15564_15863 , RIfec3750_8344, \9181_9480 );
and \U$6748 ( \15565_15864 , RIf14ff18_5369, \9183_9482 );
and \U$6749 ( \15566_15865 , RIfe923d0_8008, \9185_9484 );
and \U$6750 ( \15567_15866 , RIf14efa0_5358, \9187_9486 );
and \U$6751 ( \15568_15867 , RIf14e898_5353, \9189_9488 );
and \U$6752 ( \15569_15868 , RIf14d380_5338, \9191_9490 );
and \U$6753 ( \15570_15869 , RIfe92268_8007, \9193_9492 );
and \U$6754 ( \15571_15870 , RIe1ea650_4044, \9195_9494 );
and \U$6755 ( \15572_15871 , RIe1e7950_4012, \9197_9496 );
and \U$6756 ( \15573_15872 , RIe1e4c50_3980, \9199_9498 );
and \U$6757 ( \15574_15873 , RIe1e1f50_3948, \9201_9500 );
and \U$6758 ( \15575_15874 , RIe1df250_3916, \9203_9502 );
and \U$6759 ( \15576_15875 , RIe1dc550_3884, \9205_9504 );
and \U$6760 ( \15577_15876 , RIe1d9850_3852, \9207_9506 );
and \U$6761 ( \15578_15877 , RIe1d6b50_3820, \9209_9508 );
and \U$6762 ( \15579_15878 , RIe1d1150_3756, \9211_9510 );
and \U$6763 ( \15580_15879 , RIe1ce450_3724, \9213_9512 );
and \U$6764 ( \15581_15880 , RIe1cb750_3692, \9215_9514 );
and \U$6765 ( \15582_15881 , RIe1c8a50_3660, \9217_9516 );
and \U$6766 ( \15583_15882 , RIe1c5d50_3628, \9219_9518 );
and \U$6767 ( \15584_15883 , RIe1c3050_3596, \9221_9520 );
and \U$6768 ( \15585_15884 , RIe1c0350_3564, \9223_9522 );
and \U$6769 ( \15586_15885 , RIe1bd650_3532, \9225_9524 );
and \U$6770 ( \15587_15886 , RIfcda4e0_7506, \9227_9526 );
and \U$6771 ( \15588_15887 , RIfc9d220_6810, \9229_9528 );
and \U$6772 ( \15589_15888 , RIe1b8628_3475, \9231_9530 );
and \U$6773 ( \15590_15889 , RIe1b6738_3453, \9233_9532 );
and \U$6774 ( \15591_15890 , RIfc4f2c8_5923, \9235_9534 );
and \U$6775 ( \15592_15891 , RIfce16c8_7587, \9237_9536 );
and \U$6776 ( \15593_15892 , RIfe91cc8_8003, \9239_9538 );
and \U$6777 ( \15594_15893 , RIfe91e30_8004, \9241_9540 );
and \U$6778 ( \15595_15894 , RIf1484c0_5282, \9243_9542 );
and \U$6779 ( \15596_15895 , RIf147548_5271, \9245_9544 );
and \U$6780 ( \15597_15896 , RIfe91f98_8005, \9247_9546 );
and \U$6781 ( \15598_15897 , RIfe91b60_8002, \9249_9548 );
and \U$6782 ( \15599_15898 , RIf146b70_5264, \9251_9550 );
and \U$6783 ( \15600_15899 , RIfc9f548_6835, \9253_9552 );
and \U$6784 ( \15601_15900 , RIfe92100_8006, \9255_9554 );
and \U$6785 ( \15602_15901 , RIfe919f8_8001, \9257_9556 );
and \U$6786 ( \15603_15902 , RIe1a7990_3284, \9259_9558 );
and \U$6787 ( \15604_15903 , RIe1a4c90_3252, \9261_9560 );
and \U$6788 ( \15605_15904 , RIe1a1f90_3220, \9263_9562 );
and \U$6789 ( \15606_15905 , RIe19f290_3188, \9265_9564 );
and \U$6790 ( \15607_15906 , RIe18b790_2964, \9267_9566 );
and \U$6791 ( \15608_15907 , RIe177c90_2740, \9269_9568 );
and \U$6792 ( \15609_15908 , RIe2255e8_4715, \9271_9570 );
and \U$6793 ( \15610_15909 , RIe21a1e8_4587, \9273_9572 );
and \U$6794 ( \15611_15910 , RIe2039e8_4331, \9275_9574 );
and \U$6795 ( \15612_15911 , RIe1fda48_4263, \9277_9576 );
and \U$6796 ( \15613_15912 , RIe1f6e00_4186, \9279_9578 );
and \U$6797 ( \15614_15913 , RIe1ef948_4103, \9281_9580 );
and \U$6798 ( \15615_15914 , RIe1d3e50_3788, \9283_9582 );
and \U$6799 ( \15616_15915 , RIe1ba950_3500, \9285_9584 );
and \U$6800 ( \15617_15916 , RIe1ad7c8_3351, \9287_9586 );
and \U$6801 ( \15618_15917 , RIe16fe00_2650, \9289_9588 );
or \U$6802 ( \15619_15918 , \15555_15854 , \15556_15855 , \15557_15856 , \15558_15857 , \15559_15858 , \15560_15859 , \15561_15860 , \15562_15861 , \15563_15862 , \15564_15863 , \15565_15864 , \15566_15865 , \15567_15866 , \15568_15867 , \15569_15868 , \15570_15869 , \15571_15870 , \15572_15871 , \15573_15872 , \15574_15873 , \15575_15874 , \15576_15875 , \15577_15876 , \15578_15877 , \15579_15878 , \15580_15879 , \15581_15880 , \15582_15881 , \15583_15882 , \15584_15883 , \15585_15884 , \15586_15885 , \15587_15886 , \15588_15887 , \15589_15888 , \15590_15889 , \15591_15890 , \15592_15891 , \15593_15892 , \15594_15893 , \15595_15894 , \15596_15895 , \15597_15896 , \15598_15897 , \15599_15898 , \15600_15899 , \15601_15900 , \15602_15901 , \15603_15902 , \15604_15903 , \15605_15904 , \15606_15905 , \15607_15906 , \15608_15907 , \15609_15908 , \15610_15909 , \15611_15910 , \15612_15911 , \15613_15912 , \15614_15913 , \15615_15914 , \15616_15915 , \15617_15916 , \15618_15917 );
or \U$6803 ( \15620_15919 , \15554_15853 , \15619_15918 );
_DC \g3e4b/U$1 ( \15621 , \15620_15919 , \9298_9597 );
buf \U$6804 ( \15622_15921 , \15621 );
and \U$6805 ( \15623_15922 , \15489_15788 , \15622_15921 );
and \U$6806 ( \15624_15923 , \13913_14212 , \14046_14345 );
and \U$6807 ( \15625_15924 , \14046_14345 , \14321_14620 );
and \U$6808 ( \15626_15925 , \13913_14212 , \14321_14620 );
or \U$6809 ( \15627_15926 , \15624_15923 , \15625_15924 , \15626_15925 );
and \U$6810 ( \15628_15927 , \15622_15921 , \15627_15926 );
and \U$6811 ( \15629_15928 , \15489_15788 , \15627_15926 );
or \U$6812 ( \15630_15929 , \15623_15922 , \15628_15927 , \15629_15928 );
xor \U$6813 ( \15631_15930 , \15356_15655 , \15630_15929 );
buf g4436_GF_PartitionCandidate( \15632_15931_nG4436 , \15631_15930 );
xor \U$6814 ( \15633_15932 , \15489_15788 , \15622_15921 );
xor \U$6815 ( \15634_15933 , \15633_15932 , \15627_15926 );
buf g4439_GF_PartitionCandidate( \15635_15934_nG4439 , \15634_15933 );
nand \U$6816 ( \15636_15935 , \15635_15934_nG4439 , \14323_14622_nG443c );
and \U$6817 ( \15637_15936 , \15632_15931_nG4436 , \15636_15935 );
xor \U$6818 ( \15638_15937 , \15635_15934_nG4439 , \14323_14622_nG443c );
and \U$6823 ( \15639_15941 , \15638_15937 , \10392_10694_nG9c0e );
or \U$6824 ( \15640_15942 , 1'b0 , \15639_15941 );
xor \U$6825 ( \15641_15943 , \15637_15936 , \15640_15942 );
xor \U$6826 ( \15642_15944 , \15637_15936 , \15641_15943 );
buf \U$6827 ( \15643_15945 , \15642_15944 );
buf \U$6828 ( \15644_15946 , \15643_15945 );
and \U$6829 ( \15645_15947 , \15089_15388 , \15644_15946 );
and \U$6830 ( \15646_15948 , \14733_15032 , \14749_15048 );
and \U$6831 ( \15647_15949 , \14733_15032 , \15079_15378 );
and \U$6832 ( \15648_15950 , \14749_15048 , \15079_15378 );
or \U$6833 ( \15649_15951 , \15646_15948 , \15647_15949 , \15648_15950 );
buf \U$6834 ( \15650_15952 , \15649_15951 );
and \U$6835 ( \15651_15953 , \14738_15037 , \14740_15039 );
and \U$6836 ( \15652_15954 , \14738_15037 , \14747_15046 );
and \U$6837 ( \15653_15955 , \14740_15039 , \14747_15046 );
or \U$6838 ( \15654_15956 , \15651_15953 , \15652_15954 , \15653_15955 );
buf \U$6839 ( \15655_15957 , \15654_15956 );
and \U$6840 ( \15656_15958 , \14710_14631 , \10693_10995_nG9c0b );
and \U$6841 ( \15657_15959 , \14329_14628 , \10981_11283_nG9c08 );
or \U$6842 ( \15658_15960 , \15656_15958 , \15657_15959 );
xor \U$6843 ( \15659_15961 , \14328_14627 , \15658_15960 );
buf \U$6844 ( \15660_15962 , \15659_15961 );
buf \U$6846 ( \15661_15963 , \15660_15962 );
and \U$6847 ( \15662_15964 , \13431_13370 , \11299_11598_nG9c05 );
and \U$6848 ( \15663_15965 , \13068_13367 , \12168_12470_nG9c02 );
or \U$6849 ( \15664_15966 , \15662_15964 , \15663_15965 );
xor \U$6850 ( \15665_15967 , \13067_13366 , \15664_15966 );
buf \U$6851 ( \15666_15968 , \15665_15967 );
buf \U$6853 ( \15667_15969 , \15666_15968 );
xor \U$6854 ( \15668_15970 , \15661_15963 , \15667_15969 );
buf \U$6855 ( \15669_15971 , \15668_15970 );
and \U$6856 ( \15670_15972 , \14707_15009 , \14716_15015 );
buf \U$6857 ( \15671_15973 , \15670_15972 );
xor \U$6858 ( \15672_15974 , \15669_15971 , \15671_15973 );
and \U$6859 ( \15673_15975 , \12183_12157 , \12502_12801_nG9bff );
and \U$6860 ( \15674_15976 , \11855_12154 , \13403_13705_nG9bfc );
or \U$6861 ( \15675_15977 , \15673_15975 , \15674_15976 );
xor \U$6862 ( \15676_15978 , \11854_12153 , \15675_15977 );
buf \U$6863 ( \15677_15979 , \15676_15978 );
buf \U$6865 ( \15678_15980 , \15677_15979 );
xor \U$6866 ( \15679_15981 , \15672_15974 , \15678_15980 );
buf \U$6867 ( \15680_15982 , \15679_15981 );
xor \U$6868 ( \15681_15983 , \15655_15957 , \15680_15982 );
and \U$6869 ( \15682_15984 , \14718_15017 , \14724_15023 );
and \U$6870 ( \15683_15985 , \14718_15017 , \14731_15030 );
and \U$6871 ( \15684_15986 , \14724_15023 , \14731_15030 );
or \U$6872 ( \15685_15987 , \15682_15984 , \15683_15985 , \15684_15986 );
buf \U$6873 ( \15686_15988 , \15685_15987 );
and \U$6874 ( \15687_15989 , \10996_10421 , \13771_14070_nG9bf9 );
and \U$6875 ( \15688_15990 , \10119_10418 , \14682_14984_nG9bf6 );
or \U$6876 ( \15689_15991 , \15687_15989 , \15688_15990 );
xor \U$6877 ( \15690_15992 , \10118_10417 , \15689_15991 );
buf \U$6878 ( \15691_15993 , \15690_15992 );
buf \U$6880 ( \15692_15994 , \15691_15993 );
xor \U$6881 ( \15693_15995 , \15686_15988 , \15692_15994 );
and \U$6882 ( \15694_15996 , \10411_10707 , \15074_15373_nG9bf3 );
and \U$6883 ( \15695_15997 , \15053_15352 , \15057_15356 );
and \U$6884 ( \15696_15998 , \15057_15356 , \15062_15361 );
and \U$6885 ( \15697_15999 , \15053_15352 , \15062_15361 );
or \U$6886 ( \15698_16000 , \15695_15997 , \15696_15998 , \15697_15999 );
and \U$6887 ( \15699_16001 , \15022_15321 , \10681_10983 );
and \U$6888 ( \15700_16002 , RIdec42f8_696, \9034_9333 );
and \U$6889 ( \15701_16003 , RIdec15f8_664, \9036_9335 );
and \U$6890 ( \15702_16004 , RIfcc6cb0_7284, \9038_9337 );
and \U$6891 ( \15703_16005 , RIdebe8f8_632, \9040_9339 );
and \U$6892 ( \15704_16006 , RIfe93780_8022, \9042_9341 );
and \U$6893 ( \15705_16007 , RIdebbbf8_600, \9044_9343 );
and \U$6894 ( \15706_16008 , RIdeb8ef8_568, \9046_9345 );
and \U$6895 ( \15707_16009 , RIdeb61f8_536, \9048_9347 );
and \U$6896 ( \15708_16010 , RIee1ea00_4807, \9050_9349 );
and \U$6897 ( \15709_16011 , RIdeb07f8_472, \9052_9351 );
and \U$6898 ( \15710_16012 , RIee1e2f8_4802, \9054_9353 );
and \U$6899 ( \15711_16013 , RIdeadaf8_440, \9056_9355 );
and \U$6900 ( \15712_16014 , RIfc5d3c8_6083, \9058_9357 );
and \U$6901 ( \15713_16015 , RIdea7cc0_408, \9060_9359 );
and \U$6902 ( \15714_16016 , RIdea13c0_376, \9062_9361 );
and \U$6903 ( \15715_16017 , RIde9aac0_344, \9064_9363 );
and \U$6904 ( \15716_16018 , RIfc58238_6025, \9066_9365 );
and \U$6905 ( \15717_16019 , RIfcc3b78_7249, \9068_9367 );
and \U$6906 ( \15718_16020 , RIfc7d0d8_6445, \9070_9369 );
and \U$6907 ( \15719_16021 , RIfc59750_6040, \9072_9371 );
and \U$6908 ( \15720_16022 , RIfe93a50_8024, \9074_9373 );
and \U$6909 ( \15721_16023 , RIfe938e8_8023, \9076_9375 );
and \U$6910 ( \15722_16024 , RIde88370_254, \9078_9377 );
and \U$6911 ( \15723_16025 , RIde83e88_233, \9080_9379 );
and \U$6912 ( \15724_16026 , RIfc5f420_6106, \9082_9381 );
and \U$6913 ( \15725_16027 , RIfc976b8_6745, \9084_9383 );
and \U$6914 ( \15726_16028 , RIfc90a70_6668, \9086_9385 );
and \U$6915 ( \15727_16029 , RIfc60500_6118, \9088_9387 );
and \U$6916 ( \15728_16030 , RIee38a40_5103, \9090_9389 );
and \U$6917 ( \15729_16031 , RIe16ab08_2591, \9092_9391 );
and \U$6918 ( \15730_16032 , RIe169488_2575, \9094_9393 );
and \U$6919 ( \15731_16033 , RIe166ff8_2549, \9096_9395 );
and \U$6920 ( \15732_16034 , RIe1642f8_2517, \9098_9397 );
and \U$6921 ( \15733_16035 , RIe1615f8_2485, \9100_9399 );
and \U$6922 ( \15734_16036 , RIee369e8_5080, \9102_9401 );
and \U$6923 ( \15735_16037 , RIe15e8f8_2453, \9104_9403 );
and \U$6924 ( \15736_16038 , RIee35bd8_5070, \9106_9405 );
and \U$6925 ( \15737_16039 , RIe15bbf8_2421, \9108_9407 );
and \U$6926 ( \15738_16040 , RIe1561f8_2357, \9110_9409 );
and \U$6927 ( \15739_16041 , RIe1534f8_2325, \9112_9411 );
and \U$6928 ( \15740_16042 , RIfc3ee28_5741, \9114_9413 );
and \U$6929 ( \15741_16043 , RIe1507f8_2293, \9116_9415 );
and \U$6930 ( \15742_16044 , RIfce6c90_7648, \9118_9417 );
and \U$6931 ( \15743_16045 , RIe14daf8_2261, \9120_9419 );
and \U$6932 ( \15744_16046 , RIfcca7c0_7326, \9122_9421 );
and \U$6933 ( \15745_16047 , RIe14adf8_2229, \9124_9423 );
and \U$6934 ( \15746_16048 , RIe1480f8_2197, \9126_9425 );
and \U$6935 ( \15747_16049 , RIe1453f8_2165, \9128_9427 );
and \U$6936 ( \15748_16050 , RIee33b80_5047, \9130_9429 );
and \U$6937 ( \15749_16051 , RIee32938_5034, \9132_9431 );
and \U$6938 ( \15750_16052 , RIee316f0_5021, \9134_9433 );
and \U$6939 ( \15751_16053 , RIee30bb0_5013, \9136_9435 );
and \U$6940 ( \15752_16054 , RIe1403d0_2108, \9138_9437 );
and \U$6941 ( \15753_16055 , RIfe93618_8021, \9140_9439 );
and \U$6942 ( \15754_16056 , RIdf3bfb0_2059, \9142_9441 );
and \U$6943 ( \15755_16057 , RIfe934b0_8020, \9144_9443 );
and \U$6944 ( \15756_16058 , RIfcd0d00_7398, \9146_9445 );
and \U$6945 ( \15757_16059 , RIee2ecc0_4991, \9148_9447 );
and \U$6946 ( \15758_16060 , RIee2e720_4987, \9150_9449 );
and \U$6947 ( \15759_16061 , RIee2cb00_4967, \9152_9451 );
and \U$6948 ( \15760_16062 , RIfe93bb8_8025, \9154_9453 );
and \U$6949 ( \15761_16063 , RIdf32938_1952, \9156_9455 );
and \U$6950 ( \15762_16064 , RIdf30340_1925, \9158_9457 );
and \U$6951 ( \15763_16065 , RIdf2e450_1903, \9160_9459 );
or \U$6952 ( \15764_16066 , \15700_16002 , \15701_16003 , \15702_16004 , \15703_16005 , \15704_16006 , \15705_16007 , \15706_16008 , \15707_16009 , \15708_16010 , \15709_16011 , \15710_16012 , \15711_16013 , \15712_16014 , \15713_16015 , \15714_16016 , \15715_16017 , \15716_16018 , \15717_16019 , \15718_16020 , \15719_16021 , \15720_16022 , \15721_16023 , \15722_16024 , \15723_16025 , \15724_16026 , \15725_16027 , \15726_16028 , \15727_16029 , \15728_16030 , \15729_16031 , \15730_16032 , \15731_16033 , \15732_16034 , \15733_16035 , \15734_16036 , \15735_16037 , \15736_16038 , \15737_16039 , \15738_16040 , \15739_16041 , \15740_16042 , \15741_16043 , \15742_16044 , \15743_16045 , \15744_16046 , \15745_16047 , \15746_16048 , \15747_16049 , \15748_16050 , \15749_16051 , \15750_16052 , \15751_16053 , \15752_16054 , \15753_16055 , \15754_16056 , \15755_16057 , \15756_16058 , \15757_16059 , \15758_16060 , \15759_16061 , \15760_16062 , \15761_16063 , \15762_16064 , \15763_16065 );
and \U$6953 ( \15765_16067 , RIee2b048_4948, \9163_9462 );
and \U$6954 ( \15766_16068 , RIee29b30_4933, \9165_9464 );
and \U$6955 ( \15767_16069 , RIfc67148_6195, \9167_9466 );
and \U$6956 ( \15768_16070 , RIfc6fb18_6293, \9169_9468 );
and \U$6957 ( \15769_16071 , RIdf29860_1849, \9171_9470 );
and \U$6958 ( \15770_16072 , RIfe931e0_8018, \9173_9472 );
and \U$6959 ( \15771_16073 , RIfe93348_8019, \9175_9474 );
and \U$6960 ( \15772_16074 , RIfe93078_8017, \9177_9476 );
and \U$6961 ( \15773_16075 , RIfc672b0_6196, \9179_9478 );
and \U$6962 ( \15774_16076 , RIfca8788_6939, \9181_9480 );
and \U$6963 ( \15775_16077 , RIdf22510_1767, \9183_9482 );
and \U$6964 ( \15776_16078 , RIfcea7a0_7690, \9185_9484 );
and \U$6965 ( \15777_16079 , RIdf20ff8_1752, \9187_9486 );
and \U$6966 ( \15778_16080 , RIdf1ecd0_1727, \9189_9488 );
and \U$6967 ( \15779_16081 , RIdf1aab8_1680, \9191_9490 );
and \U$6968 ( \15780_16082 , RIfea7c58_8225, \9193_9492 );
and \U$6969 ( \15781_16083 , RIdf15ec8_1626, \9195_9494 );
and \U$6970 ( \15782_16084 , RIdf131c8_1594, \9197_9496 );
and \U$6971 ( \15783_16085 , RIdf104c8_1562, \9199_9498 );
and \U$6972 ( \15784_16086 , RIdf0d7c8_1530, \9201_9500 );
and \U$6973 ( \15785_16087 , RIdf0aac8_1498, \9203_9502 );
and \U$6974 ( \15786_16088 , RIdf07dc8_1466, \9205_9504 );
and \U$6975 ( \15787_16089 , RIdf050c8_1434, \9207_9506 );
and \U$6976 ( \15788_16090 , RIdf023c8_1402, \9209_9508 );
and \U$6977 ( \15789_16091 , RIdefc9c8_1338, \9211_9510 );
and \U$6978 ( \15790_16092 , RIdef9cc8_1306, \9213_9512 );
and \U$6979 ( \15791_16093 , RIdef6fc8_1274, \9215_9514 );
and \U$6980 ( \15792_16094 , RIdef42c8_1242, \9217_9516 );
and \U$6981 ( \15793_16095 , RIdef15c8_1210, \9219_9518 );
and \U$6982 ( \15794_16096 , RIdeee8c8_1178, \9221_9520 );
and \U$6983 ( \15795_16097 , RIdeebbc8_1146, \9223_9522 );
and \U$6984 ( \15796_16098 , RIdee8ec8_1114, \9225_9524 );
and \U$6985 ( \15797_16099 , RIee24f40_4879, \9227_9526 );
and \U$6986 ( \15798_16100 , RIee24130_4869, \9229_9528 );
and \U$6987 ( \15799_16101 , RIee235f0_4861, \9231_9530 );
and \U$6988 ( \15800_16102 , RIee22c18_4854, \9233_9532 );
and \U$6989 ( \15801_16103 , RIfe93d20_8026, \9235_9534 );
and \U$6990 ( \15802_16104 , RIdee1fb0_1035, \9237_9536 );
and \U$6991 ( \15803_16105 , RIdee0228_1014, \9239_9538 );
and \U$6992 ( \15804_16106 , RIdeddc30_987, \9241_9540 );
and \U$6993 ( \15805_16107 , RIfc684f8_6209, \9243_9542 );
and \U$6994 ( \15806_16108 , RIee21ca0_4843, \9245_9544 );
and \U$6995 ( \15807_16109 , RIfc68390_6208, \9247_9546 );
and \U$6996 ( \15808_16110 , RIee20d28_4832, \9249_9548 );
and \U$6997 ( \15809_16111 , RIded8aa0_929, \9251_9550 );
and \U$6998 ( \15810_16112 , RIfe93ff0_8028, \9253_9552 );
and \U$6999 ( \15811_16113 , RIded45b8_880, \9255_9554 );
and \U$7000 ( \15812_16114 , RIfe93e88_8027, \9257_9556 );
and \U$7001 ( \15813_16115 , RIdecf6f8_824, \9259_9558 );
and \U$7002 ( \15814_16116 , RIdecc9f8_792, \9261_9560 );
and \U$7003 ( \15815_16117 , RIdec9cf8_760, \9263_9562 );
and \U$7004 ( \15816_16118 , RIdec6ff8_728, \9265_9564 );
and \U$7005 ( \15817_16119 , RIdeb34f8_504, \9267_9566 );
and \U$7006 ( \15818_16120 , RIde941c0_312, \9269_9568 );
and \U$7007 ( \15819_16121 , RIe16d100_2618, \9271_9570 );
and \U$7008 ( \15820_16122 , RIe158ef8_2389, \9273_9572 );
and \U$7009 ( \15821_16123 , RIe1426f8_2133, \9275_9574 );
and \U$7010 ( \15822_16124 , RIdf370f0_2003, \9277_9576 );
and \U$7011 ( \15823_16125 , RIdf2b750_1871, \9279_9578 );
and \U$7012 ( \15824_16126 , RIdf1bfd0_1695, \9281_9580 );
and \U$7013 ( \15825_16127 , RIdeff6c8_1370, \9283_9582 );
and \U$7014 ( \15826_16128 , RIdee61c8_1082, \9285_9584 );
and \U$7015 ( \15827_16129 , RIdedaf30_955, \9287_9586 );
and \U$7016 ( \15828_16130 , RIde7a108_185, \9289_9588 );
or \U$7017 ( \15829_16131 , \15765_16067 , \15766_16068 , \15767_16069 , \15768_16070 , \15769_16071 , \15770_16072 , \15771_16073 , \15772_16074 , \15773_16075 , \15774_16076 , \15775_16077 , \15776_16078 , \15777_16079 , \15778_16080 , \15779_16081 , \15780_16082 , \15781_16083 , \15782_16084 , \15783_16085 , \15784_16086 , \15785_16087 , \15786_16088 , \15787_16089 , \15788_16090 , \15789_16091 , \15790_16092 , \15791_16093 , \15792_16094 , \15793_16095 , \15794_16096 , \15795_16097 , \15796_16098 , \15797_16099 , \15798_16100 , \15799_16101 , \15800_16102 , \15801_16103 , \15802_16104 , \15803_16105 , \15804_16106 , \15805_16107 , \15806_16108 , \15807_16109 , \15808_16110 , \15809_16111 , \15810_16112 , \15811_16113 , \15812_16114 , \15813_16115 , \15814_16116 , \15815_16117 , \15816_16118 , \15817_16119 , \15818_16120 , \15819_16121 , \15820_16122 , \15821_16123 , \15822_16124 , \15823_16125 , \15824_16126 , \15825_16127 , \15826_16128 , \15827_16129 , \15828_16130 );
or \U$7018 ( \15830_16132 , \15764_16066 , \15829_16131 );
_DC \g6595/U$1 ( \15831 , \15830_16132 , \9298_9597 );
and \U$7019 ( \15832_16134 , RIe19c590_3156, \8760_9059 );
and \U$7020 ( \15833_16135 , RIe199890_3124, \8762_9061 );
and \U$7021 ( \15834_16136 , RIf144f50_5244, \8764_9063 );
and \U$7022 ( \15835_16137 , RIe196b90_3092, \8766_9065 );
and \U$7023 ( \15836_16138 , RIfc76058_6365, \8768_9067 );
and \U$7024 ( \15837_16139 , RIe193e90_3060, \8770_9069 );
and \U$7025 ( \15838_16140 , RIe191190_3028, \8772_9071 );
and \U$7026 ( \15839_16141 , RIe18e490_2996, \8774_9073 );
and \U$7027 ( \15840_16142 , RIe188a90_2932, \8776_9075 );
and \U$7028 ( \15841_16143 , RIe185d90_2900, \8778_9077 );
and \U$7029 ( \15842_16144 , RIfccd8f8_7361, \8780_9079 );
and \U$7030 ( \15843_16145 , RIe183090_2868, \8782_9081 );
and \U$7031 ( \15844_16146 , RIfc76e68_6375, \8784_9083 );
and \U$7032 ( \15845_16147 , RIe180390_2836, \8786_9085 );
and \U$7033 ( \15846_16148 , RIe17d690_2804, \8788_9087 );
and \U$7034 ( \15847_16149 , RIe17a990_2772, \8790_9089 );
and \U$7035 ( \15848_16150 , RIf1419e0_5206, \8792_9091 );
and \U$7036 ( \15849_16151 , RIf140630_5192, \8794_9093 );
and \U$7037 ( \15850_16152 , RIe176bb0_2728, \8796_9095 );
and \U$7038 ( \15851_16153 , RIe1750f8_2709, \8798_9097 );
and \U$7039 ( \15852_16154 , RIfcd1840_7406, \8800_9099 );
and \U$7040 ( \15853_16155 , RIfc5f6f0_6108, \8802_9101 );
and \U$7041 ( \15854_16156 , RIee3dd38_5162, \8804_9103 );
and \U$7042 ( \15855_16157 , RIee3cc58_5150, \8806_9105 );
and \U$7043 ( \15856_16158 , RIee3b8a8_5136, \8808_9107 );
and \U$7044 ( \15857_16159 , RIee3a7c8_5124, \8810_9109 );
and \U$7045 ( \15858_16160 , RIee39580_5111, \8812_9111 );
and \U$7046 ( \15859_16161 , RIfea9008_8239, \8814_9113 );
and \U$7047 ( \15860_16162 , RIf16f7f0_5728, \8816_9115 );
and \U$7048 ( \15861_16163 , RIf16ecb0_5720, \8818_9117 );
and \U$7049 ( \15862_16164 , RIf16d900_5706, \8820_9119 );
and \U$7050 ( \15863_16165 , RIfc78ec0_6398, \8822_9121 );
and \U$7051 ( \15864_16166 , RIfcc8060_7298, \8824_9123 );
and \U$7052 ( \15865_16167 , RIe2228e8_4683, \8826_9125 );
and \U$7053 ( \15866_16168 , RIfc5a3f8_6049, \8828_9127 );
and \U$7054 ( \15867_16169 , RIe21fbe8_4651, \8830_9129 );
and \U$7055 ( \15868_16170 , RIfc74000_6342, \8832_9131 );
and \U$7056 ( \15869_16171 , RIe21cee8_4619, \8834_9133 );
and \U$7057 ( \15870_16172 , RIe2174e8_4555, \8836_9135 );
and \U$7058 ( \15871_16173 , RIe2147e8_4523, \8838_9137 );
and \U$7059 ( \15872_16174 , RIfca2c20_6874, \8840_9139 );
and \U$7060 ( \15873_16175 , RIe211ae8_4491, \8842_9141 );
and \U$7061 ( \15874_16176 , RIfca2950_6872, \8844_9143 );
and \U$7062 ( \15875_16177 , RIe20ede8_4459, \8846_9145 );
and \U$7063 ( \15876_16178 , RIfcc24f8_7233, \8848_9147 );
and \U$7064 ( \15877_16179 , RIe20c0e8_4427, \8850_9149 );
and \U$7065 ( \15878_16180 , RIe2093e8_4395, \8852_9151 );
and \U$7066 ( \15879_16181 , RIe2066e8_4363, \8854_9153 );
and \U$7067 ( \15880_16182 , RIfc45110_5808, \8856_9155 );
and \U$7068 ( \15881_16183 , RIfcc6f80_7286, \8858_9157 );
and \U$7069 ( \15882_16184 , RIfe92f10_8016, \8860_9159 );
and \U$7070 ( \15883_16185 , RIfe92970_8012, \8862_9161 );
and \U$7071 ( \15884_16186 , RIf164af8_5605, \8864_9163 );
and \U$7072 ( \15885_16187 , RIf163a18_5593, \8866_9165 );
and \U$7073 ( \15886_16188 , RIf162aa0_5582, \8868_9167 );
and \U$7074 ( \15887_16189 , RIfe92ad8_8013, \8870_9169 );
and \U$7075 ( \15888_16190 , RIf15f3c8_5543, \8872_9171 );
and \U$7076 ( \15889_16191 , RIf15d640_5522, \8874_9173 );
and \U$7077 ( \15890_16192 , RIfe92808_8011, \8876_9175 );
and \U$7078 ( \15891_16193 , RIfe92c40_8014, \8878_9177 );
and \U$7079 ( \15892_16194 , RIfe926a0_8010, \8880_9179 );
and \U$7080 ( \15893_16195 , RIfe92da8_8015, \8882_9181 );
and \U$7081 ( \15894_16196 , RIfe92538_8009, \8884_9183 );
and \U$7082 ( \15895_16197 , RIfcb5a78_7089, \8886_9185 );
or \U$7083 ( \15896_16198 , \15832_16134 , \15833_16135 , \15834_16136 , \15835_16137 , \15836_16138 , \15837_16139 , \15838_16140 , \15839_16141 , \15840_16142 , \15841_16143 , \15842_16144 , \15843_16145 , \15844_16146 , \15845_16147 , \15846_16148 , \15847_16149 , \15848_16150 , \15849_16151 , \15850_16152 , \15851_16153 , \15852_16154 , \15853_16155 , \15854_16156 , \15855_16157 , \15856_16158 , \15857_16159 , \15858_16160 , \15859_16161 , \15860_16162 , \15861_16163 , \15862_16164 , \15863_16165 , \15864_16166 , \15865_16167 , \15866_16168 , \15867_16169 , \15868_16170 , \15869_16171 , \15870_16172 , \15871_16173 , \15872_16174 , \15873_16175 , \15874_16176 , \15875_16177 , \15876_16178 , \15877_16179 , \15878_16180 , \15879_16181 , \15880_16182 , \15881_16183 , \15882_16184 , \15883_16185 , \15884_16186 , \15885_16187 , \15886_16188 , \15887_16189 , \15888_16190 , \15889_16191 , \15890_16192 , \15891_16193 , \15892_16194 , \15893_16195 , \15894_16196 , \15895_16197 );
and \U$7084 ( \15897_16199 , RIf158348_5463, \8889_9188 );
and \U$7085 ( \15898_16200 , RIf157100_5450, \8891_9190 );
and \U$7086 ( \15899_16201 , RIfc53be8_5975, \8893_9192 );
and \U$7087 ( \15900_16202 , RIfec38b8_8345, \8895_9194 );
and \U$7088 ( \15901_16203 , RIfcc5ea0_7274, \8897_9196 );
and \U$7089 ( \15902_16204 , RIf1550a8_5427, \8899_9198 );
and \U$7090 ( \15903_16205 , RIf153cf8_5413, \8901_9200 );
and \U$7091 ( \15904_16206 , RIfec3a20_8346, \8903_9202 );
and \U$7092 ( \15905_16207 , RIf152678_5397, \8905_9204 );
and \U$7093 ( \15906_16208 , RIfec3750_8344, \8907_9206 );
and \U$7094 ( \15907_16209 , RIf14ff18_5369, \8909_9208 );
and \U$7095 ( \15908_16210 , RIfe923d0_8008, \8911_9210 );
and \U$7096 ( \15909_16211 , RIf14efa0_5358, \8913_9212 );
and \U$7097 ( \15910_16212 , RIf14e898_5353, \8915_9214 );
and \U$7098 ( \15911_16213 , RIf14d380_5338, \8917_9216 );
and \U$7099 ( \15912_16214 , RIfe92268_8007, \8919_9218 );
and \U$7100 ( \15913_16215 , RIe1ea650_4044, \8921_9220 );
and \U$7101 ( \15914_16216 , RIe1e7950_4012, \8923_9222 );
and \U$7102 ( \15915_16217 , RIe1e4c50_3980, \8925_9224 );
and \U$7103 ( \15916_16218 , RIe1e1f50_3948, \8927_9226 );
and \U$7104 ( \15917_16219 , RIe1df250_3916, \8929_9228 );
and \U$7105 ( \15918_16220 , RIe1dc550_3884, \8931_9230 );
and \U$7106 ( \15919_16221 , RIe1d9850_3852, \8933_9232 );
and \U$7107 ( \15920_16222 , RIe1d6b50_3820, \8935_9234 );
and \U$7108 ( \15921_16223 , RIe1d1150_3756, \8937_9236 );
and \U$7109 ( \15922_16224 , RIe1ce450_3724, \8939_9238 );
and \U$7110 ( \15923_16225 , RIe1cb750_3692, \8941_9240 );
and \U$7111 ( \15924_16226 , RIe1c8a50_3660, \8943_9242 );
and \U$7112 ( \15925_16227 , RIe1c5d50_3628, \8945_9244 );
and \U$7113 ( \15926_16228 , RIe1c3050_3596, \8947_9246 );
and \U$7114 ( \15927_16229 , RIe1c0350_3564, \8949_9248 );
and \U$7115 ( \15928_16230 , RIe1bd650_3532, \8951_9250 );
and \U$7116 ( \15929_16231 , RIfcda4e0_7506, \8953_9252 );
and \U$7117 ( \15930_16232 , RIfc9d220_6810, \8955_9254 );
and \U$7118 ( \15931_16233 , RIe1b8628_3475, \8957_9256 );
and \U$7119 ( \15932_16234 , RIe1b6738_3453, \8959_9258 );
and \U$7120 ( \15933_16235 , RIfc4f2c8_5923, \8961_9260 );
and \U$7121 ( \15934_16236 , RIfce16c8_7587, \8963_9262 );
and \U$7122 ( \15935_16237 , RIfe91cc8_8003, \8965_9264 );
and \U$7123 ( \15936_16238 , RIfe91e30_8004, \8967_9266 );
and \U$7124 ( \15937_16239 , RIf1484c0_5282, \8969_9268 );
and \U$7125 ( \15938_16240 , RIf147548_5271, \8971_9270 );
and \U$7126 ( \15939_16241 , RIfe91f98_8005, \8973_9272 );
and \U$7127 ( \15940_16242 , RIfe91b60_8002, \8975_9274 );
and \U$7128 ( \15941_16243 , RIf146b70_5264, \8977_9276 );
and \U$7129 ( \15942_16244 , RIfc9f548_6835, \8979_9278 );
and \U$7130 ( \15943_16245 , RIfe92100_8006, \8981_9280 );
and \U$7131 ( \15944_16246 , RIfe919f8_8001, \8983_9282 );
and \U$7132 ( \15945_16247 , RIe1a7990_3284, \8985_9284 );
and \U$7133 ( \15946_16248 , RIe1a4c90_3252, \8987_9286 );
and \U$7134 ( \15947_16249 , RIe1a1f90_3220, \8989_9288 );
and \U$7135 ( \15948_16250 , RIe19f290_3188, \8991_9290 );
and \U$7136 ( \15949_16251 , RIe18b790_2964, \8993_9292 );
and \U$7137 ( \15950_16252 , RIe177c90_2740, \8995_9294 );
and \U$7138 ( \15951_16253 , RIe2255e8_4715, \8997_9296 );
and \U$7139 ( \15952_16254 , RIe21a1e8_4587, \8999_9298 );
and \U$7140 ( \15953_16255 , RIe2039e8_4331, \9001_9300 );
and \U$7141 ( \15954_16256 , RIe1fda48_4263, \9003_9302 );
and \U$7142 ( \15955_16257 , RIe1f6e00_4186, \9005_9304 );
and \U$7143 ( \15956_16258 , RIe1ef948_4103, \9007_9306 );
and \U$7144 ( \15957_16259 , RIe1d3e50_3788, \9009_9308 );
and \U$7145 ( \15958_16260 , RIe1ba950_3500, \9011_9310 );
and \U$7146 ( \15959_16261 , RIe1ad7c8_3351, \9013_9312 );
and \U$7147 ( \15960_16262 , RIe16fe00_2650, \9015_9314 );
or \U$7148 ( \15961_16263 , \15897_16199 , \15898_16200 , \15899_16201 , \15900_16202 , \15901_16203 , \15902_16204 , \15903_16205 , \15904_16206 , \15905_16207 , \15906_16208 , \15907_16209 , \15908_16210 , \15909_16211 , \15910_16212 , \15911_16213 , \15912_16214 , \15913_16215 , \15914_16216 , \15915_16217 , \15916_16218 , \15917_16219 , \15918_16220 , \15919_16221 , \15920_16222 , \15921_16223 , \15922_16224 , \15923_16225 , \15924_16226 , \15925_16227 , \15926_16228 , \15927_16229 , \15928_16230 , \15929_16231 , \15930_16232 , \15931_16233 , \15932_16234 , \15933_16235 , \15934_16236 , \15935_16237 , \15936_16238 , \15937_16239 , \15938_16240 , \15939_16241 , \15940_16242 , \15941_16243 , \15942_16244 , \15943_16245 , \15944_16246 , \15945_16247 , \15946_16248 , \15947_16249 , \15948_16250 , \15949_16251 , \15950_16252 , \15951_16253 , \15952_16254 , \15953_16255 , \15954_16256 , \15955_16257 , \15956_16258 , \15957_16259 , \15958_16260 , \15959_16261 , \15960_16262 );
or \U$7149 ( \15962_16264 , \15896_16198 , \15961_16263 );
_DC \g6596/U$1 ( \15963 , \15962_16264 , \9024_9323 );
and g6597_GF_PartitionCandidate( \15964_16266_nG6597 , \15831 , \15963 );
buf \U$7150 ( \15965_16267 , \15964_16266_nG6597 );
and \U$7151 ( \15966_16268 , \15965_16267 , \10389_10691 );
nor \U$7152 ( \15967_16269 , \15699_16001 , \15966_16268 );
xnor \U$7153 ( \15968_16270 , \15967_16269 , \10678_10980 );
and \U$7154 ( \15969_16271 , \12470_12769 , \12491_12790 );
and \U$7155 ( \15970_16272 , \13377_13679 , \12159_12461 );
nor \U$7156 ( \15971_16273 , \15969_16271 , \15970_16272 );
xnor \U$7157 ( \15972_16274 , \15971_16273 , \12481_12780 );
xor \U$7158 ( \15973_16275 , \15968_16270 , \15972_16274 );
and \U$7159 ( \15974_16276 , \10686_10988 , \15037_15336 );
and \U$7160 ( \15975_16277 , \10968_11270 , \14661_14963 );
nor \U$7161 ( \15976_16278 , \15974_16276 , \15975_16277 );
xnor \U$7162 ( \15977_16279 , \15976_16278 , \15043_15342 );
xor \U$7163 ( \15978_16280 , \15973_16275 , \15977_16279 );
xor \U$7164 ( \15979_16281 , \15698_16000 , \15978_16280 );
and \U$7165 ( \15980_16282 , \15025_15324 , \15029_15328 );
and \U$7166 ( \15981_16283 , \15029_15328 , \15044_15343 );
and \U$7167 ( \15982_16284 , \15025_15324 , \15044_15343 );
or \U$7168 ( \15983_16285 , \15980_16282 , \15981_16283 , \15982_16284 );
and \U$7169 ( \15984_16286 , \15050_15349 , \15052_15351 );
xor \U$7170 ( \15985_16287 , \15983_16285 , \15984_16286 );
and \U$7171 ( \15986_16288 , \13725_14024 , \11275_11574 );
and \U$7172 ( \15987_16289 , \14648_14950 , \10976_11278 );
nor \U$7173 ( \15988_16290 , \15986_16288 , \15987_16289 );
xnor \U$7174 ( \15989_16291 , \15988_16290 , \11281_11580 );
and \U$7175 ( \15990_16292 , \11287_11586 , \13755_14054 );
and \U$7176 ( \15991_16293 , \12146_12448 , \13390_13692 );
nor \U$7177 ( \15992_16294 , \15990_16292 , \15991_16293 );
xnor \U$7178 ( \15993_16295 , \15992_16294 , \13736_14035 );
xor \U$7179 ( \15994_16296 , \15989_16291 , \15993_16295 );
_DC \g4f34/U$1 ( \15995 , \15830_16132 , \9298_9597 );
_DC \g4fb8/U$1 ( \15996 , \15962_16264 , \9024_9323 );
xor g4fb9_GF_PartitionCandidate( \15997_16299_nG4fb9 , \15995 , \15996 );
buf \U$7180 ( \15998_16300 , \15997_16299_nG4fb9 );
xor \U$7181 ( \15999_16301 , \15998_16300 , \15034_15333 );
and \U$7182 ( \16000_16302 , \10385_10687 , \15999_16301 );
xor \U$7183 ( \16001_16303 , \15994_16296 , \16000_16302 );
xor \U$7184 ( \16002_16304 , \15985_16287 , \16001_16303 );
xor \U$7185 ( \16003_16305 , \15979_16281 , \16002_16304 );
and \U$7186 ( \16004_16306 , \14755_15054 , \15045_15344 );
and \U$7187 ( \16005_16307 , \15045_15344 , \15063_15362 );
and \U$7188 ( \16006_16308 , \14755_15054 , \15063_15362 );
or \U$7189 ( \16007_16309 , \16004_16306 , \16005_16307 , \16006_16308 );
xor \U$7190 ( \16008_16310 , \16003_16305 , \16007_16309 );
and \U$7191 ( \16009_16311 , \15064_15363 , \15068_15367 );
and \U$7192 ( \16010_16312 , \15069_15368 , \15072_15371 );
or \U$7193 ( \16011_16313 , \16009_16311 , \16010_16312 );
xor \U$7194 ( \16012_16314 , \16008_16310 , \16011_16313 );
buf g9bf0_GF_PartitionCandidate( \16013_16315_nG9bf0 , \16012_16314 );
and \U$7195 ( \16014_16316 , \10402_10704 , \16013_16315_nG9bf0 );
or \U$7196 ( \16015_16317 , \15694_15996 , \16014_16316 );
xor \U$7197 ( \16016_16318 , \10399_10703 , \16015_16317 );
buf \U$7198 ( \16017_16319 , \16016_16318 );
buf \U$7200 ( \16018_16320 , \16017_16319 );
xor \U$7201 ( \16019_16321 , \15693_15995 , \16018_16320 );
buf \U$7202 ( \16020_16322 , \16019_16321 );
xor \U$7203 ( \16021_16323 , \15681_15983 , \16020_16322 );
buf \U$7204 ( \16022_16324 , \16021_16323 );
xor \U$7205 ( \16023_16325 , \15650_15952 , \16022_16324 );
and \U$7206 ( \16024_16326 , \14704_15006 , \15081_15380 );
and \U$7207 ( \16025_16327 , \14704_15006 , \15087_15386 );
and \U$7208 ( \16026_16328 , \15081_15380 , \15087_15386 );
or \U$7209 ( \16027_16329 , \16024_16326 , \16025_16327 , \16026_16328 );
buf \U$7210 ( \16028_16330 , \16027_16329 );
xor \U$7211 ( \16029_16331 , \16023_16325 , \16028_16330 );
and \U$7212 ( \16030_16332 , \15089_15388 , \16029_16331 );
and \U$7213 ( \16031_16333 , \15644_15946 , \16029_16331 );
or \U$7214 ( \16032_16334 , \15645_15947 , \16030_16332 , \16031_16333 );
and \U$7215 ( \16033_16335 , \15669_15971 , \15671_15973 );
and \U$7216 ( \16034_16336 , \15669_15971 , \15678_15980 );
and \U$7217 ( \16035_16337 , \15671_15973 , \15678_15980 );
or \U$7218 ( \16036_16338 , \16033_16335 , \16034_16336 , \16035_16337 );
buf \U$7219 ( \16037_16339 , \16036_16338 );
and \U$7220 ( \16038_16340 , \10996_10421 , \14682_14984_nG9bf6 );
and \U$7221 ( \16039_16341 , \10119_10418 , \15074_15373_nG9bf3 );
or \U$7222 ( \16040_16342 , \16038_16340 , \16039_16341 );
xor \U$7223 ( \16041_16343 , \10118_10417 , \16040_16342 );
buf \U$7224 ( \16042_16344 , \16041_16343 );
buf \U$7226 ( \16043_16345 , \16042_16344 );
xor \U$7227 ( \16044_16346 , \16037_16339 , \16043_16345 );
and \U$7228 ( \16045_16347 , \10411_10707 , \16013_16315_nG9bf0 );
and \U$7229 ( \16046_16348 , \15983_16285 , \15984_16286 );
and \U$7230 ( \16047_16349 , \15984_16286 , \16001_16303 );
and \U$7231 ( \16048_16350 , \15983_16285 , \16001_16303 );
or \U$7232 ( \16049_16351 , \16046_16348 , \16047_16349 , \16048_16350 );
and \U$7233 ( \16050_16352 , \14648_14950 , \11275_11574 );
and \U$7234 ( \16051_16353 , \15022_15321 , \10976_11278 );
nor \U$7235 ( \16052_16354 , \16050_16352 , \16051_16353 );
xnor \U$7236 ( \16053_16355 , \16052_16354 , \11281_11580 );
not \U$7237 ( \16054_16356 , \16000_16302 );
and \U$7238 ( \16055_16357 , RIdec4460_697, \9034_9333 );
and \U$7239 ( \16056_16358 , RIdec1760_665, \9036_9335 );
and \U$7240 ( \16057_16359 , RIee1fae0_4819, \9038_9337 );
and \U$7241 ( \16058_16360 , RIdebea60_633, \9040_9339 );
and \U$7242 ( \16059_16361 , RIee1f108_4812, \9042_9341 );
and \U$7243 ( \16060_16362 , RIdebbd60_601, \9044_9343 );
and \U$7244 ( \16061_16363 , RIdeb9060_569, \9046_9345 );
and \U$7245 ( \16062_16364 , RIdeb6360_537, \9048_9347 );
and \U$7246 ( \16063_16365 , RIee1eb68_4808, \9050_9349 );
and \U$7247 ( \16064_16366 , RIdeb0960_473, \9052_9351 );
and \U$7248 ( \16065_16367 , RIee1e460_4803, \9054_9353 );
and \U$7249 ( \16066_16368 , RIdeadc60_441, \9056_9355 );
and \U$7250 ( \16067_16369 , RIee1d7b8_4794, \9058_9357 );
and \U$7251 ( \16068_16370 , RIdea8008_409, \9060_9359 );
and \U$7252 ( \16069_16371 , RIdea1708_377, \9062_9361 );
and \U$7253 ( \16070_16372 , RIde9ae08_345, \9064_9363 );
and \U$7254 ( \16071_16373 , RIfe957d8_8045, \9066_9365 );
and \U$7255 ( \16072_16374 , RIfe95508_8043, \9068_9367 );
and \U$7256 ( \16073_16375 , RIfe95670_8044, \9070_9369 );
and \U$7257 ( \16074_16376 , RIee1a7e8_4760, \9072_9371 );
and \U$7258 ( \16075_16377 , RIfe95aa8_8047, \9074_9373 );
and \U$7259 ( \16076_16378 , RIfe95238_8041, \9076_9375 );
and \U$7260 ( \16077_16379 , RIfe95940_8046, \9078_9377 );
and \U$7261 ( \16078_16380 , RIfe953a0_8042, \9080_9379 );
and \U$7262 ( \16079_16381 , RIee1a0e0_4755, \9082_9381 );
and \U$7263 ( \16080_16382 , RIee19ca8_4752, \9084_9383 );
and \U$7264 ( \16081_16383 , RIee19870_4749, \9086_9385 );
and \U$7265 ( \16082_16384 , RIee19438_4746, \9088_9387 );
and \U$7266 ( \16083_16385 , RIee38ba8_5104, \9090_9389 );
and \U$7267 ( \16084_16386 , RIfe95c10_8048, \9092_9391 );
and \U$7268 ( \16085_16387 , RIee384a0_5099, \9094_9393 );
and \U$7269 ( \16086_16388 , RIfea9440_8242, \9096_9395 );
and \U$7270 ( \16087_16389 , RIe164460_2518, \9098_9397 );
and \U$7271 ( \16088_16390 , RIe161760_2486, \9100_9399 );
and \U$7272 ( \16089_16391 , RIfe942c0_8030, \9102_9401 );
and \U$7273 ( \16090_16392 , RIe15ea60_2454, \9104_9403 );
and \U$7274 ( \16091_16393 , RIfe94158_8029, \9106_9405 );
and \U$7275 ( \16092_16394 , RIe15bd60_2422, \9108_9407 );
and \U$7276 ( \16093_16395 , RIe156360_2358, \9110_9409 );
and \U$7277 ( \16094_16396 , RIe153660_2326, \9112_9411 );
and \U$7278 ( \16095_16397 , RIfe94428_8031, \9114_9413 );
and \U$7279 ( \16096_16398 , RIe150960_2294, \9116_9415 );
and \U$7280 ( \16097_16399 , RIfe94590_8032, \9118_9417 );
and \U$7281 ( \16098_16400 , RIe14dc60_2262, \9120_9419 );
and \U$7282 ( \16099_16401 , RIfc5c2e8_6071, \9122_9421 );
and \U$7283 ( \16100_16402 , RIe14af60_2230, \9124_9423 );
and \U$7284 ( \16101_16403 , RIe148260_2198, \9126_9425 );
and \U$7285 ( \16102_16404 , RIe145560_2166, \9128_9427 );
and \U$7286 ( \16103_16405 , RIee33ce8_5048, \9130_9429 );
and \U$7287 ( \16104_16406 , RIee32aa0_5035, \9132_9431 );
and \U$7288 ( \16105_16407 , RIee31858_5022, \9134_9433 );
and \U$7289 ( \16106_16408 , RIfc5d530_6084, \9136_9435 );
and \U$7290 ( \16107_16409 , RIe140538_2109, \9138_9437 );
and \U$7291 ( \16108_16410 , RIdf3e2d8_2084, \9140_9439 );
and \U$7292 ( \16109_16411 , RIdf3c118_2060, \9142_9441 );
and \U$7293 ( \16110_16412 , RIdf39df0_2035, \9144_9443 );
and \U$7294 ( \16111_16413 , RIfcdd780_7542, \9146_9445 );
and \U$7295 ( \16112_16414 , RIee2ee28_4992, \9148_9447 );
and \U$7296 ( \16113_16415 , RIfcc88d0_7304, \9150_9449 );
and \U$7297 ( \16114_16416 , RIee2cc68_4968, \9152_9451 );
and \U$7298 ( \16115_16417 , RIdf34990_1975, \9154_9453 );
and \U$7299 ( \16116_16418 , RIdf32aa0_1953, \9156_9455 );
and \U$7300 ( \16117_16419 , RIdf304a8_1926, \9158_9457 );
and \U$7301 ( \16118_16420 , RIdf2e5b8_1904, \9160_9459 );
or \U$7302 ( \16119_16421 , \16055_16357 , \16056_16358 , \16057_16359 , \16058_16360 , \16059_16361 , \16060_16362 , \16061_16363 , \16062_16364 , \16063_16365 , \16064_16366 , \16065_16367 , \16066_16368 , \16067_16369 , \16068_16370 , \16069_16371 , \16070_16372 , \16071_16373 , \16072_16374 , \16073_16375 , \16074_16376 , \16075_16377 , \16076_16378 , \16077_16379 , \16078_16380 , \16079_16381 , \16080_16382 , \16081_16383 , \16082_16384 , \16083_16385 , \16084_16386 , \16085_16387 , \16086_16388 , \16087_16389 , \16088_16390 , \16089_16391 , \16090_16392 , \16091_16393 , \16092_16394 , \16093_16395 , \16094_16396 , \16095_16397 , \16096_16398 , \16097_16399 , \16098_16400 , \16099_16401 , \16100_16402 , \16101_16403 , \16102_16404 , \16103_16405 , \16104_16406 , \16105_16407 , \16106_16408 , \16107_16409 , \16108_16410 , \16109_16411 , \16110_16412 , \16111_16413 , \16112_16414 , \16113_16415 , \16114_16416 , \16115_16417 , \16116_16418 , \16117_16419 , \16118_16420 );
and \U$7303 ( \16120_16422 , RIee2b1b0_4949, \9163_9462 );
and \U$7304 ( \16121_16423 , RIfe946f8_8033, \9165_9464 );
and \U$7305 ( \16122_16424 , RIfcb2940_7054, \9167_9466 );
and \U$7306 ( \16123_16425 , RIee273d0_4905, \9169_9468 );
and \U$7307 ( \16124_16426 , RIfe949c8_8035, \9171_9470 );
and \U$7308 ( \16125_16427 , RIdf27538_1824, \9173_9472 );
and \U$7309 ( \16126_16428 , RIfe94b30_8036, \9175_9474 );
and \U$7310 ( \16127_16429 , RIfe94860_8034, \9177_9476 );
and \U$7311 ( \16128_16430 , RIee26f98_4902, \9179_9478 );
and \U$7312 ( \16129_16431 , RIee269f8_4898, \9181_9480 );
and \U$7313 ( \16130_16432 , RIee26728_4896, \9183_9482 );
and \U$7314 ( \16131_16433 , RIee26458_4894, \9185_9484 );
and \U$7315 ( \16132_16434 , RIee26188_4892, \9187_9486 );
and \U$7316 ( \16133_16435 , RIfe94c98_8037, \9189_9488 );
and \U$7317 ( \16134_16436 , RIee25d50_4889, \9191_9490 );
and \U$7318 ( \16135_16437 , RIfea9170_8240, \9193_9492 );
and \U$7319 ( \16136_16438 , RIdf16030_1627, \9195_9494 );
and \U$7320 ( \16137_16439 , RIdf13330_1595, \9197_9496 );
and \U$7321 ( \16138_16440 , RIdf10630_1563, \9199_9498 );
and \U$7322 ( \16139_16441 , RIdf0d930_1531, \9201_9500 );
and \U$7323 ( \16140_16442 , RIdf0ac30_1499, \9203_9502 );
and \U$7324 ( \16141_16443 , RIdf07f30_1467, \9205_9504 );
and \U$7325 ( \16142_16444 , RIdf05230_1435, \9207_9506 );
and \U$7326 ( \16143_16445 , RIdf02530_1403, \9209_9508 );
and \U$7327 ( \16144_16446 , RIdefcb30_1339, \9211_9510 );
and \U$7328 ( \16145_16447 , RIdef9e30_1307, \9213_9512 );
and \U$7329 ( \16146_16448 , RIdef7130_1275, \9215_9514 );
and \U$7330 ( \16147_16449 , RIdef4430_1243, \9217_9516 );
and \U$7331 ( \16148_16450 , RIdef1730_1211, \9219_9518 );
and \U$7332 ( \16149_16451 , RIdeeea30_1179, \9221_9520 );
and \U$7333 ( \16150_16452 , RIdeebd30_1147, \9223_9522 );
and \U$7334 ( \16151_16453 , RIdee9030_1115, \9225_9524 );
and \U$7335 ( \16152_16454 , RIee250a8_4880, \9227_9526 );
and \U$7336 ( \16153_16455 , RIee24298_4870, \9229_9528 );
and \U$7337 ( \16154_16456 , RIee23758_4862, \9231_9530 );
and \U$7338 ( \16155_16457 , RIee22d80_4855, \9233_9532 );
and \U$7339 ( \16156_16458 , RIfe950d0_8040, \9235_9534 );
and \U$7340 ( \16157_16459 , RIfe94f68_8039, \9237_9536 );
and \U$7341 ( \16158_16460 , RIfe94e00_8038, \9239_9538 );
and \U$7342 ( \16159_16461 , RIdeddd98_988, \9241_9540 );
and \U$7343 ( \16160_16462 , RIee22ab0_4853, \9243_9542 );
and \U$7344 ( \16161_16463 , RIee21e08_4844, \9245_9544 );
and \U$7345 ( \16162_16464 , RIfca46d8_6893, \9247_9546 );
and \U$7346 ( \16163_16465 , RIfc5dad0_6088, \9249_9548 );
and \U$7347 ( \16164_16466 , RIfeaa250_8252, \9251_9550 );
and \U$7348 ( \16165_16467 , RIfe96048_8051, \9253_9552 );
and \U$7349 ( \16166_16468 , RIfe95d78_8049, \9255_9554 );
and \U$7350 ( \16167_16469 , RIfe95ee0_8050, \9257_9556 );
and \U$7351 ( \16168_16470 , RIdecf860_825, \9259_9558 );
and \U$7352 ( \16169_16471 , RIdeccb60_793, \9261_9560 );
and \U$7353 ( \16170_16472 , RIdec9e60_761, \9263_9562 );
and \U$7354 ( \16171_16473 , RIdec7160_729, \9265_9564 );
and \U$7355 ( \16172_16474 , RIdeb3660_505, \9267_9566 );
and \U$7356 ( \16173_16475 , RIde94508_313, \9269_9568 );
and \U$7357 ( \16174_16476 , RIe16d268_2619, \9271_9570 );
and \U$7358 ( \16175_16477 , RIe159060_2390, \9273_9572 );
and \U$7359 ( \16176_16478 , RIe142860_2134, \9275_9574 );
and \U$7360 ( \16177_16479 , RIdf37258_2004, \9277_9576 );
and \U$7361 ( \16178_16480 , RIdf2b8b8_1872, \9279_9578 );
and \U$7362 ( \16179_16481 , RIdf1c138_1696, \9281_9580 );
and \U$7363 ( \16180_16482 , RIdeff830_1371, \9283_9582 );
and \U$7364 ( \16181_16483 , RIdee6330_1083, \9285_9584 );
and \U$7365 ( \16182_16484 , RIdedb098_956, \9287_9586 );
and \U$7366 ( \16183_16485 , RIde7a450_186, \9289_9588 );
or \U$7367 ( \16184_16486 , \16120_16422 , \16121_16423 , \16122_16424 , \16123_16425 , \16124_16426 , \16125_16427 , \16126_16428 , \16127_16429 , \16128_16430 , \16129_16431 , \16130_16432 , \16131_16433 , \16132_16434 , \16133_16435 , \16134_16436 , \16135_16437 , \16136_16438 , \16137_16439 , \16138_16440 , \16139_16441 , \16140_16442 , \16141_16443 , \16142_16444 , \16143_16445 , \16144_16446 , \16145_16447 , \16146_16448 , \16147_16449 , \16148_16450 , \16149_16451 , \16150_16452 , \16151_16453 , \16152_16454 , \16153_16455 , \16154_16456 , \16155_16457 , \16156_16458 , \16157_16459 , \16158_16460 , \16159_16461 , \16160_16462 , \16161_16463 , \16162_16464 , \16163_16465 , \16164_16466 , \16165_16467 , \16166_16468 , \16167_16469 , \16168_16470 , \16169_16471 , \16170_16472 , \16171_16473 , \16172_16474 , \16173_16475 , \16174_16476 , \16175_16477 , \16176_16478 , \16177_16479 , \16178_16480 , \16179_16481 , \16180_16482 , \16181_16483 , \16182_16484 , \16183_16485 );
or \U$7368 ( \16185_16487 , \16119_16421 , \16184_16486 );
_DC \g503d/U$1 ( \16186 , \16185_16487 , \9298_9597 );
and \U$7369 ( \16187_16489 , RIe19c6f8_3157, \8760_9059 );
and \U$7370 ( \16188_16490 , RIe1999f8_3125, \8762_9061 );
and \U$7371 ( \16189_16491 , RIf1450b8_5245, \8764_9063 );
and \U$7372 ( \16190_16492 , RIe196cf8_3093, \8766_9065 );
and \U$7373 ( \16191_16493 , RIf143fd8_5233, \8768_9067 );
and \U$7374 ( \16192_16494 , RIe193ff8_3061, \8770_9069 );
and \U$7375 ( \16193_16495 , RIe1912f8_3029, \8772_9071 );
and \U$7376 ( \16194_16496 , RIe18e5f8_2997, \8774_9073 );
and \U$7377 ( \16195_16497 , RIe188bf8_2933, \8776_9075 );
and \U$7378 ( \16196_16498 , RIe185ef8_2901, \8778_9077 );
and \U$7379 ( \16197_16499 , RIfe973f8_8065, \8780_9079 );
and \U$7380 ( \16198_16500 , RIe1831f8_2869, \8782_9081 );
and \U$7381 ( \16199_16501 , RIf142958_5217, \8784_9083 );
and \U$7382 ( \16200_16502 , RIe1804f8_2837, \8786_9085 );
and \U$7383 ( \16201_16503 , RIe17d7f8_2805, \8788_9087 );
and \U$7384 ( \16202_16504 , RIe17aaf8_2773, \8790_9089 );
and \U$7385 ( \16203_16505 , RIf141b48_5207, \8792_9091 );
and \U$7386 ( \16204_16506 , RIfc542f0_5980, \8794_9093 );
and \U$7387 ( \16205_16507 , RIfc800a8_6479, \8796_9095 );
and \U$7388 ( \16206_16508 , RIe175260_2710, \8798_9097 );
and \U$7389 ( \16207_16509 , RIfca0bc8_6851, \8800_9099 );
and \U$7390 ( \16208_16510 , RIfc48680_5846, \8802_9101 );
and \U$7391 ( \16209_16511 , RIee3dea0_5163, \8804_9103 );
and \U$7392 ( \16210_16512 , RIfcc6878_7281, \8806_9105 );
and \U$7393 ( \16211_16513 , RIee3ba10_5137, \8808_9107 );
and \U$7394 ( \16212_16514 , RIee3a930_5125, \8810_9109 );
and \U$7395 ( \16213_16515 , RIfe97290_8064, \8812_9111 );
and \U$7396 ( \16214_16516 , RIe172b00_2682, \8814_9113 );
and \U$7397 ( \16215_16517 , RIf16f958_5729, \8816_9115 );
and \U$7398 ( \16216_16518 , RIf16ee18_5721, \8818_9117 );
and \U$7399 ( \16217_16519 , RIf16da68_5707, \8820_9119 );
and \U$7400 ( \16218_16520 , RIf16d360_5702, \8822_9121 );
and \U$7401 ( \16219_16521 , RIfe96e58_8061, \8824_9123 );
and \U$7402 ( \16220_16522 , RIe222a50_4684, \8826_9125 );
and \U$7403 ( \16221_16523 , RIfe96cf0_8060, \8828_9127 );
and \U$7404 ( \16222_16524 , RIe21fd50_4652, \8830_9129 );
and \U$7405 ( \16223_16525 , RIf16a660_5670, \8832_9131 );
and \U$7406 ( \16224_16526 , RIe21d050_4620, \8834_9133 );
and \U$7407 ( \16225_16527 , RIe217650_4556, \8836_9135 );
and \U$7408 ( \16226_16528 , RIe214950_4524, \8838_9137 );
and \U$7409 ( \16227_16529 , RIf169f58_5665, \8840_9139 );
and \U$7410 ( \16228_16530 , RIe211c50_4492, \8842_9141 );
and \U$7411 ( \16229_16531 , RIf168770_5648, \8844_9143 );
and \U$7412 ( \16230_16532 , RIe20ef50_4460, \8846_9145 );
and \U$7413 ( \16231_16533 , RIf1677f8_5637, \8848_9147 );
and \U$7414 ( \16232_16534 , RIe20c250_4428, \8850_9149 );
and \U$7415 ( \16233_16535 , RIe209550_4396, \8852_9151 );
and \U$7416 ( \16234_16536 , RIe206850_4364, \8854_9153 );
and \U$7417 ( \16235_16537 , RIf166880_5626, \8856_9155 );
and \U$7418 ( \16236_16538 , RIf1657a0_5614, \8858_9157 );
and \U$7419 ( \16237_16539 , RIe201dc8_4311, \8860_9159 );
and \U$7420 ( \16238_16540 , RIe2005e0_4294, \8862_9161 );
and \U$7421 ( \16239_16541 , RIfe96b88_8059, \8864_9163 );
and \U$7422 ( \16240_16542 , RIf163b80_5594, \8866_9165 );
and \U$7423 ( \16241_16543 , RIf162c08_5583, \8868_9167 );
and \U$7424 ( \16242_16544 , RIf161420_5566, \8870_9169 );
and \U$7425 ( \16243_16545 , RIf15f530_5544, \8872_9171 );
and \U$7426 ( \16244_16546 , RIf15d7a8_5523, \8874_9173 );
and \U$7427 ( \16245_16547 , RIfe968b8_8057, \8876_9175 );
and \U$7428 ( \16246_16548 , RIfe96a20_8058, \8878_9177 );
and \U$7429 ( \16247_16549 , RIfcb3fc0_7070, \8880_9179 );
and \U$7430 ( \16248_16550 , RIfc7cf70_6444, \8882_9181 );
and \U$7431 ( \16249_16551 , RIfc579c8_6019, \8884_9183 );
and \U$7432 ( \16250_16552 , RIf159590_5476, \8886_9185 );
or \U$7433 ( \16251_16553 , \16187_16489 , \16188_16490 , \16189_16491 , \16190_16492 , \16191_16493 , \16192_16494 , \16193_16495 , \16194_16496 , \16195_16497 , \16196_16498 , \16197_16499 , \16198_16500 , \16199_16501 , \16200_16502 , \16201_16503 , \16202_16504 , \16203_16505 , \16204_16506 , \16205_16507 , \16206_16508 , \16207_16509 , \16208_16510 , \16209_16511 , \16210_16512 , \16211_16513 , \16212_16514 , \16213_16515 , \16214_16516 , \16215_16517 , \16216_16518 , \16217_16519 , \16218_16520 , \16219_16521 , \16220_16522 , \16221_16523 , \16222_16524 , \16223_16525 , \16224_16526 , \16225_16527 , \16226_16528 , \16227_16529 , \16228_16530 , \16229_16531 , \16230_16532 , \16231_16533 , \16232_16534 , \16233_16535 , \16234_16536 , \16235_16537 , \16236_16538 , \16237_16539 , \16238_16540 , \16239_16541 , \16240_16542 , \16241_16543 , \16242_16544 , \16243_16545 , \16244_16546 , \16245_16547 , \16246_16548 , \16247_16549 , \16248_16550 , \16249_16551 , \16250_16552 );
and \U$7434 ( \16252_16554 , RIf1584b0_5464, \8889_9188 );
and \U$7435 ( \16253_16555 , RIf157268_5451, \8891_9190 );
and \U$7436 ( \16254_16556 , RIf1569f8_5445, \8893_9192 );
and \U$7437 ( \16255_16557 , RIfe965e8_8055, \8895_9194 );
and \U$7438 ( \16256_16558 , RIf155d50_5436, \8897_9196 );
and \U$7439 ( \16257_16559 , RIf155210_5428, \8899_9198 );
and \U$7440 ( \16258_16560 , RIf153e60_5414, \8901_9200 );
and \U$7441 ( \16259_16561 , RIfe96750_8056, \8903_9202 );
and \U$7442 ( \16260_16562 , RIf1527e0_5398, \8905_9204 );
and \U$7443 ( \16261_16563 , RIf151430_5384, \8907_9206 );
and \U$7444 ( \16262_16564 , RIfcd2650_7416, \8909_9208 );
and \U$7445 ( \16263_16565 , RIe1f2648_4135, \8911_9210 );
and \U$7446 ( \16264_16566 , RIf14f108_5359, \8913_9212 );
and \U$7447 ( \16265_16567 , RIfc7f298_6469, \8915_9214 );
and \U$7448 ( \16266_16568 , RIf14d4e8_5339, \8917_9216 );
and \U$7449 ( \16267_16569 , RIe1ed350_4076, \8919_9218 );
and \U$7450 ( \16268_16570 , RIe1ea7b8_4045, \8921_9220 );
and \U$7451 ( \16269_16571 , RIe1e7ab8_4013, \8923_9222 );
and \U$7452 ( \16270_16572 , RIe1e4db8_3981, \8925_9224 );
and \U$7453 ( \16271_16573 , RIe1e20b8_3949, \8927_9226 );
and \U$7454 ( \16272_16574 , RIe1df3b8_3917, \8929_9228 );
and \U$7455 ( \16273_16575 , RIe1dc6b8_3885, \8931_9230 );
and \U$7456 ( \16274_16576 , RIe1d99b8_3853, \8933_9232 );
and \U$7457 ( \16275_16577 , RIe1d6cb8_3821, \8935_9234 );
and \U$7458 ( \16276_16578 , RIe1d12b8_3757, \8937_9236 );
and \U$7459 ( \16277_16579 , RIe1ce5b8_3725, \8939_9238 );
and \U$7460 ( \16278_16580 , RIe1cb8b8_3693, \8941_9240 );
and \U$7461 ( \16279_16581 , RIe1c8bb8_3661, \8943_9242 );
and \U$7462 ( \16280_16582 , RIe1c5eb8_3629, \8945_9244 );
and \U$7463 ( \16281_16583 , RIe1c31b8_3597, \8947_9246 );
and \U$7464 ( \16282_16584 , RIe1c04b8_3565, \8949_9248 );
and \U$7465 ( \16283_16585 , RIe1bd7b8_3533, \8951_9250 );
and \U$7466 ( \16284_16586 , RIf14c138_5325, \8953_9252 );
and \U$7467 ( \16285_16587 , RIf14ad88_5311, \8955_9254 );
and \U$7468 ( \16286_16588 , RIe1b8790_3476, \8957_9256 );
and \U$7469 ( \16287_16589 , RIfe96480_8054, \8959_9258 );
and \U$7470 ( \16288_16590 , RIf14a0e0_5302, \8961_9260 );
and \U$7471 ( \16289_16591 , RIf149870_5296, \8963_9262 );
and \U$7472 ( \16290_16592 , RIfe97128_8063, \8965_9264 );
and \U$7473 ( \16291_16593 , RIfe96318_8053, \8967_9266 );
and \U$7474 ( \16292_16594 , RIf148628_5283, \8969_9268 );
and \U$7475 ( \16293_16595 , RIfc58d78_6033, \8971_9270 );
and \U$7476 ( \16294_16596 , RIe1b20e8_3403, \8973_9272 );
and \U$7477 ( \16295_16597 , RIe1b04c8_3383, \8975_9274 );
and \U$7478 ( \16296_16598 , RIf146cd8_5265, \8977_9276 );
and \U$7479 ( \16297_16599 , RIfc591b0_6036, \8979_9278 );
and \U$7480 ( \16298_16600 , RIfe961b0_8052, \8981_9280 );
and \U$7481 ( \16299_16601 , RIfe96fc0_8062, \8983_9282 );
and \U$7482 ( \16300_16602 , RIe1a7af8_3285, \8985_9284 );
and \U$7483 ( \16301_16603 , RIe1a4df8_3253, \8987_9286 );
and \U$7484 ( \16302_16604 , RIe1a20f8_3221, \8989_9288 );
and \U$7485 ( \16303_16605 , RIe19f3f8_3189, \8991_9290 );
and \U$7486 ( \16304_16606 , RIe18b8f8_2965, \8993_9292 );
and \U$7487 ( \16305_16607 , RIe177df8_2741, \8995_9294 );
and \U$7488 ( \16306_16608 , RIe225750_4716, \8997_9296 );
and \U$7489 ( \16307_16609 , RIe21a350_4588, \8999_9298 );
and \U$7490 ( \16308_16610 , RIe203b50_4332, \9001_9300 );
and \U$7491 ( \16309_16611 , RIe1fdbb0_4264, \9003_9302 );
and \U$7492 ( \16310_16612 , RIe1f6f68_4187, \9005_9304 );
and \U$7493 ( \16311_16613 , RIe1efab0_4104, \9007_9306 );
and \U$7494 ( \16312_16614 , RIe1d3fb8_3789, \9009_9308 );
and \U$7495 ( \16313_16615 , RIe1baab8_3501, \9011_9310 );
and \U$7496 ( \16314_16616 , RIe1ad930_3352, \9013_9312 );
and \U$7497 ( \16315_16617 , RIe16ff68_2651, \9015_9314 );
or \U$7498 ( \16316_16618 , \16252_16554 , \16253_16555 , \16254_16556 , \16255_16557 , \16256_16558 , \16257_16559 , \16258_16560 , \16259_16561 , \16260_16562 , \16261_16563 , \16262_16564 , \16263_16565 , \16264_16566 , \16265_16567 , \16266_16568 , \16267_16569 , \16268_16570 , \16269_16571 , \16270_16572 , \16271_16573 , \16272_16574 , \16273_16575 , \16274_16576 , \16275_16577 , \16276_16578 , \16277_16579 , \16278_16580 , \16279_16581 , \16280_16582 , \16281_16583 , \16282_16584 , \16283_16585 , \16284_16586 , \16285_16587 , \16286_16588 , \16287_16589 , \16288_16590 , \16289_16591 , \16290_16592 , \16291_16593 , \16292_16594 , \16293_16595 , \16294_16596 , \16295_16597 , \16296_16598 , \16297_16599 , \16298_16600 , \16299_16601 , \16300_16602 , \16301_16603 , \16302_16604 , \16303_16605 , \16304_16606 , \16305_16607 , \16306_16608 , \16307_16609 , \16308_16610 , \16309_16611 , \16310_16612 , \16311_16613 , \16312_16614 , \16313_16615 , \16314_16616 , \16315_16617 );
or \U$7499 ( \16317_16619 , \16251_16553 , \16316_16618 );
_DC \g50c1/U$1 ( \16318 , \16317_16619 , \9024_9323 );
xor g50c2_GF_PartitionCandidate( \16319_16621_nG50c2 , \16186 , \16318 );
buf \U$7500 ( \16320_16622 , \16319_16621_nG50c2 );
and \U$7501 ( \16321_16623 , \15998_16300 , \15034_15333 );
not \U$7502 ( \16322_16624 , \16321_16623 );
and \U$7503 ( \16323_16625 , \16320_16622 , \16322_16624 );
and \U$7504 ( \16324_16626 , \16054_16356 , \16323_16625 );
xor \U$7505 ( \16325_16627 , \16053_16355 , \16324_16626 );
and \U$7506 ( \16326_16628 , \13377_13679 , \12491_12790 );
and \U$7507 ( \16327_16629 , \13725_14024 , \12159_12461 );
nor \U$7508 ( \16328_16630 , \16326_16628 , \16327_16629 );
xnor \U$7509 ( \16329_16631 , \16328_16630 , \12481_12780 );
xor \U$7510 ( \16330_16632 , \16325_16627 , \16329_16631 );
xor \U$7511 ( \16331_16633 , \16320_16622 , \15998_16300 );
not \U$7512 ( \16332_16634 , \15999_16301 );
and \U$7513 ( \16333_16635 , \16331_16633 , \16332_16634 );
and \U$7514 ( \16334_16636 , \10385_10687 , \16333_16635 );
and \U$7515 ( \16335_16637 , \10686_10988 , \15999_16301 );
nor \U$7516 ( \16336_16638 , \16334_16636 , \16335_16637 );
xnor \U$7517 ( \16337_16639 , \16336_16638 , \16323_16625 );
xor \U$7518 ( \16338_16640 , \16330_16632 , \16337_16639 );
xor \U$7519 ( \16339_16641 , \16049_16351 , \16338_16640 );
and \U$7520 ( \16340_16642 , \15989_16291 , \15993_16295 );
and \U$7521 ( \16341_16643 , \15993_16295 , \16000_16302 );
and \U$7522 ( \16342_16644 , \15989_16291 , \16000_16302 );
or \U$7523 ( \16343_16645 , \16340_16642 , \16341_16643 , \16342_16644 );
and \U$7524 ( \16344_16646 , \15968_16270 , \15972_16274 );
and \U$7525 ( \16345_16647 , \15972_16274 , \15977_16279 );
and \U$7526 ( \16346_16648 , \15968_16270 , \15977_16279 );
or \U$7527 ( \16347_16649 , \16344_16646 , \16345_16647 , \16346_16648 );
xor \U$7528 ( \16348_16650 , \16343_16645 , \16347_16649 );
and \U$7529 ( \16349_16651 , \15965_16267 , \10681_10983 );
_DC \g6598/U$1 ( \16350 , \16185_16487 , \9298_9597 );
_DC \g6599/U$1 ( \16351 , \16317_16619 , \9024_9323 );
and g659a_GF_PartitionCandidate( \16352_16654_nG659a , \16350 , \16351 );
buf \U$7530 ( \16353_16655 , \16352_16654_nG659a );
and \U$7531 ( \16354_16656 , \16353_16655 , \10389_10691 );
nor \U$7532 ( \16355_16657 , \16349_16651 , \16354_16656 );
xnor \U$7533 ( \16356_16658 , \16355_16657 , \10678_10980 );
and \U$7534 ( \16357_16659 , \12146_12448 , \13755_14054 );
and \U$7535 ( \16358_16660 , \12470_12769 , \13390_13692 );
nor \U$7536 ( \16359_16661 , \16357_16659 , \16358_16660 );
xnor \U$7537 ( \16360_16662 , \16359_16661 , \13736_14035 );
xor \U$7538 ( \16361_16663 , \16356_16658 , \16360_16662 );
and \U$7539 ( \16362_16664 , \10968_11270 , \15037_15336 );
and \U$7540 ( \16363_16665 , \11287_11586 , \14661_14963 );
nor \U$7541 ( \16364_16666 , \16362_16664 , \16363_16665 );
xnor \U$7542 ( \16365_16667 , \16364_16666 , \15043_15342 );
xor \U$7543 ( \16366_16668 , \16361_16663 , \16365_16667 );
xor \U$7544 ( \16367_16669 , \16348_16650 , \16366_16668 );
xor \U$7545 ( \16368_16670 , \16339_16641 , \16367_16669 );
and \U$7546 ( \16369_16671 , \15698_16000 , \15978_16280 );
and \U$7547 ( \16370_16672 , \15978_16280 , \16002_16304 );
and \U$7548 ( \16371_16673 , \15698_16000 , \16002_16304 );
or \U$7549 ( \16372_16674 , \16369_16671 , \16370_16672 , \16371_16673 );
xor \U$7550 ( \16373_16675 , \16368_16670 , \16372_16674 );
and \U$7551 ( \16374_16676 , \16003_16305 , \16007_16309 );
and \U$7552 ( \16375_16677 , \16008_16310 , \16011_16313 );
or \U$7553 ( \16376_16678 , \16374_16676 , \16375_16677 );
xor \U$7554 ( \16377_16679 , \16373_16675 , \16376_16678 );
buf g9bed_GF_PartitionCandidate( \16378_16680_nG9bed , \16377_16679 );
and \U$7555 ( \16379_16681 , \10402_10704 , \16378_16680_nG9bed );
or \U$7556 ( \16380_16682 , \16045_16347 , \16379_16681 );
xor \U$7557 ( \16381_16683 , \10399_10703 , \16380_16682 );
buf \U$7558 ( \16382_16684 , \16381_16683 );
buf \U$7560 ( \16383_16685 , \16382_16684 );
xor \U$7561 ( \16384_16686 , \16044_16346 , \16383_16685 );
buf \U$7562 ( \16385_16687 , \16384_16686 );
and \U$7563 ( \16386_16688 , \15686_15988 , \15692_15994 );
and \U$7564 ( \16387_16689 , \15686_15988 , \16018_16320 );
and \U$7565 ( \16388_16690 , \15692_15994 , \16018_16320 );
or \U$7566 ( \16389_16691 , \16386_16688 , \16387_16689 , \16388_16690 );
buf \U$7567 ( \16390_16692 , \16389_16691 );
xor \U$7568 ( \16391_16693 , \16385_16687 , \16390_16692 );
and \U$7569 ( \16392_16694 , \15637_15936 , \15641_15943 );
buf \U$7570 ( \16393_16695 , \16392_16694 );
buf \U$7572 ( \16394_16696 , \16393_16695 );
and \U$7573 ( \16395_16697 , \14710_14631 , \10981_11283_nG9c08 );
and \U$7574 ( \16396_16698 , \14329_14628 , \11299_11598_nG9c05 );
or \U$7575 ( \16397_16699 , \16395_16697 , \16396_16698 );
xor \U$7576 ( \16398_16700 , \14328_14627 , \16397_16699 );
buf \U$7577 ( \16399_16701 , \16398_16700 );
buf \U$7579 ( \16400_16702 , \16399_16701 );
xor \U$7580 ( \16401_16703 , \16394_16696 , \16400_16702 );
buf \U$7581 ( \16402_16704 , \16401_16703 );
not \U$6819 ( \16403_15938 , \15638_15937 );
xor \U$6820 ( \16404_15939 , \15632_15931_nG4436 , \15635_15934_nG4439 );
and \U$6821 ( \16405_15940 , \16403_15938 , \16404_15939 );
and \U$7582 ( \16406_16705 , \16405_15940 , \10392_10694_nG9c0e );
and \U$7583 ( \16407_16706 , \15638_15937 , \10693_10995_nG9c0b );
or \U$7584 ( \16408_16707 , \16406_16705 , \16407_16706 );
xor \U$7585 ( \16409_16708 , \15637_15936 , \16408_16707 );
buf \U$7586 ( \16410_16709 , \16409_16708 );
buf \U$7588 ( \16411_16710 , \16410_16709 );
xor \U$7589 ( \16412_16711 , \16402_16704 , \16411_16710 );
and \U$7590 ( \16413_16712 , \13431_13370 , \12168_12470_nG9c02 );
and \U$7591 ( \16414_16713 , \13068_13367 , \12502_12801_nG9bff );
or \U$7592 ( \16415_16714 , \16413_16712 , \16414_16713 );
xor \U$7593 ( \16416_16715 , \13067_13366 , \16415_16714 );
buf \U$7594 ( \16417_16716 , \16416_16715 );
buf \U$7596 ( \16418_16717 , \16417_16716 );
xor \U$7597 ( \16419_16718 , \16412_16711 , \16418_16717 );
buf \U$7598 ( \16420_16719 , \16419_16718 );
and \U$7599 ( \16421_16720 , \15661_15963 , \15667_15969 );
buf \U$7600 ( \16422_16721 , \16421_16720 );
xor \U$7601 ( \16423_16722 , \16420_16719 , \16422_16721 );
and \U$7602 ( \16424_16723 , \12183_12157 , \13403_13705_nG9bfc );
and \U$7603 ( \16425_16724 , \11855_12154 , \13771_14070_nG9bf9 );
or \U$7604 ( \16426_16725 , \16424_16723 , \16425_16724 );
xor \U$7605 ( \16427_16726 , \11854_12153 , \16426_16725 );
buf \U$7606 ( \16428_16727 , \16427_16726 );
buf \U$7608 ( \16429_16728 , \16428_16727 );
xor \U$7609 ( \16430_16729 , \16423_16722 , \16429_16728 );
buf \U$7610 ( \16431_16730 , \16430_16729 );
xor \U$7611 ( \16432_16731 , \16391_16693 , \16431_16730 );
buf \U$7612 ( \16433_16732 , \16432_16731 );
and \U$7613 ( \16434_16733 , \15655_15957 , \15680_15982 );
and \U$7614 ( \16435_16734 , \15655_15957 , \16020_16322 );
and \U$7615 ( \16436_16735 , \15680_15982 , \16020_16322 );
or \U$7616 ( \16437_16736 , \16434_16733 , \16435_16734 , \16436_16735 );
buf \U$7617 ( \16438_16737 , \16437_16736 );
xor \U$7618 ( \16439_16738 , \16433_16732 , \16438_16737 );
and \U$7619 ( \16440_16739 , \15650_15952 , \16022_16324 );
and \U$7620 ( \16441_16740 , \15650_15952 , \16028_16330 );
and \U$7621 ( \16442_16741 , \16022_16324 , \16028_16330 );
or \U$7622 ( \16443_16742 , \16440_16739 , \16441_16740 , \16442_16741 );
buf \U$7623 ( \16444_16743 , \16443_16742 );
xor \U$7624 ( \16445_16744 , \16439_16738 , \16444_16743 );
and \U$7625 ( \16446_16745 , \16032_16334 , \16445_16744 );
and \U$7626 ( \16447_16746 , RIdec4730_699, \8760_9059 );
and \U$7627 ( \16448_16747 , RIdec1a30_667, \8762_9061 );
and \U$7628 ( \16449_16748 , RIfce3f90_7616, \8764_9063 );
and \U$7629 ( \16450_16749 , RIdebed30_635, \8766_9065 );
and \U$7630 ( \16451_16750 , RIfcc3308_7243, \8768_9067 );
and \U$7631 ( \16452_16751 , RIdebc030_603, \8770_9069 );
and \U$7632 ( \16453_16752 , RIdeb9330_571, \8772_9071 );
and \U$7633 ( \16454_16753 , RIdeb6630_539, \8774_9073 );
and \U$7634 ( \16455_16754 , RIfc8c588_6619, \8776_9075 );
and \U$7635 ( \16456_16755 , RIdeb0c30_475, \8778_9077 );
and \U$7636 ( \16457_16756 , RIfc5a998_6053, \8780_9079 );
and \U$7637 ( \16458_16757 , RIdeadf30_443, \8782_9081 );
and \U$7638 ( \16459_16758 , RIfc99b48_6771, \8784_9083 );
and \U$7639 ( \16460_16759 , RIdea8698_411, \8786_9085 );
and \U$7640 ( \16461_16760 , RIdea1d98_379, \8788_9087 );
and \U$7641 ( \16462_16761 , RIde9b498_347, \8790_9089 );
and \U$7642 ( \16463_16762 , RIfc78bf0_6396, \8792_9091 );
and \U$7643 ( \16464_16763 , RIfcbc558_7165, \8794_9093 );
and \U$7644 ( \16465_16764 , RIfca12d0_6856, \8796_9095 );
and \U$7645 ( \16466_16765 , RIfca3fd0_6888, \8798_9097 );
and \U$7646 ( \16467_16766 , RIfec2670_8332, \8800_9099 );
and \U$7647 ( \16468_16767 , RIfec2508_8331, \8802_9101 );
and \U$7648 ( \16469_16768 , RIde88a00_256, \8804_9103 );
and \U$7649 ( \16470_16769 , RIde84518_235, \8806_9105 );
and \U$7650 ( \16471_16770 , RIfcc35d8_7245, \8808_9107 );
and \U$7651 ( \16472_16771 , RIfcb57a8_7087, \8810_9109 );
and \U$7652 ( \16473_16772 , RIfc5a290_6048, \8812_9111 );
and \U$7653 ( \16474_16773 , RIfca3058_6877, \8814_9113 );
and \U$7654 ( \16475_16774 , RIee38e78_5106, \8816_9115 );
and \U$7655 ( \16476_16775 , RIfec27d8_8333, \8818_9117 );
and \U$7656 ( \16477_16776 , RIfca3328_6879, \8820_9119 );
and \U$7657 ( \16478_16777 , RIe1672c8_2551, \8822_9121 );
and \U$7658 ( \16479_16778 , RIe164730_2520, \8824_9123 );
and \U$7659 ( \16480_16779 , RIe161a30_2488, \8826_9125 );
and \U$7660 ( \16481_16780 , RIee36cb8_5082, \8828_9127 );
and \U$7661 ( \16482_16781 , RIe15ed30_2456, \8830_9129 );
and \U$7662 ( \16483_16782 , RIfcc7250_7288, \8832_9131 );
and \U$7663 ( \16484_16783 , RIe15c030_2424, \8834_9133 );
and \U$7664 ( \16485_16784 , RIe156630_2360, \8836_9135 );
and \U$7665 ( \16486_16785 , RIe153930_2328, \8838_9137 );
and \U$7666 ( \16487_16786 , RIfcc7688_7291, \8840_9139 );
and \U$7667 ( \16488_16787 , RIe150c30_2296, \8842_9141 );
and \U$7668 ( \16489_16788 , RIfc8af08_6603, \8844_9143 );
and \U$7669 ( \16490_16789 , RIe14df30_2264, \8846_9145 );
and \U$7670 ( \16491_16790 , RIfc9a250_6776, \8848_9147 );
and \U$7671 ( \16492_16791 , RIe14b230_2232, \8850_9149 );
and \U$7672 ( \16493_16792 , RIe148530_2200, \8852_9151 );
and \U$7673 ( \16494_16793 , RIe145830_2168, \8854_9153 );
and \U$7674 ( \16495_16794 , RIfc9aac0_6782, \8856_9155 );
and \U$7675 ( \16496_16795 , RIfc56bb8_6009, \8858_9157 );
and \U$7676 ( \16497_16796 , RIfca1ca8_6863, \8860_9159 );
and \U$7677 ( \16498_16797 , RIfcec960_7714, \8862_9161 );
and \U$7678 ( \16499_16798 , RIe1406a0_2110, \8864_9163 );
and \U$7679 ( \16500_16799 , RIdf3e440_2085, \8866_9165 );
and \U$7680 ( \16501_16800 , RIdf3c280_2061, \8868_9167 );
and \U$7681 ( \16502_16801 , RIdf39f58_2036, \8870_9169 );
and \U$7682 ( \16503_16802 , RIfc9a958_6781, \8872_9171 );
and \U$7683 ( \16504_16803 , RIee2f0f8_4994, \8874_9173 );
and \U$7684 ( \16505_16804 , RIfcdb458_7517, \8876_9175 );
and \U$7685 ( \16506_16805 , RIee2cf38_4970, \8878_9177 );
and \U$7686 ( \16507_16806 , RIdf34c60_1977, \8880_9179 );
and \U$7687 ( \16508_16807 , RIfec2940_8334, \8882_9181 );
and \U$7688 ( \16509_16808 , RIdf30778_1928, \8884_9183 );
and \U$7689 ( \16510_16809 , RIdf2e888_1906, \8886_9185 );
or \U$7690 ( \16511_16810 , \16447_16746 , \16448_16747 , \16449_16748 , \16450_16749 , \16451_16750 , \16452_16751 , \16453_16752 , \16454_16753 , \16455_16754 , \16456_16755 , \16457_16756 , \16458_16757 , \16459_16758 , \16460_16759 , \16461_16760 , \16462_16761 , \16463_16762 , \16464_16763 , \16465_16764 , \16466_16765 , \16467_16766 , \16468_16767 , \16469_16768 , \16470_16769 , \16471_16770 , \16472_16771 , \16473_16772 , \16474_16773 , \16475_16774 , \16476_16775 , \16477_16776 , \16478_16777 , \16479_16778 , \16480_16779 , \16481_16780 , \16482_16781 , \16483_16782 , \16484_16783 , \16485_16784 , \16486_16785 , \16487_16786 , \16488_16787 , \16489_16788 , \16490_16789 , \16491_16790 , \16492_16791 , \16493_16792 , \16494_16793 , \16495_16794 , \16496_16795 , \16497_16796 , \16498_16797 , \16499_16798 , \16500_16799 , \16501_16800 , \16502_16801 , \16503_16802 , \16504_16803 , \16505_16804 , \16506_16805 , \16507_16806 , \16508_16807 , \16509_16808 , \16510_16809 );
and \U$7691 ( \16512_16811 , RIee2b480_4951, \8889_9188 );
and \U$7692 ( \16513_16812 , RIfec23a0_8330, \8891_9190 );
and \U$7693 ( \16514_16813 , RIee288e8_4920, \8893_9192 );
and \U$7694 ( \16515_16814 , RIfec2238_8329, \8895_9194 );
and \U$7695 ( \16516_16815 , RIdf29b30_1851, \8897_9196 );
and \U$7696 ( \16517_16816 , RIdf27808_1826, \8899_9198 );
and \U$7697 ( \16518_16817 , RIdf25a80_1805, \8901_9200 );
and \U$7698 ( \16519_16818 , RIdf23e60_1785, \8903_9202 );
and \U$7699 ( \16520_16819 , RIfc55100_5990, \8905_9204 );
and \U$7700 ( \16521_16820 , RIfcd9f40_7502, \8907_9206 );
and \U$7701 ( \16522_16821 , RIfc54f98_5989, \8909_9208 );
and \U$7702 ( \16523_16822 , RIfc54cc8_5987, \8911_9210 );
and \U$7703 ( \16524_16823 , RIfc4b218_5877, \8913_9212 );
and \U$7704 ( \16525_16824 , RIdf1efa0_1729, \8915_9214 );
and \U$7705 ( \16526_16825 , RIfcc69e0_7282, \8917_9216 );
and \U$7706 ( \16527_16826 , RIdf18bc8_1658, \8919_9218 );
and \U$7707 ( \16528_16827 , RIdf16300_1629, \8921_9220 );
and \U$7708 ( \16529_16828 , RIdf13600_1597, \8923_9222 );
and \U$7709 ( \16530_16829 , RIdf10900_1565, \8925_9224 );
and \U$7710 ( \16531_16830 , RIdf0dc00_1533, \8927_9226 );
and \U$7711 ( \16532_16831 , RIdf0af00_1501, \8929_9228 );
and \U$7712 ( \16533_16832 , RIdf08200_1469, \8931_9230 );
and \U$7713 ( \16534_16833 , RIdf05500_1437, \8933_9232 );
and \U$7714 ( \16535_16834 , RIdf02800_1405, \8935_9234 );
and \U$7715 ( \16536_16835 , RIdefce00_1341, \8937_9236 );
and \U$7716 ( \16537_16836 , RIdefa100_1309, \8939_9238 );
and \U$7717 ( \16538_16837 , RIdef7400_1277, \8941_9240 );
and \U$7718 ( \16539_16838 , RIdef4700_1245, \8943_9242 );
and \U$7719 ( \16540_16839 , RIdef1a00_1213, \8945_9244 );
and \U$7720 ( \16541_16840 , RIdeeed00_1181, \8947_9246 );
and \U$7721 ( \16542_16841 , RIdeec000_1149, \8949_9248 );
and \U$7722 ( \16543_16842 , RIdee9300_1117, \8951_9250 );
and \U$7723 ( \16544_16843 , RIfce4ad0_7624, \8953_9252 );
and \U$7724 ( \16545_16844 , RIfc9e8a0_6826, \8955_9254 );
and \U$7725 ( \16546_16845 , RIfcc46b8_7257, \8957_9256 );
and \U$7726 ( \16547_16846 , RIfcd4108_7435, \8959_9258 );
and \U$7727 ( \16548_16847 , RIdee4440_1061, \8961_9260 );
and \U$7728 ( \16549_16848 , RIdee2280_1037, \8963_9262 );
and \U$7729 ( \16550_16849 , RIdee0390_1015, \8965_9264 );
and \U$7730 ( \16551_16850 , RIdede068_990, \8967_9266 );
and \U$7731 ( \16552_16851 , RIfcda0a8_7503, \8969_9268 );
and \U$7732 ( \16553_16852 , RIfce54a8_7631, \8971_9270 );
and \U$7733 ( \16554_16853 , RIfca0790_6848, \8973_9272 );
and \U$7734 ( \16555_16854 , RIfc50ee8_5943, \8975_9274 );
and \U$7735 ( \16556_16855 , RIded8d70_931, \8977_9276 );
and \U$7736 ( \16557_16856 , RIded68e0_905, \8979_9278 );
and \U$7737 ( \16558_16857 , RIded4888_882, \8981_9280 );
and \U$7738 ( \16559_16858 , RIded2560_857, \8983_9282 );
and \U$7739 ( \16560_16859 , RIdecfb30_827, \8985_9284 );
and \U$7740 ( \16561_16860 , RIdecce30_795, \8987_9286 );
and \U$7741 ( \16562_16861 , RIdeca130_763, \8989_9288 );
and \U$7742 ( \16563_16862 , RIdec7430_731, \8991_9290 );
and \U$7743 ( \16564_16863 , RIdeb3930_507, \8993_9292 );
and \U$7744 ( \16565_16864 , RIde94b98_315, \8995_9294 );
and \U$7745 ( \16566_16865 , RIe16d538_2621, \8997_9296 );
and \U$7746 ( \16567_16866 , RIe159330_2392, \8999_9298 );
and \U$7747 ( \16568_16867 , RIe142b30_2136, \9001_9300 );
and \U$7748 ( \16569_16868 , RIdf37528_2006, \9003_9302 );
and \U$7749 ( \16570_16869 , RIdf2bb88_1874, \9005_9304 );
and \U$7750 ( \16571_16870 , RIdf1c408_1698, \9007_9306 );
and \U$7751 ( \16572_16871 , RIdeffb00_1373, \9009_9308 );
and \U$7752 ( \16573_16872 , RIdee6600_1085, \9011_9310 );
and \U$7753 ( \16574_16873 , RIdedb368_958, \9013_9312 );
and \U$7754 ( \16575_16874 , RIde7aae0_188, \9015_9314 );
or \U$7755 ( \16576_16875 , \16512_16811 , \16513_16812 , \16514_16813 , \16515_16814 , \16516_16815 , \16517_16816 , \16518_16817 , \16519_16818 , \16520_16819 , \16521_16820 , \16522_16821 , \16523_16822 , \16524_16823 , \16525_16824 , \16526_16825 , \16527_16826 , \16528_16827 , \16529_16828 , \16530_16829 , \16531_16830 , \16532_16831 , \16533_16832 , \16534_16833 , \16535_16834 , \16536_16835 , \16537_16836 , \16538_16837 , \16539_16838 , \16540_16839 , \16541_16840 , \16542_16841 , \16543_16842 , \16544_16843 , \16545_16844 , \16546_16845 , \16547_16846 , \16548_16847 , \16549_16848 , \16550_16849 , \16551_16850 , \16552_16851 , \16553_16852 , \16554_16853 , \16555_16854 , \16556_16855 , \16557_16856 , \16558_16857 , \16559_16858 , \16560_16859 , \16561_16860 , \16562_16861 , \16563_16862 , \16564_16863 , \16565_16864 , \16566_16865 , \16567_16866 , \16568_16867 , \16569_16868 , \16570_16869 , \16571_16870 , \16572_16871 , \16573_16872 , \16574_16873 , \16575_16874 );
or \U$7756 ( \16577_16876 , \16511_16810 , \16576_16875 );
_DC \g2b8f/U$1 ( \16578 , \16577_16876 , \9024_9323 );
buf \U$7757 ( \16579_16878 , \16578 );
and \U$7758 ( \16580_16879 , RIe19c9c8_3159, \9034_9333 );
and \U$7759 ( \16581_16880 , RIe199cc8_3127, \9036_9335 );
and \U$7760 ( \16582_16881 , RIfe8ea28_7967, \9038_9337 );
and \U$7761 ( \16583_16882 , RIe196fc8_3095, \9040_9339 );
and \U$7762 ( \16584_16883 , RIfec20d0_8328, \9042_9341 );
and \U$7763 ( \16585_16884 , RIe1942c8_3063, \9044_9343 );
and \U$7764 ( \16586_16885 , RIe1915c8_3031, \9046_9345 );
and \U$7765 ( \16587_16886 , RIe18e8c8_2999, \9048_9347 );
and \U$7766 ( \16588_16887 , RIe188ec8_2935, \9050_9349 );
and \U$7767 ( \16589_16888 , RIe1861c8_2903, \9052_9351 );
and \U$7768 ( \16590_16889 , RIfc68228_6207, \9054_9353 );
and \U$7769 ( \16591_16890 , RIe1834c8_2871, \9056_9355 );
and \U$7770 ( \16592_16891 , RIfccb5d0_7336, \9058_9357 );
and \U$7771 ( \16593_16892 , RIe1807c8_2839, \9060_9359 );
and \U$7772 ( \16594_16893 , RIe17dac8_2807, \9062_9361 );
and \U$7773 ( \16595_16894 , RIe17adc8_2775, \9064_9363 );
and \U$7774 ( \16596_16895 , RIf141e18_5209, \9066_9365 );
and \U$7775 ( \16597_16896 , RIf140900_5194, \9068_9367 );
and \U$7776 ( \16598_16897 , RIf140090_5188, \9070_9369 );
and \U$7777 ( \16599_16898 , RIe1753c8_2711, \9072_9371 );
and \U$7778 ( \16600_16899 , RIf13f988_5183, \9074_9373 );
and \U$7779 ( \16601_16900 , RIf13ece0_5174, \9076_9375 );
and \U$7780 ( \16602_16901 , RIee3e170_5165, \9078_9377 );
and \U$7781 ( \16603_16902 , RIee3cf28_5152, \9080_9379 );
and \U$7782 ( \16604_16903 , RIee3bce0_5139, \9082_9381 );
and \U$7783 ( \16605_16904 , RIee3ac00_5127, \9084_9383 );
and \U$7784 ( \16606_16905 , RIee39850_5113, \9086_9385 );
and \U$7785 ( \16607_16906 , RIe172dd0_2684, \9088_9387 );
and \U$7786 ( \16608_16907 , RIf16fc28_5731, \9090_9389 );
and \U$7787 ( \16609_16908 , RIf16f0e8_5723, \9092_9391 );
and \U$7788 ( \16610_16909 , RIf16dd38_5709, \9094_9393 );
and \U$7789 ( \16611_16910 , RIfce9120_7674, \9096_9395 );
and \U$7790 ( \16612_16911 , RIfc404a8_5757, \9098_9397 );
and \U$7791 ( \16613_16912 , RIe222d20_4686, \9100_9399 );
and \U$7792 ( \16614_16913 , RIf16b8a8_5683, \9102_9401 );
and \U$7793 ( \16615_16914 , RIe220020_4654, \9104_9403 );
and \U$7794 ( \16616_16915 , RIf16a930_5672, \9106_9405 );
and \U$7795 ( \16617_16916 , RIe21d320_4622, \9108_9407 );
and \U$7796 ( \16618_16917 , RIe217920_4558, \9110_9409 );
and \U$7797 ( \16619_16918 , RIe214c20_4526, \9112_9411 );
and \U$7798 ( \16620_16919 , RIfc5b910_6064, \9114_9413 );
and \U$7799 ( \16621_16920 , RIe211f20_4494, \9116_9415 );
and \U$7800 ( \16622_16921 , RIfe8e8c0_7966, \9118_9417 );
and \U$7801 ( \16623_16922 , RIe20f220_4462, \9120_9419 );
and \U$7802 ( \16624_16923 , RIfe8e758_7965, \9122_9421 );
and \U$7803 ( \16625_16924 , RIe20c520_4430, \9124_9423 );
and \U$7804 ( \16626_16925 , RIe209820_4398, \9126_9425 );
and \U$7805 ( \16627_16926 , RIe206b20_4366, \9128_9427 );
and \U$7806 ( \16628_16927 , RIf166b50_5628, \9130_9429 );
and \U$7807 ( \16629_16928 , RIf165a70_5616, \9132_9431 );
and \U$7808 ( \16630_16929 , RIfe8dd80_7958, \9134_9433 );
and \U$7809 ( \16631_16930 , RIfe8dab0_7956, \9136_9435 );
and \U$7810 ( \16632_16931 , RIf164c60_5606, \9138_9437 );
and \U$7811 ( \16633_16932 , RIf163e50_5596, \9140_9439 );
and \U$7812 ( \16634_16933 , RIf162ed8_5585, \9142_9441 );
and \U$7813 ( \16635_16934 , RIf1616f0_5568, \9144_9443 );
and \U$7814 ( \16636_16935 , RIf15f800_5546, \9146_9445 );
and \U$7815 ( \16637_16936 , RIf15da78_5525, \9148_9447 );
and \U$7816 ( \16638_16937 , RIfe8d948_7955, \9150_9449 );
and \U$7817 ( \16639_16938 , RIfe8dc18_7957, \9152_9451 );
and \U$7818 ( \16640_16939 , RIf15c560_5510, \9154_9453 );
and \U$7819 ( \16641_16940 , RIf15b048_5495, \9156_9455 );
and \U$7820 ( \16642_16941 , RIfc62828_6143, \9158_9457 );
and \U$7821 ( \16643_16942 , RIf159860_5478, \9160_9459 );
or \U$7822 ( \16644_16943 , \16580_16879 , \16581_16880 , \16582_16881 , \16583_16882 , \16584_16883 , \16585_16884 , \16586_16885 , \16587_16886 , \16588_16887 , \16589_16888 , \16590_16889 , \16591_16890 , \16592_16891 , \16593_16892 , \16594_16893 , \16595_16894 , \16596_16895 , \16597_16896 , \16598_16897 , \16599_16898 , \16600_16899 , \16601_16900 , \16602_16901 , \16603_16902 , \16604_16903 , \16605_16904 , \16606_16905 , \16607_16906 , \16608_16907 , \16609_16908 , \16610_16909 , \16611_16910 , \16612_16911 , \16613_16912 , \16614_16913 , \16615_16914 , \16616_16915 , \16617_16916 , \16618_16917 , \16619_16918 , \16620_16919 , \16621_16920 , \16622_16921 , \16623_16922 , \16624_16923 , \16625_16924 , \16626_16925 , \16627_16926 , \16628_16927 , \16629_16928 , \16630_16929 , \16631_16930 , \16632_16931 , \16633_16932 , \16634_16933 , \16635_16934 , \16636_16935 , \16637_16936 , \16638_16937 , \16639_16938 , \16640_16939 , \16641_16940 , \16642_16941 , \16643_16942 );
and \U$7823 ( \16645_16944 , RIf158780_5466, \9163_9462 );
and \U$7824 ( \16646_16945 , RIf157538_5453, \9165_9464 );
and \U$7825 ( \16647_16946 , RIfca6e38_6921, \9167_9466 );
and \U$7826 ( \16648_16947 , RIe1f9b00_4218, \9169_9468 );
and \U$7827 ( \16649_16948 , RIfc61e50_6136, \9171_9470 );
and \U$7828 ( \16650_16949 , RIfc61748_6131, \9173_9472 );
and \U$7829 ( \16651_16950 , RIf154130_5416, \9175_9474 );
and \U$7830 ( \16652_16951 , RIe1f4ad8_4161, \9177_9476 );
and \U$7831 ( \16653_16952 , RIf152ab0_5400, \9179_9478 );
and \U$7832 ( \16654_16953 , RIf151700_5386, \9181_9480 );
and \U$7833 ( \16655_16954 , RIf1501e8_5371, \9183_9482 );
and \U$7834 ( \16656_16955 , RIe1f27b0_4136, \9185_9484 );
and \U$7835 ( \16657_16956 , RIfc60ed8_6125, \9187_9486 );
and \U$7836 ( \16658_16957 , RIfc7b620_6426, \9189_9488 );
and \U$7837 ( \16659_16958 , RIf14d7b8_5341, \9191_9490 );
and \U$7838 ( \16660_16959 , RIe1ed4b8_4077, \9193_9492 );
and \U$7839 ( \16661_16960 , RIe1eaa88_4047, \9195_9494 );
and \U$7840 ( \16662_16961 , RIe1e7d88_4015, \9197_9496 );
and \U$7841 ( \16663_16962 , RIe1e5088_3983, \9199_9498 );
and \U$7842 ( \16664_16963 , RIe1e2388_3951, \9201_9500 );
and \U$7843 ( \16665_16964 , RIe1df688_3919, \9203_9502 );
and \U$7844 ( \16666_16965 , RIe1dc988_3887, \9205_9504 );
and \U$7845 ( \16667_16966 , RIe1d9c88_3855, \9207_9506 );
and \U$7846 ( \16668_16967 , RIe1d6f88_3823, \9209_9508 );
and \U$7847 ( \16669_16968 , RIe1d1588_3759, \9211_9510 );
and \U$7848 ( \16670_16969 , RIe1ce888_3727, \9213_9512 );
and \U$7849 ( \16671_16970 , RIe1cbb88_3695, \9215_9514 );
and \U$7850 ( \16672_16971 , RIe1c8e88_3663, \9217_9516 );
and \U$7851 ( \16673_16972 , RIe1c6188_3631, \9219_9518 );
and \U$7852 ( \16674_16973 , RIe1c3488_3599, \9221_9520 );
and \U$7853 ( \16675_16974 , RIe1c0788_3567, \9223_9522 );
and \U$7854 ( \16676_16975 , RIe1bda88_3535, \9225_9524 );
and \U$7855 ( \16677_16976 , RIfca4de0_6898, \9227_9526 );
and \U$7856 ( \16678_16977 , RIfc5ea48_6099, \9229_9528 );
and \U$7857 ( \16679_16978 , RIe1b8a60_3478, \9231_9530 );
and \U$7858 ( \16680_16979 , RIe1b6a08_3455, \9233_9532 );
and \U$7859 ( \16681_16980 , RIfcbd638_7177, \9235_9534 );
and \U$7860 ( \16682_16981 , RIfc44fa8_5807, \9237_9536 );
and \U$7861 ( \16683_16982 , RIfe8e5f0_7964, \9239_9538 );
and \U$7862 ( \16684_16983 , RIfe8e1b8_7961, \9241_9540 );
and \U$7863 ( \16685_16984 , RIf1488f8_5285, \9243_9542 );
and \U$7864 ( \16686_16985 , RIf147818_5273, \9245_9544 );
and \U$7865 ( \16687_16986 , RIfe8e050_7960, \9247_9546 );
and \U$7866 ( \16688_16987 , RIfe8e488_7963, \9249_9548 );
and \U$7867 ( \16689_16988 , RIf146e40_5266, \9251_9550 );
and \U$7868 ( \16690_16989 , RIf146030_5256, \9253_9552 );
and \U$7869 ( \16691_16990 , RIfe8dee8_7959, \9255_9554 );
and \U$7870 ( \16692_16991 , RIfe8e320_7962, \9257_9556 );
and \U$7871 ( \16693_16992 , RIe1a7dc8_3287, \9259_9558 );
and \U$7872 ( \16694_16993 , RIe1a50c8_3255, \9261_9560 );
and \U$7873 ( \16695_16994 , RIe1a23c8_3223, \9263_9562 );
and \U$7874 ( \16696_16995 , RIe19f6c8_3191, \9265_9564 );
and \U$7875 ( \16697_16996 , RIe18bbc8_2967, \9267_9566 );
and \U$7876 ( \16698_16997 , RIe1780c8_2743, \9269_9568 );
and \U$7877 ( \16699_16998 , RIe225a20_4718, \9271_9570 );
and \U$7878 ( \16700_16999 , RIe21a620_4590, \9273_9572 );
and \U$7879 ( \16701_17000 , RIe203e20_4334, \9275_9574 );
and \U$7880 ( \16702_17001 , RIe1fde80_4266, \9277_9576 );
and \U$7881 ( \16703_17002 , RIe1f7238_4189, \9279_9578 );
and \U$7882 ( \16704_17003 , RIe1efd80_4106, \9281_9580 );
and \U$7883 ( \16705_17004 , RIe1d4288_3791, \9283_9582 );
and \U$7884 ( \16706_17005 , RIe1bad88_3503, \9285_9584 );
and \U$7885 ( \16707_17006 , RIe1adc00_3354, \9287_9586 );
and \U$7886 ( \16708_17007 , RIe170238_2653, \9289_9588 );
or \U$7887 ( \16709_17008 , \16645_16944 , \16646_16945 , \16647_16946 , \16648_16947 , \16649_16948 , \16650_16949 , \16651_16950 , \16652_16951 , \16653_16952 , \16654_16953 , \16655_16954 , \16656_16955 , \16657_16956 , \16658_16957 , \16659_16958 , \16660_16959 , \16661_16960 , \16662_16961 , \16663_16962 , \16664_16963 , \16665_16964 , \16666_16965 , \16667_16966 , \16668_16967 , \16669_16968 , \16670_16969 , \16671_16970 , \16672_16971 , \16673_16972 , \16674_16973 , \16675_16974 , \16676_16975 , \16677_16976 , \16678_16977 , \16679_16978 , \16680_16979 , \16681_16980 , \16682_16981 , \16683_16982 , \16684_16983 , \16685_16984 , \16686_16985 , \16687_16986 , \16688_16987 , \16689_16988 , \16690_16989 , \16691_16990 , \16692_16991 , \16693_16992 , \16694_16993 , \16695_16994 , \16696_16995 , \16697_16996 , \16698_16997 , \16699_16998 , \16700_16999 , \16701_17000 , \16702_17001 , \16703_17002 , \16704_17003 , \16705_17004 , \16706_17005 , \16707_17006 , \16708_17007 );
or \U$7888 ( \16710_17009 , \16644_16943 , \16709_17008 );
_DC \g3cbc/U$1 ( \16711 , \16710_17009 , \9298_9597 );
buf \U$7889 ( \16712_17011 , \16711 );
xor \U$7890 ( \16713_17012 , \16579_16878 , \16712_17011 );
and \U$7891 ( \16714_17013 , RIdec45c8_698, \8760_9059 );
and \U$7892 ( \16715_17014 , RIdec18c8_666, \8762_9061 );
and \U$7893 ( \16716_17015 , RIfce85e0_7666, \8764_9063 );
and \U$7894 ( \16717_17016 , RIdebebc8_634, \8766_9065 );
and \U$7895 ( \16718_17017 , RIfcb8bb0_7124, \8768_9067 );
and \U$7896 ( \16719_17018 , RIdebbec8_602, \8770_9069 );
and \U$7897 ( \16720_17019 , RIdeb91c8_570, \8772_9071 );
and \U$7898 ( \16721_17020 , RIdeb64c8_538, \8774_9073 );
and \U$7899 ( \16722_17021 , RIfc85d78_6545, \8776_9075 );
and \U$7900 ( \16723_17022 , RIdeb0ac8_474, \8778_9077 );
and \U$7901 ( \16724_17023 , RIfc85aa8_6543, \8780_9079 );
and \U$7902 ( \16725_17024 , RIdeaddc8_442, \8782_9081 );
and \U$7903 ( \16726_17025 , RIfc4d3d8_5901, \8784_9083 );
and \U$7904 ( \16727_17026 , RIdea8350_410, \8786_9085 );
and \U$7905 ( \16728_17027 , RIdea1a50_378, \8788_9087 );
and \U$7906 ( \16729_17028 , RIde9b150_346, \8790_9089 );
and \U$7907 ( \16730_17029 , RIfc85ee0_6546, \8792_9091 );
and \U$7908 ( \16731_17030 , RIfc9c9b0_6804, \8794_9093 );
and \U$7909 ( \16732_17031 , RIfce13f8_7585, \8796_9095 );
and \U$7910 ( \16733_17032 , RIfcb8778_7121, \8798_9097 );
and \U$7911 ( \16734_17033 , RIfe8d510_7952, \8800_9099 );
and \U$7912 ( \16735_17034 , RIfe8d3a8_7951, \8802_9101 );
and \U$7913 ( \16736_17035 , RIde886b8_255, \8804_9103 );
and \U$7914 ( \16737_17036 , RIde841d0_234, \8806_9105 );
and \U$7915 ( \16738_17037 , RIde806c0_216, \8808_9107 );
and \U$7916 ( \16739_17038 , RIfcb8070_7116, \8810_9109 );
and \U$7917 ( \16740_17039 , RIfce1128_7583, \8812_9111 );
and \U$7918 ( \16741_17040 , RIfc9c140_6798, \8814_9113 );
and \U$7919 ( \16742_17041 , RIee38d10_5105, \8816_9115 );
and \U$7920 ( \16743_17042 , RIe16ac70_2592, \8818_9117 );
and \U$7921 ( \16744_17043 , RIfc850d0_6536, \8820_9119 );
and \U$7922 ( \16745_17044 , RIe167160_2550, \8822_9121 );
and \U$7923 ( \16746_17045 , RIe1645c8_2519, \8824_9123 );
and \U$7924 ( \16747_17046 , RIe1618c8_2487, \8826_9125 );
and \U$7925 ( \16748_17047 , RIee36b50_5081, \8828_9127 );
and \U$7926 ( \16749_17048 , RIe15ebc8_2455, \8830_9129 );
and \U$7927 ( \16750_17049 , RIee35d40_5071, \8832_9131 );
and \U$7928 ( \16751_17050 , RIe15bec8_2423, \8834_9133 );
and \U$7929 ( \16752_17051 , RIe1564c8_2359, \8836_9135 );
and \U$7930 ( \16753_17052 , RIe1537c8_2327, \8838_9137 );
and \U$7931 ( \16754_17053 , RIfc3ef90_5742, \8840_9139 );
and \U$7932 ( \16755_17054 , RIe150ac8_2295, \8842_9141 );
and \U$7933 ( \16756_17055 , RIfe8d7e0_7954, \8844_9143 );
and \U$7934 ( \16757_17056 , RIe14ddc8_2263, \8846_9145 );
and \U$7935 ( \16758_17057 , RIfce0fc0_7582, \8848_9147 );
and \U$7936 ( \16759_17058 , RIe14b0c8_2231, \8850_9149 );
and \U$7937 ( \16760_17059 , RIe1483c8_2199, \8852_9151 );
and \U$7938 ( \16761_17060 , RIe1456c8_2167, \8854_9153 );
and \U$7939 ( \16762_17061 , RIee33e50_5049, \8856_9155 );
and \U$7940 ( \16763_17062 , RIee32c08_5036, \8858_9157 );
and \U$7941 ( \16764_17063 , RIee319c0_5023, \8860_9159 );
and \U$7942 ( \16765_17064 , RIee30d18_5014, \8862_9161 );
and \U$7943 ( \16766_17065 , RIfe8cf70_7948, \8864_9163 );
and \U$7944 ( \16767_17066 , RIfe8ce08_7947, \8866_9165 );
and \U$7945 ( \16768_17067 , RIfe8d240_7950, \8868_9167 );
and \U$7946 ( \16769_17068 , RIfe8d0d8_7949, \8870_9169 );
and \U$7947 ( \16770_17069 , RIfce9dc8_7683, \8872_9171 );
and \U$7948 ( \16771_17070 , RIee2ef90_4993, \8874_9173 );
and \U$7949 ( \16772_17071 , RIfce51d8_7629, \8876_9175 );
and \U$7950 ( \16773_17072 , RIee2cdd0_4969, \8878_9177 );
and \U$7951 ( \16774_17073 , RIdf34af8_1976, \8880_9179 );
and \U$7952 ( \16775_17074 , RIfe8d678_7953, \8882_9181 );
and \U$7953 ( \16776_17075 , RIdf30610_1927, \8884_9183 );
and \U$7954 ( \16777_17076 , RIdf2e720_1905, \8886_9185 );
or \U$7955 ( \16778_17077 , \16714_17013 , \16715_17014 , \16716_17015 , \16717_17016 , \16718_17017 , \16719_17018 , \16720_17019 , \16721_17020 , \16722_17021 , \16723_17022 , \16724_17023 , \16725_17024 , \16726_17025 , \16727_17026 , \16728_17027 , \16729_17028 , \16730_17029 , \16731_17030 , \16732_17031 , \16733_17032 , \16734_17033 , \16735_17034 , \16736_17035 , \16737_17036 , \16738_17037 , \16739_17038 , \16740_17039 , \16741_17040 , \16742_17041 , \16743_17042 , \16744_17043 , \16745_17044 , \16746_17045 , \16747_17046 , \16748_17047 , \16749_17048 , \16750_17049 , \16751_17050 , \16752_17051 , \16753_17052 , \16754_17053 , \16755_17054 , \16756_17055 , \16757_17056 , \16758_17057 , \16759_17058 , \16760_17059 , \16761_17060 , \16762_17061 , \16763_17062 , \16764_17063 , \16765_17064 , \16766_17065 , \16767_17066 , \16768_17067 , \16769_17068 , \16770_17069 , \16771_17070 , \16772_17071 , \16773_17072 , \16774_17073 , \16775_17074 , \16776_17075 , \16777_17076 );
and \U$7956 ( \16779_17078 , RIee2b318_4950, \8889_9188 );
and \U$7957 ( \16780_17079 , RIee29c98_4934, \8891_9190 );
and \U$7958 ( \16781_17080 , RIee28780_4919, \8893_9192 );
and \U$7959 ( \16782_17081 , RIee27538_4906, \8895_9194 );
and \U$7960 ( \16783_17082 , RIdf299c8_1850, \8897_9196 );
and \U$7961 ( \16784_17083 , RIdf276a0_1825, \8899_9198 );
and \U$7962 ( \16785_17084 , RIdf25918_1804, \8901_9200 );
and \U$7963 ( \16786_17085 , RIdf23cf8_1784, \8903_9202 );
and \U$7964 ( \16787_17086 , RIfc83ff0_6524, \8905_9204 );
and \U$7965 ( \16788_17087 , RIfcb73c8_7107, \8907_9206 );
and \U$7966 ( \16789_17088 , RIfc51320_5946, \8909_9208 );
and \U$7967 ( \16790_17089 , RIfcdaa80_7510, \8911_9210 );
and \U$7968 ( \16791_17090 , RIfc83d20_6522, \8913_9212 );
and \U$7969 ( \16792_17091 , RIdf1ee38_1728, \8915_9214 );
and \U$7970 ( \16793_17092 , RIfc51b90_5952, \8917_9216 );
and \U$7971 ( \16794_17093 , RIdf18a60_1657, \8919_9218 );
and \U$7972 ( \16795_17094 , RIdf16198_1628, \8921_9220 );
and \U$7973 ( \16796_17095 , RIdf13498_1596, \8923_9222 );
and \U$7974 ( \16797_17096 , RIdf10798_1564, \8925_9224 );
and \U$7975 ( \16798_17097 , RIdf0da98_1532, \8927_9226 );
and \U$7976 ( \16799_17098 , RIdf0ad98_1500, \8929_9228 );
and \U$7977 ( \16800_17099 , RIdf08098_1468, \8931_9230 );
and \U$7978 ( \16801_17100 , RIdf05398_1436, \8933_9232 );
and \U$7979 ( \16802_17101 , RIdf02698_1404, \8935_9234 );
and \U$7980 ( \16803_17102 , RIdefcc98_1340, \8937_9236 );
and \U$7981 ( \16804_17103 , RIdef9f98_1308, \8939_9238 );
and \U$7982 ( \16805_17104 , RIdef7298_1276, \8941_9240 );
and \U$7983 ( \16806_17105 , RIdef4598_1244, \8943_9242 );
and \U$7984 ( \16807_17106 , RIdef1898_1212, \8945_9244 );
and \U$7985 ( \16808_17107 , RIdeeeb98_1180, \8947_9246 );
and \U$7986 ( \16809_17108 , RIdeebe98_1148, \8949_9248 );
and \U$7987 ( \16810_17109 , RIdee9198_1116, \8951_9250 );
and \U$7988 ( \16811_17110 , RIee25210_4881, \8953_9252 );
and \U$7989 ( \16812_17111 , RIee24400_4871, \8955_9254 );
and \U$7990 ( \16813_17112 , RIee238c0_4863, \8957_9256 );
and \U$7991 ( \16814_17113 , RIee22ee8_4856, \8959_9258 );
and \U$7992 ( \16815_17114 , RIfe8cca0_7946, \8961_9260 );
and \U$7993 ( \16816_17115 , RIdee2118_1036, \8963_9262 );
and \U$7994 ( \16817_17116 , RIfe8cb38_7945, \8965_9264 );
and \U$7995 ( \16818_17117 , RIdeddf00_989, \8967_9266 );
and \U$7996 ( \16819_17118 , RIfcc5a68_7271, \8969_9268 );
and \U$7997 ( \16820_17119 , RIee21f70_4845, \8971_9270 );
and \U$7998 ( \16821_17120 , RIfcb6cc0_7102, \8973_9272 );
and \U$7999 ( \16822_17121 , RIee20e90_4833, \8975_9274 );
and \U$8000 ( \16823_17122 , RIded8c08_930, \8977_9276 );
and \U$8001 ( \16824_17123 , RIded6778_904, \8979_9278 );
and \U$8002 ( \16825_17124 , RIded4720_881, \8981_9280 );
and \U$8003 ( \16826_17125 , RIded23f8_856, \8983_9282 );
and \U$8004 ( \16827_17126 , RIdecf9c8_826, \8985_9284 );
and \U$8005 ( \16828_17127 , RIdecccc8_794, \8987_9286 );
and \U$8006 ( \16829_17128 , RIdec9fc8_762, \8989_9288 );
and \U$8007 ( \16830_17129 , RIdec72c8_730, \8991_9290 );
and \U$8008 ( \16831_17130 , RIdeb37c8_506, \8993_9292 );
and \U$8009 ( \16832_17131 , RIde94850_314, \8995_9294 );
and \U$8010 ( \16833_17132 , RIe16d3d0_2620, \8997_9296 );
and \U$8011 ( \16834_17133 , RIe1591c8_2391, \8999_9298 );
and \U$8012 ( \16835_17134 , RIe1429c8_2135, \9001_9300 );
and \U$8013 ( \16836_17135 , RIdf373c0_2005, \9003_9302 );
and \U$8014 ( \16837_17136 , RIdf2ba20_1873, \9005_9304 );
and \U$8015 ( \16838_17137 , RIdf1c2a0_1697, \9007_9306 );
and \U$8016 ( \16839_17138 , RIdeff998_1372, \9009_9308 );
and \U$8017 ( \16840_17139 , RIdee6498_1084, \9011_9310 );
and \U$8018 ( \16841_17140 , RIdedb200_957, \9013_9312 );
and \U$8019 ( \16842_17141 , RIde7a798_187, \9015_9314 );
or \U$8020 ( \16843_17142 , \16779_17078 , \16780_17079 , \16781_17080 , \16782_17081 , \16783_17082 , \16784_17083 , \16785_17084 , \16786_17085 , \16787_17086 , \16788_17087 , \16789_17088 , \16790_17089 , \16791_17090 , \16792_17091 , \16793_17092 , \16794_17093 , \16795_17094 , \16796_17095 , \16797_17096 , \16798_17097 , \16799_17098 , \16800_17099 , \16801_17100 , \16802_17101 , \16803_17102 , \16804_17103 , \16805_17104 , \16806_17105 , \16807_17106 , \16808_17107 , \16809_17108 , \16810_17109 , \16811_17110 , \16812_17111 , \16813_17112 , \16814_17113 , \16815_17114 , \16816_17115 , \16817_17116 , \16818_17117 , \16819_17118 , \16820_17119 , \16821_17120 , \16822_17121 , \16823_17122 , \16824_17123 , \16825_17124 , \16826_17125 , \16827_17126 , \16828_17127 , \16829_17128 , \16830_17129 , \16831_17130 , \16832_17131 , \16833_17132 , \16834_17133 , \16835_17134 , \16836_17135 , \16837_17136 , \16838_17137 , \16839_17138 , \16840_17139 , \16841_17140 , \16842_17141 );
or \U$8021 ( \16844_17143 , \16778_17077 , \16843_17142 );
_DC \g2c14/U$1 ( \16845 , \16844_17143 , \9024_9323 );
buf \U$8022 ( \16846_17145 , \16845 );
and \U$8023 ( \16847_17146 , RIe19c860_3158, \9034_9333 );
and \U$8024 ( \16848_17147 , RIe199b60_3126, \9036_9335 );
and \U$8025 ( \16849_17148 , RIf145220_5246, \9038_9337 );
and \U$8026 ( \16850_17149 , RIe196e60_3094, \9040_9339 );
and \U$8027 ( \16851_17150 , RIf144140_5234, \9042_9341 );
and \U$8028 ( \16852_17151 , RIe194160_3062, \9044_9343 );
and \U$8029 ( \16853_17152 , RIe191460_3030, \9046_9345 );
and \U$8030 ( \16854_17153 , RIe18e760_2998, \9048_9347 );
and \U$8031 ( \16855_17154 , RIe188d60_2934, \9050_9349 );
and \U$8032 ( \16856_17155 , RIe186060_2902, \9052_9351 );
and \U$8033 ( \16857_17156 , RIf1431c8_5223, \9054_9353 );
and \U$8034 ( \16858_17157 , RIe183360_2870, \9056_9355 );
and \U$8035 ( \16859_17158 , RIf142ac0_5218, \9058_9357 );
and \U$8036 ( \16860_17159 , RIe180660_2838, \9060_9359 );
and \U$8037 ( \16861_17160 , RIe17d960_2806, \9062_9361 );
and \U$8038 ( \16862_17161 , RIe17ac60_2774, \9064_9363 );
and \U$8039 ( \16863_17162 , RIf141cb0_5208, \9066_9365 );
and \U$8040 ( \16864_17163 , RIf140798_5193, \9068_9367 );
and \U$8041 ( \16865_17164 , RIf13ff28_5187, \9070_9369 );
and \U$8042 ( \16866_17165 , RIfe8be90_7936, \9072_9371 );
and \U$8043 ( \16867_17166 , RIfceb880_7702, \9074_9373 );
and \U$8044 ( \16868_17167 , RIf13eb78_5173, \9076_9375 );
and \U$8045 ( \16869_17168 , RIee3e008_5164, \9078_9377 );
and \U$8046 ( \16870_17169 , RIee3cdc0_5151, \9080_9379 );
and \U$8047 ( \16871_17170 , RIee3bb78_5138, \9082_9381 );
and \U$8048 ( \16872_17171 , RIee3aa98_5126, \9084_9383 );
and \U$8049 ( \16873_17172 , RIee396e8_5112, \9086_9385 );
and \U$8050 ( \16874_17173 , RIe172c68_2683, \9088_9387 );
and \U$8051 ( \16875_17174 , RIf16fac0_5730, \9090_9389 );
and \U$8052 ( \16876_17175 , RIf16ef80_5722, \9092_9391 );
and \U$8053 ( \16877_17176 , RIf16dbd0_5708, \9094_9393 );
and \U$8054 ( \16878_17177 , RIfcc4af0_7260, \9096_9395 );
and \U$8055 ( \16879_17178 , RIf16c820_5694, \9098_9397 );
and \U$8056 ( \16880_17179 , RIe222bb8_4685, \9100_9399 );
and \U$8057 ( \16881_17180 , RIf16b740_5682, \9102_9401 );
and \U$8058 ( \16882_17181 , RIe21feb8_4653, \9104_9403 );
and \U$8059 ( \16883_17182 , RIf16a7c8_5671, \9106_9405 );
and \U$8060 ( \16884_17183 , RIe21d1b8_4621, \9108_9407 );
and \U$8061 ( \16885_17184 , RIe2177b8_4557, \9110_9409 );
and \U$8062 ( \16886_17185 , RIe214ab8_4525, \9112_9411 );
and \U$8063 ( \16887_17186 , RIfe8c430_7940, \9114_9413 );
and \U$8064 ( \16888_17187 , RIe211db8_4493, \9116_9415 );
and \U$8065 ( \16889_17188 , RIf1688d8_5649, \9118_9417 );
and \U$8066 ( \16890_17189 , RIe20f0b8_4461, \9120_9419 );
and \U$8067 ( \16891_17190 , RIf167960_5638, \9122_9421 );
and \U$8068 ( \16892_17191 , RIe20c3b8_4429, \9124_9423 );
and \U$8069 ( \16893_17192 , RIe2096b8_4397, \9126_9425 );
and \U$8070 ( \16894_17193 , RIe2069b8_4365, \9128_9427 );
and \U$8071 ( \16895_17194 , RIf1669e8_5627, \9130_9429 );
and \U$8072 ( \16896_17195 , RIf165908_5615, \9132_9431 );
and \U$8073 ( \16897_17196 , RIfe8c9d0_7944, \9134_9433 );
and \U$8074 ( \16898_17197 , RIfe8c700_7942, \9136_9435 );
and \U$8075 ( \16899_17198 , RIfc9c578_6801, \9138_9437 );
and \U$8076 ( \16900_17199 , RIf163ce8_5595, \9140_9439 );
and \U$8077 ( \16901_17200 , RIf162d70_5584, \9142_9441 );
and \U$8078 ( \16902_17201 , RIf161588_5567, \9144_9443 );
and \U$8079 ( \16903_17202 , RIf15f698_5545, \9146_9445 );
and \U$8080 ( \16904_17203 , RIf15d910_5524, \9148_9447 );
and \U$8081 ( \16905_17204 , RIfe8c598_7941, \9150_9449 );
and \U$8082 ( \16906_17205 , RIfe8c868_7943, \9152_9451 );
and \U$8083 ( \16907_17206 , RIf15c3f8_5509, \9154_9453 );
and \U$8084 ( \16908_17207 , RIf15aee0_5494, \9156_9455 );
and \U$8085 ( \16909_17208 , RIf15a0d0_5484, \9158_9457 );
and \U$8086 ( \16910_17209 , RIf1596f8_5477, \9160_9459 );
or \U$8087 ( \16911_17210 , \16847_17146 , \16848_17147 , \16849_17148 , \16850_17149 , \16851_17150 , \16852_17151 , \16853_17152 , \16854_17153 , \16855_17154 , \16856_17155 , \16857_17156 , \16858_17157 , \16859_17158 , \16860_17159 , \16861_17160 , \16862_17161 , \16863_17162 , \16864_17163 , \16865_17164 , \16866_17165 , \16867_17166 , \16868_17167 , \16869_17168 , \16870_17169 , \16871_17170 , \16872_17171 , \16873_17172 , \16874_17173 , \16875_17174 , \16876_17175 , \16877_17176 , \16878_17177 , \16879_17178 , \16880_17179 , \16881_17180 , \16882_17181 , \16883_17182 , \16884_17183 , \16885_17184 , \16886_17185 , \16887_17186 , \16888_17187 , \16889_17188 , \16890_17189 , \16891_17190 , \16892_17191 , \16893_17192 , \16894_17193 , \16895_17194 , \16896_17195 , \16897_17196 , \16898_17197 , \16899_17198 , \16900_17199 , \16901_17200 , \16902_17201 , \16903_17202 , \16904_17203 , \16905_17204 , \16906_17205 , \16907_17206 , \16908_17207 , \16909_17208 , \16910_17209 );
and \U$8088 ( \16912_17211 , RIf158618_5465, \9163_9462 );
and \U$8089 ( \16913_17212 , RIf1573d0_5452, \9165_9464 );
and \U$8090 ( \16914_17213 , RIf156b60_5446, \9167_9466 );
and \U$8091 ( \16915_17214 , RIfec1f68_8327, \9169_9468 );
and \U$8092 ( \16916_17215 , RIf155eb8_5437, \9171_9470 );
and \U$8093 ( \16917_17216 , RIf155378_5429, \9173_9472 );
and \U$8094 ( \16918_17217 , RIf153fc8_5415, \9175_9474 );
and \U$8095 ( \16919_17218 , RIfe8bff8_7937, \9177_9476 );
and \U$8096 ( \16920_17219 , RIf152948_5399, \9179_9478 );
and \U$8097 ( \16921_17220 , RIf151598_5385, \9181_9480 );
and \U$8098 ( \16922_17221 , RIf150080_5370, \9183_9482 );
and \U$8099 ( \16923_17222 , RIfe8c2c8_7939, \9185_9484 );
and \U$8100 ( \16924_17223 , RIf14f270_5360, \9187_9486 );
and \U$8101 ( \16925_17224 , RIfc503a8_5935, \9189_9488 );
and \U$8102 ( \16926_17225 , RIf14d650_5340, \9191_9490 );
and \U$8103 ( \16927_17226 , RIfe8c160_7938, \9193_9492 );
and \U$8104 ( \16928_17227 , RIe1ea920_4046, \9195_9494 );
and \U$8105 ( \16929_17228 , RIe1e7c20_4014, \9197_9496 );
and \U$8106 ( \16930_17229 , RIe1e4f20_3982, \9199_9498 );
and \U$8107 ( \16931_17230 , RIe1e2220_3950, \9201_9500 );
and \U$8108 ( \16932_17231 , RIe1df520_3918, \9203_9502 );
and \U$8109 ( \16933_17232 , RIe1dc820_3886, \9205_9504 );
and \U$8110 ( \16934_17233 , RIe1d9b20_3854, \9207_9506 );
and \U$8111 ( \16935_17234 , RIe1d6e20_3822, \9209_9508 );
and \U$8112 ( \16936_17235 , RIe1d1420_3758, \9211_9510 );
and \U$8113 ( \16937_17236 , RIe1ce720_3726, \9213_9512 );
and \U$8114 ( \16938_17237 , RIe1cba20_3694, \9215_9514 );
and \U$8115 ( \16939_17238 , RIe1c8d20_3662, \9217_9516 );
and \U$8116 ( \16940_17239 , RIe1c6020_3630, \9219_9518 );
and \U$8117 ( \16941_17240 , RIe1c3320_3598, \9221_9520 );
and \U$8118 ( \16942_17241 , RIe1c0620_3566, \9223_9522 );
and \U$8119 ( \16943_17242 , RIe1bd920_3534, \9225_9524 );
and \U$8120 ( \16944_17243 , RIf14c2a0_5326, \9227_9526 );
and \U$8121 ( \16945_17244 , RIf14aef0_5312, \9229_9528 );
and \U$8122 ( \16946_17245 , RIe1b88f8_3477, \9231_9530 );
and \U$8123 ( \16947_17246 , RIe1b68a0_3454, \9233_9532 );
and \U$8124 ( \16948_17247 , RIfcd4db0_7444, \9235_9534 );
and \U$8125 ( \16949_17248 , RIfc4ebc0_5918, \9237_9536 );
and \U$8126 ( \16950_17249 , RIfec1e00_8326, \9239_9538 );
and \U$8127 ( \16951_17250 , RIfe8bd28_7935, \9241_9540 );
and \U$8128 ( \16952_17251 , RIf148790_5284, \9243_9542 );
and \U$8129 ( \16953_17252 , RIf1476b0_5272, \9245_9544 );
and \U$8130 ( \16954_17253 , RIfe8ba58_7933, \9247_9546 );
and \U$8131 ( \16955_17254 , RIfec1b30_8324, \9249_9548 );
and \U$8132 ( \16956_17255 , RIfc4e788_5915, \9251_9550 );
and \U$8133 ( \16957_17256 , RIfcb8e80_7126, \9253_9552 );
and \U$8134 ( \16958_17257 , RIfe8bbc0_7934, \9255_9554 );
and \U$8135 ( \16959_17258 , RIfec1c98_8325, \9257_9556 );
and \U$8136 ( \16960_17259 , RIe1a7c60_3286, \9259_9558 );
and \U$8137 ( \16961_17260 , RIe1a4f60_3254, \9261_9560 );
and \U$8138 ( \16962_17261 , RIe1a2260_3222, \9263_9562 );
and \U$8139 ( \16963_17262 , RIe19f560_3190, \9265_9564 );
and \U$8140 ( \16964_17263 , RIe18ba60_2966, \9267_9566 );
and \U$8141 ( \16965_17264 , RIe177f60_2742, \9269_9568 );
and \U$8142 ( \16966_17265 , RIe2258b8_4717, \9271_9570 );
and \U$8143 ( \16967_17266 , RIe21a4b8_4589, \9273_9572 );
and \U$8144 ( \16968_17267 , RIe203cb8_4333, \9275_9574 );
and \U$8145 ( \16969_17268 , RIe1fdd18_4265, \9277_9576 );
and \U$8146 ( \16970_17269 , RIe1f70d0_4188, \9279_9578 );
and \U$8147 ( \16971_17270 , RIe1efc18_4105, \9281_9580 );
and \U$8148 ( \16972_17271 , RIe1d4120_3790, \9283_9582 );
and \U$8149 ( \16973_17272 , RIe1bac20_3502, \9285_9584 );
and \U$8150 ( \16974_17273 , RIe1ada98_3353, \9287_9586 );
and \U$8151 ( \16975_17274 , RIe1700d0_2652, \9289_9588 );
or \U$8152 ( \16976_17275 , \16912_17211 , \16913_17212 , \16914_17213 , \16915_17214 , \16916_17215 , \16917_17216 , \16918_17217 , \16919_17218 , \16920_17219 , \16921_17220 , \16922_17221 , \16923_17222 , \16924_17223 , \16925_17224 , \16926_17225 , \16927_17226 , \16928_17227 , \16929_17228 , \16930_17229 , \16931_17230 , \16932_17231 , \16933_17232 , \16934_17233 , \16935_17234 , \16936_17235 , \16937_17236 , \16938_17237 , \16939_17238 , \16940_17239 , \16941_17240 , \16942_17241 , \16943_17242 , \16944_17243 , \16945_17244 , \16946_17245 , \16947_17246 , \16948_17247 , \16949_17248 , \16950_17249 , \16951_17250 , \16952_17251 , \16953_17252 , \16954_17253 , \16955_17254 , \16956_17255 , \16957_17256 , \16958_17257 , \16959_17258 , \16960_17259 , \16961_17260 , \16962_17261 , \16963_17262 , \16964_17263 , \16965_17264 , \16966_17265 , \16967_17266 , \16968_17267 , \16969_17268 , \16970_17269 , \16971_17270 , \16972_17271 , \16973_17272 , \16974_17273 , \16975_17274 );
or \U$8153 ( \16977_17276 , \16911_17210 , \16976_17275 );
_DC \g3d41/U$1 ( \16978 , \16977_17276 , \9298_9597 );
buf \U$8154 ( \16979_17278 , \16978 );
and \U$8155 ( \16980_17279 , \16846_17145 , \16979_17278 );
and \U$8156 ( \16981_17280 , \15222_15521 , \15355_15654 );
and \U$8157 ( \16982_17281 , \15355_15654 , \15630_15929 );
and \U$8158 ( \16983_17282 , \15222_15521 , \15630_15929 );
or \U$8159 ( \16984_17283 , \16981_17280 , \16982_17281 , \16983_17282 );
and \U$8160 ( \16985_17284 , \16979_17278 , \16984_17283 );
and \U$8161 ( \16986_17285 , \16846_17145 , \16984_17283 );
or \U$8162 ( \16987_17286 , \16980_17279 , \16985_17284 , \16986_17285 );
xor \U$8163 ( \16988_17287 , \16713_17012 , \16987_17286 );
buf g4430_GF_PartitionCandidate( \16989_17288_nG4430 , \16988_17287 );
xor \U$8164 ( \16990_17289 , \16846_17145 , \16979_17278 );
xor \U$8165 ( \16991_17290 , \16990_17289 , \16984_17283 );
buf g4433_GF_PartitionCandidate( \16992_17291_nG4433 , \16991_17290 );
nand \U$8166 ( \16993_17292 , \16992_17291_nG4433 , \15632_15931_nG4436 );
and \U$8167 ( \16994_17293 , \16989_17288_nG4430 , \16993_17292 );
xor \U$8168 ( \16995_17294 , \16992_17291_nG4433 , \15632_15931_nG4436 );
and \U$8173 ( \16996_17298 , \16995_17294 , \10392_10694_nG9c0e );
or \U$8174 ( \16997_17299 , 1'b0 , \16996_17298 );
xor \U$8175 ( \16998_17300 , \16994_17293 , \16997_17299 );
xor \U$8176 ( \16999_17301 , \16994_17293 , \16998_17300 );
buf \U$8177 ( \17000_17302 , \16999_17301 );
buf \U$8178 ( \17001_17303 , \17000_17302 );
and \U$8179 ( \17002_17304 , \16446_16745 , \17001_17303 );
and \U$8180 ( \17003_17305 , \16420_16719 , \16422_16721 );
and \U$8181 ( \17004_17306 , \16420_16719 , \16429_16728 );
and \U$8182 ( \17005_17307 , \16422_16721 , \16429_16728 );
or \U$8183 ( \17006_17308 , \17003_17305 , \17004_17306 , \17005_17307 );
buf \U$8184 ( \17007_17309 , \17006_17308 );
and \U$8185 ( \17008_17310 , \16405_15940 , \10693_10995_nG9c0b );
and \U$8186 ( \17009_17311 , \15638_15937 , \10981_11283_nG9c08 );
or \U$8187 ( \17010_17312 , \17008_17310 , \17009_17311 );
xor \U$8188 ( \17011_17313 , \15637_15936 , \17010_17312 );
buf \U$8189 ( \17012_17314 , \17011_17313 );
buf \U$8191 ( \17013_17315 , \17012_17314 );
and \U$8192 ( \17014_17316 , \14710_14631 , \11299_11598_nG9c05 );
and \U$8193 ( \17015_17317 , \14329_14628 , \12168_12470_nG9c02 );
or \U$8194 ( \17016_17318 , \17014_17316 , \17015_17317 );
xor \U$8195 ( \17017_17319 , \14328_14627 , \17016_17318 );
buf \U$8196 ( \17018_17320 , \17017_17319 );
buf \U$8198 ( \17019_17321 , \17018_17320 );
xor \U$8199 ( \17020_17322 , \17013_17315 , \17019_17321 );
buf \U$8200 ( \17021_17323 , \17020_17322 );
and \U$8201 ( \17022_17324 , \16394_16696 , \16400_16702 );
buf \U$8202 ( \17023_17325 , \17022_17324 );
xor \U$8203 ( \17024_17326 , \17021_17323 , \17023_17325 );
and \U$8204 ( \17025_17327 , \13431_13370 , \12502_12801_nG9bff );
and \U$8205 ( \17026_17328 , \13068_13367 , \13403_13705_nG9bfc );
or \U$8206 ( \17027_17329 , \17025_17327 , \17026_17328 );
xor \U$8207 ( \17028_17330 , \13067_13366 , \17027_17329 );
buf \U$8208 ( \17029_17331 , \17028_17330 );
buf \U$8210 ( \17030_17332 , \17029_17331 );
xor \U$8211 ( \17031_17333 , \17024_17326 , \17030_17332 );
buf \U$8212 ( \17032_17334 , \17031_17333 );
xor \U$8213 ( \17033_17335 , \17007_17309 , \17032_17334 );
and \U$8214 ( \17034_17336 , \10411_10707 , \16378_16680_nG9bed );
and \U$8215 ( \17035_17337 , \16049_16351 , \16338_16640 );
and \U$8216 ( \17036_17338 , \16338_16640 , \16367_16669 );
and \U$8217 ( \17037_17339 , \16049_16351 , \16367_16669 );
or \U$8218 ( \17038_17340 , \17035_17337 , \17036_17338 , \17037_17339 );
and \U$8219 ( \17039_17341 , \16343_16645 , \16347_16649 );
and \U$8220 ( \17040_17342 , \16347_16649 , \16366_16668 );
and \U$8221 ( \17041_17343 , \16343_16645 , \16366_16668 );
or \U$8222 ( \17042_17344 , \17039_17341 , \17040_17342 , \17041_17343 );
and \U$8223 ( \17043_17345 , \16356_16658 , \16360_16662 );
and \U$8224 ( \17044_17346 , \16360_16662 , \16365_16667 );
and \U$8225 ( \17045_17347 , \16356_16658 , \16365_16667 );
or \U$8226 ( \17046_17348 , \17043_17345 , \17044_17346 , \17045_17347 );
and \U$8227 ( \17047_17349 , \16053_16355 , \16324_16626 );
xor \U$8228 ( \17048_17350 , \17046_17348 , \17047_17349 );
and \U$8229 ( \17049_17351 , \13725_14024 , \12491_12790 );
and \U$8230 ( \17050_17352 , \14648_14950 , \12159_12461 );
nor \U$8231 ( \17051_17353 , \17049_17351 , \17050_17352 );
xnor \U$8232 ( \17052_17354 , \17051_17353 , \12481_12780 );
xor \U$8233 ( \17053_17355 , \17048_17350 , \17052_17354 );
xor \U$8234 ( \17054_17356 , \17042_17344 , \17053_17355 );
and \U$8235 ( \17055_17357 , \16325_16627 , \16329_16631 );
and \U$8236 ( \17056_17358 , \16329_16631 , \16337_16639 );
and \U$8237 ( \17057_17359 , \16325_16627 , \16337_16639 );
or \U$8238 ( \17058_17360 , \17055_17357 , \17056_17358 , \17057_17359 );
and \U$8239 ( \17059_17361 , \16353_16655 , \10681_10983 );
and \U$8240 ( \17060_17362 , RIdec45c8_698, \9034_9333 );
and \U$8241 ( \17061_17363 , RIdec18c8_666, \9036_9335 );
and \U$8242 ( \17062_17364 , RIfce85e0_7666, \9038_9337 );
and \U$8243 ( \17063_17365 , RIdebebc8_634, \9040_9339 );
and \U$8244 ( \17064_17366 , RIfcb8bb0_7124, \9042_9341 );
and \U$8245 ( \17065_17367 , RIdebbec8_602, \9044_9343 );
and \U$8246 ( \17066_17368 , RIdeb91c8_570, \9046_9345 );
and \U$8247 ( \17067_17369 , RIdeb64c8_538, \9048_9347 );
and \U$8248 ( \17068_17370 , RIfc85d78_6545, \9050_9349 );
and \U$8249 ( \17069_17371 , RIdeb0ac8_474, \9052_9351 );
and \U$8250 ( \17070_17372 , RIfc85aa8_6543, \9054_9353 );
and \U$8251 ( \17071_17373 , RIdeaddc8_442, \9056_9355 );
and \U$8252 ( \17072_17374 , RIfc4d3d8_5901, \9058_9357 );
and \U$8253 ( \17073_17375 , RIdea8350_410, \9060_9359 );
and \U$8254 ( \17074_17376 , RIdea1a50_378, \9062_9361 );
and \U$8255 ( \17075_17377 , RIde9b150_346, \9064_9363 );
and \U$8256 ( \17076_17378 , RIfc85ee0_6546, \9066_9365 );
and \U$8257 ( \17077_17379 , RIfc9c9b0_6804, \9068_9367 );
and \U$8258 ( \17078_17380 , RIfce13f8_7585, \9070_9369 );
and \U$8259 ( \17079_17381 , RIfcb8778_7121, \9072_9371 );
and \U$8260 ( \17080_17382 , RIfe8d510_7952, \9074_9373 );
and \U$8261 ( \17081_17383 , RIfe8d3a8_7951, \9076_9375 );
and \U$8262 ( \17082_17384 , RIde886b8_255, \9078_9377 );
and \U$8263 ( \17083_17385 , RIde841d0_234, \9080_9379 );
and \U$8264 ( \17084_17386 , RIde806c0_216, \9082_9381 );
and \U$8265 ( \17085_17387 , RIfcb8070_7116, \9084_9383 );
and \U$8266 ( \17086_17388 , RIfce1128_7583, \9086_9385 );
and \U$8267 ( \17087_17389 , RIfc9c140_6798, \9088_9387 );
and \U$8268 ( \17088_17390 , RIee38d10_5105, \9090_9389 );
and \U$8269 ( \17089_17391 , RIe16ac70_2592, \9092_9391 );
and \U$8270 ( \17090_17392 , RIfc850d0_6536, \9094_9393 );
and \U$8271 ( \17091_17393 , RIe167160_2550, \9096_9395 );
and \U$8272 ( \17092_17394 , RIe1645c8_2519, \9098_9397 );
and \U$8273 ( \17093_17395 , RIe1618c8_2487, \9100_9399 );
and \U$8274 ( \17094_17396 , RIee36b50_5081, \9102_9401 );
and \U$8275 ( \17095_17397 , RIe15ebc8_2455, \9104_9403 );
and \U$8276 ( \17096_17398 , RIee35d40_5071, \9106_9405 );
and \U$8277 ( \17097_17399 , RIe15bec8_2423, \9108_9407 );
and \U$8278 ( \17098_17400 , RIe1564c8_2359, \9110_9409 );
and \U$8279 ( \17099_17401 , RIe1537c8_2327, \9112_9411 );
and \U$8280 ( \17100_17402 , RIfc3ef90_5742, \9114_9413 );
and \U$8281 ( \17101_17403 , RIe150ac8_2295, \9116_9415 );
and \U$8282 ( \17102_17404 , RIfe8d7e0_7954, \9118_9417 );
and \U$8283 ( \17103_17405 , RIe14ddc8_2263, \9120_9419 );
and \U$8284 ( \17104_17406 , RIfce0fc0_7582, \9122_9421 );
and \U$8285 ( \17105_17407 , RIe14b0c8_2231, \9124_9423 );
and \U$8286 ( \17106_17408 , RIe1483c8_2199, \9126_9425 );
and \U$8287 ( \17107_17409 , RIe1456c8_2167, \9128_9427 );
and \U$8288 ( \17108_17410 , RIee33e50_5049, \9130_9429 );
and \U$8289 ( \17109_17411 , RIee32c08_5036, \9132_9431 );
and \U$8290 ( \17110_17412 , RIee319c0_5023, \9134_9433 );
and \U$8291 ( \17111_17413 , RIee30d18_5014, \9136_9435 );
and \U$8292 ( \17112_17414 , RIfe8cf70_7948, \9138_9437 );
and \U$8293 ( \17113_17415 , RIfe8ce08_7947, \9140_9439 );
and \U$8294 ( \17114_17416 , RIfe8d240_7950, \9142_9441 );
and \U$8295 ( \17115_17417 , RIfe8d0d8_7949, \9144_9443 );
and \U$8296 ( \17116_17418 , RIfce9dc8_7683, \9146_9445 );
and \U$8297 ( \17117_17419 , RIee2ef90_4993, \9148_9447 );
and \U$8298 ( \17118_17420 , RIfce51d8_7629, \9150_9449 );
and \U$8299 ( \17119_17421 , RIee2cdd0_4969, \9152_9451 );
and \U$8300 ( \17120_17422 , RIdf34af8_1976, \9154_9453 );
and \U$8301 ( \17121_17423 , RIfe8d678_7953, \9156_9455 );
and \U$8302 ( \17122_17424 , RIdf30610_1927, \9158_9457 );
and \U$8303 ( \17123_17425 , RIdf2e720_1905, \9160_9459 );
or \U$8304 ( \17124_17426 , \17060_17362 , \17061_17363 , \17062_17364 , \17063_17365 , \17064_17366 , \17065_17367 , \17066_17368 , \17067_17369 , \17068_17370 , \17069_17371 , \17070_17372 , \17071_17373 , \17072_17374 , \17073_17375 , \17074_17376 , \17075_17377 , \17076_17378 , \17077_17379 , \17078_17380 , \17079_17381 , \17080_17382 , \17081_17383 , \17082_17384 , \17083_17385 , \17084_17386 , \17085_17387 , \17086_17388 , \17087_17389 , \17088_17390 , \17089_17391 , \17090_17392 , \17091_17393 , \17092_17394 , \17093_17395 , \17094_17396 , \17095_17397 , \17096_17398 , \17097_17399 , \17098_17400 , \17099_17401 , \17100_17402 , \17101_17403 , \17102_17404 , \17103_17405 , \17104_17406 , \17105_17407 , \17106_17408 , \17107_17409 , \17108_17410 , \17109_17411 , \17110_17412 , \17111_17413 , \17112_17414 , \17113_17415 , \17114_17416 , \17115_17417 , \17116_17418 , \17117_17419 , \17118_17420 , \17119_17421 , \17120_17422 , \17121_17423 , \17122_17424 , \17123_17425 );
and \U$8305 ( \17125_17427 , RIee2b318_4950, \9163_9462 );
and \U$8306 ( \17126_17428 , RIee29c98_4934, \9165_9464 );
and \U$8307 ( \17127_17429 , RIee28780_4919, \9167_9466 );
and \U$8308 ( \17128_17430 , RIee27538_4906, \9169_9468 );
and \U$8309 ( \17129_17431 , RIdf299c8_1850, \9171_9470 );
and \U$8310 ( \17130_17432 , RIdf276a0_1825, \9173_9472 );
and \U$8311 ( \17131_17433 , RIdf25918_1804, \9175_9474 );
and \U$8312 ( \17132_17434 , RIdf23cf8_1784, \9177_9476 );
and \U$8313 ( \17133_17435 , RIfc83ff0_6524, \9179_9478 );
and \U$8314 ( \17134_17436 , RIfcb73c8_7107, \9181_9480 );
and \U$8315 ( \17135_17437 , RIfc51320_5946, \9183_9482 );
and \U$8316 ( \17136_17438 , RIfcdaa80_7510, \9185_9484 );
and \U$8317 ( \17137_17439 , RIfc83d20_6522, \9187_9486 );
and \U$8318 ( \17138_17440 , RIdf1ee38_1728, \9189_9488 );
and \U$8319 ( \17139_17441 , RIfc51b90_5952, \9191_9490 );
and \U$8320 ( \17140_17442 , RIdf18a60_1657, \9193_9492 );
and \U$8321 ( \17141_17443 , RIdf16198_1628, \9195_9494 );
and \U$8322 ( \17142_17444 , RIdf13498_1596, \9197_9496 );
and \U$8323 ( \17143_17445 , RIdf10798_1564, \9199_9498 );
and \U$8324 ( \17144_17446 , RIdf0da98_1532, \9201_9500 );
and \U$8325 ( \17145_17447 , RIdf0ad98_1500, \9203_9502 );
and \U$8326 ( \17146_17448 , RIdf08098_1468, \9205_9504 );
and \U$8327 ( \17147_17449 , RIdf05398_1436, \9207_9506 );
and \U$8328 ( \17148_17450 , RIdf02698_1404, \9209_9508 );
and \U$8329 ( \17149_17451 , RIdefcc98_1340, \9211_9510 );
and \U$8330 ( \17150_17452 , RIdef9f98_1308, \9213_9512 );
and \U$8331 ( \17151_17453 , RIdef7298_1276, \9215_9514 );
and \U$8332 ( \17152_17454 , RIdef4598_1244, \9217_9516 );
and \U$8333 ( \17153_17455 , RIdef1898_1212, \9219_9518 );
and \U$8334 ( \17154_17456 , RIdeeeb98_1180, \9221_9520 );
and \U$8335 ( \17155_17457 , RIdeebe98_1148, \9223_9522 );
and \U$8336 ( \17156_17458 , RIdee9198_1116, \9225_9524 );
and \U$8337 ( \17157_17459 , RIee25210_4881, \9227_9526 );
and \U$8338 ( \17158_17460 , RIee24400_4871, \9229_9528 );
and \U$8339 ( \17159_17461 , RIee238c0_4863, \9231_9530 );
and \U$8340 ( \17160_17462 , RIee22ee8_4856, \9233_9532 );
and \U$8341 ( \17161_17463 , RIfe8cca0_7946, \9235_9534 );
and \U$8342 ( \17162_17464 , RIdee2118_1036, \9237_9536 );
and \U$8343 ( \17163_17465 , RIfe8cb38_7945, \9239_9538 );
and \U$8344 ( \17164_17466 , RIdeddf00_989, \9241_9540 );
and \U$8345 ( \17165_17467 , RIfcc5a68_7271, \9243_9542 );
and \U$8346 ( \17166_17468 , RIee21f70_4845, \9245_9544 );
and \U$8347 ( \17167_17469 , RIfcb6cc0_7102, \9247_9546 );
and \U$8348 ( \17168_17470 , RIee20e90_4833, \9249_9548 );
and \U$8349 ( \17169_17471 , RIded8c08_930, \9251_9550 );
and \U$8350 ( \17170_17472 , RIded6778_904, \9253_9552 );
and \U$8351 ( \17171_17473 , RIded4720_881, \9255_9554 );
and \U$8352 ( \17172_17474 , RIded23f8_856, \9257_9556 );
and \U$8353 ( \17173_17475 , RIdecf9c8_826, \9259_9558 );
and \U$8354 ( \17174_17476 , RIdecccc8_794, \9261_9560 );
and \U$8355 ( \17175_17477 , RIdec9fc8_762, \9263_9562 );
and \U$8356 ( \17176_17478 , RIdec72c8_730, \9265_9564 );
and \U$8357 ( \17177_17479 , RIdeb37c8_506, \9267_9566 );
and \U$8358 ( \17178_17480 , RIde94850_314, \9269_9568 );
and \U$8359 ( \17179_17481 , RIe16d3d0_2620, \9271_9570 );
and \U$8360 ( \17180_17482 , RIe1591c8_2391, \9273_9572 );
and \U$8361 ( \17181_17483 , RIe1429c8_2135, \9275_9574 );
and \U$8362 ( \17182_17484 , RIdf373c0_2005, \9277_9576 );
and \U$8363 ( \17183_17485 , RIdf2ba20_1873, \9279_9578 );
and \U$8364 ( \17184_17486 , RIdf1c2a0_1697, \9281_9580 );
and \U$8365 ( \17185_17487 , RIdeff998_1372, \9283_9582 );
and \U$8366 ( \17186_17488 , RIdee6498_1084, \9285_9584 );
and \U$8367 ( \17187_17489 , RIdedb200_957, \9287_9586 );
and \U$8368 ( \17188_17490 , RIde7a798_187, \9289_9588 );
or \U$8369 ( \17189_17491 , \17125_17427 , \17126_17428 , \17127_17429 , \17128_17430 , \17129_17431 , \17130_17432 , \17131_17433 , \17132_17434 , \17133_17435 , \17134_17436 , \17135_17437 , \17136_17438 , \17137_17439 , \17138_17440 , \17139_17441 , \17140_17442 , \17141_17443 , \17142_17444 , \17143_17445 , \17144_17446 , \17145_17447 , \17146_17448 , \17147_17449 , \17148_17450 , \17149_17451 , \17150_17452 , \17151_17453 , \17152_17454 , \17153_17455 , \17154_17456 , \17155_17457 , \17156_17458 , \17157_17459 , \17158_17460 , \17159_17461 , \17160_17462 , \17161_17463 , \17162_17464 , \17163_17465 , \17164_17466 , \17165_17467 , \17166_17468 , \17167_17469 , \17168_17470 , \17169_17471 , \17170_17472 , \17171_17473 , \17172_17474 , \17173_17475 , \17174_17476 , \17175_17477 , \17176_17478 , \17177_17479 , \17178_17480 , \17179_17481 , \17180_17482 , \17181_17483 , \17182_17484 , \17183_17485 , \17184_17486 , \17185_17487 , \17186_17488 , \17187_17489 , \17188_17490 );
or \U$8370 ( \17190_17492 , \17124_17426 , \17189_17491 );
_DC \g659b/U$1 ( \17191 , \17190_17492 , \9298_9597 );
and \U$8371 ( \17192_17494 , RIe19c860_3158, \8760_9059 );
and \U$8372 ( \17193_17495 , RIe199b60_3126, \8762_9061 );
and \U$8373 ( \17194_17496 , RIf145220_5246, \8764_9063 );
and \U$8374 ( \17195_17497 , RIe196e60_3094, \8766_9065 );
and \U$8375 ( \17196_17498 , RIf144140_5234, \8768_9067 );
and \U$8376 ( \17197_17499 , RIe194160_3062, \8770_9069 );
and \U$8377 ( \17198_17500 , RIe191460_3030, \8772_9071 );
and \U$8378 ( \17199_17501 , RIe18e760_2998, \8774_9073 );
and \U$8379 ( \17200_17502 , RIe188d60_2934, \8776_9075 );
and \U$8380 ( \17201_17503 , RIe186060_2902, \8778_9077 );
and \U$8381 ( \17202_17504 , RIf1431c8_5223, \8780_9079 );
and \U$8382 ( \17203_17505 , RIe183360_2870, \8782_9081 );
and \U$8383 ( \17204_17506 , RIf142ac0_5218, \8784_9083 );
and \U$8384 ( \17205_17507 , RIe180660_2838, \8786_9085 );
and \U$8385 ( \17206_17508 , RIe17d960_2806, \8788_9087 );
and \U$8386 ( \17207_17509 , RIe17ac60_2774, \8790_9089 );
and \U$8387 ( \17208_17510 , RIf141cb0_5208, \8792_9091 );
and \U$8388 ( \17209_17511 , RIf140798_5193, \8794_9093 );
and \U$8389 ( \17210_17512 , RIf13ff28_5187, \8796_9095 );
and \U$8390 ( \17211_17513 , RIfe8be90_7936, \8798_9097 );
and \U$8391 ( \17212_17514 , RIfceb880_7702, \8800_9099 );
and \U$8392 ( \17213_17515 , RIf13eb78_5173, \8802_9101 );
and \U$8393 ( \17214_17516 , RIee3e008_5164, \8804_9103 );
and \U$8394 ( \17215_17517 , RIee3cdc0_5151, \8806_9105 );
and \U$8395 ( \17216_17518 , RIee3bb78_5138, \8808_9107 );
and \U$8396 ( \17217_17519 , RIee3aa98_5126, \8810_9109 );
and \U$8397 ( \17218_17520 , RIee396e8_5112, \8812_9111 );
and \U$8398 ( \17219_17521 , RIe172c68_2683, \8814_9113 );
and \U$8399 ( \17220_17522 , RIf16fac0_5730, \8816_9115 );
and \U$8400 ( \17221_17523 , RIf16ef80_5722, \8818_9117 );
and \U$8401 ( \17222_17524 , RIf16dbd0_5708, \8820_9119 );
and \U$8402 ( \17223_17525 , RIfcc4af0_7260, \8822_9121 );
and \U$8403 ( \17224_17526 , RIf16c820_5694, \8824_9123 );
and \U$8404 ( \17225_17527 , RIe222bb8_4685, \8826_9125 );
and \U$8405 ( \17226_17528 , RIf16b740_5682, \8828_9127 );
and \U$8406 ( \17227_17529 , RIe21feb8_4653, \8830_9129 );
and \U$8407 ( \17228_17530 , RIf16a7c8_5671, \8832_9131 );
and \U$8408 ( \17229_17531 , RIe21d1b8_4621, \8834_9133 );
and \U$8409 ( \17230_17532 , RIe2177b8_4557, \8836_9135 );
and \U$8410 ( \17231_17533 , RIe214ab8_4525, \8838_9137 );
and \U$8411 ( \17232_17534 , RIfe8c430_7940, \8840_9139 );
and \U$8412 ( \17233_17535 , RIe211db8_4493, \8842_9141 );
and \U$8413 ( \17234_17536 , RIf1688d8_5649, \8844_9143 );
and \U$8414 ( \17235_17537 , RIe20f0b8_4461, \8846_9145 );
and \U$8415 ( \17236_17538 , RIf167960_5638, \8848_9147 );
and \U$8416 ( \17237_17539 , RIe20c3b8_4429, \8850_9149 );
and \U$8417 ( \17238_17540 , RIe2096b8_4397, \8852_9151 );
and \U$8418 ( \17239_17541 , RIe2069b8_4365, \8854_9153 );
and \U$8419 ( \17240_17542 , RIf1669e8_5627, \8856_9155 );
and \U$8420 ( \17241_17543 , RIf165908_5615, \8858_9157 );
and \U$8421 ( \17242_17544 , RIfe8c9d0_7944, \8860_9159 );
and \U$8422 ( \17243_17545 , RIfe8c700_7942, \8862_9161 );
and \U$8423 ( \17244_17546 , RIfc9c578_6801, \8864_9163 );
and \U$8424 ( \17245_17547 , RIf163ce8_5595, \8866_9165 );
and \U$8425 ( \17246_17548 , RIf162d70_5584, \8868_9167 );
and \U$8426 ( \17247_17549 , RIf161588_5567, \8870_9169 );
and \U$8427 ( \17248_17550 , RIf15f698_5545, \8872_9171 );
and \U$8428 ( \17249_17551 , RIf15d910_5524, \8874_9173 );
and \U$8429 ( \17250_17552 , RIfe8c598_7941, \8876_9175 );
and \U$8430 ( \17251_17553 , RIfe8c868_7943, \8878_9177 );
and \U$8431 ( \17252_17554 , RIf15c3f8_5509, \8880_9179 );
and \U$8432 ( \17253_17555 , RIf15aee0_5494, \8882_9181 );
and \U$8433 ( \17254_17556 , RIf15a0d0_5484, \8884_9183 );
and \U$8434 ( \17255_17557 , RIf1596f8_5477, \8886_9185 );
or \U$8435 ( \17256_17558 , \17192_17494 , \17193_17495 , \17194_17496 , \17195_17497 , \17196_17498 , \17197_17499 , \17198_17500 , \17199_17501 , \17200_17502 , \17201_17503 , \17202_17504 , \17203_17505 , \17204_17506 , \17205_17507 , \17206_17508 , \17207_17509 , \17208_17510 , \17209_17511 , \17210_17512 , \17211_17513 , \17212_17514 , \17213_17515 , \17214_17516 , \17215_17517 , \17216_17518 , \17217_17519 , \17218_17520 , \17219_17521 , \17220_17522 , \17221_17523 , \17222_17524 , \17223_17525 , \17224_17526 , \17225_17527 , \17226_17528 , \17227_17529 , \17228_17530 , \17229_17531 , \17230_17532 , \17231_17533 , \17232_17534 , \17233_17535 , \17234_17536 , \17235_17537 , \17236_17538 , \17237_17539 , \17238_17540 , \17239_17541 , \17240_17542 , \17241_17543 , \17242_17544 , \17243_17545 , \17244_17546 , \17245_17547 , \17246_17548 , \17247_17549 , \17248_17550 , \17249_17551 , \17250_17552 , \17251_17553 , \17252_17554 , \17253_17555 , \17254_17556 , \17255_17557 );
and \U$8436 ( \17257_17559 , RIf158618_5465, \8889_9188 );
and \U$8437 ( \17258_17560 , RIf1573d0_5452, \8891_9190 );
and \U$8438 ( \17259_17561 , RIf156b60_5446, \8893_9192 );
and \U$8439 ( \17260_17562 , RIfec1f68_8327, \8895_9194 );
and \U$8440 ( \17261_17563 , RIf155eb8_5437, \8897_9196 );
and \U$8441 ( \17262_17564 , RIf155378_5429, \8899_9198 );
and \U$8442 ( \17263_17565 , RIf153fc8_5415, \8901_9200 );
and \U$8443 ( \17264_17566 , RIfe8bff8_7937, \8903_9202 );
and \U$8444 ( \17265_17567 , RIf152948_5399, \8905_9204 );
and \U$8445 ( \17266_17568 , RIf151598_5385, \8907_9206 );
and \U$8446 ( \17267_17569 , RIf150080_5370, \8909_9208 );
and \U$8447 ( \17268_17570 , RIfe8c2c8_7939, \8911_9210 );
and \U$8448 ( \17269_17571 , RIf14f270_5360, \8913_9212 );
and \U$8449 ( \17270_17572 , RIfc503a8_5935, \8915_9214 );
and \U$8450 ( \17271_17573 , RIf14d650_5340, \8917_9216 );
and \U$8451 ( \17272_17574 , RIfe8c160_7938, \8919_9218 );
and \U$8452 ( \17273_17575 , RIe1ea920_4046, \8921_9220 );
and \U$8453 ( \17274_17576 , RIe1e7c20_4014, \8923_9222 );
and \U$8454 ( \17275_17577 , RIe1e4f20_3982, \8925_9224 );
and \U$8455 ( \17276_17578 , RIe1e2220_3950, \8927_9226 );
and \U$8456 ( \17277_17579 , RIe1df520_3918, \8929_9228 );
and \U$8457 ( \17278_17580 , RIe1dc820_3886, \8931_9230 );
and \U$8458 ( \17279_17581 , RIe1d9b20_3854, \8933_9232 );
and \U$8459 ( \17280_17582 , RIe1d6e20_3822, \8935_9234 );
and \U$8460 ( \17281_17583 , RIe1d1420_3758, \8937_9236 );
and \U$8461 ( \17282_17584 , RIe1ce720_3726, \8939_9238 );
and \U$8462 ( \17283_17585 , RIe1cba20_3694, \8941_9240 );
and \U$8463 ( \17284_17586 , RIe1c8d20_3662, \8943_9242 );
and \U$8464 ( \17285_17587 , RIe1c6020_3630, \8945_9244 );
and \U$8465 ( \17286_17588 , RIe1c3320_3598, \8947_9246 );
and \U$8466 ( \17287_17589 , RIe1c0620_3566, \8949_9248 );
and \U$8467 ( \17288_17590 , RIe1bd920_3534, \8951_9250 );
and \U$8468 ( \17289_17591 , RIf14c2a0_5326, \8953_9252 );
and \U$8469 ( \17290_17592 , RIf14aef0_5312, \8955_9254 );
and \U$8470 ( \17291_17593 , RIe1b88f8_3477, \8957_9256 );
and \U$8471 ( \17292_17594 , RIe1b68a0_3454, \8959_9258 );
and \U$8472 ( \17293_17595 , RIfcd4db0_7444, \8961_9260 );
and \U$8473 ( \17294_17596 , RIfc4ebc0_5918, \8963_9262 );
and \U$8474 ( \17295_17597 , RIfec1e00_8326, \8965_9264 );
and \U$8475 ( \17296_17598 , RIfe8bd28_7935, \8967_9266 );
and \U$8476 ( \17297_17599 , RIf148790_5284, \8969_9268 );
and \U$8477 ( \17298_17600 , RIf1476b0_5272, \8971_9270 );
and \U$8478 ( \17299_17601 , RIfe8ba58_7933, \8973_9272 );
and \U$8479 ( \17300_17602 , RIfec1b30_8324, \8975_9274 );
and \U$8480 ( \17301_17603 , RIfc4e788_5915, \8977_9276 );
and \U$8481 ( \17302_17604 , RIfcb8e80_7126, \8979_9278 );
and \U$8482 ( \17303_17605 , RIfe8bbc0_7934, \8981_9280 );
and \U$8483 ( \17304_17606 , RIfec1c98_8325, \8983_9282 );
and \U$8484 ( \17305_17607 , RIe1a7c60_3286, \8985_9284 );
and \U$8485 ( \17306_17608 , RIe1a4f60_3254, \8987_9286 );
and \U$8486 ( \17307_17609 , RIe1a2260_3222, \8989_9288 );
and \U$8487 ( \17308_17610 , RIe19f560_3190, \8991_9290 );
and \U$8488 ( \17309_17611 , RIe18ba60_2966, \8993_9292 );
and \U$8489 ( \17310_17612 , RIe177f60_2742, \8995_9294 );
and \U$8490 ( \17311_17613 , RIe2258b8_4717, \8997_9296 );
and \U$8491 ( \17312_17614 , RIe21a4b8_4589, \8999_9298 );
and \U$8492 ( \17313_17615 , RIe203cb8_4333, \9001_9300 );
and \U$8493 ( \17314_17616 , RIe1fdd18_4265, \9003_9302 );
and \U$8494 ( \17315_17617 , RIe1f70d0_4188, \9005_9304 );
and \U$8495 ( \17316_17618 , RIe1efc18_4105, \9007_9306 );
and \U$8496 ( \17317_17619 , RIe1d4120_3790, \9009_9308 );
and \U$8497 ( \17318_17620 , RIe1bac20_3502, \9011_9310 );
and \U$8498 ( \17319_17621 , RIe1ada98_3353, \9013_9312 );
and \U$8499 ( \17320_17622 , RIe1700d0_2652, \9015_9314 );
or \U$8500 ( \17321_17623 , \17257_17559 , \17258_17560 , \17259_17561 , \17260_17562 , \17261_17563 , \17262_17564 , \17263_17565 , \17264_17566 , \17265_17567 , \17266_17568 , \17267_17569 , \17268_17570 , \17269_17571 , \17270_17572 , \17271_17573 , \17272_17574 , \17273_17575 , \17274_17576 , \17275_17577 , \17276_17578 , \17277_17579 , \17278_17580 , \17279_17581 , \17280_17582 , \17281_17583 , \17282_17584 , \17283_17585 , \17284_17586 , \17285_17587 , \17286_17588 , \17287_17589 , \17288_17590 , \17289_17591 , \17290_17592 , \17291_17593 , \17292_17594 , \17293_17595 , \17294_17596 , \17295_17597 , \17296_17598 , \17297_17599 , \17298_17600 , \17299_17601 , \17300_17602 , \17301_17603 , \17302_17604 , \17303_17605 , \17304_17606 , \17305_17607 , \17306_17608 , \17307_17609 , \17308_17610 , \17309_17611 , \17310_17612 , \17311_17613 , \17312_17614 , \17313_17615 , \17314_17616 , \17315_17617 , \17316_17618 , \17317_17619 , \17318_17620 , \17319_17621 , \17320_17622 );
or \U$8501 ( \17322_17624 , \17256_17558 , \17321_17623 );
_DC \g659c/U$1 ( \17323 , \17322_17624 , \9024_9323 );
and g659d_GF_PartitionCandidate( \17324_17626_nG659d , \17191 , \17323 );
buf \U$8502 ( \17325_17627 , \17324_17626_nG659d );
and \U$8503 ( \17326_17628 , \17325_17627 , \10389_10691 );
nor \U$8504 ( \17327_17629 , \17059_17361 , \17326_17628 );
xnor \U$8505 ( \17328_17630 , \17327_17629 , \10678_10980 );
and \U$8506 ( \17329_17631 , \11287_11586 , \15037_15336 );
and \U$8507 ( \17330_17632 , \12146_12448 , \14661_14963 );
nor \U$8508 ( \17331_17633 , \17329_17631 , \17330_17632 );
xnor \U$8509 ( \17332_17634 , \17331_17633 , \15043_15342 );
xor \U$8510 ( \17333_17635 , \17328_17630 , \17332_17634 );
and \U$8511 ( \17334_17636 , \10686_10988 , \16333_16635 );
and \U$8512 ( \17335_17637 , \10968_11270 , \15999_16301 );
nor \U$8513 ( \17336_17638 , \17334_17636 , \17335_17637 );
xnor \U$8514 ( \17337_17639 , \17336_17638 , \16323_16625 );
xor \U$8515 ( \17338_17640 , \17333_17635 , \17337_17639 );
xor \U$8516 ( \17339_17641 , \17058_17360 , \17338_17640 );
and \U$8517 ( \17340_17642 , \15022_15321 , \11275_11574 );
and \U$8518 ( \17341_17643 , \15965_16267 , \10976_11278 );
nor \U$8519 ( \17342_17644 , \17340_17642 , \17341_17643 );
xnor \U$8520 ( \17343_17645 , \17342_17644 , \11281_11580 );
and \U$8521 ( \17344_17646 , \12470_12769 , \13755_14054 );
and \U$8522 ( \17345_17647 , \13377_13679 , \13390_13692 );
nor \U$8523 ( \17346_17648 , \17344_17646 , \17345_17647 );
xnor \U$8524 ( \17347_17649 , \17346_17648 , \13736_14035 );
xor \U$8525 ( \17348_17650 , \17343_17645 , \17347_17649 );
_DC \g5146/U$1 ( \17349 , \17190_17492 , \9298_9597 );
_DC \g51ca/U$1 ( \17350 , \17322_17624 , \9024_9323 );
xor g51cb_GF_PartitionCandidate( \17351_17653_nG51cb , \17349 , \17350 );
buf \U$8526 ( \17352_17654 , \17351_17653_nG51cb );
xor \U$8527 ( \17353_17655 , \17352_17654 , \16320_16622 );
and \U$8528 ( \17354_17656 , \10385_10687 , \17353_17655 );
xor \U$8529 ( \17355_17657 , \17348_17650 , \17354_17656 );
xor \U$8530 ( \17356_17658 , \17339_17641 , \17355_17657 );
xor \U$8531 ( \17357_17659 , \17054_17356 , \17356_17658 );
xor \U$8532 ( \17358_17660 , \17038_17340 , \17357_17659 );
and \U$8533 ( \17359_17661 , \16368_16670 , \16372_16674 );
and \U$8534 ( \17360_17662 , \16373_16675 , \16376_16678 );
or \U$8535 ( \17361_17663 , \17359_17661 , \17360_17662 );
xor \U$8536 ( \17362_17664 , \17358_17660 , \17361_17663 );
buf g9bea_GF_PartitionCandidate( \17363_17665_nG9bea , \17362_17664 );
and \U$8537 ( \17364_17666 , \10402_10704 , \17363_17665_nG9bea );
or \U$8538 ( \17365_17667 , \17034_17336 , \17364_17666 );
xor \U$8539 ( \17366_17668 , \10399_10703 , \17365_17667 );
buf \U$8540 ( \17367_17669 , \17366_17668 );
buf \U$8542 ( \17368_17670 , \17367_17669 );
xor \U$8543 ( \17369_17671 , \17033_17335 , \17368_17670 );
buf \U$8544 ( \17370_17672 , \17369_17671 );
and \U$8545 ( \17371_17673 , \16037_16339 , \16043_16345 );
and \U$8546 ( \17372_17674 , \16037_16339 , \16383_16685 );
and \U$8547 ( \17373_17675 , \16043_16345 , \16383_16685 );
or \U$8548 ( \17374_17676 , \17371_17673 , \17372_17674 , \17373_17675 );
buf \U$8549 ( \17375_17677 , \17374_17676 );
xor \U$8550 ( \17376_17678 , \17370_17672 , \17375_17677 );
and \U$8551 ( \17377_17679 , \16402_16704 , \16411_16710 );
and \U$8552 ( \17378_17680 , \16402_16704 , \16418_16717 );
and \U$8553 ( \17379_17681 , \16411_16710 , \16418_16717 );
or \U$8554 ( \17380_17682 , \17377_17679 , \17378_17680 , \17379_17681 );
buf \U$8555 ( \17381_17683 , \17380_17682 );
and \U$8556 ( \17382_17684 , \12183_12157 , \13771_14070_nG9bf9 );
and \U$8557 ( \17383_17685 , \11855_12154 , \14682_14984_nG9bf6 );
or \U$8558 ( \17384_17686 , \17382_17684 , \17383_17685 );
xor \U$8559 ( \17385_17687 , \11854_12153 , \17384_17686 );
buf \U$8560 ( \17386_17688 , \17385_17687 );
buf \U$8562 ( \17387_17689 , \17386_17688 );
xor \U$8563 ( \17388_17690 , \17381_17683 , \17387_17689 );
and \U$8564 ( \17389_17691 , \10996_10421 , \15074_15373_nG9bf3 );
and \U$8565 ( \17390_17692 , \10119_10418 , \16013_16315_nG9bf0 );
or \U$8566 ( \17391_17693 , \17389_17691 , \17390_17692 );
xor \U$8567 ( \17392_17694 , \10118_10417 , \17391_17693 );
buf \U$8568 ( \17393_17695 , \17392_17694 );
buf \U$8570 ( \17394_17696 , \17393_17695 );
xor \U$8571 ( \17395_17697 , \17388_17690 , \17394_17696 );
buf \U$8572 ( \17396_17698 , \17395_17697 );
xor \U$8573 ( \17397_17699 , \17376_17678 , \17396_17698 );
buf \U$8574 ( \17398_17700 , \17397_17699 );
and \U$8575 ( \17399_17701 , \16385_16687 , \16390_16692 );
and \U$8576 ( \17400_17702 , \16385_16687 , \16431_16730 );
and \U$8577 ( \17401_17703 , \16390_16692 , \16431_16730 );
or \U$8578 ( \17402_17704 , \17399_17701 , \17400_17702 , \17401_17703 );
buf \U$8579 ( \17403_17705 , \17402_17704 );
xor \U$8580 ( \17404_17706 , \17398_17700 , \17403_17705 );
and \U$8581 ( \17405_17707 , \16433_16732 , \16438_16737 );
and \U$8582 ( \17406_17708 , \16433_16732 , \16444_16743 );
and \U$8583 ( \17407_17709 , \16438_16737 , \16444_16743 );
or \U$8584 ( \17408_17710 , \17405_17707 , \17406_17708 , \17407_17709 );
buf \U$8585 ( \17409_17711 , \17408_17710 );
xor \U$8586 ( \17410_17712 , \17404_17706 , \17409_17711 );
and \U$8587 ( \17411_17713 , \16446_16745 , \17410_17712 );
and \U$8588 ( \17412_17714 , \17001_17303 , \17410_17712 );
or \U$8589 ( \17413_17715 , \17002_17304 , \17411_17713 , \17412_17714 );
and \U$8590 ( \17414_17716 , \17007_17309 , \17032_17334 );
and \U$8591 ( \17415_17717 , \17007_17309 , \17368_17670 );
and \U$8592 ( \17416_17718 , \17032_17334 , \17368_17670 );
or \U$8593 ( \17417_17719 , \17414_17716 , \17415_17717 , \17416_17718 );
buf \U$8594 ( \17418_17720 , \17417_17719 );
and \U$8595 ( \17419_17721 , \17381_17683 , \17387_17689 );
and \U$8596 ( \17420_17722 , \17381_17683 , \17394_17696 );
and \U$8597 ( \17421_17723 , \17387_17689 , \17394_17696 );
or \U$8598 ( \17422_17724 , \17419_17721 , \17420_17722 , \17421_17723 );
buf \U$8599 ( \17423_17725 , \17422_17724 );
and \U$8600 ( \17424_17726 , \16994_17293 , \16998_17300 );
buf \U$8601 ( \17425_17727 , \17424_17726 );
buf \U$8603 ( \17426_17728 , \17425_17727 );
and \U$8604 ( \17427_17729 , \16405_15940 , \10981_11283_nG9c08 );
and \U$8605 ( \17428_17730 , \15638_15937 , \11299_11598_nG9c05 );
or \U$8606 ( \17429_17731 , \17427_17729 , \17428_17730 );
xor \U$8607 ( \17430_17732 , \15637_15936 , \17429_17731 );
buf \U$8608 ( \17431_17733 , \17430_17732 );
buf \U$8610 ( \17432_17734 , \17431_17733 );
xor \U$8611 ( \17433_17735 , \17426_17728 , \17432_17734 );
buf \U$8612 ( \17434_17736 , \17433_17735 );
not \U$8169 ( \17435_17295 , \16995_17294 );
xor \U$8170 ( \17436_17296 , \16989_17288_nG4430 , \16992_17291_nG4433 );
and \U$8171 ( \17437_17297 , \17435_17295 , \17436_17296 );
and \U$8613 ( \17438_17737 , \17437_17297 , \10392_10694_nG9c0e );
and \U$8614 ( \17439_17738 , \16995_17294 , \10693_10995_nG9c0b );
or \U$8615 ( \17440_17739 , \17438_17737 , \17439_17738 );
xor \U$8616 ( \17441_17740 , \16994_17293 , \17440_17739 );
buf \U$8617 ( \17442_17741 , \17441_17740 );
buf \U$8619 ( \17443_17742 , \17442_17741 );
xor \U$8620 ( \17444_17743 , \17434_17736 , \17443_17742 );
and \U$8621 ( \17445_17744 , \14710_14631 , \12168_12470_nG9c02 );
and \U$8622 ( \17446_17745 , \14329_14628 , \12502_12801_nG9bff );
or \U$8623 ( \17447_17746 , \17445_17744 , \17446_17745 );
xor \U$8624 ( \17448_17747 , \14328_14627 , \17447_17746 );
buf \U$8625 ( \17449_17748 , \17448_17747 );
buf \U$8627 ( \17450_17749 , \17449_17748 );
xor \U$8628 ( \17451_17750 , \17444_17743 , \17450_17749 );
buf \U$8629 ( \17452_17751 , \17451_17750 );
and \U$8630 ( \17453_17752 , \17013_17315 , \17019_17321 );
buf \U$8631 ( \17454_17753 , \17453_17752 );
xor \U$8632 ( \17455_17754 , \17452_17751 , \17454_17753 );
and \U$8633 ( \17456_17755 , \13431_13370 , \13403_13705_nG9bfc );
and \U$8634 ( \17457_17756 , \13068_13367 , \13771_14070_nG9bf9 );
or \U$8635 ( \17458_17757 , \17456_17755 , \17457_17756 );
xor \U$8636 ( \17459_17758 , \13067_13366 , \17458_17757 );
buf \U$8637 ( \17460_17759 , \17459_17758 );
buf \U$8639 ( \17461_17760 , \17460_17759 );
xor \U$8640 ( \17462_17761 , \17455_17754 , \17461_17760 );
buf \U$8641 ( \17463_17762 , \17462_17761 );
xor \U$8642 ( \17464_17763 , \17423_17725 , \17463_17762 );
and \U$8643 ( \17465_17764 , \10411_10707 , \17363_17665_nG9bea );
and \U$8644 ( \17466_17765 , \17058_17360 , \17338_17640 );
and \U$8645 ( \17467_17766 , \17338_17640 , \17355_17657 );
and \U$8646 ( \17468_17767 , \17058_17360 , \17355_17657 );
or \U$8647 ( \17469_17768 , \17466_17765 , \17467_17766 , \17468_17767 );
and \U$8648 ( \17470_17769 , \17325_17627 , \10681_10983 );
and \U$8649 ( \17471_17770 , RIdec4730_699, \9034_9333 );
and \U$8650 ( \17472_17771 , RIdec1a30_667, \9036_9335 );
and \U$8651 ( \17473_17772 , RIfce3f90_7616, \9038_9337 );
and \U$8652 ( \17474_17773 , RIdebed30_635, \9040_9339 );
and \U$8653 ( \17475_17774 , RIfcc3308_7243, \9042_9341 );
and \U$8654 ( \17476_17775 , RIdebc030_603, \9044_9343 );
and \U$8655 ( \17477_17776 , RIdeb9330_571, \9046_9345 );
and \U$8656 ( \17478_17777 , RIdeb6630_539, \9048_9347 );
and \U$8657 ( \17479_17778 , RIfc8c588_6619, \9050_9349 );
and \U$8658 ( \17480_17779 , RIdeb0c30_475, \9052_9351 );
and \U$8659 ( \17481_17780 , RIfc5a998_6053, \9054_9353 );
and \U$8660 ( \17482_17781 , RIdeadf30_443, \9056_9355 );
and \U$8661 ( \17483_17782 , RIfc99b48_6771, \9058_9357 );
and \U$8662 ( \17484_17783 , RIdea8698_411, \9060_9359 );
and \U$8663 ( \17485_17784 , RIdea1d98_379, \9062_9361 );
and \U$8664 ( \17486_17785 , RIde9b498_347, \9064_9363 );
and \U$8665 ( \17487_17786 , RIfc78bf0_6396, \9066_9365 );
and \U$8666 ( \17488_17787 , RIfcbc558_7165, \9068_9367 );
and \U$8667 ( \17489_17788 , RIfca12d0_6856, \9070_9369 );
and \U$8668 ( \17490_17789 , RIfca3fd0_6888, \9072_9371 );
and \U$8669 ( \17491_17790 , RIfec2670_8332, \9074_9373 );
and \U$8670 ( \17492_17791 , RIfec2508_8331, \9076_9375 );
and \U$8671 ( \17493_17792 , RIde88a00_256, \9078_9377 );
and \U$8672 ( \17494_17793 , RIde84518_235, \9080_9379 );
and \U$8673 ( \17495_17794 , RIfcc35d8_7245, \9082_9381 );
and \U$8674 ( \17496_17795 , RIfcb57a8_7087, \9084_9383 );
and \U$8675 ( \17497_17796 , RIfc5a290_6048, \9086_9385 );
and \U$8676 ( \17498_17797 , RIfca3058_6877, \9088_9387 );
and \U$8677 ( \17499_17798 , RIee38e78_5106, \9090_9389 );
and \U$8678 ( \17500_17799 , RIfec27d8_8333, \9092_9391 );
and \U$8679 ( \17501_17800 , RIfca3328_6879, \9094_9393 );
and \U$8680 ( \17502_17801 , RIe1672c8_2551, \9096_9395 );
and \U$8681 ( \17503_17802 , RIe164730_2520, \9098_9397 );
and \U$8682 ( \17504_17803 , RIe161a30_2488, \9100_9399 );
and \U$8683 ( \17505_17804 , RIee36cb8_5082, \9102_9401 );
and \U$8684 ( \17506_17805 , RIe15ed30_2456, \9104_9403 );
and \U$8685 ( \17507_17806 , RIfcc7250_7288, \9106_9405 );
and \U$8686 ( \17508_17807 , RIe15c030_2424, \9108_9407 );
and \U$8687 ( \17509_17808 , RIe156630_2360, \9110_9409 );
and \U$8688 ( \17510_17809 , RIe153930_2328, \9112_9411 );
and \U$8689 ( \17511_17810 , RIfcc7688_7291, \9114_9413 );
and \U$8690 ( \17512_17811 , RIe150c30_2296, \9116_9415 );
and \U$8691 ( \17513_17812 , RIfc8af08_6603, \9118_9417 );
and \U$8692 ( \17514_17813 , RIe14df30_2264, \9120_9419 );
and \U$8693 ( \17515_17814 , RIfc9a250_6776, \9122_9421 );
and \U$8694 ( \17516_17815 , RIe14b230_2232, \9124_9423 );
and \U$8695 ( \17517_17816 , RIe148530_2200, \9126_9425 );
and \U$8696 ( \17518_17817 , RIe145830_2168, \9128_9427 );
and \U$8697 ( \17519_17818 , RIfc9aac0_6782, \9130_9429 );
and \U$8698 ( \17520_17819 , RIfc56bb8_6009, \9132_9431 );
and \U$8699 ( \17521_17820 , RIfca1ca8_6863, \9134_9433 );
and \U$8700 ( \17522_17821 , RIfcec960_7714, \9136_9435 );
and \U$8701 ( \17523_17822 , RIe1406a0_2110, \9138_9437 );
and \U$8702 ( \17524_17823 , RIdf3e440_2085, \9140_9439 );
and \U$8703 ( \17525_17824 , RIdf3c280_2061, \9142_9441 );
and \U$8704 ( \17526_17825 , RIdf39f58_2036, \9144_9443 );
and \U$8705 ( \17527_17826 , RIfc9a958_6781, \9146_9445 );
and \U$8706 ( \17528_17827 , RIee2f0f8_4994, \9148_9447 );
and \U$8707 ( \17529_17828 , RIfcdb458_7517, \9150_9449 );
and \U$8708 ( \17530_17829 , RIee2cf38_4970, \9152_9451 );
and \U$8709 ( \17531_17830 , RIdf34c60_1977, \9154_9453 );
and \U$8710 ( \17532_17831 , RIfec2940_8334, \9156_9455 );
and \U$8711 ( \17533_17832 , RIdf30778_1928, \9158_9457 );
and \U$8712 ( \17534_17833 , RIdf2e888_1906, \9160_9459 );
or \U$8713 ( \17535_17834 , \17471_17770 , \17472_17771 , \17473_17772 , \17474_17773 , \17475_17774 , \17476_17775 , \17477_17776 , \17478_17777 , \17479_17778 , \17480_17779 , \17481_17780 , \17482_17781 , \17483_17782 , \17484_17783 , \17485_17784 , \17486_17785 , \17487_17786 , \17488_17787 , \17489_17788 , \17490_17789 , \17491_17790 , \17492_17791 , \17493_17792 , \17494_17793 , \17495_17794 , \17496_17795 , \17497_17796 , \17498_17797 , \17499_17798 , \17500_17799 , \17501_17800 , \17502_17801 , \17503_17802 , \17504_17803 , \17505_17804 , \17506_17805 , \17507_17806 , \17508_17807 , \17509_17808 , \17510_17809 , \17511_17810 , \17512_17811 , \17513_17812 , \17514_17813 , \17515_17814 , \17516_17815 , \17517_17816 , \17518_17817 , \17519_17818 , \17520_17819 , \17521_17820 , \17522_17821 , \17523_17822 , \17524_17823 , \17525_17824 , \17526_17825 , \17527_17826 , \17528_17827 , \17529_17828 , \17530_17829 , \17531_17830 , \17532_17831 , \17533_17832 , \17534_17833 );
and \U$8714 ( \17536_17835 , RIee2b480_4951, \9163_9462 );
and \U$8715 ( \17537_17836 , RIfec23a0_8330, \9165_9464 );
and \U$8716 ( \17538_17837 , RIee288e8_4920, \9167_9466 );
and \U$8717 ( \17539_17838 , RIfec2238_8329, \9169_9468 );
and \U$8718 ( \17540_17839 , RIdf29b30_1851, \9171_9470 );
and \U$8719 ( \17541_17840 , RIdf27808_1826, \9173_9472 );
and \U$8720 ( \17542_17841 , RIdf25a80_1805, \9175_9474 );
and \U$8721 ( \17543_17842 , RIdf23e60_1785, \9177_9476 );
and \U$8722 ( \17544_17843 , RIfc55100_5990, \9179_9478 );
and \U$8723 ( \17545_17844 , RIfcd9f40_7502, \9181_9480 );
and \U$8724 ( \17546_17845 , RIfc54f98_5989, \9183_9482 );
and \U$8725 ( \17547_17846 , RIfc54cc8_5987, \9185_9484 );
and \U$8726 ( \17548_17847 , RIfc4b218_5877, \9187_9486 );
and \U$8727 ( \17549_17848 , RIdf1efa0_1729, \9189_9488 );
and \U$8728 ( \17550_17849 , RIfcc69e0_7282, \9191_9490 );
and \U$8729 ( \17551_17850 , RIdf18bc8_1658, \9193_9492 );
and \U$8730 ( \17552_17851 , RIdf16300_1629, \9195_9494 );
and \U$8731 ( \17553_17852 , RIdf13600_1597, \9197_9496 );
and \U$8732 ( \17554_17853 , RIdf10900_1565, \9199_9498 );
and \U$8733 ( \17555_17854 , RIdf0dc00_1533, \9201_9500 );
and \U$8734 ( \17556_17855 , RIdf0af00_1501, \9203_9502 );
and \U$8735 ( \17557_17856 , RIdf08200_1469, \9205_9504 );
and \U$8736 ( \17558_17857 , RIdf05500_1437, \9207_9506 );
and \U$8737 ( \17559_17858 , RIdf02800_1405, \9209_9508 );
and \U$8738 ( \17560_17859 , RIdefce00_1341, \9211_9510 );
and \U$8739 ( \17561_17860 , RIdefa100_1309, \9213_9512 );
and \U$8740 ( \17562_17861 , RIdef7400_1277, \9215_9514 );
and \U$8741 ( \17563_17862 , RIdef4700_1245, \9217_9516 );
and \U$8742 ( \17564_17863 , RIdef1a00_1213, \9219_9518 );
and \U$8743 ( \17565_17864 , RIdeeed00_1181, \9221_9520 );
and \U$8744 ( \17566_17865 , RIdeec000_1149, \9223_9522 );
and \U$8745 ( \17567_17866 , RIdee9300_1117, \9225_9524 );
and \U$8746 ( \17568_17867 , RIfce4ad0_7624, \9227_9526 );
and \U$8747 ( \17569_17868 , RIfc9e8a0_6826, \9229_9528 );
and \U$8748 ( \17570_17869 , RIfcc46b8_7257, \9231_9530 );
and \U$8749 ( \17571_17870 , RIfcd4108_7435, \9233_9532 );
and \U$8750 ( \17572_17871 , RIdee4440_1061, \9235_9534 );
and \U$8751 ( \17573_17872 , RIdee2280_1037, \9237_9536 );
and \U$8752 ( \17574_17873 , RIdee0390_1015, \9239_9538 );
and \U$8753 ( \17575_17874 , RIdede068_990, \9241_9540 );
and \U$8754 ( \17576_17875 , RIfcda0a8_7503, \9243_9542 );
and \U$8755 ( \17577_17876 , RIfce54a8_7631, \9245_9544 );
and \U$8756 ( \17578_17877 , RIfca0790_6848, \9247_9546 );
and \U$8757 ( \17579_17878 , RIfc50ee8_5943, \9249_9548 );
and \U$8758 ( \17580_17879 , RIded8d70_931, \9251_9550 );
and \U$8759 ( \17581_17880 , RIded68e0_905, \9253_9552 );
and \U$8760 ( \17582_17881 , RIded4888_882, \9255_9554 );
and \U$8761 ( \17583_17882 , RIded2560_857, \9257_9556 );
and \U$8762 ( \17584_17883 , RIdecfb30_827, \9259_9558 );
and \U$8763 ( \17585_17884 , RIdecce30_795, \9261_9560 );
and \U$8764 ( \17586_17885 , RIdeca130_763, \9263_9562 );
and \U$8765 ( \17587_17886 , RIdec7430_731, \9265_9564 );
and \U$8766 ( \17588_17887 , RIdeb3930_507, \9267_9566 );
and \U$8767 ( \17589_17888 , RIde94b98_315, \9269_9568 );
and \U$8768 ( \17590_17889 , RIe16d538_2621, \9271_9570 );
and \U$8769 ( \17591_17890 , RIe159330_2392, \9273_9572 );
and \U$8770 ( \17592_17891 , RIe142b30_2136, \9275_9574 );
and \U$8771 ( \17593_17892 , RIdf37528_2006, \9277_9576 );
and \U$8772 ( \17594_17893 , RIdf2bb88_1874, \9279_9578 );
and \U$8773 ( \17595_17894 , RIdf1c408_1698, \9281_9580 );
and \U$8774 ( \17596_17895 , RIdeffb00_1373, \9283_9582 );
and \U$8775 ( \17597_17896 , RIdee6600_1085, \9285_9584 );
and \U$8776 ( \17598_17897 , RIdedb368_958, \9287_9586 );
and \U$8777 ( \17599_17898 , RIde7aae0_188, \9289_9588 );
or \U$8778 ( \17600_17899 , \17536_17835 , \17537_17836 , \17538_17837 , \17539_17838 , \17540_17839 , \17541_17840 , \17542_17841 , \17543_17842 , \17544_17843 , \17545_17844 , \17546_17845 , \17547_17846 , \17548_17847 , \17549_17848 , \17550_17849 , \17551_17850 , \17552_17851 , \17553_17852 , \17554_17853 , \17555_17854 , \17556_17855 , \17557_17856 , \17558_17857 , \17559_17858 , \17560_17859 , \17561_17860 , \17562_17861 , \17563_17862 , \17564_17863 , \17565_17864 , \17566_17865 , \17567_17866 , \17568_17867 , \17569_17868 , \17570_17869 , \17571_17870 , \17572_17871 , \17573_17872 , \17574_17873 , \17575_17874 , \17576_17875 , \17577_17876 , \17578_17877 , \17579_17878 , \17580_17879 , \17581_17880 , \17582_17881 , \17583_17882 , \17584_17883 , \17585_17884 , \17586_17885 , \17587_17886 , \17588_17887 , \17589_17888 , \17590_17889 , \17591_17890 , \17592_17891 , \17593_17892 , \17594_17893 , \17595_17894 , \17596_17895 , \17597_17896 , \17598_17897 , \17599_17898 );
or \U$8779 ( \17601_17900 , \17535_17834 , \17600_17899 );
_DC \g659e/U$1 ( \17602 , \17601_17900 , \9298_9597 );
and \U$8780 ( \17603_17902 , RIe19c9c8_3159, \8760_9059 );
and \U$8781 ( \17604_17903 , RIe199cc8_3127, \8762_9061 );
and \U$8782 ( \17605_17904 , RIfe8ea28_7967, \8764_9063 );
and \U$8783 ( \17606_17905 , RIe196fc8_3095, \8766_9065 );
and \U$8784 ( \17607_17906 , RIfec20d0_8328, \8768_9067 );
and \U$8785 ( \17608_17907 , RIe1942c8_3063, \8770_9069 );
and \U$8786 ( \17609_17908 , RIe1915c8_3031, \8772_9071 );
and \U$8787 ( \17610_17909 , RIe18e8c8_2999, \8774_9073 );
and \U$8788 ( \17611_17910 , RIe188ec8_2935, \8776_9075 );
and \U$8789 ( \17612_17911 , RIe1861c8_2903, \8778_9077 );
and \U$8790 ( \17613_17912 , RIfc68228_6207, \8780_9079 );
and \U$8791 ( \17614_17913 , RIe1834c8_2871, \8782_9081 );
and \U$8792 ( \17615_17914 , RIfccb5d0_7336, \8784_9083 );
and \U$8793 ( \17616_17915 , RIe1807c8_2839, \8786_9085 );
and \U$8794 ( \17617_17916 , RIe17dac8_2807, \8788_9087 );
and \U$8795 ( \17618_17917 , RIe17adc8_2775, \8790_9089 );
and \U$8796 ( \17619_17918 , RIf141e18_5209, \8792_9091 );
and \U$8797 ( \17620_17919 , RIf140900_5194, \8794_9093 );
and \U$8798 ( \17621_17920 , RIf140090_5188, \8796_9095 );
and \U$8799 ( \17622_17921 , RIe1753c8_2711, \8798_9097 );
and \U$8800 ( \17623_17922 , RIf13f988_5183, \8800_9099 );
and \U$8801 ( \17624_17923 , RIf13ece0_5174, \8802_9101 );
and \U$8802 ( \17625_17924 , RIee3e170_5165, \8804_9103 );
and \U$8803 ( \17626_17925 , RIee3cf28_5152, \8806_9105 );
and \U$8804 ( \17627_17926 , RIee3bce0_5139, \8808_9107 );
and \U$8805 ( \17628_17927 , RIee3ac00_5127, \8810_9109 );
and \U$8806 ( \17629_17928 , RIee39850_5113, \8812_9111 );
and \U$8807 ( \17630_17929 , RIe172dd0_2684, \8814_9113 );
and \U$8808 ( \17631_17930 , RIf16fc28_5731, \8816_9115 );
and \U$8809 ( \17632_17931 , RIf16f0e8_5723, \8818_9117 );
and \U$8810 ( \17633_17932 , RIf16dd38_5709, \8820_9119 );
and \U$8811 ( \17634_17933 , RIfce9120_7674, \8822_9121 );
and \U$8812 ( \17635_17934 , RIfc404a8_5757, \8824_9123 );
and \U$8813 ( \17636_17935 , RIe222d20_4686, \8826_9125 );
and \U$8814 ( \17637_17936 , RIf16b8a8_5683, \8828_9127 );
and \U$8815 ( \17638_17937 , RIe220020_4654, \8830_9129 );
and \U$8816 ( \17639_17938 , RIf16a930_5672, \8832_9131 );
and \U$8817 ( \17640_17939 , RIe21d320_4622, \8834_9133 );
and \U$8818 ( \17641_17940 , RIe217920_4558, \8836_9135 );
and \U$8819 ( \17642_17941 , RIe214c20_4526, \8838_9137 );
and \U$8820 ( \17643_17942 , RIfc5b910_6064, \8840_9139 );
and \U$8821 ( \17644_17943 , RIe211f20_4494, \8842_9141 );
and \U$8822 ( \17645_17944 , RIfe8e8c0_7966, \8844_9143 );
and \U$8823 ( \17646_17945 , RIe20f220_4462, \8846_9145 );
and \U$8824 ( \17647_17946 , RIfe8e758_7965, \8848_9147 );
and \U$8825 ( \17648_17947 , RIe20c520_4430, \8850_9149 );
and \U$8826 ( \17649_17948 , RIe209820_4398, \8852_9151 );
and \U$8827 ( \17650_17949 , RIe206b20_4366, \8854_9153 );
and \U$8828 ( \17651_17950 , RIf166b50_5628, \8856_9155 );
and \U$8829 ( \17652_17951 , RIf165a70_5616, \8858_9157 );
and \U$8830 ( \17653_17952 , RIfe8dd80_7958, \8860_9159 );
and \U$8831 ( \17654_17953 , RIfe8dab0_7956, \8862_9161 );
and \U$8832 ( \17655_17954 , RIf164c60_5606, \8864_9163 );
and \U$8833 ( \17656_17955 , RIf163e50_5596, \8866_9165 );
and \U$8834 ( \17657_17956 , RIf162ed8_5585, \8868_9167 );
and \U$8835 ( \17658_17957 , RIf1616f0_5568, \8870_9169 );
and \U$8836 ( \17659_17958 , RIf15f800_5546, \8872_9171 );
and \U$8837 ( \17660_17959 , RIf15da78_5525, \8874_9173 );
and \U$8838 ( \17661_17960 , RIfe8d948_7955, \8876_9175 );
and \U$8839 ( \17662_17961 , RIfe8dc18_7957, \8878_9177 );
and \U$8840 ( \17663_17962 , RIf15c560_5510, \8880_9179 );
and \U$8841 ( \17664_17963 , RIf15b048_5495, \8882_9181 );
and \U$8842 ( \17665_17964 , RIfc62828_6143, \8884_9183 );
and \U$8843 ( \17666_17965 , RIf159860_5478, \8886_9185 );
or \U$8844 ( \17667_17966 , \17603_17902 , \17604_17903 , \17605_17904 , \17606_17905 , \17607_17906 , \17608_17907 , \17609_17908 , \17610_17909 , \17611_17910 , \17612_17911 , \17613_17912 , \17614_17913 , \17615_17914 , \17616_17915 , \17617_17916 , \17618_17917 , \17619_17918 , \17620_17919 , \17621_17920 , \17622_17921 , \17623_17922 , \17624_17923 , \17625_17924 , \17626_17925 , \17627_17926 , \17628_17927 , \17629_17928 , \17630_17929 , \17631_17930 , \17632_17931 , \17633_17932 , \17634_17933 , \17635_17934 , \17636_17935 , \17637_17936 , \17638_17937 , \17639_17938 , \17640_17939 , \17641_17940 , \17642_17941 , \17643_17942 , \17644_17943 , \17645_17944 , \17646_17945 , \17647_17946 , \17648_17947 , \17649_17948 , \17650_17949 , \17651_17950 , \17652_17951 , \17653_17952 , \17654_17953 , \17655_17954 , \17656_17955 , \17657_17956 , \17658_17957 , \17659_17958 , \17660_17959 , \17661_17960 , \17662_17961 , \17663_17962 , \17664_17963 , \17665_17964 , \17666_17965 );
and \U$8845 ( \17668_17967 , RIf158780_5466, \8889_9188 );
and \U$8846 ( \17669_17968 , RIf157538_5453, \8891_9190 );
and \U$8847 ( \17670_17969 , RIfca6e38_6921, \8893_9192 );
and \U$8848 ( \17671_17970 , RIe1f9b00_4218, \8895_9194 );
and \U$8849 ( \17672_17971 , RIfc61e50_6136, \8897_9196 );
and \U$8850 ( \17673_17972 , RIfc61748_6131, \8899_9198 );
and \U$8851 ( \17674_17973 , RIf154130_5416, \8901_9200 );
and \U$8852 ( \17675_17974 , RIe1f4ad8_4161, \8903_9202 );
and \U$8853 ( \17676_17975 , RIf152ab0_5400, \8905_9204 );
and \U$8854 ( \17677_17976 , RIf151700_5386, \8907_9206 );
and \U$8855 ( \17678_17977 , RIf1501e8_5371, \8909_9208 );
and \U$8856 ( \17679_17978 , RIe1f27b0_4136, \8911_9210 );
and \U$8857 ( \17680_17979 , RIfc60ed8_6125, \8913_9212 );
and \U$8858 ( \17681_17980 , RIfc7b620_6426, \8915_9214 );
and \U$8859 ( \17682_17981 , RIf14d7b8_5341, \8917_9216 );
and \U$8860 ( \17683_17982 , RIe1ed4b8_4077, \8919_9218 );
and \U$8861 ( \17684_17983 , RIe1eaa88_4047, \8921_9220 );
and \U$8862 ( \17685_17984 , RIe1e7d88_4015, \8923_9222 );
and \U$8863 ( \17686_17985 , RIe1e5088_3983, \8925_9224 );
and \U$8864 ( \17687_17986 , RIe1e2388_3951, \8927_9226 );
and \U$8865 ( \17688_17987 , RIe1df688_3919, \8929_9228 );
and \U$8866 ( \17689_17988 , RIe1dc988_3887, \8931_9230 );
and \U$8867 ( \17690_17989 , RIe1d9c88_3855, \8933_9232 );
and \U$8868 ( \17691_17990 , RIe1d6f88_3823, \8935_9234 );
and \U$8869 ( \17692_17991 , RIe1d1588_3759, \8937_9236 );
and \U$8870 ( \17693_17992 , RIe1ce888_3727, \8939_9238 );
and \U$8871 ( \17694_17993 , RIe1cbb88_3695, \8941_9240 );
and \U$8872 ( \17695_17994 , RIe1c8e88_3663, \8943_9242 );
and \U$8873 ( \17696_17995 , RIe1c6188_3631, \8945_9244 );
and \U$8874 ( \17697_17996 , RIe1c3488_3599, \8947_9246 );
and \U$8875 ( \17698_17997 , RIe1c0788_3567, \8949_9248 );
and \U$8876 ( \17699_17998 , RIe1bda88_3535, \8951_9250 );
and \U$8877 ( \17700_17999 , RIfca4de0_6898, \8953_9252 );
and \U$8878 ( \17701_18000 , RIfc5ea48_6099, \8955_9254 );
and \U$8879 ( \17702_18001 , RIe1b8a60_3478, \8957_9256 );
and \U$8880 ( \17703_18002 , RIe1b6a08_3455, \8959_9258 );
and \U$8881 ( \17704_18003 , RIfcbd638_7177, \8961_9260 );
and \U$8882 ( \17705_18004 , RIfc44fa8_5807, \8963_9262 );
and \U$8883 ( \17706_18005 , RIfe8e5f0_7964, \8965_9264 );
and \U$8884 ( \17707_18006 , RIfe8e1b8_7961, \8967_9266 );
and \U$8885 ( \17708_18007 , RIf1488f8_5285, \8969_9268 );
and \U$8886 ( \17709_18008 , RIf147818_5273, \8971_9270 );
and \U$8887 ( \17710_18009 , RIfe8e050_7960, \8973_9272 );
and \U$8888 ( \17711_18010 , RIfe8e488_7963, \8975_9274 );
and \U$8889 ( \17712_18011 , RIf146e40_5266, \8977_9276 );
and \U$8890 ( \17713_18012 , RIf146030_5256, \8979_9278 );
and \U$8891 ( \17714_18013 , RIfe8dee8_7959, \8981_9280 );
and \U$8892 ( \17715_18014 , RIfe8e320_7962, \8983_9282 );
and \U$8893 ( \17716_18015 , RIe1a7dc8_3287, \8985_9284 );
and \U$8894 ( \17717_18016 , RIe1a50c8_3255, \8987_9286 );
and \U$8895 ( \17718_18017 , RIe1a23c8_3223, \8989_9288 );
and \U$8896 ( \17719_18018 , RIe19f6c8_3191, \8991_9290 );
and \U$8897 ( \17720_18019 , RIe18bbc8_2967, \8993_9292 );
and \U$8898 ( \17721_18020 , RIe1780c8_2743, \8995_9294 );
and \U$8899 ( \17722_18021 , RIe225a20_4718, \8997_9296 );
and \U$8900 ( \17723_18022 , RIe21a620_4590, \8999_9298 );
and \U$8901 ( \17724_18023 , RIe203e20_4334, \9001_9300 );
and \U$8902 ( \17725_18024 , RIe1fde80_4266, \9003_9302 );
and \U$8903 ( \17726_18025 , RIe1f7238_4189, \9005_9304 );
and \U$8904 ( \17727_18026 , RIe1efd80_4106, \9007_9306 );
and \U$8905 ( \17728_18027 , RIe1d4288_3791, \9009_9308 );
and \U$8906 ( \17729_18028 , RIe1bad88_3503, \9011_9310 );
and \U$8907 ( \17730_18029 , RIe1adc00_3354, \9013_9312 );
and \U$8908 ( \17731_18030 , RIe170238_2653, \9015_9314 );
or \U$8909 ( \17732_18031 , \17668_17967 , \17669_17968 , \17670_17969 , \17671_17970 , \17672_17971 , \17673_17972 , \17674_17973 , \17675_17974 , \17676_17975 , \17677_17976 , \17678_17977 , \17679_17978 , \17680_17979 , \17681_17980 , \17682_17981 , \17683_17982 , \17684_17983 , \17685_17984 , \17686_17985 , \17687_17986 , \17688_17987 , \17689_17988 , \17690_17989 , \17691_17990 , \17692_17991 , \17693_17992 , \17694_17993 , \17695_17994 , \17696_17995 , \17697_17996 , \17698_17997 , \17699_17998 , \17700_17999 , \17701_18000 , \17702_18001 , \17703_18002 , \17704_18003 , \17705_18004 , \17706_18005 , \17707_18006 , \17708_18007 , \17709_18008 , \17710_18009 , \17711_18010 , \17712_18011 , \17713_18012 , \17714_18013 , \17715_18014 , \17716_18015 , \17717_18016 , \17718_18017 , \17719_18018 , \17720_18019 , \17721_18020 , \17722_18021 , \17723_18022 , \17724_18023 , \17725_18024 , \17726_18025 , \17727_18026 , \17728_18027 , \17729_18028 , \17730_18029 , \17731_18030 );
or \U$8910 ( \17733_18032 , \17667_17966 , \17732_18031 );
_DC \g659f/U$1 ( \17734 , \17733_18032 , \9024_9323 );
and g65a0_GF_PartitionCandidate( \17735_18034_nG65a0 , \17602 , \17734 );
buf \U$8911 ( \17736_18035 , \17735_18034_nG65a0 );
and \U$8912 ( \17737_18036 , \17736_18035 , \10389_10691 );
nor \U$8913 ( \17738_18037 , \17470_17769 , \17737_18036 );
xnor \U$8914 ( \17739_18038 , \17738_18037 , \10678_10980 );
not \U$8915 ( \17740_18039 , \17354_17656 );
_DC \g524f/U$1 ( \17741 , \17601_17900 , \9298_9597 );
_DC \g52d3/U$1 ( \17742 , \17733_18032 , \9024_9323 );
xor g52d4_GF_PartitionCandidate( \17743_18042_nG52d4 , \17741 , \17742 );
buf \U$8916 ( \17744_18043 , \17743_18042_nG52d4 );
and \U$8917 ( \17745_18044 , \17352_17654 , \16320_16622 );
not \U$8918 ( \17746_18045 , \17745_18044 );
and \U$8919 ( \17747_18046 , \17744_18043 , \17746_18045 );
and \U$8920 ( \17748_18047 , \17740_18039 , \17747_18046 );
xor \U$8921 ( \17749_18048 , \17739_18038 , \17748_18047 );
and \U$8922 ( \17750_18049 , \17328_17630 , \17332_17634 );
and \U$8923 ( \17751_18050 , \17332_17634 , \17337_17639 );
and \U$8924 ( \17752_18051 , \17328_17630 , \17337_17639 );
or \U$8925 ( \17753_18052 , \17750_18049 , \17751_18050 , \17752_18051 );
xor \U$8926 ( \17754_18053 , \17749_18048 , \17753_18052 );
and \U$8927 ( \17755_18054 , \17343_17645 , \17347_17649 );
and \U$8928 ( \17756_18055 , \17347_17649 , \17354_17656 );
and \U$8929 ( \17757_18056 , \17343_17645 , \17354_17656 );
or \U$8930 ( \17758_18057 , \17755_18054 , \17756_18055 , \17757_18056 );
xor \U$8931 ( \17759_18058 , \17754_18053 , \17758_18057 );
xor \U$8932 ( \17760_18059 , \17469_17768 , \17759_18058 );
and \U$8933 ( \17761_18060 , \17046_17348 , \17047_17349 );
and \U$8934 ( \17762_18061 , \17047_17349 , \17052_17354 );
and \U$8935 ( \17763_18062 , \17046_17348 , \17052_17354 );
or \U$8936 ( \17764_18063 , \17761_18060 , \17762_18061 , \17763_18062 );
and \U$8937 ( \17765_18064 , \15965_16267 , \11275_11574 );
and \U$8938 ( \17766_18065 , \16353_16655 , \10976_11278 );
nor \U$8939 ( \17767_18066 , \17765_18064 , \17766_18065 );
xnor \U$8940 ( \17768_18067 , \17767_18066 , \11281_11580 );
and \U$8941 ( \17769_18068 , \13377_13679 , \13755_14054 );
and \U$8942 ( \17770_18069 , \13725_14024 , \13390_13692 );
nor \U$8943 ( \17771_18070 , \17769_18068 , \17770_18069 );
xnor \U$8944 ( \17772_18071 , \17771_18070 , \13736_14035 );
xor \U$8945 ( \17773_18072 , \17768_18067 , \17772_18071 );
and \U$8946 ( \17774_18073 , \12146_12448 , \15037_15336 );
and \U$8947 ( \17775_18074 , \12470_12769 , \14661_14963 );
nor \U$8948 ( \17776_18075 , \17774_18073 , \17775_18074 );
xnor \U$8949 ( \17777_18076 , \17776_18075 , \15043_15342 );
xor \U$8950 ( \17778_18077 , \17773_18072 , \17777_18076 );
xor \U$8951 ( \17779_18078 , \17764_18063 , \17778_18077 );
and \U$8952 ( \17780_18079 , \14648_14950 , \12491_12790 );
and \U$8953 ( \17781_18080 , \15022_15321 , \12159_12461 );
nor \U$8954 ( \17782_18081 , \17780_18079 , \17781_18080 );
xnor \U$8955 ( \17783_18082 , \17782_18081 , \12481_12780 );
and \U$8956 ( \17784_18083 , \10968_11270 , \16333_16635 );
and \U$8957 ( \17785_18084 , \11287_11586 , \15999_16301 );
nor \U$8958 ( \17786_18085 , \17784_18083 , \17785_18084 );
xnor \U$8959 ( \17787_18086 , \17786_18085 , \16323_16625 );
xor \U$8960 ( \17788_18087 , \17783_18082 , \17787_18086 );
xor \U$8961 ( \17789_18088 , \17744_18043 , \17352_17654 );
not \U$8962 ( \17790_18089 , \17353_17655 );
and \U$8963 ( \17791_18090 , \17789_18088 , \17790_18089 );
and \U$8964 ( \17792_18091 , \10385_10687 , \17791_18090 );
and \U$8965 ( \17793_18092 , \10686_10988 , \17353_17655 );
nor \U$8966 ( \17794_18093 , \17792_18091 , \17793_18092 );
xnor \U$8967 ( \17795_18094 , \17794_18093 , \17747_18046 );
xor \U$8968 ( \17796_18095 , \17788_18087 , \17795_18094 );
xor \U$8969 ( \17797_18096 , \17779_18078 , \17796_18095 );
xor \U$8970 ( \17798_18097 , \17760_18059 , \17797_18096 );
and \U$8971 ( \17799_18098 , \17042_17344 , \17053_17355 );
and \U$8972 ( \17800_18099 , \17053_17355 , \17356_17658 );
and \U$8973 ( \17801_18100 , \17042_17344 , \17356_17658 );
or \U$8974 ( \17802_18101 , \17799_18098 , \17800_18099 , \17801_18100 );
xor \U$8975 ( \17803_18102 , \17798_18097 , \17802_18101 );
and \U$8976 ( \17804_18103 , \17038_17340 , \17357_17659 );
and \U$8977 ( \17805_18104 , \17358_17660 , \17361_17663 );
or \U$8978 ( \17806_18105 , \17804_18103 , \17805_18104 );
xor \U$8979 ( \17807_18106 , \17803_18102 , \17806_18105 );
buf g9be7_GF_PartitionCandidate( \17808_18107_nG9be7 , \17807_18106 );
and \U$8980 ( \17809_18108 , \10402_10704 , \17808_18107_nG9be7 );
or \U$8981 ( \17810_18109 , \17465_17764 , \17809_18108 );
xor \U$8982 ( \17811_18110 , \10399_10703 , \17810_18109 );
buf \U$8983 ( \17812_18111 , \17811_18110 );
buf \U$8985 ( \17813_18112 , \17812_18111 );
xor \U$8986 ( \17814_18113 , \17464_17763 , \17813_18112 );
buf \U$8987 ( \17815_18114 , \17814_18113 );
xor \U$8988 ( \17816_18115 , \17418_17720 , \17815_18114 );
and \U$8989 ( \17817_18116 , \17021_17323 , \17023_17325 );
and \U$8990 ( \17818_18117 , \17021_17323 , \17030_17332 );
and \U$8991 ( \17819_18118 , \17023_17325 , \17030_17332 );
or \U$8992 ( \17820_18119 , \17817_18116 , \17818_18117 , \17819_18118 );
buf \U$8993 ( \17821_18120 , \17820_18119 );
and \U$8994 ( \17822_18121 , \12183_12157 , \14682_14984_nG9bf6 );
and \U$8995 ( \17823_18122 , \11855_12154 , \15074_15373_nG9bf3 );
or \U$8996 ( \17824_18123 , \17822_18121 , \17823_18122 );
xor \U$8997 ( \17825_18124 , \11854_12153 , \17824_18123 );
buf \U$8998 ( \17826_18125 , \17825_18124 );
buf \U$9000 ( \17827_18126 , \17826_18125 );
xor \U$9001 ( \17828_18127 , \17821_18120 , \17827_18126 );
and \U$9002 ( \17829_18128 , \10996_10421 , \16013_16315_nG9bf0 );
and \U$9003 ( \17830_18129 , \10119_10418 , \16378_16680_nG9bed );
or \U$9004 ( \17831_18130 , \17829_18128 , \17830_18129 );
xor \U$9005 ( \17832_18131 , \10118_10417 , \17831_18130 );
buf \U$9006 ( \17833_18132 , \17832_18131 );
buf \U$9008 ( \17834_18133 , \17833_18132 );
xor \U$9009 ( \17835_18134 , \17828_18127 , \17834_18133 );
buf \U$9010 ( \17836_18135 , \17835_18134 );
xor \U$9011 ( \17837_18136 , \17816_18115 , \17836_18135 );
buf \U$9012 ( \17838_18137 , \17837_18136 );
and \U$9013 ( \17839_18138 , \17370_17672 , \17375_17677 );
and \U$9014 ( \17840_18139 , \17370_17672 , \17396_17698 );
and \U$9015 ( \17841_18140 , \17375_17677 , \17396_17698 );
or \U$9016 ( \17842_18141 , \17839_18138 , \17840_18139 , \17841_18140 );
buf \U$9017 ( \17843_18142 , \17842_18141 );
xor \U$9018 ( \17844_18143 , \17838_18137 , \17843_18142 );
and \U$9019 ( \17845_18144 , \17398_17700 , \17403_17705 );
and \U$9020 ( \17846_18145 , \17398_17700 , \17409_17711 );
and \U$9021 ( \17847_18146 , \17403_17705 , \17409_17711 );
or \U$9022 ( \17848_18147 , \17845_18144 , \17846_18145 , \17847_18146 );
buf \U$9023 ( \17849_18148 , \17848_18147 );
xor \U$9024 ( \17850_18149 , \17844_18143 , \17849_18148 );
and \U$9025 ( \17851_18150 , \17413_17715 , \17850_18149 );
and \U$9026 ( \17852_18151 , RIdec4a00_701, \8760_9059 );
and \U$9027 ( \17853_18152 , RIdec1d00_669, \8762_9061 );
and \U$9028 ( \17854_18153 , RIfcad7b0_6996, \8764_9063 );
and \U$9029 ( \17855_18154 , RIdebf000_637, \8766_9065 );
and \U$9030 ( \17856_18155 , RIfc64cb8_6169, \8768_9067 );
and \U$9031 ( \17857_18156 , RIdebc300_605, \8770_9069 );
and \U$9032 ( \17858_18157 , RIdeb9600_573, \8772_9071 );
and \U$9033 ( \17859_18158 , RIdeb6900_541, \8774_9073 );
and \U$9034 ( \17860_18159 , RIfc6f9b0_6292, \8776_9075 );
and \U$9035 ( \17861_18160 , RIdeb0f00_477, \8778_9077 );
and \U$9036 ( \17862_18161 , RIfc657f8_6177, \8780_9079 );
and \U$9037 ( \17863_18162 , RIdeae200_445, \8782_9081 );
and \U$9038 ( \17864_18163 , RIfce69c0_7646, \8784_9083 );
and \U$9039 ( \17865_18164 , RIdea8d28_413, \8786_9085 );
and \U$9040 ( \17866_18165 , RIdea2428_381, \8788_9087 );
and \U$9041 ( \17867_18166 , RIde9bb28_349, \8790_9089 );
and \U$9042 ( \17868_18167 , RIfc6fc80_6294, \8792_9091 );
and \U$9043 ( \17869_18168 , RIee1b760_4771, \8794_9093 );
and \U$9044 ( \17870_18169 , RIfca8080_6934, \8796_9095 );
and \U$9045 ( \17871_18170 , RIfe8b8f0_7932, \8798_9097 );
and \U$9046 ( \17872_18171 , RIde90020_292, \8800_9099 );
and \U$9047 ( \17873_18172 , RIde8c510_274, \8802_9101 );
and \U$9048 ( \17874_18173 , RIde89090_258, \8804_9103 );
and \U$9049 ( \17875_18174 , RIde84ba8_237, \8806_9105 );
and \U$9050 ( \17876_18175 , RIfc65ac8_6179, \8808_9107 );
and \U$9051 ( \17877_18176 , RIfcad210_6992, \8810_9109 );
and \U$9052 ( \17878_18177 , RIfcce168_7367, \8812_9111 );
and \U$9053 ( \17879_18178 , RIfcce2d0_7368, \8814_9113 );
and \U$9054 ( \17880_18179 , RIfc51488_5947, \8816_9115 );
and \U$9055 ( \17881_18180 , RIe16af40_2594, \8818_9117 );
and \U$9056 ( \17882_18181 , RIfc65c30_6180, \8820_9119 );
and \U$9057 ( \17883_18182 , RIe167598_2553, \8822_9121 );
and \U$9058 ( \17884_18183 , RIe164a00_2522, \8824_9123 );
and \U$9059 ( \17885_18184 , RIe161d00_2490, \8826_9125 );
and \U$9060 ( \17886_18185 , RIfc66e78_6193, \8828_9127 );
and \U$9061 ( \17887_18186 , RIe15f000_2458, \8830_9129 );
and \U$9062 ( \17888_18187 , RIfc6e498_6277, \8832_9131 );
and \U$9063 ( \17889_18188 , RIe15c300_2426, \8834_9133 );
and \U$9064 ( \17890_18189 , RIe156900_2362, \8836_9135 );
and \U$9065 ( \17891_18190 , RIe153c00_2330, \8838_9137 );
and \U$9066 ( \17892_18191 , RIfc6e330_6276, \8840_9139 );
and \U$9067 ( \17893_18192 , RIe150f00_2298, \8842_9141 );
and \U$9068 ( \17894_18193 , RIfccda60_7362, \8844_9143 );
and \U$9069 ( \17895_18194 , RIe14e200_2266, \8846_9145 );
and \U$9070 ( \17896_18195 , RIfc6e1c8_6275, \8848_9147 );
and \U$9071 ( \17897_18196 , RIe14b500_2234, \8850_9149 );
and \U$9072 ( \17898_18197 , RIe148800_2202, \8852_9151 );
and \U$9073 ( \17899_18198 , RIe145b00_2170, \8854_9153 );
and \U$9074 ( \17900_18199 , RIee33fb8_5050, \8856_9155 );
and \U$9075 ( \17901_18200 , RIee32d70_5037, \8858_9157 );
and \U$9076 ( \17902_18201 , RIee31c90_5025, \8860_9159 );
and \U$9077 ( \17903_18202 , RIee30fe8_5016, \8862_9161 );
and \U$9078 ( \17904_18203 , RIfea8630_8232, \8864_9163 );
and \U$9079 ( \17905_18204 , RIdf3e5a8_2086, \8866_9165 );
and \U$9080 ( \17906_18205 , RIdf3c550_2063, \8868_9167 );
and \U$9081 ( \17907_18206 , RIfea8798_8233, \8870_9169 );
and \U$9082 ( \17908_18207 , RIfc6e060_6274, \8872_9171 );
and \U$9083 ( \17909_18208 , RIfcac6d0_6984, \8874_9173 );
and \U$9084 ( \17910_18209 , RIfc56078_6001, \8876_9175 );
and \U$9085 ( \17911_18210 , RIfc6e600_6278, \8878_9177 );
and \U$9086 ( \17912_18211 , RIdf34dc8_1978, \8880_9179 );
and \U$9087 ( \17913_18212 , RIdf32d70_1955, \8882_9181 );
and \U$9088 ( \17914_18213 , RIfea84c8_8231, \8884_9183 );
and \U$9089 ( \17915_18214 , RIdf2eb58_1908, \8886_9185 );
or \U$9090 ( \17916_18215 , \17852_18151 , \17853_18152 , \17854_18153 , \17855_18154 , \17856_18155 , \17857_18156 , \17858_18157 , \17859_18158 , \17860_18159 , \17861_18160 , \17862_18161 , \17863_18162 , \17864_18163 , \17865_18164 , \17866_18165 , \17867_18166 , \17868_18167 , \17869_18168 , \17870_18169 , \17871_18170 , \17872_18171 , \17873_18172 , \17874_18173 , \17875_18174 , \17876_18175 , \17877_18176 , \17878_18177 , \17879_18178 , \17880_18179 , \17881_18180 , \17882_18181 , \17883_18182 , \17884_18183 , \17885_18184 , \17886_18185 , \17887_18186 , \17888_18187 , \17889_18188 , \17890_18189 , \17891_18190 , \17892_18191 , \17893_18192 , \17894_18193 , \17895_18194 , \17896_18195 , \17897_18196 , \17898_18197 , \17899_18198 , \17900_18199 , \17901_18200 , \17902_18201 , \17903_18202 , \17904_18203 , \17905_18204 , \17906_18205 , \17907_18206 , \17908_18207 , \17909_18208 , \17910_18209 , \17911_18210 , \17912_18211 , \17913_18212 , \17914_18213 , \17915_18214 );
and \U$9091 ( \17917_18216 , RIee2b750_4953, \8889_9188 );
and \U$9092 ( \17918_18217 , RIfc6ee70_6284, \8891_9190 );
and \U$9093 ( \17919_18218 , RIfc6efd8_6285, \8893_9192 );
and \U$9094 ( \17920_18219 , RIee27808_4908, \8895_9194 );
and \U$9095 ( \17921_18220 , RIfe8b788_7931, \8897_9196 );
and \U$9096 ( \17922_18221 , RIdf27ad8_1828, \8899_9198 );
and \U$9097 ( \17923_18222 , RIdf25d50_1807, \8901_9200 );
and \U$9098 ( \17924_18223 , RIdf24130_1787, \8903_9202 );
and \U$9099 ( \17925_18224 , RIfc66608_6187, \8905_9204 );
and \U$9100 ( \17926_18225 , RIfccde98_7365, \8907_9206 );
and \U$9101 ( \17927_18226 , RIfc66a40_6190, \8909_9208 );
and \U$9102 ( \17928_18227 , RIfc668d8_6189, \8911_9210 );
and \U$9103 ( \17929_18228 , RIfcacf40_6990, \8913_9212 );
and \U$9104 ( \17930_18229 , RIfeaaef8_8261, \8915_9214 );
and \U$9105 ( \17931_18230 , RIfc6e8d0_6280, \8917_9216 );
and \U$9106 ( \17932_18231 , RIdf18d30_1659, \8919_9218 );
and \U$9107 ( \17933_18232 , RIdf165d0_1631, \8921_9220 );
and \U$9108 ( \17934_18233 , RIdf138d0_1599, \8923_9222 );
and \U$9109 ( \17935_18234 , RIdf10bd0_1567, \8925_9224 );
and \U$9110 ( \17936_18235 , RIdf0ded0_1535, \8927_9226 );
and \U$9111 ( \17937_18236 , RIdf0b1d0_1503, \8929_9228 );
and \U$9112 ( \17938_18237 , RIdf084d0_1471, \8931_9230 );
and \U$9113 ( \17939_18238 , RIdf057d0_1439, \8933_9232 );
and \U$9114 ( \17940_18239 , RIdf02ad0_1407, \8935_9234 );
and \U$9115 ( \17941_18240 , RIdefd0d0_1343, \8937_9236 );
and \U$9116 ( \17942_18241 , RIdefa3d0_1311, \8939_9238 );
and \U$9117 ( \17943_18242 , RIdef76d0_1279, \8941_9240 );
and \U$9118 ( \17944_18243 , RIdef49d0_1247, \8943_9242 );
and \U$9119 ( \17945_18244 , RIdef1cd0_1215, \8945_9244 );
and \U$9120 ( \17946_18245 , RIdeeefd0_1183, \8947_9246 );
and \U$9121 ( \17947_18246 , RIdeec2d0_1151, \8949_9248 );
and \U$9122 ( \17948_18247 , RIdee95d0_1119, \8951_9250 );
and \U$9123 ( \17949_18248 , RIfc6dc28_6271, \8953_9252 );
and \U$9124 ( \17950_18249 , RIfc67c88_6203, \8955_9254 );
and \U$9125 ( \17951_18250 , RIfccb300_7334, \8957_9256 );
and \U$9126 ( \17952_18251 , RIfccd4c0_7358, \8959_9258 );
and \U$9127 ( \17953_18252 , RIfea81f8_8229, \8961_9260 );
and \U$9128 ( \17954_18253 , RIfea8360_8230, \8963_9262 );
and \U$9129 ( \17955_18254 , RIdee04f8_1016, \8965_9264 );
and \U$9130 ( \17956_18255 , RIdede338_992, \8967_9266 );
and \U$9131 ( \17957_18256 , RIfc6def8_6273, \8969_9268 );
and \U$9132 ( \17958_18257 , RIfcac130_6980, \8971_9270 );
and \U$9133 ( \17959_18258 , RIfc67b20_6202, \8973_9272 );
and \U$9134 ( \17960_18259 , RIfc67df0_6204, \8975_9274 );
and \U$9135 ( \17961_18260 , RIded9040_933, \8977_9276 );
and \U$9136 ( \17962_18261 , RIded6a48_906, \8979_9278 );
and \U$9137 ( \17963_18262 , RIded4b58_884, \8981_9280 );
and \U$9138 ( \17964_18263 , RIded26c8_858, \8983_9282 );
and \U$9139 ( \17965_18264 , RIdecfe00_829, \8985_9284 );
and \U$9140 ( \17966_18265 , RIdecd100_797, \8987_9286 );
and \U$9141 ( \17967_18266 , RIdeca400_765, \8989_9288 );
and \U$9142 ( \17968_18267 , RIdec7700_733, \8991_9290 );
and \U$9143 ( \17969_18268 , RIdeb3c00_509, \8993_9292 );
and \U$9144 ( \17970_18269 , RIde95228_317, \8995_9294 );
and \U$9145 ( \17971_18270 , RIe16d808_2623, \8997_9296 );
and \U$9146 ( \17972_18271 , RIe159600_2394, \8999_9298 );
and \U$9147 ( \17973_18272 , RIe142e00_2138, \9001_9300 );
and \U$9148 ( \17974_18273 , RIdf377f8_2008, \9003_9302 );
and \U$9149 ( \17975_18274 , RIdf2be58_1876, \9005_9304 );
and \U$9150 ( \17976_18275 , RIdf1c6d8_1700, \9007_9306 );
and \U$9151 ( \17977_18276 , RIdeffdd0_1375, \9009_9308 );
and \U$9152 ( \17978_18277 , RIdee68d0_1087, \9011_9310 );
and \U$9153 ( \17979_18278 , RIdedb638_960, \9013_9312 );
and \U$9154 ( \17980_18279 , RIde7b170_190, \9015_9314 );
or \U$9155 ( \17981_18280 , \17917_18216 , \17918_18217 , \17919_18218 , \17920_18219 , \17921_18220 , \17922_18221 , \17923_18222 , \17924_18223 , \17925_18224 , \17926_18225 , \17927_18226 , \17928_18227 , \17929_18228 , \17930_18229 , \17931_18230 , \17932_18231 , \17933_18232 , \17934_18233 , \17935_18234 , \17936_18235 , \17937_18236 , \17938_18237 , \17939_18238 , \17940_18239 , \17941_18240 , \17942_18241 , \17943_18242 , \17944_18243 , \17945_18244 , \17946_18245 , \17947_18246 , \17948_18247 , \17949_18248 , \17950_18249 , \17951_18250 , \17952_18251 , \17953_18252 , \17954_18253 , \17955_18254 , \17956_18255 , \17957_18256 , \17958_18257 , \17959_18258 , \17960_18259 , \17961_18260 , \17962_18261 , \17963_18262 , \17964_18263 , \17965_18264 , \17966_18265 , \17967_18266 , \17968_18267 , \17969_18268 , \17970_18269 , \17971_18270 , \17972_18271 , \17973_18272 , \17974_18273 , \17975_18274 , \17976_18275 , \17977_18276 , \17978_18277 , \17979_18278 , \17980_18279 );
or \U$9156 ( \17982_18281 , \17916_18215 , \17981_18280 );
_DC \g2a85/U$1 ( \17983 , \17982_18281 , \9024_9323 );
buf \U$9157 ( \17984_18283 , \17983 );
and \U$9158 ( \17985_18284 , RIe19cc98_3161, \9034_9333 );
and \U$9159 ( \17986_18285 , RIe199f98_3129, \9036_9335 );
and \U$9160 ( \17987_18286 , RIfc73088_6331, \9038_9337 );
and \U$9161 ( \17988_18287 , RIe197298_3097, \9040_9339 );
and \U$9162 ( \17989_18288 , RIf1442a8_5235, \9042_9341 );
and \U$9163 ( \17990_18289 , RIe194598_3065, \9044_9343 );
and \U$9164 ( \17991_18290 , RIe191898_3033, \9046_9345 );
and \U$9165 ( \17992_18291 , RIe18eb98_3001, \9048_9347 );
and \U$9166 ( \17993_18292 , RIe189198_2937, \9050_9349 );
and \U$9167 ( \17994_18293 , RIe186498_2905, \9052_9351 );
and \U$9168 ( \17995_18294 , RIfc72278_6321, \9054_9353 );
and \U$9169 ( \17996_18295 , RIe183798_2873, \9056_9355 );
and \U$9170 ( \17997_18296 , RIfc61ce8_6135, \9058_9357 );
and \U$9171 ( \17998_18297 , RIe180a98_2841, \9060_9359 );
and \U$9172 ( \17999_18298 , RIe17dd98_2809, \9062_9361 );
and \U$9173 ( \18000_18299 , RIe17b098_2777, \9064_9363 );
and \U$9174 ( \18001_18300 , RIfcaf268_7015, \9066_9365 );
and \U$9175 ( \18002_18301 , RIfca6a00_6918, \9068_9367 );
and \U$9176 ( \18003_18302 , RIfcc9b18_7317, \9070_9369 );
and \U$9177 ( \18004_18303 , RIe175530_2712, \9072_9371 );
and \U$9178 ( \18005_18304 , RIfc72818_6325, \9074_9373 );
and \U$9179 ( \18006_18305 , RIfc726b0_6324, \9076_9375 );
and \U$9180 ( \18007_18306 , RIfccf7e8_7383, \9078_9377 );
and \U$9181 ( \18008_18307 , RIfc72548_6323, \9080_9379 );
and \U$9182 ( \18009_18308 , RIee3be48_5140, \9082_9381 );
and \U$9183 ( \18010_18309 , RIee3ad68_5128, \9084_9383 );
and \U$9184 ( \18011_18310 , RIfc71fa8_6319, \9086_9385 );
and \U$9185 ( \18012_18311 , RIe1730a0_2686, \9088_9387 );
and \U$9186 ( \18013_18312 , RIfcaef98_7013, \9090_9389 );
and \U$9187 ( \18014_18313 , RIfccf518_7381, \9092_9391 );
and \U$9188 ( \18015_18314 , RIfc71e40_6318, \9094_9393 );
and \U$9189 ( \18016_18315 , RIfc62120_6138, \9096_9395 );
and \U$9190 ( \18017_18316 , RIfe8b350_7928, \9098_9397 );
and \U$9191 ( \18018_18317 , RIe222ff0_4688, \9100_9399 );
and \U$9192 ( \18019_18318 , RIfcc9f50_7320, \9102_9401 );
and \U$9193 ( \18020_18319 , RIe2202f0_4656, \9104_9403 );
and \U$9194 ( \18021_18320 , RIfc4a570_5868, \9106_9405 );
and \U$9195 ( \18022_18321 , RIe21d5f0_4624, \9108_9407 );
and \U$9196 ( \18023_18322 , RIe217bf0_4560, \9110_9409 );
and \U$9197 ( \18024_18323 , RIe214ef0_4528, \9112_9411 );
and \U$9198 ( \18025_18324 , RIfccf3b0_7380, \9114_9413 );
and \U$9199 ( \18026_18325 , RIe2121f0_4496, \9116_9415 );
and \U$9200 ( \18027_18326 , RIf168ba8_5651, \9118_9417 );
and \U$9201 ( \18028_18327 , RIe20f4f0_4464, \9120_9419 );
and \U$9202 ( \18029_18328 , RIfc71300_6310, \9122_9421 );
and \U$9203 ( \18030_18329 , RIe20c7f0_4432, \9124_9423 );
and \U$9204 ( \18031_18330 , RIe209af0_4400, \9126_9425 );
and \U$9205 ( \18032_18331 , RIe206df0_4368, \9128_9427 );
and \U$9206 ( \18033_18332 , RIfc718a0_6314, \9130_9429 );
and \U$9207 ( \18034_18333 , RIfc71a08_6315, \9132_9431 );
and \U$9208 ( \18035_18334 , RIe202098_4313, \9134_9433 );
and \U$9209 ( \18036_18335 , RIfe8b1e8_7927, \9136_9435 );
and \U$9210 ( \18037_18336 , RIfc715d0_6312, \9138_9437 );
and \U$9211 ( \18038_18337 , RIfce6588_7643, \9140_9439 );
and \U$9212 ( \18039_18338 , RIfc62c60_6146, \9142_9441 );
and \U$9213 ( \18040_18339 , RIf161858_5569, \9144_9443 );
and \U$9214 ( \18041_18340 , RIf15fad0_5548, \9146_9445 );
and \U$9215 ( \18042_18341 , RIf15dbe0_5526, \9148_9447 );
and \U$9216 ( \18043_18342 , RIe1fc698_4249, \9150_9449 );
and \U$9217 ( \18044_18343 , RIfe8b4b8_7929, \9152_9451 );
and \U$9218 ( \18045_18344 , RIfcae5c0_7006, \9154_9453 );
and \U$9219 ( \18046_18345 , RIfc63098_6149, \9156_9455 );
and \U$9220 ( \18047_18346 , RIfc63200_6150, \9158_9457 );
and \U$9221 ( \18048_18347 , RIfc71198_6309, \9160_9459 );
or \U$9222 ( \18049_18348 , \17985_18284 , \17986_18285 , \17987_18286 , \17988_18287 , \17989_18288 , \17990_18289 , \17991_18290 , \17992_18291 , \17993_18292 , \17994_18293 , \17995_18294 , \17996_18295 , \17997_18296 , \17998_18297 , \17999_18298 , \18000_18299 , \18001_18300 , \18002_18301 , \18003_18302 , \18004_18303 , \18005_18304 , \18006_18305 , \18007_18306 , \18008_18307 , \18009_18308 , \18010_18309 , \18011_18310 , \18012_18311 , \18013_18312 , \18014_18313 , \18015_18314 , \18016_18315 , \18017_18316 , \18018_18317 , \18019_18318 , \18020_18319 , \18021_18320 , \18022_18321 , \18023_18322 , \18024_18323 , \18025_18324 , \18026_18325 , \18027_18326 , \18028_18327 , \18029_18328 , \18030_18329 , \18031_18330 , \18032_18331 , \18033_18332 , \18034_18333 , \18035_18334 , \18036_18335 , \18037_18336 , \18038_18337 , \18039_18338 , \18040_18339 , \18041_18340 , \18042_18341 , \18043_18342 , \18044_18343 , \18045_18344 , \18046_18345 , \18047_18346 , \18048_18347 );
and \U$9223 ( \18050_18349 , RIf158a50_5468, \9163_9462 );
and \U$9224 ( \18051_18350 , RIf1576a0_5454, \9165_9464 );
and \U$9225 ( \18052_18351 , RIfcdc808_7531, \9167_9466 );
and \U$9226 ( \18053_18352 , RIfe8b620_7930, \9169_9468 );
and \U$9227 ( \18054_18353 , RIfc634d0_6152, \9171_9470 );
and \U$9228 ( \18055_18354 , RIfcceb40_7374, \9173_9472 );
and \U$9229 ( \18056_18355 , RIf154400_5418, \9175_9474 );
and \U$9230 ( \18057_18356 , RIe1f4da8_4163, \9177_9476 );
and \U$9231 ( \18058_18357 , RIf152c18_5401, \9179_9478 );
and \U$9232 ( \18059_18358 , RIf151868_5387, \9181_9480 );
and \U$9233 ( \18060_18359 , RIfc4d108_5899, \9183_9482 );
and \U$9234 ( \18061_18360 , RIe1f2a80_4138, \9185_9484 );
and \U$9235 ( \18062_18361 , RIfc70a90_6304, \9187_9486 );
and \U$9236 ( \18063_18362 , RIfc63bd8_6157, \9189_9488 );
and \U$9237 ( \18064_18363 , RIfca7810_6928, \9191_9490 );
and \U$9238 ( \18065_18364 , RIe1ed788_4079, \9193_9492 );
and \U$9239 ( \18066_18365 , RIe1ead58_4049, \9195_9494 );
and \U$9240 ( \18067_18366 , RIe1e8058_4017, \9197_9496 );
and \U$9241 ( \18068_18367 , RIe1e5358_3985, \9199_9498 );
and \U$9242 ( \18069_18368 , RIe1e2658_3953, \9201_9500 );
and \U$9243 ( \18070_18369 , RIe1df958_3921, \9203_9502 );
and \U$9244 ( \18071_18370 , RIe1dcc58_3889, \9205_9504 );
and \U$9245 ( \18072_18371 , RIe1d9f58_3857, \9207_9506 );
and \U$9246 ( \18073_18372 , RIe1d7258_3825, \9209_9508 );
and \U$9247 ( \18074_18373 , RIe1d1858_3761, \9211_9510 );
and \U$9248 ( \18075_18374 , RIe1ceb58_3729, \9213_9512 );
and \U$9249 ( \18076_18375 , RIe1cbe58_3697, \9215_9514 );
and \U$9250 ( \18077_18376 , RIe1c9158_3665, \9217_9516 );
and \U$9251 ( \18078_18377 , RIe1c6458_3633, \9219_9518 );
and \U$9252 ( \18079_18378 , RIe1c3758_3601, \9221_9520 );
and \U$9253 ( \18080_18379 , RIe1c0a58_3569, \9223_9522 );
and \U$9254 ( \18081_18380 , RIe1bdd58_3537, \9225_9524 );
and \U$9255 ( \18082_18381 , RIf14c408_5327, \9227_9526 );
and \U$9256 ( \18083_18382 , RIf14b1c0_5314, \9229_9528 );
and \U$9257 ( \18084_18383 , RIe1b8d30_3480, \9231_9530 );
and \U$9258 ( \18085_18384 , RIe1b6cd8_3457, \9233_9532 );
and \U$9259 ( \18086_18385 , RIfc707c0_6302, \9235_9534 );
and \U$9260 ( \18087_18386 , RIfca7c48_6931, \9237_9536 );
and \U$9261 ( \18088_18387 , RIe1b4de8_3435, \9239_9538 );
and \U$9262 ( \18089_18388 , RIe1b3a38_3421, \9241_9540 );
and \U$9263 ( \18090_18389 , RIfc70220_6298, \9243_9542 );
and \U$9264 ( \18091_18390 , RIfcce870_7372, \9245_9544 );
and \U$9265 ( \18092_18391 , RIe1b23b8_3405, \9247_9546 );
and \U$9266 ( \18093_18392 , RIe1b0630_3384, \9249_9548 );
and \U$9267 ( \18094_18393 , RIfc645b0_6164, \9251_9550 );
and \U$9268 ( \18095_18394 , RIfc700b8_6297, \9253_9552 );
and \U$9269 ( \18096_18395 , RIfeaac28_8259, \9255_9554 );
and \U$9270 ( \18097_18396 , RIe1aa690_3316, \9257_9556 );
and \U$9271 ( \18098_18397 , RIe1a8098_3289, \9259_9558 );
and \U$9272 ( \18099_18398 , RIe1a5398_3257, \9261_9560 );
and \U$9273 ( \18100_18399 , RIe1a2698_3225, \9263_9562 );
and \U$9274 ( \18101_18400 , RIe19f998_3193, \9265_9564 );
and \U$9275 ( \18102_18401 , RIe18be98_2969, \9267_9566 );
and \U$9276 ( \18103_18402 , RIe178398_2745, \9269_9568 );
and \U$9277 ( \18104_18403 , RIe225cf0_4720, \9271_9570 );
and \U$9278 ( \18105_18404 , RIe21a8f0_4592, \9273_9572 );
and \U$9279 ( \18106_18405 , RIe2040f0_4336, \9275_9574 );
and \U$9280 ( \18107_18406 , RIe1fe150_4268, \9277_9576 );
and \U$9281 ( \18108_18407 , RIe1f7508_4191, \9279_9578 );
and \U$9282 ( \18109_18408 , RIe1f0050_4108, \9281_9580 );
and \U$9283 ( \18110_18409 , RIe1d4558_3793, \9283_9582 );
and \U$9284 ( \18111_18410 , RIe1bb058_3505, \9285_9584 );
and \U$9285 ( \18112_18411 , RIe1aded0_3356, \9287_9586 );
and \U$9286 ( \18113_18412 , RIe170508_2655, \9289_9588 );
or \U$9287 ( \18114_18413 , \18050_18349 , \18051_18350 , \18052_18351 , \18053_18352 , \18054_18353 , \18055_18354 , \18056_18355 , \18057_18356 , \18058_18357 , \18059_18358 , \18060_18359 , \18061_18360 , \18062_18361 , \18063_18362 , \18064_18363 , \18065_18364 , \18066_18365 , \18067_18366 , \18068_18367 , \18069_18368 , \18070_18369 , \18071_18370 , \18072_18371 , \18073_18372 , \18074_18373 , \18075_18374 , \18076_18375 , \18077_18376 , \18078_18377 , \18079_18378 , \18080_18379 , \18081_18380 , \18082_18381 , \18083_18382 , \18084_18383 , \18085_18384 , \18086_18385 , \18087_18386 , \18088_18387 , \18089_18388 , \18090_18389 , \18091_18390 , \18092_18391 , \18093_18392 , \18094_18393 , \18095_18394 , \18096_18395 , \18097_18396 , \18098_18397 , \18099_18398 , \18100_18399 , \18101_18400 , \18102_18401 , \18103_18402 , \18104_18403 , \18105_18404 , \18106_18405 , \18107_18406 , \18108_18407 , \18109_18408 , \18110_18409 , \18111_18410 , \18112_18411 , \18113_18412 );
or \U$9288 ( \18115_18414 , \18049_18348 , \18114_18413 );
_DC \g3bb2/U$1 ( \18116 , \18115_18414 , \9298_9597 );
buf \U$9289 ( \18117_18416 , \18116 );
xor \U$9290 ( \18118_18417 , \17984_18283 , \18117_18416 );
and \U$9291 ( \18119_18418 , RIdec4898_700, \8760_9059 );
and \U$9292 ( \18120_18419 , RIdec1b98_668, \8762_9061 );
and \U$9293 ( \18121_18420 , RIfc661d0_6184, \8764_9063 );
and \U$9294 ( \18122_18421 , RIdebee98_636, \8766_9065 );
and \U$9295 ( \18123_18422 , RIfce6b28_7647, \8768_9067 );
and \U$9296 ( \18124_18423 , RIdebc198_604, \8770_9069 );
and \U$9297 ( \18125_18424 , RIdeb9498_572, \8772_9071 );
and \U$9298 ( \18126_18425 , RIdeb6798_540, \8774_9073 );
and \U$9299 ( \18127_18426 , RIfc40d18_5763, \8776_9075 );
and \U$9300 ( \18128_18427 , RIdeb0d98_476, \8778_9077 );
and \U$9301 ( \18129_18428 , RIfcad648_6995, \8780_9079 );
and \U$9302 ( \18130_18429 , RIdeae098_444, \8782_9081 );
and \U$9303 ( \18131_18430 , RIfcaa510_6960, \8784_9083 );
and \U$9304 ( \18132_18431 , RIdea89e0_412, \8786_9085 );
and \U$9305 ( \18133_18432 , RIdea20e0_380, \8788_9087 );
and \U$9306 ( \18134_18433 , RIde9b7e0_348, \8790_9089 );
and \U$9307 ( \18135_18434 , RIfcab320_6970, \8792_9091 );
and \U$9308 ( \18136_18435 , RIfca8350_6936, \8794_9093 );
and \U$9309 ( \18137_18436 , RIfc6f6e0_6290, \8796_9095 );
and \U$9310 ( \18138_18437 , RIfcaa240_6958, \8798_9097 );
and \U$9311 ( \18139_18438 , RIde8fcd8_291, \8800_9099 );
and \U$9312 ( \18140_18439 , RIfe8aae0_7922, \8802_9101 );
and \U$9313 ( \18141_18440 , RIde88d48_257, \8804_9103 );
and \U$9314 ( \18142_18441 , RIde84860_236, \8806_9105 );
and \U$9315 ( \18143_18442 , RIde80a08_217, \8808_9107 );
and \U$9316 ( \18144_18443 , RIfc64718_6165, \8810_9109 );
and \U$9317 ( \18145_18444 , RIfcae020_7002, \8812_9111 );
and \U$9318 ( \18146_18445 , RIfcadeb8_7001, \8814_9113 );
and \U$9319 ( \18147_18446 , RIee38fe0_5107, \8816_9115 );
and \U$9320 ( \18148_18447 , RIe16add8_2593, \8818_9117 );
and \U$9321 ( \18149_18448 , RIe1695f0_2576, \8820_9119 );
and \U$9322 ( \18150_18449 , RIe167430_2552, \8822_9121 );
and \U$9323 ( \18151_18450 , RIe164898_2521, \8824_9123 );
and \U$9324 ( \18152_18451 , RIe161b98_2489, \8826_9125 );
and \U$9325 ( \18153_18452 , RIfe8a3d8_7917, \8828_9127 );
and \U$9326 ( \18154_18453 , RIe15ee98_2457, \8830_9129 );
and \U$9327 ( \18155_18454 , RIfe8a270_7916, \8832_9131 );
and \U$9328 ( \18156_18455 , RIe15c198_2425, \8834_9133 );
and \U$9329 ( \18157_18456 , RIe156798_2361, \8836_9135 );
and \U$9330 ( \18158_18457 , RIe153a98_2329, \8838_9137 );
and \U$9331 ( \18159_18458 , RIfc3f0f8_5743, \8840_9139 );
and \U$9332 ( \18160_18459 , RIe150d98_2297, \8842_9141 );
and \U$9333 ( \18161_18460 , RIfcab050_6968, \8844_9143 );
and \U$9334 ( \18162_18461 , RIe14e098_2265, \8846_9145 );
and \U$9335 ( \18163_18462 , RIfcca658_7325, \8848_9147 );
and \U$9336 ( \18164_18463 , RIe14b398_2233, \8850_9149 );
and \U$9337 ( \18165_18464 , RIe148698_2201, \8852_9151 );
and \U$9338 ( \18166_18465 , RIe145998_2169, \8854_9153 );
and \U$9339 ( \18167_18466 , RIfe8a810_7920, \8856_9155 );
and \U$9340 ( \18168_18467 , RIfe8a6a8_7919, \8858_9157 );
and \U$9341 ( \18169_18468 , RIee31b28_5024, \8860_9159 );
and \U$9342 ( \18170_18469 , RIee30e80_5015, \8862_9161 );
and \U$9343 ( \18171_18470 , RIe140808_2111, \8864_9163 );
and \U$9344 ( \18172_18471 , RIfe8a540_7918, \8866_9165 );
and \U$9345 ( \18173_18472 , RIdf3c3e8_2062, \8868_9167 );
and \U$9346 ( \18174_18473 , RIdf3a0c0_2037, \8870_9169 );
and \U$9347 ( \18175_18474 , RIfc6b1f8_6241, \8872_9171 );
and \U$9348 ( \18176_18475 , RIee2f260_4995, \8874_9173 );
and \U$9349 ( \18177_18476 , RIfc70d60_6306, \8876_9175 );
and \U$9350 ( \18178_18477 , RIee2d0a0_4971, \8878_9177 );
and \U$9351 ( \18179_18478 , RIfe8a978_7921, \8880_9179 );
and \U$9352 ( \18180_18479 , RIdf32c08_1954, \8882_9181 );
and \U$9353 ( \18181_18480 , RIdf308e0_1929, \8884_9183 );
and \U$9354 ( \18182_18481 , RIdf2e9f0_1907, \8886_9185 );
or \U$9355 ( \18183_18482 , \18119_18418 , \18120_18419 , \18121_18420 , \18122_18421 , \18123_18422 , \18124_18423 , \18125_18424 , \18126_18425 , \18127_18426 , \18128_18427 , \18129_18428 , \18130_18429 , \18131_18430 , \18132_18431 , \18133_18432 , \18134_18433 , \18135_18434 , \18136_18435 , \18137_18436 , \18138_18437 , \18139_18438 , \18140_18439 , \18141_18440 , \18142_18441 , \18143_18442 , \18144_18443 , \18145_18444 , \18146_18445 , \18147_18446 , \18148_18447 , \18149_18448 , \18150_18449 , \18151_18450 , \18152_18451 , \18153_18452 , \18154_18453 , \18155_18454 , \18156_18455 , \18157_18456 , \18158_18457 , \18159_18458 , \18160_18459 , \18161_18460 , \18162_18461 , \18163_18462 , \18164_18463 , \18165_18464 , \18166_18465 , \18167_18466 , \18168_18467 , \18169_18468 , \18170_18469 , \18171_18470 , \18172_18471 , \18173_18472 , \18174_18473 , \18175_18474 , \18176_18475 , \18177_18476 , \18178_18477 , \18179_18478 , \18180_18479 , \18181_18480 , \18182_18481 );
and \U$9356 ( \18184_18483 , RIee2b5e8_4952, \8889_9188 );
and \U$9357 ( \18185_18484 , RIee29e00_4935, \8891_9190 );
and \U$9358 ( \18186_18485 , RIee28a50_4921, \8893_9192 );
and \U$9359 ( \18187_18486 , RIee276a0_4907, \8895_9194 );
and \U$9360 ( \18188_18487 , RIdf29c98_1852, \8897_9196 );
and \U$9361 ( \18189_18488 , RIdf27970_1827, \8899_9198 );
and \U$9362 ( \18190_18489 , RIdf25be8_1806, \8901_9200 );
and \U$9363 ( \18191_18490 , RIdf23fc8_1786, \8903_9202 );
and \U$9364 ( \18192_18491 , RIfc6aaf0_6236, \8905_9204 );
and \U$9365 ( \18193_18492 , RIfc6ac58_6237, \8907_9206 );
and \U$9366 ( \18194_18493 , RIdf22678_1768, \8909_9208 );
and \U$9367 ( \18195_18494 , RIfcdd4b0_7540, \8911_9210 );
and \U$9368 ( \18196_18495 , RIdf21160_1753, \8913_9212 );
and \U$9369 ( \18197_18496 , RIdf1f108_1730, \8915_9214 );
and \U$9370 ( \18198_18497 , RIdf1ac20_1681, \8917_9216 );
and \U$9371 ( \18199_18498 , RIfeaa7f0_8256, \8919_9218 );
and \U$9372 ( \18200_18499 , RIdf16468_1630, \8921_9220 );
and \U$9373 ( \18201_18500 , RIdf13768_1598, \8923_9222 );
and \U$9374 ( \18202_18501 , RIdf10a68_1566, \8925_9224 );
and \U$9375 ( \18203_18502 , RIdf0dd68_1534, \8927_9226 );
and \U$9376 ( \18204_18503 , RIdf0b068_1502, \8929_9228 );
and \U$9377 ( \18205_18504 , RIdf08368_1470, \8931_9230 );
and \U$9378 ( \18206_18505 , RIdf05668_1438, \8933_9232 );
and \U$9379 ( \18207_18506 , RIdf02968_1406, \8935_9234 );
and \U$9380 ( \18208_18507 , RIdefcf68_1342, \8937_9236 );
and \U$9381 ( \18209_18508 , RIdefa268_1310, \8939_9238 );
and \U$9382 ( \18210_18509 , RIdef7568_1278, \8941_9240 );
and \U$9383 ( \18211_18510 , RIdef4868_1246, \8943_9242 );
and \U$9384 ( \18212_18511 , RIdef1b68_1214, \8945_9244 );
and \U$9385 ( \18213_18512 , RIdeeee68_1182, \8947_9246 );
and \U$9386 ( \18214_18513 , RIdeec168_1150, \8949_9248 );
and \U$9387 ( \18215_18514 , RIdee9468_1118, \8951_9250 );
and \U$9388 ( \18216_18515 , RIee25378_4882, \8953_9252 );
and \U$9389 ( \18217_18516 , RIee24568_4872, \8955_9254 );
and \U$9390 ( \18218_18517 , RIee23a28_4864, \8957_9256 );
and \U$9391 ( \18219_18518 , RIee23050_4857, \8959_9258 );
and \U$9392 ( \18220_18519 , RIfe8adb0_7924, \8961_9260 );
and \U$9393 ( \18221_18520 , RIdee23e8_1038, \8963_9262 );
and \U$9394 ( \18222_18521 , RIfe8ac48_7923, \8965_9264 );
and \U$9395 ( \18223_18522 , RIdede1d0_991, \8967_9266 );
and \U$9396 ( \18224_18523 , RIfca5650_6904, \8969_9268 );
and \U$9397 ( \18225_18524 , RIee220d8_4846, \8971_9270 );
and \U$9398 ( \18226_18525 , RIfceeb20_7738, \8973_9272 );
and \U$9399 ( \18227_18526 , RIee20ff8_4834, \8975_9274 );
and \U$9400 ( \18228_18527 , RIded8ed8_932, \8977_9276 );
and \U$9401 ( \18229_18528 , RIfe8af18_7925, \8979_9278 );
and \U$9402 ( \18230_18529 , RIded49f0_883, \8981_9280 );
and \U$9403 ( \18231_18530 , RIfe8b080_7926, \8983_9282 );
and \U$9404 ( \18232_18531 , RIdecfc98_828, \8985_9284 );
and \U$9405 ( \18233_18532 , RIdeccf98_796, \8987_9286 );
and \U$9406 ( \18234_18533 , RIdeca298_764, \8989_9288 );
and \U$9407 ( \18235_18534 , RIdec7598_732, \8991_9290 );
and \U$9408 ( \18236_18535 , RIdeb3a98_508, \8993_9292 );
and \U$9409 ( \18237_18536 , RIde94ee0_316, \8995_9294 );
and \U$9410 ( \18238_18537 , RIe16d6a0_2622, \8997_9296 );
and \U$9411 ( \18239_18538 , RIe159498_2393, \8999_9298 );
and \U$9412 ( \18240_18539 , RIe142c98_2137, \9001_9300 );
and \U$9413 ( \18241_18540 , RIdf37690_2007, \9003_9302 );
and \U$9414 ( \18242_18541 , RIdf2bcf0_1875, \9005_9304 );
and \U$9415 ( \18243_18542 , RIdf1c570_1699, \9007_9306 );
and \U$9416 ( \18244_18543 , RIdeffc68_1374, \9009_9308 );
and \U$9417 ( \18245_18544 , RIdee6768_1086, \9011_9310 );
and \U$9418 ( \18246_18545 , RIdedb4d0_959, \9013_9312 );
and \U$9419 ( \18247_18546 , RIde7ae28_189, \9015_9314 );
or \U$9420 ( \18248_18547 , \18184_18483 , \18185_18484 , \18186_18485 , \18187_18486 , \18188_18487 , \18189_18488 , \18190_18489 , \18191_18490 , \18192_18491 , \18193_18492 , \18194_18493 , \18195_18494 , \18196_18495 , \18197_18496 , \18198_18497 , \18199_18498 , \18200_18499 , \18201_18500 , \18202_18501 , \18203_18502 , \18204_18503 , \18205_18504 , \18206_18505 , \18207_18506 , \18208_18507 , \18209_18508 , \18210_18509 , \18211_18510 , \18212_18511 , \18213_18512 , \18214_18513 , \18215_18514 , \18216_18515 , \18217_18516 , \18218_18517 , \18219_18518 , \18220_18519 , \18221_18520 , \18222_18521 , \18223_18522 , \18224_18523 , \18225_18524 , \18226_18525 , \18227_18526 , \18228_18527 , \18229_18528 , \18230_18529 , \18231_18530 , \18232_18531 , \18233_18532 , \18234_18533 , \18235_18534 , \18236_18535 , \18237_18536 , \18238_18537 , \18239_18538 , \18240_18539 , \18241_18540 , \18242_18541 , \18243_18542 , \18244_18543 , \18245_18544 , \18246_18545 , \18247_18546 );
or \U$9421 ( \18249_18548 , \18183_18482 , \18248_18547 );
_DC \g2b0a/U$1 ( \18250 , \18249_18548 , \9024_9323 );
buf \U$9422 ( \18251_18550 , \18250 );
and \U$9423 ( \18252_18551 , RIe19cb30_3160, \9034_9333 );
and \U$9424 ( \18253_18552 , RIe199e30_3128, \9036_9335 );
and \U$9425 ( \18254_18553 , RIf145388_5247, \9038_9337 );
and \U$9426 ( \18255_18554 , RIe197130_3096, \9040_9339 );
and \U$9427 ( \18256_18555 , RIfe8a108_7915, \9042_9341 );
and \U$9428 ( \18257_18556 , RIe194430_3064, \9044_9343 );
and \U$9429 ( \18258_18557 , RIe191730_3032, \9046_9345 );
and \U$9430 ( \18259_18558 , RIe18ea30_3000, \9048_9347 );
and \U$9431 ( \18260_18559 , RIe189030_2936, \9050_9349 );
and \U$9432 ( \18261_18560 , RIe186330_2904, \9052_9351 );
and \U$9433 ( \18262_18561 , RIfc6c878_6257, \9054_9353 );
and \U$9434 ( \18263_18562 , RIe183630_2872, \9056_9355 );
and \U$9435 ( \18264_18563 , RIfcabcf8_6977, \9058_9357 );
and \U$9436 ( \18265_18564 , RIe180930_2840, \9060_9359 );
and \U$9437 ( \18266_18565 , RIe17dc30_2808, \9062_9361 );
and \U$9438 ( \18267_18566 , RIe17af30_2776, \9064_9363 );
and \U$9439 ( \18268_18567 , RIfcccc50_7352, \9066_9365 );
and \U$9440 ( \18269_18568 , RIfcccdb8_7353, \9068_9367 );
and \U$9441 ( \18270_18569 , RIe176d18_2729, \9070_9369 );
and \U$9442 ( \18271_18570 , RIfea7af0_8224, \9072_9371 );
and \U$9443 ( \18272_18571 , RIfe89fa0_7914, \9074_9373 );
and \U$9444 ( \18273_18572 , RIfe89e38_7913, \9076_9375 );
and \U$9445 ( \18274_18573 , RIfcdd078_7537, \9078_9377 );
and \U$9446 ( \18275_18574 , RIfccb738_7337, \9080_9379 );
and \U$9447 ( \18276_18575 , RIfca9868_6951, \9082_9381 );
and \U$9448 ( \18277_18576 , RIfcabb90_6976, \9084_9383 );
and \U$9449 ( \18278_18577 , RIfca99d0_6952, \9086_9385 );
and \U$9450 ( \18279_18578 , RIe172f38_2685, \9088_9387 );
and \U$9451 ( \18280_18579 , RIf16fd90_5732, \9090_9389 );
and \U$9452 ( \18281_18580 , RIf16f250_5724, \9092_9391 );
and \U$9453 ( \18282_18581 , RIfc6c440_6254, \9094_9393 );
and \U$9454 ( \18283_18582 , RIfcaba28_6975, \9096_9395 );
and \U$9455 ( \18284_18583 , RIfc40610_5758, \9098_9397 );
and \U$9456 ( \18285_18584 , RIe222e88_4687, \9100_9399 );
and \U$9457 ( \18286_18585 , RIfc5d260_6082, \9102_9401 );
and \U$9458 ( \18287_18586 , RIe220188_4655, \9104_9403 );
and \U$9459 ( \18288_18587 , RIfcab758_6973, \9106_9405 );
and \U$9460 ( \18289_18588 , RIe21d488_4623, \9108_9407 );
and \U$9461 ( \18290_18589 , RIe217a88_4559, \9110_9409 );
and \U$9462 ( \18291_18590 , RIe214d88_4527, \9112_9411 );
and \U$9463 ( \18292_18591 , RIfe892f8_7905, \9114_9413 );
and \U$9464 ( \18293_18592 , RIe212088_4495, \9116_9415 );
and \U$9465 ( \18294_18593 , RIf168a40_5650, \9118_9417 );
and \U$9466 ( \18295_18594 , RIe20f388_4463, \9120_9419 );
and \U$9467 ( \18296_18595 , RIf167ac8_5639, \9122_9421 );
and \U$9468 ( \18297_18596 , RIe20c688_4431, \9124_9423 );
and \U$9469 ( \18298_18597 , RIe209988_4399, \9126_9425 );
and \U$9470 ( \18299_18598 , RIe206c88_4367, \9128_9427 );
and \U$9471 ( \18300_18599 , RIfc6c2d8_6253, \9130_9429 );
and \U$9472 ( \18301_18600 , RIfceec88_7739, \9132_9431 );
and \U$9473 ( \18302_18601 , RIe201f30_4312, \9134_9433 );
and \U$9474 ( \18303_18602 , RIe200748_4295, \9136_9435 );
and \U$9475 ( \18304_18603 , RIf164dc8_5607, \9138_9437 );
and \U$9476 ( \18305_18604 , RIf163fb8_5597, \9140_9439 );
and \U$9477 ( \18306_18605 , RIf163040_5586, \9142_9441 );
and \U$9478 ( \18307_18606 , RIfe895c8_7907, \9144_9443 );
and \U$9479 ( \18308_18607 , RIf15f968_5547, \9146_9445 );
and \U$9480 ( \18309_18608 , RIfe89898_7909, \9148_9447 );
and \U$9481 ( \18310_18609 , RIfe89460_7906, \9150_9449 );
and \U$9482 ( \18311_18610 , RIe1fb5b8_4237, \9152_9451 );
and \U$9483 ( \18312_18611 , RIf15c6c8_5511, \9154_9453 );
and \U$9484 ( \18313_18612 , RIfe89730_7908, \9156_9455 );
and \U$9485 ( \18314_18613 , RIf15a238_5485, \9158_9457 );
and \U$9486 ( \18315_18614 , RIf1599c8_5479, \9160_9459 );
or \U$9487 ( \18316_18615 , \18252_18551 , \18253_18552 , \18254_18553 , \18255_18554 , \18256_18555 , \18257_18556 , \18258_18557 , \18259_18558 , \18260_18559 , \18261_18560 , \18262_18561 , \18263_18562 , \18264_18563 , \18265_18564 , \18266_18565 , \18267_18566 , \18268_18567 , \18269_18568 , \18270_18569 , \18271_18570 , \18272_18571 , \18273_18572 , \18274_18573 , \18275_18574 , \18276_18575 , \18277_18576 , \18278_18577 , \18279_18578 , \18280_18579 , \18281_18580 , \18282_18581 , \18283_18582 , \18284_18583 , \18285_18584 , \18286_18585 , \18287_18586 , \18288_18587 , \18289_18588 , \18290_18589 , \18291_18590 , \18292_18591 , \18293_18592 , \18294_18593 , \18295_18594 , \18296_18595 , \18297_18596 , \18298_18597 , \18299_18598 , \18300_18599 , \18301_18600 , \18302_18601 , \18303_18602 , \18304_18603 , \18305_18604 , \18306_18605 , \18307_18606 , \18308_18607 , \18309_18608 , \18310_18609 , \18311_18610 , \18312_18611 , \18313_18612 , \18314_18613 , \18315_18614 );
and \U$9488 ( \18317_18616 , RIf1588e8_5467, \9163_9462 );
and \U$9489 ( \18318_18617 , RIfe89cd0_7912, \9165_9464 );
and \U$9490 ( \18319_18618 , RIfc5ba78_6065, \9167_9466 );
and \U$9491 ( \18320_18619 , RIe1f9c68_4219, \9169_9468 );
and \U$9492 ( \18321_18620 , RIfc5bd48_6067, \9171_9470 );
and \U$9493 ( \18322_18621 , RIf1554e0_5430, \9173_9472 );
and \U$9494 ( \18323_18622 , RIf154298_5417, \9175_9474 );
and \U$9495 ( \18324_18623 , RIe1f4c40_4162, \9177_9476 );
and \U$9496 ( \18325_18624 , RIfe89b68_7911, \9179_9478 );
and \U$9497 ( \18326_18625 , RIfe89a00_7910, \9181_9480 );
and \U$9498 ( \18327_18626 , RIf150350_5372, \9183_9482 );
and \U$9499 ( \18328_18627 , RIe1f2918_4137, \9185_9484 );
and \U$9500 ( \18329_18628 , RIf14f3d8_5361, \9187_9486 );
and \U$9501 ( \18330_18629 , RIfccc818_7349, \9189_9488 );
and \U$9502 ( \18331_18630 , RIf14d920_5342, \9191_9490 );
and \U$9503 ( \18332_18631 , RIe1ed620_4078, \9193_9492 );
and \U$9504 ( \18333_18632 , RIe1eabf0_4048, \9195_9494 );
and \U$9505 ( \18334_18633 , RIe1e7ef0_4016, \9197_9496 );
and \U$9506 ( \18335_18634 , RIe1e51f0_3984, \9199_9498 );
and \U$9507 ( \18336_18635 , RIe1e24f0_3952, \9201_9500 );
and \U$9508 ( \18337_18636 , RIe1df7f0_3920, \9203_9502 );
and \U$9509 ( \18338_18637 , RIe1dcaf0_3888, \9205_9504 );
and \U$9510 ( \18339_18638 , RIe1d9df0_3856, \9207_9506 );
and \U$9511 ( \18340_18639 , RIe1d70f0_3824, \9209_9508 );
and \U$9512 ( \18341_18640 , RIe1d16f0_3760, \9211_9510 );
and \U$9513 ( \18342_18641 , RIe1ce9f0_3728, \9213_9512 );
and \U$9514 ( \18343_18642 , RIe1cbcf0_3696, \9215_9514 );
and \U$9515 ( \18344_18643 , RIe1c8ff0_3664, \9217_9516 );
and \U$9516 ( \18345_18644 , RIe1c62f0_3632, \9219_9518 );
and \U$9517 ( \18346_18645 , RIe1c35f0_3600, \9221_9520 );
and \U$9518 ( \18347_18646 , RIe1c08f0_3568, \9223_9522 );
and \U$9519 ( \18348_18647 , RIe1bdbf0_3536, \9225_9524 );
and \U$9520 ( \18349_18648 , RIfc680c0_6206, \9227_9526 );
and \U$9521 ( \18350_18649 , RIf14b058_5313, \9229_9528 );
and \U$9522 ( \18351_18650 , RIe1b8bc8_3479, \9231_9530 );
and \U$9523 ( \18352_18651 , RIe1b6b70_3456, \9233_9532 );
and \U$9524 ( \18353_18652 , RIfcac298_6981, \9235_9534 );
and \U$9525 ( \18354_18653 , RIf1499d8_5297, \9237_9536 );
and \U$9526 ( \18355_18654 , RIfe89190_7904, \9239_9538 );
and \U$9527 ( \18356_18655 , RIfec19c8_8323, \9241_9540 );
and \U$9528 ( \18357_18656 , RIf148a60_5286, \9243_9542 );
and \U$9529 ( \18358_18657 , RIfccdd30_7364, \9245_9544 );
and \U$9530 ( \18359_18658 , RIe1b2250_3404, \9247_9546 );
and \U$9531 ( \18360_18659 , RIfec1860_8322, \9249_9548 );
and \U$9532 ( \18361_18660 , RIfc6e768_6279, \9251_9550 );
and \U$9533 ( \18362_18661 , RIfc54728_5983, \9253_9552 );
and \U$9534 ( \18363_18662 , RIe1abfe0_3334, \9255_9554 );
and \U$9535 ( \18364_18663 , RIe1aa528_3315, \9257_9556 );
and \U$9536 ( \18365_18664 , RIe1a7f30_3288, \9259_9558 );
and \U$9537 ( \18366_18665 , RIe1a5230_3256, \9261_9560 );
and \U$9538 ( \18367_18666 , RIe1a2530_3224, \9263_9562 );
and \U$9539 ( \18368_18667 , RIe19f830_3192, \9265_9564 );
and \U$9540 ( \18369_18668 , RIe18bd30_2968, \9267_9566 );
and \U$9541 ( \18370_18669 , RIe178230_2744, \9269_9568 );
and \U$9542 ( \18371_18670 , RIe225b88_4719, \9271_9570 );
and \U$9543 ( \18372_18671 , RIe21a788_4591, \9273_9572 );
and \U$9544 ( \18373_18672 , RIe203f88_4335, \9275_9574 );
and \U$9545 ( \18374_18673 , RIe1fdfe8_4267, \9277_9576 );
and \U$9546 ( \18375_18674 , RIe1f73a0_4190, \9279_9578 );
and \U$9547 ( \18376_18675 , RIe1efee8_4107, \9281_9580 );
and \U$9548 ( \18377_18676 , RIe1d43f0_3792, \9283_9582 );
and \U$9549 ( \18378_18677 , RIe1baef0_3504, \9285_9584 );
and \U$9550 ( \18379_18678 , RIe1add68_3355, \9287_9586 );
and \U$9551 ( \18380_18679 , RIe1703a0_2654, \9289_9588 );
or \U$9552 ( \18381_18680 , \18317_18616 , \18318_18617 , \18319_18618 , \18320_18619 , \18321_18620 , \18322_18621 , \18323_18622 , \18324_18623 , \18325_18624 , \18326_18625 , \18327_18626 , \18328_18627 , \18329_18628 , \18330_18629 , \18331_18630 , \18332_18631 , \18333_18632 , \18334_18633 , \18335_18634 , \18336_18635 , \18337_18636 , \18338_18637 , \18339_18638 , \18340_18639 , \18341_18640 , \18342_18641 , \18343_18642 , \18344_18643 , \18345_18644 , \18346_18645 , \18347_18646 , \18348_18647 , \18349_18648 , \18350_18649 , \18351_18650 , \18352_18651 , \18353_18652 , \18354_18653 , \18355_18654 , \18356_18655 , \18357_18656 , \18358_18657 , \18359_18658 , \18360_18659 , \18361_18660 , \18362_18661 , \18363_18662 , \18364_18663 , \18365_18664 , \18366_18665 , \18367_18666 , \18368_18667 , \18369_18668 , \18370_18669 , \18371_18670 , \18372_18671 , \18373_18672 , \18374_18673 , \18375_18674 , \18376_18675 , \18377_18676 , \18378_18677 , \18379_18678 , \18380_18679 );
or \U$9553 ( \18382_18681 , \18316_18615 , \18381_18680 );
_DC \g3c37/U$1 ( \18383 , \18382_18681 , \9298_9597 );
buf \U$9554 ( \18384_18683 , \18383 );
and \U$9555 ( \18385_18684 , \18251_18550 , \18384_18683 );
and \U$9556 ( \18386_18685 , \16579_16878 , \16712_17011 );
and \U$9557 ( \18387_18686 , \16712_17011 , \16987_17286 );
and \U$9558 ( \18388_18687 , \16579_16878 , \16987_17286 );
or \U$9559 ( \18389_18688 , \18386_18685 , \18387_18686 , \18388_18687 );
and \U$9560 ( \18390_18689 , \18384_18683 , \18389_18688 );
and \U$9561 ( \18391_18690 , \18251_18550 , \18389_18688 );
or \U$9562 ( \18392_18691 , \18385_18684 , \18390_18689 , \18391_18690 );
xor \U$9563 ( \18393_18692 , \18118_18417 , \18392_18691 );
buf g442a_GF_PartitionCandidate( \18394_18693_nG442a , \18393_18692 );
xor \U$9564 ( \18395_18694 , \18251_18550 , \18384_18683 );
xor \U$9565 ( \18396_18695 , \18395_18694 , \18389_18688 );
buf g442d_GF_PartitionCandidate( \18397_18696_nG442d , \18396_18695 );
nand \U$9566 ( \18398_18697 , \18397_18696_nG442d , \16989_17288_nG4430 );
and \U$9567 ( \18399_18698 , \18394_18693_nG442a , \18398_18697 );
xor \U$9568 ( \18400_18699 , \18397_18696_nG442d , \16989_17288_nG4430 );
and \U$9573 ( \18401_18703 , \18400_18699 , \10392_10694_nG9c0e );
or \U$9574 ( \18402_18704 , 1'b0 , \18401_18703 );
xor \U$9575 ( \18403_18705 , \18399_18698 , \18402_18704 );
xor \U$9576 ( \18404_18706 , \18399_18698 , \18403_18705 );
buf \U$9577 ( \18405_18707 , \18404_18706 );
buf \U$9578 ( \18406_18708 , \18405_18707 );
and \U$9579 ( \18407_18709 , \17851_18150 , \18406_18708 );
and \U$9580 ( \18408_18710 , \17838_18137 , \17843_18142 );
and \U$9581 ( \18409_18711 , \17838_18137 , \17849_18148 );
and \U$9582 ( \18410_18712 , \17843_18142 , \17849_18148 );
or \U$9583 ( \18411_18713 , \18408_18710 , \18409_18711 , \18410_18712 );
buf \U$9584 ( \18412_18714 , \18411_18713 );
and \U$9585 ( \18413_18715 , \17423_17725 , \17463_17762 );
and \U$9586 ( \18414_18716 , \17423_17725 , \17813_18112 );
and \U$9587 ( \18415_18717 , \17463_17762 , \17813_18112 );
or \U$9588 ( \18416_18718 , \18413_18715 , \18414_18716 , \18415_18717 );
buf \U$9589 ( \18417_18719 , \18416_18718 );
and \U$9590 ( \18418_18720 , \17437_17297 , \10693_10995_nG9c0b );
and \U$9591 ( \18419_18721 , \16995_17294 , \10981_11283_nG9c08 );
or \U$9592 ( \18420_18722 , \18418_18720 , \18419_18721 );
xor \U$9593 ( \18421_18723 , \16994_17293 , \18420_18722 );
buf \U$9594 ( \18422_18724 , \18421_18723 );
buf \U$9596 ( \18423_18725 , \18422_18724 );
and \U$9597 ( \18424_18726 , \16405_15940 , \11299_11598_nG9c05 );
and \U$9598 ( \18425_18727 , \15638_15937 , \12168_12470_nG9c02 );
or \U$9599 ( \18426_18728 , \18424_18726 , \18425_18727 );
xor \U$9600 ( \18427_18729 , \15637_15936 , \18426_18728 );
buf \U$9601 ( \18428_18730 , \18427_18729 );
buf \U$9603 ( \18429_18731 , \18428_18730 );
xor \U$9604 ( \18430_18732 , \18423_18725 , \18429_18731 );
buf \U$9605 ( \18431_18733 , \18430_18732 );
and \U$9606 ( \18432_18734 , \17426_17728 , \17432_17734 );
buf \U$9607 ( \18433_18735 , \18432_18734 );
xor \U$9608 ( \18434_18736 , \18431_18733 , \18433_18735 );
and \U$9609 ( \18435_18737 , \14710_14631 , \12502_12801_nG9bff );
and \U$9610 ( \18436_18738 , \14329_14628 , \13403_13705_nG9bfc );
or \U$9611 ( \18437_18739 , \18435_18737 , \18436_18738 );
xor \U$9612 ( \18438_18740 , \14328_14627 , \18437_18739 );
buf \U$9613 ( \18439_18741 , \18438_18740 );
buf \U$9615 ( \18440_18742 , \18439_18741 );
xor \U$9616 ( \18441_18743 , \18434_18736 , \18440_18742 );
buf \U$9617 ( \18442_18744 , \18441_18743 );
and \U$9618 ( \18443_18745 , \10996_10421 , \16378_16680_nG9bed );
and \U$9619 ( \18444_18746 , \10119_10418 , \17363_17665_nG9bea );
or \U$9620 ( \18445_18747 , \18443_18745 , \18444_18746 );
xor \U$9621 ( \18446_18748 , \10118_10417 , \18445_18747 );
buf \U$9622 ( \18447_18749 , \18446_18748 );
buf \U$9624 ( \18448_18750 , \18447_18749 );
xor \U$9625 ( \18449_18751 , \18442_18744 , \18448_18750 );
and \U$9626 ( \18450_18752 , \10411_10707 , \17808_18107_nG9be7 );
and \U$9627 ( \18451_18753 , \17764_18063 , \17778_18077 );
and \U$9628 ( \18452_18754 , \17778_18077 , \17796_18095 );
and \U$9629 ( \18453_18755 , \17764_18063 , \17796_18095 );
or \U$9630 ( \18454_18756 , \18451_18753 , \18452_18754 , \18453_18755 );
and \U$9631 ( \18455_18757 , \17768_18067 , \17772_18071 );
and \U$9632 ( \18456_18758 , \17772_18071 , \17777_18076 );
and \U$9633 ( \18457_18759 , \17768_18067 , \17777_18076 );
or \U$9634 ( \18458_18760 , \18455_18757 , \18456_18758 , \18457_18759 );
and \U$9635 ( \18459_18761 , \17783_18082 , \17787_18086 );
and \U$9636 ( \18460_18762 , \17787_18086 , \17795_18094 );
and \U$9637 ( \18461_18763 , \17783_18082 , \17795_18094 );
or \U$9638 ( \18462_18764 , \18459_18761 , \18460_18762 , \18461_18763 );
xor \U$9639 ( \18463_18765 , \18458_18760 , \18462_18764 );
and \U$9640 ( \18464_18766 , \17736_18035 , \10681_10983 );
and \U$9641 ( \18465_18767 , RIdec4898_700, \9034_9333 );
and \U$9642 ( \18466_18768 , RIdec1b98_668, \9036_9335 );
and \U$9643 ( \18467_18769 , RIfc661d0_6184, \9038_9337 );
and \U$9644 ( \18468_18770 , RIdebee98_636, \9040_9339 );
and \U$9645 ( \18469_18771 , RIfce6b28_7647, \9042_9341 );
and \U$9646 ( \18470_18772 , RIdebc198_604, \9044_9343 );
and \U$9647 ( \18471_18773 , RIdeb9498_572, \9046_9345 );
and \U$9648 ( \18472_18774 , RIdeb6798_540, \9048_9347 );
and \U$9649 ( \18473_18775 , RIfc40d18_5763, \9050_9349 );
and \U$9650 ( \18474_18776 , RIdeb0d98_476, \9052_9351 );
and \U$9651 ( \18475_18777 , RIfcad648_6995, \9054_9353 );
and \U$9652 ( \18476_18778 , RIdeae098_444, \9056_9355 );
and \U$9653 ( \18477_18779 , RIfcaa510_6960, \9058_9357 );
and \U$9654 ( \18478_18780 , RIdea89e0_412, \9060_9359 );
and \U$9655 ( \18479_18781 , RIdea20e0_380, \9062_9361 );
and \U$9656 ( \18480_18782 , RIde9b7e0_348, \9064_9363 );
and \U$9657 ( \18481_18783 , RIfcab320_6970, \9066_9365 );
and \U$9658 ( \18482_18784 , RIfca8350_6936, \9068_9367 );
and \U$9659 ( \18483_18785 , RIfc6f6e0_6290, \9070_9369 );
and \U$9660 ( \18484_18786 , RIfcaa240_6958, \9072_9371 );
and \U$9661 ( \18485_18787 , RIde8fcd8_291, \9074_9373 );
and \U$9662 ( \18486_18788 , RIfe8aae0_7922, \9076_9375 );
and \U$9663 ( \18487_18789 , RIde88d48_257, \9078_9377 );
and \U$9664 ( \18488_18790 , RIde84860_236, \9080_9379 );
and \U$9665 ( \18489_18791 , RIde80a08_217, \9082_9381 );
and \U$9666 ( \18490_18792 , RIfc64718_6165, \9084_9383 );
and \U$9667 ( \18491_18793 , RIfcae020_7002, \9086_9385 );
and \U$9668 ( \18492_18794 , RIfcadeb8_7001, \9088_9387 );
and \U$9669 ( \18493_18795 , RIee38fe0_5107, \9090_9389 );
and \U$9670 ( \18494_18796 , RIe16add8_2593, \9092_9391 );
and \U$9671 ( \18495_18797 , RIe1695f0_2576, \9094_9393 );
and \U$9672 ( \18496_18798 , RIe167430_2552, \9096_9395 );
and \U$9673 ( \18497_18799 , RIe164898_2521, \9098_9397 );
and \U$9674 ( \18498_18800 , RIe161b98_2489, \9100_9399 );
and \U$9675 ( \18499_18801 , RIfe8a3d8_7917, \9102_9401 );
and \U$9676 ( \18500_18802 , RIe15ee98_2457, \9104_9403 );
and \U$9677 ( \18501_18803 , RIfe8a270_7916, \9106_9405 );
and \U$9678 ( \18502_18804 , RIe15c198_2425, \9108_9407 );
and \U$9679 ( \18503_18805 , RIe156798_2361, \9110_9409 );
and \U$9680 ( \18504_18806 , RIe153a98_2329, \9112_9411 );
and \U$9681 ( \18505_18807 , RIfc3f0f8_5743, \9114_9413 );
and \U$9682 ( \18506_18808 , RIe150d98_2297, \9116_9415 );
and \U$9683 ( \18507_18809 , RIfcab050_6968, \9118_9417 );
and \U$9684 ( \18508_18810 , RIe14e098_2265, \9120_9419 );
and \U$9685 ( \18509_18811 , RIfcca658_7325, \9122_9421 );
and \U$9686 ( \18510_18812 , RIe14b398_2233, \9124_9423 );
and \U$9687 ( \18511_18813 , RIe148698_2201, \9126_9425 );
and \U$9688 ( \18512_18814 , RIe145998_2169, \9128_9427 );
and \U$9689 ( \18513_18815 , RIfe8a810_7920, \9130_9429 );
and \U$9690 ( \18514_18816 , RIfe8a6a8_7919, \9132_9431 );
and \U$9691 ( \18515_18817 , RIee31b28_5024, \9134_9433 );
and \U$9692 ( \18516_18818 , RIee30e80_5015, \9136_9435 );
and \U$9693 ( \18517_18819 , RIe140808_2111, \9138_9437 );
and \U$9694 ( \18518_18820 , RIfe8a540_7918, \9140_9439 );
and \U$9695 ( \18519_18821 , RIdf3c3e8_2062, \9142_9441 );
and \U$9696 ( \18520_18822 , RIdf3a0c0_2037, \9144_9443 );
and \U$9697 ( \18521_18823 , RIfc6b1f8_6241, \9146_9445 );
and \U$9698 ( \18522_18824 , RIee2f260_4995, \9148_9447 );
and \U$9699 ( \18523_18825 , RIfc70d60_6306, \9150_9449 );
and \U$9700 ( \18524_18826 , RIee2d0a0_4971, \9152_9451 );
and \U$9701 ( \18525_18827 , RIfe8a978_7921, \9154_9453 );
and \U$9702 ( \18526_18828 , RIdf32c08_1954, \9156_9455 );
and \U$9703 ( \18527_18829 , RIdf308e0_1929, \9158_9457 );
and \U$9704 ( \18528_18830 , RIdf2e9f0_1907, \9160_9459 );
or \U$9705 ( \18529_18831 , \18465_18767 , \18466_18768 , \18467_18769 , \18468_18770 , \18469_18771 , \18470_18772 , \18471_18773 , \18472_18774 , \18473_18775 , \18474_18776 , \18475_18777 , \18476_18778 , \18477_18779 , \18478_18780 , \18479_18781 , \18480_18782 , \18481_18783 , \18482_18784 , \18483_18785 , \18484_18786 , \18485_18787 , \18486_18788 , \18487_18789 , \18488_18790 , \18489_18791 , \18490_18792 , \18491_18793 , \18492_18794 , \18493_18795 , \18494_18796 , \18495_18797 , \18496_18798 , \18497_18799 , \18498_18800 , \18499_18801 , \18500_18802 , \18501_18803 , \18502_18804 , \18503_18805 , \18504_18806 , \18505_18807 , \18506_18808 , \18507_18809 , \18508_18810 , \18509_18811 , \18510_18812 , \18511_18813 , \18512_18814 , \18513_18815 , \18514_18816 , \18515_18817 , \18516_18818 , \18517_18819 , \18518_18820 , \18519_18821 , \18520_18822 , \18521_18823 , \18522_18824 , \18523_18825 , \18524_18826 , \18525_18827 , \18526_18828 , \18527_18829 , \18528_18830 );
and \U$9706 ( \18530_18832 , RIee2b5e8_4952, \9163_9462 );
and \U$9707 ( \18531_18833 , RIee29e00_4935, \9165_9464 );
and \U$9708 ( \18532_18834 , RIee28a50_4921, \9167_9466 );
and \U$9709 ( \18533_18835 , RIee276a0_4907, \9169_9468 );
and \U$9710 ( \18534_18836 , RIdf29c98_1852, \9171_9470 );
and \U$9711 ( \18535_18837 , RIdf27970_1827, \9173_9472 );
and \U$9712 ( \18536_18838 , RIdf25be8_1806, \9175_9474 );
and \U$9713 ( \18537_18839 , RIdf23fc8_1786, \9177_9476 );
and \U$9714 ( \18538_18840 , RIfc6aaf0_6236, \9179_9478 );
and \U$9715 ( \18539_18841 , RIfc6ac58_6237, \9181_9480 );
and \U$9716 ( \18540_18842 , RIdf22678_1768, \9183_9482 );
and \U$9717 ( \18541_18843 , RIfcdd4b0_7540, \9185_9484 );
and \U$9718 ( \18542_18844 , RIdf21160_1753, \9187_9486 );
and \U$9719 ( \18543_18845 , RIdf1f108_1730, \9189_9488 );
and \U$9720 ( \18544_18846 , RIdf1ac20_1681, \9191_9490 );
and \U$9721 ( \18545_18847 , RIfeaa7f0_8256, \9193_9492 );
and \U$9722 ( \18546_18848 , RIdf16468_1630, \9195_9494 );
and \U$9723 ( \18547_18849 , RIdf13768_1598, \9197_9496 );
and \U$9724 ( \18548_18850 , RIdf10a68_1566, \9199_9498 );
and \U$9725 ( \18549_18851 , RIdf0dd68_1534, \9201_9500 );
and \U$9726 ( \18550_18852 , RIdf0b068_1502, \9203_9502 );
and \U$9727 ( \18551_18853 , RIdf08368_1470, \9205_9504 );
and \U$9728 ( \18552_18854 , RIdf05668_1438, \9207_9506 );
and \U$9729 ( \18553_18855 , RIdf02968_1406, \9209_9508 );
and \U$9730 ( \18554_18856 , RIdefcf68_1342, \9211_9510 );
and \U$9731 ( \18555_18857 , RIdefa268_1310, \9213_9512 );
and \U$9732 ( \18556_18858 , RIdef7568_1278, \9215_9514 );
and \U$9733 ( \18557_18859 , RIdef4868_1246, \9217_9516 );
and \U$9734 ( \18558_18860 , RIdef1b68_1214, \9219_9518 );
and \U$9735 ( \18559_18861 , RIdeeee68_1182, \9221_9520 );
and \U$9736 ( \18560_18862 , RIdeec168_1150, \9223_9522 );
and \U$9737 ( \18561_18863 , RIdee9468_1118, \9225_9524 );
and \U$9738 ( \18562_18864 , RIee25378_4882, \9227_9526 );
and \U$9739 ( \18563_18865 , RIee24568_4872, \9229_9528 );
and \U$9740 ( \18564_18866 , RIee23a28_4864, \9231_9530 );
and \U$9741 ( \18565_18867 , RIee23050_4857, \9233_9532 );
and \U$9742 ( \18566_18868 , RIfe8adb0_7924, \9235_9534 );
and \U$9743 ( \18567_18869 , RIdee23e8_1038, \9237_9536 );
and \U$9744 ( \18568_18870 , RIfe8ac48_7923, \9239_9538 );
and \U$9745 ( \18569_18871 , RIdede1d0_991, \9241_9540 );
and \U$9746 ( \18570_18872 , RIfca5650_6904, \9243_9542 );
and \U$9747 ( \18571_18873 , RIee220d8_4846, \9245_9544 );
and \U$9748 ( \18572_18874 , RIfceeb20_7738, \9247_9546 );
and \U$9749 ( \18573_18875 , RIee20ff8_4834, \9249_9548 );
and \U$9750 ( \18574_18876 , RIded8ed8_932, \9251_9550 );
and \U$9751 ( \18575_18877 , RIfe8af18_7925, \9253_9552 );
and \U$9752 ( \18576_18878 , RIded49f0_883, \9255_9554 );
and \U$9753 ( \18577_18879 , RIfe8b080_7926, \9257_9556 );
and \U$9754 ( \18578_18880 , RIdecfc98_828, \9259_9558 );
and \U$9755 ( \18579_18881 , RIdeccf98_796, \9261_9560 );
and \U$9756 ( \18580_18882 , RIdeca298_764, \9263_9562 );
and \U$9757 ( \18581_18883 , RIdec7598_732, \9265_9564 );
and \U$9758 ( \18582_18884 , RIdeb3a98_508, \9267_9566 );
and \U$9759 ( \18583_18885 , RIde94ee0_316, \9269_9568 );
and \U$9760 ( \18584_18886 , RIe16d6a0_2622, \9271_9570 );
and \U$9761 ( \18585_18887 , RIe159498_2393, \9273_9572 );
and \U$9762 ( \18586_18888 , RIe142c98_2137, \9275_9574 );
and \U$9763 ( \18587_18889 , RIdf37690_2007, \9277_9576 );
and \U$9764 ( \18588_18890 , RIdf2bcf0_1875, \9279_9578 );
and \U$9765 ( \18589_18891 , RIdf1c570_1699, \9281_9580 );
and \U$9766 ( \18590_18892 , RIdeffc68_1374, \9283_9582 );
and \U$9767 ( \18591_18893 , RIdee6768_1086, \9285_9584 );
and \U$9768 ( \18592_18894 , RIdedb4d0_959, \9287_9586 );
and \U$9769 ( \18593_18895 , RIde7ae28_189, \9289_9588 );
or \U$9770 ( \18594_18896 , \18530_18832 , \18531_18833 , \18532_18834 , \18533_18835 , \18534_18836 , \18535_18837 , \18536_18838 , \18537_18839 , \18538_18840 , \18539_18841 , \18540_18842 , \18541_18843 , \18542_18844 , \18543_18845 , \18544_18846 , \18545_18847 , \18546_18848 , \18547_18849 , \18548_18850 , \18549_18851 , \18550_18852 , \18551_18853 , \18552_18854 , \18553_18855 , \18554_18856 , \18555_18857 , \18556_18858 , \18557_18859 , \18558_18860 , \18559_18861 , \18560_18862 , \18561_18863 , \18562_18864 , \18563_18865 , \18564_18866 , \18565_18867 , \18566_18868 , \18567_18869 , \18568_18870 , \18569_18871 , \18570_18872 , \18571_18873 , \18572_18874 , \18573_18875 , \18574_18876 , \18575_18877 , \18576_18878 , \18577_18879 , \18578_18880 , \18579_18881 , \18580_18882 , \18581_18883 , \18582_18884 , \18583_18885 , \18584_18886 , \18585_18887 , \18586_18888 , \18587_18889 , \18588_18890 , \18589_18891 , \18590_18892 , \18591_18893 , \18592_18894 , \18593_18895 );
or \U$9771 ( \18595_18897 , \18529_18831 , \18594_18896 );
_DC \g65a1/U$1 ( \18596 , \18595_18897 , \9298_9597 );
and \U$9772 ( \18597_18899 , RIe19cb30_3160, \8760_9059 );
and \U$9773 ( \18598_18900 , RIe199e30_3128, \8762_9061 );
and \U$9774 ( \18599_18901 , RIf145388_5247, \8764_9063 );
and \U$9775 ( \18600_18902 , RIe197130_3096, \8766_9065 );
and \U$9776 ( \18601_18903 , RIfe8a108_7915, \8768_9067 );
and \U$9777 ( \18602_18904 , RIe194430_3064, \8770_9069 );
and \U$9778 ( \18603_18905 , RIe191730_3032, \8772_9071 );
and \U$9779 ( \18604_18906 , RIe18ea30_3000, \8774_9073 );
and \U$9780 ( \18605_18907 , RIe189030_2936, \8776_9075 );
and \U$9781 ( \18606_18908 , RIe186330_2904, \8778_9077 );
and \U$9782 ( \18607_18909 , RIfc6c878_6257, \8780_9079 );
and \U$9783 ( \18608_18910 , RIe183630_2872, \8782_9081 );
and \U$9784 ( \18609_18911 , RIfcabcf8_6977, \8784_9083 );
and \U$9785 ( \18610_18912 , RIe180930_2840, \8786_9085 );
and \U$9786 ( \18611_18913 , RIe17dc30_2808, \8788_9087 );
and \U$9787 ( \18612_18914 , RIe17af30_2776, \8790_9089 );
and \U$9788 ( \18613_18915 , RIfcccc50_7352, \8792_9091 );
and \U$9789 ( \18614_18916 , RIfcccdb8_7353, \8794_9093 );
and \U$9790 ( \18615_18917 , RIe176d18_2729, \8796_9095 );
and \U$9791 ( \18616_18918 , RIfea7af0_8224, \8798_9097 );
and \U$9792 ( \18617_18919 , RIfe89fa0_7914, \8800_9099 );
and \U$9793 ( \18618_18920 , RIfe89e38_7913, \8802_9101 );
and \U$9794 ( \18619_18921 , RIfcdd078_7537, \8804_9103 );
and \U$9795 ( \18620_18922 , RIfccb738_7337, \8806_9105 );
and \U$9796 ( \18621_18923 , RIfca9868_6951, \8808_9107 );
and \U$9797 ( \18622_18924 , RIfcabb90_6976, \8810_9109 );
and \U$9798 ( \18623_18925 , RIfca99d0_6952, \8812_9111 );
and \U$9799 ( \18624_18926 , RIe172f38_2685, \8814_9113 );
and \U$9800 ( \18625_18927 , RIf16fd90_5732, \8816_9115 );
and \U$9801 ( \18626_18928 , RIf16f250_5724, \8818_9117 );
and \U$9802 ( \18627_18929 , RIfc6c440_6254, \8820_9119 );
and \U$9803 ( \18628_18930 , RIfcaba28_6975, \8822_9121 );
and \U$9804 ( \18629_18931 , RIfc40610_5758, \8824_9123 );
and \U$9805 ( \18630_18932 , RIe222e88_4687, \8826_9125 );
and \U$9806 ( \18631_18933 , RIfc5d260_6082, \8828_9127 );
and \U$9807 ( \18632_18934 , RIe220188_4655, \8830_9129 );
and \U$9808 ( \18633_18935 , RIfcab758_6973, \8832_9131 );
and \U$9809 ( \18634_18936 , RIe21d488_4623, \8834_9133 );
and \U$9810 ( \18635_18937 , RIe217a88_4559, \8836_9135 );
and \U$9811 ( \18636_18938 , RIe214d88_4527, \8838_9137 );
and \U$9812 ( \18637_18939 , RIfe892f8_7905, \8840_9139 );
and \U$9813 ( \18638_18940 , RIe212088_4495, \8842_9141 );
and \U$9814 ( \18639_18941 , RIf168a40_5650, \8844_9143 );
and \U$9815 ( \18640_18942 , RIe20f388_4463, \8846_9145 );
and \U$9816 ( \18641_18943 , RIf167ac8_5639, \8848_9147 );
and \U$9817 ( \18642_18944 , RIe20c688_4431, \8850_9149 );
and \U$9818 ( \18643_18945 , RIe209988_4399, \8852_9151 );
and \U$9819 ( \18644_18946 , RIe206c88_4367, \8854_9153 );
and \U$9820 ( \18645_18947 , RIfc6c2d8_6253, \8856_9155 );
and \U$9821 ( \18646_18948 , RIfceec88_7739, \8858_9157 );
and \U$9822 ( \18647_18949 , RIe201f30_4312, \8860_9159 );
and \U$9823 ( \18648_18950 , RIe200748_4295, \8862_9161 );
and \U$9824 ( \18649_18951 , RIf164dc8_5607, \8864_9163 );
and \U$9825 ( \18650_18952 , RIf163fb8_5597, \8866_9165 );
and \U$9826 ( \18651_18953 , RIf163040_5586, \8868_9167 );
and \U$9827 ( \18652_18954 , RIfe895c8_7907, \8870_9169 );
and \U$9828 ( \18653_18955 , RIf15f968_5547, \8872_9171 );
and \U$9829 ( \18654_18956 , RIfe89898_7909, \8874_9173 );
and \U$9830 ( \18655_18957 , RIfe89460_7906, \8876_9175 );
and \U$9831 ( \18656_18958 , RIe1fb5b8_4237, \8878_9177 );
and \U$9832 ( \18657_18959 , RIf15c6c8_5511, \8880_9179 );
and \U$9833 ( \18658_18960 , RIfe89730_7908, \8882_9181 );
and \U$9834 ( \18659_18961 , RIf15a238_5485, \8884_9183 );
and \U$9835 ( \18660_18962 , RIf1599c8_5479, \8886_9185 );
or \U$9836 ( \18661_18963 , \18597_18899 , \18598_18900 , \18599_18901 , \18600_18902 , \18601_18903 , \18602_18904 , \18603_18905 , \18604_18906 , \18605_18907 , \18606_18908 , \18607_18909 , \18608_18910 , \18609_18911 , \18610_18912 , \18611_18913 , \18612_18914 , \18613_18915 , \18614_18916 , \18615_18917 , \18616_18918 , \18617_18919 , \18618_18920 , \18619_18921 , \18620_18922 , \18621_18923 , \18622_18924 , \18623_18925 , \18624_18926 , \18625_18927 , \18626_18928 , \18627_18929 , \18628_18930 , \18629_18931 , \18630_18932 , \18631_18933 , \18632_18934 , \18633_18935 , \18634_18936 , \18635_18937 , \18636_18938 , \18637_18939 , \18638_18940 , \18639_18941 , \18640_18942 , \18641_18943 , \18642_18944 , \18643_18945 , \18644_18946 , \18645_18947 , \18646_18948 , \18647_18949 , \18648_18950 , \18649_18951 , \18650_18952 , \18651_18953 , \18652_18954 , \18653_18955 , \18654_18956 , \18655_18957 , \18656_18958 , \18657_18959 , \18658_18960 , \18659_18961 , \18660_18962 );
and \U$9837 ( \18662_18964 , RIf1588e8_5467, \8889_9188 );
and \U$9838 ( \18663_18965 , RIfe89cd0_7912, \8891_9190 );
and \U$9839 ( \18664_18966 , RIfc5ba78_6065, \8893_9192 );
and \U$9840 ( \18665_18967 , RIe1f9c68_4219, \8895_9194 );
and \U$9841 ( \18666_18968 , RIfc5bd48_6067, \8897_9196 );
and \U$9842 ( \18667_18969 , RIf1554e0_5430, \8899_9198 );
and \U$9843 ( \18668_18970 , RIf154298_5417, \8901_9200 );
and \U$9844 ( \18669_18971 , RIe1f4c40_4162, \8903_9202 );
and \U$9845 ( \18670_18972 , RIfe89b68_7911, \8905_9204 );
and \U$9846 ( \18671_18973 , RIfe89a00_7910, \8907_9206 );
and \U$9847 ( \18672_18974 , RIf150350_5372, \8909_9208 );
and \U$9848 ( \18673_18975 , RIe1f2918_4137, \8911_9210 );
and \U$9849 ( \18674_18976 , RIf14f3d8_5361, \8913_9212 );
and \U$9850 ( \18675_18977 , RIfccc818_7349, \8915_9214 );
and \U$9851 ( \18676_18978 , RIf14d920_5342, \8917_9216 );
and \U$9852 ( \18677_18979 , RIe1ed620_4078, \8919_9218 );
and \U$9853 ( \18678_18980 , RIe1eabf0_4048, \8921_9220 );
and \U$9854 ( \18679_18981 , RIe1e7ef0_4016, \8923_9222 );
and \U$9855 ( \18680_18982 , RIe1e51f0_3984, \8925_9224 );
and \U$9856 ( \18681_18983 , RIe1e24f0_3952, \8927_9226 );
and \U$9857 ( \18682_18984 , RIe1df7f0_3920, \8929_9228 );
and \U$9858 ( \18683_18985 , RIe1dcaf0_3888, \8931_9230 );
and \U$9859 ( \18684_18986 , RIe1d9df0_3856, \8933_9232 );
and \U$9860 ( \18685_18987 , RIe1d70f0_3824, \8935_9234 );
and \U$9861 ( \18686_18988 , RIe1d16f0_3760, \8937_9236 );
and \U$9862 ( \18687_18989 , RIe1ce9f0_3728, \8939_9238 );
and \U$9863 ( \18688_18990 , RIe1cbcf0_3696, \8941_9240 );
and \U$9864 ( \18689_18991 , RIe1c8ff0_3664, \8943_9242 );
and \U$9865 ( \18690_18992 , RIe1c62f0_3632, \8945_9244 );
and \U$9866 ( \18691_18993 , RIe1c35f0_3600, \8947_9246 );
and \U$9867 ( \18692_18994 , RIe1c08f0_3568, \8949_9248 );
and \U$9868 ( \18693_18995 , RIe1bdbf0_3536, \8951_9250 );
and \U$9869 ( \18694_18996 , RIfc680c0_6206, \8953_9252 );
and \U$9870 ( \18695_18997 , RIf14b058_5313, \8955_9254 );
and \U$9871 ( \18696_18998 , RIe1b8bc8_3479, \8957_9256 );
and \U$9872 ( \18697_18999 , RIe1b6b70_3456, \8959_9258 );
and \U$9873 ( \18698_19000 , RIfcac298_6981, \8961_9260 );
and \U$9874 ( \18699_19001 , RIf1499d8_5297, \8963_9262 );
and \U$9875 ( \18700_19002 , RIfe89190_7904, \8965_9264 );
and \U$9876 ( \18701_19003 , RIfec19c8_8323, \8967_9266 );
and \U$9877 ( \18702_19004 , RIf148a60_5286, \8969_9268 );
and \U$9878 ( \18703_19005 , RIfccdd30_7364, \8971_9270 );
and \U$9879 ( \18704_19006 , RIe1b2250_3404, \8973_9272 );
and \U$9880 ( \18705_19007 , RIfec1860_8322, \8975_9274 );
and \U$9881 ( \18706_19008 , RIfc6e768_6279, \8977_9276 );
and \U$9882 ( \18707_19009 , RIfc54728_5983, \8979_9278 );
and \U$9883 ( \18708_19010 , RIe1abfe0_3334, \8981_9280 );
and \U$9884 ( \18709_19011 , RIe1aa528_3315, \8983_9282 );
and \U$9885 ( \18710_19012 , RIe1a7f30_3288, \8985_9284 );
and \U$9886 ( \18711_19013 , RIe1a5230_3256, \8987_9286 );
and \U$9887 ( \18712_19014 , RIe1a2530_3224, \8989_9288 );
and \U$9888 ( \18713_19015 , RIe19f830_3192, \8991_9290 );
and \U$9889 ( \18714_19016 , RIe18bd30_2968, \8993_9292 );
and \U$9890 ( \18715_19017 , RIe178230_2744, \8995_9294 );
and \U$9891 ( \18716_19018 , RIe225b88_4719, \8997_9296 );
and \U$9892 ( \18717_19019 , RIe21a788_4591, \8999_9298 );
and \U$9893 ( \18718_19020 , RIe203f88_4335, \9001_9300 );
and \U$9894 ( \18719_19021 , RIe1fdfe8_4267, \9003_9302 );
and \U$9895 ( \18720_19022 , RIe1f73a0_4190, \9005_9304 );
and \U$9896 ( \18721_19023 , RIe1efee8_4107, \9007_9306 );
and \U$9897 ( \18722_19024 , RIe1d43f0_3792, \9009_9308 );
and \U$9898 ( \18723_19025 , RIe1baef0_3504, \9011_9310 );
and \U$9899 ( \18724_19026 , RIe1add68_3355, \9013_9312 );
and \U$9900 ( \18725_19027 , RIe1703a0_2654, \9015_9314 );
or \U$9901 ( \18726_19028 , \18662_18964 , \18663_18965 , \18664_18966 , \18665_18967 , \18666_18968 , \18667_18969 , \18668_18970 , \18669_18971 , \18670_18972 , \18671_18973 , \18672_18974 , \18673_18975 , \18674_18976 , \18675_18977 , \18676_18978 , \18677_18979 , \18678_18980 , \18679_18981 , \18680_18982 , \18681_18983 , \18682_18984 , \18683_18985 , \18684_18986 , \18685_18987 , \18686_18988 , \18687_18989 , \18688_18990 , \18689_18991 , \18690_18992 , \18691_18993 , \18692_18994 , \18693_18995 , \18694_18996 , \18695_18997 , \18696_18998 , \18697_18999 , \18698_19000 , \18699_19001 , \18700_19002 , \18701_19003 , \18702_19004 , \18703_19005 , \18704_19006 , \18705_19007 , \18706_19008 , \18707_19009 , \18708_19010 , \18709_19011 , \18710_19012 , \18711_19013 , \18712_19014 , \18713_19015 , \18714_19016 , \18715_19017 , \18716_19018 , \18717_19019 , \18718_19020 , \18719_19021 , \18720_19022 , \18721_19023 , \18722_19024 , \18723_19025 , \18724_19026 , \18725_19027 );
or \U$9902 ( \18727_19029 , \18661_18963 , \18726_19028 );
_DC \g65a2/U$1 ( \18728 , \18727_19029 , \9024_9323 );
and g65a3_GF_PartitionCandidate( \18729_19031_nG65a3 , \18596 , \18728 );
buf \U$9903 ( \18730_19032 , \18729_19031_nG65a3 );
and \U$9904 ( \18731_19033 , \18730_19032 , \10389_10691 );
nor \U$9905 ( \18732_19034 , \18464_18766 , \18731_19033 );
xnor \U$9906 ( \18733_19035 , \18732_19034 , \10678_10980 );
and \U$9907 ( \18734_19036 , \16353_16655 , \11275_11574 );
and \U$9908 ( \18735_19037 , \17325_17627 , \10976_11278 );
nor \U$9909 ( \18736_19038 , \18734_19036 , \18735_19037 );
xnor \U$9910 ( \18737_19039 , \18736_19038 , \11281_11580 );
xor \U$9911 ( \18738_19040 , \18733_19035 , \18737_19039 );
_DC \g5358/U$1 ( \18739 , \18595_18897 , \9298_9597 );
_DC \g53dc/U$1 ( \18740 , \18727_19029 , \9024_9323 );
xor g53dd_GF_PartitionCandidate( \18741_19043_nG53dd , \18739 , \18740 );
buf \U$9912 ( \18742_19044 , \18741_19043_nG53dd );
xor \U$9913 ( \18743_19045 , \18742_19044 , \17744_18043 );
and \U$9914 ( \18744_19046 , \10385_10687 , \18743_19045 );
xor \U$9915 ( \18745_19047 , \18738_19040 , \18744_19046 );
xor \U$9916 ( \18746_19048 , \18463_18765 , \18745_19047 );
xor \U$9917 ( \18747_19049 , \18454_18756 , \18746_19048 );
and \U$9918 ( \18748_19050 , \17749_18048 , \17753_18052 );
and \U$9919 ( \18749_19051 , \17753_18052 , \17758_18057 );
and \U$9920 ( \18750_19052 , \17749_18048 , \17758_18057 );
or \U$9921 ( \18751_19053 , \18748_19050 , \18749_19051 , \18750_19052 );
and \U$9922 ( \18752_19054 , \15022_15321 , \12491_12790 );
and \U$9923 ( \18753_19055 , \15965_16267 , \12159_12461 );
nor \U$9924 ( \18754_19056 , \18752_19054 , \18753_19055 );
xnor \U$9925 ( \18755_19057 , \18754_19056 , \12481_12780 );
and \U$9926 ( \18756_19058 , \13725_14024 , \13755_14054 );
and \U$9927 ( \18757_19059 , \14648_14950 , \13390_13692 );
nor \U$9928 ( \18758_19060 , \18756_19058 , \18757_19059 );
xnor \U$9929 ( \18759_19061 , \18758_19060 , \13736_14035 );
xor \U$9930 ( \18760_19062 , \18755_19057 , \18759_19061 );
and \U$9931 ( \18761_19063 , \12470_12769 , \15037_15336 );
and \U$9932 ( \18762_19064 , \13377_13679 , \14661_14963 );
nor \U$9933 ( \18763_19065 , \18761_19063 , \18762_19064 );
xnor \U$9934 ( \18764_19066 , \18763_19065 , \15043_15342 );
xor \U$9935 ( \18765_19067 , \18760_19062 , \18764_19066 );
xor \U$9936 ( \18766_19068 , \18751_19053 , \18765_19067 );
and \U$9937 ( \18767_19069 , \17739_18038 , \17748_18047 );
and \U$9938 ( \18768_19070 , \11287_11586 , \16333_16635 );
and \U$9939 ( \18769_19071 , \12146_12448 , \15999_16301 );
nor \U$9940 ( \18770_19072 , \18768_19070 , \18769_19071 );
xnor \U$9941 ( \18771_19073 , \18770_19072 , \16323_16625 );
xor \U$9942 ( \18772_19074 , \18767_19069 , \18771_19073 );
and \U$9943 ( \18773_19075 , \10686_10988 , \17791_18090 );
and \U$9944 ( \18774_19076 , \10968_11270 , \17353_17655 );
nor \U$9945 ( \18775_19077 , \18773_19075 , \18774_19076 );
xnor \U$9946 ( \18776_19078 , \18775_19077 , \17747_18046 );
xor \U$9947 ( \18777_19079 , \18772_19074 , \18776_19078 );
xor \U$9948 ( \18778_19080 , \18766_19068 , \18777_19079 );
xor \U$9949 ( \18779_19081 , \18747_19049 , \18778_19080 );
and \U$9950 ( \18780_19082 , \17469_17768 , \17759_18058 );
and \U$9951 ( \18781_19083 , \17759_18058 , \17797_18096 );
and \U$9952 ( \18782_19084 , \17469_17768 , \17797_18096 );
or \U$9953 ( \18783_19085 , \18780_19082 , \18781_19083 , \18782_19084 );
xor \U$9954 ( \18784_19086 , \18779_19081 , \18783_19085 );
and \U$9955 ( \18785_19087 , \17798_18097 , \17802_18101 );
and \U$9956 ( \18786_19088 , \17803_18102 , \17806_18105 );
or \U$9957 ( \18787_19089 , \18785_19087 , \18786_19088 );
xor \U$9958 ( \18788_19090 , \18784_19086 , \18787_19089 );
buf g9be4_GF_PartitionCandidate( \18789_19091_nG9be4 , \18788_19090 );
and \U$9959 ( \18790_19092 , \10402_10704 , \18789_19091_nG9be4 );
or \U$9960 ( \18791_19093 , \18450_18752 , \18790_19092 );
xor \U$9961 ( \18792_19094 , \10399_10703 , \18791_19093 );
buf \U$9962 ( \18793_19095 , \18792_19094 );
buf \U$9964 ( \18794_19096 , \18793_19095 );
xor \U$9965 ( \18795_19097 , \18449_18751 , \18794_19096 );
buf \U$9966 ( \18796_19098 , \18795_19097 );
xor \U$9967 ( \18797_19099 , \18417_18719 , \18796_19098 );
and \U$9968 ( \18798_19100 , \17821_18120 , \17827_18126 );
and \U$9969 ( \18799_19101 , \17821_18120 , \17834_18133 );
and \U$9970 ( \18800_19102 , \17827_18126 , \17834_18133 );
or \U$9971 ( \18801_19103 , \18798_19100 , \18799_19101 , \18800_19102 );
buf \U$9972 ( \18802_19104 , \18801_19103 );
and \U$9973 ( \18803_19105 , \17434_17736 , \17443_17742 );
and \U$9974 ( \18804_19106 , \17434_17736 , \17450_17749 );
and \U$9975 ( \18805_19107 , \17443_17742 , \17450_17749 );
or \U$9976 ( \18806_19108 , \18803_19105 , \18804_19106 , \18805_19107 );
buf \U$9977 ( \18807_19109 , \18806_19108 );
and \U$9978 ( \18808_19110 , \13431_13370 , \13771_14070_nG9bf9 );
and \U$9979 ( \18809_19111 , \13068_13367 , \14682_14984_nG9bf6 );
or \U$9980 ( \18810_19112 , \18808_19110 , \18809_19111 );
xor \U$9981 ( \18811_19113 , \13067_13366 , \18810_19112 );
buf \U$9982 ( \18812_19114 , \18811_19113 );
buf \U$9984 ( \18813_19115 , \18812_19114 );
xor \U$9985 ( \18814_19116 , \18807_19109 , \18813_19115 );
and \U$9986 ( \18815_19117 , \12183_12157 , \15074_15373_nG9bf3 );
and \U$9987 ( \18816_19118 , \11855_12154 , \16013_16315_nG9bf0 );
or \U$9988 ( \18817_19119 , \18815_19117 , \18816_19118 );
xor \U$9989 ( \18818_19120 , \11854_12153 , \18817_19119 );
buf \U$9990 ( \18819_19121 , \18818_19120 );
buf \U$9992 ( \18820_19122 , \18819_19121 );
xor \U$9993 ( \18821_19123 , \18814_19116 , \18820_19122 );
buf \U$9994 ( \18822_19124 , \18821_19123 );
xor \U$9995 ( \18823_19125 , \18802_19104 , \18822_19124 );
and \U$9996 ( \18824_19126 , \17452_17751 , \17454_17753 );
and \U$9997 ( \18825_19127 , \17452_17751 , \17461_17760 );
and \U$9998 ( \18826_19128 , \17454_17753 , \17461_17760 );
or \U$9999 ( \18827_19129 , \18824_19126 , \18825_19127 , \18826_19128 );
buf \U$10000 ( \18828_19130 , \18827_19129 );
xor \U$10001 ( \18829_19131 , \18823_19125 , \18828_19130 );
buf \U$10002 ( \18830_19132 , \18829_19131 );
xor \U$10003 ( \18831_19133 , \18797_19099 , \18830_19132 );
buf \U$10004 ( \18832_19134 , \18831_19133 );
xor \U$10005 ( \18833_19135 , \18412_18714 , \18832_19134 );
and \U$10006 ( \18834_19136 , \17418_17720 , \17815_18114 );
and \U$10007 ( \18835_19137 , \17418_17720 , \17836_18135 );
and \U$10008 ( \18836_19138 , \17815_18114 , \17836_18135 );
or \U$10009 ( \18837_19139 , \18834_19136 , \18835_19137 , \18836_19138 );
buf \U$10010 ( \18838_19140 , \18837_19139 );
xor \U$10011 ( \18839_19141 , \18833_19135 , \18838_19140 );
and \U$10012 ( \18840_19142 , \17851_18150 , \18839_19141 );
and \U$10013 ( \18841_19143 , \18406_18708 , \18839_19141 );
or \U$10014 ( \18842_19144 , \18407_18709 , \18840_19142 , \18841_19143 );
and \U$10015 ( \18843_19145 , \18412_18714 , \18832_19134 );
and \U$10016 ( \18844_19146 , \18412_18714 , \18838_19140 );
and \U$10017 ( \18845_19147 , \18832_19134 , \18838_19140 );
or \U$10018 ( \18846_19148 , \18843_19145 , \18844_19146 , \18845_19147 );
buf \U$10019 ( \18847_19149 , \18846_19148 );
and \U$10020 ( \18848_19150 , \18802_19104 , \18822_19124 );
and \U$10021 ( \18849_19151 , \18802_19104 , \18828_19130 );
and \U$10022 ( \18850_19152 , \18822_19124 , \18828_19130 );
or \U$10023 ( \18851_19153 , \18848_19150 , \18849_19151 , \18850_19152 );
buf \U$10024 ( \18852_19154 , \18851_19153 );
and \U$10025 ( \18853_19155 , \18807_19109 , \18813_19115 );
and \U$10026 ( \18854_19156 , \18807_19109 , \18820_19122 );
and \U$10027 ( \18855_19157 , \18813_19115 , \18820_19122 );
or \U$10028 ( \18856_19158 , \18853_19155 , \18854_19156 , \18855_19157 );
buf \U$10029 ( \18857_19159 , \18856_19158 );
and \U$10030 ( \18858_19160 , \18423_18725 , \18429_18731 );
buf \U$10031 ( \18859_19161 , \18858_19160 );
and \U$10032 ( \18860_19162 , \14710_14631 , \13403_13705_nG9bfc );
and \U$10033 ( \18861_19163 , \14329_14628 , \13771_14070_nG9bf9 );
or \U$10034 ( \18862_19164 , \18860_19162 , \18861_19163 );
xor \U$10035 ( \18863_19165 , \14328_14627 , \18862_19164 );
buf \U$10036 ( \18864_19166 , \18863_19165 );
buf \U$10038 ( \18865_19167 , \18864_19166 );
xor \U$10039 ( \18866_19168 , \18859_19161 , \18865_19167 );
and \U$10040 ( \18867_19169 , \13431_13370 , \14682_14984_nG9bf6 );
and \U$10041 ( \18868_19170 , \13068_13367 , \15074_15373_nG9bf3 );
or \U$10042 ( \18869_19171 , \18867_19169 , \18868_19170 );
xor \U$10043 ( \18870_19172 , \13067_13366 , \18869_19171 );
buf \U$10044 ( \18871_19173 , \18870_19172 );
buf \U$10046 ( \18872_19174 , \18871_19173 );
xor \U$10047 ( \18873_19175 , \18866_19168 , \18872_19174 );
buf \U$10048 ( \18874_19176 , \18873_19175 );
xor \U$10049 ( \18875_19177 , \18857_19159 , \18874_19176 );
and \U$10050 ( \18876_19178 , \10996_10421 , \17363_17665_nG9bea );
and \U$10051 ( \18877_19179 , \10119_10418 , \17808_18107_nG9be7 );
or \U$10052 ( \18878_19180 , \18876_19178 , \18877_19179 );
xor \U$10053 ( \18879_19181 , \10118_10417 , \18878_19180 );
buf \U$10054 ( \18880_19182 , \18879_19181 );
buf \U$10056 ( \18881_19183 , \18880_19182 );
xor \U$10057 ( \18882_19184 , \18875_19177 , \18881_19183 );
buf \U$10058 ( \18883_19185 , \18882_19184 );
xor \U$10059 ( \18884_19186 , \18852_19154 , \18883_19185 );
and \U$10060 ( \18885_19187 , \18442_18744 , \18448_18750 );
and \U$10061 ( \18886_19188 , \18442_18744 , \18794_19096 );
and \U$10062 ( \18887_19189 , \18448_18750 , \18794_19096 );
or \U$10063 ( \18888_19190 , \18885_19187 , \18886_19188 , \18887_19189 );
buf \U$10064 ( \18889_19191 , \18888_19190 );
and \U$10065 ( \18890_19192 , \18431_18733 , \18433_18735 );
and \U$10066 ( \18891_19193 , \18431_18733 , \18440_18742 );
and \U$10067 ( \18892_19194 , \18433_18735 , \18440_18742 );
or \U$10068 ( \18893_19195 , \18890_19192 , \18891_19193 , \18892_19194 );
buf \U$10069 ( \18894_19196 , \18893_19195 );
and \U$10070 ( \18895_19197 , \18399_18698 , \18403_18705 );
buf \U$10071 ( \18896_19198 , \18895_19197 );
buf \U$10073 ( \18897_19199 , \18896_19198 );
and \U$10074 ( \18898_19200 , \17437_17297 , \10981_11283_nG9c08 );
and \U$10075 ( \18899_19201 , \16995_17294 , \11299_11598_nG9c05 );
or \U$10076 ( \18900_19202 , \18898_19200 , \18899_19201 );
xor \U$10077 ( \18901_19203 , \16994_17293 , \18900_19202 );
buf \U$10078 ( \18902_19204 , \18901_19203 );
buf \U$10080 ( \18903_19205 , \18902_19204 );
xor \U$10081 ( \18904_19206 , \18897_19199 , \18903_19205 );
buf \U$10082 ( \18905_19207 , \18904_19206 );
not \U$9569 ( \18906_18700 , \18400_18699 );
xor \U$9570 ( \18907_18701 , \18394_18693_nG442a , \18397_18696_nG442d );
and \U$9571 ( \18908_18702 , \18906_18700 , \18907_18701 );
and \U$10083 ( \18909_19208 , \18908_18702 , \10392_10694_nG9c0e );
and \U$10084 ( \18910_19209 , \18400_18699 , \10693_10995_nG9c0b );
or \U$10085 ( \18911_19210 , \18909_19208 , \18910_19209 );
xor \U$10086 ( \18912_19211 , \18399_18698 , \18911_19210 );
buf \U$10087 ( \18913_19212 , \18912_19211 );
buf \U$10089 ( \18914_19213 , \18913_19212 );
xor \U$10090 ( \18915_19214 , \18905_19207 , \18914_19213 );
and \U$10091 ( \18916_19215 , \16405_15940 , \12168_12470_nG9c02 );
and \U$10092 ( \18917_19216 , \15638_15937 , \12502_12801_nG9bff );
or \U$10093 ( \18918_19217 , \18916_19215 , \18917_19216 );
xor \U$10094 ( \18919_19218 , \15637_15936 , \18918_19217 );
buf \U$10095 ( \18920_19219 , \18919_19218 );
buf \U$10097 ( \18921_19220 , \18920_19219 );
xor \U$10098 ( \18922_19221 , \18915_19214 , \18921_19220 );
buf \U$10099 ( \18923_19222 , \18922_19221 );
xor \U$10100 ( \18924_19223 , \18894_19196 , \18923_19222 );
and \U$10101 ( \18925_19224 , \12183_12157 , \16013_16315_nG9bf0 );
and \U$10102 ( \18926_19225 , \11855_12154 , \16378_16680_nG9bed );
or \U$10103 ( \18927_19226 , \18925_19224 , \18926_19225 );
xor \U$10104 ( \18928_19227 , \11854_12153 , \18927_19226 );
buf \U$10105 ( \18929_19228 , \18928_19227 );
buf \U$10107 ( \18930_19229 , \18929_19228 );
xor \U$10108 ( \18931_19230 , \18924_19223 , \18930_19229 );
buf \U$10109 ( \18932_19231 , \18931_19230 );
xor \U$10110 ( \18933_19232 , \18889_19191 , \18932_19231 );
and \U$10111 ( \18934_19233 , \10411_10707 , \18789_19091_nG9be4 );
and \U$10112 ( \18935_19234 , \18751_19053 , \18765_19067 );
and \U$10113 ( \18936_19235 , \18765_19067 , \18777_19079 );
and \U$10114 ( \18937_19236 , \18751_19053 , \18777_19079 );
or \U$10115 ( \18938_19237 , \18935_19234 , \18936_19235 , \18937_19236 );
and \U$10116 ( \18939_19238 , \18755_19057 , \18759_19061 );
and \U$10117 ( \18940_19239 , \18759_19061 , \18764_19066 );
and \U$10118 ( \18941_19240 , \18755_19057 , \18764_19066 );
or \U$10119 ( \18942_19241 , \18939_19238 , \18940_19239 , \18941_19240 );
and \U$10120 ( \18943_19242 , \15965_16267 , \12491_12790 );
and \U$10121 ( \18944_19243 , \16353_16655 , \12159_12461 );
nor \U$10122 ( \18945_19244 , \18943_19242 , \18944_19243 );
xnor \U$10123 ( \18946_19245 , \18945_19244 , \12481_12780 );
and \U$10124 ( \18947_19246 , \13377_13679 , \15037_15336 );
and \U$10125 ( \18948_19247 , \13725_14024 , \14661_14963 );
nor \U$10126 ( \18949_19248 , \18947_19246 , \18948_19247 );
xnor \U$10127 ( \18950_19249 , \18949_19248 , \15043_15342 );
xor \U$10128 ( \18951_19250 , \18946_19245 , \18950_19249 );
and \U$10129 ( \18952_19251 , \12146_12448 , \16333_16635 );
and \U$10130 ( \18953_19252 , \12470_12769 , \15999_16301 );
nor \U$10131 ( \18954_19253 , \18952_19251 , \18953_19252 );
xnor \U$10132 ( \18955_19254 , \18954_19253 , \16323_16625 );
xor \U$10133 ( \18956_19255 , \18951_19250 , \18955_19254 );
xor \U$10134 ( \18957_19256 , \18942_19241 , \18956_19255 );
and \U$10135 ( \18958_19257 , \17325_17627 , \11275_11574 );
and \U$10136 ( \18959_19258 , \17736_18035 , \10976_11278 );
nor \U$10137 ( \18960_19259 , \18958_19257 , \18959_19258 );
xnor \U$10138 ( \18961_19260 , \18960_19259 , \11281_11580 );
and \U$10139 ( \18962_19261 , \14648_14950 , \13755_14054 );
and \U$10140 ( \18963_19262 , \15022_15321 , \13390_13692 );
nor \U$10141 ( \18964_19263 , \18962_19261 , \18963_19262 );
xnor \U$10142 ( \18965_19264 , \18964_19263 , \13736_14035 );
xor \U$10143 ( \18966_19265 , \18961_19260 , \18965_19264 );
and \U$10144 ( \18967_19266 , RIdec4a00_701, \9034_9333 );
and \U$10145 ( \18968_19267 , RIdec1d00_669, \9036_9335 );
and \U$10146 ( \18969_19268 , RIfcad7b0_6996, \9038_9337 );
and \U$10147 ( \18970_19269 , RIdebf000_637, \9040_9339 );
and \U$10148 ( \18971_19270 , RIfc64cb8_6169, \9042_9341 );
and \U$10149 ( \18972_19271 , RIdebc300_605, \9044_9343 );
and \U$10150 ( \18973_19272 , RIdeb9600_573, \9046_9345 );
and \U$10151 ( \18974_19273 , RIdeb6900_541, \9048_9347 );
and \U$10152 ( \18975_19274 , RIfc6f9b0_6292, \9050_9349 );
and \U$10153 ( \18976_19275 , RIdeb0f00_477, \9052_9351 );
and \U$10154 ( \18977_19276 , RIfc657f8_6177, \9054_9353 );
and \U$10155 ( \18978_19277 , RIdeae200_445, \9056_9355 );
and \U$10156 ( \18979_19278 , RIfce69c0_7646, \9058_9357 );
and \U$10157 ( \18980_19279 , RIdea8d28_413, \9060_9359 );
and \U$10158 ( \18981_19280 , RIdea2428_381, \9062_9361 );
and \U$10159 ( \18982_19281 , RIde9bb28_349, \9064_9363 );
and \U$10160 ( \18983_19282 , RIfc6fc80_6294, \9066_9365 );
and \U$10161 ( \18984_19283 , RIee1b760_4771, \9068_9367 );
and \U$10162 ( \18985_19284 , RIfca8080_6934, \9070_9369 );
and \U$10163 ( \18986_19285 , RIfe8b8f0_7932, \9072_9371 );
and \U$10164 ( \18987_19286 , RIde90020_292, \9074_9373 );
and \U$10165 ( \18988_19287 , RIde8c510_274, \9076_9375 );
and \U$10166 ( \18989_19288 , RIde89090_258, \9078_9377 );
and \U$10167 ( \18990_19289 , RIde84ba8_237, \9080_9379 );
and \U$10168 ( \18991_19290 , RIfc65ac8_6179, \9082_9381 );
and \U$10169 ( \18992_19291 , RIfcad210_6992, \9084_9383 );
and \U$10170 ( \18993_19292 , RIfcce168_7367, \9086_9385 );
and \U$10171 ( \18994_19293 , RIfcce2d0_7368, \9088_9387 );
and \U$10172 ( \18995_19294 , RIfc51488_5947, \9090_9389 );
and \U$10173 ( \18996_19295 , RIe16af40_2594, \9092_9391 );
and \U$10174 ( \18997_19296 , RIfc65c30_6180, \9094_9393 );
and \U$10175 ( \18998_19297 , RIe167598_2553, \9096_9395 );
and \U$10176 ( \18999_19298 , RIe164a00_2522, \9098_9397 );
and \U$10177 ( \19000_19299 , RIe161d00_2490, \9100_9399 );
and \U$10178 ( \19001_19300 , RIfc66e78_6193, \9102_9401 );
and \U$10179 ( \19002_19301 , RIe15f000_2458, \9104_9403 );
and \U$10180 ( \19003_19302 , RIfc6e498_6277, \9106_9405 );
and \U$10181 ( \19004_19303 , RIe15c300_2426, \9108_9407 );
and \U$10182 ( \19005_19304 , RIe156900_2362, \9110_9409 );
and \U$10183 ( \19006_19305 , RIe153c00_2330, \9112_9411 );
and \U$10184 ( \19007_19306 , RIfc6e330_6276, \9114_9413 );
and \U$10185 ( \19008_19307 , RIe150f00_2298, \9116_9415 );
and \U$10186 ( \19009_19308 , RIfccda60_7362, \9118_9417 );
and \U$10187 ( \19010_19309 , RIe14e200_2266, \9120_9419 );
and \U$10188 ( \19011_19310 , RIfc6e1c8_6275, \9122_9421 );
and \U$10189 ( \19012_19311 , RIe14b500_2234, \9124_9423 );
and \U$10190 ( \19013_19312 , RIe148800_2202, \9126_9425 );
and \U$10191 ( \19014_19313 , RIe145b00_2170, \9128_9427 );
and \U$10192 ( \19015_19314 , RIee33fb8_5050, \9130_9429 );
and \U$10193 ( \19016_19315 , RIee32d70_5037, \9132_9431 );
and \U$10194 ( \19017_19316 , RIee31c90_5025, \9134_9433 );
and \U$10195 ( \19018_19317 , RIee30fe8_5016, \9136_9435 );
and \U$10196 ( \19019_19318 , RIfea8630_8232, \9138_9437 );
and \U$10197 ( \19020_19319 , RIdf3e5a8_2086, \9140_9439 );
and \U$10198 ( \19021_19320 , RIdf3c550_2063, \9142_9441 );
and \U$10199 ( \19022_19321 , RIfea8798_8233, \9144_9443 );
and \U$10200 ( \19023_19322 , RIfc6e060_6274, \9146_9445 );
and \U$10201 ( \19024_19323 , RIfcac6d0_6984, \9148_9447 );
and \U$10202 ( \19025_19324 , RIfc56078_6001, \9150_9449 );
and \U$10203 ( \19026_19325 , RIfc6e600_6278, \9152_9451 );
and \U$10204 ( \19027_19326 , RIdf34dc8_1978, \9154_9453 );
and \U$10205 ( \19028_19327 , RIdf32d70_1955, \9156_9455 );
and \U$10206 ( \19029_19328 , RIfea84c8_8231, \9158_9457 );
and \U$10207 ( \19030_19329 , RIdf2eb58_1908, \9160_9459 );
or \U$10208 ( \19031_19330 , \18967_19266 , \18968_19267 , \18969_19268 , \18970_19269 , \18971_19270 , \18972_19271 , \18973_19272 , \18974_19273 , \18975_19274 , \18976_19275 , \18977_19276 , \18978_19277 , \18979_19278 , \18980_19279 , \18981_19280 , \18982_19281 , \18983_19282 , \18984_19283 , \18985_19284 , \18986_19285 , \18987_19286 , \18988_19287 , \18989_19288 , \18990_19289 , \18991_19290 , \18992_19291 , \18993_19292 , \18994_19293 , \18995_19294 , \18996_19295 , \18997_19296 , \18998_19297 , \18999_19298 , \19000_19299 , \19001_19300 , \19002_19301 , \19003_19302 , \19004_19303 , \19005_19304 , \19006_19305 , \19007_19306 , \19008_19307 , \19009_19308 , \19010_19309 , \19011_19310 , \19012_19311 , \19013_19312 , \19014_19313 , \19015_19314 , \19016_19315 , \19017_19316 , \19018_19317 , \19019_19318 , \19020_19319 , \19021_19320 , \19022_19321 , \19023_19322 , \19024_19323 , \19025_19324 , \19026_19325 , \19027_19326 , \19028_19327 , \19029_19328 , \19030_19329 );
and \U$10209 ( \19032_19331 , RIee2b750_4953, \9163_9462 );
and \U$10210 ( \19033_19332 , RIfc6ee70_6284, \9165_9464 );
and \U$10211 ( \19034_19333 , RIfc6efd8_6285, \9167_9466 );
and \U$10212 ( \19035_19334 , RIee27808_4908, \9169_9468 );
and \U$10213 ( \19036_19335 , RIfe8b788_7931, \9171_9470 );
and \U$10214 ( \19037_19336 , RIdf27ad8_1828, \9173_9472 );
and \U$10215 ( \19038_19337 , RIdf25d50_1807, \9175_9474 );
and \U$10216 ( \19039_19338 , RIdf24130_1787, \9177_9476 );
and \U$10217 ( \19040_19339 , RIfc66608_6187, \9179_9478 );
and \U$10218 ( \19041_19340 , RIfccde98_7365, \9181_9480 );
and \U$10219 ( \19042_19341 , RIfc66a40_6190, \9183_9482 );
and \U$10220 ( \19043_19342 , RIfc668d8_6189, \9185_9484 );
and \U$10221 ( \19044_19343 , RIfcacf40_6990, \9187_9486 );
and \U$10222 ( \19045_19344 , RIfeaaef8_8261, \9189_9488 );
and \U$10223 ( \19046_19345 , RIfc6e8d0_6280, \9191_9490 );
and \U$10224 ( \19047_19346 , RIdf18d30_1659, \9193_9492 );
and \U$10225 ( \19048_19347 , RIdf165d0_1631, \9195_9494 );
and \U$10226 ( \19049_19348 , RIdf138d0_1599, \9197_9496 );
and \U$10227 ( \19050_19349 , RIdf10bd0_1567, \9199_9498 );
and \U$10228 ( \19051_19350 , RIdf0ded0_1535, \9201_9500 );
and \U$10229 ( \19052_19351 , RIdf0b1d0_1503, \9203_9502 );
and \U$10230 ( \19053_19352 , RIdf084d0_1471, \9205_9504 );
and \U$10231 ( \19054_19353 , RIdf057d0_1439, \9207_9506 );
and \U$10232 ( \19055_19354 , RIdf02ad0_1407, \9209_9508 );
and \U$10233 ( \19056_19355 , RIdefd0d0_1343, \9211_9510 );
and \U$10234 ( \19057_19356 , RIdefa3d0_1311, \9213_9512 );
and \U$10235 ( \19058_19357 , RIdef76d0_1279, \9215_9514 );
and \U$10236 ( \19059_19358 , RIdef49d0_1247, \9217_9516 );
and \U$10237 ( \19060_19359 , RIdef1cd0_1215, \9219_9518 );
and \U$10238 ( \19061_19360 , RIdeeefd0_1183, \9221_9520 );
and \U$10239 ( \19062_19361 , RIdeec2d0_1151, \9223_9522 );
and \U$10240 ( \19063_19362 , RIdee95d0_1119, \9225_9524 );
and \U$10241 ( \19064_19363 , RIfc6dc28_6271, \9227_9526 );
and \U$10242 ( \19065_19364 , RIfc67c88_6203, \9229_9528 );
and \U$10243 ( \19066_19365 , RIfccb300_7334, \9231_9530 );
and \U$10244 ( \19067_19366 , RIfccd4c0_7358, \9233_9532 );
and \U$10245 ( \19068_19367 , RIfea81f8_8229, \9235_9534 );
and \U$10246 ( \19069_19368 , RIfea8360_8230, \9237_9536 );
and \U$10247 ( \19070_19369 , RIdee04f8_1016, \9239_9538 );
and \U$10248 ( \19071_19370 , RIdede338_992, \9241_9540 );
and \U$10249 ( \19072_19371 , RIfc6def8_6273, \9243_9542 );
and \U$10250 ( \19073_19372 , RIfcac130_6980, \9245_9544 );
and \U$10251 ( \19074_19373 , RIfc67b20_6202, \9247_9546 );
and \U$10252 ( \19075_19374 , RIfc67df0_6204, \9249_9548 );
and \U$10253 ( \19076_19375 , RIded9040_933, \9251_9550 );
and \U$10254 ( \19077_19376 , RIded6a48_906, \9253_9552 );
and \U$10255 ( \19078_19377 , RIded4b58_884, \9255_9554 );
and \U$10256 ( \19079_19378 , RIded26c8_858, \9257_9556 );
and \U$10257 ( \19080_19379 , RIdecfe00_829, \9259_9558 );
and \U$10258 ( \19081_19380 , RIdecd100_797, \9261_9560 );
and \U$10259 ( \19082_19381 , RIdeca400_765, \9263_9562 );
and \U$10260 ( \19083_19382 , RIdec7700_733, \9265_9564 );
and \U$10261 ( \19084_19383 , RIdeb3c00_509, \9267_9566 );
and \U$10262 ( \19085_19384 , RIde95228_317, \9269_9568 );
and \U$10263 ( \19086_19385 , RIe16d808_2623, \9271_9570 );
and \U$10264 ( \19087_19386 , RIe159600_2394, \9273_9572 );
and \U$10265 ( \19088_19387 , RIe142e00_2138, \9275_9574 );
and \U$10266 ( \19089_19388 , RIdf377f8_2008, \9277_9576 );
and \U$10267 ( \19090_19389 , RIdf2be58_1876, \9279_9578 );
and \U$10268 ( \19091_19390 , RIdf1c6d8_1700, \9281_9580 );
and \U$10269 ( \19092_19391 , RIdeffdd0_1375, \9283_9582 );
and \U$10270 ( \19093_19392 , RIdee68d0_1087, \9285_9584 );
and \U$10271 ( \19094_19393 , RIdedb638_960, \9287_9586 );
and \U$10272 ( \19095_19394 , RIde7b170_190, \9289_9588 );
or \U$10273 ( \19096_19395 , \19032_19331 , \19033_19332 , \19034_19333 , \19035_19334 , \19036_19335 , \19037_19336 , \19038_19337 , \19039_19338 , \19040_19339 , \19041_19340 , \19042_19341 , \19043_19342 , \19044_19343 , \19045_19344 , \19046_19345 , \19047_19346 , \19048_19347 , \19049_19348 , \19050_19349 , \19051_19350 , \19052_19351 , \19053_19352 , \19054_19353 , \19055_19354 , \19056_19355 , \19057_19356 , \19058_19357 , \19059_19358 , \19060_19359 , \19061_19360 , \19062_19361 , \19063_19362 , \19064_19363 , \19065_19364 , \19066_19365 , \19067_19366 , \19068_19367 , \19069_19368 , \19070_19369 , \19071_19370 , \19072_19371 , \19073_19372 , \19074_19373 , \19075_19374 , \19076_19375 , \19077_19376 , \19078_19377 , \19079_19378 , \19080_19379 , \19081_19380 , \19082_19381 , \19083_19382 , \19084_19383 , \19085_19384 , \19086_19385 , \19087_19386 , \19088_19387 , \19089_19388 , \19090_19389 , \19091_19390 , \19092_19391 , \19093_19392 , \19094_19393 , \19095_19394 );
or \U$10274 ( \19097_19396 , \19031_19330 , \19096_19395 );
_DC \g5461/U$1 ( \19098 , \19097_19396 , \9298_9597 );
and \U$10275 ( \19099_19398 , RIe19cc98_3161, \8760_9059 );
and \U$10276 ( \19100_19399 , RIe199f98_3129, \8762_9061 );
and \U$10277 ( \19101_19400 , RIfc73088_6331, \8764_9063 );
and \U$10278 ( \19102_19401 , RIe197298_3097, \8766_9065 );
and \U$10279 ( \19103_19402 , RIf1442a8_5235, \8768_9067 );
and \U$10280 ( \19104_19403 , RIe194598_3065, \8770_9069 );
and \U$10281 ( \19105_19404 , RIe191898_3033, \8772_9071 );
and \U$10282 ( \19106_19405 , RIe18eb98_3001, \8774_9073 );
and \U$10283 ( \19107_19406 , RIe189198_2937, \8776_9075 );
and \U$10284 ( \19108_19407 , RIe186498_2905, \8778_9077 );
and \U$10285 ( \19109_19408 , RIfc72278_6321, \8780_9079 );
and \U$10286 ( \19110_19409 , RIe183798_2873, \8782_9081 );
and \U$10287 ( \19111_19410 , RIfc61ce8_6135, \8784_9083 );
and \U$10288 ( \19112_19411 , RIe180a98_2841, \8786_9085 );
and \U$10289 ( \19113_19412 , RIe17dd98_2809, \8788_9087 );
and \U$10290 ( \19114_19413 , RIe17b098_2777, \8790_9089 );
and \U$10291 ( \19115_19414 , RIfcaf268_7015, \8792_9091 );
and \U$10292 ( \19116_19415 , RIfca6a00_6918, \8794_9093 );
and \U$10293 ( \19117_19416 , RIfcc9b18_7317, \8796_9095 );
and \U$10294 ( \19118_19417 , RIe175530_2712, \8798_9097 );
and \U$10295 ( \19119_19418 , RIfc72818_6325, \8800_9099 );
and \U$10296 ( \19120_19419 , RIfc726b0_6324, \8802_9101 );
and \U$10297 ( \19121_19420 , RIfccf7e8_7383, \8804_9103 );
and \U$10298 ( \19122_19421 , RIfc72548_6323, \8806_9105 );
and \U$10299 ( \19123_19422 , RIee3be48_5140, \8808_9107 );
and \U$10300 ( \19124_19423 , RIee3ad68_5128, \8810_9109 );
and \U$10301 ( \19125_19424 , RIfc71fa8_6319, \8812_9111 );
and \U$10302 ( \19126_19425 , RIe1730a0_2686, \8814_9113 );
and \U$10303 ( \19127_19426 , RIfcaef98_7013, \8816_9115 );
and \U$10304 ( \19128_19427 , RIfccf518_7381, \8818_9117 );
and \U$10305 ( \19129_19428 , RIfc71e40_6318, \8820_9119 );
and \U$10306 ( \19130_19429 , RIfc62120_6138, \8822_9121 );
and \U$10307 ( \19131_19430 , RIfe8b350_7928, \8824_9123 );
and \U$10308 ( \19132_19431 , RIe222ff0_4688, \8826_9125 );
and \U$10309 ( \19133_19432 , RIfcc9f50_7320, \8828_9127 );
and \U$10310 ( \19134_19433 , RIe2202f0_4656, \8830_9129 );
and \U$10311 ( \19135_19434 , RIfc4a570_5868, \8832_9131 );
and \U$10312 ( \19136_19435 , RIe21d5f0_4624, \8834_9133 );
and \U$10313 ( \19137_19436 , RIe217bf0_4560, \8836_9135 );
and \U$10314 ( \19138_19437 , RIe214ef0_4528, \8838_9137 );
and \U$10315 ( \19139_19438 , RIfccf3b0_7380, \8840_9139 );
and \U$10316 ( \19140_19439 , RIe2121f0_4496, \8842_9141 );
and \U$10317 ( \19141_19440 , RIf168ba8_5651, \8844_9143 );
and \U$10318 ( \19142_19441 , RIe20f4f0_4464, \8846_9145 );
and \U$10319 ( \19143_19442 , RIfc71300_6310, \8848_9147 );
and \U$10320 ( \19144_19443 , RIe20c7f0_4432, \8850_9149 );
and \U$10321 ( \19145_19444 , RIe209af0_4400, \8852_9151 );
and \U$10322 ( \19146_19445 , RIe206df0_4368, \8854_9153 );
and \U$10323 ( \19147_19446 , RIfc718a0_6314, \8856_9155 );
and \U$10324 ( \19148_19447 , RIfc71a08_6315, \8858_9157 );
and \U$10325 ( \19149_19448 , RIe202098_4313, \8860_9159 );
and \U$10326 ( \19150_19449 , RIfe8b1e8_7927, \8862_9161 );
and \U$10327 ( \19151_19450 , RIfc715d0_6312, \8864_9163 );
and \U$10328 ( \19152_19451 , RIfce6588_7643, \8866_9165 );
and \U$10329 ( \19153_19452 , RIfc62c60_6146, \8868_9167 );
and \U$10330 ( \19154_19453 , RIf161858_5569, \8870_9169 );
and \U$10331 ( \19155_19454 , RIf15fad0_5548, \8872_9171 );
and \U$10332 ( \19156_19455 , RIf15dbe0_5526, \8874_9173 );
and \U$10333 ( \19157_19456 , RIe1fc698_4249, \8876_9175 );
and \U$10334 ( \19158_19457 , RIfe8b4b8_7929, \8878_9177 );
and \U$10335 ( \19159_19458 , RIfcae5c0_7006, \8880_9179 );
and \U$10336 ( \19160_19459 , RIfc63098_6149, \8882_9181 );
and \U$10337 ( \19161_19460 , RIfc63200_6150, \8884_9183 );
and \U$10338 ( \19162_19461 , RIfc71198_6309, \8886_9185 );
or \U$10339 ( \19163_19462 , \19099_19398 , \19100_19399 , \19101_19400 , \19102_19401 , \19103_19402 , \19104_19403 , \19105_19404 , \19106_19405 , \19107_19406 , \19108_19407 , \19109_19408 , \19110_19409 , \19111_19410 , \19112_19411 , \19113_19412 , \19114_19413 , \19115_19414 , \19116_19415 , \19117_19416 , \19118_19417 , \19119_19418 , \19120_19419 , \19121_19420 , \19122_19421 , \19123_19422 , \19124_19423 , \19125_19424 , \19126_19425 , \19127_19426 , \19128_19427 , \19129_19428 , \19130_19429 , \19131_19430 , \19132_19431 , \19133_19432 , \19134_19433 , \19135_19434 , \19136_19435 , \19137_19436 , \19138_19437 , \19139_19438 , \19140_19439 , \19141_19440 , \19142_19441 , \19143_19442 , \19144_19443 , \19145_19444 , \19146_19445 , \19147_19446 , \19148_19447 , \19149_19448 , \19150_19449 , \19151_19450 , \19152_19451 , \19153_19452 , \19154_19453 , \19155_19454 , \19156_19455 , \19157_19456 , \19158_19457 , \19159_19458 , \19160_19459 , \19161_19460 , \19162_19461 );
and \U$10340 ( \19164_19463 , RIf158a50_5468, \8889_9188 );
and \U$10341 ( \19165_19464 , RIf1576a0_5454, \8891_9190 );
and \U$10342 ( \19166_19465 , RIfcdc808_7531, \8893_9192 );
and \U$10343 ( \19167_19466 , RIfe8b620_7930, \8895_9194 );
and \U$10344 ( \19168_19467 , RIfc634d0_6152, \8897_9196 );
and \U$10345 ( \19169_19468 , RIfcceb40_7374, \8899_9198 );
and \U$10346 ( \19170_19469 , RIf154400_5418, \8901_9200 );
and \U$10347 ( \19171_19470 , RIe1f4da8_4163, \8903_9202 );
and \U$10348 ( \19172_19471 , RIf152c18_5401, \8905_9204 );
and \U$10349 ( \19173_19472 , RIf151868_5387, \8907_9206 );
and \U$10350 ( \19174_19473 , RIfc4d108_5899, \8909_9208 );
and \U$10351 ( \19175_19474 , RIe1f2a80_4138, \8911_9210 );
and \U$10352 ( \19176_19475 , RIfc70a90_6304, \8913_9212 );
and \U$10353 ( \19177_19476 , RIfc63bd8_6157, \8915_9214 );
and \U$10354 ( \19178_19477 , RIfca7810_6928, \8917_9216 );
and \U$10355 ( \19179_19478 , RIe1ed788_4079, \8919_9218 );
and \U$10356 ( \19180_19479 , RIe1ead58_4049, \8921_9220 );
and \U$10357 ( \19181_19480 , RIe1e8058_4017, \8923_9222 );
and \U$10358 ( \19182_19481 , RIe1e5358_3985, \8925_9224 );
and \U$10359 ( \19183_19482 , RIe1e2658_3953, \8927_9226 );
and \U$10360 ( \19184_19483 , RIe1df958_3921, \8929_9228 );
and \U$10361 ( \19185_19484 , RIe1dcc58_3889, \8931_9230 );
and \U$10362 ( \19186_19485 , RIe1d9f58_3857, \8933_9232 );
and \U$10363 ( \19187_19486 , RIe1d7258_3825, \8935_9234 );
and \U$10364 ( \19188_19487 , RIe1d1858_3761, \8937_9236 );
and \U$10365 ( \19189_19488 , RIe1ceb58_3729, \8939_9238 );
and \U$10366 ( \19190_19489 , RIe1cbe58_3697, \8941_9240 );
and \U$10367 ( \19191_19490 , RIe1c9158_3665, \8943_9242 );
and \U$10368 ( \19192_19491 , RIe1c6458_3633, \8945_9244 );
and \U$10369 ( \19193_19492 , RIe1c3758_3601, \8947_9246 );
and \U$10370 ( \19194_19493 , RIe1c0a58_3569, \8949_9248 );
and \U$10371 ( \19195_19494 , RIe1bdd58_3537, \8951_9250 );
and \U$10372 ( \19196_19495 , RIf14c408_5327, \8953_9252 );
and \U$10373 ( \19197_19496 , RIf14b1c0_5314, \8955_9254 );
and \U$10374 ( \19198_19497 , RIe1b8d30_3480, \8957_9256 );
and \U$10375 ( \19199_19498 , RIe1b6cd8_3457, \8959_9258 );
and \U$10376 ( \19200_19499 , RIfc707c0_6302, \8961_9260 );
and \U$10377 ( \19201_19500 , RIfca7c48_6931, \8963_9262 );
and \U$10378 ( \19202_19501 , RIe1b4de8_3435, \8965_9264 );
and \U$10379 ( \19203_19502 , RIe1b3a38_3421, \8967_9266 );
and \U$10380 ( \19204_19503 , RIfc70220_6298, \8969_9268 );
and \U$10381 ( \19205_19504 , RIfcce870_7372, \8971_9270 );
and \U$10382 ( \19206_19505 , RIe1b23b8_3405, \8973_9272 );
and \U$10383 ( \19207_19506 , RIe1b0630_3384, \8975_9274 );
and \U$10384 ( \19208_19507 , RIfc645b0_6164, \8977_9276 );
and \U$10385 ( \19209_19508 , RIfc700b8_6297, \8979_9278 );
and \U$10386 ( \19210_19509 , RIfeaac28_8259, \8981_9280 );
and \U$10387 ( \19211_19510 , RIe1aa690_3316, \8983_9282 );
and \U$10388 ( \19212_19511 , RIe1a8098_3289, \8985_9284 );
and \U$10389 ( \19213_19512 , RIe1a5398_3257, \8987_9286 );
and \U$10390 ( \19214_19513 , RIe1a2698_3225, \8989_9288 );
and \U$10391 ( \19215_19514 , RIe19f998_3193, \8991_9290 );
and \U$10392 ( \19216_19515 , RIe18be98_2969, \8993_9292 );
and \U$10393 ( \19217_19516 , RIe178398_2745, \8995_9294 );
and \U$10394 ( \19218_19517 , RIe225cf0_4720, \8997_9296 );
and \U$10395 ( \19219_19518 , RIe21a8f0_4592, \8999_9298 );
and \U$10396 ( \19220_19519 , RIe2040f0_4336, \9001_9300 );
and \U$10397 ( \19221_19520 , RIe1fe150_4268, \9003_9302 );
and \U$10398 ( \19222_19521 , RIe1f7508_4191, \9005_9304 );
and \U$10399 ( \19223_19522 , RIe1f0050_4108, \9007_9306 );
and \U$10400 ( \19224_19523 , RIe1d4558_3793, \9009_9308 );
and \U$10401 ( \19225_19524 , RIe1bb058_3505, \9011_9310 );
and \U$10402 ( \19226_19525 , RIe1aded0_3356, \9013_9312 );
and \U$10403 ( \19227_19526 , RIe170508_2655, \9015_9314 );
or \U$10404 ( \19228_19527 , \19164_19463 , \19165_19464 , \19166_19465 , \19167_19466 , \19168_19467 , \19169_19468 , \19170_19469 , \19171_19470 , \19172_19471 , \19173_19472 , \19174_19473 , \19175_19474 , \19176_19475 , \19177_19476 , \19178_19477 , \19179_19478 , \19180_19479 , \19181_19480 , \19182_19481 , \19183_19482 , \19184_19483 , \19185_19484 , \19186_19485 , \19187_19486 , \19188_19487 , \19189_19488 , \19190_19489 , \19191_19490 , \19192_19491 , \19193_19492 , \19194_19493 , \19195_19494 , \19196_19495 , \19197_19496 , \19198_19497 , \19199_19498 , \19200_19499 , \19201_19500 , \19202_19501 , \19203_19502 , \19204_19503 , \19205_19504 , \19206_19505 , \19207_19506 , \19208_19507 , \19209_19508 , \19210_19509 , \19211_19510 , \19212_19511 , \19213_19512 , \19214_19513 , \19215_19514 , \19216_19515 , \19217_19516 , \19218_19517 , \19219_19518 , \19220_19519 , \19221_19520 , \19222_19521 , \19223_19522 , \19224_19523 , \19225_19524 , \19226_19525 , \19227_19526 );
or \U$10405 ( \19229_19528 , \19163_19462 , \19228_19527 );
_DC \g54e5/U$1 ( \19230 , \19229_19528 , \9024_9323 );
xor g54e6_GF_PartitionCandidate( \19231_19530_nG54e6 , \19098 , \19230 );
buf \U$10406 ( \19232_19531 , \19231_19530_nG54e6 );
xor \U$10407 ( \19233_19532 , \19232_19531 , \18742_19044 );
not \U$10408 ( \19234_19533 , \18743_19045 );
and \U$10409 ( \19235_19534 , \19233_19532 , \19234_19533 );
and \U$10410 ( \19236_19535 , \10385_10687 , \19235_19534 );
and \U$10411 ( \19237_19536 , \10686_10988 , \18743_19045 );
nor \U$10412 ( \19238_19537 , \19236_19535 , \19237_19536 );
and \U$10413 ( \19239_19538 , \18742_19044 , \17744_18043 );
not \U$10414 ( \19240_19539 , \19239_19538 );
and \U$10415 ( \19241_19540 , \19232_19531 , \19240_19539 );
xnor \U$10416 ( \19242_19541 , \19238_19537 , \19241_19540 );
xor \U$10417 ( \19243_19542 , \18966_19265 , \19242_19541 );
xor \U$10418 ( \19244_19543 , \18957_19256 , \19243_19542 );
xor \U$10419 ( \19245_19544 , \18938_19237 , \19244_19543 );
and \U$10420 ( \19246_19545 , \18767_19069 , \18771_19073 );
and \U$10421 ( \19247_19546 , \18771_19073 , \18776_19078 );
and \U$10422 ( \19248_19547 , \18767_19069 , \18776_19078 );
or \U$10423 ( \19249_19548 , \19246_19545 , \19247_19546 , \19248_19547 );
and \U$10424 ( \19250_19549 , \18458_18760 , \18462_18764 );
and \U$10425 ( \19251_19550 , \18462_18764 , \18745_19047 );
and \U$10426 ( \19252_19551 , \18458_18760 , \18745_19047 );
or \U$10427 ( \19253_19552 , \19250_19549 , \19251_19550 , \19252_19551 );
xor \U$10428 ( \19254_19553 , \19249_19548 , \19253_19552 );
and \U$10429 ( \19255_19554 , \18730_19032 , \10681_10983 );
_DC \g65a4/U$1 ( \19256 , \19097_19396 , \9298_9597 );
_DC \g65a5/U$1 ( \19257 , \19229_19528 , \9024_9323 );
and g65a6_GF_PartitionCandidate( \19258_19557_nG65a6 , \19256 , \19257 );
buf \U$10430 ( \19259_19558 , \19258_19557_nG65a6 );
and \U$10431 ( \19260_19559 , \19259_19558 , \10389_10691 );
nor \U$10432 ( \19261_19560 , \19255_19554 , \19260_19559 );
xnor \U$10433 ( \19262_19561 , \19261_19560 , \10678_10980 );
not \U$10434 ( \19263_19562 , \18744_19046 );
and \U$10435 ( \19264_19563 , \19263_19562 , \19241_19540 );
xor \U$10436 ( \19265_19564 , \19262_19561 , \19264_19563 );
and \U$10437 ( \19266_19565 , \18733_19035 , \18737_19039 );
and \U$10438 ( \19267_19566 , \18737_19039 , \18744_19046 );
and \U$10439 ( \19268_19567 , \18733_19035 , \18744_19046 );
or \U$10440 ( \19269_19568 , \19266_19565 , \19267_19566 , \19268_19567 );
xor \U$10441 ( \19270_19569 , \19265_19564 , \19269_19568 );
and \U$10442 ( \19271_19570 , \10968_11270 , \17791_18090 );
and \U$10443 ( \19272_19571 , \11287_11586 , \17353_17655 );
nor \U$10444 ( \19273_19572 , \19271_19570 , \19272_19571 );
xnor \U$10445 ( \19274_19573 , \19273_19572 , \17747_18046 );
xor \U$10446 ( \19275_19574 , \19270_19569 , \19274_19573 );
xor \U$10447 ( \19276_19575 , \19254_19553 , \19275_19574 );
xor \U$10448 ( \19277_19576 , \19245_19544 , \19276_19575 );
and \U$10449 ( \19278_19577 , \18454_18756 , \18746_19048 );
and \U$10450 ( \19279_19578 , \18746_19048 , \18778_19080 );
and \U$10451 ( \19280_19579 , \18454_18756 , \18778_19080 );
or \U$10452 ( \19281_19580 , \19278_19577 , \19279_19578 , \19280_19579 );
xor \U$10453 ( \19282_19581 , \19277_19576 , \19281_19580 );
and \U$10454 ( \19283_19582 , \18779_19081 , \18783_19085 );
and \U$10455 ( \19284_19583 , \18784_19086 , \18787_19089 );
or \U$10456 ( \19285_19584 , \19283_19582 , \19284_19583 );
xor \U$10457 ( \19286_19585 , \19282_19581 , \19285_19584 );
buf g9be1_GF_PartitionCandidate( \19287_19586_nG9be1 , \19286_19585 );
and \U$10458 ( \19288_19587 , \10402_10704 , \19287_19586_nG9be1 );
or \U$10459 ( \19289_19588 , \18934_19233 , \19288_19587 );
xor \U$10460 ( \19290_19589 , \10399_10703 , \19289_19588 );
buf \U$10461 ( \19291_19590 , \19290_19589 );
buf \U$10463 ( \19292_19591 , \19291_19590 );
xor \U$10464 ( \19293_19592 , \18933_19232 , \19292_19591 );
buf \U$10465 ( \19294_19593 , \19293_19592 );
xor \U$10466 ( \19295_19594 , \18884_19186 , \19294_19593 );
buf \U$10467 ( \19296_19595 , \19295_19594 );
xor \U$10468 ( \19297_19596 , \18847_19149 , \19296_19595 );
and \U$10469 ( \19298_19597 , \18417_18719 , \18796_19098 );
and \U$10470 ( \19299_19598 , \18417_18719 , \18830_19132 );
and \U$10471 ( \19300_19599 , \18796_19098 , \18830_19132 );
or \U$10472 ( \19301_19600 , \19298_19597 , \19299_19598 , \19300_19599 );
buf \U$10473 ( \19302_19601 , \19301_19600 );
xor \U$10474 ( \19303_19602 , \19297_19596 , \19302_19601 );
and \U$10475 ( \19304_19603 , \18842_19144 , \19303_19602 );
and \U$10476 ( \19305_19604 , RIdec4cd0_703, \8760_9059 );
and \U$10477 ( \19306_19605 , RIdec1fd0_671, \8762_9061 );
and \U$10478 ( \19307_19606 , RIfc7b4b8_6425, \8764_9063 );
and \U$10479 ( \19308_19607 , RIdebf2d0_639, \8766_9065 );
and \U$10480 ( \19309_19608 , RIfc7b1e8_6423, \8768_9067 );
and \U$10481 ( \19310_19609 , RIdebc5d0_607, \8770_9069 );
and \U$10482 ( \19311_19610 , RIdeb98d0_575, \8772_9071 );
and \U$10483 ( \19312_19611 , RIdeb6bd0_543, \8774_9073 );
and \U$10484 ( \19313_19612 , RIfe83358_7837, \8776_9075 );
and \U$10485 ( \19314_19613 , RIdeb11d0_479, \8778_9077 );
and \U$10486 ( \19315_19614 , RIee1e5c8_4804, \8780_9079 );
and \U$10487 ( \19316_19615 , RIdeae4d0_447, \8782_9081 );
and \U$10488 ( \19317_19616 , RIfc437c0_5790, \8784_9083 );
and \U$10489 ( \19318_19617 , RIdea93b8_415, \8786_9085 );
and \U$10490 ( \19319_19618 , RIdea2ab8_383, \8788_9087 );
and \U$10491 ( \19320_19619 , RIde9c1b8_351, \8790_9089 );
and \U$10492 ( \19321_19620 , RIfc90ea8_6671, \8792_9091 );
and \U$10493 ( \19322_19621 , RIfc7af18_6421, \8794_9093 );
and \U$10494 ( \19323_19622 , RIfe83088_7835, \8796_9095 );
and \U$10495 ( \19324_19623 , RIee1a950_4761, \8798_9097 );
and \U$10496 ( \19325_19624 , RIde906b0_294, \8800_9099 );
and \U$10497 ( \19326_19625 , RIde8cba0_276, \8802_9101 );
and \U$10498 ( \19327_19626 , RIfe82f20_7834, \8804_9103 );
and \U$10499 ( \19328_19627 , RIfe82db8_7833, \8806_9105 );
and \U$10500 ( \19329_19628 , RIee1a248_4756, \8808_9107 );
and \U$10501 ( \19330_19629 , RIfe831f0_7836, \8810_9109 );
and \U$10502 ( \19331_19630 , RIfcc2390_7232, \8812_9111 );
and \U$10503 ( \19332_19631 , RIee195a0_4747, \8814_9113 );
and \U$10504 ( \19333_19632 , RIfcbe718_7189, \8816_9115 );
and \U$10505 ( \19334_19633 , RIfea9e18_8249, \8818_9117 );
and \U$10506 ( \19335_19634 , RIfc43220_5786, \8820_9119 );
and \U$10507 ( \19336_19635 , RIe167868_2555, \8822_9121 );
and \U$10508 ( \19337_19636 , RIe164cd0_2524, \8824_9123 );
and \U$10509 ( \19338_19637 , RIe161fd0_2492, \8826_9125 );
and \U$10510 ( \19339_19638 , RIee36f88_5084, \8828_9127 );
and \U$10511 ( \19340_19639 , RIe15f2d0_2460, \8830_9129 );
and \U$10512 ( \19341_19640 , RIee35ea8_5072, \8832_9131 );
and \U$10513 ( \19342_19641 , RIe15c5d0_2428, \8834_9133 );
and \U$10514 ( \19343_19642 , RIe156bd0_2364, \8836_9135 );
and \U$10515 ( \19344_19643 , RIe153ed0_2332, \8838_9137 );
and \U$10516 ( \19345_19644 , RIfe83628_7839, \8840_9139 );
and \U$10517 ( \19346_19645 , RIe1511d0_2300, \8842_9141 );
and \U$10518 ( \19347_19646 , RIfebfda8_8303, \8844_9143 );
and \U$10519 ( \19348_19647 , RIe14e4d0_2268, \8846_9145 );
and \U$10520 ( \19349_19648 , RIfebfc40_8302, \8848_9147 );
and \U$10521 ( \19350_19649 , RIe14b7d0_2236, \8850_9149 );
and \U$10522 ( \19351_19650 , RIe148ad0_2204, \8852_9151 );
and \U$10523 ( \19352_19651 , RIe145dd0_2172, \8854_9153 );
and \U$10524 ( \19353_19652 , RIee34120_5051, \8856_9155 );
and \U$10525 ( \19354_19653 , RIee32ed8_5038, \8858_9157 );
and \U$10526 ( \19355_19654 , RIee31df8_5026, \8860_9159 );
and \U$10527 ( \19356_19655 , RIfcc1f58_7229, \8862_9161 );
and \U$10528 ( \19357_19656 , RIe140ad8_2113, \8864_9163 );
and \U$10529 ( \19358_19657 , RIdf3e878_2088, \8866_9165 );
and \U$10530 ( \19359_19658 , RIfe834c0_7838, \8868_9167 );
and \U$10531 ( \19360_19659 , RIdf3a390_2039, \8870_9169 );
and \U$10532 ( \19361_19660 , RIfc5a6c8_6051, \8872_9171 );
and \U$10533 ( \19362_19661 , RIfc91e20_6682, \8874_9173 );
and \U$10534 ( \19363_19662 , RIee2e888_4988, \8876_9175 );
and \U$10535 ( \19364_19663 , RIfc96a10_6736, \8878_9177 );
and \U$10536 ( \19365_19664 , RIdf35098_1980, \8880_9179 );
and \U$10537 ( \19366_19665 , RIfeab600_8266, \8882_9181 );
and \U$10538 ( \19367_19666 , RIdf30bb0_1931, \8884_9183 );
and \U$10539 ( \19368_19667 , RIfeab768_8267, \8886_9185 );
or \U$10540 ( \19369_19668 , \19305_19604 , \19306_19605 , \19307_19606 , \19308_19607 , \19309_19608 , \19310_19609 , \19311_19610 , \19312_19611 , \19313_19612 , \19314_19613 , \19315_19614 , \19316_19615 , \19317_19616 , \19318_19617 , \19319_19618 , \19320_19619 , \19321_19620 , \19322_19621 , \19323_19622 , \19324_19623 , \19325_19624 , \19326_19625 , \19327_19626 , \19328_19627 , \19329_19628 , \19330_19629 , \19331_19630 , \19332_19631 , \19333_19632 , \19334_19633 , \19335_19634 , \19336_19635 , \19337_19636 , \19338_19637 , \19339_19638 , \19340_19639 , \19341_19640 , \19342_19641 , \19343_19642 , \19344_19643 , \19345_19644 , \19346_19645 , \19347_19646 , \19348_19647 , \19349_19648 , \19350_19649 , \19351_19650 , \19352_19651 , \19353_19652 , \19354_19653 , \19355_19654 , \19356_19655 , \19357_19656 , \19358_19657 , \19359_19658 , \19360_19659 , \19361_19660 , \19362_19661 , \19363_19662 , \19364_19663 , \19365_19664 , \19366_19665 , \19367_19666 , \19368_19667 );
and \U$10541 ( \19370_19669 , RIfcbe9e8_7191, \8889_9188 );
and \U$10542 ( \19371_19670 , RIfc79fa0_6410, \8891_9190 );
and \U$10543 ( \19372_19671 , RIfc96740_6734, \8893_9192 );
and \U$10544 ( \19373_19672 , RIfc92258_6685, \8895_9194 );
and \U$10545 ( \19374_19673 , RIfea7118_8217, \8897_9196 );
and \U$10546 ( \19375_19674 , RIfea95a8_8243, \8899_9198 );
and \U$10547 ( \19376_19675 , RIdf26020_1809, \8901_9200 );
and \U$10548 ( \19377_19676 , RIdf24400_1789, \8903_9202 );
and \U$10549 ( \19378_19677 , RIfc79a00_6406, \8905_9204 );
and \U$10550 ( \19379_19678 , RIfc5add0_6056, \8907_9206 );
and \U$10551 ( \19380_19679 , RIfce5d18_7637, \8909_9208 );
and \U$10552 ( \19381_19680 , RIfc92690_6688, \8911_9210 );
and \U$10553 ( \19382_19681 , RIfce3018_7605, \8913_9212 );
and \U$10554 ( \19383_19682 , RIdf1f270_1731, \8915_9214 );
and \U$10555 ( \19384_19683 , RIfc79730_6404, \8917_9216 );
and \U$10556 ( \19385_19684 , RIdf19000_1661, \8919_9218 );
and \U$10557 ( \19386_19685 , RIdf168a0_1633, \8921_9220 );
and \U$10558 ( \19387_19686 , RIdf13ba0_1601, \8923_9222 );
and \U$10559 ( \19388_19687 , RIdf10ea0_1569, \8925_9224 );
and \U$10560 ( \19389_19688 , RIdf0e1a0_1537, \8927_9226 );
and \U$10561 ( \19390_19689 , RIdf0b4a0_1505, \8929_9228 );
and \U$10562 ( \19391_19690 , RIdf087a0_1473, \8931_9230 );
and \U$10563 ( \19392_19691 , RIdf05aa0_1441, \8933_9232 );
and \U$10564 ( \19393_19692 , RIdf02da0_1409, \8935_9234 );
and \U$10565 ( \19394_19693 , RIdefd3a0_1345, \8937_9236 );
and \U$10566 ( \19395_19694 , RIdefa6a0_1313, \8939_9238 );
and \U$10567 ( \19396_19695 , RIdef79a0_1281, \8941_9240 );
and \U$10568 ( \19397_19696 , RIdef4ca0_1249, \8943_9242 );
and \U$10569 ( \19398_19697 , RIdef1fa0_1217, \8945_9244 );
and \U$10570 ( \19399_19698 , RIdeef2a0_1185, \8947_9246 );
and \U$10571 ( \19400_19699 , RIdeec5a0_1153, \8949_9248 );
and \U$10572 ( \19401_19700 , RIdee98a0_1121, \8951_9250 );
and \U$10573 ( \19402_19701 , RIfc5b7a8_6063, \8953_9252 );
and \U$10574 ( \19403_19702 , RIfc5b640_6062, \8955_9254 );
and \U$10575 ( \19404_19703 , RIfc931d0_6696, \8957_9256 );
and \U$10576 ( \19405_19704 , RIfcecac8_7715, \8959_9258 );
and \U$10577 ( \19406_19705 , RIdee4710_1063, \8961_9260 );
and \U$10578 ( \19407_19706 , RIdee26b8_1040, \8963_9262 );
and \U$10579 ( \19408_19707 , RIdee07c8_1018, \8965_9264 );
and \U$10580 ( \19409_19708 , RIdede4a0_993, \8967_9266 );
and \U$10581 ( \19410_19709 , RIfcbf0f0_7196, \8969_9268 );
and \U$10582 ( \19411_19710 , RIfcbf528_7199, \8971_9270 );
and \U$10583 ( \19412_19711 , RIfc792f8_6401, \8973_9272 );
and \U$10584 ( \19413_19712 , RIfc93068_6695, \8975_9274 );
and \U$10585 ( \19414_19713 , RIded91a8_934, \8977_9276 );
and \U$10586 ( \19415_19714 , RIded6d18_908, \8979_9278 );
and \U$10587 ( \19416_19715 , RIded4e28_886, \8981_9280 );
and \U$10588 ( \19417_19716 , RIded2998_860, \8983_9282 );
and \U$10589 ( \19418_19717 , RIded00d0_831, \8985_9284 );
and \U$10590 ( \19419_19718 , RIdecd3d0_799, \8987_9286 );
and \U$10591 ( \19420_19719 , RIdeca6d0_767, \8989_9288 );
and \U$10592 ( \19421_19720 , RIdec79d0_735, \8991_9290 );
and \U$10593 ( \19422_19721 , RIdeb3ed0_511, \8993_9292 );
and \U$10594 ( \19423_19722 , RIde958b8_319, \8995_9294 );
and \U$10595 ( \19424_19723 , RIe16dad8_2625, \8997_9296 );
and \U$10596 ( \19425_19724 , RIe1598d0_2396, \8999_9298 );
and \U$10597 ( \19426_19725 , RIe1430d0_2140, \9001_9300 );
and \U$10598 ( \19427_19726 , RIdf37ac8_2010, \9003_9302 );
and \U$10599 ( \19428_19727 , RIdf2c128_1878, \9005_9304 );
and \U$10600 ( \19429_19728 , RIdf1c9a8_1702, \9007_9306 );
and \U$10601 ( \19430_19729 , RIdf000a0_1377, \9009_9308 );
and \U$10602 ( \19431_19730 , RIdee6ba0_1089, \9011_9310 );
and \U$10603 ( \19432_19731 , RIdedb908_962, \9013_9312 );
and \U$10604 ( \19433_19732 , RIde7b800_192, \9015_9314 );
or \U$10605 ( \19434_19733 , \19370_19669 , \19371_19670 , \19372_19671 , \19373_19672 , \19374_19673 , \19375_19674 , \19376_19675 , \19377_19676 , \19378_19677 , \19379_19678 , \19380_19679 , \19381_19680 , \19382_19681 , \19383_19682 , \19384_19683 , \19385_19684 , \19386_19685 , \19387_19686 , \19388_19687 , \19389_19688 , \19390_19689 , \19391_19690 , \19392_19691 , \19393_19692 , \19394_19693 , \19395_19694 , \19396_19695 , \19397_19696 , \19398_19697 , \19399_19698 , \19400_19699 , \19401_19700 , \19402_19701 , \19403_19702 , \19404_19703 , \19405_19704 , \19406_19705 , \19407_19706 , \19408_19707 , \19409_19708 , \19410_19709 , \19411_19710 , \19412_19711 , \19413_19712 , \19414_19713 , \19415_19714 , \19416_19715 , \19417_19716 , \19418_19717 , \19419_19718 , \19420_19719 , \19421_19720 , \19422_19721 , \19423_19722 , \19424_19723 , \19425_19724 , \19426_19725 , \19427_19726 , \19428_19727 , \19429_19728 , \19430_19729 , \19431_19730 , \19432_19731 , \19433_19732 );
or \U$10606 ( \19435_19734 , \19369_19668 , \19434_19733 );
_DC \g297b/U$1 ( \19436 , \19435_19734 , \9024_9323 );
buf \U$10607 ( \19437_19736 , \19436 );
and \U$10608 ( \19438_19737 , RIe19cf68_3163, \9034_9333 );
and \U$10609 ( \19439_19738 , RIe19a268_3131, \9036_9335 );
and \U$10610 ( \19440_19739 , RIfc8d7d0_6632, \9038_9337 );
and \U$10611 ( \19441_19740 , RIe197568_3099, \9040_9339 );
and \U$10612 ( \19442_19741 , RIfc561e0_6002, \9042_9341 );
and \U$10613 ( \19443_19742 , RIe194868_3067, \9044_9343 );
and \U$10614 ( \19444_19743 , RIe191b68_3035, \9046_9345 );
and \U$10615 ( \19445_19744 , RIe18ee68_3003, \9048_9347 );
and \U$10616 ( \19446_19745 , RIe189468_2939, \9050_9349 );
and \U$10617 ( \19447_19746 , RIe186768_2907, \9052_9351 );
and \U$10618 ( \19448_19747 , RIf143330_5224, \9054_9353 );
and \U$10619 ( \19449_19748 , RIe183a68_2875, \9056_9355 );
and \U$10620 ( \19450_19749 , RIfc7d948_6451, \9058_9357 );
and \U$10621 ( \19451_19750 , RIe180d68_2843, \9060_9359 );
and \U$10622 ( \19452_19751 , RIe17e068_2811, \9062_9361 );
and \U$10623 ( \19453_19752 , RIe17b368_2779, \9064_9363 );
and \U$10624 ( \19454_19753 , RIfc564b0_6004, \9066_9365 );
and \U$10625 ( \19455_19754 , RIfcd6700_7462, \9068_9367 );
and \U$10626 ( \19456_19755 , RIfc461f0_5820, \9070_9369 );
and \U$10627 ( \19457_19756 , RIe175698_2713, \9072_9371 );
and \U$10628 ( \19458_19757 , RIfc46088_5819, \9074_9373 );
and \U$10629 ( \19459_19758 , RIfc45f20_5818, \9076_9375 );
and \U$10630 ( \19460_19759 , RIfc7dc18_6453, \9078_9377 );
and \U$10631 ( \19461_19760 , RIfcd69d0_7464, \9080_9379 );
and \U$10632 ( \19462_19761 , RIfc98630_6756, \9082_9381 );
and \U$10633 ( \19463_19762 , RIfcc2a98_7237, \9084_9383 );
and \U$10634 ( \19464_19763 , RIfc7d510_6448, \9086_9385 );
and \U$10635 ( \19465_19764 , RIe173208_2687, \9088_9387 );
and \U$10636 ( \19466_19765 , RIfc8e478_6641, \9090_9389 );
and \U$10637 ( \19467_19766 , RIfc45ae8_5815, \9092_9391 );
and \U$10638 ( \19468_19767 , RIfc8e8b0_6644, \9094_9393 );
and \U$10639 ( \19469_19768 , RIfc45980_5814, \9096_9395 );
and \U$10640 ( \19470_19769 , RIfe82ae8_7831, \9098_9397 );
and \U$10641 ( \19471_19770 , RIe2232c0_4690, \9100_9399 );
and \U$10642 ( \19472_19771 , RIf16ba10_5684, \9102_9401 );
and \U$10643 ( \19473_19772 , RIe2205c0_4658, \9104_9403 );
and \U$10644 ( \19474_19773 , RIfcd24e8_7415, \9106_9405 );
and \U$10645 ( \19475_19774 , RIe21d8c0_4626, \9108_9407 );
and \U$10646 ( \19476_19775 , RIe217ec0_4562, \9110_9409 );
and \U$10647 ( \19477_19776 , RIe2151c0_4530, \9112_9411 );
and \U$10648 ( \19478_19777 , RIfebf268_8295, \9114_9413 );
and \U$10649 ( \19479_19778 , RIe2124c0_4498, \9116_9415 );
and \U$10650 ( \19480_19779 , RIf168d10_5652, \9118_9417 );
and \U$10651 ( \19481_19780 , RIe20f7c0_4466, \9120_9419 );
and \U$10652 ( \19482_19781 , RIfc7d240_6446, \9122_9421 );
and \U$10653 ( \19483_19782 , RIe20cac0_4434, \9124_9423 );
and \U$10654 ( \19484_19783 , RIe209dc0_4402, \9126_9425 );
and \U$10655 ( \19485_19784 , RIe2070c0_4370, \9128_9427 );
and \U$10656 ( \19486_19785 , RIf166e20_5630, \9130_9429 );
and \U$10657 ( \19487_19786 , RIfebf6a0_8298, \9132_9431 );
and \U$10658 ( \19488_19787 , RIfebf808_8299, \9134_9433 );
and \U$10659 ( \19489_19788 , RIfebf538_8297, \9136_9435 );
and \U$10660 ( \19490_19789 , RIfc8eb80_6646, \9138_9437 );
and \U$10661 ( \19491_19790 , RIf164120_5598, \9140_9439 );
and \U$10662 ( \19492_19791 , RIfc453e0_5810, \9142_9441 );
and \U$10663 ( \19493_19792 , RIf161b28_5571, \9144_9443 );
and \U$10664 ( \19494_19793 , RIf15fc38_5549, \9146_9445 );
and \U$10665 ( \19495_19794 , RIf15dd48_5527, \9148_9447 );
and \U$10666 ( \19496_19795 , RIe1fc968_4251, \9150_9449 );
and \U$10667 ( \19497_19796 , RIe1fb888_4239, \9152_9451 );
and \U$10668 ( \19498_19797 , RIfebf3d0_8296, \9154_9453 );
and \U$10669 ( \19499_19798 , RIf15b318_5497, \9156_9455 );
and \U$10670 ( \19500_19799 , RIfca2518_6869, \9158_9457 );
and \U$10671 ( \19501_19800 , RIfc8f120_6650, \9160_9459 );
or \U$10672 ( \19502_19801 , \19438_19737 , \19439_19738 , \19440_19739 , \19441_19740 , \19442_19741 , \19443_19742 , \19444_19743 , \19445_19744 , \19446_19745 , \19447_19746 , \19448_19747 , \19449_19748 , \19450_19749 , \19451_19750 , \19452_19751 , \19453_19752 , \19454_19753 , \19455_19754 , \19456_19755 , \19457_19756 , \19458_19757 , \19459_19758 , \19460_19759 , \19461_19760 , \19462_19761 , \19463_19762 , \19464_19763 , \19465_19764 , \19466_19765 , \19467_19766 , \19468_19767 , \19469_19768 , \19470_19769 , \19471_19770 , \19472_19771 , \19473_19772 , \19474_19773 , \19475_19774 , \19476_19775 , \19477_19776 , \19478_19777 , \19479_19778 , \19480_19779 , \19481_19780 , \19482_19781 , \19483_19782 , \19484_19783 , \19485_19784 , \19486_19785 , \19487_19786 , \19488_19787 , \19489_19788 , \19490_19789 , \19491_19790 , \19492_19791 , \19493_19792 , \19494_19793 , \19495_19794 , \19496_19795 , \19497_19796 , \19498_19797 , \19499_19798 , \19500_19799 , \19501_19800 );
and \U$10673 ( \19503_19802 , RIfebfad8_8301, \9163_9462 );
and \U$10674 ( \19504_19803 , RIfebf970_8300, \9165_9464 );
and \U$10675 ( \19505_19804 , RIfc7cca0_6442, \9167_9466 );
and \U$10676 ( \19506_19805 , RIe1f9dd0_4220, \9169_9468 );
and \U$10677 ( \19507_19806 , RIfe82c50_7832, \9171_9470 );
and \U$10678 ( \19508_19807 , RIf155648_5431, \9173_9472 );
and \U$10679 ( \19509_19808 , RIfc8f288_6651, \9175_9474 );
and \U$10680 ( \19510_19809 , RIe1f4f10_4164, \9177_9476 );
and \U$10681 ( \19511_19810 , RIf152d80_5402, \9179_9478 );
and \U$10682 ( \19512_19811 , RIfc8f828_6655, \9181_9480 );
and \U$10683 ( \19513_19812 , RIfcb3b88_7067, \9183_9482 );
and \U$10684 ( \19514_19813 , RIe1f2d50_4140, \9185_9484 );
and \U$10685 ( \19515_19814 , RIfc445d0_5800, \9187_9486 );
and \U$10686 ( \19516_19815 , RIfc8faf8_6657, \9189_9488 );
and \U$10687 ( \19517_19816 , RIf14da88_5343, \9191_9490 );
and \U$10688 ( \19518_19817 , RIe1eda58_4081, \9193_9492 );
and \U$10689 ( \19519_19818 , RIe1eb028_4051, \9195_9494 );
and \U$10690 ( \19520_19819 , RIe1e8328_4019, \9197_9496 );
and \U$10691 ( \19521_19820 , RIe1e5628_3987, \9199_9498 );
and \U$10692 ( \19522_19821 , RIe1e2928_3955, \9201_9500 );
and \U$10693 ( \19523_19822 , RIe1dfc28_3923, \9203_9502 );
and \U$10694 ( \19524_19823 , RIe1dcf28_3891, \9205_9504 );
and \U$10695 ( \19525_19824 , RIe1da228_3859, \9207_9506 );
and \U$10696 ( \19526_19825 , RIe1d7528_3827, \9209_9508 );
and \U$10697 ( \19527_19826 , RIe1d1b28_3763, \9211_9510 );
and \U$10698 ( \19528_19827 , RIe1cee28_3731, \9213_9512 );
and \U$10699 ( \19529_19828 , RIe1cc128_3699, \9215_9514 );
and \U$10700 ( \19530_19829 , RIe1c9428_3667, \9217_9516 );
and \U$10701 ( \19531_19830 , RIe1c6728_3635, \9219_9518 );
and \U$10702 ( \19532_19831 , RIe1c3a28_3603, \9221_9520 );
and \U$10703 ( \19533_19832 , RIe1c0d28_3571, \9223_9522 );
and \U$10704 ( \19534_19833 , RIe1be028_3539, \9225_9524 );
and \U$10705 ( \19535_19834 , RIfc7bff8_6433, \9227_9526 );
and \U$10706 ( \19536_19835 , RIfc44030_5796, \9229_9528 );
and \U$10707 ( \19537_19836 , RIe1b9000_3482, \9231_9530 );
and \U$10708 ( \19538_19837 , RIe1b6fa8_3459, \9233_9532 );
and \U$10709 ( \19539_19838 , RIfcbdd40_7182, \9235_9534 );
and \U$10710 ( \19540_19839 , RIfc8ff30_6660, \9237_9536 );
and \U$10711 ( \19541_19840 , RIe1b50b8_3437, \9239_9538 );
and \U$10712 ( \19542_19841 , RIe1b3d08_3423, \9241_9540 );
and \U$10713 ( \19543_19842 , RIfcbe178_7185, \9243_9542 );
and \U$10714 ( \19544_19843 , RIfc43d60_5794, \9245_9544 );
and \U$10715 ( \19545_19844 , RIe1b2520_3406, \9247_9546 );
and \U$10716 ( \19546_19845 , RIe1b0798_3385, \9249_9548 );
and \U$10717 ( \19547_19846 , RIfcdb5c0_7518, \9251_9550 );
and \U$10718 ( \19548_19847 , RIfc7ba58_6429, \9253_9552 );
and \U$10719 ( \19549_19848 , RIe1ac148_3335, \9255_9554 );
and \U$10720 ( \19550_19849 , RIe1aa960_3318, \9257_9556 );
and \U$10721 ( \19551_19850 , RIe1a8368_3291, \9259_9558 );
and \U$10722 ( \19552_19851 , RIe1a5668_3259, \9261_9560 );
and \U$10723 ( \19553_19852 , RIe1a2968_3227, \9263_9562 );
and \U$10724 ( \19554_19853 , RIe19fc68_3195, \9265_9564 );
and \U$10725 ( \19555_19854 , RIe18c168_2971, \9267_9566 );
and \U$10726 ( \19556_19855 , RIe178668_2747, \9269_9568 );
and \U$10727 ( \19557_19856 , RIe225fc0_4722, \9271_9570 );
and \U$10728 ( \19558_19857 , RIe21abc0_4594, \9273_9572 );
and \U$10729 ( \19559_19858 , RIe2043c0_4338, \9275_9574 );
and \U$10730 ( \19560_19859 , RIe1fe420_4270, \9277_9576 );
and \U$10731 ( \19561_19860 , RIe1f77d8_4193, \9279_9578 );
and \U$10732 ( \19562_19861 , RIe1f0320_4110, \9281_9580 );
and \U$10733 ( \19563_19862 , RIe1d4828_3795, \9283_9582 );
and \U$10734 ( \19564_19863 , RIe1bb328_3507, \9285_9584 );
and \U$10735 ( \19565_19864 , RIe1ae1a0_3358, \9287_9586 );
and \U$10736 ( \19566_19865 , RIe1707d8_2657, \9289_9588 );
or \U$10737 ( \19567_19866 , \19503_19802 , \19504_19803 , \19505_19804 , \19506_19805 , \19507_19806 , \19508_19807 , \19509_19808 , \19510_19809 , \19511_19810 , \19512_19811 , \19513_19812 , \19514_19813 , \19515_19814 , \19516_19815 , \19517_19816 , \19518_19817 , \19519_19818 , \19520_19819 , \19521_19820 , \19522_19821 , \19523_19822 , \19524_19823 , \19525_19824 , \19526_19825 , \19527_19826 , \19528_19827 , \19529_19828 , \19530_19829 , \19531_19830 , \19532_19831 , \19533_19832 , \19534_19833 , \19535_19834 , \19536_19835 , \19537_19836 , \19538_19837 , \19539_19838 , \19540_19839 , \19541_19840 , \19542_19841 , \19543_19842 , \19544_19843 , \19545_19844 , \19546_19845 , \19547_19846 , \19548_19847 , \19549_19848 , \19550_19849 , \19551_19850 , \19552_19851 , \19553_19852 , \19554_19853 , \19555_19854 , \19556_19855 , \19557_19856 , \19558_19857 , \19559_19858 , \19560_19859 , \19561_19860 , \19562_19861 , \19563_19862 , \19564_19863 , \19565_19864 , \19566_19865 );
or \U$10738 ( \19568_19867 , \19502_19801 , \19567_19866 );
_DC \g3aa8/U$1 ( \19569 , \19568_19867 , \9298_9597 );
buf \U$10739 ( \19570_19869 , \19569 );
xor \U$10740 ( \19571_19870 , \19437_19736 , \19570_19869 );
and \U$10741 ( \19572_19871 , RIdec4b68_702, \8760_9059 );
and \U$10742 ( \19573_19872 , RIdec1e68_670, \8762_9061 );
and \U$10743 ( \19574_19873 , RIfc5df08_6091, \8764_9063 );
and \U$10744 ( \19575_19874 , RIdebf168_638, \8766_9065 );
and \U$10745 ( \19576_19875 , RIfce6df8_7649, \8768_9067 );
and \U$10746 ( \19577_19876 , RIdebc468_606, \8770_9069 );
and \U$10747 ( \19578_19877 , RIdeb9768_574, \8772_9071 );
and \U$10748 ( \19579_19878 , RIdeb6a68_542, \8774_9073 );
and \U$10749 ( \19580_19879 , RIfc75ef0_6364, \8776_9075 );
and \U$10750 ( \19581_19880 , RIdeb1068_478, \8778_9077 );
and \U$10751 ( \19582_19881 , RIfcc12b0_7220, \8780_9079 );
and \U$10752 ( \19583_19882 , RIdeae368_446, \8782_9081 );
and \U$10753 ( \19584_19883 , RIfc5e340_6094, \8784_9083 );
and \U$10754 ( \19585_19884 , RIdea9070_414, \8786_9085 );
and \U$10755 ( \19586_19885 , RIdea2770_382, \8788_9087 );
and \U$10756 ( \19587_19886 , RIde9be70_350, \8790_9089 );
and \U$10757 ( \19588_19887 , RIfced4a0_7722, \8792_9091 );
and \U$10758 ( \19589_19888 , RIfcc1418_7221, \8794_9093 );
and \U$10759 ( \19590_19889 , RIfc95930_6724, \8796_9095 );
and \U$10760 ( \19591_19890 , RIfcec0f0_7708, \8798_9097 );
and \U$10761 ( \19592_19891 , RIde90368_293, \8800_9099 );
and \U$10762 ( \19593_19892 , RIde8c858_275, \8802_9101 );
and \U$10763 ( \19594_19893 , RIde893d8_259, \8804_9103 );
and \U$10764 ( \19595_19894 , RIde84ef0_238, \8806_9105 );
and \U$10765 ( \19596_19895 , RIde80d50_218, \8808_9107 );
and \U$10766 ( \19597_19896 , RIfc95a98_6725, \8810_9109 );
and \U$10767 ( \19598_19897 , RIfced068_7719, \8812_9111 );
and \U$10768 ( \19599_19898 , RIfced1d0_7720, \8814_9113 );
and \U$10769 ( \19600_19899 , RIfcedfe0_7730, \8816_9115 );
and \U$10770 ( \19601_19900 , RIe16b0a8_2595, \8818_9117 );
and \U$10771 ( \19602_19901 , RIe169758_2577, \8820_9119 );
and \U$10772 ( \19603_19902 , RIe167700_2554, \8822_9121 );
and \U$10773 ( \19604_19903 , RIe164b68_2523, \8824_9123 );
and \U$10774 ( \19605_19904 , RIe161e68_2491, \8826_9125 );
and \U$10775 ( \19606_19905 , RIee36e20_5083, \8828_9127 );
and \U$10776 ( \19607_19906 , RIe15f168_2459, \8830_9129 );
and \U$10777 ( \19608_19907 , RIfc426e0_5778, \8832_9131 );
and \U$10778 ( \19609_19908 , RIe15c468_2427, \8834_9133 );
and \U$10779 ( \19610_19909 , RIe156a68_2363, \8836_9135 );
and \U$10780 ( \19611_19910 , RIe153d68_2331, \8838_9137 );
and \U$10781 ( \19612_19911 , RIfe82818_7829, \8840_9139 );
and \U$10782 ( \19613_19912 , RIe151068_2299, \8842_9141 );
and \U$10783 ( \19614_19913 , RIee34c60_5059, \8844_9143 );
and \U$10784 ( \19615_19914 , RIe14e368_2267, \8846_9145 );
and \U$10785 ( \19616_19915 , RIfc5f9c0_6110, \8848_9147 );
and \U$10786 ( \19617_19916 , RIe14b668_2235, \8850_9149 );
and \U$10787 ( \19618_19917 , RIe148968_2203, \8852_9151 );
and \U$10788 ( \19619_19918 , RIe145c68_2171, \8854_9153 );
and \U$10789 ( \19620_19919 , RIfccfef0_7388, \8856_9155 );
and \U$10790 ( \19621_19920 , RIfca57b8_6905, \8858_9157 );
and \U$10791 ( \19622_19921 , RIfc600c8_6115, \8860_9159 );
and \U$10792 ( \19623_19922 , RIfcafda8_7023, \8862_9161 );
and \U$10793 ( \19624_19923 , RIe140970_2112, \8864_9163 );
and \U$10794 ( \19625_19924 , RIdf3e710_2087, \8866_9165 );
and \U$10795 ( \19626_19925 , RIdf3c6b8_2064, \8868_9167 );
and \U$10796 ( \19627_19926 , RIdf3a228_2038, \8870_9169 );
and \U$10797 ( \19628_19927 , RIfc5fc90_6112, \8872_9171 );
and \U$10798 ( \19629_19928 , RIee2f3c8_4996, \8874_9173 );
and \U$10799 ( \19630_19929 , RIfc742d0_6344, \8876_9175 );
and \U$10800 ( \19631_19930 , RIee2d208_4972, \8878_9177 );
and \U$10801 ( \19632_19931 , RIdf34f30_1979, \8880_9179 );
and \U$10802 ( \19633_19932 , RIfebf100_8294, \8882_9181 );
and \U$10803 ( \19634_19933 , RIdf30a48_1930, \8884_9183 );
and \U$10804 ( \19635_19934 , RIdf2ecc0_1909, \8886_9185 );
or \U$10805 ( \19636_19935 , \19572_19871 , \19573_19872 , \19574_19873 , \19575_19874 , \19576_19875 , \19577_19876 , \19578_19877 , \19579_19878 , \19580_19879 , \19581_19880 , \19582_19881 , \19583_19882 , \19584_19883 , \19585_19884 , \19586_19885 , \19587_19886 , \19588_19887 , \19589_19888 , \19590_19889 , \19591_19890 , \19592_19891 , \19593_19892 , \19594_19893 , \19595_19894 , \19596_19895 , \19597_19896 , \19598_19897 , \19599_19898 , \19600_19899 , \19601_19900 , \19602_19901 , \19603_19902 , \19604_19903 , \19605_19904 , \19606_19905 , \19607_19906 , \19608_19907 , \19609_19908 , \19610_19909 , \19611_19910 , \19612_19911 , \19613_19912 , \19614_19913 , \19615_19914 , \19616_19915 , \19617_19916 , \19618_19917 , \19619_19918 , \19620_19919 , \19621_19920 , \19622_19921 , \19623_19922 , \19624_19923 , \19625_19924 , \19626_19925 , \19627_19926 , \19628_19927 , \19629_19928 , \19630_19929 , \19631_19930 , \19632_19931 , \19633_19932 , \19634_19933 , \19635_19934 );
and \U$10806 ( \19637_19936 , RIfcb08e8_7031, \8889_9188 );
and \U$10807 ( \19638_19937 , RIfcee418_7733, \8891_9190 );
and \U$10808 ( \19639_19938 , RIfc95ed0_6728, \8893_9192 );
and \U$10809 ( \19640_19939 , RIfcdef68_7559, \8895_9194 );
and \U$10810 ( \19641_19940 , RIdf29e00_1853, \8897_9196 );
and \U$10811 ( \19642_19941 , RIdf27c40_1829, \8899_9198 );
and \U$10812 ( \19643_19942 , RIdf25eb8_1808, \8901_9200 );
and \U$10813 ( \19644_19943 , RIdf24298_1788, \8903_9202 );
and \U$10814 ( \19645_19944 , RIfc5ed18_6101, \8905_9204 );
and \U$10815 ( \19646_19945 , RIfcee850_7736, \8907_9206 );
and \U$10816 ( \19647_19946 , RIdf227e0_1769, \8909_9208 );
and \U$10817 ( \19648_19947 , RIfc5efe8_6103, \8911_9210 );
and \U$10818 ( \19649_19948 , RIdf212c8_1754, \8913_9212 );
and \U$10819 ( \19650_19949 , RIfeaa520_8254, \8915_9214 );
and \U$10820 ( \19651_19950 , RIdf1ad88_1682, \8917_9216 );
and \U$10821 ( \19652_19951 , RIdf18e98_1660, \8919_9218 );
and \U$10822 ( \19653_19952 , RIdf16738_1632, \8921_9220 );
and \U$10823 ( \19654_19953 , RIdf13a38_1600, \8923_9222 );
and \U$10824 ( \19655_19954 , RIdf10d38_1568, \8925_9224 );
and \U$10825 ( \19656_19955 , RIdf0e038_1536, \8927_9226 );
and \U$10826 ( \19657_19956 , RIdf0b338_1504, \8929_9228 );
and \U$10827 ( \19658_19957 , RIdf08638_1472, \8931_9230 );
and \U$10828 ( \19659_19958 , RIdf05938_1440, \8933_9232 );
and \U$10829 ( \19660_19959 , RIdf02c38_1408, \8935_9234 );
and \U$10830 ( \19661_19960 , RIdefd238_1344, \8937_9236 );
and \U$10831 ( \19662_19961 , RIdefa538_1312, \8939_9238 );
and \U$10832 ( \19663_19962 , RIdef7838_1280, \8941_9240 );
and \U$10833 ( \19664_19963 , RIdef4b38_1248, \8943_9242 );
and \U$10834 ( \19665_19964 , RIdef1e38_1216, \8945_9244 );
and \U$10835 ( \19666_19965 , RIdeef138_1184, \8947_9246 );
and \U$10836 ( \19667_19966 , RIdeec438_1152, \8949_9248 );
and \U$10837 ( \19668_19967 , RIdee9738_1120, \8951_9250 );
and \U$10838 ( \19669_19968 , RIfcc96e0_7314, \8953_9252 );
and \U$10839 ( \19670_19969 , RIfccfd88_7387, \8955_9254 );
and \U$10840 ( \19671_19970 , RIfc60aa0_6122, \8957_9256 );
and \U$10841 ( \19672_19971 , RIfca5ec0_6910, \8959_9258 );
and \U$10842 ( \19673_19972 , RIdee45a8_1062, \8961_9260 );
and \U$10843 ( \19674_19973 , RIdee2550_1039, \8963_9262 );
and \U$10844 ( \19675_19974 , RIdee0660_1017, \8965_9264 );
and \U$10845 ( \19676_19975 , RIfe826b0_7828, \8967_9266 );
and \U$10846 ( \19677_19976 , RIfcdeb30_7556, \8969_9268 );
and \U$10847 ( \19678_19977 , RIfc73bc8_6339, \8971_9270 );
and \U$10848 ( \19679_19978 , RIfca5bf0_6908, \8973_9272 );
and \U$10849 ( \19680_19979 , RIfc73a60_6338, \8975_9274 );
and \U$10850 ( \19681_19980 , RIfe82980_7830, \8977_9276 );
and \U$10851 ( \19682_19981 , RIded6bb0_907, \8979_9278 );
and \U$10852 ( \19683_19982 , RIded4cc0_885, \8981_9280 );
and \U$10853 ( \19684_19983 , RIded2830_859, \8983_9282 );
and \U$10854 ( \19685_19984 , RIdecff68_830, \8985_9284 );
and \U$10855 ( \19686_19985 , RIdecd268_798, \8987_9286 );
and \U$10856 ( \19687_19986 , RIdeca568_766, \8989_9288 );
and \U$10857 ( \19688_19987 , RIdec7868_734, \8991_9290 );
and \U$10858 ( \19689_19988 , RIdeb3d68_510, \8993_9292 );
and \U$10859 ( \19690_19989 , RIde95570_318, \8995_9294 );
and \U$10860 ( \19691_19990 , RIe16d970_2624, \8997_9296 );
and \U$10861 ( \19692_19991 , RIe159768_2395, \8999_9298 );
and \U$10862 ( \19693_19992 , RIe142f68_2139, \9001_9300 );
and \U$10863 ( \19694_19993 , RIdf37960_2009, \9003_9302 );
and \U$10864 ( \19695_19994 , RIdf2bfc0_1877, \9005_9304 );
and \U$10865 ( \19696_19995 , RIdf1c840_1701, \9007_9306 );
and \U$10866 ( \19697_19996 , RIdefff38_1376, \9009_9308 );
and \U$10867 ( \19698_19997 , RIdee6a38_1088, \9011_9310 );
and \U$10868 ( \19699_19998 , RIdedb7a0_961, \9013_9312 );
and \U$10869 ( \19700_19999 , RIde7b4b8_191, \9015_9314 );
or \U$10870 ( \19701_20000 , \19637_19936 , \19638_19937 , \19639_19938 , \19640_19939 , \19641_19940 , \19642_19941 , \19643_19942 , \19644_19943 , \19645_19944 , \19646_19945 , \19647_19946 , \19648_19947 , \19649_19948 , \19650_19949 , \19651_19950 , \19652_19951 , \19653_19952 , \19654_19953 , \19655_19954 , \19656_19955 , \19657_19956 , \19658_19957 , \19659_19958 , \19660_19959 , \19661_19960 , \19662_19961 , \19663_19962 , \19664_19963 , \19665_19964 , \19666_19965 , \19667_19966 , \19668_19967 , \19669_19968 , \19670_19969 , \19671_19970 , \19672_19971 , \19673_19972 , \19674_19973 , \19675_19974 , \19676_19975 , \19677_19976 , \19678_19977 , \19679_19978 , \19680_19979 , \19681_19980 , \19682_19981 , \19683_19982 , \19684_19983 , \19685_19984 , \19686_19985 , \19687_19986 , \19688_19987 , \19689_19988 , \19690_19989 , \19691_19990 , \19692_19991 , \19693_19992 , \19694_19993 , \19695_19994 , \19696_19995 , \19697_19996 , \19698_19997 , \19699_19998 , \19700_19999 );
or \U$10871 ( \19702_20001 , \19636_19935 , \19701_20000 );
_DC \g2a00/U$1 ( \19703 , \19702_20001 , \9024_9323 );
buf \U$10872 ( \19704_20003 , \19703 );
and \U$10873 ( \19705_20004 , RIe19ce00_3162, \9034_9333 );
and \U$10874 ( \19706_20005 , RIe19a100_3130, \9036_9335 );
and \U$10875 ( \19707_20006 , RIfce96c0_7678, \9038_9337 );
and \U$10876 ( \19708_20007 , RIe197400_3098, \9040_9339 );
and \U$10877 ( \19709_20008 , RIf144410_5236, \9042_9341 );
and \U$10878 ( \19710_20009 , RIe194700_3066, \9044_9343 );
and \U$10879 ( \19711_20010 , RIe191a00_3034, \9046_9345 );
and \U$10880 ( \19712_20011 , RIe18ed00_3002, \9048_9347 );
and \U$10881 ( \19713_20012 , RIe189300_2938, \9050_9349 );
and \U$10882 ( \19714_20013 , RIe186600_2906, \9052_9351 );
and \U$10883 ( \19715_20014 , RIfebee30_8292, \9054_9353 );
and \U$10884 ( \19716_20015 , RIe183900_2874, \9056_9355 );
and \U$10885 ( \19717_20016 , RIfcdbcc8_7523, \9058_9357 );
and \U$10886 ( \19718_20017 , RIe180c00_2842, \9060_9359 );
and \U$10887 ( \19719_20018 , RIe17df00_2810, \9062_9361 );
and \U$10888 ( \19720_20019 , RIe17b200_2778, \9064_9363 );
and \U$10889 ( \19721_20020 , RIf141f80_5210, \9066_9365 );
and \U$10890 ( \19722_20021 , RIfce7398_7653, \9068_9367 );
and \U$10891 ( \19723_20022 , RIfcb1e00_7046, \9070_9369 );
and \U$10892 ( \19724_20023 , RIfe82548_7827, \9072_9371 );
and \U$10893 ( \19725_20024 , RIfca42a0_6890, \9074_9373 );
and \U$10894 ( \19726_20025 , RIfcbff00_7206, \9076_9375 );
and \U$10895 ( \19727_20026 , RIfcaaee8_6967, \9078_9377 );
and \U$10896 ( \19728_20027 , RIee3d090_5153, \9080_9379 );
and \U$10897 ( \19729_20028 , RIfc5c180_6070, \9082_9381 );
and \U$10898 ( \19730_20029 , RIfce35b8_7609, \9084_9383 );
and \U$10899 ( \19731_20030 , RIee399b8_5114, \9086_9385 );
and \U$10900 ( \19732_20031 , RIfea8a68_8235, \9088_9387 );
and \U$10901 ( \19733_20032 , RIf16fef8_5733, \9090_9389 );
and \U$10902 ( \19734_20033 , RIfebecc8_8291, \9092_9391 );
and \U$10903 ( \19735_20034 , RIfc5c450_6072, \9094_9393 );
and \U$10904 ( \19736_20035 , RIfce9288_7675, \9096_9395 );
and \U$10905 ( \19737_20036 , RIfc40778_5759, \9098_9397 );
and \U$10906 ( \19738_20037 , RIe223158_4689, \9100_9399 );
and \U$10907 ( \19739_20038 , RIfce77d0_7656, \9102_9401 );
and \U$10908 ( \19740_20039 , RIe220458_4657, \9104_9403 );
and \U$10909 ( \19741_20040 , RIfce24d8_7597, \9106_9405 );
and \U$10910 ( \19742_20041 , RIe21d758_4625, \9108_9407 );
and \U$10911 ( \19743_20042 , RIe217d58_4561, \9110_9409 );
and \U$10912 ( \19744_20043 , RIe215058_4529, \9112_9411 );
and \U$10913 ( \19745_20044 , RIfce8a18_7669, \9114_9413 );
and \U$10914 ( \19746_20045 , RIe212358_4497, \9116_9415 );
and \U$10915 ( \19747_20046 , RIfce1998_7589, \9118_9417 );
and \U$10916 ( \19748_20047 , RIe20f658_4465, \9120_9419 );
and \U$10917 ( \19749_20048 , RIfc77840_6382, \9122_9421 );
and \U$10918 ( \19750_20049 , RIe20c958_4433, \9124_9423 );
and \U$10919 ( \19751_20050 , RIe209c58_4401, \9126_9425 );
and \U$10920 ( \19752_20051 , RIe206f58_4369, \9128_9427 );
and \U$10921 ( \19753_20052 , RIf166cb8_5629, \9130_9429 );
and \U$10922 ( \19754_20053 , RIf165bd8_5617, \9132_9431 );
and \U$10923 ( \19755_20054 , RIfe81fa8_7823, \9134_9433 );
and \U$10924 ( \19756_20055 , RIfe81e40_7822, \9136_9435 );
and \U$10925 ( \19757_20056 , RIfc5c888_6075, \9138_9437 );
and \U$10926 ( \19758_20057 , RIfceb178_7697, \9140_9439 );
and \U$10927 ( \19759_20058 , RIf1631a8_5587, \9142_9441 );
and \U$10928 ( \19760_20059 , RIf1619c0_5570, \9144_9443 );
and \U$10929 ( \19761_20060 , RIfccf248_7379, \9146_9445 );
and \U$10930 ( \19762_20061 , RIfc77570_6380, \9148_9447 );
and \U$10931 ( \19763_20062 , RIe1fc800_4250, \9150_9449 );
and \U$10932 ( \19764_20063 , RIe1fb720_4238, \9152_9451 );
and \U$10933 ( \19765_20064 , RIf15c830_5512, \9154_9453 );
and \U$10934 ( \19766_20065 , RIf15b1b0_5496, \9156_9455 );
and \U$10935 ( \19767_20066 , RIfcd0fd0_7400, \9158_9457 );
and \U$10936 ( \19768_20067 , RIfccc6b0_7348, \9160_9459 );
or \U$10937 ( \19769_20068 , \19705_20004 , \19706_20005 , \19707_20006 , \19708_20007 , \19709_20008 , \19710_20009 , \19711_20010 , \19712_20011 , \19713_20012 , \19714_20013 , \19715_20014 , \19716_20015 , \19717_20016 , \19718_20017 , \19719_20018 , \19720_20019 , \19721_20020 , \19722_20021 , \19723_20022 , \19724_20023 , \19725_20024 , \19726_20025 , \19727_20026 , \19728_20027 , \19729_20028 , \19730_20029 , \19731_20030 , \19732_20031 , \19733_20032 , \19734_20033 , \19735_20034 , \19736_20035 , \19737_20036 , \19738_20037 , \19739_20038 , \19740_20039 , \19741_20040 , \19742_20041 , \19743_20042 , \19744_20043 , \19745_20044 , \19746_20045 , \19747_20046 , \19748_20047 , \19749_20048 , \19750_20049 , \19751_20050 , \19752_20051 , \19753_20052 , \19754_20053 , \19755_20054 , \19756_20055 , \19757_20056 , \19758_20057 , \19759_20058 , \19760_20059 , \19761_20060 , \19762_20061 , \19763_20062 , \19764_20063 , \19765_20064 , \19766_20065 , \19767_20066 , \19768_20067 );
and \U$10938 ( \19770_20069 , RIf158bb8_5469, \9163_9462 );
and \U$10939 ( \19771_20070 , RIf157808_5455, \9165_9464 );
and \U$10940 ( \19772_20071 , RIfc5d0f8_6081, \9167_9466 );
and \U$10941 ( \19773_20072 , RIfebef98_8293, \9169_9468 );
and \U$10942 ( \19774_20073 , RIfcc8a38_7305, \9171_9470 );
and \U$10943 ( \19775_20074 , RIfcd7ab0_7476, \9173_9472 );
and \U$10944 ( \19776_20075 , RIfcb1428_7039, \9175_9474 );
and \U$10945 ( \19777_20076 , RIfeaa0e8_8251, \9177_9476 );
and \U$10946 ( \19778_20077 , RIfccc548_7347, \9179_9478 );
and \U$10947 ( \19779_20078 , RIfce3450_7608, \9181_9480 );
and \U$10948 ( \19780_20079 , RIf1504b8_5373, \9183_9482 );
and \U$10949 ( \19781_20080 , RIe1f2be8_4139, \9185_9484 );
and \U$10950 ( \19782_20081 , RIf14f540_5362, \9187_9486 );
and \U$10951 ( \19783_20082 , RIfc772a0_6378, \9189_9488 );
and \U$10952 ( \19784_20083 , RIfcec258_7709, \9191_9490 );
and \U$10953 ( \19785_20084 , RIe1ed8f0_4080, \9193_9492 );
and \U$10954 ( \19786_20085 , RIe1eaec0_4050, \9195_9494 );
and \U$10955 ( \19787_20086 , RIe1e81c0_4018, \9197_9496 );
and \U$10956 ( \19788_20087 , RIe1e54c0_3986, \9199_9498 );
and \U$10957 ( \19789_20088 , RIe1e27c0_3954, \9201_9500 );
and \U$10958 ( \19790_20089 , RIe1dfac0_3922, \9203_9502 );
and \U$10959 ( \19791_20090 , RIe1dcdc0_3890, \9205_9504 );
and \U$10960 ( \19792_20091 , RIe1da0c0_3858, \9207_9506 );
and \U$10961 ( \19793_20092 , RIe1d73c0_3826, \9209_9508 );
and \U$10962 ( \19794_20093 , RIe1d19c0_3762, \9211_9510 );
and \U$10963 ( \19795_20094 , RIe1cecc0_3730, \9213_9512 );
and \U$10964 ( \19796_20095 , RIe1cbfc0_3698, \9215_9514 );
and \U$10965 ( \19797_20096 , RIe1c92c0_3666, \9217_9516 );
and \U$10966 ( \19798_20097 , RIe1c65c0_3634, \9219_9518 );
and \U$10967 ( \19799_20098 , RIe1c38c0_3602, \9221_9520 );
and \U$10968 ( \19800_20099 , RIe1c0bc0_3570, \9223_9522 );
and \U$10969 ( \19801_20100 , RIe1bdec0_3538, \9225_9524 );
and \U$10970 ( \19802_20101 , RIf14c570_5328, \9227_9526 );
and \U$10971 ( \19803_20102 , RIf14b328_5315, \9229_9528 );
and \U$10972 ( \19804_20103 , RIe1b8e98_3481, \9231_9530 );
and \U$10973 ( \19805_20104 , RIe1b6e40_3458, \9233_9532 );
and \U$10974 ( \19806_20105 , RIfc76760_6370, \9235_9534 );
and \U$10975 ( \19807_20106 , RIfc94b20_6714, \9237_9536 );
and \U$10976 ( \19808_20107 , RIe1b4f50_3436, \9239_9538 );
and \U$10977 ( \19809_20108 , RIe1b3ba0_3422, \9241_9540 );
and \U$10978 ( \19810_20109 , RIfcec3c0_7710, \9243_9542 );
and \U$10979 ( \19811_20110 , RIfceb010_7696, \9245_9544 );
and \U$10980 ( \19812_20111 , RIfe823e0_7826, \9247_9546 );
and \U$10981 ( \19813_20112 , RIfe82110_7824, \9249_9548 );
and \U$10982 ( \19814_20113 , RIfcdd8e8_7543, \9251_9550 );
and \U$10983 ( \19815_20114 , RIfcc0ba8_7215, \9253_9552 );
and \U$10984 ( \19816_20115 , RIfe82278_7825, \9255_9554 );
and \U$10985 ( \19817_20116 , RIe1aa7f8_3317, \9257_9556 );
and \U$10986 ( \19818_20117 , RIe1a8200_3290, \9259_9558 );
and \U$10987 ( \19819_20118 , RIe1a5500_3258, \9261_9560 );
and \U$10988 ( \19820_20119 , RIe1a2800_3226, \9263_9562 );
and \U$10989 ( \19821_20120 , RIe19fb00_3194, \9265_9564 );
and \U$10990 ( \19822_20121 , RIe18c000_2970, \9267_9566 );
and \U$10991 ( \19823_20122 , RIe178500_2746, \9269_9568 );
and \U$10992 ( \19824_20123 , RIe225e58_4721, \9271_9570 );
and \U$10993 ( \19825_20124 , RIe21aa58_4593, \9273_9572 );
and \U$10994 ( \19826_20125 , RIe204258_4337, \9275_9574 );
and \U$10995 ( \19827_20126 , RIe1fe2b8_4269, \9277_9576 );
and \U$10996 ( \19828_20127 , RIe1f7670_4192, \9279_9578 );
and \U$10997 ( \19829_20128 , RIe1f01b8_4109, \9281_9580 );
and \U$10998 ( \19830_20129 , RIe1d46c0_3794, \9283_9582 );
and \U$10999 ( \19831_20130 , RIe1bb1c0_3506, \9285_9584 );
and \U$11000 ( \19832_20131 , RIe1ae038_3357, \9287_9586 );
and \U$11001 ( \19833_20132 , RIe170670_2656, \9289_9588 );
or \U$11002 ( \19834_20133 , \19770_20069 , \19771_20070 , \19772_20071 , \19773_20072 , \19774_20073 , \19775_20074 , \19776_20075 , \19777_20076 , \19778_20077 , \19779_20078 , \19780_20079 , \19781_20080 , \19782_20081 , \19783_20082 , \19784_20083 , \19785_20084 , \19786_20085 , \19787_20086 , \19788_20087 , \19789_20088 , \19790_20089 , \19791_20090 , \19792_20091 , \19793_20092 , \19794_20093 , \19795_20094 , \19796_20095 , \19797_20096 , \19798_20097 , \19799_20098 , \19800_20099 , \19801_20100 , \19802_20101 , \19803_20102 , \19804_20103 , \19805_20104 , \19806_20105 , \19807_20106 , \19808_20107 , \19809_20108 , \19810_20109 , \19811_20110 , \19812_20111 , \19813_20112 , \19814_20113 , \19815_20114 , \19816_20115 , \19817_20116 , \19818_20117 , \19819_20118 , \19820_20119 , \19821_20120 , \19822_20121 , \19823_20122 , \19824_20123 , \19825_20124 , \19826_20125 , \19827_20126 , \19828_20127 , \19829_20128 , \19830_20129 , \19831_20130 , \19832_20131 , \19833_20132 );
or \U$11003 ( \19835_20134 , \19769_20068 , \19834_20133 );
_DC \g3b2d/U$1 ( \19836 , \19835_20134 , \9298_9597 );
buf \U$11004 ( \19837_20136 , \19836 );
and \U$11005 ( \19838_20137 , \19704_20003 , \19837_20136 );
and \U$11006 ( \19839_20138 , \17984_18283 , \18117_18416 );
and \U$11007 ( \19840_20139 , \18117_18416 , \18392_18691 );
and \U$11008 ( \19841_20140 , \17984_18283 , \18392_18691 );
or \U$11009 ( \19842_20141 , \19839_20138 , \19840_20139 , \19841_20140 );
and \U$11010 ( \19843_20142 , \19837_20136 , \19842_20141 );
and \U$11011 ( \19844_20143 , \19704_20003 , \19842_20141 );
or \U$11012 ( \19845_20144 , \19838_20137 , \19843_20142 , \19844_20143 );
xor \U$11013 ( \19846_20145 , \19571_19870 , \19845_20144 );
buf g4424_GF_PartitionCandidate( \19847_20146_nG4424 , \19846_20145 );
xor \U$11014 ( \19848_20147 , \19704_20003 , \19837_20136 );
xor \U$11015 ( \19849_20148 , \19848_20147 , \19842_20141 );
buf g4427_GF_PartitionCandidate( \19850_20149_nG4427 , \19849_20148 );
nand \U$11016 ( \19851_20150 , \19850_20149_nG4427 , \18394_18693_nG442a );
and \U$11017 ( \19852_20151 , \19847_20146_nG4424 , \19851_20150 );
xor \U$11018 ( \19853_20152 , \19850_20149_nG4427 , \18394_18693_nG442a );
and \U$11023 ( \19854_20156 , \19853_20152 , \10392_10694_nG9c0e );
or \U$11024 ( \19855_20157 , 1'b0 , \19854_20156 );
xor \U$11025 ( \19856_20158 , \19852_20151 , \19855_20157 );
xor \U$11026 ( \19857_20159 , \19852_20151 , \19856_20158 );
buf \U$11027 ( \19858_20160 , \19857_20159 );
buf \U$11028 ( \19859_20161 , \19858_20160 );
and \U$11029 ( \19860_20162 , \19304_19603 , \19859_20161 );
and \U$11030 ( \19861_20163 , \18847_19149 , \19296_19595 );
and \U$11031 ( \19862_20164 , \18847_19149 , \19302_19601 );
and \U$11032 ( \19863_20165 , \19296_19595 , \19302_19601 );
or \U$11033 ( \19864_20166 , \19861_20163 , \19862_20164 , \19863_20165 );
buf \U$11034 ( \19865_20167 , \19864_20166 );
and \U$11035 ( \19866_20168 , \18852_19154 , \18883_19185 );
and \U$11036 ( \19867_20169 , \18852_19154 , \19294_19593 );
and \U$11037 ( \19868_20170 , \18883_19185 , \19294_19593 );
or \U$11038 ( \19869_20171 , \19866_20168 , \19867_20169 , \19868_20170 );
buf \U$11039 ( \19870_20172 , \19869_20171 );
xor \U$11040 ( \19871_20173 , \19865_20167 , \19870_20172 );
and \U$11041 ( \19872_20174 , \18889_19191 , \18932_19231 );
and \U$11042 ( \19873_20175 , \18889_19191 , \19292_19591 );
and \U$11043 ( \19874_20176 , \18932_19231 , \19292_19591 );
or \U$11044 ( \19875_20177 , \19872_20174 , \19873_20175 , \19874_20176 );
buf \U$11045 ( \19876_20178 , \19875_20177 );
and \U$11046 ( \19877_20179 , \18857_19159 , \18874_19176 );
and \U$11047 ( \19878_20180 , \18857_19159 , \18881_19183 );
and \U$11048 ( \19879_20181 , \18874_19176 , \18881_19183 );
or \U$11049 ( \19880_20182 , \19877_20179 , \19878_20180 , \19879_20181 );
buf \U$11050 ( \19881_20183 , \19880_20182 );
and \U$11051 ( \19882_20184 , \18859_19161 , \18865_19167 );
and \U$11052 ( \19883_20185 , \18859_19161 , \18872_19174 );
and \U$11053 ( \19884_20186 , \18865_19167 , \18872_19174 );
or \U$11054 ( \19885_20187 , \19882_20184 , \19883_20185 , \19884_20186 );
buf \U$11055 ( \19886_20188 , \19885_20187 );
and \U$11056 ( \19887_20189 , \18897_19199 , \18903_19205 );
buf \U$11057 ( \19888_20190 , \19887_20189 );
and \U$11058 ( \19889_20191 , \18908_18702 , \10693_10995_nG9c0b );
and \U$11059 ( \19890_20192 , \18400_18699 , \10981_11283_nG9c08 );
or \U$11060 ( \19891_20193 , \19889_20191 , \19890_20192 );
xor \U$11061 ( \19892_20194 , \18399_18698 , \19891_20193 );
buf \U$11062 ( \19893_20195 , \19892_20194 );
buf \U$11064 ( \19894_20196 , \19893_20195 );
and \U$11065 ( \19895_20197 , \17437_17297 , \11299_11598_nG9c05 );
and \U$11066 ( \19896_20198 , \16995_17294 , \12168_12470_nG9c02 );
or \U$11067 ( \19897_20199 , \19895_20197 , \19896_20198 );
xor \U$11068 ( \19898_20200 , \16994_17293 , \19897_20199 );
buf \U$11069 ( \19899_20201 , \19898_20200 );
buf \U$11071 ( \19900_20202 , \19899_20201 );
xor \U$11072 ( \19901_20203 , \19894_20196 , \19900_20202 );
buf \U$11073 ( \19902_20204 , \19901_20203 );
xor \U$11074 ( \19903_20205 , \19888_20190 , \19902_20204 );
and \U$11075 ( \19904_20206 , \16405_15940 , \12502_12801_nG9bff );
and \U$11076 ( \19905_20207 , \15638_15937 , \13403_13705_nG9bfc );
or \U$11077 ( \19906_20208 , \19904_20206 , \19905_20207 );
xor \U$11078 ( \19907_20209 , \15637_15936 , \19906_20208 );
buf \U$11079 ( \19908_20210 , \19907_20209 );
buf \U$11081 ( \19909_20211 , \19908_20210 );
xor \U$11082 ( \19910_20212 , \19903_20205 , \19909_20211 );
buf \U$11083 ( \19911_20213 , \19910_20212 );
xor \U$11084 ( \19912_20214 , \19886_20188 , \19911_20213 );
and \U$11085 ( \19913_20215 , \12183_12157 , \16378_16680_nG9bed );
and \U$11086 ( \19914_20216 , \11855_12154 , \17363_17665_nG9bea );
or \U$11087 ( \19915_20217 , \19913_20215 , \19914_20216 );
xor \U$11088 ( \19916_20218 , \11854_12153 , \19915_20217 );
buf \U$11089 ( \19917_20219 , \19916_20218 );
buf \U$11091 ( \19918_20220 , \19917_20219 );
xor \U$11092 ( \19919_20221 , \19912_20214 , \19918_20220 );
buf \U$11093 ( \19920_20222 , \19919_20221 );
xor \U$11094 ( \19921_20223 , \19881_20183 , \19920_20222 );
and \U$11095 ( \19922_20224 , \18894_19196 , \18923_19222 );
and \U$11096 ( \19923_20225 , \18894_19196 , \18930_19229 );
and \U$11097 ( \19924_20226 , \18923_19222 , \18930_19229 );
or \U$11098 ( \19925_20227 , \19922_20224 , \19923_20225 , \19924_20226 );
buf \U$11099 ( \19926_20228 , \19925_20227 );
xor \U$11100 ( \19927_20229 , \19921_20223 , \19926_20228 );
buf \U$11101 ( \19928_20230 , \19927_20229 );
xor \U$11102 ( \19929_20231 , \19876_20178 , \19928_20230 );
and \U$11103 ( \19930_20232 , \18905_19207 , \18914_19213 );
and \U$11104 ( \19931_20233 , \18905_19207 , \18921_19220 );
and \U$11105 ( \19932_20234 , \18914_19213 , \18921_19220 );
or \U$11106 ( \19933_20235 , \19930_20232 , \19931_20233 , \19932_20234 );
buf \U$11107 ( \19934_20236 , \19933_20235 );
and \U$11108 ( \19935_20237 , \14710_14631 , \13771_14070_nG9bf9 );
and \U$11109 ( \19936_20238 , \14329_14628 , \14682_14984_nG9bf6 );
or \U$11110 ( \19937_20239 , \19935_20237 , \19936_20238 );
xor \U$11111 ( \19938_20240 , \14328_14627 , \19937_20239 );
buf \U$11112 ( \19939_20241 , \19938_20240 );
buf \U$11114 ( \19940_20242 , \19939_20241 );
xor \U$11115 ( \19941_20243 , \19934_20236 , \19940_20242 );
and \U$11116 ( \19942_20244 , \13431_13370 , \15074_15373_nG9bf3 );
and \U$11117 ( \19943_20245 , \13068_13367 , \16013_16315_nG9bf0 );
or \U$11118 ( \19944_20246 , \19942_20244 , \19943_20245 );
xor \U$11119 ( \19945_20247 , \13067_13366 , \19944_20246 );
buf \U$11120 ( \19946_20248 , \19945_20247 );
buf \U$11122 ( \19947_20249 , \19946_20248 );
xor \U$11123 ( \19948_20250 , \19941_20243 , \19947_20249 );
buf \U$11124 ( \19949_20251 , \19948_20250 );
and \U$11125 ( \19950_20252 , \10996_10421 , \17808_18107_nG9be7 );
and \U$11126 ( \19951_20253 , \10119_10418 , \18789_19091_nG9be4 );
or \U$11127 ( \19952_20254 , \19950_20252 , \19951_20253 );
xor \U$11128 ( \19953_20255 , \10118_10417 , \19952_20254 );
buf \U$11129 ( \19954_20256 , \19953_20255 );
buf \U$11131 ( \19955_20257 , \19954_20256 );
xor \U$11132 ( \19956_20258 , \19949_20251 , \19955_20257 );
and \U$11133 ( \19957_20259 , \10411_10707 , \19287_19586_nG9be1 );
and \U$11134 ( \19958_20260 , \19249_19548 , \19253_19552 );
and \U$11135 ( \19959_20261 , \19253_19552 , \19275_19574 );
and \U$11136 ( \19960_20262 , \19249_19548 , \19275_19574 );
or \U$11137 ( \19961_20263 , \19958_20260 , \19959_20261 , \19960_20262 );
and \U$11138 ( \19962_20264 , \15022_15321 , \13755_14054 );
and \U$11139 ( \19963_20265 , \15965_16267 , \13390_13692 );
nor \U$11140 ( \19964_20266 , \19962_20264 , \19963_20265 );
xnor \U$11141 ( \19965_20267 , \19964_20266 , \13736_14035 );
and \U$11142 ( \19966_20268 , \13725_14024 , \15037_15336 );
and \U$11143 ( \19967_20269 , \14648_14950 , \14661_14963 );
nor \U$11144 ( \19968_20270 , \19966_20268 , \19967_20269 );
xnor \U$11145 ( \19969_20271 , \19968_20270 , \15043_15342 );
xor \U$11146 ( \19970_20272 , \19965_20267 , \19969_20271 );
and \U$11147 ( \19971_20273 , \10686_10988 , \19235_19534 );
and \U$11148 ( \19972_20274 , \10968_11270 , \18743_19045 );
nor \U$11149 ( \19973_20275 , \19971_20273 , \19972_20274 );
xnor \U$11150 ( \19974_20276 , \19973_20275 , \19241_19540 );
xor \U$11151 ( \19975_20277 , \19970_20272 , \19974_20276 );
and \U$11152 ( \19976_20278 , \19259_19558 , \10681_10983 );
and \U$11153 ( \19977_20279 , RIdec4b68_702, \9034_9333 );
and \U$11154 ( \19978_20280 , RIdec1e68_670, \9036_9335 );
and \U$11155 ( \19979_20281 , RIfc5df08_6091, \9038_9337 );
and \U$11156 ( \19980_20282 , RIdebf168_638, \9040_9339 );
and \U$11157 ( \19981_20283 , RIfce6df8_7649, \9042_9341 );
and \U$11158 ( \19982_20284 , RIdebc468_606, \9044_9343 );
and \U$11159 ( \19983_20285 , RIdeb9768_574, \9046_9345 );
and \U$11160 ( \19984_20286 , RIdeb6a68_542, \9048_9347 );
and \U$11161 ( \19985_20287 , RIfc75ef0_6364, \9050_9349 );
and \U$11162 ( \19986_20288 , RIdeb1068_478, \9052_9351 );
and \U$11163 ( \19987_20289 , RIfcc12b0_7220, \9054_9353 );
and \U$11164 ( \19988_20290 , RIdeae368_446, \9056_9355 );
and \U$11165 ( \19989_20291 , RIfc5e340_6094, \9058_9357 );
and \U$11166 ( \19990_20292 , RIdea9070_414, \9060_9359 );
and \U$11167 ( \19991_20293 , RIdea2770_382, \9062_9361 );
and \U$11168 ( \19992_20294 , RIde9be70_350, \9064_9363 );
and \U$11169 ( \19993_20295 , RIfced4a0_7722, \9066_9365 );
and \U$11170 ( \19994_20296 , RIfcc1418_7221, \9068_9367 );
and \U$11171 ( \19995_20297 , RIfc95930_6724, \9070_9369 );
and \U$11172 ( \19996_20298 , RIfcec0f0_7708, \9072_9371 );
and \U$11173 ( \19997_20299 , RIde90368_293, \9074_9373 );
and \U$11174 ( \19998_20300 , RIde8c858_275, \9076_9375 );
and \U$11175 ( \19999_20301 , RIde893d8_259, \9078_9377 );
and \U$11176 ( \20000_20302 , RIde84ef0_238, \9080_9379 );
and \U$11177 ( \20001_20303 , RIde80d50_218, \9082_9381 );
and \U$11178 ( \20002_20304 , RIfc95a98_6725, \9084_9383 );
and \U$11179 ( \20003_20305 , RIfced068_7719, \9086_9385 );
and \U$11180 ( \20004_20306 , RIfced1d0_7720, \9088_9387 );
and \U$11181 ( \20005_20307 , RIfcedfe0_7730, \9090_9389 );
and \U$11182 ( \20006_20308 , RIe16b0a8_2595, \9092_9391 );
and \U$11183 ( \20007_20309 , RIe169758_2577, \9094_9393 );
and \U$11184 ( \20008_20310 , RIe167700_2554, \9096_9395 );
and \U$11185 ( \20009_20311 , RIe164b68_2523, \9098_9397 );
and \U$11186 ( \20010_20312 , RIe161e68_2491, \9100_9399 );
and \U$11187 ( \20011_20313 , RIee36e20_5083, \9102_9401 );
and \U$11188 ( \20012_20314 , RIe15f168_2459, \9104_9403 );
and \U$11189 ( \20013_20315 , RIfc426e0_5778, \9106_9405 );
and \U$11190 ( \20014_20316 , RIe15c468_2427, \9108_9407 );
and \U$11191 ( \20015_20317 , RIe156a68_2363, \9110_9409 );
and \U$11192 ( \20016_20318 , RIe153d68_2331, \9112_9411 );
and \U$11193 ( \20017_20319 , RIfe82818_7829, \9114_9413 );
and \U$11194 ( \20018_20320 , RIe151068_2299, \9116_9415 );
and \U$11195 ( \20019_20321 , RIee34c60_5059, \9118_9417 );
and \U$11196 ( \20020_20322 , RIe14e368_2267, \9120_9419 );
and \U$11197 ( \20021_20323 , RIfc5f9c0_6110, \9122_9421 );
and \U$11198 ( \20022_20324 , RIe14b668_2235, \9124_9423 );
and \U$11199 ( \20023_20325 , RIe148968_2203, \9126_9425 );
and \U$11200 ( \20024_20326 , RIe145c68_2171, \9128_9427 );
and \U$11201 ( \20025_20327 , RIfccfef0_7388, \9130_9429 );
and \U$11202 ( \20026_20328 , RIfca57b8_6905, \9132_9431 );
and \U$11203 ( \20027_20329 , RIfc600c8_6115, \9134_9433 );
and \U$11204 ( \20028_20330 , RIfcafda8_7023, \9136_9435 );
and \U$11205 ( \20029_20331 , RIe140970_2112, \9138_9437 );
and \U$11206 ( \20030_20332 , RIdf3e710_2087, \9140_9439 );
and \U$11207 ( \20031_20333 , RIdf3c6b8_2064, \9142_9441 );
and \U$11208 ( \20032_20334 , RIdf3a228_2038, \9144_9443 );
and \U$11209 ( \20033_20335 , RIfc5fc90_6112, \9146_9445 );
and \U$11210 ( \20034_20336 , RIee2f3c8_4996, \9148_9447 );
and \U$11211 ( \20035_20337 , RIfc742d0_6344, \9150_9449 );
and \U$11212 ( \20036_20338 , RIee2d208_4972, \9152_9451 );
and \U$11213 ( \20037_20339 , RIdf34f30_1979, \9154_9453 );
and \U$11214 ( \20038_20340 , RIfebf100_8294, \9156_9455 );
and \U$11215 ( \20039_20341 , RIdf30a48_1930, \9158_9457 );
and \U$11216 ( \20040_20342 , RIdf2ecc0_1909, \9160_9459 );
or \U$11217 ( \20041_20343 , \19977_20279 , \19978_20280 , \19979_20281 , \19980_20282 , \19981_20283 , \19982_20284 , \19983_20285 , \19984_20286 , \19985_20287 , \19986_20288 , \19987_20289 , \19988_20290 , \19989_20291 , \19990_20292 , \19991_20293 , \19992_20294 , \19993_20295 , \19994_20296 , \19995_20297 , \19996_20298 , \19997_20299 , \19998_20300 , \19999_20301 , \20000_20302 , \20001_20303 , \20002_20304 , \20003_20305 , \20004_20306 , \20005_20307 , \20006_20308 , \20007_20309 , \20008_20310 , \20009_20311 , \20010_20312 , \20011_20313 , \20012_20314 , \20013_20315 , \20014_20316 , \20015_20317 , \20016_20318 , \20017_20319 , \20018_20320 , \20019_20321 , \20020_20322 , \20021_20323 , \20022_20324 , \20023_20325 , \20024_20326 , \20025_20327 , \20026_20328 , \20027_20329 , \20028_20330 , \20029_20331 , \20030_20332 , \20031_20333 , \20032_20334 , \20033_20335 , \20034_20336 , \20035_20337 , \20036_20338 , \20037_20339 , \20038_20340 , \20039_20341 , \20040_20342 );
and \U$11218 ( \20042_20344 , RIfcb08e8_7031, \9163_9462 );
and \U$11219 ( \20043_20345 , RIfcee418_7733, \9165_9464 );
and \U$11220 ( \20044_20346 , RIfc95ed0_6728, \9167_9466 );
and \U$11221 ( \20045_20347 , RIfcdef68_7559, \9169_9468 );
and \U$11222 ( \20046_20348 , RIdf29e00_1853, \9171_9470 );
and \U$11223 ( \20047_20349 , RIdf27c40_1829, \9173_9472 );
and \U$11224 ( \20048_20350 , RIdf25eb8_1808, \9175_9474 );
and \U$11225 ( \20049_20351 , RIdf24298_1788, \9177_9476 );
and \U$11226 ( \20050_20352 , RIfc5ed18_6101, \9179_9478 );
and \U$11227 ( \20051_20353 , RIfcee850_7736, \9181_9480 );
and \U$11228 ( \20052_20354 , RIdf227e0_1769, \9183_9482 );
and \U$11229 ( \20053_20355 , RIfc5efe8_6103, \9185_9484 );
and \U$11230 ( \20054_20356 , RIdf212c8_1754, \9187_9486 );
and \U$11231 ( \20055_20357 , RIfeaa520_8254, \9189_9488 );
and \U$11232 ( \20056_20358 , RIdf1ad88_1682, \9191_9490 );
and \U$11233 ( \20057_20359 , RIdf18e98_1660, \9193_9492 );
and \U$11234 ( \20058_20360 , RIdf16738_1632, \9195_9494 );
and \U$11235 ( \20059_20361 , RIdf13a38_1600, \9197_9496 );
and \U$11236 ( \20060_20362 , RIdf10d38_1568, \9199_9498 );
and \U$11237 ( \20061_20363 , RIdf0e038_1536, \9201_9500 );
and \U$11238 ( \20062_20364 , RIdf0b338_1504, \9203_9502 );
and \U$11239 ( \20063_20365 , RIdf08638_1472, \9205_9504 );
and \U$11240 ( \20064_20366 , RIdf05938_1440, \9207_9506 );
and \U$11241 ( \20065_20367 , RIdf02c38_1408, \9209_9508 );
and \U$11242 ( \20066_20368 , RIdefd238_1344, \9211_9510 );
and \U$11243 ( \20067_20369 , RIdefa538_1312, \9213_9512 );
and \U$11244 ( \20068_20370 , RIdef7838_1280, \9215_9514 );
and \U$11245 ( \20069_20371 , RIdef4b38_1248, \9217_9516 );
and \U$11246 ( \20070_20372 , RIdef1e38_1216, \9219_9518 );
and \U$11247 ( \20071_20373 , RIdeef138_1184, \9221_9520 );
and \U$11248 ( \20072_20374 , RIdeec438_1152, \9223_9522 );
and \U$11249 ( \20073_20375 , RIdee9738_1120, \9225_9524 );
and \U$11250 ( \20074_20376 , RIfcc96e0_7314, \9227_9526 );
and \U$11251 ( \20075_20377 , RIfccfd88_7387, \9229_9528 );
and \U$11252 ( \20076_20378 , RIfc60aa0_6122, \9231_9530 );
and \U$11253 ( \20077_20379 , RIfca5ec0_6910, \9233_9532 );
and \U$11254 ( \20078_20380 , RIdee45a8_1062, \9235_9534 );
and \U$11255 ( \20079_20381 , RIdee2550_1039, \9237_9536 );
and \U$11256 ( \20080_20382 , RIdee0660_1017, \9239_9538 );
and \U$11257 ( \20081_20383 , RIfe826b0_7828, \9241_9540 );
and \U$11258 ( \20082_20384 , RIfcdeb30_7556, \9243_9542 );
and \U$11259 ( \20083_20385 , RIfc73bc8_6339, \9245_9544 );
and \U$11260 ( \20084_20386 , RIfca5bf0_6908, \9247_9546 );
and \U$11261 ( \20085_20387 , RIfc73a60_6338, \9249_9548 );
and \U$11262 ( \20086_20388 , RIfe82980_7830, \9251_9550 );
and \U$11263 ( \20087_20389 , RIded6bb0_907, \9253_9552 );
and \U$11264 ( \20088_20390 , RIded4cc0_885, \9255_9554 );
and \U$11265 ( \20089_20391 , RIded2830_859, \9257_9556 );
and \U$11266 ( \20090_20392 , RIdecff68_830, \9259_9558 );
and \U$11267 ( \20091_20393 , RIdecd268_798, \9261_9560 );
and \U$11268 ( \20092_20394 , RIdeca568_766, \9263_9562 );
and \U$11269 ( \20093_20395 , RIdec7868_734, \9265_9564 );
and \U$11270 ( \20094_20396 , RIdeb3d68_510, \9267_9566 );
and \U$11271 ( \20095_20397 , RIde95570_318, \9269_9568 );
and \U$11272 ( \20096_20398 , RIe16d970_2624, \9271_9570 );
and \U$11273 ( \20097_20399 , RIe159768_2395, \9273_9572 );
and \U$11274 ( \20098_20400 , RIe142f68_2139, \9275_9574 );
and \U$11275 ( \20099_20401 , RIdf37960_2009, \9277_9576 );
and \U$11276 ( \20100_20402 , RIdf2bfc0_1877, \9279_9578 );
and \U$11277 ( \20101_20403 , RIdf1c840_1701, \9281_9580 );
and \U$11278 ( \20102_20404 , RIdefff38_1376, \9283_9582 );
and \U$11279 ( \20103_20405 , RIdee6a38_1088, \9285_9584 );
and \U$11280 ( \20104_20406 , RIdedb7a0_961, \9287_9586 );
and \U$11281 ( \20105_20407 , RIde7b4b8_191, \9289_9588 );
or \U$11282 ( \20106_20408 , \20042_20344 , \20043_20345 , \20044_20346 , \20045_20347 , \20046_20348 , \20047_20349 , \20048_20350 , \20049_20351 , \20050_20352 , \20051_20353 , \20052_20354 , \20053_20355 , \20054_20356 , \20055_20357 , \20056_20358 , \20057_20359 , \20058_20360 , \20059_20361 , \20060_20362 , \20061_20363 , \20062_20364 , \20063_20365 , \20064_20366 , \20065_20367 , \20066_20368 , \20067_20369 , \20068_20370 , \20069_20371 , \20070_20372 , \20071_20373 , \20072_20374 , \20073_20375 , \20074_20376 , \20075_20377 , \20076_20378 , \20077_20379 , \20078_20380 , \20079_20381 , \20080_20382 , \20081_20383 , \20082_20384 , \20083_20385 , \20084_20386 , \20085_20387 , \20086_20388 , \20087_20389 , \20088_20390 , \20089_20391 , \20090_20392 , \20091_20393 , \20092_20394 , \20093_20395 , \20094_20396 , \20095_20397 , \20096_20398 , \20097_20399 , \20098_20400 , \20099_20401 , \20100_20402 , \20101_20403 , \20102_20404 , \20103_20405 , \20104_20406 , \20105_20407 );
or \U$11283 ( \20107_20409 , \20041_20343 , \20106_20408 );
_DC \g65a7/U$1 ( \20108 , \20107_20409 , \9298_9597 );
and \U$11284 ( \20109_20411 , RIe19ce00_3162, \8760_9059 );
and \U$11285 ( \20110_20412 , RIe19a100_3130, \8762_9061 );
and \U$11286 ( \20111_20413 , RIfce96c0_7678, \8764_9063 );
and \U$11287 ( \20112_20414 , RIe197400_3098, \8766_9065 );
and \U$11288 ( \20113_20415 , RIf144410_5236, \8768_9067 );
and \U$11289 ( \20114_20416 , RIe194700_3066, \8770_9069 );
and \U$11290 ( \20115_20417 , RIe191a00_3034, \8772_9071 );
and \U$11291 ( \20116_20418 , RIe18ed00_3002, \8774_9073 );
and \U$11292 ( \20117_20419 , RIe189300_2938, \8776_9075 );
and \U$11293 ( \20118_20420 , RIe186600_2906, \8778_9077 );
and \U$11294 ( \20119_20421 , RIfebee30_8292, \8780_9079 );
and \U$11295 ( \20120_20422 , RIe183900_2874, \8782_9081 );
and \U$11296 ( \20121_20423 , RIfcdbcc8_7523, \8784_9083 );
and \U$11297 ( \20122_20424 , RIe180c00_2842, \8786_9085 );
and \U$11298 ( \20123_20425 , RIe17df00_2810, \8788_9087 );
and \U$11299 ( \20124_20426 , RIe17b200_2778, \8790_9089 );
and \U$11300 ( \20125_20427 , RIf141f80_5210, \8792_9091 );
and \U$11301 ( \20126_20428 , RIfce7398_7653, \8794_9093 );
and \U$11302 ( \20127_20429 , RIfcb1e00_7046, \8796_9095 );
and \U$11303 ( \20128_20430 , RIfe82548_7827, \8798_9097 );
and \U$11304 ( \20129_20431 , RIfca42a0_6890, \8800_9099 );
and \U$11305 ( \20130_20432 , RIfcbff00_7206, \8802_9101 );
and \U$11306 ( \20131_20433 , RIfcaaee8_6967, \8804_9103 );
and \U$11307 ( \20132_20434 , RIee3d090_5153, \8806_9105 );
and \U$11308 ( \20133_20435 , RIfc5c180_6070, \8808_9107 );
and \U$11309 ( \20134_20436 , RIfce35b8_7609, \8810_9109 );
and \U$11310 ( \20135_20437 , RIee399b8_5114, \8812_9111 );
and \U$11311 ( \20136_20438 , RIfea8a68_8235, \8814_9113 );
and \U$11312 ( \20137_20439 , RIf16fef8_5733, \8816_9115 );
and \U$11313 ( \20138_20440 , RIfebecc8_8291, \8818_9117 );
and \U$11314 ( \20139_20441 , RIfc5c450_6072, \8820_9119 );
and \U$11315 ( \20140_20442 , RIfce9288_7675, \8822_9121 );
and \U$11316 ( \20141_20443 , RIfc40778_5759, \8824_9123 );
and \U$11317 ( \20142_20444 , RIe223158_4689, \8826_9125 );
and \U$11318 ( \20143_20445 , RIfce77d0_7656, \8828_9127 );
and \U$11319 ( \20144_20446 , RIe220458_4657, \8830_9129 );
and \U$11320 ( \20145_20447 , RIfce24d8_7597, \8832_9131 );
and \U$11321 ( \20146_20448 , RIe21d758_4625, \8834_9133 );
and \U$11322 ( \20147_20449 , RIe217d58_4561, \8836_9135 );
and \U$11323 ( \20148_20450 , RIe215058_4529, \8838_9137 );
and \U$11324 ( \20149_20451 , RIfce8a18_7669, \8840_9139 );
and \U$11325 ( \20150_20452 , RIe212358_4497, \8842_9141 );
and \U$11326 ( \20151_20453 , RIfce1998_7589, \8844_9143 );
and \U$11327 ( \20152_20454 , RIe20f658_4465, \8846_9145 );
and \U$11328 ( \20153_20455 , RIfc77840_6382, \8848_9147 );
and \U$11329 ( \20154_20456 , RIe20c958_4433, \8850_9149 );
and \U$11330 ( \20155_20457 , RIe209c58_4401, \8852_9151 );
and \U$11331 ( \20156_20458 , RIe206f58_4369, \8854_9153 );
and \U$11332 ( \20157_20459 , RIf166cb8_5629, \8856_9155 );
and \U$11333 ( \20158_20460 , RIf165bd8_5617, \8858_9157 );
and \U$11334 ( \20159_20461 , RIfe81fa8_7823, \8860_9159 );
and \U$11335 ( \20160_20462 , RIfe81e40_7822, \8862_9161 );
and \U$11336 ( \20161_20463 , RIfc5c888_6075, \8864_9163 );
and \U$11337 ( \20162_20464 , RIfceb178_7697, \8866_9165 );
and \U$11338 ( \20163_20465 , RIf1631a8_5587, \8868_9167 );
and \U$11339 ( \20164_20466 , RIf1619c0_5570, \8870_9169 );
and \U$11340 ( \20165_20467 , RIfccf248_7379, \8872_9171 );
and \U$11341 ( \20166_20468 , RIfc77570_6380, \8874_9173 );
and \U$11342 ( \20167_20469 , RIe1fc800_4250, \8876_9175 );
and \U$11343 ( \20168_20470 , RIe1fb720_4238, \8878_9177 );
and \U$11344 ( \20169_20471 , RIf15c830_5512, \8880_9179 );
and \U$11345 ( \20170_20472 , RIf15b1b0_5496, \8882_9181 );
and \U$11346 ( \20171_20473 , RIfcd0fd0_7400, \8884_9183 );
and \U$11347 ( \20172_20474 , RIfccc6b0_7348, \8886_9185 );
or \U$11348 ( \20173_20475 , \20109_20411 , \20110_20412 , \20111_20413 , \20112_20414 , \20113_20415 , \20114_20416 , \20115_20417 , \20116_20418 , \20117_20419 , \20118_20420 , \20119_20421 , \20120_20422 , \20121_20423 , \20122_20424 , \20123_20425 , \20124_20426 , \20125_20427 , \20126_20428 , \20127_20429 , \20128_20430 , \20129_20431 , \20130_20432 , \20131_20433 , \20132_20434 , \20133_20435 , \20134_20436 , \20135_20437 , \20136_20438 , \20137_20439 , \20138_20440 , \20139_20441 , \20140_20442 , \20141_20443 , \20142_20444 , \20143_20445 , \20144_20446 , \20145_20447 , \20146_20448 , \20147_20449 , \20148_20450 , \20149_20451 , \20150_20452 , \20151_20453 , \20152_20454 , \20153_20455 , \20154_20456 , \20155_20457 , \20156_20458 , \20157_20459 , \20158_20460 , \20159_20461 , \20160_20462 , \20161_20463 , \20162_20464 , \20163_20465 , \20164_20466 , \20165_20467 , \20166_20468 , \20167_20469 , \20168_20470 , \20169_20471 , \20170_20472 , \20171_20473 , \20172_20474 );
and \U$11349 ( \20174_20476 , RIf158bb8_5469, \8889_9188 );
and \U$11350 ( \20175_20477 , RIf157808_5455, \8891_9190 );
and \U$11351 ( \20176_20478 , RIfc5d0f8_6081, \8893_9192 );
and \U$11352 ( \20177_20479 , RIfebef98_8293, \8895_9194 );
and \U$11353 ( \20178_20480 , RIfcc8a38_7305, \8897_9196 );
and \U$11354 ( \20179_20481 , RIfcd7ab0_7476, \8899_9198 );
and \U$11355 ( \20180_20482 , RIfcb1428_7039, \8901_9200 );
and \U$11356 ( \20181_20483 , RIfeaa0e8_8251, \8903_9202 );
and \U$11357 ( \20182_20484 , RIfccc548_7347, \8905_9204 );
and \U$11358 ( \20183_20485 , RIfce3450_7608, \8907_9206 );
and \U$11359 ( \20184_20486 , RIf1504b8_5373, \8909_9208 );
and \U$11360 ( \20185_20487 , RIe1f2be8_4139, \8911_9210 );
and \U$11361 ( \20186_20488 , RIf14f540_5362, \8913_9212 );
and \U$11362 ( \20187_20489 , RIfc772a0_6378, \8915_9214 );
and \U$11363 ( \20188_20490 , RIfcec258_7709, \8917_9216 );
and \U$11364 ( \20189_20491 , RIe1ed8f0_4080, \8919_9218 );
and \U$11365 ( \20190_20492 , RIe1eaec0_4050, \8921_9220 );
and \U$11366 ( \20191_20493 , RIe1e81c0_4018, \8923_9222 );
and \U$11367 ( \20192_20494 , RIe1e54c0_3986, \8925_9224 );
and \U$11368 ( \20193_20495 , RIe1e27c0_3954, \8927_9226 );
and \U$11369 ( \20194_20496 , RIe1dfac0_3922, \8929_9228 );
and \U$11370 ( \20195_20497 , RIe1dcdc0_3890, \8931_9230 );
and \U$11371 ( \20196_20498 , RIe1da0c0_3858, \8933_9232 );
and \U$11372 ( \20197_20499 , RIe1d73c0_3826, \8935_9234 );
and \U$11373 ( \20198_20500 , RIe1d19c0_3762, \8937_9236 );
and \U$11374 ( \20199_20501 , RIe1cecc0_3730, \8939_9238 );
and \U$11375 ( \20200_20502 , RIe1cbfc0_3698, \8941_9240 );
and \U$11376 ( \20201_20503 , RIe1c92c0_3666, \8943_9242 );
and \U$11377 ( \20202_20504 , RIe1c65c0_3634, \8945_9244 );
and \U$11378 ( \20203_20505 , RIe1c38c0_3602, \8947_9246 );
and \U$11379 ( \20204_20506 , RIe1c0bc0_3570, \8949_9248 );
and \U$11380 ( \20205_20507 , RIe1bdec0_3538, \8951_9250 );
and \U$11381 ( \20206_20508 , RIf14c570_5328, \8953_9252 );
and \U$11382 ( \20207_20509 , RIf14b328_5315, \8955_9254 );
and \U$11383 ( \20208_20510 , RIe1b8e98_3481, \8957_9256 );
and \U$11384 ( \20209_20511 , RIe1b6e40_3458, \8959_9258 );
and \U$11385 ( \20210_20512 , RIfc76760_6370, \8961_9260 );
and \U$11386 ( \20211_20513 , RIfc94b20_6714, \8963_9262 );
and \U$11387 ( \20212_20514 , RIe1b4f50_3436, \8965_9264 );
and \U$11388 ( \20213_20515 , RIe1b3ba0_3422, \8967_9266 );
and \U$11389 ( \20214_20516 , RIfcec3c0_7710, \8969_9268 );
and \U$11390 ( \20215_20517 , RIfceb010_7696, \8971_9270 );
and \U$11391 ( \20216_20518 , RIfe823e0_7826, \8973_9272 );
and \U$11392 ( \20217_20519 , RIfe82110_7824, \8975_9274 );
and \U$11393 ( \20218_20520 , RIfcdd8e8_7543, \8977_9276 );
and \U$11394 ( \20219_20521 , RIfcc0ba8_7215, \8979_9278 );
and \U$11395 ( \20220_20522 , RIfe82278_7825, \8981_9280 );
and \U$11396 ( \20221_20523 , RIe1aa7f8_3317, \8983_9282 );
and \U$11397 ( \20222_20524 , RIe1a8200_3290, \8985_9284 );
and \U$11398 ( \20223_20525 , RIe1a5500_3258, \8987_9286 );
and \U$11399 ( \20224_20526 , RIe1a2800_3226, \8989_9288 );
and \U$11400 ( \20225_20527 , RIe19fb00_3194, \8991_9290 );
and \U$11401 ( \20226_20528 , RIe18c000_2970, \8993_9292 );
and \U$11402 ( \20227_20529 , RIe178500_2746, \8995_9294 );
and \U$11403 ( \20228_20530 , RIe225e58_4721, \8997_9296 );
and \U$11404 ( \20229_20531 , RIe21aa58_4593, \8999_9298 );
and \U$11405 ( \20230_20532 , RIe204258_4337, \9001_9300 );
and \U$11406 ( \20231_20533 , RIe1fe2b8_4269, \9003_9302 );
and \U$11407 ( \20232_20534 , RIe1f7670_4192, \9005_9304 );
and \U$11408 ( \20233_20535 , RIe1f01b8_4109, \9007_9306 );
and \U$11409 ( \20234_20536 , RIe1d46c0_3794, \9009_9308 );
and \U$11410 ( \20235_20537 , RIe1bb1c0_3506, \9011_9310 );
and \U$11411 ( \20236_20538 , RIe1ae038_3357, \9013_9312 );
and \U$11412 ( \20237_20539 , RIe170670_2656, \9015_9314 );
or \U$11413 ( \20238_20540 , \20174_20476 , \20175_20477 , \20176_20478 , \20177_20479 , \20178_20480 , \20179_20481 , \20180_20482 , \20181_20483 , \20182_20484 , \20183_20485 , \20184_20486 , \20185_20487 , \20186_20488 , \20187_20489 , \20188_20490 , \20189_20491 , \20190_20492 , \20191_20493 , \20192_20494 , \20193_20495 , \20194_20496 , \20195_20497 , \20196_20498 , \20197_20499 , \20198_20500 , \20199_20501 , \20200_20502 , \20201_20503 , \20202_20504 , \20203_20505 , \20204_20506 , \20205_20507 , \20206_20508 , \20207_20509 , \20208_20510 , \20209_20511 , \20210_20512 , \20211_20513 , \20212_20514 , \20213_20515 , \20214_20516 , \20215_20517 , \20216_20518 , \20217_20519 , \20218_20520 , \20219_20521 , \20220_20522 , \20221_20523 , \20222_20524 , \20223_20525 , \20224_20526 , \20225_20527 , \20226_20528 , \20227_20529 , \20228_20530 , \20229_20531 , \20230_20532 , \20231_20533 , \20232_20534 , \20233_20535 , \20234_20536 , \20235_20537 , \20236_20538 , \20237_20539 );
or \U$11414 ( \20239_20541 , \20173_20475 , \20238_20540 );
_DC \g65a8/U$1 ( \20240 , \20239_20541 , \9024_9323 );
and g65a9_GF_PartitionCandidate( \20241_20543_nG65a9 , \20108 , \20240 );
buf \U$11415 ( \20242_20544 , \20241_20543_nG65a9 );
and \U$11416 ( \20243_20545 , \20242_20544 , \10389_10691 );
nor \U$11417 ( \20244_20546 , \19976_20278 , \20243_20545 );
xnor \U$11418 ( \20245_20547 , \20244_20546 , \10678_10980 );
and \U$11419 ( \20246_20548 , \17736_18035 , \11275_11574 );
and \U$11420 ( \20247_20549 , \18730_19032 , \10976_11278 );
nor \U$11421 ( \20248_20550 , \20246_20548 , \20247_20549 );
xnor \U$11422 ( \20249_20551 , \20248_20550 , \11281_11580 );
xor \U$11423 ( \20250_20552 , \20245_20547 , \20249_20551 );
_DC \g556a/U$1 ( \20251 , \20107_20409 , \9298_9597 );
_DC \g55ee/U$1 ( \20252 , \20239_20541 , \9024_9323 );
xor g55ef_GF_PartitionCandidate( \20253_20555_nG55ef , \20251 , \20252 );
buf \U$11424 ( \20254_20556 , \20253_20555_nG55ef );
xor \U$11425 ( \20255_20557 , \20254_20556 , \19232_19531 );
and \U$11426 ( \20256_20558 , \10385_10687 , \20255_20557 );
xor \U$11427 ( \20257_20559 , \20250_20552 , \20256_20558 );
xor \U$11428 ( \20258_20560 , \19975_20277 , \20257_20559 );
and \U$11429 ( \20259_20561 , \16353_16655 , \12491_12790 );
and \U$11430 ( \20260_20562 , \17325_17627 , \12159_12461 );
nor \U$11431 ( \20261_20563 , \20259_20561 , \20260_20562 );
xnor \U$11432 ( \20262_20564 , \20261_20563 , \12481_12780 );
and \U$11433 ( \20263_20565 , \12470_12769 , \16333_16635 );
and \U$11434 ( \20264_20566 , \13377_13679 , \15999_16301 );
nor \U$11435 ( \20265_20567 , \20263_20565 , \20264_20566 );
xnor \U$11436 ( \20266_20568 , \20265_20567 , \16323_16625 );
xor \U$11437 ( \20267_20569 , \20262_20564 , \20266_20568 );
and \U$11438 ( \20268_20570 , \11287_11586 , \17791_18090 );
and \U$11439 ( \20269_20571 , \12146_12448 , \17353_17655 );
nor \U$11440 ( \20270_20572 , \20268_20570 , \20269_20571 );
xnor \U$11441 ( \20271_20573 , \20270_20572 , \17747_18046 );
xor \U$11442 ( \20272_20574 , \20267_20569 , \20271_20573 );
xor \U$11443 ( \20273_20575 , \20258_20560 , \20272_20574 );
xor \U$11444 ( \20274_20576 , \19961_20263 , \20273_20575 );
and \U$11445 ( \20275_20577 , \19265_19564 , \19269_19568 );
and \U$11446 ( \20276_20578 , \19269_19568 , \19274_19573 );
and \U$11447 ( \20277_20579 , \19265_19564 , \19274_19573 );
or \U$11448 ( \20278_20580 , \20275_20577 , \20276_20578 , \20277_20579 );
and \U$11449 ( \20279_20581 , \18942_19241 , \18956_19255 );
and \U$11450 ( \20280_20582 , \18956_19255 , \19243_19542 );
and \U$11451 ( \20281_20583 , \18942_19241 , \19243_19542 );
or \U$11452 ( \20282_20584 , \20279_20581 , \20280_20582 , \20281_20583 );
xor \U$11453 ( \20283_20585 , \20278_20580 , \20282_20584 );
and \U$11454 ( \20284_20586 , \18946_19245 , \18950_19249 );
and \U$11455 ( \20285_20587 , \18950_19249 , \18955_19254 );
and \U$11456 ( \20286_20588 , \18946_19245 , \18955_19254 );
or \U$11457 ( \20287_20589 , \20284_20586 , \20285_20587 , \20286_20588 );
and \U$11458 ( \20288_20590 , \18961_19260 , \18965_19264 );
and \U$11459 ( \20289_20591 , \18965_19264 , \19242_19541 );
and \U$11460 ( \20290_20592 , \18961_19260 , \19242_19541 );
or \U$11461 ( \20291_20593 , \20288_20590 , \20289_20591 , \20290_20592 );
xor \U$11462 ( \20292_20594 , \20287_20589 , \20291_20593 );
and \U$11463 ( \20293_20595 , \19262_19561 , \19264_19563 );
xor \U$11464 ( \20294_20596 , \20292_20594 , \20293_20595 );
xor \U$11465 ( \20295_20597 , \20283_20585 , \20294_20596 );
xor \U$11466 ( \20296_20598 , \20274_20576 , \20295_20597 );
and \U$11467 ( \20297_20599 , \18938_19237 , \19244_19543 );
and \U$11468 ( \20298_20600 , \19244_19543 , \19276_19575 );
and \U$11469 ( \20299_20601 , \18938_19237 , \19276_19575 );
or \U$11470 ( \20300_20602 , \20297_20599 , \20298_20600 , \20299_20601 );
xor \U$11471 ( \20301_20603 , \20296_20598 , \20300_20602 );
and \U$11472 ( \20302_20604 , \19277_19576 , \19281_19580 );
and \U$11473 ( \20303_20605 , \19282_19581 , \19285_19584 );
or \U$11474 ( \20304_20606 , \20302_20604 , \20303_20605 );
xor \U$11475 ( \20305_20607 , \20301_20603 , \20304_20606 );
buf g9bde_GF_PartitionCandidate( \20306_20608_nG9bde , \20305_20607 );
and \U$11476 ( \20307_20609 , \10402_10704 , \20306_20608_nG9bde );
or \U$11477 ( \20308_20610 , \19957_20259 , \20307_20609 );
xor \U$11478 ( \20309_20611 , \10399_10703 , \20308_20610 );
buf \U$11479 ( \20310_20612 , \20309_20611 );
buf \U$11481 ( \20311_20613 , \20310_20612 );
xor \U$11482 ( \20312_20614 , \19956_20258 , \20311_20613 );
buf \U$11483 ( \20313_20615 , \20312_20614 );
xor \U$11484 ( \20314_20616 , \19929_20231 , \20313_20615 );
buf \U$11485 ( \20315_20617 , \20314_20616 );
xor \U$11486 ( \20316_20618 , \19871_20173 , \20315_20617 );
and \U$11487 ( \20317_20619 , \19304_19603 , \20316_20618 );
and \U$11488 ( \20318_20620 , \19859_20161 , \20316_20618 );
or \U$11489 ( \20319_20621 , \19860_20162 , \20317_20619 , \20318_20620 );
and \U$11490 ( \20320_20622 , \19865_20167 , \19870_20172 );
and \U$11491 ( \20321_20623 , \19865_20167 , \20315_20617 );
and \U$11492 ( \20322_20624 , \19870_20172 , \20315_20617 );
or \U$11493 ( \20323_20625 , \20320_20622 , \20321_20623 , \20322_20624 );
xor \U$11494 ( \20324_20626 , \20319_20621 , \20323_20625 );
and \U$11495 ( \20325_20627 , \19876_20178 , \19928_20230 );
and \U$11496 ( \20326_20628 , \19876_20178 , \20313_20615 );
and \U$11497 ( \20327_20629 , \19928_20230 , \20313_20615 );
or \U$11498 ( \20328_20630 , \20325_20627 , \20326_20628 , \20327_20629 );
xor \U$11499 ( \20329_20631 , \20324_20626 , \20328_20630 );
and \U$11500 ( \20330_20632 , \19949_20251 , \19955_20257 );
and \U$11501 ( \20331_20633 , \19949_20251 , \20311_20613 );
and \U$11502 ( \20332_20634 , \19955_20257 , \20311_20613 );
or \U$11503 ( \20333_20635 , \20330_20632 , \20331_20633 , \20332_20634 );
buf \U$11504 ( \20334_20636 , \20333_20635 );
and \U$11505 ( \20335_20637 , \19934_20236 , \19940_20242 );
and \U$11506 ( \20336_20638 , \19934_20236 , \19947_20249 );
and \U$11507 ( \20337_20639 , \19940_20242 , \19947_20249 );
or \U$11508 ( \20338_20640 , \20335_20637 , \20336_20638 , \20337_20639 );
buf \U$11509 ( \20339_20641 , \20338_20640 );
and \U$11510 ( \20340_20642 , \19852_20151 , \19856_20158 );
buf \U$11511 ( \20341_20643 , \20340_20642 );
buf \U$11513 ( \20342_20644 , \20341_20643 );
and \U$11514 ( \20343_20645 , \18908_18702 , \10981_11283_nG9c08 );
and \U$11515 ( \20344_20646 , \18400_18699 , \11299_11598_nG9c05 );
or \U$11516 ( \20345_20647 , \20343_20645 , \20344_20646 );
xor \U$11517 ( \20346_20648 , \18399_18698 , \20345_20647 );
buf \U$11518 ( \20347_20649 , \20346_20648 );
buf \U$11520 ( \20348_20650 , \20347_20649 );
xor \U$11521 ( \20349_20651 , \20342_20644 , \20348_20650 );
buf \U$11522 ( \20350_20652 , \20349_20651 );
not \U$11019 ( \20351_20153 , \19853_20152 );
xor \U$11020 ( \20352_20154 , \19847_20146_nG4424 , \19850_20149_nG4427 );
and \U$11021 ( \20353_20155 , \20351_20153 , \20352_20154 );
and \U$11523 ( \20354_20653 , \20353_20155 , \10392_10694_nG9c0e );
and \U$11524 ( \20355_20654 , \19853_20152 , \10693_10995_nG9c0b );
or \U$11525 ( \20356_20655 , \20354_20653 , \20355_20654 );
xor \U$11526 ( \20357_20656 , \19852_20151 , \20356_20655 );
buf \U$11527 ( \20358_20657 , \20357_20656 );
buf \U$11529 ( \20359_20658 , \20358_20657 );
xor \U$11530 ( \20360_20659 , \20350_20652 , \20359_20658 );
and \U$11531 ( \20361_20660 , \17437_17297 , \12168_12470_nG9c02 );
and \U$11532 ( \20362_20661 , \16995_17294 , \12502_12801_nG9bff );
or \U$11533 ( \20363_20662 , \20361_20660 , \20362_20661 );
xor \U$11534 ( \20364_20663 , \16994_17293 , \20363_20662 );
buf \U$11535 ( \20365_20664 , \20364_20663 );
buf \U$11537 ( \20366_20665 , \20365_20664 );
xor \U$11538 ( \20367_20666 , \20360_20659 , \20366_20665 );
buf \U$11539 ( \20368_20667 , \20367_20666 );
and \U$11540 ( \20369_20668 , \19894_20196 , \19900_20202 );
buf \U$11541 ( \20370_20669 , \20369_20668 );
xor \U$11542 ( \20371_20670 , \20368_20667 , \20370_20669 );
and \U$11543 ( \20372_20671 , \16405_15940 , \13403_13705_nG9bfc );
and \U$11544 ( \20373_20672 , \15638_15937 , \13771_14070_nG9bf9 );
or \U$11545 ( \20374_20673 , \20372_20671 , \20373_20672 );
xor \U$11546 ( \20375_20674 , \15637_15936 , \20374_20673 );
buf \U$11547 ( \20376_20675 , \20375_20674 );
buf \U$11549 ( \20377_20676 , \20376_20675 );
xor \U$11550 ( \20378_20677 , \20371_20670 , \20377_20676 );
buf \U$11551 ( \20379_20678 , \20378_20677 );
xor \U$11552 ( \20380_20679 , \20339_20641 , \20379_20678 );
and \U$11553 ( \20381_20680 , \12183_12157 , \17363_17665_nG9bea );
and \U$11554 ( \20382_20681 , \11855_12154 , \17808_18107_nG9be7 );
or \U$11555 ( \20383_20682 , \20381_20680 , \20382_20681 );
xor \U$11556 ( \20384_20683 , \11854_12153 , \20383_20682 );
buf \U$11557 ( \20385_20684 , \20384_20683 );
buf \U$11559 ( \20386_20685 , \20385_20684 );
xor \U$11560 ( \20387_20686 , \20380_20679 , \20386_20685 );
buf \U$11561 ( \20388_20687 , \20387_20686 );
xor \U$11562 ( \20389_20688 , \20334_20636 , \20388_20687 );
and \U$11563 ( \20390_20689 , \19886_20188 , \19911_20213 );
and \U$11564 ( \20391_20690 , \19886_20188 , \19918_20220 );
and \U$11565 ( \20392_20691 , \19911_20213 , \19918_20220 );
or \U$11566 ( \20393_20692 , \20390_20689 , \20391_20690 , \20392_20691 );
buf \U$11567 ( \20394_20693 , \20393_20692 );
xor \U$11568 ( \20395_20694 , \20389_20688 , \20394_20693 );
buf \U$11569 ( \20396_20695 , \20395_20694 );
and \U$11570 ( \20397_20696 , \19888_20190 , \19902_20204 );
and \U$11571 ( \20398_20697 , \19888_20190 , \19909_20211 );
and \U$11572 ( \20399_20698 , \19902_20204 , \19909_20211 );
or \U$11573 ( \20400_20699 , \20397_20696 , \20398_20697 , \20399_20698 );
buf \U$11574 ( \20401_20700 , \20400_20699 );
and \U$11575 ( \20402_20701 , \14710_14631 , \14682_14984_nG9bf6 );
and \U$11576 ( \20403_20702 , \14329_14628 , \15074_15373_nG9bf3 );
or \U$11577 ( \20404_20703 , \20402_20701 , \20403_20702 );
xor \U$11578 ( \20405_20704 , \14328_14627 , \20404_20703 );
buf \U$11579 ( \20406_20705 , \20405_20704 );
buf \U$11581 ( \20407_20706 , \20406_20705 );
xor \U$11582 ( \20408_20707 , \20401_20700 , \20407_20706 );
and \U$11583 ( \20409_20708 , \13431_13370 , \16013_16315_nG9bf0 );
and \U$11584 ( \20410_20709 , \13068_13367 , \16378_16680_nG9bed );
or \U$11585 ( \20411_20710 , \20409_20708 , \20410_20709 );
xor \U$11586 ( \20412_20711 , \13067_13366 , \20411_20710 );
buf \U$11587 ( \20413_20712 , \20412_20711 );
buf \U$11589 ( \20414_20713 , \20413_20712 );
xor \U$11590 ( \20415_20714 , \20408_20707 , \20414_20713 );
buf \U$11591 ( \20416_20715 , \20415_20714 );
and \U$11592 ( \20417_20716 , \10996_10421 , \18789_19091_nG9be4 );
and \U$11593 ( \20418_20717 , \10119_10418 , \19287_19586_nG9be1 );
or \U$11594 ( \20419_20718 , \20417_20716 , \20418_20717 );
xor \U$11595 ( \20420_20719 , \10118_10417 , \20419_20718 );
buf \U$11596 ( \20421_20720 , \20420_20719 );
buf \U$11598 ( \20422_20721 , \20421_20720 );
xor \U$11599 ( \20423_20722 , \20416_20715 , \20422_20721 );
and \U$11600 ( \20424_20723 , \10411_10707 , \20306_20608_nG9bde );
and \U$11601 ( \20425_20724 , \20278_20580 , \20282_20584 );
and \U$11602 ( \20426_20725 , \20282_20584 , \20294_20596 );
and \U$11603 ( \20427_20726 , \20278_20580 , \20294_20596 );
or \U$11604 ( \20428_20727 , \20425_20724 , \20426_20725 , \20427_20726 );
and \U$11605 ( \20429_20728 , \15965_16267 , \13755_14054 );
and \U$11606 ( \20430_20729 , \16353_16655 , \13390_13692 );
nor \U$11607 ( \20431_20730 , \20429_20728 , \20430_20729 );
xnor \U$11608 ( \20432_20731 , \20431_20730 , \13736_14035 );
and \U$11609 ( \20433_20732 , \10968_11270 , \19235_19534 );
and \U$11610 ( \20434_20733 , \11287_11586 , \18743_19045 );
nor \U$11611 ( \20435_20734 , \20433_20732 , \20434_20733 );
xnor \U$11612 ( \20436_20735 , \20435_20734 , \19241_19540 );
xor \U$11613 ( \20437_20736 , \20432_20731 , \20436_20735 );
and \U$11614 ( \20438_20737 , RIdec4cd0_703, \9034_9333 );
and \U$11615 ( \20439_20738 , RIdec1fd0_671, \9036_9335 );
and \U$11616 ( \20440_20739 , RIfc7b4b8_6425, \9038_9337 );
and \U$11617 ( \20441_20740 , RIdebf2d0_639, \9040_9339 );
and \U$11618 ( \20442_20741 , RIfc7b1e8_6423, \9042_9341 );
and \U$11619 ( \20443_20742 , RIdebc5d0_607, \9044_9343 );
and \U$11620 ( \20444_20743 , RIdeb98d0_575, \9046_9345 );
and \U$11621 ( \20445_20744 , RIdeb6bd0_543, \9048_9347 );
and \U$11622 ( \20446_20745 , RIfe83358_7837, \9050_9349 );
and \U$11623 ( \20447_20746 , RIdeb11d0_479, \9052_9351 );
and \U$11624 ( \20448_20747 , RIee1e5c8_4804, \9054_9353 );
and \U$11625 ( \20449_20748 , RIdeae4d0_447, \9056_9355 );
and \U$11626 ( \20450_20749 , RIfc437c0_5790, \9058_9357 );
and \U$11627 ( \20451_20750 , RIdea93b8_415, \9060_9359 );
and \U$11628 ( \20452_20751 , RIdea2ab8_383, \9062_9361 );
and \U$11629 ( \20453_20752 , RIde9c1b8_351, \9064_9363 );
and \U$11630 ( \20454_20753 , RIfc90ea8_6671, \9066_9365 );
and \U$11631 ( \20455_20754 , RIfc7af18_6421, \9068_9367 );
and \U$11632 ( \20456_20755 , RIfe83088_7835, \9070_9369 );
and \U$11633 ( \20457_20756 , RIee1a950_4761, \9072_9371 );
and \U$11634 ( \20458_20757 , RIde906b0_294, \9074_9373 );
and \U$11635 ( \20459_20758 , RIde8cba0_276, \9076_9375 );
and \U$11636 ( \20460_20759 , RIfe82f20_7834, \9078_9377 );
and \U$11637 ( \20461_20760 , RIfe82db8_7833, \9080_9379 );
and \U$11638 ( \20462_20761 , RIee1a248_4756, \9082_9381 );
and \U$11639 ( \20463_20762 , RIfe831f0_7836, \9084_9383 );
and \U$11640 ( \20464_20763 , RIfcc2390_7232, \9086_9385 );
and \U$11641 ( \20465_20764 , RIee195a0_4747, \9088_9387 );
and \U$11642 ( \20466_20765 , RIfcbe718_7189, \9090_9389 );
and \U$11643 ( \20467_20766 , RIfea9e18_8249, \9092_9391 );
and \U$11644 ( \20468_20767 , RIfc43220_5786, \9094_9393 );
and \U$11645 ( \20469_20768 , RIe167868_2555, \9096_9395 );
and \U$11646 ( \20470_20769 , RIe164cd0_2524, \9098_9397 );
and \U$11647 ( \20471_20770 , RIe161fd0_2492, \9100_9399 );
and \U$11648 ( \20472_20771 , RIee36f88_5084, \9102_9401 );
and \U$11649 ( \20473_20772 , RIe15f2d0_2460, \9104_9403 );
and \U$11650 ( \20474_20773 , RIee35ea8_5072, \9106_9405 );
and \U$11651 ( \20475_20774 , RIe15c5d0_2428, \9108_9407 );
and \U$11652 ( \20476_20775 , RIe156bd0_2364, \9110_9409 );
and \U$11653 ( \20477_20776 , RIe153ed0_2332, \9112_9411 );
and \U$11654 ( \20478_20777 , RIfe83628_7839, \9114_9413 );
and \U$11655 ( \20479_20778 , RIe1511d0_2300, \9116_9415 );
and \U$11656 ( \20480_20779 , RIfebfda8_8303, \9118_9417 );
and \U$11657 ( \20481_20780 , RIe14e4d0_2268, \9120_9419 );
and \U$11658 ( \20482_20781 , RIfebfc40_8302, \9122_9421 );
and \U$11659 ( \20483_20782 , RIe14b7d0_2236, \9124_9423 );
and \U$11660 ( \20484_20783 , RIe148ad0_2204, \9126_9425 );
and \U$11661 ( \20485_20784 , RIe145dd0_2172, \9128_9427 );
and \U$11662 ( \20486_20785 , RIee34120_5051, \9130_9429 );
and \U$11663 ( \20487_20786 , RIee32ed8_5038, \9132_9431 );
and \U$11664 ( \20488_20787 , RIee31df8_5026, \9134_9433 );
and \U$11665 ( \20489_20788 , RIfcc1f58_7229, \9136_9435 );
and \U$11666 ( \20490_20789 , RIe140ad8_2113, \9138_9437 );
and \U$11667 ( \20491_20790 , RIdf3e878_2088, \9140_9439 );
and \U$11668 ( \20492_20791 , RIfe834c0_7838, \9142_9441 );
and \U$11669 ( \20493_20792 , RIdf3a390_2039, \9144_9443 );
and \U$11670 ( \20494_20793 , RIfc5a6c8_6051, \9146_9445 );
and \U$11671 ( \20495_20794 , RIfc91e20_6682, \9148_9447 );
and \U$11672 ( \20496_20795 , RIee2e888_4988, \9150_9449 );
and \U$11673 ( \20497_20796 , RIfc96a10_6736, \9152_9451 );
and \U$11674 ( \20498_20797 , RIdf35098_1980, \9154_9453 );
and \U$11675 ( \20499_20798 , RIfeab600_8266, \9156_9455 );
and \U$11676 ( \20500_20799 , RIdf30bb0_1931, \9158_9457 );
and \U$11677 ( \20501_20800 , RIfeab768_8267, \9160_9459 );
or \U$11678 ( \20502_20801 , \20438_20737 , \20439_20738 , \20440_20739 , \20441_20740 , \20442_20741 , \20443_20742 , \20444_20743 , \20445_20744 , \20446_20745 , \20447_20746 , \20448_20747 , \20449_20748 , \20450_20749 , \20451_20750 , \20452_20751 , \20453_20752 , \20454_20753 , \20455_20754 , \20456_20755 , \20457_20756 , \20458_20757 , \20459_20758 , \20460_20759 , \20461_20760 , \20462_20761 , \20463_20762 , \20464_20763 , \20465_20764 , \20466_20765 , \20467_20766 , \20468_20767 , \20469_20768 , \20470_20769 , \20471_20770 , \20472_20771 , \20473_20772 , \20474_20773 , \20475_20774 , \20476_20775 , \20477_20776 , \20478_20777 , \20479_20778 , \20480_20779 , \20481_20780 , \20482_20781 , \20483_20782 , \20484_20783 , \20485_20784 , \20486_20785 , \20487_20786 , \20488_20787 , \20489_20788 , \20490_20789 , \20491_20790 , \20492_20791 , \20493_20792 , \20494_20793 , \20495_20794 , \20496_20795 , \20497_20796 , \20498_20797 , \20499_20798 , \20500_20799 , \20501_20800 );
and \U$11679 ( \20503_20802 , RIfcbe9e8_7191, \9163_9462 );
and \U$11680 ( \20504_20803 , RIfc79fa0_6410, \9165_9464 );
and \U$11681 ( \20505_20804 , RIfc96740_6734, \9167_9466 );
and \U$11682 ( \20506_20805 , RIfc92258_6685, \9169_9468 );
and \U$11683 ( \20507_20806 , RIfea7118_8217, \9171_9470 );
and \U$11684 ( \20508_20807 , RIfea95a8_8243, \9173_9472 );
and \U$11685 ( \20509_20808 , RIdf26020_1809, \9175_9474 );
and \U$11686 ( \20510_20809 , RIdf24400_1789, \9177_9476 );
and \U$11687 ( \20511_20810 , RIfc79a00_6406, \9179_9478 );
and \U$11688 ( \20512_20811 , RIfc5add0_6056, \9181_9480 );
and \U$11689 ( \20513_20812 , RIfce5d18_7637, \9183_9482 );
and \U$11690 ( \20514_20813 , RIfc92690_6688, \9185_9484 );
and \U$11691 ( \20515_20814 , RIfce3018_7605, \9187_9486 );
and \U$11692 ( \20516_20815 , RIdf1f270_1731, \9189_9488 );
and \U$11693 ( \20517_20816 , RIfc79730_6404, \9191_9490 );
and \U$11694 ( \20518_20817 , RIdf19000_1661, \9193_9492 );
and \U$11695 ( \20519_20818 , RIdf168a0_1633, \9195_9494 );
and \U$11696 ( \20520_20819 , RIdf13ba0_1601, \9197_9496 );
and \U$11697 ( \20521_20820 , RIdf10ea0_1569, \9199_9498 );
and \U$11698 ( \20522_20821 , RIdf0e1a0_1537, \9201_9500 );
and \U$11699 ( \20523_20822 , RIdf0b4a0_1505, \9203_9502 );
and \U$11700 ( \20524_20823 , RIdf087a0_1473, \9205_9504 );
and \U$11701 ( \20525_20824 , RIdf05aa0_1441, \9207_9506 );
and \U$11702 ( \20526_20825 , RIdf02da0_1409, \9209_9508 );
and \U$11703 ( \20527_20826 , RIdefd3a0_1345, \9211_9510 );
and \U$11704 ( \20528_20827 , RIdefa6a0_1313, \9213_9512 );
and \U$11705 ( \20529_20828 , RIdef79a0_1281, \9215_9514 );
and \U$11706 ( \20530_20829 , RIdef4ca0_1249, \9217_9516 );
and \U$11707 ( \20531_20830 , RIdef1fa0_1217, \9219_9518 );
and \U$11708 ( \20532_20831 , RIdeef2a0_1185, \9221_9520 );
and \U$11709 ( \20533_20832 , RIdeec5a0_1153, \9223_9522 );
and \U$11710 ( \20534_20833 , RIdee98a0_1121, \9225_9524 );
and \U$11711 ( \20535_20834 , RIfc5b7a8_6063, \9227_9526 );
and \U$11712 ( \20536_20835 , RIfc5b640_6062, \9229_9528 );
and \U$11713 ( \20537_20836 , RIfc931d0_6696, \9231_9530 );
and \U$11714 ( \20538_20837 , RIfcecac8_7715, \9233_9532 );
and \U$11715 ( \20539_20838 , RIdee4710_1063, \9235_9534 );
and \U$11716 ( \20540_20839 , RIdee26b8_1040, \9237_9536 );
and \U$11717 ( \20541_20840 , RIdee07c8_1018, \9239_9538 );
and \U$11718 ( \20542_20841 , RIdede4a0_993, \9241_9540 );
and \U$11719 ( \20543_20842 , RIfcbf0f0_7196, \9243_9542 );
and \U$11720 ( \20544_20843 , RIfcbf528_7199, \9245_9544 );
and \U$11721 ( \20545_20844 , RIfc792f8_6401, \9247_9546 );
and \U$11722 ( \20546_20845 , RIfc93068_6695, \9249_9548 );
and \U$11723 ( \20547_20846 , RIded91a8_934, \9251_9550 );
and \U$11724 ( \20548_20847 , RIded6d18_908, \9253_9552 );
and \U$11725 ( \20549_20848 , RIded4e28_886, \9255_9554 );
and \U$11726 ( \20550_20849 , RIded2998_860, \9257_9556 );
and \U$11727 ( \20551_20850 , RIded00d0_831, \9259_9558 );
and \U$11728 ( \20552_20851 , RIdecd3d0_799, \9261_9560 );
and \U$11729 ( \20553_20852 , RIdeca6d0_767, \9263_9562 );
and \U$11730 ( \20554_20853 , RIdec79d0_735, \9265_9564 );
and \U$11731 ( \20555_20854 , RIdeb3ed0_511, \9267_9566 );
and \U$11732 ( \20556_20855 , RIde958b8_319, \9269_9568 );
and \U$11733 ( \20557_20856 , RIe16dad8_2625, \9271_9570 );
and \U$11734 ( \20558_20857 , RIe1598d0_2396, \9273_9572 );
and \U$11735 ( \20559_20858 , RIe1430d0_2140, \9275_9574 );
and \U$11736 ( \20560_20859 , RIdf37ac8_2010, \9277_9576 );
and \U$11737 ( \20561_20860 , RIdf2c128_1878, \9279_9578 );
and \U$11738 ( \20562_20861 , RIdf1c9a8_1702, \9281_9580 );
and \U$11739 ( \20563_20862 , RIdf000a0_1377, \9283_9582 );
and \U$11740 ( \20564_20863 , RIdee6ba0_1089, \9285_9584 );
and \U$11741 ( \20565_20864 , RIdedb908_962, \9287_9586 );
and \U$11742 ( \20566_20865 , RIde7b800_192, \9289_9588 );
or \U$11743 ( \20567_20866 , \20503_20802 , \20504_20803 , \20505_20804 , \20506_20805 , \20507_20806 , \20508_20807 , \20509_20808 , \20510_20809 , \20511_20810 , \20512_20811 , \20513_20812 , \20514_20813 , \20515_20814 , \20516_20815 , \20517_20816 , \20518_20817 , \20519_20818 , \20520_20819 , \20521_20820 , \20522_20821 , \20523_20822 , \20524_20823 , \20525_20824 , \20526_20825 , \20527_20826 , \20528_20827 , \20529_20828 , \20530_20829 , \20531_20830 , \20532_20831 , \20533_20832 , \20534_20833 , \20535_20834 , \20536_20835 , \20537_20836 , \20538_20837 , \20539_20838 , \20540_20839 , \20541_20840 , \20542_20841 , \20543_20842 , \20544_20843 , \20545_20844 , \20546_20845 , \20547_20846 , \20548_20847 , \20549_20848 , \20550_20849 , \20551_20850 , \20552_20851 , \20553_20852 , \20554_20853 , \20555_20854 , \20556_20855 , \20557_20856 , \20558_20857 , \20559_20858 , \20560_20859 , \20561_20860 , \20562_20861 , \20563_20862 , \20564_20863 , \20565_20864 , \20566_20865 );
or \U$11744 ( \20568_20867 , \20502_20801 , \20567_20866 );
_DC \g5673/U$1 ( \20569 , \20568_20867 , \9298_9597 );
and \U$11745 ( \20570_20869 , RIe19cf68_3163, \8760_9059 );
and \U$11746 ( \20571_20870 , RIe19a268_3131, \8762_9061 );
and \U$11747 ( \20572_20871 , RIfc8d7d0_6632, \8764_9063 );
and \U$11748 ( \20573_20872 , RIe197568_3099, \8766_9065 );
and \U$11749 ( \20574_20873 , RIfc561e0_6002, \8768_9067 );
and \U$11750 ( \20575_20874 , RIe194868_3067, \8770_9069 );
and \U$11751 ( \20576_20875 , RIe191b68_3035, \8772_9071 );
and \U$11752 ( \20577_20876 , RIe18ee68_3003, \8774_9073 );
and \U$11753 ( \20578_20877 , RIe189468_2939, \8776_9075 );
and \U$11754 ( \20579_20878 , RIe186768_2907, \8778_9077 );
and \U$11755 ( \20580_20879 , RIf143330_5224, \8780_9079 );
and \U$11756 ( \20581_20880 , RIe183a68_2875, \8782_9081 );
and \U$11757 ( \20582_20881 , RIfc7d948_6451, \8784_9083 );
and \U$11758 ( \20583_20882 , RIe180d68_2843, \8786_9085 );
and \U$11759 ( \20584_20883 , RIe17e068_2811, \8788_9087 );
and \U$11760 ( \20585_20884 , RIe17b368_2779, \8790_9089 );
and \U$11761 ( \20586_20885 , RIfc564b0_6004, \8792_9091 );
and \U$11762 ( \20587_20886 , RIfcd6700_7462, \8794_9093 );
and \U$11763 ( \20588_20887 , RIfc461f0_5820, \8796_9095 );
and \U$11764 ( \20589_20888 , RIe175698_2713, \8798_9097 );
and \U$11765 ( \20590_20889 , RIfc46088_5819, \8800_9099 );
and \U$11766 ( \20591_20890 , RIfc45f20_5818, \8802_9101 );
and \U$11767 ( \20592_20891 , RIfc7dc18_6453, \8804_9103 );
and \U$11768 ( \20593_20892 , RIfcd69d0_7464, \8806_9105 );
and \U$11769 ( \20594_20893 , RIfc98630_6756, \8808_9107 );
and \U$11770 ( \20595_20894 , RIfcc2a98_7237, \8810_9109 );
and \U$11771 ( \20596_20895 , RIfc7d510_6448, \8812_9111 );
and \U$11772 ( \20597_20896 , RIe173208_2687, \8814_9113 );
and \U$11773 ( \20598_20897 , RIfc8e478_6641, \8816_9115 );
and \U$11774 ( \20599_20898 , RIfc45ae8_5815, \8818_9117 );
and \U$11775 ( \20600_20899 , RIfc8e8b0_6644, \8820_9119 );
and \U$11776 ( \20601_20900 , RIfc45980_5814, \8822_9121 );
and \U$11777 ( \20602_20901 , RIfe82ae8_7831, \8824_9123 );
and \U$11778 ( \20603_20902 , RIe2232c0_4690, \8826_9125 );
and \U$11779 ( \20604_20903 , RIf16ba10_5684, \8828_9127 );
and \U$11780 ( \20605_20904 , RIe2205c0_4658, \8830_9129 );
and \U$11781 ( \20606_20905 , RIfcd24e8_7415, \8832_9131 );
and \U$11782 ( \20607_20906 , RIe21d8c0_4626, \8834_9133 );
and \U$11783 ( \20608_20907 , RIe217ec0_4562, \8836_9135 );
and \U$11784 ( \20609_20908 , RIe2151c0_4530, \8838_9137 );
and \U$11785 ( \20610_20909 , RIfebf268_8295, \8840_9139 );
and \U$11786 ( \20611_20910 , RIe2124c0_4498, \8842_9141 );
and \U$11787 ( \20612_20911 , RIf168d10_5652, \8844_9143 );
and \U$11788 ( \20613_20912 , RIe20f7c0_4466, \8846_9145 );
and \U$11789 ( \20614_20913 , RIfc7d240_6446, \8848_9147 );
and \U$11790 ( \20615_20914 , RIe20cac0_4434, \8850_9149 );
and \U$11791 ( \20616_20915 , RIe209dc0_4402, \8852_9151 );
and \U$11792 ( \20617_20916 , RIe2070c0_4370, \8854_9153 );
and \U$11793 ( \20618_20917 , RIf166e20_5630, \8856_9155 );
and \U$11794 ( \20619_20918 , RIfebf6a0_8298, \8858_9157 );
and \U$11795 ( \20620_20919 , RIfebf808_8299, \8860_9159 );
and \U$11796 ( \20621_20920 , RIfebf538_8297, \8862_9161 );
and \U$11797 ( \20622_20921 , RIfc8eb80_6646, \8864_9163 );
and \U$11798 ( \20623_20922 , RIf164120_5598, \8866_9165 );
and \U$11799 ( \20624_20923 , RIfc453e0_5810, \8868_9167 );
and \U$11800 ( \20625_20924 , RIf161b28_5571, \8870_9169 );
and \U$11801 ( \20626_20925 , RIf15fc38_5549, \8872_9171 );
and \U$11802 ( \20627_20926 , RIf15dd48_5527, \8874_9173 );
and \U$11803 ( \20628_20927 , RIe1fc968_4251, \8876_9175 );
and \U$11804 ( \20629_20928 , RIe1fb888_4239, \8878_9177 );
and \U$11805 ( \20630_20929 , RIfebf3d0_8296, \8880_9179 );
and \U$11806 ( \20631_20930 , RIf15b318_5497, \8882_9181 );
and \U$11807 ( \20632_20931 , RIfca2518_6869, \8884_9183 );
and \U$11808 ( \20633_20932 , RIfc8f120_6650, \8886_9185 );
or \U$11809 ( \20634_20933 , \20570_20869 , \20571_20870 , \20572_20871 , \20573_20872 , \20574_20873 , \20575_20874 , \20576_20875 , \20577_20876 , \20578_20877 , \20579_20878 , \20580_20879 , \20581_20880 , \20582_20881 , \20583_20882 , \20584_20883 , \20585_20884 , \20586_20885 , \20587_20886 , \20588_20887 , \20589_20888 , \20590_20889 , \20591_20890 , \20592_20891 , \20593_20892 , \20594_20893 , \20595_20894 , \20596_20895 , \20597_20896 , \20598_20897 , \20599_20898 , \20600_20899 , \20601_20900 , \20602_20901 , \20603_20902 , \20604_20903 , \20605_20904 , \20606_20905 , \20607_20906 , \20608_20907 , \20609_20908 , \20610_20909 , \20611_20910 , \20612_20911 , \20613_20912 , \20614_20913 , \20615_20914 , \20616_20915 , \20617_20916 , \20618_20917 , \20619_20918 , \20620_20919 , \20621_20920 , \20622_20921 , \20623_20922 , \20624_20923 , \20625_20924 , \20626_20925 , \20627_20926 , \20628_20927 , \20629_20928 , \20630_20929 , \20631_20930 , \20632_20931 , \20633_20932 );
and \U$11810 ( \20635_20934 , RIfebfad8_8301, \8889_9188 );
and \U$11811 ( \20636_20935 , RIfebf970_8300, \8891_9190 );
and \U$11812 ( \20637_20936 , RIfc7cca0_6442, \8893_9192 );
and \U$11813 ( \20638_20937 , RIe1f9dd0_4220, \8895_9194 );
and \U$11814 ( \20639_20938 , RIfe82c50_7832, \8897_9196 );
and \U$11815 ( \20640_20939 , RIf155648_5431, \8899_9198 );
and \U$11816 ( \20641_20940 , RIfc8f288_6651, \8901_9200 );
and \U$11817 ( \20642_20941 , RIe1f4f10_4164, \8903_9202 );
and \U$11818 ( \20643_20942 , RIf152d80_5402, \8905_9204 );
and \U$11819 ( \20644_20943 , RIfc8f828_6655, \8907_9206 );
and \U$11820 ( \20645_20944 , RIfcb3b88_7067, \8909_9208 );
and \U$11821 ( \20646_20945 , RIe1f2d50_4140, \8911_9210 );
and \U$11822 ( \20647_20946 , RIfc445d0_5800, \8913_9212 );
and \U$11823 ( \20648_20947 , RIfc8faf8_6657, \8915_9214 );
and \U$11824 ( \20649_20948 , RIf14da88_5343, \8917_9216 );
and \U$11825 ( \20650_20949 , RIe1eda58_4081, \8919_9218 );
and \U$11826 ( \20651_20950 , RIe1eb028_4051, \8921_9220 );
and \U$11827 ( \20652_20951 , RIe1e8328_4019, \8923_9222 );
and \U$11828 ( \20653_20952 , RIe1e5628_3987, \8925_9224 );
and \U$11829 ( \20654_20953 , RIe1e2928_3955, \8927_9226 );
and \U$11830 ( \20655_20954 , RIe1dfc28_3923, \8929_9228 );
and \U$11831 ( \20656_20955 , RIe1dcf28_3891, \8931_9230 );
and \U$11832 ( \20657_20956 , RIe1da228_3859, \8933_9232 );
and \U$11833 ( \20658_20957 , RIe1d7528_3827, \8935_9234 );
and \U$11834 ( \20659_20958 , RIe1d1b28_3763, \8937_9236 );
and \U$11835 ( \20660_20959 , RIe1cee28_3731, \8939_9238 );
and \U$11836 ( \20661_20960 , RIe1cc128_3699, \8941_9240 );
and \U$11837 ( \20662_20961 , RIe1c9428_3667, \8943_9242 );
and \U$11838 ( \20663_20962 , RIe1c6728_3635, \8945_9244 );
and \U$11839 ( \20664_20963 , RIe1c3a28_3603, \8947_9246 );
and \U$11840 ( \20665_20964 , RIe1c0d28_3571, \8949_9248 );
and \U$11841 ( \20666_20965 , RIe1be028_3539, \8951_9250 );
and \U$11842 ( \20667_20966 , RIfc7bff8_6433, \8953_9252 );
and \U$11843 ( \20668_20967 , RIfc44030_5796, \8955_9254 );
and \U$11844 ( \20669_20968 , RIe1b9000_3482, \8957_9256 );
and \U$11845 ( \20670_20969 , RIe1b6fa8_3459, \8959_9258 );
and \U$11846 ( \20671_20970 , RIfcbdd40_7182, \8961_9260 );
and \U$11847 ( \20672_20971 , RIfc8ff30_6660, \8963_9262 );
and \U$11848 ( \20673_20972 , RIe1b50b8_3437, \8965_9264 );
and \U$11849 ( \20674_20973 , RIe1b3d08_3423, \8967_9266 );
and \U$11850 ( \20675_20974 , RIfcbe178_7185, \8969_9268 );
and \U$11851 ( \20676_20975 , RIfc43d60_5794, \8971_9270 );
and \U$11852 ( \20677_20976 , RIe1b2520_3406, \8973_9272 );
and \U$11853 ( \20678_20977 , RIe1b0798_3385, \8975_9274 );
and \U$11854 ( \20679_20978 , RIfcdb5c0_7518, \8977_9276 );
and \U$11855 ( \20680_20979 , RIfc7ba58_6429, \8979_9278 );
and \U$11856 ( \20681_20980 , RIe1ac148_3335, \8981_9280 );
and \U$11857 ( \20682_20981 , RIe1aa960_3318, \8983_9282 );
and \U$11858 ( \20683_20982 , RIe1a8368_3291, \8985_9284 );
and \U$11859 ( \20684_20983 , RIe1a5668_3259, \8987_9286 );
and \U$11860 ( \20685_20984 , RIe1a2968_3227, \8989_9288 );
and \U$11861 ( \20686_20985 , RIe19fc68_3195, \8991_9290 );
and \U$11862 ( \20687_20986 , RIe18c168_2971, \8993_9292 );
and \U$11863 ( \20688_20987 , RIe178668_2747, \8995_9294 );
and \U$11864 ( \20689_20988 , RIe225fc0_4722, \8997_9296 );
and \U$11865 ( \20690_20989 , RIe21abc0_4594, \8999_9298 );
and \U$11866 ( \20691_20990 , RIe2043c0_4338, \9001_9300 );
and \U$11867 ( \20692_20991 , RIe1fe420_4270, \9003_9302 );
and \U$11868 ( \20693_20992 , RIe1f77d8_4193, \9005_9304 );
and \U$11869 ( \20694_20993 , RIe1f0320_4110, \9007_9306 );
and \U$11870 ( \20695_20994 , RIe1d4828_3795, \9009_9308 );
and \U$11871 ( \20696_20995 , RIe1bb328_3507, \9011_9310 );
and \U$11872 ( \20697_20996 , RIe1ae1a0_3358, \9013_9312 );
and \U$11873 ( \20698_20997 , RIe1707d8_2657, \9015_9314 );
or \U$11874 ( \20699_20998 , \20635_20934 , \20636_20935 , \20637_20936 , \20638_20937 , \20639_20938 , \20640_20939 , \20641_20940 , \20642_20941 , \20643_20942 , \20644_20943 , \20645_20944 , \20646_20945 , \20647_20946 , \20648_20947 , \20649_20948 , \20650_20949 , \20651_20950 , \20652_20951 , \20653_20952 , \20654_20953 , \20655_20954 , \20656_20955 , \20657_20956 , \20658_20957 , \20659_20958 , \20660_20959 , \20661_20960 , \20662_20961 , \20663_20962 , \20664_20963 , \20665_20964 , \20666_20965 , \20667_20966 , \20668_20967 , \20669_20968 , \20670_20969 , \20671_20970 , \20672_20971 , \20673_20972 , \20674_20973 , \20675_20974 , \20676_20975 , \20677_20976 , \20678_20977 , \20679_20978 , \20680_20979 , \20681_20980 , \20682_20981 , \20683_20982 , \20684_20983 , \20685_20984 , \20686_20985 , \20687_20986 , \20688_20987 , \20689_20988 , \20690_20989 , \20691_20990 , \20692_20991 , \20693_20992 , \20694_20993 , \20695_20994 , \20696_20995 , \20697_20996 , \20698_20997 );
or \U$11875 ( \20700_20999 , \20634_20933 , \20699_20998 );
_DC \g56f7/U$1 ( \20701 , \20700_20999 , \9024_9323 );
xor g56f8_GF_PartitionCandidate( \20702_21001_nG56f8 , \20569 , \20701 );
buf \U$11876 ( \20703_21002 , \20702_21001_nG56f8 );
xor \U$11877 ( \20704_21003 , \20703_21002 , \20254_20556 );
not \U$11878 ( \20705_21004 , \20255_20557 );
and \U$11879 ( \20706_21005 , \20704_21003 , \20705_21004 );
and \U$11880 ( \20707_21006 , \10385_10687 , \20706_21005 );
and \U$11881 ( \20708_21007 , \10686_10988 , \20255_20557 );
nor \U$11882 ( \20709_21008 , \20707_21006 , \20708_21007 );
and \U$11883 ( \20710_21009 , \20254_20556 , \19232_19531 );
not \U$11884 ( \20711_21010 , \20710_21009 );
and \U$11885 ( \20712_21011 , \20703_21002 , \20711_21010 );
xnor \U$11886 ( \20713_21012 , \20709_21008 , \20712_21011 );
xor \U$11887 ( \20714_21013 , \20437_20736 , \20713_21012 );
and \U$11888 ( \20715_21014 , \18730_19032 , \11275_11574 );
and \U$11889 ( \20716_21015 , \19259_19558 , \10976_11278 );
nor \U$11890 ( \20717_21016 , \20715_21014 , \20716_21015 );
xnor \U$11891 ( \20718_21017 , \20717_21016 , \11281_11580 );
and \U$11892 ( \20719_21018 , \17325_17627 , \12491_12790 );
and \U$11893 ( \20720_21019 , \17736_18035 , \12159_12461 );
nor \U$11894 ( \20721_21020 , \20719_21018 , \20720_21019 );
xnor \U$11895 ( \20722_21021 , \20721_21020 , \12481_12780 );
xor \U$11896 ( \20723_21022 , \20718_21017 , \20722_21021 );
and \U$11897 ( \20724_21023 , \14648_14950 , \15037_15336 );
and \U$11898 ( \20725_21024 , \15022_15321 , \14661_14963 );
nor \U$11899 ( \20726_21025 , \20724_21023 , \20725_21024 );
xnor \U$11900 ( \20727_21026 , \20726_21025 , \15043_15342 );
xor \U$11901 ( \20728_21027 , \20723_21022 , \20727_21026 );
xor \U$11902 ( \20729_21028 , \20714_21013 , \20728_21027 );
and \U$11903 ( \20730_21029 , \20242_20544 , \10681_10983 );
_DC \g65aa/U$1 ( \20731 , \20568_20867 , \9298_9597 );
_DC \g65ab/U$1 ( \20732 , \20700_20999 , \9024_9323 );
and g65ac_GF_PartitionCandidate( \20733_21032_nG65ac , \20731 , \20732 );
buf \U$11904 ( \20734_21033 , \20733_21032_nG65ac );
and \U$11905 ( \20735_21034 , \20734_21033 , \10389_10691 );
nor \U$11906 ( \20736_21035 , \20730_21029 , \20735_21034 );
xnor \U$11907 ( \20737_21036 , \20736_21035 , \10678_10980 );
not \U$11908 ( \20738_21037 , \20256_20558 );
and \U$11909 ( \20739_21038 , \20738_21037 , \20712_21011 );
xor \U$11910 ( \20740_21039 , \20737_21036 , \20739_21038 );
and \U$11911 ( \20741_21040 , \13377_13679 , \16333_16635 );
and \U$11912 ( \20742_21041 , \13725_14024 , \15999_16301 );
nor \U$11913 ( \20743_21042 , \20741_21040 , \20742_21041 );
xnor \U$11914 ( \20744_21043 , \20743_21042 , \16323_16625 );
xor \U$11915 ( \20745_21044 , \20740_21039 , \20744_21043 );
and \U$11916 ( \20746_21045 , \12146_12448 , \17791_18090 );
and \U$11917 ( \20747_21046 , \12470_12769 , \17353_17655 );
nor \U$11918 ( \20748_21047 , \20746_21045 , \20747_21046 );
xnor \U$11919 ( \20749_21048 , \20748_21047 , \17747_18046 );
xor \U$11920 ( \20750_21049 , \20745_21044 , \20749_21048 );
xor \U$11921 ( \20751_21050 , \20729_21028 , \20750_21049 );
xor \U$11922 ( \20752_21051 , \20428_20727 , \20751_21050 );
and \U$11923 ( \20753_21052 , \20287_20589 , \20291_20593 );
and \U$11924 ( \20754_21053 , \20291_20593 , \20293_20595 );
and \U$11925 ( \20755_21054 , \20287_20589 , \20293_20595 );
or \U$11926 ( \20756_21055 , \20753_21052 , \20754_21053 , \20755_21054 );
and \U$11927 ( \20757_21056 , \19975_20277 , \20257_20559 );
and \U$11928 ( \20758_21057 , \20257_20559 , \20272_20574 );
and \U$11929 ( \20759_21058 , \19975_20277 , \20272_20574 );
or \U$11930 ( \20760_21059 , \20757_21056 , \20758_21057 , \20759_21058 );
xor \U$11931 ( \20761_21060 , \20756_21055 , \20760_21059 );
and \U$11932 ( \20762_21061 , \19965_20267 , \19969_20271 );
and \U$11933 ( \20763_21062 , \19969_20271 , \19974_20276 );
and \U$11934 ( \20764_21063 , \19965_20267 , \19974_20276 );
or \U$11935 ( \20765_21064 , \20762_21061 , \20763_21062 , \20764_21063 );
and \U$11936 ( \20766_21065 , \20245_20547 , \20249_20551 );
and \U$11937 ( \20767_21066 , \20249_20551 , \20256_20558 );
and \U$11938 ( \20768_21067 , \20245_20547 , \20256_20558 );
or \U$11939 ( \20769_21068 , \20766_21065 , \20767_21066 , \20768_21067 );
xor \U$11940 ( \20770_21069 , \20765_21064 , \20769_21068 );
and \U$11941 ( \20771_21070 , \20262_20564 , \20266_20568 );
and \U$11942 ( \20772_21071 , \20266_20568 , \20271_20573 );
and \U$11943 ( \20773_21072 , \20262_20564 , \20271_20573 );
or \U$11944 ( \20774_21073 , \20771_21070 , \20772_21071 , \20773_21072 );
xor \U$11945 ( \20775_21074 , \20770_21069 , \20774_21073 );
xor \U$11946 ( \20776_21075 , \20761_21060 , \20775_21074 );
xor \U$11947 ( \20777_21076 , \20752_21051 , \20776_21075 );
and \U$11948 ( \20778_21077 , \19961_20263 , \20273_20575 );
and \U$11949 ( \20779_21078 , \20273_20575 , \20295_20597 );
and \U$11950 ( \20780_21079 , \19961_20263 , \20295_20597 );
or \U$11951 ( \20781_21080 , \20778_21077 , \20779_21078 , \20780_21079 );
xor \U$11952 ( \20782_21081 , \20777_21076 , \20781_21080 );
and \U$11953 ( \20783_21082 , \20296_20598 , \20300_20602 );
and \U$11954 ( \20784_21083 , \20301_20603 , \20304_20606 );
or \U$11955 ( \20785_21084 , \20783_21082 , \20784_21083 );
xor \U$11956 ( \20786_21085 , \20782_21081 , \20785_21084 );
buf g9bdb_GF_PartitionCandidate( \20787_21086_nG9bdb , \20786_21085 );
and \U$11957 ( \20788_21087 , \10402_10704 , \20787_21086_nG9bdb );
or \U$11958 ( \20789_21088 , \20424_20723 , \20788_21087 );
xor \U$11959 ( \20790_21089 , \10399_10703 , \20789_21088 );
buf \U$11960 ( \20791_21090 , \20790_21089 );
buf \U$11962 ( \20792_21091 , \20791_21090 );
xor \U$11963 ( \20793_21092 , \20423_20722 , \20792_21091 );
buf \U$11964 ( \20794_21093 , \20793_21092 );
xor \U$11965 ( \20795_21094 , \20396_20695 , \20794_21093 );
and \U$11966 ( \20796_21095 , \19881_20183 , \19920_20222 );
and \U$11967 ( \20797_21096 , \19881_20183 , \19926_20228 );
and \U$11968 ( \20798_21097 , \19920_20222 , \19926_20228 );
or \U$11969 ( \20799_21098 , \20796_21095 , \20797_21096 , \20798_21097 );
buf \U$11970 ( \20800_21099 , \20799_21098 );
xor \U$11971 ( \20801_21100 , \20795_21094 , \20800_21099 );
and \U$11972 ( \20802_21101 , \20329_20631 , \20801_21100 );
and \U$11973 ( \20803_21102 , \20319_20621 , \20323_20625 );
and \U$11974 ( \20804_21103 , \20319_20621 , \20328_20630 );
and \U$11975 ( \20805_21104 , \20323_20625 , \20328_20630 );
or \U$11976 ( \20806_21105 , \20803_21102 , \20804_21103 , \20805_21104 );
xor \U$11977 ( \20807_21106 , \20802_21101 , \20806_21105 );
and \U$11978 ( \20808_21107 , RIdec4fa0_705, \8760_9059 );
and \U$11979 ( \20809_21108 , RIdec22a0_673, \8762_9061 );
and \U$11980 ( \20810_21109 , RIee1fdb0_4821, \8764_9063 );
and \U$11981 ( \20811_21110 , RIdebf5a0_641, \8766_9065 );
and \U$11982 ( \20812_21111 , RIee1f270_4813, \8768_9067 );
and \U$11983 ( \20813_21112 , RIdebc8a0_609, \8770_9069 );
and \U$11984 ( \20814_21113 , RIdeb9ba0_577, \8772_9071 );
and \U$11985 ( \20815_21114 , RIdeb6ea0_545, \8774_9073 );
and \U$11986 ( \20816_21115 , RIee1ecd0_4809, \8776_9075 );
and \U$11987 ( \20817_21116 , RIdeb14a0_481, \8778_9077 );
and \U$11988 ( \20818_21117 , RIee1e730_4805, \8780_9079 );
and \U$11989 ( \20819_21118 , RIdeae7a0_449, \8782_9081 );
and \U$11990 ( \20820_21119 , RIee1d920_4795, \8784_9083 );
and \U$11991 ( \20821_21120 , RIdea9a48_417, \8786_9085 );
and \U$11992 ( \20822_21121 , RIdea3148_385, \8788_9087 );
and \U$11993 ( \20823_21122 , RIde9c848_353, \8790_9089 );
and \U$11994 ( \20824_21123 , RIee1cb10_4785, \8792_9091 );
and \U$11995 ( \20825_21124 , RIee1ba30_4773, \8794_9093 );
and \U$11996 ( \20826_21125 , RIee1b1c0_4767, \8796_9095 );
and \U$11997 ( \20827_21126 , RIfec04b0_8308, \8798_9097 );
and \U$11998 ( \20828_21127 , RIfe850e0_7858, \8800_9099 );
and \U$11999 ( \20829_21128 , RIde8d230_278, \8802_9101 );
and \U$12000 ( \20830_21129 , RIfea9cb0_8248, \8804_9103 );
and \U$12001 ( \20831_21130 , RIfe84f78_7857, \8806_9105 );
and \U$12002 ( \20832_21131 , RIee1a3b0_4757, \8808_9107 );
and \U$12003 ( \20833_21132 , RIfe853b0_7860, \8810_9109 );
and \U$12004 ( \20834_21133 , RIee199d8_4750, \8812_9111 );
and \U$12005 ( \20835_21134 , RIfe85248_7859, \8814_9113 );
and \U$12006 ( \20836_21135 , RIee39148_5108, \8816_9115 );
and \U$12007 ( \20837_21136 , RIe16b378_2597, \8818_9117 );
and \U$12008 ( \20838_21137 , RIee38608_5100, \8820_9119 );
and \U$12009 ( \20839_21138 , RIe167b38_2557, \8822_9121 );
and \U$12010 ( \20840_21139 , RIe164fa0_2526, \8824_9123 );
and \U$12011 ( \20841_21140 , RIe1622a0_2494, \8826_9125 );
and \U$12012 ( \20842_21141 , RIfe85950_7864, \8828_9127 );
and \U$12013 ( \20843_21142 , RIe15f5a0_2462, \8830_9129 );
and \U$12014 ( \20844_21143 , RIee36010_5073, \8832_9131 );
and \U$12015 ( \20845_21144 , RIe15c8a0_2430, \8834_9133 );
and \U$12016 ( \20846_21145 , RIe156ea0_2366, \8836_9135 );
and \U$12017 ( \20847_21146 , RIe1541a0_2334, \8838_9137 );
and \U$12018 ( \20848_21147 , RIfe85c20_7866, \8840_9139 );
and \U$12019 ( \20849_21148 , RIe1514a0_2302, \8842_9141 );
and \U$12020 ( \20850_21149 , RIee34dc8_5060, \8844_9143 );
and \U$12021 ( \20851_21150 , RIe14e7a0_2270, \8846_9145 );
and \U$12022 ( \20852_21151 , RIfc861b0_6548, \8848_9147 );
and \U$12023 ( \20853_21152 , RIe14baa0_2238, \8850_9149 );
and \U$12024 ( \20854_21153 , RIe148da0_2206, \8852_9151 );
and \U$12025 ( \20855_21154 , RIe1460a0_2174, \8854_9153 );
and \U$12026 ( \20856_21155 , RIee343f0_5053, \8856_9155 );
and \U$12027 ( \20857_21156 , RIfe85518_7861, \8858_9157 );
and \U$12028 ( \20858_21157 , RIfe857e8_7863, \8860_9159 );
and \U$12029 ( \20859_21158 , RIfe85680_7862, \8862_9161 );
and \U$12030 ( \20860_21159 , RIe140c40_2114, \8864_9163 );
and \U$12031 ( \20861_21160 , RIdf3eb48_2090, \8866_9165 );
and \U$12032 ( \20862_21161 , RIdf3c820_2065, \8868_9167 );
and \U$12033 ( \20863_21162 , RIdf3a660_2041, \8870_9169 );
and \U$12034 ( \20864_21163 , RIfc9d4f0_6812, \8872_9171 );
and \U$12035 ( \20865_21164 , RIee2f698_4998, \8874_9173 );
and \U$12036 ( \20866_21165 , RIfc52298_5957, \8876_9175 );
and \U$12037 ( \20867_21166 , RIee2d4d8_4974, \8878_9177 );
and \U$12038 ( \20868_21167 , RIdf35368_1982, \8880_9179 );
and \U$12039 ( \20869_21168 , RIdf32ed8_1956, \8882_9181 );
and \U$12040 ( \20870_21169 , RIdf30e80_1933, \8884_9183 );
and \U$12041 ( \20871_21170 , RIfe85ab8_7865, \8886_9185 );
or \U$12042 ( \20872_21171 , \20808_21107 , \20809_21108 , \20810_21109 , \20811_21110 , \20812_21111 , \20813_21112 , \20814_21113 , \20815_21114 , \20816_21115 , \20817_21116 , \20818_21117 , \20819_21118 , \20820_21119 , \20821_21120 , \20822_21121 , \20823_21122 , \20824_21123 , \20825_21124 , \20826_21125 , \20827_21126 , \20828_21127 , \20829_21128 , \20830_21129 , \20831_21130 , \20832_21131 , \20833_21132 , \20834_21133 , \20835_21134 , \20836_21135 , \20837_21136 , \20838_21137 , \20839_21138 , \20840_21139 , \20841_21140 , \20842_21141 , \20843_21142 , \20844_21143 , \20845_21144 , \20846_21145 , \20847_21146 , \20848_21147 , \20849_21148 , \20850_21149 , \20851_21150 , \20852_21151 , \20853_21152 , \20854_21153 , \20855_21154 , \20856_21155 , \20857_21156 , \20858_21157 , \20859_21158 , \20860_21159 , \20861_21160 , \20862_21161 , \20863_21162 , \20864_21163 , \20865_21164 , \20866_21165 , \20867_21166 , \20868_21167 , \20869_21168 , \20870_21169 , \20871_21170 );
and \U$12043 ( \20873_21172 , RIee2b8b8_4954, \8889_9188 );
and \U$12044 ( \20874_21173 , RIee29f68_4936, \8891_9190 );
and \U$12045 ( \20875_21174 , RIee28bb8_4922, \8893_9192 );
and \U$12046 ( \20876_21175 , RIee27970_4909, \8895_9194 );
and \U$12047 ( \20877_21176 , RIdf2a0d0_1855, \8897_9196 );
and \U$12048 ( \20878_21177 , RIfe84e10_7856, \8899_9198 );
and \U$12049 ( \20879_21178 , RIdf262f0_1811, \8901_9200 );
and \U$12050 ( \20880_21179 , RIfe84ca8_7855, \8903_9202 );
and \U$12051 ( \20881_21180 , RIee27100_4903, \8905_9204 );
and \U$12052 ( \20882_21181 , RIee26b60_4899, \8907_9206 );
and \U$12053 ( \20883_21182 , RIfcd32f8_7425, \8909_9208 );
and \U$12054 ( \20884_21183 , RIee265c0_4895, \8911_9210 );
and \U$12055 ( \20885_21184 , RIfc9e300_6822, \8913_9212 );
and \U$12056 ( \20886_21185 , RIdf1f540_1733, \8915_9214 );
and \U$12057 ( \20887_21186 , RIee25eb8_4890, \8917_9216 );
and \U$12058 ( \20888_21187 , RIfe84b40_7854, \8919_9218 );
and \U$12059 ( \20889_21188 , RIdf16b70_1635, \8921_9220 );
and \U$12060 ( \20890_21189 , RIdf13e70_1603, \8923_9222 );
and \U$12061 ( \20891_21190 , RIdf11170_1571, \8925_9224 );
and \U$12062 ( \20892_21191 , RIdf0e470_1539, \8927_9226 );
and \U$12063 ( \20893_21192 , RIdf0b770_1507, \8929_9228 );
and \U$12064 ( \20894_21193 , RIdf08a70_1475, \8931_9230 );
and \U$12065 ( \20895_21194 , RIdf05d70_1443, \8933_9232 );
and \U$12066 ( \20896_21195 , RIdf03070_1411, \8935_9234 );
and \U$12067 ( \20897_21196 , RIdefd670_1347, \8937_9236 );
and \U$12068 ( \20898_21197 , RIdefa970_1315, \8939_9238 );
and \U$12069 ( \20899_21198 , RIdef7c70_1283, \8941_9240 );
and \U$12070 ( \20900_21199 , RIdef4f70_1251, \8943_9242 );
and \U$12071 ( \20901_21200 , RIdef2270_1219, \8945_9244 );
and \U$12072 ( \20902_21201 , RIdeef570_1187, \8947_9246 );
and \U$12073 ( \20903_21202 , RIdeec870_1155, \8949_9248 );
and \U$12074 ( \20904_21203 , RIdee9b70_1123, \8951_9250 );
and \U$12075 ( \20905_21204 , RIfec0348_8307, \8953_9252 );
and \U$12076 ( \20906_21205 , RIfcb54d8_7085, \8955_9254 );
and \U$12077 ( \20907_21206 , RIee23cf8_4866, \8957_9256 );
and \U$12078 ( \20908_21207 , RIfc54e30_5988, \8959_9258 );
and \U$12079 ( \20909_21208 , RIfec0078_8305, \8961_9260 );
and \U$12080 ( \20910_21209 , RIdee2988_1042, \8963_9262 );
and \U$12081 ( \20911_21210 , RIfec01e0_8306, \8965_9264 );
and \U$12082 ( \20912_21211 , RIdede770_995, \8967_9266 );
and \U$12083 ( \20913_21212 , RIfcd7ee8_7479, \8969_9268 );
and \U$12084 ( \20914_21213 , RIfcd43d8_7437, \8971_9270 );
and \U$12085 ( \20915_21214 , RIfc88eb0_6580, \8973_9272 );
and \U$12086 ( \20916_21215 , RIfc9e5d0_6824, \8975_9274 );
and \U$12087 ( \20917_21216 , RIded9478_936, \8977_9276 );
and \U$12088 ( \20918_21217 , RIded6fe8_910, \8979_9278 );
and \U$12089 ( \20919_21218 , RIded50f8_888, \8981_9280 );
and \U$12090 ( \20920_21219 , RIfeab330_8264, \8983_9282 );
and \U$12091 ( \20921_21220 , RIded03a0_833, \8985_9284 );
and \U$12092 ( \20922_21221 , RIdecd6a0_801, \8987_9286 );
and \U$12093 ( \20923_21222 , RIdeca9a0_769, \8989_9288 );
and \U$12094 ( \20924_21223 , RIdec7ca0_737, \8991_9290 );
and \U$12095 ( \20925_21224 , RIdeb41a0_513, \8993_9292 );
and \U$12096 ( \20926_21225 , RIde95f48_321, \8995_9294 );
and \U$12097 ( \20927_21226 , RIe16dda8_2627, \8997_9296 );
and \U$12098 ( \20928_21227 , RIe159ba0_2398, \8999_9298 );
and \U$12099 ( \20929_21228 , RIe1433a0_2142, \9001_9300 );
and \U$12100 ( \20930_21229 , RIdf37d98_2012, \9003_9302 );
and \U$12101 ( \20931_21230 , RIdf2c3f8_1880, \9005_9304 );
and \U$12102 ( \20932_21231 , RIdf1cc78_1704, \9007_9306 );
and \U$12103 ( \20933_21232 , RIdf00370_1379, \9009_9308 );
and \U$12104 ( \20934_21233 , RIdee6e70_1091, \9011_9310 );
and \U$12105 ( \20935_21234 , RIdedbbd8_964, \9013_9312 );
and \U$12106 ( \20936_21235 , RIde7be90_194, \9015_9314 );
or \U$12107 ( \20937_21236 , \20873_21172 , \20874_21173 , \20875_21174 , \20876_21175 , \20877_21176 , \20878_21177 , \20879_21178 , \20880_21179 , \20881_21180 , \20882_21181 , \20883_21182 , \20884_21183 , \20885_21184 , \20886_21185 , \20887_21186 , \20888_21187 , \20889_21188 , \20890_21189 , \20891_21190 , \20892_21191 , \20893_21192 , \20894_21193 , \20895_21194 , \20896_21195 , \20897_21196 , \20898_21197 , \20899_21198 , \20900_21199 , \20901_21200 , \20902_21201 , \20903_21202 , \20904_21203 , \20905_21204 , \20906_21205 , \20907_21206 , \20908_21207 , \20909_21208 , \20910_21209 , \20911_21210 , \20912_21211 , \20913_21212 , \20914_21213 , \20915_21214 , \20916_21215 , \20917_21216 , \20918_21217 , \20919_21218 , \20920_21219 , \20921_21220 , \20922_21221 , \20923_21222 , \20924_21223 , \20925_21224 , \20926_21225 , \20927_21226 , \20928_21227 , \20929_21228 , \20930_21229 , \20931_21230 , \20932_21231 , \20933_21232 , \20934_21233 , \20935_21234 , \20936_21235 );
or \U$12108 ( \20938_21237 , \20872_21171 , \20937_21236 );
_DC \g2871/U$1 ( \20939 , \20938_21237 , \9024_9323 );
buf \U$12109 ( \20940_21239 , \20939 );
and \U$12110 ( \20941_21240 , RIe19d238_3165, \9034_9333 );
and \U$12111 ( \20942_21241 , RIe19a538_3133, \9036_9335 );
and \U$12112 ( \20943_21242 , RIf145658_5249, \9038_9337 );
and \U$12113 ( \20944_21243 , RIe197838_3101, \9040_9339 );
and \U$12114 ( \20945_21244 , RIf1446e0_5238, \9042_9341 );
and \U$12115 ( \20946_21245 , RIe194b38_3069, \9044_9343 );
and \U$12116 ( \20947_21246 , RIe191e38_3037, \9046_9345 );
and \U$12117 ( \20948_21247 , RIe18f138_3005, \9048_9347 );
and \U$12118 ( \20949_21248 , RIe189738_2941, \9050_9349 );
and \U$12119 ( \20950_21249 , RIe186a38_2909, \9052_9351 );
and \U$12120 ( \20951_21250 , RIf143600_5226, \9054_9353 );
and \U$12121 ( \20952_21251 , RIe183d38_2877, \9056_9355 );
and \U$12122 ( \20953_21252 , RIf142c28_5219, \9058_9357 );
and \U$12123 ( \20954_21253 , RIe181038_2845, \9060_9359 );
and \U$12124 ( \20955_21254 , RIe17e338_2813, \9062_9361 );
and \U$12125 ( \20956_21255 , RIe17b638_2781, \9064_9363 );
and \U$12126 ( \20957_21256 , RIf1420e8_5211, \9066_9365 );
and \U$12127 ( \20958_21257 , RIf140a68_5195, \9068_9367 );
and \U$12128 ( \20959_21258 , RIf1401f8_5189, \9070_9369 );
and \U$12129 ( \20960_21259 , RIfebff10_8304, \9072_9371 );
and \U$12130 ( \20961_21260 , RIf13faf0_5184, \9074_9373 );
and \U$12131 ( \20962_21261 , RIf13ee48_5175, \9076_9375 );
and \U$12132 ( \20963_21262 , RIee3e2d8_5166, \9078_9377 );
and \U$12133 ( \20964_21263 , RIee3d1f8_5154, \9080_9379 );
and \U$12134 ( \20965_21264 , RIee3c118_5142, \9082_9381 );
and \U$12135 ( \20966_21265 , RIee3b038_5130, \9084_9383 );
and \U$12136 ( \20967_21266 , RIee39c88_5116, \9086_9385 );
and \U$12137 ( \20968_21267 , RIfe838f8_7841, \9088_9387 );
and \U$12138 ( \20969_21268 , RIf1701c8_5735, \9090_9389 );
and \U$12139 ( \20970_21269 , RIfc5ab00_6054, \9092_9391 );
and \U$12140 ( \20971_21270 , RIf16e008_5711, \9094_9393 );
and \U$12141 ( \20972_21271 , RIfcb0e88_7035, \9096_9395 );
and \U$12142 ( \20973_21272 , RIf16caf0_5696, \9098_9397 );
and \U$12143 ( \20974_21273 , RIe223590_4692, \9100_9399 );
and \U$12144 ( \20975_21274 , RIf16bce0_5686, \9102_9401 );
and \U$12145 ( \20976_21275 , RIe220890_4660, \9104_9403 );
and \U$12146 ( \20977_21276 , RIf16ac00_5674, \9106_9405 );
and \U$12147 ( \20978_21277 , RIe21db90_4628, \9108_9407 );
and \U$12148 ( \20979_21278 , RIe218190_4564, \9110_9409 );
and \U$12149 ( \20980_21279 , RIe215490_4532, \9112_9411 );
and \U$12150 ( \20981_21280 , RIf16a228_5667, \9114_9413 );
and \U$12151 ( \20982_21281 , RIe212790_4500, \9116_9415 );
and \U$12152 ( \20983_21282 , RIf168fe0_5654, \9118_9417 );
and \U$12153 ( \20984_21283 , RIe20fa90_4468, \9120_9419 );
and \U$12154 ( \20985_21284 , RIf167d98_5641, \9122_9421 );
and \U$12155 ( \20986_21285 , RIe20cd90_4436, \9124_9423 );
and \U$12156 ( \20987_21286 , RIe20a090_4404, \9126_9425 );
and \U$12157 ( \20988_21287 , RIe207390_4372, \9128_9427 );
and \U$12158 ( \20989_21288 , RIf1670f0_5632, \9130_9429 );
and \U$12159 ( \20990_21289 , RIf165ea8_5619, \9132_9431 );
and \U$12160 ( \20991_21290 , RIe202200_4314, \9134_9433 );
and \U$12161 ( \20992_21291 , RIfe83e98_7845, \9136_9435 );
and \U$12162 ( \20993_21292 , RIf164f30_5608, \9138_9437 );
and \U$12163 ( \20994_21293 , RIf1643f0_5600, \9140_9439 );
and \U$12164 ( \20995_21294 , RIfce8310_7664, \9142_9441 );
and \U$12165 ( \20996_21295 , RIf161df8_5573, \9144_9443 );
and \U$12166 ( \20997_21296 , RIf15ff08_5551, \9146_9445 );
and \U$12167 ( \20998_21297 , RIf15e018_5529, \9148_9447 );
and \U$12168 ( \20999_21298 , RIfe83d30_7844, \9150_9449 );
and \U$12169 ( \21000_21299 , RIfe84000_7846, \9152_9451 );
and \U$12170 ( \21001_21300 , RIf15cb00_5514, \9154_9453 );
and \U$12171 ( \21002_21301 , RIf15b5e8_5499, \9156_9455 );
and \U$12172 ( \21003_21302 , RIf15a508_5487, \9158_9457 );
and \U$12173 ( \21004_21303 , RIfc887a8_6575, \9160_9459 );
or \U$12174 ( \21005_21304 , \20941_21240 , \20942_21241 , \20943_21242 , \20944_21243 , \20945_21244 , \20946_21245 , \20947_21246 , \20948_21247 , \20949_21248 , \20950_21249 , \20951_21250 , \20952_21251 , \20953_21252 , \20954_21253 , \20955_21254 , \20956_21255 , \20957_21256 , \20958_21257 , \20959_21258 , \20960_21259 , \20961_21260 , \20962_21261 , \20963_21262 , \20964_21263 , \20965_21264 , \20966_21265 , \20967_21266 , \20968_21267 , \20969_21268 , \20970_21269 , \20971_21270 , \20972_21271 , \20973_21272 , \20974_21273 , \20975_21274 , \20976_21275 , \20977_21276 , \20978_21277 , \20979_21278 , \20980_21279 , \20981_21280 , \20982_21281 , \20983_21282 , \20984_21283 , \20985_21284 , \20986_21285 , \20987_21286 , \20988_21287 , \20989_21288 , \20990_21289 , \20991_21290 , \20992_21291 , \20993_21292 , \20994_21293 , \20995_21294 , \20996_21295 , \20997_21296 , \20998_21297 , \20999_21298 , \21000_21299 , \21001_21300 , \21002_21301 , \21003_21302 , \21004_21303 );
and \U$12175 ( \21006_21305 , RIf158d20_5470, \9163_9462 );
and \U$12176 ( \21007_21306 , RIf157970_5456, \9165_9464 );
and \U$12177 ( \21008_21307 , RIf156cc8_5447, \9167_9466 );
and \U$12178 ( \21009_21308 , RIfe84438_7849, \9169_9468 );
and \U$12179 ( \21010_21309 , RIf156020_5438, \9171_9470 );
and \U$12180 ( \21011_21310 , RIfc51fc8_5955, \9173_9472 );
and \U$12181 ( \21012_21311 , RIf154568_5419, \9175_9474 );
and \U$12182 ( \21013_21312 , RIe1f51e0_4166, \9177_9476 );
and \U$12183 ( \21014_21313 , RIf153050_5404, \9179_9478 );
and \U$12184 ( \21015_21314 , RIf1519d0_5388, \9181_9480 );
and \U$12185 ( \21016_21315 , RIf150788_5375, \9183_9482 );
and \U$12186 ( \21017_21316 , RIfe842d0_7848, \9185_9484 );
and \U$12187 ( \21018_21317 , RIf14f810_5364, \9187_9486 );
and \U$12188 ( \21019_21318 , RIf14eb68_5355, \9189_9488 );
and \U$12189 ( \21020_21319 , RIf14dd58_5345, \9191_9490 );
and \U$12190 ( \21021_21320 , RIfe84168_7847, \9193_9492 );
and \U$12191 ( \21022_21321 , RIe1eb2f8_4053, \9195_9494 );
and \U$12192 ( \21023_21322 , RIe1e85f8_4021, \9197_9496 );
and \U$12193 ( \21024_21323 , RIe1e58f8_3989, \9199_9498 );
and \U$12194 ( \21025_21324 , RIe1e2bf8_3957, \9201_9500 );
and \U$12195 ( \21026_21325 , RIe1dfef8_3925, \9203_9502 );
and \U$12196 ( \21027_21326 , RIe1dd1f8_3893, \9205_9504 );
and \U$12197 ( \21028_21327 , RIe1da4f8_3861, \9207_9506 );
and \U$12198 ( \21029_21328 , RIe1d77f8_3829, \9209_9508 );
and \U$12199 ( \21030_21329 , RIe1d1df8_3765, \9211_9510 );
and \U$12200 ( \21031_21330 , RIe1cf0f8_3733, \9213_9512 );
and \U$12201 ( \21032_21331 , RIe1cc3f8_3701, \9215_9514 );
and \U$12202 ( \21033_21332 , RIe1c96f8_3669, \9217_9516 );
and \U$12203 ( \21034_21333 , RIe1c69f8_3637, \9219_9518 );
and \U$12204 ( \21035_21334 , RIe1c3cf8_3605, \9221_9520 );
and \U$12205 ( \21036_21335 , RIe1c0ff8_3573, \9223_9522 );
and \U$12206 ( \21037_21336 , RIe1be2f8_3541, \9225_9524 );
and \U$12207 ( \21038_21337 , RIf14c840_5330, \9227_9526 );
and \U$12208 ( \21039_21338 , RIf14b5f8_5317, \9229_9528 );
and \U$12209 ( \21040_21339 , RIfe83a60_7842, \9231_9530 );
and \U$12210 ( \21041_21340 , RIfe849d8_7853, \9233_9532 );
and \U$12211 ( \21042_21341 , RIfc74168_6343, \9235_9534 );
and \U$12212 ( \21043_21342 , RIf149b40_5298, \9237_9536 );
and \U$12213 ( \21044_21343 , RIfe83bc8_7843, \9239_9538 );
and \U$12214 ( \21045_21344 , RIfe84708_7851, \9241_9540 );
and \U$12215 ( \21046_21345 , RIf148d30_5288, \9243_9542 );
and \U$12216 ( \21047_21346 , RIf147ae8_5275, \9245_9544 );
and \U$12217 ( \21048_21347 , RIfe84870_7852, \9247_9546 );
and \U$12218 ( \21049_21348 , RIe1b0900_3386, \9249_9548 );
and \U$12219 ( \21050_21349 , RIf146fa8_5267, \9251_9550 );
and \U$12220 ( \21051_21350 , RIf146300_5258, \9253_9552 );
and \U$12221 ( \21052_21351 , RIfe845a0_7850, \9255_9554 );
and \U$12222 ( \21053_21352 , RIfe83790_7840, \9257_9556 );
and \U$12223 ( \21054_21353 , RIe1a8638_3293, \9259_9558 );
and \U$12224 ( \21055_21354 , RIe1a5938_3261, \9261_9560 );
and \U$12225 ( \21056_21355 , RIe1a2c38_3229, \9263_9562 );
and \U$12226 ( \21057_21356 , RIe19ff38_3197, \9265_9564 );
and \U$12227 ( \21058_21357 , RIe18c438_2973, \9267_9566 );
and \U$12228 ( \21059_21358 , RIe178938_2749, \9269_9568 );
and \U$12229 ( \21060_21359 , RIe226290_4724, \9271_9570 );
and \U$12230 ( \21061_21360 , RIe21ae90_4596, \9273_9572 );
and \U$12231 ( \21062_21361 , RIe204690_4340, \9275_9574 );
and \U$12232 ( \21063_21362 , RIe1fe6f0_4272, \9277_9576 );
and \U$12233 ( \21064_21363 , RIe1f7aa8_4195, \9279_9578 );
and \U$12234 ( \21065_21364 , RIe1f05f0_4112, \9281_9580 );
and \U$12235 ( \21066_21365 , RIe1d4af8_3797, \9283_9582 );
and \U$12236 ( \21067_21366 , RIe1bb5f8_3509, \9285_9584 );
and \U$12237 ( \21068_21367 , RIe1ae470_3360, \9287_9586 );
and \U$12238 ( \21069_21368 , RIe170aa8_2659, \9289_9588 );
or \U$12239 ( \21070_21369 , \21006_21305 , \21007_21306 , \21008_21307 , \21009_21308 , \21010_21309 , \21011_21310 , \21012_21311 , \21013_21312 , \21014_21313 , \21015_21314 , \21016_21315 , \21017_21316 , \21018_21317 , \21019_21318 , \21020_21319 , \21021_21320 , \21022_21321 , \21023_21322 , \21024_21323 , \21025_21324 , \21026_21325 , \21027_21326 , \21028_21327 , \21029_21328 , \21030_21329 , \21031_21330 , \21032_21331 , \21033_21332 , \21034_21333 , \21035_21334 , \21036_21335 , \21037_21336 , \21038_21337 , \21039_21338 , \21040_21339 , \21041_21340 , \21042_21341 , \21043_21342 , \21044_21343 , \21045_21344 , \21046_21345 , \21047_21346 , \21048_21347 , \21049_21348 , \21050_21349 , \21051_21350 , \21052_21351 , \21053_21352 , \21054_21353 , \21055_21354 , \21056_21355 , \21057_21356 , \21058_21357 , \21059_21358 , \21060_21359 , \21061_21360 , \21062_21361 , \21063_21362 , \21064_21363 , \21065_21364 , \21066_21365 , \21067_21366 , \21068_21367 , \21069_21368 );
or \U$12240 ( \21071_21370 , \21005_21304 , \21070_21369 );
_DC \g399e/U$1 ( \21072 , \21071_21370 , \9298_9597 );
buf \U$12241 ( \21073_21372 , \21072 );
xor \U$12242 ( \21074_21373 , \20940_21239 , \21073_21372 );
and \U$12243 ( \21075_21374 , RIdec4e38_704, \8760_9059 );
and \U$12244 ( \21076_21375 , RIdec2138_672, \8762_9061 );
and \U$12245 ( \21077_21376 , RIee1fc48_4820, \8764_9063 );
and \U$12246 ( \21078_21377 , RIdebf438_640, \8766_9065 );
and \U$12247 ( \21079_21378 , RIfc49490_5856, \8768_9067 );
and \U$12248 ( \21080_21379 , RIdebc738_608, \8770_9069 );
and \U$12249 ( \21081_21380 , RIdeb9a38_576, \8772_9071 );
and \U$12250 ( \21082_21381 , RIdeb6d38_544, \8774_9073 );
and \U$12251 ( \21083_21382 , RIfc48ef0_5852, \8776_9075 );
and \U$12252 ( \21084_21383 , RIdeb1338_480, \8778_9077 );
and \U$12253 ( \21085_21384 , RIfcd9b08_7499, \8780_9079 );
and \U$12254 ( \21086_21385 , RIdeae638_448, \8782_9081 );
and \U$12255 ( \21087_21386 , RIfc8b610_6608, \8784_9083 );
and \U$12256 ( \21088_21387 , RIdea9700_416, \8786_9085 );
and \U$12257 ( \21089_21388 , RIdea2e00_384, \8788_9087 );
and \U$12258 ( \21090_21389 , RIde9c500_352, \8790_9089 );
and \U$12259 ( \21091_21390 , RIee1c9a8_4784, \8792_9091 );
and \U$12260 ( \21092_21391 , RIee1b8c8_4772, \8794_9093 );
and \U$12261 ( \21093_21392 , RIfc80918_6485, \8796_9095 );
and \U$12262 ( \21094_21393 , RIfcdad50_7512, \8798_9097 );
and \U$12263 ( \21095_21394 , RIfe86e68_7879, \8800_9099 );
and \U$12264 ( \21096_21395 , RIde8cee8_277, \8802_9101 );
and \U$12265 ( \21097_21396 , RIfe86d00_7878, \8804_9103 );
and \U$12266 ( \21098_21397 , RIfec0d20_8314, \8806_9105 );
and \U$12267 ( \21099_21398 , RIde81098_219, \8808_9107 );
and \U$12268 ( \21100_21399 , RIfc8b8e0_6610, \8810_9109 );
and \U$12269 ( \21101_21400 , RIfcd2d58_7421, \8812_9111 );
and \U$12270 ( \21102_21401 , RIfce4530_7620, \8814_9113 );
and \U$12271 ( \21103_21402 , RIfc8ba48_6611, \8816_9115 );
and \U$12272 ( \21104_21403 , RIe16b210_2596, \8818_9117 );
and \U$12273 ( \21105_21404 , RIe1698c0_2578, \8820_9119 );
and \U$12274 ( \21106_21405 , RIe1679d0_2556, \8822_9121 );
and \U$12275 ( \21107_21406 , RIe164e38_2525, \8824_9123 );
and \U$12276 ( \21108_21407 , RIe162138_2493, \8826_9125 );
and \U$12277 ( \21109_21408 , RIee370f0_5085, \8828_9127 );
and \U$12278 ( \21110_21409 , RIe15f438_2461, \8830_9129 );
and \U$12279 ( \21111_21410 , RIfc999e0_6770, \8832_9131 );
and \U$12280 ( \21112_21411 , RIe15c738_2429, \8834_9133 );
and \U$12281 ( \21113_21412 , RIe156d38_2365, \8836_9135 );
and \U$12282 ( \21114_21413 , RIe154038_2333, \8838_9137 );
and \U$12283 ( \21115_21414 , RIfc3f260_5744, \8840_9139 );
and \U$12284 ( \21116_21415 , RIe151338_2301, \8842_9141 );
and \U$12285 ( \21117_21416 , RIfc48518_5845, \8844_9143 );
and \U$12286 ( \21118_21417 , RIe14e638_2269, \8846_9145 );
and \U$12287 ( \21119_21418 , RIfc99e18_6773, \8848_9147 );
and \U$12288 ( \21120_21419 , RIe14b938_2237, \8850_9149 );
and \U$12289 ( \21121_21420 , RIe148c38_2205, \8852_9151 );
and \U$12290 ( \21122_21421 , RIe145f38_2173, \8854_9153 );
and \U$12291 ( \21123_21422 , RIee34288_5052, \8856_9155 );
and \U$12292 ( \21124_21423 , RIee33040_5039, \8858_9157 );
and \U$12293 ( \21125_21424 , RIee31f60_5027, \8860_9159 );
and \U$12294 ( \21126_21425 , RIfcd99a0_7498, \8862_9161 );
and \U$12295 ( \21127_21426 , RIfe86b98_7877, \8864_9163 );
and \U$12296 ( \21128_21427 , RIdf3e9e0_2089, \8866_9165 );
and \U$12297 ( \21129_21428 , RIfe86a30_7876, \8868_9167 );
and \U$12298 ( \21130_21429 , RIdf3a4f8_2040, \8870_9169 );
and \U$12299 ( \21131_21430 , RIfcc3470_7244, \8872_9171 );
and \U$12300 ( \21132_21431 , RIee2f530_4997, \8874_9173 );
and \U$12301 ( \21133_21432 , RIfc7fdd8_6477, \8876_9175 );
and \U$12302 ( \21134_21433 , RIee2d370_4973, \8878_9177 );
and \U$12303 ( \21135_21434 , RIdf35200_1981, \8880_9179 );
and \U$12304 ( \21136_21435 , RIfec0ff0_8316, \8882_9181 );
and \U$12305 ( \21137_21436 , RIdf30d18_1932, \8884_9183 );
and \U$12306 ( \21138_21437 , RIfec0e88_8315, \8886_9185 );
or \U$12307 ( \21139_21438 , \21075_21374 , \21076_21375 , \21077_21376 , \21078_21377 , \21079_21378 , \21080_21379 , \21081_21380 , \21082_21381 , \21083_21382 , \21084_21383 , \21085_21384 , \21086_21385 , \21087_21386 , \21088_21387 , \21089_21388 , \21090_21389 , \21091_21390 , \21092_21391 , \21093_21392 , \21094_21393 , \21095_21394 , \21096_21395 , \21097_21396 , \21098_21397 , \21099_21398 , \21100_21399 , \21101_21400 , \21102_21401 , \21103_21402 , \21104_21403 , \21105_21404 , \21106_21405 , \21107_21406 , \21108_21407 , \21109_21408 , \21110_21409 , \21111_21410 , \21112_21411 , \21113_21412 , \21114_21413 , \21115_21414 , \21116_21415 , \21117_21416 , \21118_21417 , \21119_21418 , \21120_21419 , \21121_21420 , \21122_21421 , \21123_21422 , \21124_21423 , \21125_21424 , \21126_21425 , \21127_21426 , \21128_21427 , \21129_21428 , \21130_21429 , \21131_21430 , \21132_21431 , \21133_21432 , \21134_21433 , \21135_21434 , \21136_21435 , \21137_21436 , \21138_21437 );
and \U$12308 ( \21140_21439 , RIfcd2a88_7419, \8889_9188 );
and \U$12309 ( \21141_21440 , RIfc8c858_6621, \8891_9190 );
and \U$12310 ( \21142_21441 , RIfc47ca8_5839, \8893_9192 );
and \U$12311 ( \21143_21442 , RIfcd6430_7460, \8895_9194 );
and \U$12312 ( \21144_21443 , RIdf29f68_1854, \8897_9196 );
and \U$12313 ( \21145_21444 , RIdf27da8_1830, \8899_9198 );
and \U$12314 ( \21146_21445 , RIdf26188_1810, \8901_9200 );
and \U$12315 ( \21147_21446 , RIdf24568_1790, \8903_9202 );
and \U$12316 ( \21148_21447 , RIfc8cb28_6623, \8905_9204 );
and \U$12317 ( \21149_21448 , RIfcdb188_7515, \8907_9206 );
and \U$12318 ( \21150_21449 , RIdf22948_1770, \8909_9208 );
and \U$12319 ( \21151_21450 , RIfc475a0_5834, \8911_9210 );
and \U$12320 ( \21152_21451 , RIdf21430_1755, \8913_9212 );
and \U$12321 ( \21153_21452 , RIdf1f3d8_1732, \8915_9214 );
and \U$12322 ( \21154_21453 , RIfec0bb8_8313, \8917_9216 );
and \U$12323 ( \21155_21454 , RIfe868c8_7875, \8919_9218 );
and \U$12324 ( \21156_21455 , RIdf16a08_1634, \8921_9220 );
and \U$12325 ( \21157_21456 , RIdf13d08_1602, \8923_9222 );
and \U$12326 ( \21158_21457 , RIdf11008_1570, \8925_9224 );
and \U$12327 ( \21159_21458 , RIdf0e308_1538, \8927_9226 );
and \U$12328 ( \21160_21459 , RIdf0b608_1506, \8929_9228 );
and \U$12329 ( \21161_21460 , RIdf08908_1474, \8931_9230 );
and \U$12330 ( \21162_21461 , RIdf05c08_1442, \8933_9232 );
and \U$12331 ( \21163_21462 , RIdf02f08_1410, \8935_9234 );
and \U$12332 ( \21164_21463 , RIdefd508_1346, \8937_9236 );
and \U$12333 ( \21165_21464 , RIdefa808_1314, \8939_9238 );
and \U$12334 ( \21166_21465 , RIdef7b08_1282, \8941_9240 );
and \U$12335 ( \21167_21466 , RIdef4e08_1250, \8943_9242 );
and \U$12336 ( \21168_21467 , RIdef2108_1218, \8945_9244 );
and \U$12337 ( \21169_21468 , RIdeef408_1186, \8947_9246 );
and \U$12338 ( \21170_21469 , RIdeec708_1154, \8949_9248 );
and \U$12339 ( \21171_21470 , RIdee9a08_1122, \8951_9250 );
and \U$12340 ( \21172_21471 , RIee254e0_4883, \8953_9252 );
and \U$12341 ( \21173_21472 , RIee246d0_4873, \8955_9254 );
and \U$12342 ( \21174_21473 , RIee23b90_4865, \8957_9256 );
and \U$12343 ( \21175_21474 , RIee231b8_4858, \8959_9258 );
and \U$12344 ( \21176_21475 , RIfe86fd0_7880, \8961_9260 );
and \U$12345 ( \21177_21476 , RIdee2820_1041, \8963_9262 );
and \U$12346 ( \21178_21477 , RIdee0930_1019, \8965_9264 );
and \U$12347 ( \21179_21478 , RIdede608_994, \8967_9266 );
and \U$12348 ( \21180_21479 , RIfc55da8_5999, \8969_9268 );
and \U$12349 ( \21181_21480 , RIfc98a68_6759, \8971_9270 );
and \U$12350 ( \21182_21481 , RIfcc3038_7241, \8973_9272 );
and \U$12351 ( \21183_21482 , RIfc464c0_5822, \8975_9274 );
and \U$12352 ( \21184_21483 , RIded9310_935, \8977_9276 );
and \U$12353 ( \21185_21484 , RIded6e80_909, \8979_9278 );
and \U$12354 ( \21186_21485 , RIded4f90_887, \8981_9280 );
and \U$12355 ( \21187_21486 , RIded2b00_861, \8983_9282 );
and \U$12356 ( \21188_21487 , RIded0238_832, \8985_9284 );
and \U$12357 ( \21189_21488 , RIdecd538_800, \8987_9286 );
and \U$12358 ( \21190_21489 , RIdeca838_768, \8989_9288 );
and \U$12359 ( \21191_21490 , RIdec7b38_736, \8991_9290 );
and \U$12360 ( \21192_21491 , RIdeb4038_512, \8993_9292 );
and \U$12361 ( \21193_21492 , RIde95c00_320, \8995_9294 );
and \U$12362 ( \21194_21493 , RIe16dc40_2626, \8997_9296 );
and \U$12363 ( \21195_21494 , RIe159a38_2397, \8999_9298 );
and \U$12364 ( \21196_21495 , RIe143238_2141, \9001_9300 );
and \U$12365 ( \21197_21496 , RIdf37c30_2011, \9003_9302 );
and \U$12366 ( \21198_21497 , RIdf2c290_1879, \9005_9304 );
and \U$12367 ( \21199_21498 , RIdf1cb10_1703, \9007_9306 );
and \U$12368 ( \21200_21499 , RIdf00208_1378, \9009_9308 );
and \U$12369 ( \21201_21500 , RIdee6d08_1090, \9011_9310 );
and \U$12370 ( \21202_21501 , RIdedba70_963, \9013_9312 );
and \U$12371 ( \21203_21502 , RIde7bb48_193, \9015_9314 );
or \U$12372 ( \21204_21503 , \21140_21439 , \21141_21440 , \21142_21441 , \21143_21442 , \21144_21443 , \21145_21444 , \21146_21445 , \21147_21446 , \21148_21447 , \21149_21448 , \21150_21449 , \21151_21450 , \21152_21451 , \21153_21452 , \21154_21453 , \21155_21454 , \21156_21455 , \21157_21456 , \21158_21457 , \21159_21458 , \21160_21459 , \21161_21460 , \21162_21461 , \21163_21462 , \21164_21463 , \21165_21464 , \21166_21465 , \21167_21466 , \21168_21467 , \21169_21468 , \21170_21469 , \21171_21470 , \21172_21471 , \21173_21472 , \21174_21473 , \21175_21474 , \21176_21475 , \21177_21476 , \21178_21477 , \21179_21478 , \21180_21479 , \21181_21480 , \21182_21481 , \21183_21482 , \21184_21483 , \21185_21484 , \21186_21485 , \21187_21486 , \21188_21487 , \21189_21488 , \21190_21489 , \21191_21490 , \21192_21491 , \21193_21492 , \21194_21493 , \21195_21494 , \21196_21495 , \21197_21496 , \21198_21497 , \21199_21498 , \21200_21499 , \21201_21500 , \21202_21501 , \21203_21502 );
or \U$12373 ( \21205_21504 , \21139_21438 , \21204_21503 );
_DC \g28f6/U$1 ( \21206 , \21205_21504 , \9024_9323 );
buf \U$12374 ( \21207_21506 , \21206 );
and \U$12375 ( \21208_21507 , RIe19d0d0_3164, \9034_9333 );
and \U$12376 ( \21209_21508 , RIe19a3d0_3132, \9036_9335 );
and \U$12377 ( \21210_21509 , RIf1454f0_5248, \9038_9337 );
and \U$12378 ( \21211_21510 , RIe1976d0_3100, \9040_9339 );
and \U$12379 ( \21212_21511 , RIf144578_5237, \9042_9341 );
and \U$12380 ( \21213_21512 , RIe1949d0_3068, \9044_9343 );
and \U$12381 ( \21214_21513 , RIe191cd0_3036, \9046_9345 );
and \U$12382 ( \21215_21514 , RIe18efd0_3004, \9048_9347 );
and \U$12383 ( \21216_21515 , RIe1895d0_2940, \9050_9349 );
and \U$12384 ( \21217_21516 , RIe1868d0_2908, \9052_9351 );
and \U$12385 ( \21218_21517 , RIf143498_5225, \9054_9353 );
and \U$12386 ( \21219_21518 , RIe183bd0_2876, \9056_9355 );
and \U$12387 ( \21220_21519 , RIfc51758_5949, \9058_9357 );
and \U$12388 ( \21221_21520 , RIe180ed0_2844, \9060_9359 );
and \U$12389 ( \21222_21521 , RIe17e1d0_2812, \9062_9361 );
and \U$12390 ( \21223_21522 , RIe17b4d0_2780, \9064_9363 );
and \U$12391 ( \21224_21523 , RIfc9b060_6786, \9066_9365 );
and \U$12392 ( \21225_21524 , RIfc9ee40_6830, \9068_9367 );
and \U$12393 ( \21226_21525 , RIe176e80_2730, \9070_9369 );
and \U$12394 ( \21227_21526 , RIe175800_2714, \9072_9371 );
and \U$12395 ( \21228_21527 , RIfcb70f8_7105, \9074_9373 );
and \U$12396 ( \21229_21528 , RIfce0cf0_7580, \9076_9375 );
and \U$12397 ( \21230_21529 , RIfcc4280_7254, \9078_9377 );
and \U$12398 ( \21231_21530 , RIfcba7d0_7144, \9080_9379 );
and \U$12399 ( \21232_21531 , RIee3bfb0_5141, \9082_9381 );
and \U$12400 ( \21233_21532 , RIee3aed0_5129, \9084_9383 );
and \U$12401 ( \21234_21533 , RIee39b20_5115, \9086_9385 );
and \U$12402 ( \21235_21534 , RIe173370_2688, \9088_9387 );
and \U$12403 ( \21236_21535 , RIf170060_5734, \9090_9389 );
and \U$12404 ( \21237_21536 , RIf16f3b8_5725, \9092_9391 );
and \U$12405 ( \21238_21537 , RIf16dea0_5710, \9094_9393 );
and \U$12406 ( \21239_21538 , RIf16d4c8_5703, \9096_9395 );
and \U$12407 ( \21240_21539 , RIf16c988_5695, \9098_9397 );
and \U$12408 ( \21241_21540 , RIe223428_4691, \9100_9399 );
and \U$12409 ( \21242_21541 , RIf16bb78_5685, \9102_9401 );
and \U$12410 ( \21243_21542 , RIe220728_4659, \9104_9403 );
and \U$12411 ( \21244_21543 , RIf16aa98_5673, \9106_9405 );
and \U$12412 ( \21245_21544 , RIe21da28_4627, \9108_9407 );
and \U$12413 ( \21246_21545 , RIe218028_4563, \9110_9409 );
and \U$12414 ( \21247_21546 , RIe215328_4531, \9112_9411 );
and \U$12415 ( \21248_21547 , RIf16a0c0_5666, \9114_9413 );
and \U$12416 ( \21249_21548 , RIe212628_4499, \9116_9415 );
and \U$12417 ( \21250_21549 , RIf168e78_5653, \9118_9417 );
and \U$12418 ( \21251_21550 , RIe20f928_4467, \9120_9419 );
and \U$12419 ( \21252_21551 , RIf167c30_5640, \9122_9421 );
and \U$12420 ( \21253_21552 , RIe20cc28_4435, \9124_9423 );
and \U$12421 ( \21254_21553 , RIe209f28_4403, \9126_9425 );
and \U$12422 ( \21255_21554 , RIe207228_4371, \9128_9427 );
and \U$12423 ( \21256_21555 , RIf166f88_5631, \9130_9429 );
and \U$12424 ( \21257_21556 , RIf165d40_5618, \9132_9431 );
and \U$12425 ( \21258_21557 , RIfec0618_8309, \9134_9433 );
and \U$12426 ( \21259_21558 , RIfe86760_7874, \9136_9435 );
and \U$12427 ( \21260_21559 , RIfc52b08_5963, \9138_9437 );
and \U$12428 ( \21261_21560 , RIf164288_5599, \9140_9439 );
and \U$12429 ( \21262_21561 , RIf163310_5588, \9142_9441 );
and \U$12430 ( \21263_21562 , RIf161c90_5572, \9144_9443 );
and \U$12431 ( \21264_21563 , RIf15fda0_5550, \9146_9445 );
and \U$12432 ( \21265_21564 , RIf15deb0_5528, \9148_9447 );
and \U$12433 ( \21266_21565 , RIfe865f8_7873, \9150_9449 );
and \U$12434 ( \21267_21566 , RIfe85d88_7867, \9152_9451 );
and \U$12435 ( \21268_21567 , RIf15c998_5513, \9154_9453 );
and \U$12436 ( \21269_21568 , RIf15b480_5498, \9156_9455 );
and \U$12437 ( \21270_21569 , RIf15a3a0_5486, \9158_9457 );
and \U$12438 ( \21271_21570 , RIf159b30_5480, \9160_9459 );
or \U$12439 ( \21272_21571 , \21208_21507 , \21209_21508 , \21210_21509 , \21211_21510 , \21212_21511 , \21213_21512 , \21214_21513 , \21215_21514 , \21216_21515 , \21217_21516 , \21218_21517 , \21219_21518 , \21220_21519 , \21221_21520 , \21222_21521 , \21223_21522 , \21224_21523 , \21225_21524 , \21226_21525 , \21227_21526 , \21228_21527 , \21229_21528 , \21230_21529 , \21231_21530 , \21232_21531 , \21233_21532 , \21234_21533 , \21235_21534 , \21236_21535 , \21237_21536 , \21238_21537 , \21239_21538 , \21240_21539 , \21241_21540 , \21242_21541 , \21243_21542 , \21244_21543 , \21245_21544 , \21246_21545 , \21247_21546 , \21248_21547 , \21249_21548 , \21250_21549 , \21251_21550 , \21252_21551 , \21253_21552 , \21254_21553 , \21255_21554 , \21256_21555 , \21257_21556 , \21258_21557 , \21259_21558 , \21260_21559 , \21261_21560 , \21262_21561 , \21263_21562 , \21264_21563 , \21265_21564 , \21266_21565 , \21267_21566 , \21268_21567 , \21269_21568 , \21270_21569 , \21271_21570 );
and \U$12440 ( \21273_21572 , RIfc83348_6515, \9163_9462 );
and \U$12441 ( \21274_21573 , RIfc4ade0_5874, \9165_9464 );
and \U$12442 ( \21275_21574 , RIfc89720_6586, \9167_9466 );
and \U$12443 ( \21276_21575 , RIe1f9f38_4221, \9169_9468 );
and \U$12444 ( \21277_21576 , RIfc4ac78_5873, \9171_9470 );
and \U$12445 ( \21278_21577 , RIfc9f110_6832, \9173_9472 );
and \U$12446 ( \21279_21578 , RIfc4ab10_5872, \9175_9474 );
and \U$12447 ( \21280_21579 , RIe1f5078_4165, \9177_9476 );
and \U$12448 ( \21281_21580 , RIf152ee8_5403, \9179_9478 );
and \U$12449 ( \21282_21581 , RIfc899f0_6588, \9181_9480 );
and \U$12450 ( \21283_21582 , RIf150620_5374, \9183_9482 );
and \U$12451 ( \21284_21583 , RIe1f2eb8_4141, \9185_9484 );
and \U$12452 ( \21285_21584 , RIf14f6a8_5363, \9187_9486 );
and \U$12453 ( \21286_21585 , RIf14ea00_5354, \9189_9488 );
and \U$12454 ( \21287_21586 , RIf14dbf0_5344, \9191_9490 );
and \U$12455 ( \21288_21587 , RIe1edbc0_4082, \9193_9492 );
and \U$12456 ( \21289_21588 , RIe1eb190_4052, \9195_9494 );
and \U$12457 ( \21290_21589 , RIe1e8490_4020, \9197_9496 );
and \U$12458 ( \21291_21590 , RIe1e5790_3988, \9199_9498 );
and \U$12459 ( \21292_21591 , RIe1e2a90_3956, \9201_9500 );
and \U$12460 ( \21293_21592 , RIe1dfd90_3924, \9203_9502 );
and \U$12461 ( \21294_21593 , RIe1dd090_3892, \9205_9504 );
and \U$12462 ( \21295_21594 , RIe1da390_3860, \9207_9506 );
and \U$12463 ( \21296_21595 , RIe1d7690_3828, \9209_9508 );
and \U$12464 ( \21297_21596 , RIe1d1c90_3764, \9211_9510 );
and \U$12465 ( \21298_21597 , RIe1cef90_3732, \9213_9512 );
and \U$12466 ( \21299_21598 , RIe1cc290_3700, \9215_9514 );
and \U$12467 ( \21300_21599 , RIe1c9590_3668, \9217_9516 );
and \U$12468 ( \21301_21600 , RIe1c6890_3636, \9219_9518 );
and \U$12469 ( \21302_21601 , RIe1c3b90_3604, \9221_9520 );
and \U$12470 ( \21303_21602 , RIe1c0e90_3572, \9223_9522 );
and \U$12471 ( \21304_21603 , RIe1be190_3540, \9225_9524 );
and \U$12472 ( \21305_21604 , RIf14c6d8_5329, \9227_9526 );
and \U$12473 ( \21306_21605 , RIf14b490_5316, \9229_9528 );
and \U$12474 ( \21307_21606 , RIfe85ef0_7868, \9231_9530 );
and \U$12475 ( \21308_21607 , RIfe86490_7872, \9233_9532 );
and \U$12476 ( \21309_21608 , RIf14a248_5303, \9235_9534 );
and \U$12477 ( \21310_21609 , RIfc819f8_6497, \9237_9536 );
and \U$12478 ( \21311_21610 , RIfec0a50_8312, \9239_9538 );
and \U$12479 ( \21312_21611 , RIfe861c0_7870, \9241_9540 );
and \U$12480 ( \21313_21612 , RIf148bc8_5287, \9243_9542 );
and \U$12481 ( \21314_21613 , RIf147980_5274, \9245_9544 );
and \U$12482 ( \21315_21614 , RIfe86328_7871, \9247_9546 );
and \U$12483 ( \21316_21615 , RIfec0780_8310, \9249_9548 );
and \U$12484 ( \21317_21616 , RIfcbb478_7153, \9251_9550 );
and \U$12485 ( \21318_21617 , RIf146198_5257, \9253_9552 );
and \U$12486 ( \21319_21618 , RIfe86058_7869, \9255_9554 );
and \U$12487 ( \21320_21619 , RIfec08e8_8311, \9257_9556 );
and \U$12488 ( \21321_21620 , RIe1a84d0_3292, \9259_9558 );
and \U$12489 ( \21322_21621 , RIe1a57d0_3260, \9261_9560 );
and \U$12490 ( \21323_21622 , RIe1a2ad0_3228, \9263_9562 );
and \U$12491 ( \21324_21623 , RIe19fdd0_3196, \9265_9564 );
and \U$12492 ( \21325_21624 , RIe18c2d0_2972, \9267_9566 );
and \U$12493 ( \21326_21625 , RIe1787d0_2748, \9269_9568 );
and \U$12494 ( \21327_21626 , RIe226128_4723, \9271_9570 );
and \U$12495 ( \21328_21627 , RIe21ad28_4595, \9273_9572 );
and \U$12496 ( \21329_21628 , RIe204528_4339, \9275_9574 );
and \U$12497 ( \21330_21629 , RIe1fe588_4271, \9277_9576 );
and \U$12498 ( \21331_21630 , RIe1f7940_4194, \9279_9578 );
and \U$12499 ( \21332_21631 , RIe1f0488_4111, \9281_9580 );
and \U$12500 ( \21333_21632 , RIe1d4990_3796, \9283_9582 );
and \U$12501 ( \21334_21633 , RIe1bb490_3508, \9285_9584 );
and \U$12502 ( \21335_21634 , RIe1ae308_3359, \9287_9586 );
and \U$12503 ( \21336_21635 , RIe170940_2658, \9289_9588 );
or \U$12504 ( \21337_21636 , \21273_21572 , \21274_21573 , \21275_21574 , \21276_21575 , \21277_21576 , \21278_21577 , \21279_21578 , \21280_21579 , \21281_21580 , \21282_21581 , \21283_21582 , \21284_21583 , \21285_21584 , \21286_21585 , \21287_21586 , \21288_21587 , \21289_21588 , \21290_21589 , \21291_21590 , \21292_21591 , \21293_21592 , \21294_21593 , \21295_21594 , \21296_21595 , \21297_21596 , \21298_21597 , \21299_21598 , \21300_21599 , \21301_21600 , \21302_21601 , \21303_21602 , \21304_21603 , \21305_21604 , \21306_21605 , \21307_21606 , \21308_21607 , \21309_21608 , \21310_21609 , \21311_21610 , \21312_21611 , \21313_21612 , \21314_21613 , \21315_21614 , \21316_21615 , \21317_21616 , \21318_21617 , \21319_21618 , \21320_21619 , \21321_21620 , \21322_21621 , \21323_21622 , \21324_21623 , \21325_21624 , \21326_21625 , \21327_21626 , \21328_21627 , \21329_21628 , \21330_21629 , \21331_21630 , \21332_21631 , \21333_21632 , \21334_21633 , \21335_21634 , \21336_21635 );
or \U$12505 ( \21338_21637 , \21272_21571 , \21337_21636 );
_DC \g3a23/U$1 ( \21339 , \21338_21637 , \9298_9597 );
buf \U$12506 ( \21340_21639 , \21339 );
and \U$12507 ( \21341_21640 , \21207_21506 , \21340_21639 );
and \U$12508 ( \21342_21641 , \19437_19736 , \19570_19869 );
and \U$12509 ( \21343_21642 , \19570_19869 , \19845_20144 );
and \U$12510 ( \21344_21643 , \19437_19736 , \19845_20144 );
or \U$12511 ( \21345_21644 , \21342_21641 , \21343_21642 , \21344_21643 );
and \U$12512 ( \21346_21645 , \21340_21639 , \21345_21644 );
and \U$12513 ( \21347_21646 , \21207_21506 , \21345_21644 );
or \U$12514 ( \21348_21647 , \21341_21640 , \21346_21645 , \21347_21646 );
xor \U$12515 ( \21349_21648 , \21074_21373 , \21348_21647 );
buf g441e_GF_PartitionCandidate( \21350_21649_nG441e , \21349_21648 );
xor \U$12516 ( \21351_21650 , \21207_21506 , \21340_21639 );
xor \U$12517 ( \21352_21651 , \21351_21650 , \21345_21644 );
buf g4421_GF_PartitionCandidate( \21353_21652_nG4421 , \21352_21651 );
nand \U$12518 ( \21354_21653 , \21353_21652_nG4421 , \19847_20146_nG4424 );
and \U$12519 ( \21355_21654 , \21350_21649_nG441e , \21354_21653 );
xor \U$12520 ( \21356_21655 , \21353_21652_nG4421 , \19847_20146_nG4424 );
and \U$12525 ( \21357_21659 , \21356_21655 , \10392_10694_nG9c0e );
or \U$12526 ( \21358_21660 , 1'b0 , \21357_21659 );
xor \U$12527 ( \21359_21661 , \21355_21654 , \21358_21660 );
xor \U$12528 ( \21360_21662 , \21355_21654 , \21359_21661 );
buf \U$12529 ( \21361_21663 , \21360_21662 );
buf \U$12530 ( \21362_21664 , \21361_21663 );
xor \U$12531 ( \21363_21665 , \20807_21106 , \21362_21664 );
and \U$12532 ( \21364_21666 , \20396_20695 , \20794_21093 );
and \U$12533 ( \21365_21667 , \20396_20695 , \20800_21099 );
and \U$12534 ( \21366_21668 , \20794_21093 , \20800_21099 );
or \U$12535 ( \21367_21669 , \21364_21666 , \21365_21667 , \21366_21668 );
and \U$12536 ( \21368_21670 , \21363_21665 , \21367_21669 );
and \U$12537 ( \21369_21671 , \20416_20715 , \20422_20721 );
and \U$12538 ( \21370_21672 , \20416_20715 , \20792_21091 );
and \U$12539 ( \21371_21673 , \20422_20721 , \20792_21091 );
or \U$12540 ( \21372_21674 , \21369_21671 , \21370_21672 , \21371_21673 );
buf \U$12541 ( \21373_21675 , \21372_21674 );
and \U$12542 ( \21374_21676 , \20350_20652 , \20359_20658 );
and \U$12543 ( \21375_21677 , \20350_20652 , \20366_20665 );
and \U$12544 ( \21376_21678 , \20359_20658 , \20366_20665 );
or \U$12545 ( \21377_21679 , \21374_21676 , \21375_21677 , \21376_21678 );
buf \U$12546 ( \21378_21680 , \21377_21679 );
and \U$12547 ( \21379_21681 , \16405_15940 , \13771_14070_nG9bf9 );
and \U$12548 ( \21380_21682 , \15638_15937 , \14682_14984_nG9bf6 );
or \U$12549 ( \21381_21683 , \21379_21681 , \21380_21682 );
xor \U$12550 ( \21382_21684 , \15637_15936 , \21381_21683 );
buf \U$12551 ( \21383_21685 , \21382_21684 );
buf \U$12553 ( \21384_21686 , \21383_21685 );
xor \U$12554 ( \21385_21687 , \21378_21680 , \21384_21686 );
and \U$12555 ( \21386_21688 , \14710_14631 , \15074_15373_nG9bf3 );
and \U$12556 ( \21387_21689 , \14329_14628 , \16013_16315_nG9bf0 );
or \U$12557 ( \21388_21690 , \21386_21688 , \21387_21689 );
xor \U$12558 ( \21389_21691 , \14328_14627 , \21388_21690 );
buf \U$12559 ( \21390_21692 , \21389_21691 );
buf \U$12561 ( \21391_21693 , \21390_21692 );
xor \U$12562 ( \21392_21694 , \21385_21687 , \21391_21693 );
buf \U$12563 ( \21393_21695 , \21392_21694 );
and \U$12564 ( \21394_21696 , \20368_20667 , \20370_20669 );
and \U$12565 ( \21395_21697 , \20368_20667 , \20377_20676 );
and \U$12566 ( \21396_21698 , \20370_20669 , \20377_20676 );
or \U$12567 ( \21397_21699 , \21394_21696 , \21395_21697 , \21396_21698 );
buf \U$12568 ( \21398_21700 , \21397_21699 );
xor \U$12569 ( \21399_21701 , \21393_21695 , \21398_21700 );
and \U$12570 ( \21400_21702 , \10996_10421 , \19287_19586_nG9be1 );
and \U$12571 ( \21401_21703 , \10119_10418 , \20306_20608_nG9bde );
or \U$12572 ( \21402_21704 , \21400_21702 , \21401_21703 );
xor \U$12573 ( \21403_21705 , \10118_10417 , \21402_21704 );
buf \U$12574 ( \21404_21706 , \21403_21705 );
buf \U$12576 ( \21405_21707 , \21404_21706 );
xor \U$12577 ( \21406_21708 , \21399_21701 , \21405_21707 );
buf \U$12578 ( \21407_21709 , \21406_21708 );
xor \U$12579 ( \21408_21710 , \21373_21675 , \21407_21709 );
and \U$12580 ( \21409_21711 , \20353_20155 , \10693_10995_nG9c0b );
and \U$12581 ( \21410_21712 , \19853_20152 , \10981_11283_nG9c08 );
or \U$12582 ( \21411_21713 , \21409_21711 , \21410_21712 );
xor \U$12583 ( \21412_21714 , \19852_20151 , \21411_21713 );
buf \U$12584 ( \21413_21715 , \21412_21714 );
buf \U$12586 ( \21414_21716 , \21413_21715 );
and \U$12587 ( \21415_21717 , \18908_18702 , \11299_11598_nG9c05 );
and \U$12588 ( \21416_21718 , \18400_18699 , \12168_12470_nG9c02 );
or \U$12589 ( \21417_21719 , \21415_21717 , \21416_21718 );
xor \U$12590 ( \21418_21720 , \18399_18698 , \21417_21719 );
buf \U$12591 ( \21419_21721 , \21418_21720 );
buf \U$12593 ( \21420_21722 , \21419_21721 );
xor \U$12594 ( \21421_21723 , \21414_21716 , \21420_21722 );
buf \U$12595 ( \21422_21724 , \21421_21723 );
and \U$12596 ( \21423_21725 , \20342_20644 , \20348_20650 );
buf \U$12597 ( \21424_21726 , \21423_21725 );
xor \U$12598 ( \21425_21727 , \21422_21724 , \21424_21726 );
and \U$12599 ( \21426_21728 , \17437_17297 , \12502_12801_nG9bff );
and \U$12600 ( \21427_21729 , \16995_17294 , \13403_13705_nG9bfc );
or \U$12601 ( \21428_21730 , \21426_21728 , \21427_21729 );
xor \U$12602 ( \21429_21731 , \16994_17293 , \21428_21730 );
buf \U$12603 ( \21430_21732 , \21429_21731 );
buf \U$12605 ( \21431_21733 , \21430_21732 );
xor \U$12606 ( \21432_21734 , \21425_21727 , \21431_21733 );
buf \U$12607 ( \21433_21735 , \21432_21734 );
and \U$12608 ( \21434_21736 , \13431_13370 , \16378_16680_nG9bed );
and \U$12609 ( \21435_21737 , \13068_13367 , \17363_17665_nG9bea );
or \U$12610 ( \21436_21738 , \21434_21736 , \21435_21737 );
xor \U$12611 ( \21437_21739 , \13067_13366 , \21436_21738 );
buf \U$12612 ( \21438_21740 , \21437_21739 );
buf \U$12614 ( \21439_21741 , \21438_21740 );
xor \U$12615 ( \21440_21742 , \21433_21735 , \21439_21741 );
and \U$12616 ( \21441_21743 , \12183_12157 , \17808_18107_nG9be7 );
and \U$12617 ( \21442_21744 , \11855_12154 , \18789_19091_nG9be4 );
or \U$12618 ( \21443_21745 , \21441_21743 , \21442_21744 );
xor \U$12619 ( \21444_21746 , \11854_12153 , \21443_21745 );
buf \U$12620 ( \21445_21747 , \21444_21746 );
buf \U$12622 ( \21446_21748 , \21445_21747 );
xor \U$12623 ( \21447_21749 , \21440_21742 , \21446_21748 );
buf \U$12624 ( \21448_21750 , \21447_21749 );
xor \U$12625 ( \21449_21751 , \21408_21710 , \21448_21750 );
buf \U$12626 ( \21450_21752 , \21449_21751 );
and \U$12627 ( \21451_21753 , \20334_20636 , \20388_20687 );
and \U$12628 ( \21452_21754 , \20334_20636 , \20394_20693 );
and \U$12629 ( \21453_21755 , \20388_20687 , \20394_20693 );
or \U$12630 ( \21454_21756 , \21451_21753 , \21452_21754 , \21453_21755 );
buf \U$12631 ( \21455_21757 , \21454_21756 );
xor \U$12632 ( \21456_21758 , \21450_21752 , \21455_21757 );
and \U$12633 ( \21457_21759 , \20339_20641 , \20379_20678 );
and \U$12634 ( \21458_21760 , \20339_20641 , \20386_20685 );
and \U$12635 ( \21459_21761 , \20379_20678 , \20386_20685 );
or \U$12636 ( \21460_21762 , \21457_21759 , \21458_21760 , \21459_21761 );
buf \U$12637 ( \21461_21763 , \21460_21762 );
and \U$12638 ( \21462_21764 , \20401_20700 , \20407_20706 );
and \U$12639 ( \21463_21765 , \20401_20700 , \20414_20713 );
and \U$12640 ( \21464_21766 , \20407_20706 , \20414_20713 );
or \U$12641 ( \21465_21767 , \21462_21764 , \21463_21765 , \21464_21766 );
buf \U$12642 ( \21466_21768 , \21465_21767 );
xor \U$12643 ( \21467_21769 , \21461_21763 , \21466_21768 );
and \U$12644 ( \21468_21770 , \10411_10707 , \20787_21086_nG9bdb );
and \U$12645 ( \21469_21771 , \20428_20727 , \20751_21050 );
and \U$12646 ( \21470_21772 , \20751_21050 , \20776_21075 );
and \U$12647 ( \21471_21773 , \20428_20727 , \20776_21075 );
or \U$12648 ( \21472_21774 , \21469_21771 , \21470_21772 , \21471_21773 );
and \U$12649 ( \21473_21775 , \20756_21055 , \20760_21059 );
and \U$12650 ( \21474_21776 , \20760_21059 , \20775_21074 );
and \U$12651 ( \21475_21777 , \20756_21055 , \20775_21074 );
or \U$12652 ( \21476_21778 , \21473_21775 , \21474_21776 , \21475_21777 );
and \U$12653 ( \21477_21779 , \20740_21039 , \20744_21043 );
and \U$12654 ( \21478_21780 , \20744_21043 , \20749_21048 );
and \U$12655 ( \21479_21781 , \20740_21039 , \20749_21048 );
or \U$12656 ( \21480_21782 , \21477_21779 , \21478_21780 , \21479_21781 );
and \U$12657 ( \21481_21783 , \19259_19558 , \11275_11574 );
and \U$12658 ( \21482_21784 , \20242_20544 , \10976_11278 );
nor \U$12659 ( \21483_21785 , \21481_21783 , \21482_21784 );
xnor \U$12660 ( \21484_21786 , \21483_21785 , \11281_11580 );
and \U$12661 ( \21485_21787 , \11287_11586 , \19235_19534 );
and \U$12662 ( \21486_21788 , \12146_12448 , \18743_19045 );
nor \U$12663 ( \21487_21789 , \21485_21787 , \21486_21788 );
xnor \U$12664 ( \21488_21790 , \21487_21789 , \19241_19540 );
xor \U$12665 ( \21489_21791 , \21484_21786 , \21488_21790 );
and \U$12666 ( \21490_21792 , \10686_10988 , \20706_21005 );
and \U$12667 ( \21491_21793 , \10968_11270 , \20255_20557 );
nor \U$12668 ( \21492_21794 , \21490_21792 , \21491_21793 );
xnor \U$12669 ( \21493_21795 , \21492_21794 , \20712_21011 );
xor \U$12670 ( \21494_21796 , \21489_21791 , \21493_21795 );
xor \U$12671 ( \21495_21797 , \21480_21782 , \21494_21796 );
and \U$12672 ( \21496_21798 , \20432_20731 , \20436_20735 );
and \U$12673 ( \21497_21799 , \20436_20735 , \20713_21012 );
and \U$12674 ( \21498_21800 , \20432_20731 , \20713_21012 );
or \U$12675 ( \21499_21801 , \21496_21798 , \21497_21799 , \21498_21800 );
and \U$12676 ( \21500_21802 , \20737_21036 , \20739_21038 );
xor \U$12677 ( \21501_21803 , \21499_21801 , \21500_21802 );
and \U$12678 ( \21502_21804 , \12470_12769 , \17791_18090 );
and \U$12679 ( \21503_21805 , \13377_13679 , \17353_17655 );
nor \U$12680 ( \21504_21806 , \21502_21804 , \21503_21805 );
xnor \U$12681 ( \21505_21807 , \21504_21806 , \17747_18046 );
xor \U$12682 ( \21506_21808 , \21501_21803 , \21505_21807 );
xor \U$12683 ( \21507_21809 , \21495_21797 , \21506_21808 );
xor \U$12684 ( \21508_21810 , \21476_21778 , \21507_21809 );
and \U$12685 ( \21509_21811 , \20765_21064 , \20769_21068 );
and \U$12686 ( \21510_21812 , \20769_21068 , \20774_21073 );
and \U$12687 ( \21511_21813 , \20765_21064 , \20774_21073 );
or \U$12688 ( \21512_21814 , \21509_21811 , \21510_21812 , \21511_21813 );
and \U$12689 ( \21513_21815 , \20714_21013 , \20728_21027 );
and \U$12690 ( \21514_21816 , \20728_21027 , \20750_21049 );
and \U$12691 ( \21515_21817 , \20714_21013 , \20750_21049 );
or \U$12692 ( \21516_21818 , \21513_21815 , \21514_21816 , \21515_21817 );
xor \U$12693 ( \21517_21819 , \21512_21814 , \21516_21818 );
and \U$12694 ( \21518_21820 , \20718_21017 , \20722_21021 );
and \U$12695 ( \21519_21821 , \20722_21021 , \20727_21026 );
and \U$12696 ( \21520_21822 , \20718_21017 , \20727_21026 );
or \U$12697 ( \21521_21823 , \21518_21820 , \21519_21821 , \21520_21822 );
and \U$12698 ( \21522_21824 , \20734_21033 , \10681_10983 );
and \U$12699 ( \21523_21825 , RIdec4e38_704, \9034_9333 );
and \U$12700 ( \21524_21826 , RIdec2138_672, \9036_9335 );
and \U$12701 ( \21525_21827 , RIee1fc48_4820, \9038_9337 );
and \U$12702 ( \21526_21828 , RIdebf438_640, \9040_9339 );
and \U$12703 ( \21527_21829 , RIfc49490_5856, \9042_9341 );
and \U$12704 ( \21528_21830 , RIdebc738_608, \9044_9343 );
and \U$12705 ( \21529_21831 , RIdeb9a38_576, \9046_9345 );
and \U$12706 ( \21530_21832 , RIdeb6d38_544, \9048_9347 );
and \U$12707 ( \21531_21833 , RIfc48ef0_5852, \9050_9349 );
and \U$12708 ( \21532_21834 , RIdeb1338_480, \9052_9351 );
and \U$12709 ( \21533_21835 , RIfcd9b08_7499, \9054_9353 );
and \U$12710 ( \21534_21836 , RIdeae638_448, \9056_9355 );
and \U$12711 ( \21535_21837 , RIfc8b610_6608, \9058_9357 );
and \U$12712 ( \21536_21838 , RIdea9700_416, \9060_9359 );
and \U$12713 ( \21537_21839 , RIdea2e00_384, \9062_9361 );
and \U$12714 ( \21538_21840 , RIde9c500_352, \9064_9363 );
and \U$12715 ( \21539_21841 , RIee1c9a8_4784, \9066_9365 );
and \U$12716 ( \21540_21842 , RIee1b8c8_4772, \9068_9367 );
and \U$12717 ( \21541_21843 , RIfc80918_6485, \9070_9369 );
and \U$12718 ( \21542_21844 , RIfcdad50_7512, \9072_9371 );
and \U$12719 ( \21543_21845 , RIfe86e68_7879, \9074_9373 );
and \U$12720 ( \21544_21846 , RIde8cee8_277, \9076_9375 );
and \U$12721 ( \21545_21847 , RIfe86d00_7878, \9078_9377 );
and \U$12722 ( \21546_21848 , RIfec0d20_8314, \9080_9379 );
and \U$12723 ( \21547_21849 , RIde81098_219, \9082_9381 );
and \U$12724 ( \21548_21850 , RIfc8b8e0_6610, \9084_9383 );
and \U$12725 ( \21549_21851 , RIfcd2d58_7421, \9086_9385 );
and \U$12726 ( \21550_21852 , RIfce4530_7620, \9088_9387 );
and \U$12727 ( \21551_21853 , RIfc8ba48_6611, \9090_9389 );
and \U$12728 ( \21552_21854 , RIe16b210_2596, \9092_9391 );
and \U$12729 ( \21553_21855 , RIe1698c0_2578, \9094_9393 );
and \U$12730 ( \21554_21856 , RIe1679d0_2556, \9096_9395 );
and \U$12731 ( \21555_21857 , RIe164e38_2525, \9098_9397 );
and \U$12732 ( \21556_21858 , RIe162138_2493, \9100_9399 );
and \U$12733 ( \21557_21859 , RIee370f0_5085, \9102_9401 );
and \U$12734 ( \21558_21860 , RIe15f438_2461, \9104_9403 );
and \U$12735 ( \21559_21861 , RIfc999e0_6770, \9106_9405 );
and \U$12736 ( \21560_21862 , RIe15c738_2429, \9108_9407 );
and \U$12737 ( \21561_21863 , RIe156d38_2365, \9110_9409 );
and \U$12738 ( \21562_21864 , RIe154038_2333, \9112_9411 );
and \U$12739 ( \21563_21865 , RIfc3f260_5744, \9114_9413 );
and \U$12740 ( \21564_21866 , RIe151338_2301, \9116_9415 );
and \U$12741 ( \21565_21867 , RIfc48518_5845, \9118_9417 );
and \U$12742 ( \21566_21868 , RIe14e638_2269, \9120_9419 );
and \U$12743 ( \21567_21869 , RIfc99e18_6773, \9122_9421 );
and \U$12744 ( \21568_21870 , RIe14b938_2237, \9124_9423 );
and \U$12745 ( \21569_21871 , RIe148c38_2205, \9126_9425 );
and \U$12746 ( \21570_21872 , RIe145f38_2173, \9128_9427 );
and \U$12747 ( \21571_21873 , RIee34288_5052, \9130_9429 );
and \U$12748 ( \21572_21874 , RIee33040_5039, \9132_9431 );
and \U$12749 ( \21573_21875 , RIee31f60_5027, \9134_9433 );
and \U$12750 ( \21574_21876 , RIfcd99a0_7498, \9136_9435 );
and \U$12751 ( \21575_21877 , RIfe86b98_7877, \9138_9437 );
and \U$12752 ( \21576_21878 , RIdf3e9e0_2089, \9140_9439 );
and \U$12753 ( \21577_21879 , RIfe86a30_7876, \9142_9441 );
and \U$12754 ( \21578_21880 , RIdf3a4f8_2040, \9144_9443 );
and \U$12755 ( \21579_21881 , RIfcc3470_7244, \9146_9445 );
and \U$12756 ( \21580_21882 , RIee2f530_4997, \9148_9447 );
and \U$12757 ( \21581_21883 , RIfc7fdd8_6477, \9150_9449 );
and \U$12758 ( \21582_21884 , RIee2d370_4973, \9152_9451 );
and \U$12759 ( \21583_21885 , RIdf35200_1981, \9154_9453 );
and \U$12760 ( \21584_21886 , RIfec0ff0_8316, \9156_9455 );
and \U$12761 ( \21585_21887 , RIdf30d18_1932, \9158_9457 );
and \U$12762 ( \21586_21888 , RIfec0e88_8315, \9160_9459 );
or \U$12763 ( \21587_21889 , \21523_21825 , \21524_21826 , \21525_21827 , \21526_21828 , \21527_21829 , \21528_21830 , \21529_21831 , \21530_21832 , \21531_21833 , \21532_21834 , \21533_21835 , \21534_21836 , \21535_21837 , \21536_21838 , \21537_21839 , \21538_21840 , \21539_21841 , \21540_21842 , \21541_21843 , \21542_21844 , \21543_21845 , \21544_21846 , \21545_21847 , \21546_21848 , \21547_21849 , \21548_21850 , \21549_21851 , \21550_21852 , \21551_21853 , \21552_21854 , \21553_21855 , \21554_21856 , \21555_21857 , \21556_21858 , \21557_21859 , \21558_21860 , \21559_21861 , \21560_21862 , \21561_21863 , \21562_21864 , \21563_21865 , \21564_21866 , \21565_21867 , \21566_21868 , \21567_21869 , \21568_21870 , \21569_21871 , \21570_21872 , \21571_21873 , \21572_21874 , \21573_21875 , \21574_21876 , \21575_21877 , \21576_21878 , \21577_21879 , \21578_21880 , \21579_21881 , \21580_21882 , \21581_21883 , \21582_21884 , \21583_21885 , \21584_21886 , \21585_21887 , \21586_21888 );
and \U$12764 ( \21588_21890 , RIfcd2a88_7419, \9163_9462 );
and \U$12765 ( \21589_21891 , RIfc8c858_6621, \9165_9464 );
and \U$12766 ( \21590_21892 , RIfc47ca8_5839, \9167_9466 );
and \U$12767 ( \21591_21893 , RIfcd6430_7460, \9169_9468 );
and \U$12768 ( \21592_21894 , RIdf29f68_1854, \9171_9470 );
and \U$12769 ( \21593_21895 , RIdf27da8_1830, \9173_9472 );
and \U$12770 ( \21594_21896 , RIdf26188_1810, \9175_9474 );
and \U$12771 ( \21595_21897 , RIdf24568_1790, \9177_9476 );
and \U$12772 ( \21596_21898 , RIfc8cb28_6623, \9179_9478 );
and \U$12773 ( \21597_21899 , RIfcdb188_7515, \9181_9480 );
and \U$12774 ( \21598_21900 , RIdf22948_1770, \9183_9482 );
and \U$12775 ( \21599_21901 , RIfc475a0_5834, \9185_9484 );
and \U$12776 ( \21600_21902 , RIdf21430_1755, \9187_9486 );
and \U$12777 ( \21601_21903 , RIdf1f3d8_1732, \9189_9488 );
and \U$12778 ( \21602_21904 , RIfec0bb8_8313, \9191_9490 );
and \U$12779 ( \21603_21905 , RIfe868c8_7875, \9193_9492 );
and \U$12780 ( \21604_21906 , RIdf16a08_1634, \9195_9494 );
and \U$12781 ( \21605_21907 , RIdf13d08_1602, \9197_9496 );
and \U$12782 ( \21606_21908 , RIdf11008_1570, \9199_9498 );
and \U$12783 ( \21607_21909 , RIdf0e308_1538, \9201_9500 );
and \U$12784 ( \21608_21910 , RIdf0b608_1506, \9203_9502 );
and \U$12785 ( \21609_21911 , RIdf08908_1474, \9205_9504 );
and \U$12786 ( \21610_21912 , RIdf05c08_1442, \9207_9506 );
and \U$12787 ( \21611_21913 , RIdf02f08_1410, \9209_9508 );
and \U$12788 ( \21612_21914 , RIdefd508_1346, \9211_9510 );
and \U$12789 ( \21613_21915 , RIdefa808_1314, \9213_9512 );
and \U$12790 ( \21614_21916 , RIdef7b08_1282, \9215_9514 );
and \U$12791 ( \21615_21917 , RIdef4e08_1250, \9217_9516 );
and \U$12792 ( \21616_21918 , RIdef2108_1218, \9219_9518 );
and \U$12793 ( \21617_21919 , RIdeef408_1186, \9221_9520 );
and \U$12794 ( \21618_21920 , RIdeec708_1154, \9223_9522 );
and \U$12795 ( \21619_21921 , RIdee9a08_1122, \9225_9524 );
and \U$12796 ( \21620_21922 , RIee254e0_4883, \9227_9526 );
and \U$12797 ( \21621_21923 , RIee246d0_4873, \9229_9528 );
and \U$12798 ( \21622_21924 , RIee23b90_4865, \9231_9530 );
and \U$12799 ( \21623_21925 , RIee231b8_4858, \9233_9532 );
and \U$12800 ( \21624_21926 , RIfe86fd0_7880, \9235_9534 );
and \U$12801 ( \21625_21927 , RIdee2820_1041, \9237_9536 );
and \U$12802 ( \21626_21928 , RIdee0930_1019, \9239_9538 );
and \U$12803 ( \21627_21929 , RIdede608_994, \9241_9540 );
and \U$12804 ( \21628_21930 , RIfc55da8_5999, \9243_9542 );
and \U$12805 ( \21629_21931 , RIfc98a68_6759, \9245_9544 );
and \U$12806 ( \21630_21932 , RIfcc3038_7241, \9247_9546 );
and \U$12807 ( \21631_21933 , RIfc464c0_5822, \9249_9548 );
and \U$12808 ( \21632_21934 , RIded9310_935, \9251_9550 );
and \U$12809 ( \21633_21935 , RIded6e80_909, \9253_9552 );
and \U$12810 ( \21634_21936 , RIded4f90_887, \9255_9554 );
and \U$12811 ( \21635_21937 , RIded2b00_861, \9257_9556 );
and \U$12812 ( \21636_21938 , RIded0238_832, \9259_9558 );
and \U$12813 ( \21637_21939 , RIdecd538_800, \9261_9560 );
and \U$12814 ( \21638_21940 , RIdeca838_768, \9263_9562 );
and \U$12815 ( \21639_21941 , RIdec7b38_736, \9265_9564 );
and \U$12816 ( \21640_21942 , RIdeb4038_512, \9267_9566 );
and \U$12817 ( \21641_21943 , RIde95c00_320, \9269_9568 );
and \U$12818 ( \21642_21944 , RIe16dc40_2626, \9271_9570 );
and \U$12819 ( \21643_21945 , RIe159a38_2397, \9273_9572 );
and \U$12820 ( \21644_21946 , RIe143238_2141, \9275_9574 );
and \U$12821 ( \21645_21947 , RIdf37c30_2011, \9277_9576 );
and \U$12822 ( \21646_21948 , RIdf2c290_1879, \9279_9578 );
and \U$12823 ( \21647_21949 , RIdf1cb10_1703, \9281_9580 );
and \U$12824 ( \21648_21950 , RIdf00208_1378, \9283_9582 );
and \U$12825 ( \21649_21951 , RIdee6d08_1090, \9285_9584 );
and \U$12826 ( \21650_21952 , RIdedba70_963, \9287_9586 );
and \U$12827 ( \21651_21953 , RIde7bb48_193, \9289_9588 );
or \U$12828 ( \21652_21954 , \21588_21890 , \21589_21891 , \21590_21892 , \21591_21893 , \21592_21894 , \21593_21895 , \21594_21896 , \21595_21897 , \21596_21898 , \21597_21899 , \21598_21900 , \21599_21901 , \21600_21902 , \21601_21903 , \21602_21904 , \21603_21905 , \21604_21906 , \21605_21907 , \21606_21908 , \21607_21909 , \21608_21910 , \21609_21911 , \21610_21912 , \21611_21913 , \21612_21914 , \21613_21915 , \21614_21916 , \21615_21917 , \21616_21918 , \21617_21919 , \21618_21920 , \21619_21921 , \21620_21922 , \21621_21923 , \21622_21924 , \21623_21925 , \21624_21926 , \21625_21927 , \21626_21928 , \21627_21929 , \21628_21930 , \21629_21931 , \21630_21932 , \21631_21933 , \21632_21934 , \21633_21935 , \21634_21936 , \21635_21937 , \21636_21938 , \21637_21939 , \21638_21940 , \21639_21941 , \21640_21942 , \21641_21943 , \21642_21944 , \21643_21945 , \21644_21946 , \21645_21947 , \21646_21948 , \21647_21949 , \21648_21950 , \21649_21951 , \21650_21952 , \21651_21953 );
or \U$12829 ( \21653_21955 , \21587_21889 , \21652_21954 );
_DC \g65ad/U$1 ( \21654 , \21653_21955 , \9298_9597 );
and \U$12830 ( \21655_21957 , RIe19d0d0_3164, \8760_9059 );
and \U$12831 ( \21656_21958 , RIe19a3d0_3132, \8762_9061 );
and \U$12832 ( \21657_21959 , RIf1454f0_5248, \8764_9063 );
and \U$12833 ( \21658_21960 , RIe1976d0_3100, \8766_9065 );
and \U$12834 ( \21659_21961 , RIf144578_5237, \8768_9067 );
and \U$12835 ( \21660_21962 , RIe1949d0_3068, \8770_9069 );
and \U$12836 ( \21661_21963 , RIe191cd0_3036, \8772_9071 );
and \U$12837 ( \21662_21964 , RIe18efd0_3004, \8774_9073 );
and \U$12838 ( \21663_21965 , RIe1895d0_2940, \8776_9075 );
and \U$12839 ( \21664_21966 , RIe1868d0_2908, \8778_9077 );
and \U$12840 ( \21665_21967 , RIf143498_5225, \8780_9079 );
and \U$12841 ( \21666_21968 , RIe183bd0_2876, \8782_9081 );
and \U$12842 ( \21667_21969 , RIfc51758_5949, \8784_9083 );
and \U$12843 ( \21668_21970 , RIe180ed0_2844, \8786_9085 );
and \U$12844 ( \21669_21971 , RIe17e1d0_2812, \8788_9087 );
and \U$12845 ( \21670_21972 , RIe17b4d0_2780, \8790_9089 );
and \U$12846 ( \21671_21973 , RIfc9b060_6786, \8792_9091 );
and \U$12847 ( \21672_21974 , RIfc9ee40_6830, \8794_9093 );
and \U$12848 ( \21673_21975 , RIe176e80_2730, \8796_9095 );
and \U$12849 ( \21674_21976 , RIe175800_2714, \8798_9097 );
and \U$12850 ( \21675_21977 , RIfcb70f8_7105, \8800_9099 );
and \U$12851 ( \21676_21978 , RIfce0cf0_7580, \8802_9101 );
and \U$12852 ( \21677_21979 , RIfcc4280_7254, \8804_9103 );
and \U$12853 ( \21678_21980 , RIfcba7d0_7144, \8806_9105 );
and \U$12854 ( \21679_21981 , RIee3bfb0_5141, \8808_9107 );
and \U$12855 ( \21680_21982 , RIee3aed0_5129, \8810_9109 );
and \U$12856 ( \21681_21983 , RIee39b20_5115, \8812_9111 );
and \U$12857 ( \21682_21984 , RIe173370_2688, \8814_9113 );
and \U$12858 ( \21683_21985 , RIf170060_5734, \8816_9115 );
and \U$12859 ( \21684_21986 , RIf16f3b8_5725, \8818_9117 );
and \U$12860 ( \21685_21987 , RIf16dea0_5710, \8820_9119 );
and \U$12861 ( \21686_21988 , RIf16d4c8_5703, \8822_9121 );
and \U$12862 ( \21687_21989 , RIf16c988_5695, \8824_9123 );
and \U$12863 ( \21688_21990 , RIe223428_4691, \8826_9125 );
and \U$12864 ( \21689_21991 , RIf16bb78_5685, \8828_9127 );
and \U$12865 ( \21690_21992 , RIe220728_4659, \8830_9129 );
and \U$12866 ( \21691_21993 , RIf16aa98_5673, \8832_9131 );
and \U$12867 ( \21692_21994 , RIe21da28_4627, \8834_9133 );
and \U$12868 ( \21693_21995 , RIe218028_4563, \8836_9135 );
and \U$12869 ( \21694_21996 , RIe215328_4531, \8838_9137 );
and \U$12870 ( \21695_21997 , RIf16a0c0_5666, \8840_9139 );
and \U$12871 ( \21696_21998 , RIe212628_4499, \8842_9141 );
and \U$12872 ( \21697_21999 , RIf168e78_5653, \8844_9143 );
and \U$12873 ( \21698_22000 , RIe20f928_4467, \8846_9145 );
and \U$12874 ( \21699_22001 , RIf167c30_5640, \8848_9147 );
and \U$12875 ( \21700_22002 , RIe20cc28_4435, \8850_9149 );
and \U$12876 ( \21701_22003 , RIe209f28_4403, \8852_9151 );
and \U$12877 ( \21702_22004 , RIe207228_4371, \8854_9153 );
and \U$12878 ( \21703_22005 , RIf166f88_5631, \8856_9155 );
and \U$12879 ( \21704_22006 , RIf165d40_5618, \8858_9157 );
and \U$12880 ( \21705_22007 , RIfec0618_8309, \8860_9159 );
and \U$12881 ( \21706_22008 , RIfe86760_7874, \8862_9161 );
and \U$12882 ( \21707_22009 , RIfc52b08_5963, \8864_9163 );
and \U$12883 ( \21708_22010 , RIf164288_5599, \8866_9165 );
and \U$12884 ( \21709_22011 , RIf163310_5588, \8868_9167 );
and \U$12885 ( \21710_22012 , RIf161c90_5572, \8870_9169 );
and \U$12886 ( \21711_22013 , RIf15fda0_5550, \8872_9171 );
and \U$12887 ( \21712_22014 , RIf15deb0_5528, \8874_9173 );
and \U$12888 ( \21713_22015 , RIfe865f8_7873, \8876_9175 );
and \U$12889 ( \21714_22016 , RIfe85d88_7867, \8878_9177 );
and \U$12890 ( \21715_22017 , RIf15c998_5513, \8880_9179 );
and \U$12891 ( \21716_22018 , RIf15b480_5498, \8882_9181 );
and \U$12892 ( \21717_22019 , RIf15a3a0_5486, \8884_9183 );
and \U$12893 ( \21718_22020 , RIf159b30_5480, \8886_9185 );
or \U$12894 ( \21719_22021 , \21655_21957 , \21656_21958 , \21657_21959 , \21658_21960 , \21659_21961 , \21660_21962 , \21661_21963 , \21662_21964 , \21663_21965 , \21664_21966 , \21665_21967 , \21666_21968 , \21667_21969 , \21668_21970 , \21669_21971 , \21670_21972 , \21671_21973 , \21672_21974 , \21673_21975 , \21674_21976 , \21675_21977 , \21676_21978 , \21677_21979 , \21678_21980 , \21679_21981 , \21680_21982 , \21681_21983 , \21682_21984 , \21683_21985 , \21684_21986 , \21685_21987 , \21686_21988 , \21687_21989 , \21688_21990 , \21689_21991 , \21690_21992 , \21691_21993 , \21692_21994 , \21693_21995 , \21694_21996 , \21695_21997 , \21696_21998 , \21697_21999 , \21698_22000 , \21699_22001 , \21700_22002 , \21701_22003 , \21702_22004 , \21703_22005 , \21704_22006 , \21705_22007 , \21706_22008 , \21707_22009 , \21708_22010 , \21709_22011 , \21710_22012 , \21711_22013 , \21712_22014 , \21713_22015 , \21714_22016 , \21715_22017 , \21716_22018 , \21717_22019 , \21718_22020 );
and \U$12895 ( \21720_22022 , RIfc83348_6515, \8889_9188 );
and \U$12896 ( \21721_22023 , RIfc4ade0_5874, \8891_9190 );
and \U$12897 ( \21722_22024 , RIfc89720_6586, \8893_9192 );
and \U$12898 ( \21723_22025 , RIe1f9f38_4221, \8895_9194 );
and \U$12899 ( \21724_22026 , RIfc4ac78_5873, \8897_9196 );
and \U$12900 ( \21725_22027 , RIfc9f110_6832, \8899_9198 );
and \U$12901 ( \21726_22028 , RIfc4ab10_5872, \8901_9200 );
and \U$12902 ( \21727_22029 , RIe1f5078_4165, \8903_9202 );
and \U$12903 ( \21728_22030 , RIf152ee8_5403, \8905_9204 );
and \U$12904 ( \21729_22031 , RIfc899f0_6588, \8907_9206 );
and \U$12905 ( \21730_22032 , RIf150620_5374, \8909_9208 );
and \U$12906 ( \21731_22033 , RIe1f2eb8_4141, \8911_9210 );
and \U$12907 ( \21732_22034 , RIf14f6a8_5363, \8913_9212 );
and \U$12908 ( \21733_22035 , RIf14ea00_5354, \8915_9214 );
and \U$12909 ( \21734_22036 , RIf14dbf0_5344, \8917_9216 );
and \U$12910 ( \21735_22037 , RIe1edbc0_4082, \8919_9218 );
and \U$12911 ( \21736_22038 , RIe1eb190_4052, \8921_9220 );
and \U$12912 ( \21737_22039 , RIe1e8490_4020, \8923_9222 );
and \U$12913 ( \21738_22040 , RIe1e5790_3988, \8925_9224 );
and \U$12914 ( \21739_22041 , RIe1e2a90_3956, \8927_9226 );
and \U$12915 ( \21740_22042 , RIe1dfd90_3924, \8929_9228 );
and \U$12916 ( \21741_22043 , RIe1dd090_3892, \8931_9230 );
and \U$12917 ( \21742_22044 , RIe1da390_3860, \8933_9232 );
and \U$12918 ( \21743_22045 , RIe1d7690_3828, \8935_9234 );
and \U$12919 ( \21744_22046 , RIe1d1c90_3764, \8937_9236 );
and \U$12920 ( \21745_22047 , RIe1cef90_3732, \8939_9238 );
and \U$12921 ( \21746_22048 , RIe1cc290_3700, \8941_9240 );
and \U$12922 ( \21747_22049 , RIe1c9590_3668, \8943_9242 );
and \U$12923 ( \21748_22050 , RIe1c6890_3636, \8945_9244 );
and \U$12924 ( \21749_22051 , RIe1c3b90_3604, \8947_9246 );
and \U$12925 ( \21750_22052 , RIe1c0e90_3572, \8949_9248 );
and \U$12926 ( \21751_22053 , RIe1be190_3540, \8951_9250 );
and \U$12927 ( \21752_22054 , RIf14c6d8_5329, \8953_9252 );
and \U$12928 ( \21753_22055 , RIf14b490_5316, \8955_9254 );
and \U$12929 ( \21754_22056 , RIfe85ef0_7868, \8957_9256 );
and \U$12930 ( \21755_22057 , RIfe86490_7872, \8959_9258 );
and \U$12931 ( \21756_22058 , RIf14a248_5303, \8961_9260 );
and \U$12932 ( \21757_22059 , RIfc819f8_6497, \8963_9262 );
and \U$12933 ( \21758_22060 , RIfec0a50_8312, \8965_9264 );
and \U$12934 ( \21759_22061 , RIfe861c0_7870, \8967_9266 );
and \U$12935 ( \21760_22062 , RIf148bc8_5287, \8969_9268 );
and \U$12936 ( \21761_22063 , RIf147980_5274, \8971_9270 );
and \U$12937 ( \21762_22064 , RIfe86328_7871, \8973_9272 );
and \U$12938 ( \21763_22065 , RIfec0780_8310, \8975_9274 );
and \U$12939 ( \21764_22066 , RIfcbb478_7153, \8977_9276 );
and \U$12940 ( \21765_22067 , RIf146198_5257, \8979_9278 );
and \U$12941 ( \21766_22068 , RIfe86058_7869, \8981_9280 );
and \U$12942 ( \21767_22069 , RIfec08e8_8311, \8983_9282 );
and \U$12943 ( \21768_22070 , RIe1a84d0_3292, \8985_9284 );
and \U$12944 ( \21769_22071 , RIe1a57d0_3260, \8987_9286 );
and \U$12945 ( \21770_22072 , RIe1a2ad0_3228, \8989_9288 );
and \U$12946 ( \21771_22073 , RIe19fdd0_3196, \8991_9290 );
and \U$12947 ( \21772_22074 , RIe18c2d0_2972, \8993_9292 );
and \U$12948 ( \21773_22075 , RIe1787d0_2748, \8995_9294 );
and \U$12949 ( \21774_22076 , RIe226128_4723, \8997_9296 );
and \U$12950 ( \21775_22077 , RIe21ad28_4595, \8999_9298 );
and \U$12951 ( \21776_22078 , RIe204528_4339, \9001_9300 );
and \U$12952 ( \21777_22079 , RIe1fe588_4271, \9003_9302 );
and \U$12953 ( \21778_22080 , RIe1f7940_4194, \9005_9304 );
and \U$12954 ( \21779_22081 , RIe1f0488_4111, \9007_9306 );
and \U$12955 ( \21780_22082 , RIe1d4990_3796, \9009_9308 );
and \U$12956 ( \21781_22083 , RIe1bb490_3508, \9011_9310 );
and \U$12957 ( \21782_22084 , RIe1ae308_3359, \9013_9312 );
and \U$12958 ( \21783_22085 , RIe170940_2658, \9015_9314 );
or \U$12959 ( \21784_22086 , \21720_22022 , \21721_22023 , \21722_22024 , \21723_22025 , \21724_22026 , \21725_22027 , \21726_22028 , \21727_22029 , \21728_22030 , \21729_22031 , \21730_22032 , \21731_22033 , \21732_22034 , \21733_22035 , \21734_22036 , \21735_22037 , \21736_22038 , \21737_22039 , \21738_22040 , \21739_22041 , \21740_22042 , \21741_22043 , \21742_22044 , \21743_22045 , \21744_22046 , \21745_22047 , \21746_22048 , \21747_22049 , \21748_22050 , \21749_22051 , \21750_22052 , \21751_22053 , \21752_22054 , \21753_22055 , \21754_22056 , \21755_22057 , \21756_22058 , \21757_22059 , \21758_22060 , \21759_22061 , \21760_22062 , \21761_22063 , \21762_22064 , \21763_22065 , \21764_22066 , \21765_22067 , \21766_22068 , \21767_22069 , \21768_22070 , \21769_22071 , \21770_22072 , \21771_22073 , \21772_22074 , \21773_22075 , \21774_22076 , \21775_22077 , \21776_22078 , \21777_22079 , \21778_22080 , \21779_22081 , \21780_22082 , \21781_22083 , \21782_22084 , \21783_22085 );
or \U$12960 ( \21785_22087 , \21719_22021 , \21784_22086 );
_DC \g65ae/U$1 ( \21786 , \21785_22087 , \9024_9323 );
and g65af_GF_PartitionCandidate( \21787_22089_nG65af , \21654 , \21786 );
buf \U$12961 ( \21788_22090 , \21787_22089_nG65af );
and \U$12962 ( \21789_22091 , \21788_22090 , \10389_10691 );
nor \U$12963 ( \21790_22092 , \21522_21824 , \21789_22091 );
xnor \U$12964 ( \21791_22093 , \21790_22092 , \10678_10980 );
and \U$12965 ( \21792_22094 , \16353_16655 , \13755_14054 );
and \U$12966 ( \21793_22095 , \17325_17627 , \13390_13692 );
nor \U$12967 ( \21794_22096 , \21792_22094 , \21793_22095 );
xnor \U$12968 ( \21795_22097 , \21794_22096 , \13736_14035 );
xor \U$12969 ( \21796_22098 , \21791_22093 , \21795_22097 );
_DC \g577c/U$1 ( \21797 , \21653_21955 , \9298_9597 );
_DC \g5800/U$1 ( \21798 , \21785_22087 , \9024_9323 );
xor g5801_GF_PartitionCandidate( \21799_22101_nG5801 , \21797 , \21798 );
buf \U$12970 ( \21800_22102 , \21799_22101_nG5801 );
xor \U$12971 ( \21801_22103 , \21800_22102 , \20703_21002 );
and \U$12972 ( \21802_22104 , \10385_10687 , \21801_22103 );
xor \U$12973 ( \21803_22105 , \21796_22098 , \21802_22104 );
xor \U$12974 ( \21804_22106 , \21521_21823 , \21803_22105 );
and \U$12975 ( \21805_22107 , \17736_18035 , \12491_12790 );
and \U$12976 ( \21806_22108 , \18730_19032 , \12159_12461 );
nor \U$12977 ( \21807_22109 , \21805_22107 , \21806_22108 );
xnor \U$12978 ( \21808_22110 , \21807_22109 , \12481_12780 );
and \U$12979 ( \21809_22111 , \15022_15321 , \15037_15336 );
and \U$12980 ( \21810_22112 , \15965_16267 , \14661_14963 );
nor \U$12981 ( \21811_22113 , \21809_22111 , \21810_22112 );
xnor \U$12982 ( \21812_22114 , \21811_22113 , \15043_15342 );
xor \U$12983 ( \21813_22115 , \21808_22110 , \21812_22114 );
and \U$12984 ( \21814_22116 , \13725_14024 , \16333_16635 );
and \U$12985 ( \21815_22117 , \14648_14950 , \15999_16301 );
nor \U$12986 ( \21816_22118 , \21814_22116 , \21815_22117 );
xnor \U$12987 ( \21817_22119 , \21816_22118 , \16323_16625 );
xor \U$12988 ( \21818_22120 , \21813_22115 , \21817_22119 );
xor \U$12989 ( \21819_22121 , \21804_22106 , \21818_22120 );
xor \U$12990 ( \21820_22122 , \21517_21819 , \21819_22121 );
xor \U$12991 ( \21821_22123 , \21508_21810 , \21820_22122 );
xor \U$12992 ( \21822_22124 , \21472_21774 , \21821_22123 );
and \U$12993 ( \21823_22125 , \20777_21076 , \20781_21080 );
and \U$12994 ( \21824_22126 , \20782_21081 , \20785_21084 );
or \U$12995 ( \21825_22127 , \21823_22125 , \21824_22126 );
xor \U$12996 ( \21826_22128 , \21822_22124 , \21825_22127 );
buf g9bd8_GF_PartitionCandidate( \21827_22129_nG9bd8 , \21826_22128 );
and \U$12997 ( \21828_22130 , \10402_10704 , \21827_22129_nG9bd8 );
or \U$12998 ( \21829_22131 , \21468_21770 , \21828_22130 );
xor \U$12999 ( \21830_22132 , \10399_10703 , \21829_22131 );
buf \U$13000 ( \21831_22133 , \21830_22132 );
buf \U$13002 ( \21832_22134 , \21831_22133 );
xor \U$13003 ( \21833_22135 , \21467_21769 , \21832_22134 );
buf \U$13004 ( \21834_22136 , \21833_22135 );
xor \U$13005 ( \21835_22137 , \21456_21758 , \21834_22136 );
and \U$13006 ( \21836_22138 , \21363_21665 , \21835_22137 );
and \U$13007 ( \21837_22139 , \21367_21669 , \21835_22137 );
or \U$13008 ( \21838_22140 , \21368_21670 , \21836_22138 , \21837_22139 );
and \U$13009 ( \21839_22141 , \20802_21101 , \20806_21105 );
and \U$13010 ( \21840_22142 , \20802_21101 , \21362_21664 );
and \U$13011 ( \21841_22143 , \20806_21105 , \21362_21664 );
or \U$13012 ( \21842_22144 , \21839_22141 , \21840_22142 , \21841_22143 );
xor \U$13013 ( \21843_22145 , \21838_22140 , \21842_22144 );
and \U$13014 ( \21844_22146 , \21450_21752 , \21455_21757 );
and \U$13015 ( \21845_22147 , \21450_21752 , \21834_22136 );
and \U$13016 ( \21846_22148 , \21455_21757 , \21834_22136 );
or \U$13017 ( \21847_22149 , \21844_22146 , \21845_22147 , \21846_22148 );
xor \U$13018 ( \21848_22150 , \21843_22145 , \21847_22149 );
and \U$13019 ( \21849_22151 , \21461_21763 , \21466_21768 );
and \U$13020 ( \21850_22152 , \21461_21763 , \21832_22134 );
and \U$13021 ( \21851_22153 , \21466_21768 , \21832_22134 );
or \U$13022 ( \21852_22154 , \21849_22151 , \21850_22152 , \21851_22153 );
buf \U$13023 ( \21853_22155 , \21852_22154 );
and \U$13024 ( \21854_22156 , \21422_21724 , \21424_21726 );
and \U$13025 ( \21855_22157 , \21422_21724 , \21431_21733 );
and \U$13026 ( \21856_22158 , \21424_21726 , \21431_21733 );
or \U$13027 ( \21857_22159 , \21854_22156 , \21855_22157 , \21856_22158 );
buf \U$13028 ( \21858_22160 , \21857_22159 );
and \U$13029 ( \21859_22161 , \16405_15940 , \14682_14984_nG9bf6 );
and \U$13030 ( \21860_22162 , \15638_15937 , \15074_15373_nG9bf3 );
or \U$13031 ( \21861_22163 , \21859_22161 , \21860_22162 );
xor \U$13032 ( \21862_22164 , \15637_15936 , \21861_22163 );
buf \U$13033 ( \21863_22165 , \21862_22164 );
buf \U$13035 ( \21864_22166 , \21863_22165 );
xor \U$13036 ( \21865_22167 , \21858_22160 , \21864_22166 );
and \U$13037 ( \21866_22168 , \14710_14631 , \16013_16315_nG9bf0 );
and \U$13038 ( \21867_22169 , \14329_14628 , \16378_16680_nG9bed );
or \U$13039 ( \21868_22170 , \21866_22168 , \21867_22169 );
xor \U$13040 ( \21869_22171 , \14328_14627 , \21868_22170 );
buf \U$13041 ( \21870_22172 , \21869_22171 );
buf \U$13043 ( \21871_22173 , \21870_22172 );
xor \U$13044 ( \21872_22174 , \21865_22167 , \21871_22173 );
buf \U$13045 ( \21873_22175 , \21872_22174 );
and \U$13046 ( \21874_22176 , \12183_12157 , \18789_19091_nG9be4 );
and \U$13047 ( \21875_22177 , \11855_12154 , \19287_19586_nG9be1 );
or \U$13048 ( \21876_22178 , \21874_22176 , \21875_22177 );
xor \U$13049 ( \21877_22179 , \11854_12153 , \21876_22178 );
buf \U$13050 ( \21878_22180 , \21877_22179 );
buf \U$13052 ( \21879_22181 , \21878_22180 );
xor \U$13053 ( \21880_22182 , \21873_22175 , \21879_22181 );
and \U$13054 ( \21881_22183 , \10996_10421 , \20306_20608_nG9bde );
and \U$13055 ( \21882_22184 , \10119_10418 , \20787_21086_nG9bdb );
or \U$13056 ( \21883_22185 , \21881_22183 , \21882_22184 );
xor \U$13057 ( \21884_22186 , \10118_10417 , \21883_22185 );
buf \U$13058 ( \21885_22187 , \21884_22186 );
buf \U$13060 ( \21886_22188 , \21885_22187 );
xor \U$13061 ( \21887_22189 , \21880_22182 , \21886_22188 );
buf \U$13062 ( \21888_22190 , \21887_22189 );
xor \U$13063 ( \21889_22191 , \21853_22155 , \21888_22190 );
and \U$13064 ( \21890_22192 , \21378_21680 , \21384_21686 );
and \U$13065 ( \21891_22193 , \21378_21680 , \21391_21693 );
and \U$13066 ( \21892_22194 , \21384_21686 , \21391_21693 );
or \U$13067 ( \21893_22195 , \21890_22192 , \21891_22193 , \21892_22194 );
buf \U$13068 ( \21894_22196 , \21893_22195 );
and \U$13069 ( \21895_22197 , \21355_21654 , \21359_21661 );
buf \U$13070 ( \21896_22198 , \21895_22197 );
buf \U$13072 ( \21897_22199 , \21896_22198 );
and \U$13073 ( \21898_22200 , \20353_20155 , \10981_11283_nG9c08 );
and \U$13074 ( \21899_22201 , \19853_20152 , \11299_11598_nG9c05 );
or \U$13075 ( \21900_22202 , \21898_22200 , \21899_22201 );
xor \U$13076 ( \21901_22203 , \19852_20151 , \21900_22202 );
buf \U$13077 ( \21902_22204 , \21901_22203 );
buf \U$13079 ( \21903_22205 , \21902_22204 );
xor \U$13080 ( \21904_22206 , \21897_22199 , \21903_22205 );
buf \U$13081 ( \21905_22207 , \21904_22206 );
not \U$12521 ( \21906_21656 , \21356_21655 );
xor \U$12522 ( \21907_21657 , \21350_21649_nG441e , \21353_21652_nG4421 );
and \U$12523 ( \21908_21658 , \21906_21656 , \21907_21657 );
and \U$13082 ( \21909_22208 , \21908_21658 , \10392_10694_nG9c0e );
and \U$13083 ( \21910_22209 , \21356_21655 , \10693_10995_nG9c0b );
or \U$13084 ( \21911_22210 , \21909_22208 , \21910_22209 );
xor \U$13085 ( \21912_22211 , \21355_21654 , \21911_22210 );
buf \U$13086 ( \21913_22212 , \21912_22211 );
buf \U$13088 ( \21914_22213 , \21913_22212 );
xor \U$13089 ( \21915_22214 , \21905_22207 , \21914_22213 );
and \U$13090 ( \21916_22215 , \18908_18702 , \12168_12470_nG9c02 );
and \U$13091 ( \21917_22216 , \18400_18699 , \12502_12801_nG9bff );
or \U$13092 ( \21918_22217 , \21916_22215 , \21917_22216 );
xor \U$13093 ( \21919_22218 , \18399_18698 , \21918_22217 );
buf \U$13094 ( \21920_22219 , \21919_22218 );
buf \U$13096 ( \21921_22220 , \21920_22219 );
xor \U$13097 ( \21922_22221 , \21915_22214 , \21921_22220 );
buf \U$13098 ( \21923_22222 , \21922_22221 );
and \U$13099 ( \21924_22223 , \21414_21716 , \21420_21722 );
buf \U$13100 ( \21925_22224 , \21924_22223 );
xor \U$13101 ( \21926_22225 , \21923_22222 , \21925_22224 );
and \U$13102 ( \21927_22226 , \17437_17297 , \13403_13705_nG9bfc );
and \U$13103 ( \21928_22227 , \16995_17294 , \13771_14070_nG9bf9 );
or \U$13104 ( \21929_22228 , \21927_22226 , \21928_22227 );
xor \U$13105 ( \21930_22229 , \16994_17293 , \21929_22228 );
buf \U$13106 ( \21931_22230 , \21930_22229 );
buf \U$13108 ( \21932_22231 , \21931_22230 );
xor \U$13109 ( \21933_22232 , \21926_22225 , \21932_22231 );
buf \U$13110 ( \21934_22233 , \21933_22232 );
xor \U$13111 ( \21935_22234 , \21894_22196 , \21934_22233 );
and \U$13112 ( \21936_22235 , \13431_13370 , \17363_17665_nG9bea );
and \U$13113 ( \21937_22236 , \13068_13367 , \17808_18107_nG9be7 );
or \U$13114 ( \21938_22237 , \21936_22235 , \21937_22236 );
xor \U$13115 ( \21939_22238 , \13067_13366 , \21938_22237 );
buf \U$13116 ( \21940_22239 , \21939_22238 );
buf \U$13118 ( \21941_22240 , \21940_22239 );
xor \U$13119 ( \21942_22241 , \21935_22234 , \21941_22240 );
buf \U$13120 ( \21943_22242 , \21942_22241 );
xor \U$13121 ( \21944_22243 , \21889_22191 , \21943_22242 );
buf \U$13122 ( \21945_22244 , \21944_22243 );
and \U$13123 ( \21946_22245 , \21393_21695 , \21398_21700 );
and \U$13124 ( \21947_22246 , \21393_21695 , \21405_21707 );
and \U$13125 ( \21948_22247 , \21398_21700 , \21405_21707 );
or \U$13126 ( \21949_22248 , \21946_22245 , \21947_22246 , \21948_22247 );
buf \U$13127 ( \21950_22249 , \21949_22248 );
and \U$13128 ( \21951_22250 , \21433_21735 , \21439_21741 );
and \U$13129 ( \21952_22251 , \21433_21735 , \21446_21748 );
and \U$13130 ( \21953_22252 , \21439_21741 , \21446_21748 );
or \U$13131 ( \21954_22253 , \21951_22250 , \21952_22251 , \21953_22252 );
buf \U$13132 ( \21955_22254 , \21954_22253 );
xor \U$13133 ( \21956_22255 , \21950_22249 , \21955_22254 );
and \U$13134 ( \21957_22256 , \10411_10707 , \21827_22129_nG9bd8 );
and \U$13135 ( \21958_22257 , \21512_21814 , \21516_21818 );
and \U$13136 ( \21959_22258 , \21516_21818 , \21819_22121 );
and \U$13137 ( \21960_22259 , \21512_21814 , \21819_22121 );
or \U$13138 ( \21961_22260 , \21958_22257 , \21959_22258 , \21960_22259 );
and \U$13139 ( \21962_22261 , \21499_21801 , \21500_21802 );
and \U$13140 ( \21963_22262 , \21500_21802 , \21505_21807 );
and \U$13141 ( \21964_22263 , \21499_21801 , \21505_21807 );
or \U$13142 ( \21965_22264 , \21962_22261 , \21963_22262 , \21964_22263 );
and \U$13143 ( \21966_22265 , \20242_20544 , \11275_11574 );
and \U$13144 ( \21967_22266 , \20734_21033 , \10976_11278 );
nor \U$13145 ( \21968_22267 , \21966_22265 , \21967_22266 );
xnor \U$13146 ( \21969_22268 , \21968_22267 , \11281_11580 );
and \U$13147 ( \21970_22269 , \15965_16267 , \15037_15336 );
and \U$13148 ( \21971_22270 , \16353_16655 , \14661_14963 );
nor \U$13149 ( \21972_22271 , \21970_22269 , \21971_22270 );
xnor \U$13150 ( \21973_22272 , \21972_22271 , \15043_15342 );
xor \U$13151 ( \21974_22273 , \21969_22268 , \21973_22272 );
and \U$13152 ( \21975_22274 , RIdec4fa0_705, \9034_9333 );
and \U$13153 ( \21976_22275 , RIdec22a0_673, \9036_9335 );
and \U$13154 ( \21977_22276 , RIee1fdb0_4821, \9038_9337 );
and \U$13155 ( \21978_22277 , RIdebf5a0_641, \9040_9339 );
and \U$13156 ( \21979_22278 , RIee1f270_4813, \9042_9341 );
and \U$13157 ( \21980_22279 , RIdebc8a0_609, \9044_9343 );
and \U$13158 ( \21981_22280 , RIdeb9ba0_577, \9046_9345 );
and \U$13159 ( \21982_22281 , RIdeb6ea0_545, \9048_9347 );
and \U$13160 ( \21983_22282 , RIee1ecd0_4809, \9050_9349 );
and \U$13161 ( \21984_22283 , RIdeb14a0_481, \9052_9351 );
and \U$13162 ( \21985_22284 , RIee1e730_4805, \9054_9353 );
and \U$13163 ( \21986_22285 , RIdeae7a0_449, \9056_9355 );
and \U$13164 ( \21987_22286 , RIee1d920_4795, \9058_9357 );
and \U$13165 ( \21988_22287 , RIdea9a48_417, \9060_9359 );
and \U$13166 ( \21989_22288 , RIdea3148_385, \9062_9361 );
and \U$13167 ( \21990_22289 , RIde9c848_353, \9064_9363 );
and \U$13168 ( \21991_22290 , RIee1cb10_4785, \9066_9365 );
and \U$13169 ( \21992_22291 , RIee1ba30_4773, \9068_9367 );
and \U$13170 ( \21993_22292 , RIee1b1c0_4767, \9070_9369 );
and \U$13171 ( \21994_22293 , RIfec04b0_8308, \9072_9371 );
and \U$13172 ( \21995_22294 , RIfe850e0_7858, \9074_9373 );
and \U$13173 ( \21996_22295 , RIde8d230_278, \9076_9375 );
and \U$13174 ( \21997_22296 , RIfea9cb0_8248, \9078_9377 );
and \U$13175 ( \21998_22297 , RIfe84f78_7857, \9080_9379 );
and \U$13176 ( \21999_22298 , RIee1a3b0_4757, \9082_9381 );
and \U$13177 ( \22000_22299 , RIfe853b0_7860, \9084_9383 );
and \U$13178 ( \22001_22300 , RIee199d8_4750, \9086_9385 );
and \U$13179 ( \22002_22301 , RIfe85248_7859, \9088_9387 );
and \U$13180 ( \22003_22302 , RIee39148_5108, \9090_9389 );
and \U$13181 ( \22004_22303 , RIe16b378_2597, \9092_9391 );
and \U$13182 ( \22005_22304 , RIee38608_5100, \9094_9393 );
and \U$13183 ( \22006_22305 , RIe167b38_2557, \9096_9395 );
and \U$13184 ( \22007_22306 , RIe164fa0_2526, \9098_9397 );
and \U$13185 ( \22008_22307 , RIe1622a0_2494, \9100_9399 );
and \U$13186 ( \22009_22308 , RIfe85950_7864, \9102_9401 );
and \U$13187 ( \22010_22309 , RIe15f5a0_2462, \9104_9403 );
and \U$13188 ( \22011_22310 , RIee36010_5073, \9106_9405 );
and \U$13189 ( \22012_22311 , RIe15c8a0_2430, \9108_9407 );
and \U$13190 ( \22013_22312 , RIe156ea0_2366, \9110_9409 );
and \U$13191 ( \22014_22313 , RIe1541a0_2334, \9112_9411 );
and \U$13192 ( \22015_22314 , RIfe85c20_7866, \9114_9413 );
and \U$13193 ( \22016_22315 , RIe1514a0_2302, \9116_9415 );
and \U$13194 ( \22017_22316 , RIee34dc8_5060, \9118_9417 );
and \U$13195 ( \22018_22317 , RIe14e7a0_2270, \9120_9419 );
and \U$13196 ( \22019_22318 , RIfc861b0_6548, \9122_9421 );
and \U$13197 ( \22020_22319 , RIe14baa0_2238, \9124_9423 );
and \U$13198 ( \22021_22320 , RIe148da0_2206, \9126_9425 );
and \U$13199 ( \22022_22321 , RIe1460a0_2174, \9128_9427 );
and \U$13200 ( \22023_22322 , RIee343f0_5053, \9130_9429 );
and \U$13201 ( \22024_22323 , RIfe85518_7861, \9132_9431 );
and \U$13202 ( \22025_22324 , RIfe857e8_7863, \9134_9433 );
and \U$13203 ( \22026_22325 , RIfe85680_7862, \9136_9435 );
and \U$13204 ( \22027_22326 , RIe140c40_2114, \9138_9437 );
and \U$13205 ( \22028_22327 , RIdf3eb48_2090, \9140_9439 );
and \U$13206 ( \22029_22328 , RIdf3c820_2065, \9142_9441 );
and \U$13207 ( \22030_22329 , RIdf3a660_2041, \9144_9443 );
and \U$13208 ( \22031_22330 , RIfc9d4f0_6812, \9146_9445 );
and \U$13209 ( \22032_22331 , RIee2f698_4998, \9148_9447 );
and \U$13210 ( \22033_22332 , RIfc52298_5957, \9150_9449 );
and \U$13211 ( \22034_22333 , RIee2d4d8_4974, \9152_9451 );
and \U$13212 ( \22035_22334 , RIdf35368_1982, \9154_9453 );
and \U$13213 ( \22036_22335 , RIdf32ed8_1956, \9156_9455 );
and \U$13214 ( \22037_22336 , RIdf30e80_1933, \9158_9457 );
and \U$13215 ( \22038_22337 , RIfe85ab8_7865, \9160_9459 );
or \U$13216 ( \22039_22338 , \21975_22274 , \21976_22275 , \21977_22276 , \21978_22277 , \21979_22278 , \21980_22279 , \21981_22280 , \21982_22281 , \21983_22282 , \21984_22283 , \21985_22284 , \21986_22285 , \21987_22286 , \21988_22287 , \21989_22288 , \21990_22289 , \21991_22290 , \21992_22291 , \21993_22292 , \21994_22293 , \21995_22294 , \21996_22295 , \21997_22296 , \21998_22297 , \21999_22298 , \22000_22299 , \22001_22300 , \22002_22301 , \22003_22302 , \22004_22303 , \22005_22304 , \22006_22305 , \22007_22306 , \22008_22307 , \22009_22308 , \22010_22309 , \22011_22310 , \22012_22311 , \22013_22312 , \22014_22313 , \22015_22314 , \22016_22315 , \22017_22316 , \22018_22317 , \22019_22318 , \22020_22319 , \22021_22320 , \22022_22321 , \22023_22322 , \22024_22323 , \22025_22324 , \22026_22325 , \22027_22326 , \22028_22327 , \22029_22328 , \22030_22329 , \22031_22330 , \22032_22331 , \22033_22332 , \22034_22333 , \22035_22334 , \22036_22335 , \22037_22336 , \22038_22337 );
and \U$13217 ( \22040_22339 , RIee2b8b8_4954, \9163_9462 );
and \U$13218 ( \22041_22340 , RIee29f68_4936, \9165_9464 );
and \U$13219 ( \22042_22341 , RIee28bb8_4922, \9167_9466 );
and \U$13220 ( \22043_22342 , RIee27970_4909, \9169_9468 );
and \U$13221 ( \22044_22343 , RIdf2a0d0_1855, \9171_9470 );
and \U$13222 ( \22045_22344 , RIfe84e10_7856, \9173_9472 );
and \U$13223 ( \22046_22345 , RIdf262f0_1811, \9175_9474 );
and \U$13224 ( \22047_22346 , RIfe84ca8_7855, \9177_9476 );
and \U$13225 ( \22048_22347 , RIee27100_4903, \9179_9478 );
and \U$13226 ( \22049_22348 , RIee26b60_4899, \9181_9480 );
and \U$13227 ( \22050_22349 , RIfcd32f8_7425, \9183_9482 );
and \U$13228 ( \22051_22350 , RIee265c0_4895, \9185_9484 );
and \U$13229 ( \22052_22351 , RIfc9e300_6822, \9187_9486 );
and \U$13230 ( \22053_22352 , RIdf1f540_1733, \9189_9488 );
and \U$13231 ( \22054_22353 , RIee25eb8_4890, \9191_9490 );
and \U$13232 ( \22055_22354 , RIfe84b40_7854, \9193_9492 );
and \U$13233 ( \22056_22355 , RIdf16b70_1635, \9195_9494 );
and \U$13234 ( \22057_22356 , RIdf13e70_1603, \9197_9496 );
and \U$13235 ( \22058_22357 , RIdf11170_1571, \9199_9498 );
and \U$13236 ( \22059_22358 , RIdf0e470_1539, \9201_9500 );
and \U$13237 ( \22060_22359 , RIdf0b770_1507, \9203_9502 );
and \U$13238 ( \22061_22360 , RIdf08a70_1475, \9205_9504 );
and \U$13239 ( \22062_22361 , RIdf05d70_1443, \9207_9506 );
and \U$13240 ( \22063_22362 , RIdf03070_1411, \9209_9508 );
and \U$13241 ( \22064_22363 , RIdefd670_1347, \9211_9510 );
and \U$13242 ( \22065_22364 , RIdefa970_1315, \9213_9512 );
and \U$13243 ( \22066_22365 , RIdef7c70_1283, \9215_9514 );
and \U$13244 ( \22067_22366 , RIdef4f70_1251, \9217_9516 );
and \U$13245 ( \22068_22367 , RIdef2270_1219, \9219_9518 );
and \U$13246 ( \22069_22368 , RIdeef570_1187, \9221_9520 );
and \U$13247 ( \22070_22369 , RIdeec870_1155, \9223_9522 );
and \U$13248 ( \22071_22370 , RIdee9b70_1123, \9225_9524 );
and \U$13249 ( \22072_22371 , RIfec0348_8307, \9227_9526 );
and \U$13250 ( \22073_22372 , RIfcb54d8_7085, \9229_9528 );
and \U$13251 ( \22074_22373 , RIee23cf8_4866, \9231_9530 );
and \U$13252 ( \22075_22374 , RIfc54e30_5988, \9233_9532 );
and \U$13253 ( \22076_22375 , RIfec0078_8305, \9235_9534 );
and \U$13254 ( \22077_22376 , RIdee2988_1042, \9237_9536 );
and \U$13255 ( \22078_22377 , RIfec01e0_8306, \9239_9538 );
and \U$13256 ( \22079_22378 , RIdede770_995, \9241_9540 );
and \U$13257 ( \22080_22379 , RIfcd7ee8_7479, \9243_9542 );
and \U$13258 ( \22081_22380 , RIfcd43d8_7437, \9245_9544 );
and \U$13259 ( \22082_22381 , RIfc88eb0_6580, \9247_9546 );
and \U$13260 ( \22083_22382 , RIfc9e5d0_6824, \9249_9548 );
and \U$13261 ( \22084_22383 , RIded9478_936, \9251_9550 );
and \U$13262 ( \22085_22384 , RIded6fe8_910, \9253_9552 );
and \U$13263 ( \22086_22385 , RIded50f8_888, \9255_9554 );
and \U$13264 ( \22087_22386 , RIfeab330_8264, \9257_9556 );
and \U$13265 ( \22088_22387 , RIded03a0_833, \9259_9558 );
and \U$13266 ( \22089_22388 , RIdecd6a0_801, \9261_9560 );
and \U$13267 ( \22090_22389 , RIdeca9a0_769, \9263_9562 );
and \U$13268 ( \22091_22390 , RIdec7ca0_737, \9265_9564 );
and \U$13269 ( \22092_22391 , RIdeb41a0_513, \9267_9566 );
and \U$13270 ( \22093_22392 , RIde95f48_321, \9269_9568 );
and \U$13271 ( \22094_22393 , RIe16dda8_2627, \9271_9570 );
and \U$13272 ( \22095_22394 , RIe159ba0_2398, \9273_9572 );
and \U$13273 ( \22096_22395 , RIe1433a0_2142, \9275_9574 );
and \U$13274 ( \22097_22396 , RIdf37d98_2012, \9277_9576 );
and \U$13275 ( \22098_22397 , RIdf2c3f8_1880, \9279_9578 );
and \U$13276 ( \22099_22398 , RIdf1cc78_1704, \9281_9580 );
and \U$13277 ( \22100_22399 , RIdf00370_1379, \9283_9582 );
and \U$13278 ( \22101_22400 , RIdee6e70_1091, \9285_9584 );
and \U$13279 ( \22102_22401 , RIdedbbd8_964, \9287_9586 );
and \U$13280 ( \22103_22402 , RIde7be90_194, \9289_9588 );
or \U$13281 ( \22104_22403 , \22040_22339 , \22041_22340 , \22042_22341 , \22043_22342 , \22044_22343 , \22045_22344 , \22046_22345 , \22047_22346 , \22048_22347 , \22049_22348 , \22050_22349 , \22051_22350 , \22052_22351 , \22053_22352 , \22054_22353 , \22055_22354 , \22056_22355 , \22057_22356 , \22058_22357 , \22059_22358 , \22060_22359 , \22061_22360 , \22062_22361 , \22063_22362 , \22064_22363 , \22065_22364 , \22066_22365 , \22067_22366 , \22068_22367 , \22069_22368 , \22070_22369 , \22071_22370 , \22072_22371 , \22073_22372 , \22074_22373 , \22075_22374 , \22076_22375 , \22077_22376 , \22078_22377 , \22079_22378 , \22080_22379 , \22081_22380 , \22082_22381 , \22083_22382 , \22084_22383 , \22085_22384 , \22086_22385 , \22087_22386 , \22088_22387 , \22089_22388 , \22090_22389 , \22091_22390 , \22092_22391 , \22093_22392 , \22094_22393 , \22095_22394 , \22096_22395 , \22097_22396 , \22098_22397 , \22099_22398 , \22100_22399 , \22101_22400 , \22102_22401 , \22103_22402 );
or \U$13282 ( \22105_22404 , \22039_22338 , \22104_22403 );
_DC \g5885/U$1 ( \22106 , \22105_22404 , \9298_9597 );
and \U$13283 ( \22107_22406 , RIe19d238_3165, \8760_9059 );
and \U$13284 ( \22108_22407 , RIe19a538_3133, \8762_9061 );
and \U$13285 ( \22109_22408 , RIf145658_5249, \8764_9063 );
and \U$13286 ( \22110_22409 , RIe197838_3101, \8766_9065 );
and \U$13287 ( \22111_22410 , RIf1446e0_5238, \8768_9067 );
and \U$13288 ( \22112_22411 , RIe194b38_3069, \8770_9069 );
and \U$13289 ( \22113_22412 , RIe191e38_3037, \8772_9071 );
and \U$13290 ( \22114_22413 , RIe18f138_3005, \8774_9073 );
and \U$13291 ( \22115_22414 , RIe189738_2941, \8776_9075 );
and \U$13292 ( \22116_22415 , RIe186a38_2909, \8778_9077 );
and \U$13293 ( \22117_22416 , RIf143600_5226, \8780_9079 );
and \U$13294 ( \22118_22417 , RIe183d38_2877, \8782_9081 );
and \U$13295 ( \22119_22418 , RIf142c28_5219, \8784_9083 );
and \U$13296 ( \22120_22419 , RIe181038_2845, \8786_9085 );
and \U$13297 ( \22121_22420 , RIe17e338_2813, \8788_9087 );
and \U$13298 ( \22122_22421 , RIe17b638_2781, \8790_9089 );
and \U$13299 ( \22123_22422 , RIf1420e8_5211, \8792_9091 );
and \U$13300 ( \22124_22423 , RIf140a68_5195, \8794_9093 );
and \U$13301 ( \22125_22424 , RIf1401f8_5189, \8796_9095 );
and \U$13302 ( \22126_22425 , RIfebff10_8304, \8798_9097 );
and \U$13303 ( \22127_22426 , RIf13faf0_5184, \8800_9099 );
and \U$13304 ( \22128_22427 , RIf13ee48_5175, \8802_9101 );
and \U$13305 ( \22129_22428 , RIee3e2d8_5166, \8804_9103 );
and \U$13306 ( \22130_22429 , RIee3d1f8_5154, \8806_9105 );
and \U$13307 ( \22131_22430 , RIee3c118_5142, \8808_9107 );
and \U$13308 ( \22132_22431 , RIee3b038_5130, \8810_9109 );
and \U$13309 ( \22133_22432 , RIee39c88_5116, \8812_9111 );
and \U$13310 ( \22134_22433 , RIfe838f8_7841, \8814_9113 );
and \U$13311 ( \22135_22434 , RIf1701c8_5735, \8816_9115 );
and \U$13312 ( \22136_22435 , RIfc5ab00_6054, \8818_9117 );
and \U$13313 ( \22137_22436 , RIf16e008_5711, \8820_9119 );
and \U$13314 ( \22138_22437 , RIfcb0e88_7035, \8822_9121 );
and \U$13315 ( \22139_22438 , RIf16caf0_5696, \8824_9123 );
and \U$13316 ( \22140_22439 , RIe223590_4692, \8826_9125 );
and \U$13317 ( \22141_22440 , RIf16bce0_5686, \8828_9127 );
and \U$13318 ( \22142_22441 , RIe220890_4660, \8830_9129 );
and \U$13319 ( \22143_22442 , RIf16ac00_5674, \8832_9131 );
and \U$13320 ( \22144_22443 , RIe21db90_4628, \8834_9133 );
and \U$13321 ( \22145_22444 , RIe218190_4564, \8836_9135 );
and \U$13322 ( \22146_22445 , RIe215490_4532, \8838_9137 );
and \U$13323 ( \22147_22446 , RIf16a228_5667, \8840_9139 );
and \U$13324 ( \22148_22447 , RIe212790_4500, \8842_9141 );
and \U$13325 ( \22149_22448 , RIf168fe0_5654, \8844_9143 );
and \U$13326 ( \22150_22449 , RIe20fa90_4468, \8846_9145 );
and \U$13327 ( \22151_22450 , RIf167d98_5641, \8848_9147 );
and \U$13328 ( \22152_22451 , RIe20cd90_4436, \8850_9149 );
and \U$13329 ( \22153_22452 , RIe20a090_4404, \8852_9151 );
and \U$13330 ( \22154_22453 , RIe207390_4372, \8854_9153 );
and \U$13331 ( \22155_22454 , RIf1670f0_5632, \8856_9155 );
and \U$13332 ( \22156_22455 , RIf165ea8_5619, \8858_9157 );
and \U$13333 ( \22157_22456 , RIe202200_4314, \8860_9159 );
and \U$13334 ( \22158_22457 , RIfe83e98_7845, \8862_9161 );
and \U$13335 ( \22159_22458 , RIf164f30_5608, \8864_9163 );
and \U$13336 ( \22160_22459 , RIf1643f0_5600, \8866_9165 );
and \U$13337 ( \22161_22460 , RIfce8310_7664, \8868_9167 );
and \U$13338 ( \22162_22461 , RIf161df8_5573, \8870_9169 );
and \U$13339 ( \22163_22462 , RIf15ff08_5551, \8872_9171 );
and \U$13340 ( \22164_22463 , RIf15e018_5529, \8874_9173 );
and \U$13341 ( \22165_22464 , RIfe83d30_7844, \8876_9175 );
and \U$13342 ( \22166_22465 , RIfe84000_7846, \8878_9177 );
and \U$13343 ( \22167_22466 , RIf15cb00_5514, \8880_9179 );
and \U$13344 ( \22168_22467 , RIf15b5e8_5499, \8882_9181 );
and \U$13345 ( \22169_22468 , RIf15a508_5487, \8884_9183 );
and \U$13346 ( \22170_22469 , RIfc887a8_6575, \8886_9185 );
or \U$13347 ( \22171_22470 , \22107_22406 , \22108_22407 , \22109_22408 , \22110_22409 , \22111_22410 , \22112_22411 , \22113_22412 , \22114_22413 , \22115_22414 , \22116_22415 , \22117_22416 , \22118_22417 , \22119_22418 , \22120_22419 , \22121_22420 , \22122_22421 , \22123_22422 , \22124_22423 , \22125_22424 , \22126_22425 , \22127_22426 , \22128_22427 , \22129_22428 , \22130_22429 , \22131_22430 , \22132_22431 , \22133_22432 , \22134_22433 , \22135_22434 , \22136_22435 , \22137_22436 , \22138_22437 , \22139_22438 , \22140_22439 , \22141_22440 , \22142_22441 , \22143_22442 , \22144_22443 , \22145_22444 , \22146_22445 , \22147_22446 , \22148_22447 , \22149_22448 , \22150_22449 , \22151_22450 , \22152_22451 , \22153_22452 , \22154_22453 , \22155_22454 , \22156_22455 , \22157_22456 , \22158_22457 , \22159_22458 , \22160_22459 , \22161_22460 , \22162_22461 , \22163_22462 , \22164_22463 , \22165_22464 , \22166_22465 , \22167_22466 , \22168_22467 , \22169_22468 , \22170_22469 );
and \U$13348 ( \22172_22471 , RIf158d20_5470, \8889_9188 );
and \U$13349 ( \22173_22472 , RIf157970_5456, \8891_9190 );
and \U$13350 ( \22174_22473 , RIf156cc8_5447, \8893_9192 );
and \U$13351 ( \22175_22474 , RIfe84438_7849, \8895_9194 );
and \U$13352 ( \22176_22475 , RIf156020_5438, \8897_9196 );
and \U$13353 ( \22177_22476 , RIfc51fc8_5955, \8899_9198 );
and \U$13354 ( \22178_22477 , RIf154568_5419, \8901_9200 );
and \U$13355 ( \22179_22478 , RIe1f51e0_4166, \8903_9202 );
and \U$13356 ( \22180_22479 , RIf153050_5404, \8905_9204 );
and \U$13357 ( \22181_22480 , RIf1519d0_5388, \8907_9206 );
and \U$13358 ( \22182_22481 , RIf150788_5375, \8909_9208 );
and \U$13359 ( \22183_22482 , RIfe842d0_7848, \8911_9210 );
and \U$13360 ( \22184_22483 , RIf14f810_5364, \8913_9212 );
and \U$13361 ( \22185_22484 , RIf14eb68_5355, \8915_9214 );
and \U$13362 ( \22186_22485 , RIf14dd58_5345, \8917_9216 );
and \U$13363 ( \22187_22486 , RIfe84168_7847, \8919_9218 );
and \U$13364 ( \22188_22487 , RIe1eb2f8_4053, \8921_9220 );
and \U$13365 ( \22189_22488 , RIe1e85f8_4021, \8923_9222 );
and \U$13366 ( \22190_22489 , RIe1e58f8_3989, \8925_9224 );
and \U$13367 ( \22191_22490 , RIe1e2bf8_3957, \8927_9226 );
and \U$13368 ( \22192_22491 , RIe1dfef8_3925, \8929_9228 );
and \U$13369 ( \22193_22492 , RIe1dd1f8_3893, \8931_9230 );
and \U$13370 ( \22194_22493 , RIe1da4f8_3861, \8933_9232 );
and \U$13371 ( \22195_22494 , RIe1d77f8_3829, \8935_9234 );
and \U$13372 ( \22196_22495 , RIe1d1df8_3765, \8937_9236 );
and \U$13373 ( \22197_22496 , RIe1cf0f8_3733, \8939_9238 );
and \U$13374 ( \22198_22497 , RIe1cc3f8_3701, \8941_9240 );
and \U$13375 ( \22199_22498 , RIe1c96f8_3669, \8943_9242 );
and \U$13376 ( \22200_22499 , RIe1c69f8_3637, \8945_9244 );
and \U$13377 ( \22201_22500 , RIe1c3cf8_3605, \8947_9246 );
and \U$13378 ( \22202_22501 , RIe1c0ff8_3573, \8949_9248 );
and \U$13379 ( \22203_22502 , RIe1be2f8_3541, \8951_9250 );
and \U$13380 ( \22204_22503 , RIf14c840_5330, \8953_9252 );
and \U$13381 ( \22205_22504 , RIf14b5f8_5317, \8955_9254 );
and \U$13382 ( \22206_22505 , RIfe83a60_7842, \8957_9256 );
and \U$13383 ( \22207_22506 , RIfe849d8_7853, \8959_9258 );
and \U$13384 ( \22208_22507 , RIfc74168_6343, \8961_9260 );
and \U$13385 ( \22209_22508 , RIf149b40_5298, \8963_9262 );
and \U$13386 ( \22210_22509 , RIfe83bc8_7843, \8965_9264 );
and \U$13387 ( \22211_22510 , RIfe84708_7851, \8967_9266 );
and \U$13388 ( \22212_22511 , RIf148d30_5288, \8969_9268 );
and \U$13389 ( \22213_22512 , RIf147ae8_5275, \8971_9270 );
and \U$13390 ( \22214_22513 , RIfe84870_7852, \8973_9272 );
and \U$13391 ( \22215_22514 , RIe1b0900_3386, \8975_9274 );
and \U$13392 ( \22216_22515 , RIf146fa8_5267, \8977_9276 );
and \U$13393 ( \22217_22516 , RIf146300_5258, \8979_9278 );
and \U$13394 ( \22218_22517 , RIfe845a0_7850, \8981_9280 );
and \U$13395 ( \22219_22518 , RIfe83790_7840, \8983_9282 );
and \U$13396 ( \22220_22519 , RIe1a8638_3293, \8985_9284 );
and \U$13397 ( \22221_22520 , RIe1a5938_3261, \8987_9286 );
and \U$13398 ( \22222_22521 , RIe1a2c38_3229, \8989_9288 );
and \U$13399 ( \22223_22522 , RIe19ff38_3197, \8991_9290 );
and \U$13400 ( \22224_22523 , RIe18c438_2973, \8993_9292 );
and \U$13401 ( \22225_22524 , RIe178938_2749, \8995_9294 );
and \U$13402 ( \22226_22525 , RIe226290_4724, \8997_9296 );
and \U$13403 ( \22227_22526 , RIe21ae90_4596, \8999_9298 );
and \U$13404 ( \22228_22527 , RIe204690_4340, \9001_9300 );
and \U$13405 ( \22229_22528 , RIe1fe6f0_4272, \9003_9302 );
and \U$13406 ( \22230_22529 , RIe1f7aa8_4195, \9005_9304 );
and \U$13407 ( \22231_22530 , RIe1f05f0_4112, \9007_9306 );
and \U$13408 ( \22232_22531 , RIe1d4af8_3797, \9009_9308 );
and \U$13409 ( \22233_22532 , RIe1bb5f8_3509, \9011_9310 );
and \U$13410 ( \22234_22533 , RIe1ae470_3360, \9013_9312 );
and \U$13411 ( \22235_22534 , RIe170aa8_2659, \9015_9314 );
or \U$13412 ( \22236_22535 , \22172_22471 , \22173_22472 , \22174_22473 , \22175_22474 , \22176_22475 , \22177_22476 , \22178_22477 , \22179_22478 , \22180_22479 , \22181_22480 , \22182_22481 , \22183_22482 , \22184_22483 , \22185_22484 , \22186_22485 , \22187_22486 , \22188_22487 , \22189_22488 , \22190_22489 , \22191_22490 , \22192_22491 , \22193_22492 , \22194_22493 , \22195_22494 , \22196_22495 , \22197_22496 , \22198_22497 , \22199_22498 , \22200_22499 , \22201_22500 , \22202_22501 , \22203_22502 , \22204_22503 , \22205_22504 , \22206_22505 , \22207_22506 , \22208_22507 , \22209_22508 , \22210_22509 , \22211_22510 , \22212_22511 , \22213_22512 , \22214_22513 , \22215_22514 , \22216_22515 , \22217_22516 , \22218_22517 , \22219_22518 , \22220_22519 , \22221_22520 , \22222_22521 , \22223_22522 , \22224_22523 , \22225_22524 , \22226_22525 , \22227_22526 , \22228_22527 , \22229_22528 , \22230_22529 , \22231_22530 , \22232_22531 , \22233_22532 , \22234_22533 , \22235_22534 );
or \U$13413 ( \22237_22536 , \22171_22470 , \22236_22535 );
_DC \g5909/U$1 ( \22238 , \22237_22536 , \9024_9323 );
xor g590a_GF_PartitionCandidate( \22239_22538_nG590a , \22106 , \22238 );
buf \U$13414 ( \22240_22539 , \22239_22538_nG590a );
xor \U$13415 ( \22241_22540 , \22240_22539 , \21800_22102 );
not \U$13416 ( \22242_22541 , \21801_22103 );
and \U$13417 ( \22243_22542 , \22241_22540 , \22242_22541 );
and \U$13418 ( \22244_22543 , \10385_10687 , \22243_22542 );
and \U$13419 ( \22245_22544 , \10686_10988 , \21801_22103 );
nor \U$13420 ( \22246_22545 , \22244_22543 , \22245_22544 );
and \U$13421 ( \22247_22546 , \21800_22102 , \20703_21002 );
not \U$13422 ( \22248_22547 , \22247_22546 );
and \U$13423 ( \22249_22548 , \22240_22539 , \22248_22547 );
xnor \U$13424 ( \22250_22549 , \22246_22545 , \22249_22548 );
xor \U$13425 ( \22251_22550 , \21974_22273 , \22250_22549 );
xor \U$13426 ( \22252_22551 , \21965_22264 , \22251_22550 );
and \U$13427 ( \22253_22552 , \21788_22090 , \10681_10983 );
_DC \g65b0/U$1 ( \22254 , \22105_22404 , \9298_9597 );
_DC \g65b1/U$1 ( \22255 , \22237_22536 , \9024_9323 );
and g65b2_GF_PartitionCandidate( \22256_22555_nG65b2 , \22254 , \22255 );
buf \U$13428 ( \22257_22556 , \22256_22555_nG65b2 );
and \U$13429 ( \22258_22557 , \22257_22556 , \10389_10691 );
nor \U$13430 ( \22259_22558 , \22253_22552 , \22258_22557 );
xnor \U$13431 ( \22260_22559 , \22259_22558 , \10678_10980 );
not \U$13432 ( \22261_22560 , \21802_22104 );
and \U$13433 ( \22262_22561 , \22261_22560 , \22249_22548 );
xor \U$13434 ( \22263_22562 , \22260_22559 , \22262_22561 );
and \U$13435 ( \22264_22563 , \21791_22093 , \21795_22097 );
and \U$13436 ( \22265_22564 , \21795_22097 , \21802_22104 );
and \U$13437 ( \22266_22565 , \21791_22093 , \21802_22104 );
or \U$13438 ( \22267_22566 , \22264_22563 , \22265_22564 , \22266_22565 );
xor \U$13439 ( \22268_22567 , \22263_22562 , \22267_22566 );
and \U$13440 ( \22269_22568 , \21484_21786 , \21488_21790 );
and \U$13441 ( \22270_22569 , \21488_21790 , \21493_21795 );
and \U$13442 ( \22271_22570 , \21484_21786 , \21493_21795 );
or \U$13443 ( \22272_22571 , \22269_22568 , \22270_22569 , \22271_22570 );
xor \U$13444 ( \22273_22572 , \22268_22567 , \22272_22571 );
xor \U$13445 ( \22274_22573 , \22252_22551 , \22273_22572 );
xor \U$13446 ( \22275_22574 , \21961_22260 , \22274_22573 );
and \U$13447 ( \22276_22575 , \21521_21823 , \21803_22105 );
and \U$13448 ( \22277_22576 , \21803_22105 , \21818_22120 );
and \U$13449 ( \22278_22577 , \21521_21823 , \21818_22120 );
or \U$13450 ( \22279_22578 , \22276_22575 , \22277_22576 , \22278_22577 );
and \U$13451 ( \22280_22579 , \21480_21782 , \21494_21796 );
and \U$13452 ( \22281_22580 , \21494_21796 , \21506_21808 );
and \U$13453 ( \22282_22581 , \21480_21782 , \21506_21808 );
or \U$13454 ( \22283_22582 , \22280_22579 , \22281_22580 , \22282_22581 );
xor \U$13455 ( \22284_22583 , \22279_22578 , \22283_22582 );
and \U$13456 ( \22285_22584 , \21808_22110 , \21812_22114 );
and \U$13457 ( \22286_22585 , \21812_22114 , \21817_22119 );
and \U$13458 ( \22287_22586 , \21808_22110 , \21817_22119 );
or \U$13459 ( \22288_22587 , \22285_22584 , \22286_22585 , \22287_22586 );
and \U$13460 ( \22289_22588 , \18730_19032 , \12491_12790 );
and \U$13461 ( \22290_22589 , \19259_19558 , \12159_12461 );
nor \U$13462 ( \22291_22590 , \22289_22588 , \22290_22589 );
xnor \U$13463 ( \22292_22591 , \22291_22590 , \12481_12780 );
and \U$13464 ( \22293_22592 , \14648_14950 , \16333_16635 );
and \U$13465 ( \22294_22593 , \15022_15321 , \15999_16301 );
nor \U$13466 ( \22295_22594 , \22293_22592 , \22294_22593 );
xnor \U$13467 ( \22296_22595 , \22295_22594 , \16323_16625 );
xor \U$13468 ( \22297_22596 , \22292_22591 , \22296_22595 );
and \U$13469 ( \22298_22597 , \13377_13679 , \17791_18090 );
and \U$13470 ( \22299_22598 , \13725_14024 , \17353_17655 );
nor \U$13471 ( \22300_22599 , \22298_22597 , \22299_22598 );
xnor \U$13472 ( \22301_22600 , \22300_22599 , \17747_18046 );
xor \U$13473 ( \22302_22601 , \22297_22596 , \22301_22600 );
xor \U$13474 ( \22303_22602 , \22288_22587 , \22302_22601 );
and \U$13475 ( \22304_22603 , \17325_17627 , \13755_14054 );
and \U$13476 ( \22305_22604 , \17736_18035 , \13390_13692 );
nor \U$13477 ( \22306_22605 , \22304_22603 , \22305_22604 );
xnor \U$13478 ( \22307_22606 , \22306_22605 , \13736_14035 );
and \U$13479 ( \22308_22607 , \12146_12448 , \19235_19534 );
and \U$13480 ( \22309_22608 , \12470_12769 , \18743_19045 );
nor \U$13481 ( \22310_22609 , \22308_22607 , \22309_22608 );
xnor \U$13482 ( \22311_22610 , \22310_22609 , \19241_19540 );
xor \U$13483 ( \22312_22611 , \22307_22606 , \22311_22610 );
and \U$13484 ( \22313_22612 , \10968_11270 , \20706_21005 );
and \U$13485 ( \22314_22613 , \11287_11586 , \20255_20557 );
nor \U$13486 ( \22315_22614 , \22313_22612 , \22314_22613 );
xnor \U$13487 ( \22316_22615 , \22315_22614 , \20712_21011 );
xor \U$13488 ( \22317_22616 , \22312_22611 , \22316_22615 );
xor \U$13489 ( \22318_22617 , \22303_22602 , \22317_22616 );
xor \U$13490 ( \22319_22618 , \22284_22583 , \22318_22617 );
xor \U$13491 ( \22320_22619 , \22275_22574 , \22319_22618 );
and \U$13492 ( \22321_22620 , \21476_21778 , \21507_21809 );
and \U$13493 ( \22322_22621 , \21507_21809 , \21820_22122 );
and \U$13494 ( \22323_22622 , \21476_21778 , \21820_22122 );
or \U$13495 ( \22324_22623 , \22321_22620 , \22322_22621 , \22323_22622 );
xor \U$13496 ( \22325_22624 , \22320_22619 , \22324_22623 );
and \U$13497 ( \22326_22625 , \21472_21774 , \21821_22123 );
and \U$13498 ( \22327_22626 , \21822_22124 , \21825_22127 );
or \U$13499 ( \22328_22627 , \22326_22625 , \22327_22626 );
xor \U$13500 ( \22329_22628 , \22325_22624 , \22328_22627 );
buf g9bd5_GF_PartitionCandidate( \22330_22629_nG9bd5 , \22329_22628 );
and \U$13501 ( \22331_22630 , \10402_10704 , \22330_22629_nG9bd5 );
or \U$13502 ( \22332_22631 , \21957_22256 , \22331_22630 );
xor \U$13503 ( \22333_22632 , \10399_10703 , \22332_22631 );
buf \U$13504 ( \22334_22633 , \22333_22632 );
buf \U$13506 ( \22335_22634 , \22334_22633 );
xor \U$13507 ( \22336_22635 , \21956_22255 , \22335_22634 );
buf \U$13508 ( \22337_22636 , \22336_22635 );
xor \U$13509 ( \22338_22637 , \21945_22244 , \22337_22636 );
and \U$13510 ( \22339_22638 , \21373_21675 , \21407_21709 );
and \U$13511 ( \22340_22639 , \21373_21675 , \21448_21750 );
and \U$13512 ( \22341_22640 , \21407_21709 , \21448_21750 );
or \U$13513 ( \22342_22641 , \22339_22638 , \22340_22639 , \22341_22640 );
buf \U$13514 ( \22343_22642 , \22342_22641 );
xor \U$13515 ( \22344_22643 , \22338_22637 , \22343_22642 );
and \U$13516 ( \22345_22644 , \21848_22150 , \22344_22643 );
and \U$13517 ( \22346_22645 , \21838_22140 , \21842_22144 );
and \U$13518 ( \22347_22646 , \21838_22140 , \21847_22149 );
and \U$13519 ( \22348_22647 , \21842_22144 , \21847_22149 );
or \U$13520 ( \22349_22648 , \22346_22645 , \22347_22646 , \22348_22647 );
xor \U$13521 ( \22350_22649 , \22345_22644 , \22349_22648 );
and \U$13522 ( \22351_22650 , RIdec53d8_708, \8760_9059 );
and \U$13523 ( \22352_22651 , RIdec26d8_676, \8762_9061 );
and \U$13524 ( \22353_22652 , RIee20080_4823, \8764_9063 );
and \U$13525 ( \22354_22653 , RIdebf9d8_644, \8766_9065 );
and \U$13526 ( \22355_22654 , RIee1f3d8_4814, \8768_9067 );
and \U$13527 ( \22356_22655 , RIdebccd8_612, \8770_9069 );
and \U$13528 ( \22357_22656 , RIdeb9fd8_580, \8772_9071 );
and \U$13529 ( \22358_22657 , RIdeb72d8_548, \8774_9073 );
and \U$13530 ( \22359_22658 , RIee1ee38_4810, \8776_9075 );
and \U$13531 ( \22360_22659 , RIdeb18d8_484, \8778_9077 );
and \U$13532 ( \22361_22660 , RIee1e898_4806, \8780_9079 );
and \U$13533 ( \22362_22661 , RIdeaebd8_452, \8782_9081 );
and \U$13534 ( \22363_22662 , RIee1da88_4796, \8784_9083 );
and \U$13535 ( \22364_22663 , RIdeaa420_420, \8786_9085 );
and \U$13536 ( \22365_22664 , RIdea3b20_388, \8788_9087 );
and \U$13537 ( \22366_22665 , RIde9d220_356, \8790_9089 );
and \U$13538 ( \22367_22666 , RIee1cde0_4787, \8792_9091 );
and \U$13539 ( \22368_22667 , RIee1bd00_4775, \8794_9093 );
and \U$13540 ( \22369_22668 , RIee1b490_4769, \8796_9095 );
and \U$13541 ( \22370_22669 , RIfcd8a28_7487, \8798_9097 );
and \U$13542 ( \22371_22670 , RIde91088_297, \8800_9099 );
and \U$13543 ( \22372_22671 , RIde8d8c0_280, \8802_9101 );
and \U$13544 ( \22373_22672 , RIfe7dac0_7774, \8804_9103 );
and \U$13545 ( \22374_22673 , RIfe7d958_7773, \8806_9105 );
and \U$13546 ( \22375_22674 , RIee1a518_4758, \8808_9107 );
and \U$13547 ( \22376_22675 , RIee19e10_4753, \8810_9109 );
and \U$13548 ( \22377_22676 , RIee19b40_4751, \8812_9111 );
and \U$13549 ( \22378_22677 , RIfc768c8_6371, \8814_9113 );
and \U$13550 ( \22379_22678 , RIfcd05f8_7393, \8816_9115 );
and \U$13551 ( \22380_22679 , RIfe7dd90_7776, \8818_9117 );
and \U$13552 ( \22381_22680 , RIee38770_5101, \8820_9119 );
and \U$13553 ( \22382_22681 , RIfe7dc28_7775, \8822_9121 );
and \U$13554 ( \22383_22682 , RIe1653d8_2529, \8824_9123 );
and \U$13555 ( \22384_22683 , RIe1626d8_2497, \8826_9125 );
and \U$13556 ( \22385_22684 , RIee373c0_5087, \8828_9127 );
and \U$13557 ( \22386_22685 , RIe15f9d8_2465, \8830_9129 );
and \U$13558 ( \22387_22686 , RIee362e0_5075, \8832_9131 );
and \U$13559 ( \22388_22687 , RIe15ccd8_2433, \8834_9133 );
and \U$13560 ( \22389_22688 , RIe1572d8_2369, \8836_9135 );
and \U$13561 ( \22390_22689 , RIe1545d8_2337, \8838_9137 );
and \U$13562 ( \22391_22690 , RIfe7def8_7777, \8840_9139 );
and \U$13563 ( \22392_22691 , RIe1518d8_2305, \8842_9141 );
and \U$13564 ( \22393_22692 , RIfebdeb8_8281, \8844_9143 );
and \U$13565 ( \22394_22693 , RIe14ebd8_2273, \8846_9145 );
and \U$13566 ( \22395_22694 , RIfc649e8_6167, \8848_9147 );
and \U$13567 ( \22396_22695 , RIe14bed8_2241, \8850_9149 );
and \U$13568 ( \22397_22696 , RIe1491d8_2209, \8852_9151 );
and \U$13569 ( \22398_22697 , RIe1464d8_2177, \8854_9153 );
and \U$13570 ( \22399_22698 , RIfe7d7f0_7772, \8856_9155 );
and \U$13571 ( \22400_22699 , RIfe7d688_7771, \8858_9157 );
and \U$13572 ( \22401_22700 , RIee32230_5029, \8860_9159 );
and \U$13573 ( \22402_22701 , RIfceb9e8_7703, \8862_9161 );
and \U$13574 ( \22403_22702 , RIfebdd50_8280, \8864_9163 );
and \U$13575 ( \22404_22703 , RIfe7d520_7770, \8866_9165 );
and \U$13576 ( \22405_22704 , RIfebdbe8_8279, \8868_9167 );
and \U$13577 ( \22406_22705 , RIfe7d3b8_7769, \8870_9169 );
and \U$13578 ( \22407_22706 , RIfc734c0_6334, \8872_9171 );
and \U$13579 ( \22408_22707 , RIee2f968_5000, \8874_9173 );
and \U$13580 ( \22409_22708 , RIfccfab8_7385, \8876_9175 );
and \U$13581 ( \22410_22709 , RIee2d7a8_4976, \8878_9177 );
and \U$13582 ( \22411_22710 , RIdf357a0_1985, \8880_9179 );
and \U$13583 ( \22412_22711 , RIdf33310_1959, \8882_9181 );
and \U$13584 ( \22413_22712 , RIdf312b8_1936, \8884_9183 );
and \U$13585 ( \22414_22713 , RIdf2f0f8_1912, \8886_9185 );
or \U$13586 ( \22415_22714 , \22351_22650 , \22352_22651 , \22353_22652 , \22354_22653 , \22355_22654 , \22356_22655 , \22357_22656 , \22358_22657 , \22359_22658 , \22360_22659 , \22361_22660 , \22362_22661 , \22363_22662 , \22364_22663 , \22365_22664 , \22366_22665 , \22367_22666 , \22368_22667 , \22369_22668 , \22370_22669 , \22371_22670 , \22372_22671 , \22373_22672 , \22374_22673 , \22375_22674 , \22376_22675 , \22377_22676 , \22378_22677 , \22379_22678 , \22380_22679 , \22381_22680 , \22382_22681 , \22383_22682 , \22384_22683 , \22385_22684 , \22386_22685 , \22387_22686 , \22388_22687 , \22389_22688 , \22390_22689 , \22391_22690 , \22392_22691 , \22393_22692 , \22394_22693 , \22395_22694 , \22396_22695 , \22397_22696 , \22398_22697 , \22399_22698 , \22400_22699 , \22401_22700 , \22402_22701 , \22403_22702 , \22404_22703 , \22405_22704 , \22406_22705 , \22407_22706 , \22408_22707 , \22409_22708 , \22410_22709 , \22411_22710 , \22412_22711 , \22413_22712 , \22414_22713 );
and \U$13587 ( \22416_22715 , RIee2bcf0_4957, \8889_9188 );
and \U$13588 ( \22417_22716 , RIee2a238_4938, \8891_9190 );
and \U$13589 ( \22418_22717 , RIee28e88_4924, \8893_9192 );
and \U$13590 ( \22419_22718 , RIee27c40_4911, \8895_9194 );
and \U$13591 ( \22420_22719 , RIfe7ce18_7765, \8897_9196 );
and \U$13592 ( \22421_22720 , RIfe7ccb0_7764, \8899_9198 );
and \U$13593 ( \22422_22721 , RIfe7cf80_7766, \8901_9200 );
and \U$13594 ( \22423_22722 , RIfe7cb48_7763, \8903_9202 );
and \U$13595 ( \22424_22723 , RIee27268_4904, \8905_9204 );
and \U$13596 ( \22425_22724 , RIee26e30_4901, \8907_9206 );
and \U$13597 ( \22426_22725 , RIee26890_4897, \8909_9208 );
and \U$13598 ( \22427_22726 , RIfcaa0d8_6957, \8911_9210 );
and \U$13599 ( \22428_22727 , RIee262f0_4893, \8913_9212 );
and \U$13600 ( \22429_22728 , RIfe7d250_7768, \8915_9214 );
and \U$13601 ( \22430_22729 , RIee26020_4891, \8917_9216 );
and \U$13602 ( \22431_22730 , RIfe7d0e8_7767, \8919_9218 );
and \U$13603 ( \22432_22731 , RIdf16fa8_1638, \8921_9220 );
and \U$13604 ( \22433_22732 , RIdf142a8_1606, \8923_9222 );
and \U$13605 ( \22434_22733 , RIdf115a8_1574, \8925_9224 );
and \U$13606 ( \22435_22734 , RIdf0e8a8_1542, \8927_9226 );
and \U$13607 ( \22436_22735 , RIdf0bba8_1510, \8929_9228 );
and \U$13608 ( \22437_22736 , RIdf08ea8_1478, \8931_9230 );
and \U$13609 ( \22438_22737 , RIdf061a8_1446, \8933_9232 );
and \U$13610 ( \22439_22738 , RIdf034a8_1414, \8935_9234 );
and \U$13611 ( \22440_22739 , RIdefdaa8_1350, \8937_9236 );
and \U$13612 ( \22441_22740 , RIdefada8_1318, \8939_9238 );
and \U$13613 ( \22442_22741 , RIdef80a8_1286, \8941_9240 );
and \U$13614 ( \22443_22742 , RIdef53a8_1254, \8943_9242 );
and \U$13615 ( \22444_22743 , RIdef26a8_1222, \8945_9244 );
and \U$13616 ( \22445_22744 , RIdeef9a8_1190, \8947_9246 );
and \U$13617 ( \22446_22745 , RIdeecca8_1158, \8949_9248 );
and \U$13618 ( \22447_22746 , RIdee9fa8_1126, \8951_9250 );
and \U$13619 ( \22448_22747 , RIee25648_4884, \8953_9252 );
and \U$13620 ( \22449_22748 , RIee249a0_4875, \8955_9254 );
and \U$13621 ( \22450_22749 , RIfebe020_8282, \8957_9256 );
and \U$13622 ( \22451_22750 , RIee23488_4860, \8959_9258 );
and \U$13623 ( \22452_22751 , RIfebe2f0_8284, \8961_9260 );
and \U$13624 ( \22453_22752 , RIfebe188_8283, \8963_9262 );
and \U$13625 ( \22454_22753 , RIfe7e1c8_7779, \8965_9264 );
and \U$13626 ( \22455_22754 , RIfe7e060_7778, \8967_9266 );
and \U$13627 ( \22456_22755 , RIfcbf7f8_7201, \8969_9268 );
and \U$13628 ( \22457_22756 , RIfc7aae0_6418, \8971_9270 );
and \U$13629 ( \22458_22757 , RIfc787b8_6393, \8973_9272 );
and \U$13630 ( \22459_22758 , RIfc618b0_6132, \8975_9274 );
and \U$13631 ( \22460_22759 , RIded98b0_939, \8977_9276 );
and \U$13632 ( \22461_22760 , RIded72b8_912, \8979_9278 );
and \U$13633 ( \22462_22761 , RIded5530_891, \8981_9280 );
and \U$13634 ( \22463_22762 , RIded2dd0_863, \8983_9282 );
and \U$13635 ( \22464_22763 , RIded07d8_836, \8985_9284 );
and \U$13636 ( \22465_22764 , RIdecdad8_804, \8987_9286 );
and \U$13637 ( \22466_22765 , RIdecadd8_772, \8989_9288 );
and \U$13638 ( \22467_22766 , RIdec80d8_740, \8991_9290 );
and \U$13639 ( \22468_22767 , RIdeb45d8_516, \8993_9292 );
and \U$13640 ( \22469_22768 , RIde96920_324, \8995_9294 );
and \U$13641 ( \22470_22769 , RIe16e1e0_2630, \8997_9296 );
and \U$13642 ( \22471_22770 , RIe159fd8_2401, \8999_9298 );
and \U$13643 ( \22472_22771 , RIe1437d8_2145, \9001_9300 );
and \U$13644 ( \22473_22772 , RIdf381d0_2015, \9003_9302 );
and \U$13645 ( \22474_22773 , RIdf2c830_1883, \9005_9304 );
and \U$13646 ( \22475_22774 , RIdf1d0b0_1707, \9007_9306 );
and \U$13647 ( \22476_22775 , RIdf007a8_1382, \9009_9308 );
and \U$13648 ( \22477_22776 , RIdee72a8_1094, \9011_9310 );
and \U$13649 ( \22478_22777 , RIdedc010_967, \9013_9312 );
and \U$13650 ( \22479_22778 , RIde7c868_197, \9015_9314 );
or \U$13651 ( \22480_22779 , \22416_22715 , \22417_22716 , \22418_22717 , \22419_22718 , \22420_22719 , \22421_22720 , \22422_22721 , \22423_22722 , \22424_22723 , \22425_22724 , \22426_22725 , \22427_22726 , \22428_22727 , \22429_22728 , \22430_22729 , \22431_22730 , \22432_22731 , \22433_22732 , \22434_22733 , \22435_22734 , \22436_22735 , \22437_22736 , \22438_22737 , \22439_22738 , \22440_22739 , \22441_22740 , \22442_22741 , \22443_22742 , \22444_22743 , \22445_22744 , \22446_22745 , \22447_22746 , \22448_22747 , \22449_22748 , \22450_22749 , \22451_22750 , \22452_22751 , \22453_22752 , \22454_22753 , \22455_22754 , \22456_22755 , \22457_22756 , \22458_22757 , \22459_22758 , \22460_22759 , \22461_22760 , \22462_22761 , \22463_22762 , \22464_22763 , \22465_22764 , \22466_22765 , \22467_22766 , \22468_22767 , \22469_22768 , \22470_22769 , \22471_22770 , \22472_22771 , \22473_22772 , \22474_22773 , \22475_22774 , \22476_22775 , \22477_22776 , \22478_22777 , \22479_22778 );
or \U$13652 ( \22481_22780 , \22415_22714 , \22480_22779 );
_DC \g2767/U$1 ( \22482 , \22481_22780 , \9024_9323 );
buf \U$13653 ( \22483_22782 , \22482 );
and \U$13654 ( \22484_22783 , RIe19d670_3168, \9034_9333 );
and \U$13655 ( \22485_22784 , RIe19a970_3136, \9036_9335 );
and \U$13656 ( \22486_22785 , RIfe7b630_7748, \9038_9337 );
and \U$13657 ( \22487_22786 , RIe197c70_3104, \9040_9339 );
and \U$13658 ( \22488_22787 , RIfe7b4c8_7747, \9042_9341 );
and \U$13659 ( \22489_22788 , RIe194f70_3072, \9044_9343 );
and \U$13660 ( \22490_22789 , RIe192270_3040, \9046_9345 );
and \U$13661 ( \22491_22790 , RIe18f570_3008, \9048_9347 );
and \U$13662 ( \22492_22791 , RIe189b70_2944, \9050_9349 );
and \U$13663 ( \22493_22792 , RIe186e70_2912, \9052_9351 );
and \U$13664 ( \22494_22793 , RIfe7b360_7746, \9054_9353 );
and \U$13665 ( \22495_22794 , RIe184170_2880, \9056_9355 );
and \U$13666 ( \22496_22795 , RIfe7b1f8_7745, \9058_9357 );
and \U$13667 ( \22497_22796 , RIe181470_2848, \9060_9359 );
and \U$13668 ( \22498_22797 , RIe17e770_2816, \9062_9361 );
and \U$13669 ( \22499_22798 , RIe17ba70_2784, \9064_9363 );
and \U$13670 ( \22500_22799 , RIf1423b8_5213, \9066_9365 );
and \U$13671 ( \22501_22800 , RIf140ea0_5198, \9068_9367 );
and \U$13672 ( \22502_22801 , RIf140360_5190, \9070_9369 );
and \U$13673 ( \22503_22802 , RIfe7b798_7749, \9072_9371 );
and \U$13674 ( \22504_22803 , RIf13fc58_5185, \9074_9373 );
and \U$13675 ( \22505_22804 , RIf13f280_5178, \9076_9375 );
and \U$13676 ( \22506_22805 , RIfc79460_6402, \9078_9377 );
and \U$13677 ( \22507_22806 , RIee3d4c8_5156, \9080_9379 );
and \U$13678 ( \22508_22807 , RIfe7b090_7744, \9082_9381 );
and \U$13679 ( \22509_22808 , RIfe7af28_7743, \9084_9383 );
and \U$13680 ( \22510_22809 , RIee39df0_5117, \9086_9385 );
and \U$13681 ( \22511_22810 , RIe1737a8_2691, \9088_9387 );
and \U$13682 ( \22512_22811 , RIfe7adc0_7742, \9090_9389 );
and \U$13683 ( \22513_22812 , RIfe7ac58_7741, \9092_9391 );
and \U$13684 ( \22514_22813 , RIf16e440_5714, \9094_9393 );
and \U$13685 ( \22515_22814 , RIfcb20d0_7048, \9096_9395 );
and \U$13686 ( \22516_22815 , RIfe7bd38_7753, \9098_9397 );
and \U$13687 ( \22517_22816 , RIe2239c8_4695, \9100_9399 );
and \U$13688 ( \22518_22817 , RIf16be48_5687, \9102_9401 );
and \U$13689 ( \22519_22818 , RIe220cc8_4663, \9104_9403 );
and \U$13690 ( \22520_22819 , RIf16aed0_5676, \9106_9405 );
and \U$13691 ( \22521_22820 , RIe21dfc8_4631, \9108_9407 );
and \U$13692 ( \22522_22821 , RIe2185c8_4567, \9110_9409 );
and \U$13693 ( \22523_22822 , RIe2158c8_4535, \9112_9411 );
and \U$13694 ( \22524_22823 , RIfebd7b0_8276, \9114_9413 );
and \U$13695 ( \22525_22824 , RIe212bc8_4503, \9116_9415 );
and \U$13696 ( \22526_22825 , RIfebd648_8275, \9118_9417 );
and \U$13697 ( \22527_22826 , RIe20fec8_4471, \9120_9419 );
and \U$13698 ( \22528_22827 , RIfe7b900_7750, \9122_9421 );
and \U$13699 ( \22529_22828 , RIe20d1c8_4439, \9124_9423 );
and \U$13700 ( \22530_22829 , RIe20a4c8_4407, \9126_9425 );
and \U$13701 ( \22531_22830 , RIe2077c8_4375, \9128_9427 );
and \U$13702 ( \22532_22831 , RIf167258_5633, \9130_9429 );
and \U$13703 ( \22533_22832 , RIf166178_5621, \9132_9431 );
and \U$13704 ( \22534_22833 , RIe2024d0_4316, \9134_9433 );
and \U$13705 ( \22535_22834 , RIfe7bbd0_7752, \9136_9435 );
and \U$13706 ( \22536_22835 , RIf165368_5611, \9138_9437 );
and \U$13707 ( \22537_22836 , RIf1646c0_5602, \9140_9439 );
and \U$13708 ( \22538_22837 , RIfcd0a30_7396, \9142_9441 );
and \U$13709 ( \22539_22838 , RIf1620c8_5575, \9144_9443 );
and \U$13710 ( \22540_22839 , RIf1601d8_5553, \9146_9445 );
and \U$13711 ( \22541_22840 , RIf15e2e8_5531, \9148_9447 );
and \U$13712 ( \22542_22841 , RIfe7ba68_7751, \9150_9449 );
and \U$13713 ( \22543_22842 , RIfe7bea0_7754, \9152_9451 );
and \U$13714 ( \22544_22843 , RIf15cdd0_5516, \9154_9453 );
and \U$13715 ( \22545_22844 , RIf15b8b8_5501, \9156_9455 );
and \U$13716 ( \22546_22845 , RIf15a7d8_5489, \9158_9457 );
and \U$13717 ( \22547_22846 , RIfca4840_6894, \9160_9459 );
or \U$13718 ( \22548_22847 , \22484_22783 , \22485_22784 , \22486_22785 , \22487_22786 , \22488_22787 , \22489_22788 , \22490_22789 , \22491_22790 , \22492_22791 , \22493_22792 , \22494_22793 , \22495_22794 , \22496_22795 , \22497_22796 , \22498_22797 , \22499_22798 , \22500_22799 , \22501_22800 , \22502_22801 , \22503_22802 , \22504_22803 , \22505_22804 , \22506_22805 , \22507_22806 , \22508_22807 , \22509_22808 , \22510_22809 , \22511_22810 , \22512_22811 , \22513_22812 , \22514_22813 , \22515_22814 , \22516_22815 , \22517_22816 , \22518_22817 , \22519_22818 , \22520_22819 , \22521_22820 , \22522_22821 , \22523_22822 , \22524_22823 , \22525_22824 , \22526_22825 , \22527_22826 , \22528_22827 , \22529_22828 , \22530_22829 , \22531_22830 , \22532_22831 , \22533_22832 , \22534_22833 , \22535_22834 , \22536_22835 , \22537_22836 , \22538_22837 , \22539_22838 , \22540_22839 , \22541_22840 , \22542_22841 , \22543_22842 , \22544_22843 , \22545_22844 , \22546_22845 , \22547_22846 );
and \U$13719 ( \22549_22848 , RIf158ff0_5472, \9163_9462 );
and \U$13720 ( \22550_22849 , RIf157c40_5458, \9165_9464 );
and \U$13721 ( \22551_22850 , RIf156f98_5449, \9167_9466 );
and \U$13722 ( \22552_22851 , RIfe7c170_7756, \9169_9468 );
and \U$13723 ( \22553_22852 , RIf156458_5441, \9171_9470 );
and \U$13724 ( \22554_22853 , RIf155918_5433, \9173_9472 );
and \U$13725 ( \22555_22854 , RIf1549a0_5422, \9175_9474 );
and \U$13726 ( \22556_22855 , RIe1f54b0_4168, \9177_9476 );
and \U$13727 ( \22557_22856 , RIfe7c008_7755, \9179_9478 );
and \U$13728 ( \22558_22857 , RIf151b38_5389, \9181_9480 );
and \U$13729 ( \22559_22858 , RIf150bc0_5378, \9183_9482 );
and \U$13730 ( \22560_22859 , RIe1f32f0_4144, \9185_9484 );
and \U$13731 ( \22561_22860 , RIf14fae0_5366, \9187_9486 );
and \U$13732 ( \22562_22861 , RIf14ee38_5357, \9189_9488 );
and \U$13733 ( \22563_22862 , RIf14e028_5347, \9191_9490 );
and \U$13734 ( \22564_22863 , RIe1edff8_4085, \9193_9492 );
and \U$13735 ( \22565_22864 , RIe1eb730_4056, \9195_9494 );
and \U$13736 ( \22566_22865 , RIe1e8a30_4024, \9197_9496 );
and \U$13737 ( \22567_22866 , RIe1e5d30_3992, \9199_9498 );
and \U$13738 ( \22568_22867 , RIe1e3030_3960, \9201_9500 );
and \U$13739 ( \22569_22868 , RIe1e0330_3928, \9203_9502 );
and \U$13740 ( \22570_22869 , RIe1dd630_3896, \9205_9504 );
and \U$13741 ( \22571_22870 , RIe1da930_3864, \9207_9506 );
and \U$13742 ( \22572_22871 , RIe1d7c30_3832, \9209_9508 );
and \U$13743 ( \22573_22872 , RIe1d2230_3768, \9211_9510 );
and \U$13744 ( \22574_22873 , RIe1cf530_3736, \9213_9512 );
and \U$13745 ( \22575_22874 , RIe1cc830_3704, \9215_9514 );
and \U$13746 ( \22576_22875 , RIe1c9b30_3672, \9217_9516 );
and \U$13747 ( \22577_22876 , RIe1c6e30_3640, \9219_9518 );
and \U$13748 ( \22578_22877 , RIe1c4130_3608, \9221_9520 );
and \U$13749 ( \22579_22878 , RIe1c1430_3576, \9223_9522 );
and \U$13750 ( \22580_22879 , RIe1be730_3544, \9225_9524 );
and \U$13751 ( \22581_22880 , RIf14cb10_5332, \9227_9526 );
and \U$13752 ( \22582_22881 , RIf14b8c8_5319, \9229_9528 );
and \U$13753 ( \22583_22882 , RIfebda80_8278, \9231_9530 );
and \U$13754 ( \22584_22883 , RIfe7c878_7761, \9233_9532 );
and \U$13755 ( \22585_22884 , RIf14a680_5306, \9235_9534 );
and \U$13756 ( \22586_22885 , RIfe7c2d8_7757, \9237_9536 );
and \U$13757 ( \22587_22886 , RIfe7c9e0_7762, \9239_9538 );
and \U$13758 ( \22588_22887 , RIfe7c440_7758, \9241_9540 );
and \U$13759 ( \22589_22888 , RIf149000_5290, \9243_9542 );
and \U$13760 ( \22590_22889 , RIf147db8_5277, \9245_9544 );
and \U$13761 ( \22591_22890 , RIe1b2688_3407, \9247_9546 );
and \U$13762 ( \22592_22891 , RIfebd918_8277, \9249_9548 );
and \U$13763 ( \22593_22892 , RIfe7c5a8_7759, \9251_9550 );
and \U$13764 ( \22594_22893 , RIf146738_5261, \9253_9552 );
and \U$13765 ( \22595_22894 , RIfe7c710_7760, \9255_9554 );
and \U$13766 ( \22596_22895 , RIe1aad98_3321, \9257_9556 );
and \U$13767 ( \22597_22896 , RIe1a8a70_3296, \9259_9558 );
and \U$13768 ( \22598_22897 , RIe1a5d70_3264, \9261_9560 );
and \U$13769 ( \22599_22898 , RIe1a3070_3232, \9263_9562 );
and \U$13770 ( \22600_22899 , RIe1a0370_3200, \9265_9564 );
and \U$13771 ( \22601_22900 , RIe18c870_2976, \9267_9566 );
and \U$13772 ( \22602_22901 , RIe178d70_2752, \9269_9568 );
and \U$13773 ( \22603_22902 , RIe2266c8_4727, \9271_9570 );
and \U$13774 ( \22604_22903 , RIe21b2c8_4599, \9273_9572 );
and \U$13775 ( \22605_22904 , RIe204ac8_4343, \9275_9574 );
and \U$13776 ( \22606_22905 , RIe1feb28_4275, \9277_9576 );
and \U$13777 ( \22607_22906 , RIe1f7ee0_4198, \9279_9578 );
and \U$13778 ( \22608_22907 , RIe1f0a28_4115, \9281_9580 );
and \U$13779 ( \22609_22908 , RIe1d4f30_3800, \9283_9582 );
and \U$13780 ( \22610_22909 , RIe1bba30_3512, \9285_9584 );
and \U$13781 ( \22611_22910 , RIe1ae8a8_3363, \9287_9586 );
and \U$13782 ( \22612_22911 , RIe170ee0_2662, \9289_9588 );
or \U$13783 ( \22613_22912 , \22549_22848 , \22550_22849 , \22551_22850 , \22552_22851 , \22553_22852 , \22554_22853 , \22555_22854 , \22556_22855 , \22557_22856 , \22558_22857 , \22559_22858 , \22560_22859 , \22561_22860 , \22562_22861 , \22563_22862 , \22564_22863 , \22565_22864 , \22566_22865 , \22567_22866 , \22568_22867 , \22569_22868 , \22570_22869 , \22571_22870 , \22572_22871 , \22573_22872 , \22574_22873 , \22575_22874 , \22576_22875 , \22577_22876 , \22578_22877 , \22579_22878 , \22580_22879 , \22581_22880 , \22582_22881 , \22583_22882 , \22584_22883 , \22585_22884 , \22586_22885 , \22587_22886 , \22588_22887 , \22589_22888 , \22590_22889 , \22591_22890 , \22592_22891 , \22593_22892 , \22594_22893 , \22595_22894 , \22596_22895 , \22597_22896 , \22598_22897 , \22599_22898 , \22600_22899 , \22601_22900 , \22602_22901 , \22603_22902 , \22604_22903 , \22605_22904 , \22606_22905 , \22607_22906 , \22608_22907 , \22609_22908 , \22610_22909 , \22611_22910 , \22612_22911 );
or \U$13784 ( \22614_22913 , \22548_22847 , \22613_22912 );
_DC \g3894/U$1 ( \22615 , \22614_22913 , \9298_9597 );
buf \U$13785 ( \22616_22915 , \22615 );
xor \U$13786 ( \22617_22916 , \22483_22782 , \22616_22915 );
and \U$13787 ( \22618_22917 , RIdec5270_707, \8760_9059 );
and \U$13788 ( \22619_22918 , RIdec2570_675, \8762_9061 );
and \U$13789 ( \22620_22919 , RIee1ff18_4822, \8764_9063 );
and \U$13790 ( \22621_22920 , RIdebf870_643, \8766_9065 );
and \U$13791 ( \22622_22921 , RIfe7f848_7795, \8768_9067 );
and \U$13792 ( \22623_22922 , RIdebcb70_611, \8770_9069 );
and \U$13793 ( \22624_22923 , RIdeb9e70_579, \8772_9071 );
and \U$13794 ( \22625_22924 , RIdeb7170_547, \8774_9073 );
and \U$13795 ( \22626_22925 , RIfe7fc80_7798, \8776_9075 );
and \U$13796 ( \22627_22926 , RIdeb1770_483, \8778_9077 );
and \U$13797 ( \22628_22927 , RIfca5d58_6909, \8780_9079 );
and \U$13798 ( \22629_22928 , RIdeaea70_451, \8782_9081 );
and \U$13799 ( \22630_22929 , RIfcaf808_7019, \8784_9083 );
and \U$13800 ( \22631_22930 , RIdeaa0d8_419, \8786_9085 );
and \U$13801 ( \22632_22931 , RIdea37d8_387, \8788_9087 );
and \U$13802 ( \22633_22932 , RIde9ced8_355, \8790_9089 );
and \U$13803 ( \22634_22933 , RIfcdc3d0_7528, \8792_9091 );
and \U$13804 ( \22635_22934 , RIfcce438_7369, \8794_9093 );
and \U$13805 ( \22636_22935 , RIfcb0a50_7032, \8796_9095 );
and \U$13806 ( \22637_22936 , RIfc75680_6358, \8798_9097 );
and \U$13807 ( \22638_22937 , RIde90d40_296, \8800_9099 );
and \U$13808 ( \22639_22938 , RIfe7f9b0_7796, \8802_9101 );
and \U$13809 ( \22640_22939 , RIde89720_260, \8804_9103 );
and \U$13810 ( \22641_22940 , RIde85580_240, \8806_9105 );
and \U$13811 ( \22642_22941 , RIde81728_221, \8808_9107 );
and \U$13812 ( \22643_22942 , RIfc52f40_5966, \8810_9109 );
and \U$13813 ( \22644_22943 , RIfc82100_6502, \8812_9111 );
and \U$13814 ( \22645_22944 , RIfca7108_6923, \8814_9113 );
and \U$13815 ( \22646_22945 , RIfe7fb18_7797, \8816_9115 );
and \U$13816 ( \22647_22946 , RIe16b648_2599, \8818_9117 );
and \U$13817 ( \22648_22947 , RIe169a28_2579, \8820_9119 );
and \U$13818 ( \22649_22948 , RIe167ca0_2558, \8822_9121 );
and \U$13819 ( \22650_22949 , RIe165270_2528, \8824_9123 );
and \U$13820 ( \22651_22950 , RIe162570_2496, \8826_9125 );
and \U$13821 ( \22652_22951 , RIee37258_5086, \8828_9127 );
and \U$13822 ( \22653_22952 , RIe15f870_2464, \8830_9129 );
and \U$13823 ( \22654_22953 , RIee36178_5074, \8832_9131 );
and \U$13824 ( \22655_22954 , RIe15cb70_2432, \8834_9133 );
and \U$13825 ( \22656_22955 , RIe157170_2368, \8836_9135 );
and \U$13826 ( \22657_22956 , RIe154470_2336, \8838_9137 );
and \U$13827 ( \22658_22957 , RIfc86fc0_6558, \8840_9139 );
and \U$13828 ( \22659_22958 , RIe151770_2304, \8842_9141 );
and \U$13829 ( \22660_22959 , RIfc4eff8_5921, \8844_9143 );
and \U$13830 ( \22661_22960 , RIe14ea70_2272, \8846_9145 );
and \U$13831 ( \22662_22961 , RIfce1290_7584, \8848_9147 );
and \U$13832 ( \22663_22962 , RIe14bd70_2240, \8850_9149 );
and \U$13833 ( \22664_22963 , RIe149070_2208, \8852_9151 );
and \U$13834 ( \22665_22964 , RIe146370_2176, \8854_9153 );
and \U$13835 ( \22666_22965 , RIee34558_5054, \8856_9155 );
and \U$13836 ( \22667_22966 , RIee331a8_5040, \8858_9157 );
and \U$13837 ( \22668_22967 , RIee320c8_5028, \8860_9159 );
and \U$13838 ( \22669_22968 , RIee31150_5017, \8862_9161 );
and \U$13839 ( \22670_22969 , RIfe800b8_7801, \8864_9163 );
and \U$13840 ( \22671_22970 , RIfe7ff50_7800, \8866_9165 );
and \U$13841 ( \22672_22971 , RIdf3caf0_2067, \8868_9167 );
and \U$13842 ( \22673_22972 , RIfe7fde8_7799, \8870_9169 );
and \U$13843 ( \22674_22973 , RIfcc8330_7300, \8872_9171 );
and \U$13844 ( \22675_22974 , RIee2f800_4999, \8874_9173 );
and \U$13845 ( \22676_22975 , RIfca0d30_6852, \8876_9175 );
and \U$13846 ( \22677_22976 , RIee2d640_4975, \8878_9177 );
and \U$13847 ( \22678_22977 , RIdf35638_1984, \8880_9179 );
and \U$13848 ( \22679_22978 , RIdf331a8_1958, \8882_9181 );
and \U$13849 ( \22680_22979 , RIdf31150_1935, \8884_9183 );
and \U$13850 ( \22681_22980 , RIdf2ef90_1911, \8886_9185 );
or \U$13851 ( \22682_22981 , \22618_22917 , \22619_22918 , \22620_22919 , \22621_22920 , \22622_22921 , \22623_22922 , \22624_22923 , \22625_22924 , \22626_22925 , \22627_22926 , \22628_22927 , \22629_22928 , \22630_22929 , \22631_22930 , \22632_22931 , \22633_22932 , \22634_22933 , \22635_22934 , \22636_22935 , \22637_22936 , \22638_22937 , \22639_22938 , \22640_22939 , \22641_22940 , \22642_22941 , \22643_22942 , \22644_22943 , \22645_22944 , \22646_22945 , \22647_22946 , \22648_22947 , \22649_22948 , \22650_22949 , \22651_22950 , \22652_22951 , \22653_22952 , \22654_22953 , \22655_22954 , \22656_22955 , \22657_22956 , \22658_22957 , \22659_22958 , \22660_22959 , \22661_22960 , \22662_22961 , \22663_22962 , \22664_22963 , \22665_22964 , \22666_22965 , \22667_22966 , \22668_22967 , \22669_22968 , \22670_22969 , \22671_22970 , \22672_22971 , \22673_22972 , \22674_22973 , \22675_22974 , \22676_22975 , \22677_22976 , \22678_22977 , \22679_22978 , \22680_22979 , \22681_22980 );
and \U$13852 ( \22683_22982 , RIee2bb88_4956, \8889_9188 );
and \U$13853 ( \22684_22983 , RIee2a0d0_4937, \8891_9190 );
and \U$13854 ( \22685_22984 , RIee28d20_4923, \8893_9192 );
and \U$13855 ( \22686_22985 , RIfe7f578_7793, \8895_9194 );
and \U$13856 ( \22687_22986 , RIdf2a238_1856, \8897_9196 );
and \U$13857 ( \22688_22987 , RIdf27f10_1831, \8899_9198 );
and \U$13858 ( \22689_22988 , RIfe7f6e0_7794, \8901_9200 );
and \U$13859 ( \22690_22989 , RIdf246d0_1791, \8903_9202 );
and \U$13860 ( \22691_22990 , RIfcce9d8_7373, \8905_9204 );
and \U$13861 ( \22692_22991 , RIfc63638_6153, \8907_9206 );
and \U$13862 ( \22693_22992 , RIdf22c18_1772, \8909_9208 );
and \U$13863 ( \22694_22993 , RIfc62990_6144, \8911_9210 );
and \U$13864 ( \22695_22994 , RIdf21700_1757, \8913_9212 );
and \U$13865 ( \22696_22995 , RIdf1f810_1735, \8915_9214 );
and \U$13866 ( \22697_22996 , RIfeaa958_8257, \8917_9216 );
and \U$13867 ( \22698_22997 , RIdf19168_1662, \8919_9218 );
and \U$13868 ( \22699_22998 , RIdf16e40_1637, \8921_9220 );
and \U$13869 ( \22700_22999 , RIdf14140_1605, \8923_9222 );
and \U$13870 ( \22701_23000 , RIdf11440_1573, \8925_9224 );
and \U$13871 ( \22702_23001 , RIdf0e740_1541, \8927_9226 );
and \U$13872 ( \22703_23002 , RIdf0ba40_1509, \8929_9228 );
and \U$13873 ( \22704_23003 , RIdf08d40_1477, \8931_9230 );
and \U$13874 ( \22705_23004 , RIdf06040_1445, \8933_9232 );
and \U$13875 ( \22706_23005 , RIdf03340_1413, \8935_9234 );
and \U$13876 ( \22707_23006 , RIdefd940_1349, \8937_9236 );
and \U$13877 ( \22708_23007 , RIdefac40_1317, \8939_9238 );
and \U$13878 ( \22709_23008 , RIdef7f40_1285, \8941_9240 );
and \U$13879 ( \22710_23009 , RIdef5240_1253, \8943_9242 );
and \U$13880 ( \22711_23010 , RIdef2540_1221, \8945_9244 );
and \U$13881 ( \22712_23011 , RIdeef840_1189, \8947_9246 );
and \U$13882 ( \22713_23012 , RIdeecb40_1157, \8949_9248 );
and \U$13883 ( \22714_23013 , RIdee9e40_1125, \8951_9250 );
and \U$13884 ( \22715_23014 , RIfcb7800_7110, \8953_9252 );
and \U$13885 ( \22716_23015 , RIee24838_4874, \8955_9254 );
and \U$13886 ( \22717_23016 , RIfc4cb68_5895, \8957_9256 );
and \U$13887 ( \22718_23017 , RIee23320_4859, \8959_9258 );
and \U$13888 ( \22719_23018 , RIfe80388_7803, \8961_9260 );
and \U$13889 ( \22720_23019 , RIdee2c58_1044, \8963_9262 );
and \U$13890 ( \22721_23020 , RIfe80220_7802, \8965_9264 );
and \U$13891 ( \22722_23021 , RIdedea40_997, \8967_9266 );
and \U$13892 ( \22723_23022 , RIfc98900_6758, \8969_9268 );
and \U$13893 ( \22724_23023 , RIee223a8_4848, \8971_9270 );
and \U$13894 ( \22725_23024 , RIfcc8600_7302, \8973_9272 );
and \U$13895 ( \22726_23025 , RIee212c8_4836, \8975_9274 );
and \U$13896 ( \22727_23026 , RIded9748_938, \8977_9276 );
and \U$13897 ( \22728_23027 , RIfe804f0_7804, \8979_9278 );
and \U$13898 ( \22729_23028 , RIded53c8_890, \8981_9280 );
and \U$13899 ( \22730_23029 , RIded2c68_862, \8983_9282 );
and \U$13900 ( \22731_23030 , RIded0670_835, \8985_9284 );
and \U$13901 ( \22732_23031 , RIdecd970_803, \8987_9286 );
and \U$13902 ( \22733_23032 , RIdecac70_771, \8989_9288 );
and \U$13903 ( \22734_23033 , RIdec7f70_739, \8991_9290 );
and \U$13904 ( \22735_23034 , RIdeb4470_515, \8993_9292 );
and \U$13905 ( \22736_23035 , RIde965d8_323, \8995_9294 );
and \U$13906 ( \22737_23036 , RIe16e078_2629, \8997_9296 );
and \U$13907 ( \22738_23037 , RIe159e70_2400, \8999_9298 );
and \U$13908 ( \22739_23038 , RIe143670_2144, \9001_9300 );
and \U$13909 ( \22740_23039 , RIdf38068_2014, \9003_9302 );
and \U$13910 ( \22741_23040 , RIdf2c6c8_1882, \9005_9304 );
and \U$13911 ( \22742_23041 , RIdf1cf48_1706, \9007_9306 );
and \U$13912 ( \22743_23042 , RIdf00640_1381, \9009_9308 );
and \U$13913 ( \22744_23043 , RIdee7140_1093, \9011_9310 );
and \U$13914 ( \22745_23044 , RIdedbea8_966, \9013_9312 );
and \U$13915 ( \22746_23045 , RIde7c520_196, \9015_9314 );
or \U$13916 ( \22747_23046 , \22683_22982 , \22684_22983 , \22685_22984 , \22686_22985 , \22687_22986 , \22688_22987 , \22689_22988 , \22690_22989 , \22691_22990 , \22692_22991 , \22693_22992 , \22694_22993 , \22695_22994 , \22696_22995 , \22697_22996 , \22698_22997 , \22699_22998 , \22700_22999 , \22701_23000 , \22702_23001 , \22703_23002 , \22704_23003 , \22705_23004 , \22706_23005 , \22707_23006 , \22708_23007 , \22709_23008 , \22710_23009 , \22711_23010 , \22712_23011 , \22713_23012 , \22714_23013 , \22715_23014 , \22716_23015 , \22717_23016 , \22718_23017 , \22719_23018 , \22720_23019 , \22721_23020 , \22722_23021 , \22723_23022 , \22724_23023 , \22725_23024 , \22726_23025 , \22727_23026 , \22728_23027 , \22729_23028 , \22730_23029 , \22731_23030 , \22732_23031 , \22733_23032 , \22734_23033 , \22735_23034 , \22736_23035 , \22737_23036 , \22738_23037 , \22739_23038 , \22740_23039 , \22741_23040 , \22742_23041 , \22743_23042 , \22744_23043 , \22745_23044 , \22746_23045 );
or \U$13917 ( \22748_23047 , \22682_22981 , \22747_23046 );
_DC \g27ec/U$1 ( \22749 , \22748_23047 , \9024_9323 );
buf \U$13918 ( \22750_23049 , \22749 );
and \U$13919 ( \22751_23050 , RIe19d508_3167, \9034_9333 );
and \U$13920 ( \22752_23051 , RIe19a808_3135, \9036_9335 );
and \U$13921 ( \22753_23052 , RIfe7ee70_7788, \9038_9337 );
and \U$13922 ( \22754_23053 , RIe197b08_3103, \9040_9339 );
and \U$13923 ( \22755_23054 , RIfe7efd8_7789, \9042_9341 );
and \U$13924 ( \22756_23055 , RIe194e08_3071, \9044_9343 );
and \U$13925 ( \22757_23056 , RIe192108_3039, \9046_9345 );
and \U$13926 ( \22758_23057 , RIe18f408_3007, \9048_9347 );
and \U$13927 ( \22759_23058 , RIe189a08_2943, \9050_9349 );
and \U$13928 ( \22760_23059 , RIe186d08_2911, \9052_9351 );
and \U$13929 ( \22761_23060 , RIf143768_5227, \9054_9353 );
and \U$13930 ( \22762_23061 , RIe184008_2879, \9056_9355 );
and \U$13931 ( \22763_23062 , RIfc4bbf0_5884, \9058_9357 );
and \U$13932 ( \22764_23063 , RIe181308_2847, \9060_9359 );
and \U$13933 ( \22765_23064 , RIe17e608_2815, \9062_9361 );
and \U$13934 ( \22766_23065 , RIe17b908_2783, \9064_9363 );
and \U$13935 ( \22767_23066 , RIfe7f410_7792, \9066_9365 );
and \U$13936 ( \22768_23067 , RIf140d38_5197, \9068_9367 );
and \U$13937 ( \22769_23068 , RIe176fe8_2731, \9070_9369 );
and \U$13938 ( \22770_23069 , RIe175ad0_2716, \9072_9371 );
and \U$13939 ( \22771_23070 , RIfe7f2a8_7791, \9074_9373 );
and \U$13940 ( \22772_23071 , RIf13f118_5177, \9076_9375 );
and \U$13941 ( \22773_23072 , RIee3e440_5167, \9078_9377 );
and \U$13942 ( \22774_23073 , RIee3d360_5155, \9080_9379 );
and \U$13943 ( \22775_23074 , RIee3c280_5143, \9082_9381 );
and \U$13944 ( \22776_23075 , RIee3b1a0_5131, \9084_9383 );
and \U$13945 ( \22777_23076 , RIfe7f140_7790, \9086_9385 );
and \U$13946 ( \22778_23077 , RIe173640_2690, \9088_9387 );
and \U$13947 ( \22779_23078 , RIf170330_5736, \9090_9389 );
and \U$13948 ( \22780_23079 , RIf16f520_5726, \9092_9391 );
and \U$13949 ( \22781_23080 , RIf16e2d8_5713, \9094_9393 );
and \U$13950 ( \22782_23081 , RIf16d630_5704, \9096_9395 );
and \U$13951 ( \22783_23082 , RIfe7ea38_7785, \9098_9397 );
and \U$13952 ( \22784_23083 , RIe223860_4694, \9100_9399 );
and \U$13953 ( \22785_23084 , RIfc9c410_6800, \9102_9401 );
and \U$13954 ( \22786_23085 , RIe220b60_4662, \9104_9403 );
and \U$13955 ( \22787_23086 , RIfcb8340_7118, \9106_9405 );
and \U$13956 ( \22788_23087 , RIe21de60_4630, \9108_9407 );
and \U$13957 ( \22789_23088 , RIe218460_4566, \9110_9409 );
and \U$13958 ( \22790_23089 , RIe215760_4534, \9112_9411 );
and \U$13959 ( \22791_23090 , RIfc9cc80_6806, \9114_9413 );
and \U$13960 ( \22792_23091 , RIe212a60_4502, \9116_9415 );
and \U$13961 ( \22793_23092 , RIfc4ddb0_5908, \9118_9417 );
and \U$13962 ( \22794_23093 , RIe20fd60_4470, \9120_9419 );
and \U$13963 ( \22795_23094 , RIfc873f8_6561, \9122_9421 );
and \U$13964 ( \22796_23095 , RIe20d060_4438, \9124_9423 );
and \U$13965 ( \22797_23096 , RIe20a360_4406, \9126_9425 );
and \U$13966 ( \22798_23097 , RIe207660_4374, \9128_9427 );
and \U$13967 ( \22799_23098 , RIfc86750_6552, \9130_9429 );
and \U$13968 ( \22800_23099 , RIfc4e4b8_5913, \9132_9431 );
and \U$13969 ( \22801_23100 , RIe202368_4315, \9134_9433 );
and \U$13970 ( \22802_23101 , RIe200a18_4297, \9136_9435 );
and \U$13971 ( \22803_23102 , RIf165200_5610, \9138_9437 );
and \U$13972 ( \22804_23103 , RIf164558_5601, \9140_9439 );
and \U$13973 ( \22805_23104 , RIf163478_5589, \9142_9441 );
and \U$13974 ( \22806_23105 , RIf161f60_5574, \9144_9443 );
and \U$13975 ( \22807_23106 , RIf160070_5552, \9146_9445 );
and \U$13976 ( \22808_23107 , RIf15e180_5530, \9148_9447 );
and \U$13977 ( \22809_23108 , RIe1fcc38_4253, \9150_9449 );
and \U$13978 ( \22810_23109 , RIe1fb9f0_4240, \9152_9451 );
and \U$13979 ( \22811_23110 , RIf15cc68_5515, \9154_9453 );
and \U$13980 ( \22812_23111 , RIf15b750_5500, \9156_9455 );
and \U$13981 ( \22813_23112 , RIf15a670_5488, \9158_9457 );
and \U$13982 ( \22814_23113 , RIf159c98_5481, \9160_9459 );
or \U$13983 ( \22815_23114 , \22751_23050 , \22752_23051 , \22753_23052 , \22754_23053 , \22755_23054 , \22756_23055 , \22757_23056 , \22758_23057 , \22759_23058 , \22760_23059 , \22761_23060 , \22762_23061 , \22763_23062 , \22764_23063 , \22765_23064 , \22766_23065 , \22767_23066 , \22768_23067 , \22769_23068 , \22770_23069 , \22771_23070 , \22772_23071 , \22773_23072 , \22774_23073 , \22775_23074 , \22776_23075 , \22777_23076 , \22778_23077 , \22779_23078 , \22780_23079 , \22781_23080 , \22782_23081 , \22783_23082 , \22784_23083 , \22785_23084 , \22786_23085 , \22787_23086 , \22788_23087 , \22789_23088 , \22790_23089 , \22791_23090 , \22792_23091 , \22793_23092 , \22794_23093 , \22795_23094 , \22796_23095 , \22797_23096 , \22798_23097 , \22799_23098 , \22800_23099 , \22801_23100 , \22802_23101 , \22803_23102 , \22804_23103 , \22805_23104 , \22806_23105 , \22807_23106 , \22808_23107 , \22809_23108 , \22810_23109 , \22811_23110 , \22812_23111 , \22813_23112 , \22814_23113 );
and \U$13984 ( \22816_23115 , RIf158e88_5471, \9163_9462 );
and \U$13985 ( \22817_23116 , RIf157ad8_5457, \9165_9464 );
and \U$13986 ( \22818_23117 , RIf156e30_5448, \9167_9466 );
and \U$13987 ( \22819_23118 , RIfe7e768_7783, \9169_9468 );
and \U$13988 ( \22820_23119 , RIf1562f0_5440, \9171_9470 );
and \U$13989 ( \22821_23120 , RIf1557b0_5432, \9173_9472 );
and \U$13990 ( \22822_23121 , RIf154838_5421, \9175_9474 );
and \U$13991 ( \22823_23122 , RIfe7e8d0_7784, \9177_9476 );
and \U$13992 ( \22824_23123 , RIf1531b8_5405, \9179_9478 );
and \U$13993 ( \22825_23124 , RIfc52400_5958, \9181_9480 );
and \U$13994 ( \22826_23125 , RIf150a58_5377, \9183_9482 );
and \U$13995 ( \22827_23126 , RIe1f3188_4143, \9185_9484 );
and \U$13996 ( \22828_23127 , RIf14f978_5365, \9187_9486 );
and \U$13997 ( \22829_23128 , RIf14ecd0_5356, \9189_9488 );
and \U$13998 ( \22830_23129 , RIf14dec0_5346, \9191_9490 );
and \U$13999 ( \22831_23130 , RIe1ede90_4084, \9193_9492 );
and \U$14000 ( \22832_23131 , RIe1eb5c8_4055, \9195_9494 );
and \U$14001 ( \22833_23132 , RIe1e88c8_4023, \9197_9496 );
and \U$14002 ( \22834_23133 , RIe1e5bc8_3991, \9199_9498 );
and \U$14003 ( \22835_23134 , RIe1e2ec8_3959, \9201_9500 );
and \U$14004 ( \22836_23135 , RIe1e01c8_3927, \9203_9502 );
and \U$14005 ( \22837_23136 , RIe1dd4c8_3895, \9205_9504 );
and \U$14006 ( \22838_23137 , RIe1da7c8_3863, \9207_9506 );
and \U$14007 ( \22839_23138 , RIe1d7ac8_3831, \9209_9508 );
and \U$14008 ( \22840_23139 , RIe1d20c8_3767, \9211_9510 );
and \U$14009 ( \22841_23140 , RIe1cf3c8_3735, \9213_9512 );
and \U$14010 ( \22842_23141 , RIe1cc6c8_3703, \9215_9514 );
and \U$14011 ( \22843_23142 , RIe1c99c8_3671, \9217_9516 );
and \U$14012 ( \22844_23143 , RIe1c6cc8_3639, \9219_9518 );
and \U$14013 ( \22845_23144 , RIe1c3fc8_3607, \9221_9520 );
and \U$14014 ( \22846_23145 , RIe1c12c8_3575, \9223_9522 );
and \U$14015 ( \22847_23146 , RIe1be5c8_3543, \9225_9524 );
and \U$14016 ( \22848_23147 , RIf14c9a8_5331, \9227_9526 );
and \U$14017 ( \22849_23148 , RIf14b760_5318, \9229_9528 );
and \U$14018 ( \22850_23149 , RIfe7ed08_7787, \9231_9530 );
and \U$14019 ( \22851_23150 , RIfe7e600_7782, \9233_9532 );
and \U$14020 ( \22852_23151 , RIf14a518_5305, \9235_9534 );
and \U$14021 ( \22853_23152 , RIfca1f78_6865, \9237_9536 );
and \U$14022 ( \22854_23153 , RIfe7eba0_7786, \9239_9538 );
and \U$14023 ( \22855_23154 , RIfe7e498_7781, \9241_9540 );
and \U$14024 ( \22856_23155 , RIf148e98_5289, \9243_9542 );
and \U$14025 ( \22857_23156 , RIf147c50_5276, \9245_9544 );
and \U$14026 ( \22858_23157 , RIfe7e330_7780, \9247_9546 );
and \U$14027 ( \22859_23158 , RIe1b0a68_3387, \9249_9548 );
and \U$14028 ( \22860_23159 , RIf147278_5269, \9251_9550 );
and \U$14029 ( \22861_23160 , RIf1465d0_5260, \9253_9552 );
and \U$14030 ( \22862_23161 , RIe1ac418_3337, \9255_9554 );
and \U$14031 ( \22863_23162 , RIe1aac30_3320, \9257_9556 );
and \U$14032 ( \22864_23163 , RIe1a8908_3295, \9259_9558 );
and \U$14033 ( \22865_23164 , RIe1a5c08_3263, \9261_9560 );
and \U$14034 ( \22866_23165 , RIe1a2f08_3231, \9263_9562 );
and \U$14035 ( \22867_23166 , RIe1a0208_3199, \9265_9564 );
and \U$14036 ( \22868_23167 , RIe18c708_2975, \9267_9566 );
and \U$14037 ( \22869_23168 , RIe178c08_2751, \9269_9568 );
and \U$14038 ( \22870_23169 , RIe226560_4726, \9271_9570 );
and \U$14039 ( \22871_23170 , RIe21b160_4598, \9273_9572 );
and \U$14040 ( \22872_23171 , RIe204960_4342, \9275_9574 );
and \U$14041 ( \22873_23172 , RIe1fe9c0_4274, \9277_9576 );
and \U$14042 ( \22874_23173 , RIe1f7d78_4197, \9279_9578 );
and \U$14043 ( \22875_23174 , RIe1f08c0_4114, \9281_9580 );
and \U$14044 ( \22876_23175 , RIe1d4dc8_3799, \9283_9582 );
and \U$14045 ( \22877_23176 , RIe1bb8c8_3511, \9285_9584 );
and \U$14046 ( \22878_23177 , RIe1ae740_3362, \9287_9586 );
and \U$14047 ( \22879_23178 , RIe170d78_2661, \9289_9588 );
or \U$14048 ( \22880_23179 , \22816_23115 , \22817_23116 , \22818_23117 , \22819_23118 , \22820_23119 , \22821_23120 , \22822_23121 , \22823_23122 , \22824_23123 , \22825_23124 , \22826_23125 , \22827_23126 , \22828_23127 , \22829_23128 , \22830_23129 , \22831_23130 , \22832_23131 , \22833_23132 , \22834_23133 , \22835_23134 , \22836_23135 , \22837_23136 , \22838_23137 , \22839_23138 , \22840_23139 , \22841_23140 , \22842_23141 , \22843_23142 , \22844_23143 , \22845_23144 , \22846_23145 , \22847_23146 , \22848_23147 , \22849_23148 , \22850_23149 , \22851_23150 , \22852_23151 , \22853_23152 , \22854_23153 , \22855_23154 , \22856_23155 , \22857_23156 , \22858_23157 , \22859_23158 , \22860_23159 , \22861_23160 , \22862_23161 , \22863_23162 , \22864_23163 , \22865_23164 , \22866_23165 , \22867_23166 , \22868_23167 , \22869_23168 , \22870_23169 , \22871_23170 , \22872_23171 , \22873_23172 , \22874_23173 , \22875_23174 , \22876_23175 , \22877_23176 , \22878_23177 , \22879_23178 );
or \U$14049 ( \22881_23180 , \22815_23114 , \22880_23179 );
_DC \g3919/U$1 ( \22882 , \22881_23180 , \9298_9597 );
buf \U$14050 ( \22883_23182 , \22882 );
and \U$14051 ( \22884_23183 , \22750_23049 , \22883_23182 );
and \U$14052 ( \22885_23184 , \20940_21239 , \21073_21372 );
and \U$14053 ( \22886_23185 , \21073_21372 , \21348_21647 );
and \U$14054 ( \22887_23186 , \20940_21239 , \21348_21647 );
or \U$14055 ( \22888_23187 , \22885_23184 , \22886_23185 , \22887_23186 );
and \U$14056 ( \22889_23188 , \22883_23182 , \22888_23187 );
and \U$14057 ( \22890_23189 , \22750_23049 , \22888_23187 );
or \U$14058 ( \22891_23190 , \22884_23183 , \22889_23188 , \22890_23189 );
xor \U$14059 ( \22892_23191 , \22617_22916 , \22891_23190 );
buf g4418_GF_PartitionCandidate( \22893_23192_nG4418 , \22892_23191 );
xor \U$14060 ( \22894_23193 , \22750_23049 , \22883_23182 );
xor \U$14061 ( \22895_23194 , \22894_23193 , \22888_23187 );
buf g441b_GF_PartitionCandidate( \22896_23195_nG441b , \22895_23194 );
nand \U$14062 ( \22897_23196 , \22896_23195_nG441b , \21350_21649_nG441e );
and \U$14063 ( \22898_23197 , \22893_23192_nG4418 , \22897_23196 );
xor \U$14064 ( \22899_23198 , \22896_23195_nG441b , \21350_21649_nG441e );
and \U$14069 ( \22900_23202 , \22899_23198 , \10392_10694_nG9c0e );
or \U$14070 ( \22901_23203 , 1'b0 , \22900_23202 );
xor \U$14071 ( \22902_23204 , \22898_23197 , \22901_23203 );
xor \U$14072 ( \22903_23205 , \22898_23197 , \22902_23204 );
buf \U$14073 ( \22904_23206 , \22903_23205 );
buf \U$14074 ( \22905_23207 , \22904_23206 );
xor \U$14075 ( \22906_23208 , \22350_22649 , \22905_23207 );
and \U$14076 ( \22907_23209 , \21945_22244 , \22337_22636 );
and \U$14077 ( \22908_23210 , \21945_22244 , \22343_22642 );
and \U$14078 ( \22909_23211 , \22337_22636 , \22343_22642 );
or \U$14079 ( \22910_23212 , \22907_23209 , \22908_23210 , \22909_23211 );
and \U$14080 ( \22911_23213 , \22906_23208 , \22910_23212 );
and \U$14081 ( \22912_23214 , \21873_22175 , \21879_22181 );
and \U$14082 ( \22913_23215 , \21873_22175 , \21886_22188 );
and \U$14083 ( \22914_23216 , \21879_22181 , \21886_22188 );
or \U$14084 ( \22915_23217 , \22912_23214 , \22913_23215 , \22914_23216 );
buf \U$14085 ( \22916_23218 , \22915_23217 );
and \U$14086 ( \22917_23219 , \21894_22196 , \21934_22233 );
and \U$14087 ( \22918_23220 , \21894_22196 , \21941_22240 );
and \U$14088 ( \22919_23221 , \21934_22233 , \21941_22240 );
or \U$14089 ( \22920_23222 , \22917_23219 , \22918_23220 , \22919_23221 );
buf \U$14090 ( \22921_23223 , \22920_23222 );
and \U$14091 ( \22922_23224 , \12183_12157 , \19287_19586_nG9be1 );
and \U$14092 ( \22923_23225 , \11855_12154 , \20306_20608_nG9bde );
or \U$14093 ( \22924_23226 , \22922_23224 , \22923_23225 );
xor \U$14094 ( \22925_23227 , \11854_12153 , \22924_23226 );
buf \U$14095 ( \22926_23228 , \22925_23227 );
buf \U$14097 ( \22927_23229 , \22926_23228 );
xor \U$14098 ( \22928_23230 , \22921_23223 , \22927_23229 );
and \U$14099 ( \22929_23231 , \10996_10421 , \20787_21086_nG9bdb );
and \U$14100 ( \22930_23232 , \10119_10418 , \21827_22129_nG9bd8 );
or \U$14101 ( \22931_23233 , \22929_23231 , \22930_23232 );
xor \U$14102 ( \22932_23234 , \10118_10417 , \22931_23233 );
buf \U$14103 ( \22933_23235 , \22932_23234 );
buf \U$14105 ( \22934_23236 , \22933_23235 );
xor \U$14106 ( \22935_23237 , \22928_23230 , \22934_23236 );
buf \U$14107 ( \22936_23238 , \22935_23237 );
xor \U$14108 ( \22937_23239 , \22916_23218 , \22936_23238 );
and \U$14109 ( \22938_23240 , \21950_22249 , \21955_22254 );
and \U$14110 ( \22939_23241 , \21950_22249 , \22335_22634 );
and \U$14111 ( \22940_23242 , \21955_22254 , \22335_22634 );
or \U$14112 ( \22941_23243 , \22938_23240 , \22939_23241 , \22940_23242 );
buf \U$14113 ( \22942_23244 , \22941_23243 );
xor \U$14114 ( \22943_23245 , \22937_23239 , \22942_23244 );
buf \U$14115 ( \22944_23246 , \22943_23245 );
and \U$14116 ( \22945_23247 , \21853_22155 , \21888_22190 );
and \U$14117 ( \22946_23248 , \21853_22155 , \21943_22242 );
and \U$14118 ( \22947_23249 , \21888_22190 , \21943_22242 );
or \U$14119 ( \22948_23250 , \22945_23247 , \22946_23248 , \22947_23249 );
buf \U$14120 ( \22949_23251 , \22948_23250 );
xor \U$14121 ( \22950_23252 , \22944_23246 , \22949_23251 );
and \U$14122 ( \22951_23253 , \21858_22160 , \21864_22166 );
and \U$14123 ( \22952_23254 , \21858_22160 , \21871_22173 );
and \U$14124 ( \22953_23255 , \21864_22166 , \21871_22173 );
or \U$14125 ( \22954_23256 , \22951_23253 , \22952_23254 , \22953_23255 );
buf \U$14126 ( \22955_23257 , \22954_23256 );
and \U$14127 ( \22956_23258 , \21905_22207 , \21914_22213 );
and \U$14128 ( \22957_23259 , \21905_22207 , \21921_22220 );
and \U$14129 ( \22958_23260 , \21914_22213 , \21921_22220 );
or \U$14130 ( \22959_23261 , \22956_23258 , \22957_23259 , \22958_23260 );
buf \U$14131 ( \22960_23262 , \22959_23261 );
and \U$14132 ( \22961_23263 , \21908_21658 , \10693_10995_nG9c0b );
and \U$14133 ( \22962_23264 , \21356_21655 , \10981_11283_nG9c08 );
or \U$14134 ( \22963_23265 , \22961_23263 , \22962_23264 );
xor \U$14135 ( \22964_23266 , \21355_21654 , \22963_23265 );
buf \U$14136 ( \22965_23267 , \22964_23266 );
buf \U$14138 ( \22966_23268 , \22965_23267 );
and \U$14139 ( \22967_23269 , \20353_20155 , \11299_11598_nG9c05 );
and \U$14140 ( \22968_23270 , \19853_20152 , \12168_12470_nG9c02 );
or \U$14141 ( \22969_23271 , \22967_23269 , \22968_23270 );
xor \U$14142 ( \22970_23272 , \19852_20151 , \22969_23271 );
buf \U$14143 ( \22971_23273 , \22970_23272 );
buf \U$14145 ( \22972_23274 , \22971_23273 );
xor \U$14146 ( \22973_23275 , \22966_23268 , \22972_23274 );
buf \U$14147 ( \22974_23276 , \22973_23275 );
xor \U$14148 ( \22975_23277 , \22960_23262 , \22974_23276 );
and \U$14149 ( \22976_23278 , \16405_15940 , \15074_15373_nG9bf3 );
and \U$14150 ( \22977_23279 , \15638_15937 , \16013_16315_nG9bf0 );
or \U$14151 ( \22978_23280 , \22976_23278 , \22977_23279 );
xor \U$14152 ( \22979_23281 , \15637_15936 , \22978_23280 );
buf \U$14153 ( \22980_23282 , \22979_23281 );
buf \U$14155 ( \22981_23283 , \22980_23282 );
xor \U$14156 ( \22982_23284 , \22975_23277 , \22981_23283 );
buf \U$14157 ( \22983_23285 , \22982_23284 );
xor \U$14158 ( \22984_23286 , \22955_23257 , \22983_23285 );
and \U$14159 ( \22985_23287 , \21923_22222 , \21925_22224 );
and \U$14160 ( \22986_23288 , \21923_22222 , \21932_22231 );
and \U$14161 ( \22987_23289 , \21925_22224 , \21932_22231 );
or \U$14162 ( \22988_23290 , \22985_23287 , \22986_23288 , \22987_23289 );
buf \U$14163 ( \22989_23291 , \22988_23290 );
xor \U$14164 ( \22990_23292 , \22984_23286 , \22989_23291 );
buf \U$14165 ( \22991_23293 , \22990_23292 );
and \U$14166 ( \22992_23294 , \21897_22199 , \21903_22205 );
buf \U$14167 ( \22993_23295 , \22992_23294 );
and \U$14168 ( \22994_23296 , \18908_18702 , \12502_12801_nG9bff );
and \U$14169 ( \22995_23297 , \18400_18699 , \13403_13705_nG9bfc );
or \U$14170 ( \22996_23298 , \22994_23296 , \22995_23297 );
xor \U$14171 ( \22997_23299 , \18399_18698 , \22996_23298 );
buf \U$14172 ( \22998_23300 , \22997_23299 );
buf \U$14174 ( \22999_23301 , \22998_23300 );
xor \U$14175 ( \23000_23302 , \22993_23295 , \22999_23301 );
and \U$14176 ( \23001_23303 , \17437_17297 , \13771_14070_nG9bf9 );
and \U$14177 ( \23002_23304 , \16995_17294 , \14682_14984_nG9bf6 );
or \U$14178 ( \23003_23305 , \23001_23303 , \23002_23304 );
xor \U$14179 ( \23004_23306 , \16994_17293 , \23003_23305 );
buf \U$14180 ( \23005_23307 , \23004_23306 );
buf \U$14182 ( \23006_23308 , \23005_23307 );
xor \U$14183 ( \23007_23309 , \23000_23302 , \23006_23308 );
buf \U$14184 ( \23008_23310 , \23007_23309 );
and \U$14185 ( \23009_23311 , \14710_14631 , \16378_16680_nG9bed );
and \U$14186 ( \23010_23312 , \14329_14628 , \17363_17665_nG9bea );
or \U$14187 ( \23011_23313 , \23009_23311 , \23010_23312 );
xor \U$14188 ( \23012_23314 , \14328_14627 , \23011_23313 );
buf \U$14189 ( \23013_23315 , \23012_23314 );
buf \U$14191 ( \23014_23316 , \23013_23315 );
xor \U$14192 ( \23015_23317 , \23008_23310 , \23014_23316 );
and \U$14193 ( \23016_23318 , \13431_13370 , \17808_18107_nG9be7 );
and \U$14194 ( \23017_23319 , \13068_13367 , \18789_19091_nG9be4 );
or \U$14195 ( \23018_23320 , \23016_23318 , \23017_23319 );
xor \U$14196 ( \23019_23321 , \13067_13366 , \23018_23320 );
buf \U$14197 ( \23020_23322 , \23019_23321 );
buf \U$14199 ( \23021_23323 , \23020_23322 );
xor \U$14200 ( \23022_23324 , \23015_23317 , \23021_23323 );
buf \U$14201 ( \23023_23325 , \23022_23324 );
xor \U$14202 ( \23024_23326 , \22991_23293 , \23023_23325 );
and \U$14203 ( \23025_23327 , \10411_10707 , \22330_22629_nG9bd5 );
and \U$14204 ( \23026_23328 , \21965_22264 , \22251_22550 );
and \U$14205 ( \23027_23329 , \22251_22550 , \22273_22572 );
and \U$14206 ( \23028_23330 , \21965_22264 , \22273_22572 );
or \U$14207 ( \23029_23331 , \23026_23328 , \23027_23329 , \23028_23330 );
and \U$14208 ( \23030_23332 , \22279_22578 , \22283_22582 );
and \U$14209 ( \23031_23333 , \22283_22582 , \22318_22617 );
and \U$14210 ( \23032_23334 , \22279_22578 , \22318_22617 );
or \U$14211 ( \23033_23335 , \23030_23332 , \23031_23333 , \23032_23334 );
xor \U$14212 ( \23034_23336 , \23029_23331 , \23033_23335 );
and \U$14213 ( \23035_23337 , \21969_22268 , \21973_22272 );
and \U$14214 ( \23036_23338 , \21973_22272 , \22250_22549 );
and \U$14215 ( \23037_23339 , \21969_22268 , \22250_22549 );
or \U$14216 ( \23038_23340 , \23035_23337 , \23036_23338 , \23037_23339 );
and \U$14217 ( \23039_23341 , \22292_22591 , \22296_22595 );
and \U$14218 ( \23040_23342 , \22296_22595 , \22301_22600 );
and \U$14219 ( \23041_23343 , \22292_22591 , \22301_22600 );
or \U$14220 ( \23042_23344 , \23039_23341 , \23040_23342 , \23041_23343 );
xor \U$14221 ( \23043_23345 , \23038_23340 , \23042_23344 );
and \U$14222 ( \23044_23346 , \22307_22606 , \22311_22610 );
and \U$14223 ( \23045_23347 , \22311_22610 , \22316_22615 );
and \U$14224 ( \23046_23348 , \22307_22606 , \22316_22615 );
or \U$14225 ( \23047_23349 , \23044_23346 , \23045_23347 , \23046_23348 );
xor \U$14226 ( \23048_23350 , \23043_23345 , \23047_23349 );
and \U$14227 ( \23049_23351 , \22257_22556 , \10681_10983 );
and \U$14228 ( \23050_23352 , RIdec5270_707, \9034_9333 );
and \U$14229 ( \23051_23353 , RIdec2570_675, \9036_9335 );
and \U$14230 ( \23052_23354 , RIee1ff18_4822, \9038_9337 );
and \U$14231 ( \23053_23355 , RIdebf870_643, \9040_9339 );
and \U$14232 ( \23054_23356 , RIfe7f848_7795, \9042_9341 );
and \U$14233 ( \23055_23357 , RIdebcb70_611, \9044_9343 );
and \U$14234 ( \23056_23358 , RIdeb9e70_579, \9046_9345 );
and \U$14235 ( \23057_23359 , RIdeb7170_547, \9048_9347 );
and \U$14236 ( \23058_23360 , RIfe7fc80_7798, \9050_9349 );
and \U$14237 ( \23059_23361 , RIdeb1770_483, \9052_9351 );
and \U$14238 ( \23060_23362 , RIfca5d58_6909, \9054_9353 );
and \U$14239 ( \23061_23363 , RIdeaea70_451, \9056_9355 );
and \U$14240 ( \23062_23364 , RIfcaf808_7019, \9058_9357 );
and \U$14241 ( \23063_23365 , RIdeaa0d8_419, \9060_9359 );
and \U$14242 ( \23064_23366 , RIdea37d8_387, \9062_9361 );
and \U$14243 ( \23065_23367 , RIde9ced8_355, \9064_9363 );
and \U$14244 ( \23066_23368 , RIfcdc3d0_7528, \9066_9365 );
and \U$14245 ( \23067_23369 , RIfcce438_7369, \9068_9367 );
and \U$14246 ( \23068_23370 , RIfcb0a50_7032, \9070_9369 );
and \U$14247 ( \23069_23371 , RIfc75680_6358, \9072_9371 );
and \U$14248 ( \23070_23372 , RIde90d40_296, \9074_9373 );
and \U$14249 ( \23071_23373 , RIfe7f9b0_7796, \9076_9375 );
and \U$14250 ( \23072_23374 , RIde89720_260, \9078_9377 );
and \U$14251 ( \23073_23375 , RIde85580_240, \9080_9379 );
and \U$14252 ( \23074_23376 , RIde81728_221, \9082_9381 );
and \U$14253 ( \23075_23377 , RIfc52f40_5966, \9084_9383 );
and \U$14254 ( \23076_23378 , RIfc82100_6502, \9086_9385 );
and \U$14255 ( \23077_23379 , RIfca7108_6923, \9088_9387 );
and \U$14256 ( \23078_23380 , RIfe7fb18_7797, \9090_9389 );
and \U$14257 ( \23079_23381 , RIe16b648_2599, \9092_9391 );
and \U$14258 ( \23080_23382 , RIe169a28_2579, \9094_9393 );
and \U$14259 ( \23081_23383 , RIe167ca0_2558, \9096_9395 );
and \U$14260 ( \23082_23384 , RIe165270_2528, \9098_9397 );
and \U$14261 ( \23083_23385 , RIe162570_2496, \9100_9399 );
and \U$14262 ( \23084_23386 , RIee37258_5086, \9102_9401 );
and \U$14263 ( \23085_23387 , RIe15f870_2464, \9104_9403 );
and \U$14264 ( \23086_23388 , RIee36178_5074, \9106_9405 );
and \U$14265 ( \23087_23389 , RIe15cb70_2432, \9108_9407 );
and \U$14266 ( \23088_23390 , RIe157170_2368, \9110_9409 );
and \U$14267 ( \23089_23391 , RIe154470_2336, \9112_9411 );
and \U$14268 ( \23090_23392 , RIfc86fc0_6558, \9114_9413 );
and \U$14269 ( \23091_23393 , RIe151770_2304, \9116_9415 );
and \U$14270 ( \23092_23394 , RIfc4eff8_5921, \9118_9417 );
and \U$14271 ( \23093_23395 , RIe14ea70_2272, \9120_9419 );
and \U$14272 ( \23094_23396 , RIfce1290_7584, \9122_9421 );
and \U$14273 ( \23095_23397 , RIe14bd70_2240, \9124_9423 );
and \U$14274 ( \23096_23398 , RIe149070_2208, \9126_9425 );
and \U$14275 ( \23097_23399 , RIe146370_2176, \9128_9427 );
and \U$14276 ( \23098_23400 , RIee34558_5054, \9130_9429 );
and \U$14277 ( \23099_23401 , RIee331a8_5040, \9132_9431 );
and \U$14278 ( \23100_23402 , RIee320c8_5028, \9134_9433 );
and \U$14279 ( \23101_23403 , RIee31150_5017, \9136_9435 );
and \U$14280 ( \23102_23404 , RIfe800b8_7801, \9138_9437 );
and \U$14281 ( \23103_23405 , RIfe7ff50_7800, \9140_9439 );
and \U$14282 ( \23104_23406 , RIdf3caf0_2067, \9142_9441 );
and \U$14283 ( \23105_23407 , RIfe7fde8_7799, \9144_9443 );
and \U$14284 ( \23106_23408 , RIfcc8330_7300, \9146_9445 );
and \U$14285 ( \23107_23409 , RIee2f800_4999, \9148_9447 );
and \U$14286 ( \23108_23410 , RIfca0d30_6852, \9150_9449 );
and \U$14287 ( \23109_23411 , RIee2d640_4975, \9152_9451 );
and \U$14288 ( \23110_23412 , RIdf35638_1984, \9154_9453 );
and \U$14289 ( \23111_23413 , RIdf331a8_1958, \9156_9455 );
and \U$14290 ( \23112_23414 , RIdf31150_1935, \9158_9457 );
and \U$14291 ( \23113_23415 , RIdf2ef90_1911, \9160_9459 );
or \U$14292 ( \23114_23416 , \23050_23352 , \23051_23353 , \23052_23354 , \23053_23355 , \23054_23356 , \23055_23357 , \23056_23358 , \23057_23359 , \23058_23360 , \23059_23361 , \23060_23362 , \23061_23363 , \23062_23364 , \23063_23365 , \23064_23366 , \23065_23367 , \23066_23368 , \23067_23369 , \23068_23370 , \23069_23371 , \23070_23372 , \23071_23373 , \23072_23374 , \23073_23375 , \23074_23376 , \23075_23377 , \23076_23378 , \23077_23379 , \23078_23380 , \23079_23381 , \23080_23382 , \23081_23383 , \23082_23384 , \23083_23385 , \23084_23386 , \23085_23387 , \23086_23388 , \23087_23389 , \23088_23390 , \23089_23391 , \23090_23392 , \23091_23393 , \23092_23394 , \23093_23395 , \23094_23396 , \23095_23397 , \23096_23398 , \23097_23399 , \23098_23400 , \23099_23401 , \23100_23402 , \23101_23403 , \23102_23404 , \23103_23405 , \23104_23406 , \23105_23407 , \23106_23408 , \23107_23409 , \23108_23410 , \23109_23411 , \23110_23412 , \23111_23413 , \23112_23414 , \23113_23415 );
and \U$14293 ( \23115_23417 , RIee2bb88_4956, \9163_9462 );
and \U$14294 ( \23116_23418 , RIee2a0d0_4937, \9165_9464 );
and \U$14295 ( \23117_23419 , RIee28d20_4923, \9167_9466 );
and \U$14296 ( \23118_23420 , RIfe7f578_7793, \9169_9468 );
and \U$14297 ( \23119_23421 , RIdf2a238_1856, \9171_9470 );
and \U$14298 ( \23120_23422 , RIdf27f10_1831, \9173_9472 );
and \U$14299 ( \23121_23423 , RIfe7f6e0_7794, \9175_9474 );
and \U$14300 ( \23122_23424 , RIdf246d0_1791, \9177_9476 );
and \U$14301 ( \23123_23425 , RIfcce9d8_7373, \9179_9478 );
and \U$14302 ( \23124_23426 , RIfc63638_6153, \9181_9480 );
and \U$14303 ( \23125_23427 , RIdf22c18_1772, \9183_9482 );
and \U$14304 ( \23126_23428 , RIfc62990_6144, \9185_9484 );
and \U$14305 ( \23127_23429 , RIdf21700_1757, \9187_9486 );
and \U$14306 ( \23128_23430 , RIdf1f810_1735, \9189_9488 );
and \U$14307 ( \23129_23431 , RIfeaa958_8257, \9191_9490 );
and \U$14308 ( \23130_23432 , RIdf19168_1662, \9193_9492 );
and \U$14309 ( \23131_23433 , RIdf16e40_1637, \9195_9494 );
and \U$14310 ( \23132_23434 , RIdf14140_1605, \9197_9496 );
and \U$14311 ( \23133_23435 , RIdf11440_1573, \9199_9498 );
and \U$14312 ( \23134_23436 , RIdf0e740_1541, \9201_9500 );
and \U$14313 ( \23135_23437 , RIdf0ba40_1509, \9203_9502 );
and \U$14314 ( \23136_23438 , RIdf08d40_1477, \9205_9504 );
and \U$14315 ( \23137_23439 , RIdf06040_1445, \9207_9506 );
and \U$14316 ( \23138_23440 , RIdf03340_1413, \9209_9508 );
and \U$14317 ( \23139_23441 , RIdefd940_1349, \9211_9510 );
and \U$14318 ( \23140_23442 , RIdefac40_1317, \9213_9512 );
and \U$14319 ( \23141_23443 , RIdef7f40_1285, \9215_9514 );
and \U$14320 ( \23142_23444 , RIdef5240_1253, \9217_9516 );
and \U$14321 ( \23143_23445 , RIdef2540_1221, \9219_9518 );
and \U$14322 ( \23144_23446 , RIdeef840_1189, \9221_9520 );
and \U$14323 ( \23145_23447 , RIdeecb40_1157, \9223_9522 );
and \U$14324 ( \23146_23448 , RIdee9e40_1125, \9225_9524 );
and \U$14325 ( \23147_23449 , RIfcb7800_7110, \9227_9526 );
and \U$14326 ( \23148_23450 , RIee24838_4874, \9229_9528 );
and \U$14327 ( \23149_23451 , RIfc4cb68_5895, \9231_9530 );
and \U$14328 ( \23150_23452 , RIee23320_4859, \9233_9532 );
and \U$14329 ( \23151_23453 , RIfe80388_7803, \9235_9534 );
and \U$14330 ( \23152_23454 , RIdee2c58_1044, \9237_9536 );
and \U$14331 ( \23153_23455 , RIfe80220_7802, \9239_9538 );
and \U$14332 ( \23154_23456 , RIdedea40_997, \9241_9540 );
and \U$14333 ( \23155_23457 , RIfc98900_6758, \9243_9542 );
and \U$14334 ( \23156_23458 , RIee223a8_4848, \9245_9544 );
and \U$14335 ( \23157_23459 , RIfcc8600_7302, \9247_9546 );
and \U$14336 ( \23158_23460 , RIee212c8_4836, \9249_9548 );
and \U$14337 ( \23159_23461 , RIded9748_938, \9251_9550 );
and \U$14338 ( \23160_23462 , RIfe804f0_7804, \9253_9552 );
and \U$14339 ( \23161_23463 , RIded53c8_890, \9255_9554 );
and \U$14340 ( \23162_23464 , RIded2c68_862, \9257_9556 );
and \U$14341 ( \23163_23465 , RIded0670_835, \9259_9558 );
and \U$14342 ( \23164_23466 , RIdecd970_803, \9261_9560 );
and \U$14343 ( \23165_23467 , RIdecac70_771, \9263_9562 );
and \U$14344 ( \23166_23468 , RIdec7f70_739, \9265_9564 );
and \U$14345 ( \23167_23469 , RIdeb4470_515, \9267_9566 );
and \U$14346 ( \23168_23470 , RIde965d8_323, \9269_9568 );
and \U$14347 ( \23169_23471 , RIe16e078_2629, \9271_9570 );
and \U$14348 ( \23170_23472 , RIe159e70_2400, \9273_9572 );
and \U$14349 ( \23171_23473 , RIe143670_2144, \9275_9574 );
and \U$14350 ( \23172_23474 , RIdf38068_2014, \9277_9576 );
and \U$14351 ( \23173_23475 , RIdf2c6c8_1882, \9279_9578 );
and \U$14352 ( \23174_23476 , RIdf1cf48_1706, \9281_9580 );
and \U$14353 ( \23175_23477 , RIdf00640_1381, \9283_9582 );
and \U$14354 ( \23176_23478 , RIdee7140_1093, \9285_9584 );
and \U$14355 ( \23177_23479 , RIdedbea8_966, \9287_9586 );
and \U$14356 ( \23178_23480 , RIde7c520_196, \9289_9588 );
or \U$14357 ( \23179_23481 , \23115_23417 , \23116_23418 , \23117_23419 , \23118_23420 , \23119_23421 , \23120_23422 , \23121_23423 , \23122_23424 , \23123_23425 , \23124_23426 , \23125_23427 , \23126_23428 , \23127_23429 , \23128_23430 , \23129_23431 , \23130_23432 , \23131_23433 , \23132_23434 , \23133_23435 , \23134_23436 , \23135_23437 , \23136_23438 , \23137_23439 , \23138_23440 , \23139_23441 , \23140_23442 , \23141_23443 , \23142_23444 , \23143_23445 , \23144_23446 , \23145_23447 , \23146_23448 , \23147_23449 , \23148_23450 , \23149_23451 , \23150_23452 , \23151_23453 , \23152_23454 , \23153_23455 , \23154_23456 , \23155_23457 , \23156_23458 , \23157_23459 , \23158_23460 , \23159_23461 , \23160_23462 , \23161_23463 , \23162_23464 , \23163_23465 , \23164_23466 , \23165_23467 , \23166_23468 , \23167_23469 , \23168_23470 , \23169_23471 , \23170_23472 , \23171_23473 , \23172_23474 , \23173_23475 , \23174_23476 , \23175_23477 , \23176_23478 , \23177_23479 , \23178_23480 );
or \U$14358 ( \23180_23482 , \23114_23416 , \23179_23481 );
_DC \g65b3/U$1 ( \23181 , \23180_23482 , \9298_9597 );
and \U$14359 ( \23182_23484 , RIe19d508_3167, \8760_9059 );
and \U$14360 ( \23183_23485 , RIe19a808_3135, \8762_9061 );
and \U$14361 ( \23184_23486 , RIfe7ee70_7788, \8764_9063 );
and \U$14362 ( \23185_23487 , RIe197b08_3103, \8766_9065 );
and \U$14363 ( \23186_23488 , RIfe7efd8_7789, \8768_9067 );
and \U$14364 ( \23187_23489 , RIe194e08_3071, \8770_9069 );
and \U$14365 ( \23188_23490 , RIe192108_3039, \8772_9071 );
and \U$14366 ( \23189_23491 , RIe18f408_3007, \8774_9073 );
and \U$14367 ( \23190_23492 , RIe189a08_2943, \8776_9075 );
and \U$14368 ( \23191_23493 , RIe186d08_2911, \8778_9077 );
and \U$14369 ( \23192_23494 , RIf143768_5227, \8780_9079 );
and \U$14370 ( \23193_23495 , RIe184008_2879, \8782_9081 );
and \U$14371 ( \23194_23496 , RIfc4bbf0_5884, \8784_9083 );
and \U$14372 ( \23195_23497 , RIe181308_2847, \8786_9085 );
and \U$14373 ( \23196_23498 , RIe17e608_2815, \8788_9087 );
and \U$14374 ( \23197_23499 , RIe17b908_2783, \8790_9089 );
and \U$14375 ( \23198_23500 , RIfe7f410_7792, \8792_9091 );
and \U$14376 ( \23199_23501 , RIf140d38_5197, \8794_9093 );
and \U$14377 ( \23200_23502 , RIe176fe8_2731, \8796_9095 );
and \U$14378 ( \23201_23503 , RIe175ad0_2716, \8798_9097 );
and \U$14379 ( \23202_23504 , RIfe7f2a8_7791, \8800_9099 );
and \U$14380 ( \23203_23505 , RIf13f118_5177, \8802_9101 );
and \U$14381 ( \23204_23506 , RIee3e440_5167, \8804_9103 );
and \U$14382 ( \23205_23507 , RIee3d360_5155, \8806_9105 );
and \U$14383 ( \23206_23508 , RIee3c280_5143, \8808_9107 );
and \U$14384 ( \23207_23509 , RIee3b1a0_5131, \8810_9109 );
and \U$14385 ( \23208_23510 , RIfe7f140_7790, \8812_9111 );
and \U$14386 ( \23209_23511 , RIe173640_2690, \8814_9113 );
and \U$14387 ( \23210_23512 , RIf170330_5736, \8816_9115 );
and \U$14388 ( \23211_23513 , RIf16f520_5726, \8818_9117 );
and \U$14389 ( \23212_23514 , RIf16e2d8_5713, \8820_9119 );
and \U$14390 ( \23213_23515 , RIf16d630_5704, \8822_9121 );
and \U$14391 ( \23214_23516 , RIfe7ea38_7785, \8824_9123 );
and \U$14392 ( \23215_23517 , RIe223860_4694, \8826_9125 );
and \U$14393 ( \23216_23518 , RIfc9c410_6800, \8828_9127 );
and \U$14394 ( \23217_23519 , RIe220b60_4662, \8830_9129 );
and \U$14395 ( \23218_23520 , RIfcb8340_7118, \8832_9131 );
and \U$14396 ( \23219_23521 , RIe21de60_4630, \8834_9133 );
and \U$14397 ( \23220_23522 , RIe218460_4566, \8836_9135 );
and \U$14398 ( \23221_23523 , RIe215760_4534, \8838_9137 );
and \U$14399 ( \23222_23524 , RIfc9cc80_6806, \8840_9139 );
and \U$14400 ( \23223_23525 , RIe212a60_4502, \8842_9141 );
and \U$14401 ( \23224_23526 , RIfc4ddb0_5908, \8844_9143 );
and \U$14402 ( \23225_23527 , RIe20fd60_4470, \8846_9145 );
and \U$14403 ( \23226_23528 , RIfc873f8_6561, \8848_9147 );
and \U$14404 ( \23227_23529 , RIe20d060_4438, \8850_9149 );
and \U$14405 ( \23228_23530 , RIe20a360_4406, \8852_9151 );
and \U$14406 ( \23229_23531 , RIe207660_4374, \8854_9153 );
and \U$14407 ( \23230_23532 , RIfc86750_6552, \8856_9155 );
and \U$14408 ( \23231_23533 , RIfc4e4b8_5913, \8858_9157 );
and \U$14409 ( \23232_23534 , RIe202368_4315, \8860_9159 );
and \U$14410 ( \23233_23535 , RIe200a18_4297, \8862_9161 );
and \U$14411 ( \23234_23536 , RIf165200_5610, \8864_9163 );
and \U$14412 ( \23235_23537 , RIf164558_5601, \8866_9165 );
and \U$14413 ( \23236_23538 , RIf163478_5589, \8868_9167 );
and \U$14414 ( \23237_23539 , RIf161f60_5574, \8870_9169 );
and \U$14415 ( \23238_23540 , RIf160070_5552, \8872_9171 );
and \U$14416 ( \23239_23541 , RIf15e180_5530, \8874_9173 );
and \U$14417 ( \23240_23542 , RIe1fcc38_4253, \8876_9175 );
and \U$14418 ( \23241_23543 , RIe1fb9f0_4240, \8878_9177 );
and \U$14419 ( \23242_23544 , RIf15cc68_5515, \8880_9179 );
and \U$14420 ( \23243_23545 , RIf15b750_5500, \8882_9181 );
and \U$14421 ( \23244_23546 , RIf15a670_5488, \8884_9183 );
and \U$14422 ( \23245_23547 , RIf159c98_5481, \8886_9185 );
or \U$14423 ( \23246_23548 , \23182_23484 , \23183_23485 , \23184_23486 , \23185_23487 , \23186_23488 , \23187_23489 , \23188_23490 , \23189_23491 , \23190_23492 , \23191_23493 , \23192_23494 , \23193_23495 , \23194_23496 , \23195_23497 , \23196_23498 , \23197_23499 , \23198_23500 , \23199_23501 , \23200_23502 , \23201_23503 , \23202_23504 , \23203_23505 , \23204_23506 , \23205_23507 , \23206_23508 , \23207_23509 , \23208_23510 , \23209_23511 , \23210_23512 , \23211_23513 , \23212_23514 , \23213_23515 , \23214_23516 , \23215_23517 , \23216_23518 , \23217_23519 , \23218_23520 , \23219_23521 , \23220_23522 , \23221_23523 , \23222_23524 , \23223_23525 , \23224_23526 , \23225_23527 , \23226_23528 , \23227_23529 , \23228_23530 , \23229_23531 , \23230_23532 , \23231_23533 , \23232_23534 , \23233_23535 , \23234_23536 , \23235_23537 , \23236_23538 , \23237_23539 , \23238_23540 , \23239_23541 , \23240_23542 , \23241_23543 , \23242_23544 , \23243_23545 , \23244_23546 , \23245_23547 );
and \U$14424 ( \23247_23549 , RIf158e88_5471, \8889_9188 );
and \U$14425 ( \23248_23550 , RIf157ad8_5457, \8891_9190 );
and \U$14426 ( \23249_23551 , RIf156e30_5448, \8893_9192 );
and \U$14427 ( \23250_23552 , RIfe7e768_7783, \8895_9194 );
and \U$14428 ( \23251_23553 , RIf1562f0_5440, \8897_9196 );
and \U$14429 ( \23252_23554 , RIf1557b0_5432, \8899_9198 );
and \U$14430 ( \23253_23555 , RIf154838_5421, \8901_9200 );
and \U$14431 ( \23254_23556 , RIfe7e8d0_7784, \8903_9202 );
and \U$14432 ( \23255_23557 , RIf1531b8_5405, \8905_9204 );
and \U$14433 ( \23256_23558 , RIfc52400_5958, \8907_9206 );
and \U$14434 ( \23257_23559 , RIf150a58_5377, \8909_9208 );
and \U$14435 ( \23258_23560 , RIe1f3188_4143, \8911_9210 );
and \U$14436 ( \23259_23561 , RIf14f978_5365, \8913_9212 );
and \U$14437 ( \23260_23562 , RIf14ecd0_5356, \8915_9214 );
and \U$14438 ( \23261_23563 , RIf14dec0_5346, \8917_9216 );
and \U$14439 ( \23262_23564 , RIe1ede90_4084, \8919_9218 );
and \U$14440 ( \23263_23565 , RIe1eb5c8_4055, \8921_9220 );
and \U$14441 ( \23264_23566 , RIe1e88c8_4023, \8923_9222 );
and \U$14442 ( \23265_23567 , RIe1e5bc8_3991, \8925_9224 );
and \U$14443 ( \23266_23568 , RIe1e2ec8_3959, \8927_9226 );
and \U$14444 ( \23267_23569 , RIe1e01c8_3927, \8929_9228 );
and \U$14445 ( \23268_23570 , RIe1dd4c8_3895, \8931_9230 );
and \U$14446 ( \23269_23571 , RIe1da7c8_3863, \8933_9232 );
and \U$14447 ( \23270_23572 , RIe1d7ac8_3831, \8935_9234 );
and \U$14448 ( \23271_23573 , RIe1d20c8_3767, \8937_9236 );
and \U$14449 ( \23272_23574 , RIe1cf3c8_3735, \8939_9238 );
and \U$14450 ( \23273_23575 , RIe1cc6c8_3703, \8941_9240 );
and \U$14451 ( \23274_23576 , RIe1c99c8_3671, \8943_9242 );
and \U$14452 ( \23275_23577 , RIe1c6cc8_3639, \8945_9244 );
and \U$14453 ( \23276_23578 , RIe1c3fc8_3607, \8947_9246 );
and \U$14454 ( \23277_23579 , RIe1c12c8_3575, \8949_9248 );
and \U$14455 ( \23278_23580 , RIe1be5c8_3543, \8951_9250 );
and \U$14456 ( \23279_23581 , RIf14c9a8_5331, \8953_9252 );
and \U$14457 ( \23280_23582 , RIf14b760_5318, \8955_9254 );
and \U$14458 ( \23281_23583 , RIfe7ed08_7787, \8957_9256 );
and \U$14459 ( \23282_23584 , RIfe7e600_7782, \8959_9258 );
and \U$14460 ( \23283_23585 , RIf14a518_5305, \8961_9260 );
and \U$14461 ( \23284_23586 , RIfca1f78_6865, \8963_9262 );
and \U$14462 ( \23285_23587 , RIfe7eba0_7786, \8965_9264 );
and \U$14463 ( \23286_23588 , RIfe7e498_7781, \8967_9266 );
and \U$14464 ( \23287_23589 , RIf148e98_5289, \8969_9268 );
and \U$14465 ( \23288_23590 , RIf147c50_5276, \8971_9270 );
and \U$14466 ( \23289_23591 , RIfe7e330_7780, \8973_9272 );
and \U$14467 ( \23290_23592 , RIe1b0a68_3387, \8975_9274 );
and \U$14468 ( \23291_23593 , RIf147278_5269, \8977_9276 );
and \U$14469 ( \23292_23594 , RIf1465d0_5260, \8979_9278 );
and \U$14470 ( \23293_23595 , RIe1ac418_3337, \8981_9280 );
and \U$14471 ( \23294_23596 , RIe1aac30_3320, \8983_9282 );
and \U$14472 ( \23295_23597 , RIe1a8908_3295, \8985_9284 );
and \U$14473 ( \23296_23598 , RIe1a5c08_3263, \8987_9286 );
and \U$14474 ( \23297_23599 , RIe1a2f08_3231, \8989_9288 );
and \U$14475 ( \23298_23600 , RIe1a0208_3199, \8991_9290 );
and \U$14476 ( \23299_23601 , RIe18c708_2975, \8993_9292 );
and \U$14477 ( \23300_23602 , RIe178c08_2751, \8995_9294 );
and \U$14478 ( \23301_23603 , RIe226560_4726, \8997_9296 );
and \U$14479 ( \23302_23604 , RIe21b160_4598, \8999_9298 );
and \U$14480 ( \23303_23605 , RIe204960_4342, \9001_9300 );
and \U$14481 ( \23304_23606 , RIe1fe9c0_4274, \9003_9302 );
and \U$14482 ( \23305_23607 , RIe1f7d78_4197, \9005_9304 );
and \U$14483 ( \23306_23608 , RIe1f08c0_4114, \9007_9306 );
and \U$14484 ( \23307_23609 , RIe1d4dc8_3799, \9009_9308 );
and \U$14485 ( \23308_23610 , RIe1bb8c8_3511, \9011_9310 );
and \U$14486 ( \23309_23611 , RIe1ae740_3362, \9013_9312 );
and \U$14487 ( \23310_23612 , RIe170d78_2661, \9015_9314 );
or \U$14488 ( \23311_23613 , \23247_23549 , \23248_23550 , \23249_23551 , \23250_23552 , \23251_23553 , \23252_23554 , \23253_23555 , \23254_23556 , \23255_23557 , \23256_23558 , \23257_23559 , \23258_23560 , \23259_23561 , \23260_23562 , \23261_23563 , \23262_23564 , \23263_23565 , \23264_23566 , \23265_23567 , \23266_23568 , \23267_23569 , \23268_23570 , \23269_23571 , \23270_23572 , \23271_23573 , \23272_23574 , \23273_23575 , \23274_23576 , \23275_23577 , \23276_23578 , \23277_23579 , \23278_23580 , \23279_23581 , \23280_23582 , \23281_23583 , \23282_23584 , \23283_23585 , \23284_23586 , \23285_23587 , \23286_23588 , \23287_23589 , \23288_23590 , \23289_23591 , \23290_23592 , \23291_23593 , \23292_23594 , \23293_23595 , \23294_23596 , \23295_23597 , \23296_23598 , \23297_23599 , \23298_23600 , \23299_23601 , \23300_23602 , \23301_23603 , \23302_23604 , \23303_23605 , \23304_23606 , \23305_23607 , \23306_23608 , \23307_23609 , \23308_23610 , \23309_23611 , \23310_23612 );
or \U$14489 ( \23312_23614 , \23246_23548 , \23311_23613 );
_DC \g65b4/U$1 ( \23313 , \23312_23614 , \9024_9323 );
and g65b5_GF_PartitionCandidate( \23314_23616_nG65b5 , \23181 , \23313 );
buf \U$14490 ( \23315_23617 , \23314_23616_nG65b5 );
and \U$14491 ( \23316_23618 , \23315_23617 , \10389_10691 );
nor \U$14492 ( \23317_23619 , \23049_23351 , \23316_23618 );
xnor \U$14493 ( \23318_23620 , \23317_23619 , \10678_10980 );
and \U$14494 ( \23319_23621 , \17736_18035 , \13755_14054 );
and \U$14495 ( \23320_23622 , \18730_19032 , \13390_13692 );
nor \U$14496 ( \23321_23623 , \23319_23621 , \23320_23622 );
xnor \U$14497 ( \23322_23624 , \23321_23623 , \13736_14035 );
xor \U$14498 ( \23323_23625 , \23318_23620 , \23322_23624 );
_DC \g598e/U$1 ( \23324 , \23180_23482 , \9298_9597 );
_DC \g5a12/U$1 ( \23325 , \23312_23614 , \9024_9323 );
xor g5a13_GF_PartitionCandidate( \23326_23628_nG5a13 , \23324 , \23325 );
buf \U$14499 ( \23327_23629 , \23326_23628_nG5a13 );
xor \U$14500 ( \23328_23630 , \23327_23629 , \22240_22539 );
and \U$14501 ( \23329_23631 , \10385_10687 , \23328_23630 );
xor \U$14502 ( \23330_23632 , \23323_23625 , \23329_23631 );
and \U$14503 ( \23331_23633 , \19259_19558 , \12491_12790 );
and \U$14504 ( \23332_23634 , \20242_20544 , \12159_12461 );
nor \U$14505 ( \23333_23635 , \23331_23633 , \23332_23634 );
xnor \U$14506 ( \23334_23636 , \23333_23635 , \12481_12780 );
and \U$14507 ( \23335_23637 , \16353_16655 , \15037_15336 );
and \U$14508 ( \23336_23638 , \17325_17627 , \14661_14963 );
nor \U$14509 ( \23337_23639 , \23335_23637 , \23336_23638 );
xnor \U$14510 ( \23338_23640 , \23337_23639 , \15043_15342 );
xor \U$14511 ( \23339_23641 , \23334_23636 , \23338_23640 );
and \U$14512 ( \23340_23642 , \10686_10988 , \22243_22542 );
and \U$14513 ( \23341_23643 , \10968_11270 , \21801_22103 );
nor \U$14514 ( \23342_23644 , \23340_23642 , \23341_23643 );
xnor \U$14515 ( \23343_23645 , \23342_23644 , \22249_22548 );
xor \U$14516 ( \23344_23646 , \23339_23641 , \23343_23645 );
xor \U$14517 ( \23345_23647 , \23330_23632 , \23344_23646 );
and \U$14518 ( \23346_23648 , \20734_21033 , \11275_11574 );
and \U$14519 ( \23347_23649 , \21788_22090 , \10976_11278 );
nor \U$14520 ( \23348_23650 , \23346_23648 , \23347_23649 );
xnor \U$14521 ( \23349_23651 , \23348_23650 , \11281_11580 );
and \U$14522 ( \23350_23652 , \12470_12769 , \19235_19534 );
and \U$14523 ( \23351_23653 , \13377_13679 , \18743_19045 );
nor \U$14524 ( \23352_23654 , \23350_23652 , \23351_23653 );
xnor \U$14525 ( \23353_23655 , \23352_23654 , \19241_19540 );
xor \U$14526 ( \23354_23656 , \23349_23651 , \23353_23655 );
and \U$14527 ( \23355_23657 , \11287_11586 , \20706_21005 );
and \U$14528 ( \23356_23658 , \12146_12448 , \20255_20557 );
nor \U$14529 ( \23357_23659 , \23355_23657 , \23356_23658 );
xnor \U$14530 ( \23358_23660 , \23357_23659 , \20712_21011 );
xor \U$14531 ( \23359_23661 , \23354_23656 , \23358_23660 );
xor \U$14532 ( \23360_23662 , \23345_23647 , \23359_23661 );
xor \U$14533 ( \23361_23663 , \23048_23350 , \23360_23662 );
and \U$14534 ( \23362_23664 , \22263_22562 , \22267_22566 );
and \U$14535 ( \23363_23665 , \22267_22566 , \22272_22571 );
and \U$14536 ( \23364_23666 , \22263_22562 , \22272_22571 );
or \U$14537 ( \23365_23667 , \23362_23664 , \23363_23665 , \23364_23666 );
and \U$14538 ( \23366_23668 , \22288_22587 , \22302_22601 );
and \U$14539 ( \23367_23669 , \22302_22601 , \22317_22616 );
and \U$14540 ( \23368_23670 , \22288_22587 , \22317_22616 );
or \U$14541 ( \23369_23671 , \23366_23668 , \23367_23669 , \23368_23670 );
xor \U$14542 ( \23370_23672 , \23365_23667 , \23369_23671 );
and \U$14543 ( \23371_23673 , \22260_22559 , \22262_22561 );
and \U$14544 ( \23372_23674 , \15022_15321 , \16333_16635 );
and \U$14545 ( \23373_23675 , \15965_16267 , \15999_16301 );
nor \U$14546 ( \23374_23676 , \23372_23674 , \23373_23675 );
xnor \U$14547 ( \23375_23677 , \23374_23676 , \16323_16625 );
xor \U$14548 ( \23376_23678 , \23371_23673 , \23375_23677 );
and \U$14549 ( \23377_23679 , \13725_14024 , \17791_18090 );
and \U$14550 ( \23378_23680 , \14648_14950 , \17353_17655 );
nor \U$14551 ( \23379_23681 , \23377_23679 , \23378_23680 );
xnor \U$14552 ( \23380_23682 , \23379_23681 , \17747_18046 );
xor \U$14553 ( \23381_23683 , \23376_23678 , \23380_23682 );
xor \U$14554 ( \23382_23684 , \23370_23672 , \23381_23683 );
xor \U$14555 ( \23383_23685 , \23361_23663 , \23382_23684 );
xor \U$14556 ( \23384_23686 , \23034_23336 , \23383_23685 );
and \U$14557 ( \23385_23687 , \21961_22260 , \22274_22573 );
and \U$14558 ( \23386_23688 , \22274_22573 , \22319_22618 );
and \U$14559 ( \23387_23689 , \21961_22260 , \22319_22618 );
or \U$14560 ( \23388_23690 , \23385_23687 , \23386_23688 , \23387_23689 );
xor \U$14561 ( \23389_23691 , \23384_23686 , \23388_23690 );
and \U$14562 ( \23390_23692 , \22320_22619 , \22324_22623 );
and \U$14563 ( \23391_23693 , \22325_22624 , \22328_22627 );
or \U$14564 ( \23392_23694 , \23390_23692 , \23391_23693 );
xor \U$14565 ( \23393_23695 , \23389_23691 , \23392_23694 );
buf g9bd2_GF_PartitionCandidate( \23394_23696_nG9bd2 , \23393_23695 );
and \U$14566 ( \23395_23697 , \10402_10704 , \23394_23696_nG9bd2 );
or \U$14567 ( \23396_23698 , \23025_23327 , \23395_23697 );
xor \U$14568 ( \23397_23699 , \10399_10703 , \23396_23698 );
buf \U$14569 ( \23398_23700 , \23397_23699 );
buf \U$14571 ( \23399_23701 , \23398_23700 );
xor \U$14572 ( \23400_23702 , \23024_23326 , \23399_23701 );
buf \U$14573 ( \23401_23703 , \23400_23702 );
xor \U$14574 ( \23402_23704 , \22950_23252 , \23401_23703 );
and \U$14575 ( \23403_23705 , \22906_23208 , \23402_23704 );
and \U$14576 ( \23404_23706 , \22910_23212 , \23402_23704 );
or \U$14577 ( \23405_23707 , \22911_23213 , \23403_23705 , \23404_23706 );
and \U$14578 ( \23406_23708 , \22345_22644 , \22349_22648 );
and \U$14579 ( \23407_23709 , \22345_22644 , \22905_23207 );
and \U$14580 ( \23408_23710 , \22349_22648 , \22905_23207 );
or \U$14581 ( \23409_23711 , \23406_23708 , \23407_23709 , \23408_23710 );
xor \U$14582 ( \23410_23712 , \23405_23707 , \23409_23711 );
and \U$14583 ( \23411_23713 , \22944_23246 , \22949_23251 );
and \U$14584 ( \23412_23714 , \22944_23246 , \23401_23703 );
and \U$14585 ( \23413_23715 , \22949_23251 , \23401_23703 );
or \U$14586 ( \23414_23716 , \23411_23713 , \23412_23714 , \23413_23715 );
xor \U$14587 ( \23415_23717 , \23410_23712 , \23414_23716 );
and \U$14588 ( \23416_23718 , \23008_23310 , \23014_23316 );
and \U$14589 ( \23417_23719 , \23008_23310 , \23021_23323 );
and \U$14590 ( \23418_23720 , \23014_23316 , \23021_23323 );
or \U$14591 ( \23419_23721 , \23416_23718 , \23417_23719 , \23418_23720 );
buf \U$14592 ( \23420_23722 , \23419_23721 );
and \U$14593 ( \23421_23723 , \22955_23257 , \22983_23285 );
and \U$14594 ( \23422_23724 , \22955_23257 , \22989_23291 );
and \U$14595 ( \23423_23725 , \22983_23285 , \22989_23291 );
or \U$14596 ( \23424_23726 , \23421_23723 , \23422_23724 , \23423_23725 );
buf \U$14597 ( \23425_23727 , \23424_23726 );
xor \U$14598 ( \23426_23728 , \23420_23722 , \23425_23727 );
and \U$14599 ( \23427_23729 , \10996_10421 , \21827_22129_nG9bd8 );
and \U$14600 ( \23428_23730 , \10119_10418 , \22330_22629_nG9bd5 );
or \U$14601 ( \23429_23731 , \23427_23729 , \23428_23730 );
xor \U$14602 ( \23430_23732 , \10118_10417 , \23429_23731 );
buf \U$14603 ( \23431_23733 , \23430_23732 );
buf \U$14605 ( \23432_23734 , \23431_23733 );
xor \U$14606 ( \23433_23735 , \23426_23728 , \23432_23734 );
buf \U$14607 ( \23434_23736 , \23433_23735 );
and \U$14608 ( \23435_23737 , \22991_23293 , \23023_23325 );
and \U$14609 ( \23436_23738 , \22991_23293 , \23399_23701 );
and \U$14610 ( \23437_23739 , \23023_23325 , \23399_23701 );
or \U$14611 ( \23438_23740 , \23435_23737 , \23436_23738 , \23437_23739 );
buf \U$14612 ( \23439_23741 , \23438_23740 );
xor \U$14613 ( \23440_23742 , \23434_23736 , \23439_23741 );
and \U$14614 ( \23441_23743 , \22921_23223 , \22927_23229 );
and \U$14615 ( \23442_23744 , \22921_23223 , \22934_23236 );
and \U$14616 ( \23443_23745 , \22927_23229 , \22934_23236 );
or \U$14617 ( \23444_23746 , \23441_23743 , \23442_23744 , \23443_23745 );
buf \U$14618 ( \23445_23747 , \23444_23746 );
xor \U$14619 ( \23446_23748 , \23440_23742 , \23445_23747 );
buf \U$14620 ( \23447_23749 , \23446_23748 );
and \U$14621 ( \23448_23750 , \22916_23218 , \22936_23238 );
and \U$14622 ( \23449_23751 , \22916_23218 , \22942_23244 );
and \U$14623 ( \23450_23752 , \22936_23238 , \22942_23244 );
or \U$14624 ( \23451_23753 , \23448_23750 , \23449_23751 , \23450_23752 );
buf \U$14625 ( \23452_23754 , \23451_23753 );
xor \U$14626 ( \23453_23755 , \23447_23749 , \23452_23754 );
and \U$14627 ( \23454_23756 , \22960_23262 , \22974_23276 );
and \U$14628 ( \23455_23757 , \22960_23262 , \22981_23283 );
and \U$14629 ( \23456_23758 , \22974_23276 , \22981_23283 );
or \U$14630 ( \23457_23759 , \23454_23756 , \23455_23757 , \23456_23758 );
buf \U$14631 ( \23458_23760 , \23457_23759 );
and \U$14632 ( \23459_23761 , \22966_23268 , \22972_23274 );
buf \U$14633 ( \23460_23762 , \23459_23761 );
and \U$14634 ( \23461_23763 , \18908_18702 , \13403_13705_nG9bfc );
and \U$14635 ( \23462_23764 , \18400_18699 , \13771_14070_nG9bf9 );
or \U$14636 ( \23463_23765 , \23461_23763 , \23462_23764 );
xor \U$14637 ( \23464_23766 , \18399_18698 , \23463_23765 );
buf \U$14638 ( \23465_23767 , \23464_23766 );
buf \U$14640 ( \23466_23768 , \23465_23767 );
xor \U$14641 ( \23467_23769 , \23460_23762 , \23466_23768 );
and \U$14642 ( \23468_23770 , \17437_17297 , \14682_14984_nG9bf6 );
and \U$14643 ( \23469_23771 , \16995_17294 , \15074_15373_nG9bf3 );
or \U$14644 ( \23470_23772 , \23468_23770 , \23469_23771 );
xor \U$14645 ( \23471_23773 , \16994_17293 , \23470_23772 );
buf \U$14646 ( \23472_23774 , \23471_23773 );
buf \U$14648 ( \23473_23775 , \23472_23774 );
xor \U$14649 ( \23474_23776 , \23467_23769 , \23473_23775 );
buf \U$14650 ( \23475_23777 , \23474_23776 );
xor \U$14651 ( \23476_23778 , \23458_23760 , \23475_23777 );
and \U$14652 ( \23477_23779 , \14710_14631 , \17363_17665_nG9bea );
and \U$14653 ( \23478_23780 , \14329_14628 , \17808_18107_nG9be7 );
or \U$14654 ( \23479_23781 , \23477_23779 , \23478_23780 );
xor \U$14655 ( \23480_23782 , \14328_14627 , \23479_23781 );
buf \U$14656 ( \23481_23783 , \23480_23782 );
buf \U$14658 ( \23482_23784 , \23481_23783 );
xor \U$14659 ( \23483_23785 , \23476_23778 , \23482_23784 );
buf \U$14660 ( \23484_23786 , \23483_23785 );
and \U$14661 ( \23485_23787 , \22993_23295 , \22999_23301 );
and \U$14662 ( \23486_23788 , \22993_23295 , \23006_23308 );
and \U$14663 ( \23487_23789 , \22999_23301 , \23006_23308 );
or \U$14664 ( \23488_23790 , \23485_23787 , \23486_23788 , \23487_23789 );
buf \U$14665 ( \23489_23791 , \23488_23790 );
and \U$14666 ( \23490_23792 , \22898_23197 , \22902_23204 );
buf \U$14667 ( \23491_23793 , \23490_23792 );
buf \U$14669 ( \23492_23794 , \23491_23793 );
not \U$14065 ( \23493_23199 , \22899_23198 );
xor \U$14066 ( \23494_23200 , \22893_23192_nG4418 , \22896_23195_nG441b );
and \U$14067 ( \23495_23201 , \23493_23199 , \23494_23200 );
and \U$14670 ( \23496_23795 , \23495_23201 , \10392_10694_nG9c0e );
and \U$14671 ( \23497_23796 , \22899_23198 , \10693_10995_nG9c0b );
or \U$14672 ( \23498_23797 , \23496_23795 , \23497_23796 );
xor \U$14673 ( \23499_23798 , \22898_23197 , \23498_23797 );
buf \U$14674 ( \23500_23799 , \23499_23798 );
buf \U$14676 ( \23501_23800 , \23500_23799 );
xor \U$14677 ( \23502_23801 , \23492_23794 , \23501_23800 );
buf \U$14678 ( \23503_23802 , \23502_23801 );
and \U$14679 ( \23504_23803 , \21908_21658 , \10981_11283_nG9c08 );
and \U$14680 ( \23505_23804 , \21356_21655 , \11299_11598_nG9c05 );
or \U$14681 ( \23506_23805 , \23504_23803 , \23505_23804 );
xor \U$14682 ( \23507_23806 , \21355_21654 , \23506_23805 );
buf \U$14683 ( \23508_23807 , \23507_23806 );
buf \U$14685 ( \23509_23808 , \23508_23807 );
xor \U$14686 ( \23510_23809 , \23503_23802 , \23509_23808 );
and \U$14687 ( \23511_23810 , \20353_20155 , \12168_12470_nG9c02 );
and \U$14688 ( \23512_23811 , \19853_20152 , \12502_12801_nG9bff );
or \U$14689 ( \23513_23812 , \23511_23810 , \23512_23811 );
xor \U$14690 ( \23514_23813 , \19852_20151 , \23513_23812 );
buf \U$14691 ( \23515_23814 , \23514_23813 );
buf \U$14693 ( \23516_23815 , \23515_23814 );
xor \U$14694 ( \23517_23816 , \23510_23809 , \23516_23815 );
buf \U$14695 ( \23518_23817 , \23517_23816 );
xor \U$14696 ( \23519_23818 , \23489_23791 , \23518_23817 );
and \U$14697 ( \23520_23819 , \16405_15940 , \16013_16315_nG9bf0 );
and \U$14698 ( \23521_23820 , \15638_15937 , \16378_16680_nG9bed );
or \U$14699 ( \23522_23821 , \23520_23819 , \23521_23820 );
xor \U$14700 ( \23523_23822 , \15637_15936 , \23522_23821 );
buf \U$14701 ( \23524_23823 , \23523_23822 );
buf \U$14703 ( \23525_23824 , \23524_23823 );
xor \U$14704 ( \23526_23825 , \23519_23818 , \23525_23824 );
buf \U$14705 ( \23527_23826 , \23526_23825 );
and \U$14706 ( \23528_23827 , \13431_13370 , \18789_19091_nG9be4 );
and \U$14707 ( \23529_23828 , \13068_13367 , \19287_19586_nG9be1 );
or \U$14708 ( \23530_23829 , \23528_23827 , \23529_23828 );
xor \U$14709 ( \23531_23830 , \13067_13366 , \23530_23829 );
buf \U$14710 ( \23532_23831 , \23531_23830 );
buf \U$14712 ( \23533_23832 , \23532_23831 );
xor \U$14713 ( \23534_23833 , \23527_23826 , \23533_23832 );
and \U$14714 ( \23535_23834 , \12183_12157 , \20306_20608_nG9bde );
and \U$14715 ( \23536_23835 , \11855_12154 , \20787_21086_nG9bdb );
or \U$14716 ( \23537_23836 , \23535_23834 , \23536_23835 );
xor \U$14717 ( \23538_23837 , \11854_12153 , \23537_23836 );
buf \U$14718 ( \23539_23838 , \23538_23837 );
buf \U$14720 ( \23540_23839 , \23539_23838 );
xor \U$14721 ( \23541_23840 , \23534_23833 , \23540_23839 );
buf \U$14722 ( \23542_23841 , \23541_23840 );
xor \U$14723 ( \23543_23842 , \23484_23786 , \23542_23841 );
and \U$14724 ( \23544_23843 , \10411_10707 , \23394_23696_nG9bd2 );
and \U$14725 ( \23545_23844 , \23365_23667 , \23369_23671 );
and \U$14726 ( \23546_23845 , \23369_23671 , \23381_23683 );
and \U$14727 ( \23547_23846 , \23365_23667 , \23381_23683 );
or \U$14728 ( \23548_23847 , \23545_23844 , \23546_23845 , \23547_23846 );
and \U$14729 ( \23549_23848 , \23048_23350 , \23360_23662 );
and \U$14730 ( \23550_23849 , \23360_23662 , \23382_23684 );
and \U$14731 ( \23551_23850 , \23048_23350 , \23382_23684 );
or \U$14732 ( \23552_23851 , \23549_23848 , \23550_23849 , \23551_23850 );
xor \U$14733 ( \23553_23852 , \23548_23847 , \23552_23851 );
and \U$14734 ( \23554_23853 , \23330_23632 , \23344_23646 );
and \U$14735 ( \23555_23854 , \23344_23646 , \23359_23661 );
and \U$14736 ( \23556_23855 , \23330_23632 , \23359_23661 );
or \U$14737 ( \23557_23856 , \23554_23853 , \23555_23854 , \23556_23855 );
and \U$14738 ( \23558_23857 , \23371_23673 , \23375_23677 );
and \U$14739 ( \23559_23858 , \23375_23677 , \23380_23682 );
and \U$14740 ( \23560_23859 , \23371_23673 , \23380_23682 );
or \U$14741 ( \23561_23860 , \23558_23857 , \23559_23858 , \23560_23859 );
and \U$14742 ( \23562_23861 , \17325_17627 , \15037_15336 );
and \U$14743 ( \23563_23862 , \17736_18035 , \14661_14963 );
nor \U$14744 ( \23564_23863 , \23562_23861 , \23563_23862 );
xnor \U$14745 ( \23565_23864 , \23564_23863 , \15043_15342 );
and \U$14746 ( \23566_23865 , \10968_11270 , \22243_22542 );
and \U$14747 ( \23567_23866 , \11287_11586 , \21801_22103 );
nor \U$14748 ( \23568_23867 , \23566_23865 , \23567_23866 );
xnor \U$14749 ( \23569_23868 , \23568_23867 , \22249_22548 );
xor \U$14750 ( \23570_23869 , \23565_23864 , \23569_23868 );
and \U$14751 ( \23571_23870 , RIdec53d8_708, \9034_9333 );
and \U$14752 ( \23572_23871 , RIdec26d8_676, \9036_9335 );
and \U$14753 ( \23573_23872 , RIee20080_4823, \9038_9337 );
and \U$14754 ( \23574_23873 , RIdebf9d8_644, \9040_9339 );
and \U$14755 ( \23575_23874 , RIee1f3d8_4814, \9042_9341 );
and \U$14756 ( \23576_23875 , RIdebccd8_612, \9044_9343 );
and \U$14757 ( \23577_23876 , RIdeb9fd8_580, \9046_9345 );
and \U$14758 ( \23578_23877 , RIdeb72d8_548, \9048_9347 );
and \U$14759 ( \23579_23878 , RIee1ee38_4810, \9050_9349 );
and \U$14760 ( \23580_23879 , RIdeb18d8_484, \9052_9351 );
and \U$14761 ( \23581_23880 , RIee1e898_4806, \9054_9353 );
and \U$14762 ( \23582_23881 , RIdeaebd8_452, \9056_9355 );
and \U$14763 ( \23583_23882 , RIee1da88_4796, \9058_9357 );
and \U$14764 ( \23584_23883 , RIdeaa420_420, \9060_9359 );
and \U$14765 ( \23585_23884 , RIdea3b20_388, \9062_9361 );
and \U$14766 ( \23586_23885 , RIde9d220_356, \9064_9363 );
and \U$14767 ( \23587_23886 , RIee1cde0_4787, \9066_9365 );
and \U$14768 ( \23588_23887 , RIee1bd00_4775, \9068_9367 );
and \U$14769 ( \23589_23888 , RIee1b490_4769, \9070_9369 );
and \U$14770 ( \23590_23889 , RIfcd8a28_7487, \9072_9371 );
and \U$14771 ( \23591_23890 , RIde91088_297, \9074_9373 );
and \U$14772 ( \23592_23891 , RIde8d8c0_280, \9076_9375 );
and \U$14773 ( \23593_23892 , RIfe7dac0_7774, \9078_9377 );
and \U$14774 ( \23594_23893 , RIfe7d958_7773, \9080_9379 );
and \U$14775 ( \23595_23894 , RIee1a518_4758, \9082_9381 );
and \U$14776 ( \23596_23895 , RIee19e10_4753, \9084_9383 );
and \U$14777 ( \23597_23896 , RIee19b40_4751, \9086_9385 );
and \U$14778 ( \23598_23897 , RIfc768c8_6371, \9088_9387 );
and \U$14779 ( \23599_23898 , RIfcd05f8_7393, \9090_9389 );
and \U$14780 ( \23600_23899 , RIfe7dd90_7776, \9092_9391 );
and \U$14781 ( \23601_23900 , RIee38770_5101, \9094_9393 );
and \U$14782 ( \23602_23901 , RIfe7dc28_7775, \9096_9395 );
and \U$14783 ( \23603_23902 , RIe1653d8_2529, \9098_9397 );
and \U$14784 ( \23604_23903 , RIe1626d8_2497, \9100_9399 );
and \U$14785 ( \23605_23904 , RIee373c0_5087, \9102_9401 );
and \U$14786 ( \23606_23905 , RIe15f9d8_2465, \9104_9403 );
and \U$14787 ( \23607_23906 , RIee362e0_5075, \9106_9405 );
and \U$14788 ( \23608_23907 , RIe15ccd8_2433, \9108_9407 );
and \U$14789 ( \23609_23908 , RIe1572d8_2369, \9110_9409 );
and \U$14790 ( \23610_23909 , RIe1545d8_2337, \9112_9411 );
and \U$14791 ( \23611_23910 , RIfe7def8_7777, \9114_9413 );
and \U$14792 ( \23612_23911 , RIe1518d8_2305, \9116_9415 );
and \U$14793 ( \23613_23912 , RIfebdeb8_8281, \9118_9417 );
and \U$14794 ( \23614_23913 , RIe14ebd8_2273, \9120_9419 );
and \U$14795 ( \23615_23914 , RIfc649e8_6167, \9122_9421 );
and \U$14796 ( \23616_23915 , RIe14bed8_2241, \9124_9423 );
and \U$14797 ( \23617_23916 , RIe1491d8_2209, \9126_9425 );
and \U$14798 ( \23618_23917 , RIe1464d8_2177, \9128_9427 );
and \U$14799 ( \23619_23918 , RIfe7d7f0_7772, \9130_9429 );
and \U$14800 ( \23620_23919 , RIfe7d688_7771, \9132_9431 );
and \U$14801 ( \23621_23920 , RIee32230_5029, \9134_9433 );
and \U$14802 ( \23622_23921 , RIfceb9e8_7703, \9136_9435 );
and \U$14803 ( \23623_23922 , RIfebdd50_8280, \9138_9437 );
and \U$14804 ( \23624_23923 , RIfe7d520_7770, \9140_9439 );
and \U$14805 ( \23625_23924 , RIfebdbe8_8279, \9142_9441 );
and \U$14806 ( \23626_23925 , RIfe7d3b8_7769, \9144_9443 );
and \U$14807 ( \23627_23926 , RIfc734c0_6334, \9146_9445 );
and \U$14808 ( \23628_23927 , RIee2f968_5000, \9148_9447 );
and \U$14809 ( \23629_23928 , RIfccfab8_7385, \9150_9449 );
and \U$14810 ( \23630_23929 , RIee2d7a8_4976, \9152_9451 );
and \U$14811 ( \23631_23930 , RIdf357a0_1985, \9154_9453 );
and \U$14812 ( \23632_23931 , RIdf33310_1959, \9156_9455 );
and \U$14813 ( \23633_23932 , RIdf312b8_1936, \9158_9457 );
and \U$14814 ( \23634_23933 , RIdf2f0f8_1912, \9160_9459 );
or \U$14815 ( \23635_23934 , \23571_23870 , \23572_23871 , \23573_23872 , \23574_23873 , \23575_23874 , \23576_23875 , \23577_23876 , \23578_23877 , \23579_23878 , \23580_23879 , \23581_23880 , \23582_23881 , \23583_23882 , \23584_23883 , \23585_23884 , \23586_23885 , \23587_23886 , \23588_23887 , \23589_23888 , \23590_23889 , \23591_23890 , \23592_23891 , \23593_23892 , \23594_23893 , \23595_23894 , \23596_23895 , \23597_23896 , \23598_23897 , \23599_23898 , \23600_23899 , \23601_23900 , \23602_23901 , \23603_23902 , \23604_23903 , \23605_23904 , \23606_23905 , \23607_23906 , \23608_23907 , \23609_23908 , \23610_23909 , \23611_23910 , \23612_23911 , \23613_23912 , \23614_23913 , \23615_23914 , \23616_23915 , \23617_23916 , \23618_23917 , \23619_23918 , \23620_23919 , \23621_23920 , \23622_23921 , \23623_23922 , \23624_23923 , \23625_23924 , \23626_23925 , \23627_23926 , \23628_23927 , \23629_23928 , \23630_23929 , \23631_23930 , \23632_23931 , \23633_23932 , \23634_23933 );
and \U$14816 ( \23636_23935 , RIee2bcf0_4957, \9163_9462 );
and \U$14817 ( \23637_23936 , RIee2a238_4938, \9165_9464 );
and \U$14818 ( \23638_23937 , RIee28e88_4924, \9167_9466 );
and \U$14819 ( \23639_23938 , RIee27c40_4911, \9169_9468 );
and \U$14820 ( \23640_23939 , RIfe7ce18_7765, \9171_9470 );
and \U$14821 ( \23641_23940 , RIfe7ccb0_7764, \9173_9472 );
and \U$14822 ( \23642_23941 , RIfe7cf80_7766, \9175_9474 );
and \U$14823 ( \23643_23942 , RIfe7cb48_7763, \9177_9476 );
and \U$14824 ( \23644_23943 , RIee27268_4904, \9179_9478 );
and \U$14825 ( \23645_23944 , RIee26e30_4901, \9181_9480 );
and \U$14826 ( \23646_23945 , RIee26890_4897, \9183_9482 );
and \U$14827 ( \23647_23946 , RIfcaa0d8_6957, \9185_9484 );
and \U$14828 ( \23648_23947 , RIee262f0_4893, \9187_9486 );
and \U$14829 ( \23649_23948 , RIfe7d250_7768, \9189_9488 );
and \U$14830 ( \23650_23949 , RIee26020_4891, \9191_9490 );
and \U$14831 ( \23651_23950 , RIfe7d0e8_7767, \9193_9492 );
and \U$14832 ( \23652_23951 , RIdf16fa8_1638, \9195_9494 );
and \U$14833 ( \23653_23952 , RIdf142a8_1606, \9197_9496 );
and \U$14834 ( \23654_23953 , RIdf115a8_1574, \9199_9498 );
and \U$14835 ( \23655_23954 , RIdf0e8a8_1542, \9201_9500 );
and \U$14836 ( \23656_23955 , RIdf0bba8_1510, \9203_9502 );
and \U$14837 ( \23657_23956 , RIdf08ea8_1478, \9205_9504 );
and \U$14838 ( \23658_23957 , RIdf061a8_1446, \9207_9506 );
and \U$14839 ( \23659_23958 , RIdf034a8_1414, \9209_9508 );
and \U$14840 ( \23660_23959 , RIdefdaa8_1350, \9211_9510 );
and \U$14841 ( \23661_23960 , RIdefada8_1318, \9213_9512 );
and \U$14842 ( \23662_23961 , RIdef80a8_1286, \9215_9514 );
and \U$14843 ( \23663_23962 , RIdef53a8_1254, \9217_9516 );
and \U$14844 ( \23664_23963 , RIdef26a8_1222, \9219_9518 );
and \U$14845 ( \23665_23964 , RIdeef9a8_1190, \9221_9520 );
and \U$14846 ( \23666_23965 , RIdeecca8_1158, \9223_9522 );
and \U$14847 ( \23667_23966 , RIdee9fa8_1126, \9225_9524 );
and \U$14848 ( \23668_23967 , RIee25648_4884, \9227_9526 );
and \U$14849 ( \23669_23968 , RIee249a0_4875, \9229_9528 );
and \U$14850 ( \23670_23969 , RIfebe020_8282, \9231_9530 );
and \U$14851 ( \23671_23970 , RIee23488_4860, \9233_9532 );
and \U$14852 ( \23672_23971 , RIfebe2f0_8284, \9235_9534 );
and \U$14853 ( \23673_23972 , RIfebe188_8283, \9237_9536 );
and \U$14854 ( \23674_23973 , RIfe7e1c8_7779, \9239_9538 );
and \U$14855 ( \23675_23974 , RIfe7e060_7778, \9241_9540 );
and \U$14856 ( \23676_23975 , RIfcbf7f8_7201, \9243_9542 );
and \U$14857 ( \23677_23976 , RIfc7aae0_6418, \9245_9544 );
and \U$14858 ( \23678_23977 , RIfc787b8_6393, \9247_9546 );
and \U$14859 ( \23679_23978 , RIfc618b0_6132, \9249_9548 );
and \U$14860 ( \23680_23979 , RIded98b0_939, \9251_9550 );
and \U$14861 ( \23681_23980 , RIded72b8_912, \9253_9552 );
and \U$14862 ( \23682_23981 , RIded5530_891, \9255_9554 );
and \U$14863 ( \23683_23982 , RIded2dd0_863, \9257_9556 );
and \U$14864 ( \23684_23983 , RIded07d8_836, \9259_9558 );
and \U$14865 ( \23685_23984 , RIdecdad8_804, \9261_9560 );
and \U$14866 ( \23686_23985 , RIdecadd8_772, \9263_9562 );
and \U$14867 ( \23687_23986 , RIdec80d8_740, \9265_9564 );
and \U$14868 ( \23688_23987 , RIdeb45d8_516, \9267_9566 );
and \U$14869 ( \23689_23988 , RIde96920_324, \9269_9568 );
and \U$14870 ( \23690_23989 , RIe16e1e0_2630, \9271_9570 );
and \U$14871 ( \23691_23990 , RIe159fd8_2401, \9273_9572 );
and \U$14872 ( \23692_23991 , RIe1437d8_2145, \9275_9574 );
and \U$14873 ( \23693_23992 , RIdf381d0_2015, \9277_9576 );
and \U$14874 ( \23694_23993 , RIdf2c830_1883, \9279_9578 );
and \U$14875 ( \23695_23994 , RIdf1d0b0_1707, \9281_9580 );
and \U$14876 ( \23696_23995 , RIdf007a8_1382, \9283_9582 );
and \U$14877 ( \23697_23996 , RIdee72a8_1094, \9285_9584 );
and \U$14878 ( \23698_23997 , RIdedc010_967, \9287_9586 );
and \U$14879 ( \23699_23998 , RIde7c868_197, \9289_9588 );
or \U$14880 ( \23700_23999 , \23636_23935 , \23637_23936 , \23638_23937 , \23639_23938 , \23640_23939 , \23641_23940 , \23642_23941 , \23643_23942 , \23644_23943 , \23645_23944 , \23646_23945 , \23647_23946 , \23648_23947 , \23649_23948 , \23650_23949 , \23651_23950 , \23652_23951 , \23653_23952 , \23654_23953 , \23655_23954 , \23656_23955 , \23657_23956 , \23658_23957 , \23659_23958 , \23660_23959 , \23661_23960 , \23662_23961 , \23663_23962 , \23664_23963 , \23665_23964 , \23666_23965 , \23667_23966 , \23668_23967 , \23669_23968 , \23670_23969 , \23671_23970 , \23672_23971 , \23673_23972 , \23674_23973 , \23675_23974 , \23676_23975 , \23677_23976 , \23678_23977 , \23679_23978 , \23680_23979 , \23681_23980 , \23682_23981 , \23683_23982 , \23684_23983 , \23685_23984 , \23686_23985 , \23687_23986 , \23688_23987 , \23689_23988 , \23690_23989 , \23691_23990 , \23692_23991 , \23693_23992 , \23694_23993 , \23695_23994 , \23696_23995 , \23697_23996 , \23698_23997 , \23699_23998 );
or \U$14881 ( \23701_24000 , \23635_23934 , \23700_23999 );
_DC \g5a97/U$1 ( \23702 , \23701_24000 , \9298_9597 );
and \U$14882 ( \23703_24002 , RIe19d670_3168, \8760_9059 );
and \U$14883 ( \23704_24003 , RIe19a970_3136, \8762_9061 );
and \U$14884 ( \23705_24004 , RIfe7b630_7748, \8764_9063 );
and \U$14885 ( \23706_24005 , RIe197c70_3104, \8766_9065 );
and \U$14886 ( \23707_24006 , RIfe7b4c8_7747, \8768_9067 );
and \U$14887 ( \23708_24007 , RIe194f70_3072, \8770_9069 );
and \U$14888 ( \23709_24008 , RIe192270_3040, \8772_9071 );
and \U$14889 ( \23710_24009 , RIe18f570_3008, \8774_9073 );
and \U$14890 ( \23711_24010 , RIe189b70_2944, \8776_9075 );
and \U$14891 ( \23712_24011 , RIe186e70_2912, \8778_9077 );
and \U$14892 ( \23713_24012 , RIfe7b360_7746, \8780_9079 );
and \U$14893 ( \23714_24013 , RIe184170_2880, \8782_9081 );
and \U$14894 ( \23715_24014 , RIfe7b1f8_7745, \8784_9083 );
and \U$14895 ( \23716_24015 , RIe181470_2848, \8786_9085 );
and \U$14896 ( \23717_24016 , RIe17e770_2816, \8788_9087 );
and \U$14897 ( \23718_24017 , RIe17ba70_2784, \8790_9089 );
and \U$14898 ( \23719_24018 , RIf1423b8_5213, \8792_9091 );
and \U$14899 ( \23720_24019 , RIf140ea0_5198, \8794_9093 );
and \U$14900 ( \23721_24020 , RIf140360_5190, \8796_9095 );
and \U$14901 ( \23722_24021 , RIfe7b798_7749, \8798_9097 );
and \U$14902 ( \23723_24022 , RIf13fc58_5185, \8800_9099 );
and \U$14903 ( \23724_24023 , RIf13f280_5178, \8802_9101 );
and \U$14904 ( \23725_24024 , RIfc79460_6402, \8804_9103 );
and \U$14905 ( \23726_24025 , RIee3d4c8_5156, \8806_9105 );
and \U$14906 ( \23727_24026 , RIfe7b090_7744, \8808_9107 );
and \U$14907 ( \23728_24027 , RIfe7af28_7743, \8810_9109 );
and \U$14908 ( \23729_24028 , RIee39df0_5117, \8812_9111 );
and \U$14909 ( \23730_24029 , RIe1737a8_2691, \8814_9113 );
and \U$14910 ( \23731_24030 , RIfe7adc0_7742, \8816_9115 );
and \U$14911 ( \23732_24031 , RIfe7ac58_7741, \8818_9117 );
and \U$14912 ( \23733_24032 , RIf16e440_5714, \8820_9119 );
and \U$14913 ( \23734_24033 , RIfcb20d0_7048, \8822_9121 );
and \U$14914 ( \23735_24034 , RIfe7bd38_7753, \8824_9123 );
and \U$14915 ( \23736_24035 , RIe2239c8_4695, \8826_9125 );
and \U$14916 ( \23737_24036 , RIf16be48_5687, \8828_9127 );
and \U$14917 ( \23738_24037 , RIe220cc8_4663, \8830_9129 );
and \U$14918 ( \23739_24038 , RIf16aed0_5676, \8832_9131 );
and \U$14919 ( \23740_24039 , RIe21dfc8_4631, \8834_9133 );
and \U$14920 ( \23741_24040 , RIe2185c8_4567, \8836_9135 );
and \U$14921 ( \23742_24041 , RIe2158c8_4535, \8838_9137 );
and \U$14922 ( \23743_24042 , RIfebd7b0_8276, \8840_9139 );
and \U$14923 ( \23744_24043 , RIe212bc8_4503, \8842_9141 );
and \U$14924 ( \23745_24044 , RIfebd648_8275, \8844_9143 );
and \U$14925 ( \23746_24045 , RIe20fec8_4471, \8846_9145 );
and \U$14926 ( \23747_24046 , RIfe7b900_7750, \8848_9147 );
and \U$14927 ( \23748_24047 , RIe20d1c8_4439, \8850_9149 );
and \U$14928 ( \23749_24048 , RIe20a4c8_4407, \8852_9151 );
and \U$14929 ( \23750_24049 , RIe2077c8_4375, \8854_9153 );
and \U$14930 ( \23751_24050 , RIf167258_5633, \8856_9155 );
and \U$14931 ( \23752_24051 , RIf166178_5621, \8858_9157 );
and \U$14932 ( \23753_24052 , RIe2024d0_4316, \8860_9159 );
and \U$14933 ( \23754_24053 , RIfe7bbd0_7752, \8862_9161 );
and \U$14934 ( \23755_24054 , RIf165368_5611, \8864_9163 );
and \U$14935 ( \23756_24055 , RIf1646c0_5602, \8866_9165 );
and \U$14936 ( \23757_24056 , RIfcd0a30_7396, \8868_9167 );
and \U$14937 ( \23758_24057 , RIf1620c8_5575, \8870_9169 );
and \U$14938 ( \23759_24058 , RIf1601d8_5553, \8872_9171 );
and \U$14939 ( \23760_24059 , RIf15e2e8_5531, \8874_9173 );
and \U$14940 ( \23761_24060 , RIfe7ba68_7751, \8876_9175 );
and \U$14941 ( \23762_24061 , RIfe7bea0_7754, \8878_9177 );
and \U$14942 ( \23763_24062 , RIf15cdd0_5516, \8880_9179 );
and \U$14943 ( \23764_24063 , RIf15b8b8_5501, \8882_9181 );
and \U$14944 ( \23765_24064 , RIf15a7d8_5489, \8884_9183 );
and \U$14945 ( \23766_24065 , RIfca4840_6894, \8886_9185 );
or \U$14946 ( \23767_24066 , \23703_24002 , \23704_24003 , \23705_24004 , \23706_24005 , \23707_24006 , \23708_24007 , \23709_24008 , \23710_24009 , \23711_24010 , \23712_24011 , \23713_24012 , \23714_24013 , \23715_24014 , \23716_24015 , \23717_24016 , \23718_24017 , \23719_24018 , \23720_24019 , \23721_24020 , \23722_24021 , \23723_24022 , \23724_24023 , \23725_24024 , \23726_24025 , \23727_24026 , \23728_24027 , \23729_24028 , \23730_24029 , \23731_24030 , \23732_24031 , \23733_24032 , \23734_24033 , \23735_24034 , \23736_24035 , \23737_24036 , \23738_24037 , \23739_24038 , \23740_24039 , \23741_24040 , \23742_24041 , \23743_24042 , \23744_24043 , \23745_24044 , \23746_24045 , \23747_24046 , \23748_24047 , \23749_24048 , \23750_24049 , \23751_24050 , \23752_24051 , \23753_24052 , \23754_24053 , \23755_24054 , \23756_24055 , \23757_24056 , \23758_24057 , \23759_24058 , \23760_24059 , \23761_24060 , \23762_24061 , \23763_24062 , \23764_24063 , \23765_24064 , \23766_24065 );
and \U$14947 ( \23768_24067 , RIf158ff0_5472, \8889_9188 );
and \U$14948 ( \23769_24068 , RIf157c40_5458, \8891_9190 );
and \U$14949 ( \23770_24069 , RIf156f98_5449, \8893_9192 );
and \U$14950 ( \23771_24070 , RIfe7c170_7756, \8895_9194 );
and \U$14951 ( \23772_24071 , RIf156458_5441, \8897_9196 );
and \U$14952 ( \23773_24072 , RIf155918_5433, \8899_9198 );
and \U$14953 ( \23774_24073 , RIf1549a0_5422, \8901_9200 );
and \U$14954 ( \23775_24074 , RIe1f54b0_4168, \8903_9202 );
and \U$14955 ( \23776_24075 , RIfe7c008_7755, \8905_9204 );
and \U$14956 ( \23777_24076 , RIf151b38_5389, \8907_9206 );
and \U$14957 ( \23778_24077 , RIf150bc0_5378, \8909_9208 );
and \U$14958 ( \23779_24078 , RIe1f32f0_4144, \8911_9210 );
and \U$14959 ( \23780_24079 , RIf14fae0_5366, \8913_9212 );
and \U$14960 ( \23781_24080 , RIf14ee38_5357, \8915_9214 );
and \U$14961 ( \23782_24081 , RIf14e028_5347, \8917_9216 );
and \U$14962 ( \23783_24082 , RIe1edff8_4085, \8919_9218 );
and \U$14963 ( \23784_24083 , RIe1eb730_4056, \8921_9220 );
and \U$14964 ( \23785_24084 , RIe1e8a30_4024, \8923_9222 );
and \U$14965 ( \23786_24085 , RIe1e5d30_3992, \8925_9224 );
and \U$14966 ( \23787_24086 , RIe1e3030_3960, \8927_9226 );
and \U$14967 ( \23788_24087 , RIe1e0330_3928, \8929_9228 );
and \U$14968 ( \23789_24088 , RIe1dd630_3896, \8931_9230 );
and \U$14969 ( \23790_24089 , RIe1da930_3864, \8933_9232 );
and \U$14970 ( \23791_24090 , RIe1d7c30_3832, \8935_9234 );
and \U$14971 ( \23792_24091 , RIe1d2230_3768, \8937_9236 );
and \U$14972 ( \23793_24092 , RIe1cf530_3736, \8939_9238 );
and \U$14973 ( \23794_24093 , RIe1cc830_3704, \8941_9240 );
and \U$14974 ( \23795_24094 , RIe1c9b30_3672, \8943_9242 );
and \U$14975 ( \23796_24095 , RIe1c6e30_3640, \8945_9244 );
and \U$14976 ( \23797_24096 , RIe1c4130_3608, \8947_9246 );
and \U$14977 ( \23798_24097 , RIe1c1430_3576, \8949_9248 );
and \U$14978 ( \23799_24098 , RIe1be730_3544, \8951_9250 );
and \U$14979 ( \23800_24099 , RIf14cb10_5332, \8953_9252 );
and \U$14980 ( \23801_24100 , RIf14b8c8_5319, \8955_9254 );
and \U$14981 ( \23802_24101 , RIfebda80_8278, \8957_9256 );
and \U$14982 ( \23803_24102 , RIfe7c878_7761, \8959_9258 );
and \U$14983 ( \23804_24103 , RIf14a680_5306, \8961_9260 );
and \U$14984 ( \23805_24104 , RIfe7c2d8_7757, \8963_9262 );
and \U$14985 ( \23806_24105 , RIfe7c9e0_7762, \8965_9264 );
and \U$14986 ( \23807_24106 , RIfe7c440_7758, \8967_9266 );
and \U$14987 ( \23808_24107 , RIf149000_5290, \8969_9268 );
and \U$14988 ( \23809_24108 , RIf147db8_5277, \8971_9270 );
and \U$14989 ( \23810_24109 , RIe1b2688_3407, \8973_9272 );
and \U$14990 ( \23811_24110 , RIfebd918_8277, \8975_9274 );
and \U$14991 ( \23812_24111 , RIfe7c5a8_7759, \8977_9276 );
and \U$14992 ( \23813_24112 , RIf146738_5261, \8979_9278 );
and \U$14993 ( \23814_24113 , RIfe7c710_7760, \8981_9280 );
and \U$14994 ( \23815_24114 , RIe1aad98_3321, \8983_9282 );
and \U$14995 ( \23816_24115 , RIe1a8a70_3296, \8985_9284 );
and \U$14996 ( \23817_24116 , RIe1a5d70_3264, \8987_9286 );
and \U$14997 ( \23818_24117 , RIe1a3070_3232, \8989_9288 );
and \U$14998 ( \23819_24118 , RIe1a0370_3200, \8991_9290 );
and \U$14999 ( \23820_24119 , RIe18c870_2976, \8993_9292 );
and \U$15000 ( \23821_24120 , RIe178d70_2752, \8995_9294 );
and \U$15001 ( \23822_24121 , RIe2266c8_4727, \8997_9296 );
and \U$15002 ( \23823_24122 , RIe21b2c8_4599, \8999_9298 );
and \U$15003 ( \23824_24123 , RIe204ac8_4343, \9001_9300 );
and \U$15004 ( \23825_24124 , RIe1feb28_4275, \9003_9302 );
and \U$15005 ( \23826_24125 , RIe1f7ee0_4198, \9005_9304 );
and \U$15006 ( \23827_24126 , RIe1f0a28_4115, \9007_9306 );
and \U$15007 ( \23828_24127 , RIe1d4f30_3800, \9009_9308 );
and \U$15008 ( \23829_24128 , RIe1bba30_3512, \9011_9310 );
and \U$15009 ( \23830_24129 , RIe1ae8a8_3363, \9013_9312 );
and \U$15010 ( \23831_24130 , RIe170ee0_2662, \9015_9314 );
or \U$15011 ( \23832_24131 , \23768_24067 , \23769_24068 , \23770_24069 , \23771_24070 , \23772_24071 , \23773_24072 , \23774_24073 , \23775_24074 , \23776_24075 , \23777_24076 , \23778_24077 , \23779_24078 , \23780_24079 , \23781_24080 , \23782_24081 , \23783_24082 , \23784_24083 , \23785_24084 , \23786_24085 , \23787_24086 , \23788_24087 , \23789_24088 , \23790_24089 , \23791_24090 , \23792_24091 , \23793_24092 , \23794_24093 , \23795_24094 , \23796_24095 , \23797_24096 , \23798_24097 , \23799_24098 , \23800_24099 , \23801_24100 , \23802_24101 , \23803_24102 , \23804_24103 , \23805_24104 , \23806_24105 , \23807_24106 , \23808_24107 , \23809_24108 , \23810_24109 , \23811_24110 , \23812_24111 , \23813_24112 , \23814_24113 , \23815_24114 , \23816_24115 , \23817_24116 , \23818_24117 , \23819_24118 , \23820_24119 , \23821_24120 , \23822_24121 , \23823_24122 , \23824_24123 , \23825_24124 , \23826_24125 , \23827_24126 , \23828_24127 , \23829_24128 , \23830_24129 , \23831_24130 );
or \U$15012 ( \23833_24132 , \23767_24066 , \23832_24131 );
_DC \g5b1b/U$1 ( \23834 , \23833_24132 , \9024_9323 );
xor g5b1c_GF_PartitionCandidate( \23835_24134_nG5b1c , \23702 , \23834 );
buf \U$15013 ( \23836_24135 , \23835_24134_nG5b1c );
xor \U$15014 ( \23837_24136 , \23836_24135 , \23327_23629 );
not \U$15015 ( \23838_24137 , \23328_23630 );
and \U$15016 ( \23839_24138 , \23837_24136 , \23838_24137 );
and \U$15017 ( \23840_24139 , \10385_10687 , \23839_24138 );
and \U$15018 ( \23841_24140 , \10686_10988 , \23328_23630 );
nor \U$15019 ( \23842_24141 , \23840_24139 , \23841_24140 );
and \U$15020 ( \23843_24142 , \23327_23629 , \22240_22539 );
not \U$15021 ( \23844_24143 , \23843_24142 );
and \U$15022 ( \23845_24144 , \23836_24135 , \23844_24143 );
xnor \U$15023 ( \23846_24145 , \23842_24141 , \23845_24144 );
xor \U$15024 ( \23847_24146 , \23570_23869 , \23846_24145 );
xor \U$15025 ( \23848_24147 , \23561_23860 , \23847_24146 );
and \U$15026 ( \23849_24148 , \18730_19032 , \13755_14054 );
and \U$15027 ( \23850_24149 , \19259_19558 , \13390_13692 );
nor \U$15028 ( \23851_24150 , \23849_24148 , \23850_24149 );
xnor \U$15029 ( \23852_24151 , \23851_24150 , \13736_14035 );
and \U$15030 ( \23853_24152 , \13377_13679 , \19235_19534 );
and \U$15031 ( \23854_24153 , \13725_14024 , \18743_19045 );
nor \U$15032 ( \23855_24154 , \23853_24152 , \23854_24153 );
xnor \U$15033 ( \23856_24155 , \23855_24154 , \19241_19540 );
xor \U$15034 ( \23857_24156 , \23852_24151 , \23856_24155 );
and \U$15035 ( \23858_24157 , \12146_12448 , \20706_21005 );
and \U$15036 ( \23859_24158 , \12470_12769 , \20255_20557 );
nor \U$15037 ( \23860_24159 , \23858_24157 , \23859_24158 );
xnor \U$15038 ( \23861_24160 , \23860_24159 , \20712_21011 );
xor \U$15039 ( \23862_24161 , \23857_24156 , \23861_24160 );
xor \U$15040 ( \23863_24162 , \23848_24147 , \23862_24161 );
xor \U$15041 ( \23864_24163 , \23557_23856 , \23863_24162 );
and \U$15042 ( \23865_24164 , \23038_23340 , \23042_23344 );
and \U$15043 ( \23866_24165 , \23042_23344 , \23047_23349 );
and \U$15044 ( \23867_24166 , \23038_23340 , \23047_23349 );
or \U$15045 ( \23868_24167 , \23865_24164 , \23866_24165 , \23867_24166 );
and \U$15046 ( \23869_24168 , \21788_22090 , \11275_11574 );
and \U$15047 ( \23870_24169 , \22257_22556 , \10976_11278 );
nor \U$15048 ( \23871_24170 , \23869_24168 , \23870_24169 );
xnor \U$15049 ( \23872_24171 , \23871_24170 , \11281_11580 );
not \U$15050 ( \23873_24172 , \23329_23631 );
and \U$15051 ( \23874_24173 , \23873_24172 , \23845_24144 );
xor \U$15052 ( \23875_24174 , \23872_24171 , \23874_24173 );
and \U$15053 ( \23876_24175 , \23349_23651 , \23353_23655 );
and \U$15054 ( \23877_24176 , \23353_23655 , \23358_23660 );
and \U$15055 ( \23878_24177 , \23349_23651 , \23358_23660 );
or \U$15056 ( \23879_24178 , \23876_24175 , \23877_24176 , \23878_24177 );
xor \U$15057 ( \23880_24179 , \23875_24174 , \23879_24178 );
and \U$15058 ( \23881_24180 , \14648_14950 , \17791_18090 );
and \U$15059 ( \23882_24181 , \15022_15321 , \17353_17655 );
nor \U$15060 ( \23883_24182 , \23881_24180 , \23882_24181 );
xnor \U$15061 ( \23884_24183 , \23883_24182 , \17747_18046 );
xor \U$15062 ( \23885_24184 , \23880_24179 , \23884_24183 );
xor \U$15063 ( \23886_24185 , \23868_24167 , \23885_24184 );
and \U$15064 ( \23887_24186 , \23318_23620 , \23322_23624 );
and \U$15065 ( \23888_24187 , \23322_23624 , \23329_23631 );
and \U$15066 ( \23889_24188 , \23318_23620 , \23329_23631 );
or \U$15067 ( \23890_24189 , \23887_24186 , \23888_24187 , \23889_24188 );
and \U$15068 ( \23891_24190 , \23334_23636 , \23338_23640 );
and \U$15069 ( \23892_24191 , \23338_23640 , \23343_23645 );
and \U$15070 ( \23893_24192 , \23334_23636 , \23343_23645 );
or \U$15071 ( \23894_24193 , \23891_24190 , \23892_24191 , \23893_24192 );
xor \U$15072 ( \23895_24194 , \23890_24189 , \23894_24193 );
and \U$15073 ( \23896_24195 , \23315_23617 , \10681_10983 );
_DC \g65b6/U$1 ( \23897 , \23701_24000 , \9298_9597 );
_DC \g65b7/U$1 ( \23898 , \23833_24132 , \9024_9323 );
and g65b8_GF_PartitionCandidate( \23899_24198_nG65b8 , \23897 , \23898 );
buf \U$15074 ( \23900_24199 , \23899_24198_nG65b8 );
and \U$15075 ( \23901_24200 , \23900_24199 , \10389_10691 );
nor \U$15076 ( \23902_24201 , \23896_24195 , \23901_24200 );
xnor \U$15077 ( \23903_24202 , \23902_24201 , \10678_10980 );
and \U$15078 ( \23904_24203 , \20242_20544 , \12491_12790 );
and \U$15079 ( \23905_24204 , \20734_21033 , \12159_12461 );
nor \U$15080 ( \23906_24205 , \23904_24203 , \23905_24204 );
xnor \U$15081 ( \23907_24206 , \23906_24205 , \12481_12780 );
xor \U$15082 ( \23908_24207 , \23903_24202 , \23907_24206 );
and \U$15083 ( \23909_24208 , \15965_16267 , \16333_16635 );
and \U$15084 ( \23910_24209 , \16353_16655 , \15999_16301 );
nor \U$15085 ( \23911_24210 , \23909_24208 , \23910_24209 );
xnor \U$15086 ( \23912_24211 , \23911_24210 , \16323_16625 );
xor \U$15087 ( \23913_24212 , \23908_24207 , \23912_24211 );
xor \U$15088 ( \23914_24213 , \23895_24194 , \23913_24212 );
xor \U$15089 ( \23915_24214 , \23886_24185 , \23914_24213 );
xor \U$15090 ( \23916_24215 , \23864_24163 , \23915_24214 );
xor \U$15091 ( \23917_24216 , \23553_23852 , \23916_24215 );
and \U$15092 ( \23918_24217 , \23029_23331 , \23033_23335 );
and \U$15093 ( \23919_24218 , \23033_23335 , \23383_23685 );
and \U$15094 ( \23920_24219 , \23029_23331 , \23383_23685 );
or \U$15095 ( \23921_24220 , \23918_24217 , \23919_24218 , \23920_24219 );
xor \U$15096 ( \23922_24221 , \23917_24216 , \23921_24220 );
and \U$15097 ( \23923_24222 , \23384_23686 , \23388_23690 );
and \U$15098 ( \23924_24223 , \23389_23691 , \23392_23694 );
or \U$15099 ( \23925_24224 , \23923_24222 , \23924_24223 );
xor \U$15100 ( \23926_24225 , \23922_24221 , \23925_24224 );
buf g9bcf_GF_PartitionCandidate( \23927_24226_nG9bcf , \23926_24225 );
and \U$15101 ( \23928_24227 , \10402_10704 , \23927_24226_nG9bcf );
or \U$15102 ( \23929_24228 , \23544_23843 , \23928_24227 );
xor \U$15103 ( \23930_24229 , \10399_10703 , \23929_24228 );
buf \U$15104 ( \23931_24230 , \23930_24229 );
buf \U$15106 ( \23932_24231 , \23931_24230 );
xor \U$15107 ( \23933_24232 , \23543_23842 , \23932_24231 );
buf \U$15108 ( \23934_24233 , \23933_24232 );
xor \U$15109 ( \23935_24234 , \23453_23755 , \23934_24233 );
and \U$15110 ( \23936_24235 , \23415_23717 , \23935_24234 );
and \U$15111 ( \23937_24236 , \23405_23707 , \23409_23711 );
and \U$15112 ( \23938_24237 , \23405_23707 , \23414_23716 );
and \U$15113 ( \23939_24238 , \23409_23711 , \23414_23716 );
or \U$15114 ( \23940_24239 , \23937_24236 , \23938_24237 , \23939_24238 );
xor \U$15115 ( \23941_24240 , \23936_24235 , \23940_24239 );
and \U$15116 ( \23942_24241 , RIdec56a8_710, \8760_9059 );
and \U$15117 ( \23943_24242 , RIdec29a8_678, \8762_9061 );
and \U$15118 ( \23944_24243 , RIfc54020_5978, \8764_9063 );
and \U$15119 ( \23945_24244 , RIdebfca8_646, \8766_9065 );
and \U$15120 ( \23946_24245 , RIee1f540_4815, \8768_9067 );
and \U$15121 ( \23947_24246 , RIdebcfa8_614, \8770_9069 );
and \U$15122 ( \23948_24247 , RIdeba2a8_582, \8772_9071 );
and \U$15123 ( \23949_24248 , RIdeb75a8_550, \8774_9073 );
and \U$15124 ( \23950_24249 , RIfc4fe08_5931, \8776_9075 );
and \U$15125 ( \23951_24250 , RIdeb1ba8_486, \8778_9077 );
and \U$15126 ( \23952_24251 , RIfc6b630_6244, \8780_9079 );
and \U$15127 ( \23953_24252 , RIdeaeea8_454, \8782_9081 );
and \U$15128 ( \23954_24253 , RIfc6a118_6229, \8784_9083 );
and \U$15129 ( \23955_24254 , RIdeaaab0_422, \8786_9085 );
and \U$15130 ( \23956_24255 , RIdea41b0_390, \8788_9087 );
and \U$15131 ( \23957_24256 , RIde9d8b0_358, \8790_9089 );
and \U$15132 ( \23958_24257 , RIfc69ce0_6226, \8792_9091 );
and \U$15133 ( \23959_24258 , RIee1be68_4776, \8794_9093 );
and \U$15134 ( \23960_24259 , RIfc653c0_6174, \8796_9095 );
and \U$15135 ( \23961_24260 , RIee1ac20_4763, \8798_9097 );
and \U$15136 ( \23962_24261 , RIde91718_299, \8800_9099 );
and \U$15137 ( \23963_24262 , RIde8df50_282, \8802_9101 );
and \U$15138 ( \23964_24263 , RIde89db0_262, \8804_9103 );
and \U$15139 ( \23965_24264 , RIde85c10_242, \8806_9105 );
and \U$15140 ( \23966_24265 , RIde81db8_223, \8808_9107 );
and \U$15141 ( \23967_24266 , RIfca76a8_6927, \8810_9109 );
and \U$15142 ( \23968_24267 , RIfcca4f0_7324, \8812_9111 );
and \U$15143 ( \23969_24268 , RIfc4ce38_5897, \8814_9113 );
and \U$15144 ( \23970_24269 , RIfc6b360_6242, \8816_9115 );
and \U$15145 ( \23971_24270 , RIe16b918_2601, \8818_9117 );
and \U$15146 ( \23972_24271 , RIe169cf8_2581, \8820_9119 );
and \U$15147 ( \23973_24272 , RIe167f70_2560, \8822_9121 );
and \U$15148 ( \23974_24273 , RIe1656a8_2531, \8824_9123 );
and \U$15149 ( \23975_24274 , RIe1629a8_2499, \8826_9125 );
and \U$15150 ( \23976_24275 , RIee37690_5089, \8828_9127 );
and \U$15151 ( \23977_24276 , RIe15fca8_2467, \8830_9129 );
and \U$15152 ( \23978_24277 , RIfce93f0_7676, \8832_9131 );
and \U$15153 ( \23979_24278 , RIe15cfa8_2435, \8834_9133 );
and \U$15154 ( \23980_24279 , RIe1575a8_2371, \8836_9135 );
and \U$15155 ( \23981_24280 , RIe1548a8_2339, \8838_9137 );
and \U$15156 ( \23982_24281 , RIee35908_5068, \8840_9139 );
and \U$15157 ( \23983_24282 , RIe151ba8_2307, \8842_9141 );
and \U$15158 ( \23984_24283 , RIee34f30_5061, \8844_9143 );
and \U$15159 ( \23985_24284 , RIe14eea8_2275, \8846_9145 );
and \U$15160 ( \23986_24285 , RIfce32e8_7607, \8848_9147 );
and \U$15161 ( \23987_24286 , RIe14c1a8_2243, \8850_9149 );
and \U$15162 ( \23988_24287 , RIe1494a8_2211, \8852_9151 );
and \U$15163 ( \23989_24288 , RIe1467a8_2179, \8854_9153 );
and \U$15164 ( \23990_24289 , RIfcde2c0_7550, \8856_9155 );
and \U$15165 ( \23991_24290 , RIfc687c8_6211, \8858_9157 );
and \U$15166 ( \23992_24291 , RIfca9160_6946, \8860_9159 );
and \U$15167 ( \23993_24292 , RIfcb1590_7040, \8862_9161 );
and \U$15168 ( \23994_24293 , RIe141078_2117, \8864_9163 );
and \U$15169 ( \23995_24294 , RIdf3ef80_2093, \8866_9165 );
and \U$15170 ( \23996_24295 , RIdf3cdc0_2069, \8868_9167 );
and \U$15171 ( \23997_24296 , RIfebeb60_8290, \8870_9169 );
and \U$15172 ( \23998_24297 , RIfc64448_6163, \8872_9171 );
and \U$15173 ( \23999_24298 , RIee2fad0_5001, \8874_9173 );
and \U$15174 ( \24000_24299 , RIfca7978_6929, \8876_9175 );
and \U$15175 ( \24001_24300 , RIfc676e8_6199, \8878_9177 );
and \U$15176 ( \24002_24301 , RIdf35a70_1987, \8880_9179 );
and \U$15177 ( \24003_24302 , RIdf335e0_1961, \8882_9181 );
and \U$15178 ( \24004_24303 , RIdf31420_1937, \8884_9183 );
and \U$15179 ( \24005_24304 , RIdf2f3c8_1914, \8886_9185 );
or \U$15180 ( \24006_24305 , \23942_24241 , \23943_24242 , \23944_24243 , \23945_24244 , \23946_24245 , \23947_24246 , \23948_24247 , \23949_24248 , \23950_24249 , \23951_24250 , \23952_24251 , \23953_24252 , \23954_24253 , \23955_24254 , \23956_24255 , \23957_24256 , \23958_24257 , \23959_24258 , \23960_24259 , \23961_24260 , \23962_24261 , \23963_24262 , \23964_24263 , \23965_24264 , \23966_24265 , \23967_24266 , \23968_24267 , \23969_24268 , \23970_24269 , \23971_24270 , \23972_24271 , \23973_24272 , \23974_24273 , \23975_24274 , \23976_24275 , \23977_24276 , \23978_24277 , \23979_24278 , \23980_24279 , \23981_24280 , \23982_24281 , \23983_24282 , \23984_24283 , \23985_24284 , \23986_24285 , \23987_24286 , \23988_24287 , \23989_24288 , \23990_24289 , \23991_24290 , \23992_24291 , \23993_24292 , \23994_24293 , \23995_24294 , \23996_24295 , \23997_24296 , \23998_24297 , \23999_24298 , \24000_24299 , \24001_24300 , \24002_24301 , \24003_24302 , \24004_24303 , \24005_24304 );
and \U$15181 ( \24007_24306 , RIfccef78_7377, \8889_9188 );
and \U$15182 ( \24008_24307 , RIfca6fa0_6922, \8891_9190 );
and \U$15183 ( \24009_24308 , RIfc62558_6141, \8893_9192 );
and \U$15184 ( \24010_24309 , RIfc61fb8_6137, \8895_9194 );
and \U$15185 ( \24011_24310 , RIfe81b70_7820, \8897_9196 );
and \U$15186 ( \24012_24311 , RIdf281e0_1833, \8899_9198 );
and \U$15187 ( \24013_24312 , RIfe81cd8_7821, \8901_9200 );
and \U$15188 ( \24014_24313 , RIdf249a0_1793, \8903_9202 );
and \U$15189 ( \24015_24314 , RIfc44300_5798, \8905_9204 );
and \U$15190 ( \24016_24315 , RIfcafc40_7022, \8907_9206 );
and \U$15191 ( \24017_24316 , RIdf22ee8_1774, \8909_9208 );
and \U$15192 ( \24018_24317 , RIfcaac18_6965, \8911_9210 );
and \U$15193 ( \24019_24318 , RIdf219d0_1759, \8913_9212 );
and \U$15194 ( \24020_24319 , RIdf1fae0_1737, \8915_9214 );
and \U$15195 ( \24021_24320 , RIdf1b1c0_1685, \8917_9216 );
and \U$15196 ( \24022_24321 , RIdf19438_1664, \8919_9218 );
and \U$15197 ( \24023_24322 , RIdf17278_1640, \8921_9220 );
and \U$15198 ( \24024_24323 , RIdf14578_1608, \8923_9222 );
and \U$15199 ( \24025_24324 , RIdf11878_1576, \8925_9224 );
and \U$15200 ( \24026_24325 , RIdf0eb78_1544, \8927_9226 );
and \U$15201 ( \24027_24326 , RIdf0be78_1512, \8929_9228 );
and \U$15202 ( \24028_24327 , RIdf09178_1480, \8931_9230 );
and \U$15203 ( \24029_24328 , RIdf06478_1448, \8933_9232 );
and \U$15204 ( \24030_24329 , RIdf03778_1416, \8935_9234 );
and \U$15205 ( \24031_24330 , RIdefdd78_1352, \8937_9236 );
and \U$15206 ( \24032_24331 , RIdefb078_1320, \8939_9238 );
and \U$15207 ( \24033_24332 , RIdef8378_1288, \8941_9240 );
and \U$15208 ( \24034_24333 , RIdef5678_1256, \8943_9242 );
and \U$15209 ( \24035_24334 , RIdef2978_1224, \8945_9244 );
and \U$15210 ( \24036_24335 , RIdeefc78_1192, \8947_9246 );
and \U$15211 ( \24037_24336 , RIdeecf78_1160, \8949_9248 );
and \U$15212 ( \24038_24337 , RIdeea278_1128, \8951_9250 );
and \U$15213 ( \24039_24338 , RIfc611a8_6127, \8953_9252 );
and \U$15214 ( \24040_24339 , RIfc61a18_6133, \8955_9254 );
and \U$15215 ( \24041_24340 , RIfca65c8_6915, \8957_9256 );
and \U$15216 ( \24042_24341 , RIfca6b68_6919, \8959_9258 );
and \U$15217 ( \24043_24342 , RIdee4b48_1066, \8961_9260 );
and \U$15218 ( \24044_24343 , RIdee2dc0_1045, \8963_9262 );
and \U$15219 ( \24045_24344 , RIdee0c00_1021, \8965_9264 );
and \U$15220 ( \24046_24345 , RIdedeba8_998, \8967_9266 );
and \U$15221 ( \24047_24346 , RIfc626c0_6142, \8969_9268 );
and \U$15222 ( \24048_24347 , RIfc738f8_6337, \8971_9270 );
and \U$15223 ( \24049_24348 , RIfcb31b0_7060, \8973_9272 );
and \U$15224 ( \24050_24349 , RIee21430_4837, \8975_9274 );
and \U$15225 ( \24051_24350 , RIded9a18_940, \8977_9276 );
and \U$15226 ( \24052_24351 , RIded7588_914, \8979_9278 );
and \U$15227 ( \24053_24352 , RIded5698_892, \8981_9280 );
and \U$15228 ( \24054_24353 , RIded30a0_865, \8983_9282 );
and \U$15229 ( \24055_24354 , RIded0aa8_838, \8985_9284 );
and \U$15230 ( \24056_24355 , RIdecdda8_806, \8987_9286 );
and \U$15231 ( \24057_24356 , RIdecb0a8_774, \8989_9288 );
and \U$15232 ( \24058_24357 , RIdec83a8_742, \8991_9290 );
and \U$15233 ( \24059_24358 , RIdeb48a8_518, \8993_9292 );
and \U$15234 ( \24060_24359 , RIde96fb0_326, \8995_9294 );
and \U$15235 ( \24061_24360 , RIe16e4b0_2632, \8997_9296 );
and \U$15236 ( \24062_24361 , RIe15a2a8_2403, \8999_9298 );
and \U$15237 ( \24063_24362 , RIe143aa8_2147, \9001_9300 );
and \U$15238 ( \24064_24363 , RIdf384a0_2017, \9003_9302 );
and \U$15239 ( \24065_24364 , RIdf2cb00_1885, \9005_9304 );
and \U$15240 ( \24066_24365 , RIdf1d380_1709, \9007_9306 );
and \U$15241 ( \24067_24366 , RIdf00a78_1384, \9009_9308 );
and \U$15242 ( \24068_24367 , RIdee7578_1096, \9011_9310 );
and \U$15243 ( \24069_24368 , RIdedc2e0_969, \9013_9312 );
and \U$15244 ( \24070_24369 , RIde7cef8_199, \9015_9314 );
or \U$15245 ( \24071_24370 , \24007_24306 , \24008_24307 , \24009_24308 , \24010_24309 , \24011_24310 , \24012_24311 , \24013_24312 , \24014_24313 , \24015_24314 , \24016_24315 , \24017_24316 , \24018_24317 , \24019_24318 , \24020_24319 , \24021_24320 , \24022_24321 , \24023_24322 , \24024_24323 , \24025_24324 , \24026_24325 , \24027_24326 , \24028_24327 , \24029_24328 , \24030_24329 , \24031_24330 , \24032_24331 , \24033_24332 , \24034_24333 , \24035_24334 , \24036_24335 , \24037_24336 , \24038_24337 , \24039_24338 , \24040_24339 , \24041_24340 , \24042_24341 , \24043_24342 , \24044_24343 , \24045_24344 , \24046_24345 , \24047_24346 , \24048_24347 , \24049_24348 , \24050_24349 , \24051_24350 , \24052_24351 , \24053_24352 , \24054_24353 , \24055_24354 , \24056_24355 , \24057_24356 , \24058_24357 , \24059_24358 , \24060_24359 , \24061_24360 , \24062_24361 , \24063_24362 , \24064_24363 , \24065_24364 , \24066_24365 , \24067_24366 , \24068_24367 , \24069_24368 , \24070_24369 );
or \U$15246 ( \24072_24371 , \24006_24305 , \24071_24370 );
_DC \g265d/U$1 ( \24073 , \24072_24371 , \9024_9323 );
buf \U$15247 ( \24074_24373 , \24073 );
and \U$15248 ( \24075_24374 , RIe19d940_3170, \9034_9333 );
and \U$15249 ( \24076_24375 , RIe19ac40_3138, \9036_9335 );
and \U$15250 ( \24077_24376 , RIfc64880_6166, \9038_9337 );
and \U$15251 ( \24078_24377 , RIe197f40_3106, \9040_9339 );
and \U$15252 ( \24079_24378 , RIf144848_5239, \9042_9341 );
and \U$15253 ( \24080_24379 , RIe195240_3074, \9044_9343 );
and \U$15254 ( \24081_24380 , RIe192540_3042, \9046_9345 );
and \U$15255 ( \24082_24381 , RIe18f840_3010, \9048_9347 );
and \U$15256 ( \24083_24382 , RIe189e40_2946, \9050_9349 );
and \U$15257 ( \24084_24383 , RIe187140_2914, \9052_9351 );
and \U$15258 ( \24085_24384 , RIf143a38_5229, \9054_9353 );
and \U$15259 ( \24086_24385 , RIe184440_2882, \9056_9355 );
and \U$15260 ( \24087_24386 , RIfc6f140_6286, \9058_9357 );
and \U$15261 ( \24088_24387 , RIe181740_2850, \9060_9359 );
and \U$15262 ( \24089_24388 , RIe17ea40_2818, \9062_9361 );
and \U$15263 ( \24090_24389 , RIe17bd40_2786, \9064_9363 );
and \U$15264 ( \24091_24390 , RIfc64f88_6171, \9066_9365 );
and \U$15265 ( \24092_24391 , RIf141008_5199, \9068_9367 );
and \U$15266 ( \24093_24392 , RIe177150_2732, \9070_9369 );
and \U$15267 ( \24094_24393 , RIfe81738_7817, \9072_9371 );
and \U$15268 ( \24095_24394 , RIfccabf8_7329, \9074_9373 );
and \U$15269 ( \24096_24395 , RIf13f3e8_5179, \9076_9375 );
and \U$15270 ( \24097_24396 , RIfca81e8_6935, \9078_9377 );
and \U$15271 ( \24098_24397 , RIee3d630_5157, \9080_9379 );
and \U$15272 ( \24099_24398 , RIfc66068_6183, \9082_9381 );
and \U$15273 ( \24100_24399 , RIfc6ed08_6283, \9084_9383 );
and \U$15274 ( \24101_24400 , RIfcdde88_7547, \9086_9385 );
and \U$15275 ( \24102_24401 , RIe173a78_2693, \9088_9387 );
and \U$15276 ( \24103_24402 , RIfc66338_6185, \9090_9389 );
and \U$15277 ( \24104_24403 , RIfc6eba0_6282, \9092_9391 );
and \U$15278 ( \24105_24404 , RIfc664a0_6186, \9094_9393 );
and \U$15279 ( \24106_24405 , RIfcacdd8_6989, \9096_9395 );
and \U$15280 ( \24107_24406 , RIfe81468_7815, \9098_9397 );
and \U$15281 ( \24108_24407 , RIe223c98_4697, \9100_9399 );
and \U$15282 ( \24109_24408 , RIfc66d10_6192, \9102_9401 );
and \U$15283 ( \24110_24409 , RIe220f98_4665, \9104_9403 );
and \U$15284 ( \24111_24410 , RIf16b038_5677, \9106_9405 );
and \U$15285 ( \24112_24411 , RIe21e298_4633, \9108_9407 );
and \U$15286 ( \24113_24412 , RIe218898_4569, \9110_9409 );
and \U$15287 ( \24114_24413 , RIe215b98_4537, \9112_9411 );
and \U$15288 ( \24115_24414 , RIfc3fc38_5751, \9114_9413 );
and \U$15289 ( \24116_24415 , RIe212e98_4505, \9116_9415 );
and \U$15290 ( \24117_24416 , RIfc67850_6200, \9118_9417 );
and \U$15291 ( \24118_24417 , RIe210198_4473, \9120_9419 );
and \U$15292 ( \24119_24418 , RIf167f00_5642, \9122_9421 );
and \U$15293 ( \24120_24419 , RIe20d498_4441, \9124_9423 );
and \U$15294 ( \24121_24420 , RIe20a798_4409, \9126_9425 );
and \U$15295 ( \24122_24421 , RIe207a98_4377, \9128_9427 );
and \U$15296 ( \24123_24422 , RIfcacb08_6987, \9130_9429 );
and \U$15297 ( \24124_24423 , RIfcac9a0_6986, \9132_9431 );
and \U$15298 ( \24125_24424 , RIfea8900_8234, \9134_9433 );
and \U$15299 ( \24126_24425 , RIfe818a0_7818, \9136_9435 );
and \U$15300 ( \24127_24426 , RIfca8a58_6941, \9138_9437 );
and \U$15301 ( \24128_24427 , RIfccad60_7330, \9140_9439 );
and \U$15302 ( \24129_24428 , RIfcac838_6985, \9142_9441 );
and \U$15303 ( \24130_24429 , RIfc67418_6197, \9144_9443 );
and \U$15304 ( \24131_24430 , RIf160340_5554, \9146_9445 );
and \U$15305 ( \24132_24431 , RIf15e450_5532, \9148_9447 );
and \U$15306 ( \24133_24432 , RIfe81a08_7819, \9150_9449 );
and \U$15307 ( \24134_24433 , RIfe81300_7814, \9152_9451 );
and \U$15308 ( \24135_24434 , RIfc6dac0_6270, \9154_9453 );
and \U$15309 ( \24136_24435 , RIf15ba20_5502, \9156_9455 );
and \U$15310 ( \24137_24436 , RIfc6d958_6269, \9158_9457 );
and \U$15311 ( \24138_24437 , RIfc6d7f0_6268, \9160_9459 );
or \U$15312 ( \24139_24438 , \24075_24374 , \24076_24375 , \24077_24376 , \24078_24377 , \24079_24378 , \24080_24379 , \24081_24380 , \24082_24381 , \24083_24382 , \24084_24383 , \24085_24384 , \24086_24385 , \24087_24386 , \24088_24387 , \24089_24388 , \24090_24389 , \24091_24390 , \24092_24391 , \24093_24392 , \24094_24393 , \24095_24394 , \24096_24395 , \24097_24396 , \24098_24397 , \24099_24398 , \24100_24399 , \24101_24400 , \24102_24401 , \24103_24402 , \24104_24403 , \24105_24404 , \24106_24405 , \24107_24406 , \24108_24407 , \24109_24408 , \24110_24409 , \24111_24410 , \24112_24411 , \24113_24412 , \24114_24413 , \24115_24414 , \24116_24415 , \24117_24416 , \24118_24417 , \24119_24418 , \24120_24419 , \24121_24420 , \24122_24421 , \24123_24422 , \24124_24423 , \24125_24424 , \24126_24425 , \24127_24426 , \24128_24427 , \24129_24428 , \24130_24429 , \24131_24430 , \24132_24431 , \24133_24432 , \24134_24433 , \24135_24434 , \24136_24435 , \24137_24436 , \24138_24437 );
and \U$15313 ( \24140_24439 , RIfc587d8_6029, \9163_9462 );
and \U$15314 ( \24141_24440 , RIfc6cf80_6262, \9165_9464 );
and \U$15315 ( \24142_24441 , RIfc6d3b8_6265, \9167_9466 );
and \U$15316 ( \24143_24442 , RIfe815d0_7816, \9169_9468 );
and \U$15317 ( \24144_24443 , RIfc6d520_6266, \9171_9470 );
and \U$15318 ( \24145_24444 , RIfcabe60_6978, \9173_9472 );
and \U$15319 ( \24146_24445 , RIfc6d0e8_6263, \9175_9474 );
and \U$15320 ( \24147_24446 , RIe1f5780_4170, \9177_9476 );
and \U$15321 ( \24148_24447 , RIfc6c5a8_6255, \9179_9478 );
and \U$15322 ( \24149_24448 , RIfc68d68_6215, \9181_9480 );
and \U$15323 ( \24150_24449 , RIfc68c00_6214, \9183_9482 );
and \U$15324 ( \24151_24450 , RIe1f3458_4145, \9185_9484 );
and \U$15325 ( \24152_24451 , RIfc68a98_6213, \9187_9486 );
and \U$15326 ( \24153_24452 , RIfccb8a0_7338, \9189_9488 );
and \U$15327 ( \24154_24453 , RIfca9b38_6953, \9191_9490 );
and \U$15328 ( \24155_24454 , RIe1ee160_4086, \9193_9492 );
and \U$15329 ( \24156_24455 , RIe1eba00_4058, \9195_9494 );
and \U$15330 ( \24157_24456 , RIe1e8d00_4026, \9197_9496 );
and \U$15331 ( \24158_24457 , RIe1e6000_3994, \9199_9498 );
and \U$15332 ( \24159_24458 , RIe1e3300_3962, \9201_9500 );
and \U$15333 ( \24160_24459 , RIe1e0600_3930, \9203_9502 );
and \U$15334 ( \24161_24460 , RIe1dd900_3898, \9205_9504 );
and \U$15335 ( \24162_24461 , RIe1dac00_3866, \9207_9506 );
and \U$15336 ( \24163_24462 , RIe1d7f00_3834, \9209_9508 );
and \U$15337 ( \24164_24463 , RIe1d2500_3770, \9211_9510 );
and \U$15338 ( \24165_24464 , RIe1cf800_3738, \9213_9512 );
and \U$15339 ( \24166_24465 , RIe1ccb00_3706, \9215_9514 );
and \U$15340 ( \24167_24466 , RIe1c9e00_3674, \9217_9516 );
and \U$15341 ( \24168_24467 , RIe1c7100_3642, \9219_9518 );
and \U$15342 ( \24169_24468 , RIe1c4400_3610, \9221_9520 );
and \U$15343 ( \24170_24469 , RIe1c1700_3578, \9223_9522 );
and \U$15344 ( \24171_24470 , RIe1bea00_3546, \9225_9524 );
and \U$15345 ( \24172_24471 , RIfc6bbd0_6248, \9227_9526 );
and \U$15346 ( \24173_24472 , RIfcdd348_7539, \9229_9528 );
and \U$15347 ( \24174_24473 , RIe1b9438_3485, \9231_9530 );
and \U$15348 ( \24175_24474 , RIe1b73e0_3462, \9233_9532 );
and \U$15349 ( \24176_24475 , RIfcab5f0_6972, \9235_9534 );
and \U$15350 ( \24177_24476 , RIfccbb70_7340, \9237_9536 );
and \U$15351 ( \24178_24477 , RIe1b5220_3438, \9239_9538 );
and \U$15352 ( \24179_24478 , RIe1b3e70_3424, \9241_9540 );
and \U$15353 ( \24180_24479 , RIfc6c9e0_6258, \9243_9542 );
and \U$15354 ( \24181_24480 , RIfcab488_6971, \9245_9544 );
and \U$15355 ( \24182_24481 , RIfea7dc0_8226, \9247_9546 );
and \U$15356 ( \24183_24482 , RIe1b0bd0_3388, \9249_9548 );
and \U$15357 ( \24184_24483 , RIfc6ce18_6261, \9251_9550 );
and \U$15358 ( \24185_24484 , RIfcabfc8_6979, \9253_9552 );
and \U$15359 ( \24186_24485 , RIe1ac580_3338, \9255_9554 );
and \U$15360 ( \24187_24486 , RIe1aaf00_3322, \9257_9556 );
and \U$15361 ( \24188_24487 , RIe1a8d40_3298, \9259_9558 );
and \U$15362 ( \24189_24488 , RIe1a6040_3266, \9261_9560 );
and \U$15363 ( \24190_24489 , RIe1a3340_3234, \9263_9562 );
and \U$15364 ( \24191_24490 , RIe1a0640_3202, \9265_9564 );
and \U$15365 ( \24192_24491 , RIe18cb40_2978, \9267_9566 );
and \U$15366 ( \24193_24492 , RIe179040_2754, \9269_9568 );
and \U$15367 ( \24194_24493 , RIe226998_4729, \9271_9570 );
and \U$15368 ( \24195_24494 , RIe21b598_4601, \9273_9572 );
and \U$15369 ( \24196_24495 , RIe204d98_4345, \9275_9574 );
and \U$15370 ( \24197_24496 , RIe1fedf8_4277, \9277_9576 );
and \U$15371 ( \24198_24497 , RIe1f81b0_4200, \9279_9578 );
and \U$15372 ( \24199_24498 , RIe1f0cf8_4117, \9281_9580 );
and \U$15373 ( \24200_24499 , RIe1d5200_3802, \9283_9582 );
and \U$15374 ( \24201_24500 , RIe1bbd00_3514, \9285_9584 );
and \U$15375 ( \24202_24501 , RIe1aeb78_3365, \9287_9586 );
and \U$15376 ( \24203_24502 , RIe1711b0_2664, \9289_9588 );
or \U$15377 ( \24204_24503 , \24140_24439 , \24141_24440 , \24142_24441 , \24143_24442 , \24144_24443 , \24145_24444 , \24146_24445 , \24147_24446 , \24148_24447 , \24149_24448 , \24150_24449 , \24151_24450 , \24152_24451 , \24153_24452 , \24154_24453 , \24155_24454 , \24156_24455 , \24157_24456 , \24158_24457 , \24159_24458 , \24160_24459 , \24161_24460 , \24162_24461 , \24163_24462 , \24164_24463 , \24165_24464 , \24166_24465 , \24167_24466 , \24168_24467 , \24169_24468 , \24170_24469 , \24171_24470 , \24172_24471 , \24173_24472 , \24174_24473 , \24175_24474 , \24176_24475 , \24177_24476 , \24178_24477 , \24179_24478 , \24180_24479 , \24181_24480 , \24182_24481 , \24183_24482 , \24184_24483 , \24185_24484 , \24186_24485 , \24187_24486 , \24188_24487 , \24189_24488 , \24190_24489 , \24191_24490 , \24192_24491 , \24193_24492 , \24194_24493 , \24195_24494 , \24196_24495 , \24197_24496 , \24198_24497 , \24199_24498 , \24200_24499 , \24201_24500 , \24202_24501 , \24203_24502 );
or \U$15378 ( \24205_24504 , \24139_24438 , \24204_24503 );
_DC \g378a/U$1 ( \24206 , \24205_24504 , \9298_9597 );
buf \U$15379 ( \24207_24506 , \24206 );
xor \U$15380 ( \24208_24507 , \24074_24373 , \24207_24506 );
and \U$15381 ( \24209_24508 , RIdec5540_709, \8760_9059 );
and \U$15382 ( \24210_24509 , RIdec2840_677, \8762_9061 );
and \U$15383 ( \24211_24510 , RIfcc4dc0_7262, \8764_9063 );
and \U$15384 ( \24212_24511 , RIdebfb40_645, \8766_9065 );
and \U$15385 ( \24213_24512 , RIfc9d7c0_6814, \8768_9067 );
and \U$15386 ( \24214_24513 , RIdebce40_613, \8770_9069 );
and \U$15387 ( \24215_24514 , RIdeba140_581, \8772_9071 );
and \U$15388 ( \24216_24515 , RIdeb7440_549, \8774_9073 );
and \U$15389 ( \24217_24516 , RIfc4d978_5905, \8776_9075 );
and \U$15390 ( \24218_24517 , RIdeb1a40_485, \8778_9077 );
and \U$15391 ( \24219_24518 , RIfc9dbf8_6817, \8780_9079 );
and \U$15392 ( \24220_24519 , RIdeaed40_453, \8782_9081 );
and \U$15393 ( \24221_24520 , RIfcb8610_7120, \8784_9083 );
and \U$15394 ( \24222_24521 , RIdeaa768_421, \8786_9085 );
and \U$15395 ( \24223_24522 , RIdea3e68_389, \8788_9087 );
and \U$15396 ( \24224_24523 , RIde9d568_357, \8790_9089 );
and \U$15397 ( \24225_24524 , RIfc50678_5937, \8792_9091 );
and \U$15398 ( \24226_24525 , RIfc507e0_5938, \8794_9093 );
and \U$15399 ( \24227_24526 , RIfc9dec8_6819, \8796_9095 );
and \U$15400 ( \24228_24527 , RIfc853a0_6538, \8798_9097 );
and \U$15401 ( \24229_24528 , RIde913d0_298, \8800_9099 );
and \U$15402 ( \24230_24529 , RIde8dc08_281, \8802_9101 );
and \U$15403 ( \24231_24530 , RIde89a68_261, \8804_9103 );
and \U$15404 ( \24232_24531 , RIde858c8_241, \8806_9105 );
and \U$15405 ( \24233_24532 , RIde81a70_222, \8808_9107 );
and \U$15406 ( \24234_24533 , RIfc84860_6530, \8810_9109 );
and \U$15407 ( \24235_24534 , RIfc50948_5939, \8812_9111 );
and \U$15408 ( \24236_24535 , RIfc84c98_6533, \8814_9113 );
and \U$15409 ( \24237_24536 , RIfcb7da0_7114, \8816_9115 );
and \U$15410 ( \24238_24537 , RIe16b7b0_2600, \8818_9117 );
and \U$15411 ( \24239_24538 , RIe169b90_2580, \8820_9119 );
and \U$15412 ( \24240_24539 , RIe167e08_2559, \8822_9121 );
and \U$15413 ( \24241_24540 , RIe165540_2530, \8824_9123 );
and \U$15414 ( \24242_24541 , RIe162840_2498, \8826_9125 );
and \U$15415 ( \24243_24542 , RIee37528_5088, \8828_9127 );
and \U$15416 ( \24244_24543 , RIe15fb40_2466, \8830_9129 );
and \U$15417 ( \24245_24544 , RIfcb5be0_7090, \8832_9131 );
and \U$15418 ( \24246_24545 , RIe15ce40_2434, \8834_9133 );
and \U$15419 ( \24247_24546 , RIe157440_2370, \8836_9135 );
and \U$15420 ( \24248_24547 , RIe154740_2338, \8838_9137 );
and \U$15421 ( \24249_24548 , RIfcd35c8_7427, \8840_9139 );
and \U$15422 ( \24250_24549 , RIe151a40_2306, \8842_9141 );
and \U$15423 ( \24251_24550 , RIfc53a80_5974, \8844_9143 );
and \U$15424 ( \24252_24551 , RIe14ed40_2274, \8846_9145 );
and \U$15425 ( \24253_24552 , RIfcc6170_7276, \8848_9147 );
and \U$15426 ( \24254_24553 , RIe14c040_2242, \8850_9149 );
and \U$15427 ( \24255_24554 , RIe149340_2210, \8852_9151 );
and \U$15428 ( \24256_24555 , RIe146640_2178, \8854_9153 );
and \U$15429 ( \24257_24556 , RIfc7f130_6468, \8856_9155 );
and \U$15430 ( \24258_24557 , RIee33310_5041, \8858_9157 );
and \U$15431 ( \24259_24558 , RIfcb4f38_7081, \8860_9159 );
and \U$15432 ( \24260_24559 , RIfc47f78_5841, \8862_9161 );
and \U$15433 ( \24261_24560 , RIe140f10_2116, \8864_9163 );
and \U$15434 ( \24262_24561 , RIdf3ee18_2092, \8866_9165 );
and \U$15435 ( \24263_24562 , RIdf3cc58_2068, \8868_9167 );
and \U$15436 ( \24264_24563 , RIdf3a7c8_2042, \8870_9169 );
and \U$15437 ( \24265_24564 , RIfc7fc70_6476, \8872_9171 );
and \U$15438 ( \24266_24565 , RIfcd27b8_7417, \8874_9173 );
and \U$15439 ( \24267_24566 , RIfca1000_6854, \8876_9175 );
and \U$15440 ( \24268_24567 , RIfcc6b48_7283, \8878_9177 );
and \U$15441 ( \24269_24568 , RIdf35908_1986, \8880_9179 );
and \U$15442 ( \24270_24569 , RIdf33478_1960, \8882_9181 );
and \U$15443 ( \24271_24570 , RIfebe9f8_8289, \8884_9183 );
and \U$15444 ( \24272_24571 , RIdf2f260_1913, \8886_9185 );
or \U$15445 ( \24273_24572 , \24209_24508 , \24210_24509 , \24211_24510 , \24212_24511 , \24213_24512 , \24214_24513 , \24215_24514 , \24216_24515 , \24217_24516 , \24218_24517 , \24219_24518 , \24220_24519 , \24221_24520 , \24222_24521 , \24223_24522 , \24224_24523 , \24225_24524 , \24226_24525 , \24227_24526 , \24228_24527 , \24229_24528 , \24230_24529 , \24231_24530 , \24232_24531 , \24233_24532 , \24234_24533 , \24235_24534 , \24236_24535 , \24237_24536 , \24238_24537 , \24239_24538 , \24240_24539 , \24241_24540 , \24242_24541 , \24243_24542 , \24244_24543 , \24245_24544 , \24246_24545 , \24247_24546 , \24248_24547 , \24249_24548 , \24250_24549 , \24251_24550 , \24252_24551 , \24253_24552 , \24254_24553 , \24255_24554 , \24256_24555 , \24257_24556 , \24258_24557 , \24259_24558 , \24260_24559 , \24261_24560 , \24262_24561 , \24263_24562 , \24264_24563 , \24265_24564 , \24266_24565 , \24267_24566 , \24268_24567 , \24269_24568 , \24270_24569 , \24271_24570 , \24272_24571 );
and \U$15446 ( \24274_24573 , RIfcb7968_7111, \8889_9188 );
and \U$15447 ( \24275_24574 , RIee2a3a0_4939, \8891_9190 );
and \U$15448 ( \24276_24575 , RIfc51050_5944, \8893_9192 );
and \U$15449 ( \24277_24576 , RIfcd3fa0_7434, \8895_9194 );
and \U$15450 ( \24278_24577 , RIdf2a3a0_1857, \8897_9196 );
and \U$15451 ( \24279_24578 , RIdf28078_1832, \8899_9198 );
and \U$15452 ( \24280_24579 , RIfe81198_7813, \8901_9200 );
and \U$15453 ( \24281_24580 , RIdf24838_1792, \8903_9202 );
and \U$15454 ( \24282_24581 , RIfc84428_6527, \8905_9204 );
and \U$15455 ( \24283_24582 , RIfce7ed8_7661, \8907_9206 );
and \U$15456 ( \24284_24583 , RIdf22d80_1773, \8909_9208 );
and \U$15457 ( \24285_24584 , RIfc515f0_5948, \8911_9210 );
and \U$15458 ( \24286_24585 , RIdf21868_1758, \8913_9212 );
and \U$15459 ( \24287_24586 , RIdf1f978_1736, \8915_9214 );
and \U$15460 ( \24288_24587 , RIdf1b058_1684, \8917_9216 );
and \U$15461 ( \24289_24588 , RIdf192d0_1663, \8919_9218 );
and \U$15462 ( \24290_24589 , RIdf17110_1639, \8921_9220 );
and \U$15463 ( \24291_24590 , RIdf14410_1607, \8923_9222 );
and \U$15464 ( \24292_24591 , RIdf11710_1575, \8925_9224 );
and \U$15465 ( \24293_24592 , RIdf0ea10_1543, \8927_9226 );
and \U$15466 ( \24294_24593 , RIdf0bd10_1511, \8929_9228 );
and \U$15467 ( \24295_24594 , RIdf09010_1479, \8931_9230 );
and \U$15468 ( \24296_24595 , RIdf06310_1447, \8933_9232 );
and \U$15469 ( \24297_24596 , RIdf03610_1415, \8935_9234 );
and \U$15470 ( \24298_24597 , RIdefdc10_1351, \8937_9236 );
and \U$15471 ( \24299_24598 , RIdefaf10_1319, \8939_9238 );
and \U$15472 ( \24300_24599 , RIdef8210_1287, \8941_9240 );
and \U$15473 ( \24301_24600 , RIdef5510_1255, \8943_9242 );
and \U$15474 ( \24302_24601 , RIdef2810_1223, \8945_9244 );
and \U$15475 ( \24303_24602 , RIdeefb10_1191, \8947_9246 );
and \U$15476 ( \24304_24603 , RIdeece10_1159, \8949_9248 );
and \U$15477 ( \24305_24604 , RIdeea110_1127, \8951_9250 );
and \U$15478 ( \24306_24605 , RIfc7e1b8_6457, \8953_9252 );
and \U$15479 ( \24307_24606 , RIfca19d8_6861, \8955_9254 );
and \U$15480 ( \24308_24607 , RIfc7dab0_6452, \8957_9256 );
and \U$15481 ( \24309_24608 , RIfc7e488_6459, \8959_9258 );
and \U$15482 ( \24310_24609 , RIdee49e0_1065, \8961_9260 );
and \U$15483 ( \24311_24610 , RIfe80d60_7810, \8963_9262 );
and \U$15484 ( \24312_24611 , RIfeabba0_8270, \8965_9264 );
and \U$15485 ( \24313_24612 , RIfe80bf8_7809, \8967_9266 );
and \U$15486 ( \24314_24613 , RIfcb3750_7064, \8969_9268 );
and \U$15487 ( \24315_24614 , RIfce9f30_7684, \8971_9270 );
and \U$15488 ( \24316_24615 , RIfc7e5f0_6460, \8973_9272 );
and \U$15489 ( \24317_24616 , RIfc56a50_6008, \8975_9274 );
and \U$15490 ( \24318_24617 , RIfe81030_7812, \8977_9276 );
and \U$15491 ( \24319_24618 , RIded7420_913, \8979_9278 );
and \U$15492 ( \24320_24619 , RIfe80ec8_7811, \8981_9280 );
and \U$15493 ( \24321_24620 , RIded2f38_864, \8983_9282 );
and \U$15494 ( \24322_24621 , RIded0940_837, \8985_9284 );
and \U$15495 ( \24323_24622 , RIdecdc40_805, \8987_9286 );
and \U$15496 ( \24324_24623 , RIdecaf40_773, \8989_9288 );
and \U$15497 ( \24325_24624 , RIdec8240_741, \8991_9290 );
and \U$15498 ( \24326_24625 , RIdeb4740_517, \8993_9292 );
and \U$15499 ( \24327_24626 , RIde96c68_325, \8995_9294 );
and \U$15500 ( \24328_24627 , RIe16e348_2631, \8997_9296 );
and \U$15501 ( \24329_24628 , RIe15a140_2402, \8999_9298 );
and \U$15502 ( \24330_24629 , RIe143940_2146, \9001_9300 );
and \U$15503 ( \24331_24630 , RIdf38338_2016, \9003_9302 );
and \U$15504 ( \24332_24631 , RIdf2c998_1884, \9005_9304 );
and \U$15505 ( \24333_24632 , RIdf1d218_1708, \9007_9306 );
and \U$15506 ( \24334_24633 , RIdf00910_1383, \9009_9308 );
and \U$15507 ( \24335_24634 , RIdee7410_1095, \9011_9310 );
and \U$15508 ( \24336_24635 , RIdedc178_968, \9013_9312 );
and \U$15509 ( \24337_24636 , RIde7cbb0_198, \9015_9314 );
or \U$15510 ( \24338_24637 , \24274_24573 , \24275_24574 , \24276_24575 , \24277_24576 , \24278_24577 , \24279_24578 , \24280_24579 , \24281_24580 , \24282_24581 , \24283_24582 , \24284_24583 , \24285_24584 , \24286_24585 , \24287_24586 , \24288_24587 , \24289_24588 , \24290_24589 , \24291_24590 , \24292_24591 , \24293_24592 , \24294_24593 , \24295_24594 , \24296_24595 , \24297_24596 , \24298_24597 , \24299_24598 , \24300_24599 , \24301_24600 , \24302_24601 , \24303_24602 , \24304_24603 , \24305_24604 , \24306_24605 , \24307_24606 , \24308_24607 , \24309_24608 , \24310_24609 , \24311_24610 , \24312_24611 , \24313_24612 , \24314_24613 , \24315_24614 , \24316_24615 , \24317_24616 , \24318_24617 , \24319_24618 , \24320_24619 , \24321_24620 , \24322_24621 , \24323_24622 , \24324_24623 , \24325_24624 , \24326_24625 , \24327_24626 , \24328_24627 , \24329_24628 , \24330_24629 , \24331_24630 , \24332_24631 , \24333_24632 , \24334_24633 , \24335_24634 , \24336_24635 , \24337_24636 );
or \U$15511 ( \24339_24638 , \24273_24572 , \24338_24637 );
_DC \g26e2/U$1 ( \24340 , \24339_24638 , \9024_9323 );
buf \U$15512 ( \24341_24640 , \24340 );
and \U$15513 ( \24342_24641 , RIe19d7d8_3169, \9034_9333 );
and \U$15514 ( \24343_24642 , RIe19aad8_3137, \9036_9335 );
and \U$15515 ( \24344_24643 , RIfcc2d68_7239, \9038_9337 );
and \U$15516 ( \24345_24644 , RIe197dd8_3105, \9040_9339 );
and \U$15517 ( \24346_24645 , RIfc5c5b8_6073, \9042_9341 );
and \U$15518 ( \24347_24646 , RIe1950d8_3073, \9044_9343 );
and \U$15519 ( \24348_24647 , RIe1923d8_3041, \9046_9345 );
and \U$15520 ( \24349_24648 , RIe18f6d8_3009, \9048_9347 );
and \U$15521 ( \24350_24649 , RIe189cd8_2945, \9050_9349 );
and \U$15522 ( \24351_24650 , RIe186fd8_2913, \9052_9351 );
and \U$15523 ( \24352_24651 , RIf1438d0_5228, \9054_9353 );
and \U$15524 ( \24353_24652 , RIe1842d8_2881, \9056_9355 );
and \U$15525 ( \24354_24653 , RIfc5b370_6060, \9058_9357 );
and \U$15526 ( \24355_24654 , RIe1815d8_2849, \9060_9359 );
and \U$15527 ( \24356_24655 , RIe17e8d8_2817, \9062_9361 );
and \U$15528 ( \24357_24656 , RIe17bbd8_2785, \9064_9363 );
and \U$15529 ( \24358_24657 , RIfcbb748_7155, \9066_9365 );
and \U$15530 ( \24359_24658 , RIfc59480_6038, \9068_9367 );
and \U$15531 ( \24360_24659 , RIfcbbce8_7159, \9070_9369 );
and \U$15532 ( \24361_24660 , RIe175c38_2717, \9072_9371 );
and \U$15533 ( \24362_24661 , RIfcdb890_7520, \9074_9373 );
and \U$15534 ( \24363_24662 , RIfc59b88_6043, \9076_9375 );
and \U$15535 ( \24364_24663 , RIfc8ada0_6602, \9078_9377 );
and \U$15536 ( \24365_24664 , RIfcb5eb0_7092, \9080_9379 );
and \U$15537 ( \24366_24665 , RIfc57c98_6021, \9082_9381 );
and \U$15538 ( \24367_24666 , RIfc57158_6013, \9084_9383 );
and \U$15539 ( \24368_24667 , RIfc58aa8_6031, \9086_9385 );
and \U$15540 ( \24369_24668 , RIe173910_2692, \9088_9387 );
and \U$15541 ( \24370_24669 , RIfcc62d8_7277, \9090_9389 );
and \U$15542 ( \24371_24670 , RIfc8a968_6599, \9092_9391 );
and \U$15543 ( \24372_24671 , RIfc57428_6015, \9094_9393 );
and \U$15544 ( \24373_24672 , RIfc56d20_6010, \9096_9395 );
and \U$15545 ( \24374_24673 , RIfc408e0_5760, \9098_9397 );
and \U$15546 ( \24375_24674 , RIe223b30_4696, \9100_9399 );
and \U$15547 ( \24376_24675 , RIfc82970_6508, \9102_9401 );
and \U$15548 ( \24377_24676 , RIe220e30_4664, \9104_9403 );
and \U$15549 ( \24378_24677 , RIfcecc30_7716, \9106_9405 );
and \U$15550 ( \24379_24678 , RIe21e130_4632, \9108_9407 );
and \U$15551 ( \24380_24679 , RIe218730_4568, \9110_9409 );
and \U$15552 ( \24381_24680 , RIe215a30_4536, \9112_9411 );
and \U$15553 ( \24382_24681 , RIfc3fad0_5750, \9114_9413 );
and \U$15554 ( \24383_24682 , RIe212d30_4504, \9116_9415 );
and \U$15555 ( \24384_24683 , RIf169148_5655, \9118_9417 );
and \U$15556 ( \24385_24684 , RIe210030_4472, \9120_9419 );
and \U$15557 ( \24386_24685 , RIfc545c0_5982, \9122_9421 );
and \U$15558 ( \24387_24686 , RIe20d330_4440, \9124_9423 );
and \U$15559 ( \24388_24687 , RIe20a630_4408, \9126_9425 );
and \U$15560 ( \24389_24688 , RIe207930_4376, \9128_9427 );
and \U$15561 ( \24390_24689 , RIfc88d48_6579, \9130_9429 );
and \U$15562 ( \24391_24690 , RIfc4bec0_5886, \9132_9431 );
and \U$15563 ( \24392_24691 , RIe202638_4317, \9134_9433 );
and \U$15564 ( \24393_24692 , RIe200b80_4298, \9136_9435 );
and \U$15565 ( \24394_24693 , RIfc88910_6576, \9138_9437 );
and \U$15566 ( \24395_24694 , RIfc4c190_5888, \9140_9439 );
and \U$15567 ( \24396_24695 , RIfc4c2f8_5889, \9142_9441 );
and \U$15568 ( \24397_24696 , RIfcba398_7141, \9144_9443 );
and \U$15569 ( \24398_24697 , RIfcd4270_7436, \9146_9445 );
and \U$15570 ( \24399_24698 , RIfcba0c8_7139, \9148_9447 );
and \U$15571 ( \24400_24699 , RIe1fcda0_4254, \9150_9449 );
and \U$15572 ( \24401_24700 , RIe1fbb58_4241, \9152_9451 );
and \U$15573 ( \24402_24701 , RIfc53d50_5976, \9154_9453 );
and \U$15574 ( \24403_24702 , RIfc9b768_6791, \9156_9455 );
and \U$15575 ( \24404_24703 , RIfc537b0_5972, \9158_9457 );
and \U$15576 ( \24405_24704 , RIfc4c5c8_5891, \9160_9459 );
or \U$15577 ( \24406_24705 , \24342_24641 , \24343_24642 , \24344_24643 , \24345_24644 , \24346_24645 , \24347_24646 , \24348_24647 , \24349_24648 , \24350_24649 , \24351_24650 , \24352_24651 , \24353_24652 , \24354_24653 , \24355_24654 , \24356_24655 , \24357_24656 , \24358_24657 , \24359_24658 , \24360_24659 , \24361_24660 , \24362_24661 , \24363_24662 , \24364_24663 , \24365_24664 , \24366_24665 , \24367_24666 , \24368_24667 , \24369_24668 , \24370_24669 , \24371_24670 , \24372_24671 , \24373_24672 , \24374_24673 , \24375_24674 , \24376_24675 , \24377_24676 , \24378_24677 , \24379_24678 , \24380_24679 , \24381_24680 , \24382_24681 , \24383_24682 , \24384_24683 , \24385_24684 , \24386_24685 , \24387_24686 , \24388_24687 , \24389_24688 , \24390_24689 , \24391_24690 , \24392_24691 , \24393_24692 , \24394_24693 , \24395_24694 , \24396_24695 , \24397_24696 , \24398_24697 , \24399_24698 , \24400_24699 , \24401_24700 , \24402_24701 , \24403_24702 , \24404_24703 , \24405_24704 );
and \U$15578 ( \24407_24706 , RIfc9e468_6823, \9163_9462 );
and \U$15579 ( \24408_24707 , RIf157da8_5459, \9165_9464 );
and \U$15580 ( \24409_24708 , RIfcb9f60_7138, \9167_9466 );
and \U$15581 ( \24410_24709 , RIe1fa208_4223, \9169_9468 );
and \U$15582 ( \24411_24710 , RIfc849c8_6531, \9171_9470 );
and \U$15583 ( \24412_24711 , RIfc529a0_5962, \9173_9472 );
and \U$15584 ( \24413_24712 , RIfc9f6b0_6836, \9175_9474 );
and \U$15585 ( \24414_24713 , RIe1f5618_4169, \9177_9476 );
and \U$15586 ( \24415_24714 , RIf153320_5406, \9179_9478 );
and \U$15587 ( \24416_24715 , RIfcc4988_7259, \9181_9480 );
and \U$15588 ( \24417_24716 , RIf150d28_5379, \9183_9482 );
and \U$15589 ( \24418_24717 , RIfebe458_8285, \9185_9484 );
and \U$15590 ( \24419_24718 , RIfc87f38_6569, \9187_9486 );
and \U$15591 ( \24420_24719 , RIfcb7f08_7115, \9189_9488 );
and \U$15592 ( \24421_24720 , RIf14e190_5348, \9191_9490 );
and \U$15593 ( \24422_24721 , RIfe80658_7805, \9193_9492 );
and \U$15594 ( \24423_24722 , RIe1eb898_4057, \9195_9494 );
and \U$15595 ( \24424_24723 , RIe1e8b98_4025, \9197_9496 );
and \U$15596 ( \24425_24724 , RIe1e5e98_3993, \9199_9498 );
and \U$15597 ( \24426_24725 , RIe1e3198_3961, \9201_9500 );
and \U$15598 ( \24427_24726 , RIe1e0498_3929, \9203_9502 );
and \U$15599 ( \24428_24727 , RIe1dd798_3897, \9205_9504 );
and \U$15600 ( \24429_24728 , RIe1daa98_3865, \9207_9506 );
and \U$15601 ( \24430_24729 , RIe1d7d98_3833, \9209_9508 );
and \U$15602 ( \24431_24730 , RIe1d2398_3769, \9211_9510 );
and \U$15603 ( \24432_24731 , RIe1cf698_3737, \9213_9512 );
and \U$15604 ( \24433_24732 , RIe1cc998_3705, \9215_9514 );
and \U$15605 ( \24434_24733 , RIe1c9c98_3673, \9217_9516 );
and \U$15606 ( \24435_24734 , RIe1c6f98_3641, \9219_9518 );
and \U$15607 ( \24436_24735 , RIe1c4298_3609, \9221_9520 );
and \U$15608 ( \24437_24736 , RIe1c1598_3577, \9223_9522 );
and \U$15609 ( \24438_24737 , RIe1be898_3545, \9225_9524 );
and \U$15610 ( \24439_24738 , RIf14cc78_5333, \9227_9526 );
and \U$15611 ( \24440_24739 , RIf14ba30_5320, \9229_9528 );
and \U$15612 ( \24441_24740 , RIe1b92d0_3484, \9231_9530 );
and \U$15613 ( \24442_24741 , RIe1b7278_3461, \9233_9532 );
and \U$15614 ( \24443_24742 , RIf14a7e8_5307, \9235_9534 );
and \U$15615 ( \24444_24743 , RIf149ca8_5299, \9237_9536 );
and \U$15616 ( \24445_24744 , RIfebe5c0_8286, \9239_9538 );
and \U$15617 ( \24446_24745 , RIfe807c0_7806, \9241_9540 );
and \U$15618 ( \24447_24746 , RIfc50510_5936, \9243_9542 );
and \U$15619 ( \24448_24747 , RIfce4f08_7627, \9245_9544 );
and \U$15620 ( \24449_24748 , RIfe80a90_7808, \9247_9546 );
and \U$15621 ( \24450_24749 , RIfebe890_8288, \9249_9548 );
and \U$15622 ( \24451_24750 , RIfc9cde8_6807, \9251_9550 );
and \U$15623 ( \24452_24751 , RIfc87560_6562, \9253_9552 );
and \U$15624 ( \24453_24752 , RIfe80928_7807, \9255_9554 );
and \U$15625 ( \24454_24753 , RIfebe728_8287, \9257_9556 );
and \U$15626 ( \24455_24754 , RIe1a8bd8_3297, \9259_9558 );
and \U$15627 ( \24456_24755 , RIe1a5ed8_3265, \9261_9560 );
and \U$15628 ( \24457_24756 , RIe1a31d8_3233, \9263_9562 );
and \U$15629 ( \24458_24757 , RIe1a04d8_3201, \9265_9564 );
and \U$15630 ( \24459_24758 , RIe18c9d8_2977, \9267_9566 );
and \U$15631 ( \24460_24759 , RIe178ed8_2753, \9269_9568 );
and \U$15632 ( \24461_24760 , RIe226830_4728, \9271_9570 );
and \U$15633 ( \24462_24761 , RIe21b430_4600, \9273_9572 );
and \U$15634 ( \24463_24762 , RIe204c30_4344, \9275_9574 );
and \U$15635 ( \24464_24763 , RIe1fec90_4276, \9277_9576 );
and \U$15636 ( \24465_24764 , RIe1f8048_4199, \9279_9578 );
and \U$15637 ( \24466_24765 , RIe1f0b90_4116, \9281_9580 );
and \U$15638 ( \24467_24766 , RIe1d5098_3801, \9283_9582 );
and \U$15639 ( \24468_24767 , RIe1bbb98_3513, \9285_9584 );
and \U$15640 ( \24469_24768 , RIe1aea10_3364, \9287_9586 );
and \U$15641 ( \24470_24769 , RIe171048_2663, \9289_9588 );
or \U$15642 ( \24471_24770 , \24407_24706 , \24408_24707 , \24409_24708 , \24410_24709 , \24411_24710 , \24412_24711 , \24413_24712 , \24414_24713 , \24415_24714 , \24416_24715 , \24417_24716 , \24418_24717 , \24419_24718 , \24420_24719 , \24421_24720 , \24422_24721 , \24423_24722 , \24424_24723 , \24425_24724 , \24426_24725 , \24427_24726 , \24428_24727 , \24429_24728 , \24430_24729 , \24431_24730 , \24432_24731 , \24433_24732 , \24434_24733 , \24435_24734 , \24436_24735 , \24437_24736 , \24438_24737 , \24439_24738 , \24440_24739 , \24441_24740 , \24442_24741 , \24443_24742 , \24444_24743 , \24445_24744 , \24446_24745 , \24447_24746 , \24448_24747 , \24449_24748 , \24450_24749 , \24451_24750 , \24452_24751 , \24453_24752 , \24454_24753 , \24455_24754 , \24456_24755 , \24457_24756 , \24458_24757 , \24459_24758 , \24460_24759 , \24461_24760 , \24462_24761 , \24463_24762 , \24464_24763 , \24465_24764 , \24466_24765 , \24467_24766 , \24468_24767 , \24469_24768 , \24470_24769 );
or \U$15643 ( \24472_24771 , \24406_24705 , \24471_24770 );
_DC \g380f/U$1 ( \24473 , \24472_24771 , \9298_9597 );
buf \U$15644 ( \24474_24773 , \24473 );
and \U$15645 ( \24475_24774 , \24341_24640 , \24474_24773 );
and \U$15646 ( \24476_24775 , \22483_22782 , \22616_22915 );
and \U$15647 ( \24477_24776 , \22616_22915 , \22891_23190 );
and \U$15648 ( \24478_24777 , \22483_22782 , \22891_23190 );
or \U$15649 ( \24479_24778 , \24476_24775 , \24477_24776 , \24478_24777 );
and \U$15650 ( \24480_24779 , \24474_24773 , \24479_24778 );
and \U$15651 ( \24481_24780 , \24341_24640 , \24479_24778 );
or \U$15652 ( \24482_24781 , \24475_24774 , \24480_24779 , \24481_24780 );
xor \U$15653 ( \24483_24782 , \24208_24507 , \24482_24781 );
buf g4412_GF_PartitionCandidate( \24484_24783_nG4412 , \24483_24782 );
xor \U$15654 ( \24485_24784 , \24341_24640 , \24474_24773 );
xor \U$15655 ( \24486_24785 , \24485_24784 , \24479_24778 );
buf g4415_GF_PartitionCandidate( \24487_24786_nG4415 , \24486_24785 );
nand \U$15656 ( \24488_24787 , \24487_24786_nG4415 , \22893_23192_nG4418 );
and \U$15657 ( \24489_24788 , \24484_24783_nG4412 , \24488_24787 );
xor \U$15658 ( \24490_24789 , \24487_24786_nG4415 , \22893_23192_nG4418 );
and \U$15663 ( \24491_24793 , \24490_24789 , \10392_10694_nG9c0e );
or \U$15664 ( \24492_24794 , 1'b0 , \24491_24793 );
xor \U$15665 ( \24493_24795 , \24489_24788 , \24492_24794 );
xor \U$15666 ( \24494_24796 , \24489_24788 , \24493_24795 );
buf \U$15667 ( \24495_24797 , \24494_24796 );
buf \U$15668 ( \24496_24798 , \24495_24797 );
xor \U$15669 ( \24497_24799 , \23941_24240 , \24496_24798 );
and \U$15670 ( \24498_24800 , \23434_23736 , \23439_23741 );
and \U$15671 ( \24499_24801 , \23434_23736 , \23445_23747 );
and \U$15672 ( \24500_24802 , \23439_23741 , \23445_23747 );
or \U$15673 ( \24501_24803 , \24498_24800 , \24499_24801 , \24500_24802 );
buf \U$15674 ( \24502_24804 , \24501_24803 );
and \U$15675 ( \24503_24805 , \23527_23826 , \23533_23832 );
and \U$15676 ( \24504_24806 , \23527_23826 , \23540_23839 );
and \U$15677 ( \24505_24807 , \23533_23832 , \23540_23839 );
or \U$15678 ( \24506_24808 , \24503_24805 , \24504_24806 , \24505_24807 );
buf \U$15679 ( \24507_24809 , \24506_24808 );
and \U$15680 ( \24508_24810 , \23503_23802 , \23509_23808 );
and \U$15681 ( \24509_24811 , \23503_23802 , \23516_23815 );
and \U$15682 ( \24510_24812 , \23509_23808 , \23516_23815 );
or \U$15683 ( \24511_24813 , \24508_24810 , \24509_24811 , \24510_24812 );
buf \U$15684 ( \24512_24814 , \24511_24813 );
and \U$15685 ( \24513_24815 , \23495_23201 , \10693_10995_nG9c0b );
and \U$15686 ( \24514_24816 , \22899_23198 , \10981_11283_nG9c08 );
or \U$15687 ( \24515_24817 , \24513_24815 , \24514_24816 );
xor \U$15688 ( \24516_24818 , \22898_23197 , \24515_24817 );
buf \U$15689 ( \24517_24819 , \24516_24818 );
buf \U$15691 ( \24518_24820 , \24517_24819 );
and \U$15692 ( \24519_24821 , \21908_21658 , \11299_11598_nG9c05 );
and \U$15693 ( \24520_24822 , \21356_21655 , \12168_12470_nG9c02 );
or \U$15694 ( \24521_24823 , \24519_24821 , \24520_24822 );
xor \U$15695 ( \24522_24824 , \21355_21654 , \24521_24823 );
buf \U$15696 ( \24523_24825 , \24522_24824 );
buf \U$15698 ( \24524_24826 , \24523_24825 );
xor \U$15699 ( \24525_24827 , \24518_24820 , \24524_24826 );
buf \U$15700 ( \24526_24828 , \24525_24827 );
xor \U$15701 ( \24527_24829 , \24512_24814 , \24526_24828 );
and \U$15702 ( \24528_24830 , \17437_17297 , \15074_15373_nG9bf3 );
and \U$15703 ( \24529_24831 , \16995_17294 , \16013_16315_nG9bf0 );
or \U$15704 ( \24530_24832 , \24528_24830 , \24529_24831 );
xor \U$15705 ( \24531_24833 , \16994_17293 , \24530_24832 );
buf \U$15706 ( \24532_24834 , \24531_24833 );
buf \U$15708 ( \24533_24835 , \24532_24834 );
xor \U$15709 ( \24534_24836 , \24527_24829 , \24533_24835 );
buf \U$15710 ( \24535_24837 , \24534_24836 );
and \U$15711 ( \24536_24838 , \23460_23762 , \23466_23768 );
and \U$15712 ( \24537_24839 , \23460_23762 , \23473_23775 );
and \U$15713 ( \24538_24840 , \23466_23768 , \23473_23775 );
or \U$15714 ( \24539_24841 , \24536_24838 , \24537_24839 , \24538_24840 );
buf \U$15715 ( \24540_24842 , \24539_24841 );
xor \U$15716 ( \24541_24843 , \24535_24837 , \24540_24842 );
and \U$15717 ( \24542_24844 , \12183_12157 , \20787_21086_nG9bdb );
and \U$15718 ( \24543_24845 , \11855_12154 , \21827_22129_nG9bd8 );
or \U$15719 ( \24544_24846 , \24542_24844 , \24543_24845 );
xor \U$15720 ( \24545_24847 , \11854_12153 , \24544_24846 );
buf \U$15721 ( \24546_24848 , \24545_24847 );
buf \U$15723 ( \24547_24849 , \24546_24848 );
xor \U$15724 ( \24548_24850 , \24541_24843 , \24547_24849 );
buf \U$15725 ( \24549_24851 , \24548_24850 );
xor \U$15726 ( \24550_24852 , \24507_24809 , \24549_24851 );
and \U$15727 ( \24551_24853 , \23458_23760 , \23475_23777 );
and \U$15728 ( \24552_24854 , \23458_23760 , \23482_23784 );
and \U$15729 ( \24553_24855 , \23475_23777 , \23482_23784 );
or \U$15730 ( \24554_24856 , \24551_24853 , \24552_24854 , \24553_24855 );
buf \U$15731 ( \24555_24857 , \24554_24856 );
and \U$15732 ( \24556_24858 , \23489_23791 , \23518_23817 );
and \U$15733 ( \24557_24859 , \23489_23791 , \23525_23824 );
and \U$15734 ( \24558_24860 , \23518_23817 , \23525_23824 );
or \U$15735 ( \24559_24861 , \24556_24858 , \24557_24859 , \24558_24860 );
buf \U$15736 ( \24560_24862 , \24559_24861 );
xor \U$15737 ( \24561_24863 , \24555_24857 , \24560_24862 );
and \U$15738 ( \24562_24864 , \13431_13370 , \19287_19586_nG9be1 );
and \U$15739 ( \24563_24865 , \13068_13367 , \20306_20608_nG9bde );
or \U$15740 ( \24564_24866 , \24562_24864 , \24563_24865 );
xor \U$15741 ( \24565_24867 , \13067_13366 , \24564_24866 );
buf \U$15742 ( \24566_24868 , \24565_24867 );
buf \U$15744 ( \24567_24869 , \24566_24868 );
xor \U$15745 ( \24568_24870 , \24561_24863 , \24567_24869 );
buf \U$15746 ( \24569_24871 , \24568_24870 );
xor \U$15747 ( \24570_24872 , \24550_24852 , \24569_24871 );
buf \U$15748 ( \24571_24873 , \24570_24872 );
xor \U$15749 ( \24572_24874 , \24502_24804 , \24571_24873 );
and \U$15750 ( \24573_24875 , \23420_23722 , \23425_23727 );
and \U$15751 ( \24574_24876 , \23420_23722 , \23432_23734 );
and \U$15752 ( \24575_24877 , \23425_23727 , \23432_23734 );
or \U$15753 ( \24576_24878 , \24573_24875 , \24574_24876 , \24575_24877 );
buf \U$15754 ( \24577_24879 , \24576_24878 );
and \U$15755 ( \24578_24880 , \23492_23794 , \23501_23800 );
buf \U$15756 ( \24579_24881 , \24578_24880 );
and \U$15757 ( \24580_24882 , \20353_20155 , \12502_12801_nG9bff );
and \U$15758 ( \24581_24883 , \19853_20152 , \13403_13705_nG9bfc );
or \U$15759 ( \24582_24884 , \24580_24882 , \24581_24883 );
xor \U$15760 ( \24583_24885 , \19852_20151 , \24582_24884 );
buf \U$15761 ( \24584_24886 , \24583_24885 );
buf \U$15763 ( \24585_24887 , \24584_24886 );
xor \U$15764 ( \24586_24888 , \24579_24881 , \24585_24887 );
and \U$15765 ( \24587_24889 , \18908_18702 , \13771_14070_nG9bf9 );
and \U$15766 ( \24588_24890 , \18400_18699 , \14682_14984_nG9bf6 );
or \U$15767 ( \24589_24891 , \24587_24889 , \24588_24890 );
xor \U$15768 ( \24590_24892 , \18399_18698 , \24589_24891 );
buf \U$15769 ( \24591_24893 , \24590_24892 );
buf \U$15771 ( \24592_24894 , \24591_24893 );
xor \U$15772 ( \24593_24895 , \24586_24888 , \24592_24894 );
buf \U$15773 ( \24594_24896 , \24593_24895 );
and \U$15774 ( \24595_24897 , \16405_15940 , \16378_16680_nG9bed );
and \U$15775 ( \24596_24898 , \15638_15937 , \17363_17665_nG9bea );
or \U$15776 ( \24597_24899 , \24595_24897 , \24596_24898 );
xor \U$15777 ( \24598_24900 , \15637_15936 , \24597_24899 );
buf \U$15778 ( \24599_24901 , \24598_24900 );
buf \U$15780 ( \24600_24902 , \24599_24901 );
xor \U$15781 ( \24601_24903 , \24594_24896 , \24600_24902 );
and \U$15782 ( \24602_24904 , \14710_14631 , \17808_18107_nG9be7 );
and \U$15783 ( \24603_24905 , \14329_14628 , \18789_19091_nG9be4 );
or \U$15784 ( \24604_24906 , \24602_24904 , \24603_24905 );
xor \U$15785 ( \24605_24907 , \14328_14627 , \24604_24906 );
buf \U$15786 ( \24606_24908 , \24605_24907 );
buf \U$15788 ( \24607_24909 , \24606_24908 );
xor \U$15789 ( \24608_24910 , \24601_24903 , \24607_24909 );
buf \U$15790 ( \24609_24911 , \24608_24910 );
and \U$15791 ( \24610_24912 , \10996_10421 , \22330_22629_nG9bd5 );
and \U$15792 ( \24611_24913 , \10119_10418 , \23394_23696_nG9bd2 );
or \U$15793 ( \24612_24914 , \24610_24912 , \24611_24913 );
xor \U$15794 ( \24613_24915 , \10118_10417 , \24612_24914 );
buf \U$15795 ( \24614_24916 , \24613_24915 );
buf \U$15797 ( \24615_24917 , \24614_24916 );
xor \U$15798 ( \24616_24918 , \24609_24911 , \24615_24917 );
and \U$15799 ( \24617_24919 , \10411_10707 , \23927_24226_nG9bcf );
and \U$15800 ( \24618_24920 , \23557_23856 , \23863_24162 );
and \U$15801 ( \24619_24921 , \23863_24162 , \23915_24214 );
and \U$15802 ( \24620_24922 , \23557_23856 , \23915_24214 );
or \U$15803 ( \24621_24923 , \24618_24920 , \24619_24921 , \24620_24922 );
and \U$15804 ( \24622_24924 , \23890_24189 , \23894_24193 );
and \U$15805 ( \24623_24925 , \23894_24193 , \23913_24212 );
and \U$15806 ( \24624_24926 , \23890_24189 , \23913_24212 );
or \U$15807 ( \24625_24927 , \24622_24924 , \24623_24925 , \24624_24926 );
and \U$15808 ( \24626_24928 , \23561_23860 , \23847_24146 );
and \U$15809 ( \24627_24929 , \23847_24146 , \23862_24161 );
and \U$15810 ( \24628_24930 , \23561_23860 , \23862_24161 );
or \U$15811 ( \24629_24931 , \24626_24928 , \24627_24929 , \24628_24930 );
xor \U$15812 ( \24630_24932 , \24625_24927 , \24629_24931 );
and \U$15813 ( \24631_24933 , \23903_24202 , \23907_24206 );
and \U$15814 ( \24632_24934 , \23907_24206 , \23912_24211 );
and \U$15815 ( \24633_24935 , \23903_24202 , \23912_24211 );
or \U$15816 ( \24634_24936 , \24631_24933 , \24632_24934 , \24633_24935 );
and \U$15817 ( \24635_24937 , \23565_23864 , \23569_23868 );
and \U$15818 ( \24636_24938 , \23569_23868 , \23846_24145 );
and \U$15819 ( \24637_24939 , \23565_23864 , \23846_24145 );
or \U$15820 ( \24638_24940 , \24635_24937 , \24636_24938 , \24637_24939 );
xor \U$15821 ( \24639_24941 , \24634_24936 , \24638_24940 );
and \U$15822 ( \24640_24942 , \23872_24171 , \23874_24173 );
xor \U$15823 ( \24641_24943 , \24639_24941 , \24640_24942 );
xor \U$15824 ( \24642_24944 , \24630_24932 , \24641_24943 );
xor \U$15825 ( \24643_24945 , \24621_24923 , \24642_24944 );
and \U$15826 ( \24644_24946 , \23868_24167 , \23885_24184 );
and \U$15827 ( \24645_24947 , \23885_24184 , \23914_24213 );
and \U$15828 ( \24646_24948 , \23868_24167 , \23914_24213 );
or \U$15829 ( \24647_24949 , \24644_24946 , \24645_24947 , \24646_24948 );
and \U$15830 ( \24648_24950 , \23852_24151 , \23856_24155 );
and \U$15831 ( \24649_24951 , \23856_24155 , \23861_24160 );
and \U$15832 ( \24650_24952 , \23852_24151 , \23861_24160 );
or \U$15833 ( \24651_24953 , \24648_24950 , \24649_24951 , \24650_24952 );
and \U$15834 ( \24652_24954 , \17736_18035 , \15037_15336 );
and \U$15835 ( \24653_24955 , \18730_19032 , \14661_14963 );
nor \U$15836 ( \24654_24956 , \24652_24954 , \24653_24955 );
xnor \U$15837 ( \24655_24957 , \24654_24956 , \15043_15342 );
and \U$15838 ( \24656_24958 , \13725_14024 , \19235_19534 );
and \U$15839 ( \24657_24959 , \14648_14950 , \18743_19045 );
nor \U$15840 ( \24658_24960 , \24656_24958 , \24657_24959 );
xnor \U$15841 ( \24659_24961 , \24658_24960 , \19241_19540 );
xor \U$15842 ( \24660_24962 , \24655_24957 , \24659_24961 );
and \U$15843 ( \24661_24963 , \12470_12769 , \20706_21005 );
and \U$15844 ( \24662_24964 , \13377_13679 , \20255_20557 );
nor \U$15845 ( \24663_24965 , \24661_24963 , \24662_24964 );
xnor \U$15846 ( \24664_24966 , \24663_24965 , \20712_21011 );
xor \U$15847 ( \24665_24967 , \24660_24962 , \24664_24966 );
xor \U$15848 ( \24666_24968 , \24651_24953 , \24665_24967 );
and \U$15849 ( \24667_24969 , \20734_21033 , \12491_12790 );
and \U$15850 ( \24668_24970 , \21788_22090 , \12159_12461 );
nor \U$15851 ( \24669_24971 , \24667_24969 , \24668_24970 );
xnor \U$15852 ( \24670_24972 , \24669_24971 , \12481_12780 );
and \U$15853 ( \24671_24973 , \16353_16655 , \16333_16635 );
and \U$15854 ( \24672_24974 , \17325_17627 , \15999_16301 );
nor \U$15855 ( \24673_24975 , \24671_24973 , \24672_24974 );
xnor \U$15856 ( \24674_24976 , \24673_24975 , \16323_16625 );
xor \U$15857 ( \24675_24977 , \24670_24972 , \24674_24976 );
and \U$15858 ( \24676_24978 , \15022_15321 , \17791_18090 );
and \U$15859 ( \24677_24979 , \15965_16267 , \17353_17655 );
nor \U$15860 ( \24678_24980 , \24676_24978 , \24677_24979 );
xnor \U$15861 ( \24679_24981 , \24678_24980 , \17747_18046 );
xor \U$15862 ( \24680_24982 , \24675_24977 , \24679_24981 );
xor \U$15863 ( \24681_24983 , \24666_24968 , \24680_24982 );
xor \U$15864 ( \24682_24984 , \24647_24949 , \24681_24983 );
and \U$15865 ( \24683_24985 , \23875_24174 , \23879_24178 );
and \U$15866 ( \24684_24986 , \23879_24178 , \23884_24183 );
and \U$15867 ( \24685_24987 , \23875_24174 , \23884_24183 );
or \U$15868 ( \24686_24988 , \24683_24985 , \24684_24986 , \24685_24987 );
and \U$15869 ( \24687_24989 , \22257_22556 , \11275_11574 );
and \U$15870 ( \24688_24990 , \23315_23617 , \10976_11278 );
nor \U$15871 ( \24689_24991 , \24687_24989 , \24688_24990 );
xnor \U$15872 ( \24690_24992 , \24689_24991 , \11281_11580 );
and \U$15873 ( \24691_24993 , \19259_19558 , \13755_14054 );
and \U$15874 ( \24692_24994 , \20242_20544 , \13390_13692 );
nor \U$15875 ( \24693_24995 , \24691_24993 , \24692_24994 );
xnor \U$15876 ( \24694_24996 , \24693_24995 , \13736_14035 );
xor \U$15877 ( \24695_24997 , \24690_24992 , \24694_24996 );
and \U$15878 ( \24696_24998 , RIdec5540_709, \9034_9333 );
and \U$15879 ( \24697_24999 , RIdec2840_677, \9036_9335 );
and \U$15880 ( \24698_25000 , RIfcc4dc0_7262, \9038_9337 );
and \U$15881 ( \24699_25001 , RIdebfb40_645, \9040_9339 );
and \U$15882 ( \24700_25002 , RIfc9d7c0_6814, \9042_9341 );
and \U$15883 ( \24701_25003 , RIdebce40_613, \9044_9343 );
and \U$15884 ( \24702_25004 , RIdeba140_581, \9046_9345 );
and \U$15885 ( \24703_25005 , RIdeb7440_549, \9048_9347 );
and \U$15886 ( \24704_25006 , RIfc4d978_5905, \9050_9349 );
and \U$15887 ( \24705_25007 , RIdeb1a40_485, \9052_9351 );
and \U$15888 ( \24706_25008 , RIfc9dbf8_6817, \9054_9353 );
and \U$15889 ( \24707_25009 , RIdeaed40_453, \9056_9355 );
and \U$15890 ( \24708_25010 , RIfcb8610_7120, \9058_9357 );
and \U$15891 ( \24709_25011 , RIdeaa768_421, \9060_9359 );
and \U$15892 ( \24710_25012 , RIdea3e68_389, \9062_9361 );
and \U$15893 ( \24711_25013 , RIde9d568_357, \9064_9363 );
and \U$15894 ( \24712_25014 , RIfc50678_5937, \9066_9365 );
and \U$15895 ( \24713_25015 , RIfc507e0_5938, \9068_9367 );
and \U$15896 ( \24714_25016 , RIfc9dec8_6819, \9070_9369 );
and \U$15897 ( \24715_25017 , RIfc853a0_6538, \9072_9371 );
and \U$15898 ( \24716_25018 , RIde913d0_298, \9074_9373 );
and \U$15899 ( \24717_25019 , RIde8dc08_281, \9076_9375 );
and \U$15900 ( \24718_25020 , RIde89a68_261, \9078_9377 );
and \U$15901 ( \24719_25021 , RIde858c8_241, \9080_9379 );
and \U$15902 ( \24720_25022 , RIde81a70_222, \9082_9381 );
and \U$15903 ( \24721_25023 , RIfc84860_6530, \9084_9383 );
and \U$15904 ( \24722_25024 , RIfc50948_5939, \9086_9385 );
and \U$15905 ( \24723_25025 , RIfc84c98_6533, \9088_9387 );
and \U$15906 ( \24724_25026 , RIfcb7da0_7114, \9090_9389 );
and \U$15907 ( \24725_25027 , RIe16b7b0_2600, \9092_9391 );
and \U$15908 ( \24726_25028 , RIe169b90_2580, \9094_9393 );
and \U$15909 ( \24727_25029 , RIe167e08_2559, \9096_9395 );
and \U$15910 ( \24728_25030 , RIe165540_2530, \9098_9397 );
and \U$15911 ( \24729_25031 , RIe162840_2498, \9100_9399 );
and \U$15912 ( \24730_25032 , RIee37528_5088, \9102_9401 );
and \U$15913 ( \24731_25033 , RIe15fb40_2466, \9104_9403 );
and \U$15914 ( \24732_25034 , RIfcb5be0_7090, \9106_9405 );
and \U$15915 ( \24733_25035 , RIe15ce40_2434, \9108_9407 );
and \U$15916 ( \24734_25036 , RIe157440_2370, \9110_9409 );
and \U$15917 ( \24735_25037 , RIe154740_2338, \9112_9411 );
and \U$15918 ( \24736_25038 , RIfcd35c8_7427, \9114_9413 );
and \U$15919 ( \24737_25039 , RIe151a40_2306, \9116_9415 );
and \U$15920 ( \24738_25040 , RIfc53a80_5974, \9118_9417 );
and \U$15921 ( \24739_25041 , RIe14ed40_2274, \9120_9419 );
and \U$15922 ( \24740_25042 , RIfcc6170_7276, \9122_9421 );
and \U$15923 ( \24741_25043 , RIe14c040_2242, \9124_9423 );
and \U$15924 ( \24742_25044 , RIe149340_2210, \9126_9425 );
and \U$15925 ( \24743_25045 , RIe146640_2178, \9128_9427 );
and \U$15926 ( \24744_25046 , RIfc7f130_6468, \9130_9429 );
and \U$15927 ( \24745_25047 , RIee33310_5041, \9132_9431 );
and \U$15928 ( \24746_25048 , RIfcb4f38_7081, \9134_9433 );
and \U$15929 ( \24747_25049 , RIfc47f78_5841, \9136_9435 );
and \U$15930 ( \24748_25050 , RIe140f10_2116, \9138_9437 );
and \U$15931 ( \24749_25051 , RIdf3ee18_2092, \9140_9439 );
and \U$15932 ( \24750_25052 , RIdf3cc58_2068, \9142_9441 );
and \U$15933 ( \24751_25053 , RIdf3a7c8_2042, \9144_9443 );
and \U$15934 ( \24752_25054 , RIfc7fc70_6476, \9146_9445 );
and \U$15935 ( \24753_25055 , RIfcd27b8_7417, \9148_9447 );
and \U$15936 ( \24754_25056 , RIfca1000_6854, \9150_9449 );
and \U$15937 ( \24755_25057 , RIfcc6b48_7283, \9152_9451 );
and \U$15938 ( \24756_25058 , RIdf35908_1986, \9154_9453 );
and \U$15939 ( \24757_25059 , RIdf33478_1960, \9156_9455 );
and \U$15940 ( \24758_25060 , RIfebe9f8_8289, \9158_9457 );
and \U$15941 ( \24759_25061 , RIdf2f260_1913, \9160_9459 );
or \U$15942 ( \24760_25062 , \24696_24998 , \24697_24999 , \24698_25000 , \24699_25001 , \24700_25002 , \24701_25003 , \24702_25004 , \24703_25005 , \24704_25006 , \24705_25007 , \24706_25008 , \24707_25009 , \24708_25010 , \24709_25011 , \24710_25012 , \24711_25013 , \24712_25014 , \24713_25015 , \24714_25016 , \24715_25017 , \24716_25018 , \24717_25019 , \24718_25020 , \24719_25021 , \24720_25022 , \24721_25023 , \24722_25024 , \24723_25025 , \24724_25026 , \24725_25027 , \24726_25028 , \24727_25029 , \24728_25030 , \24729_25031 , \24730_25032 , \24731_25033 , \24732_25034 , \24733_25035 , \24734_25036 , \24735_25037 , \24736_25038 , \24737_25039 , \24738_25040 , \24739_25041 , \24740_25042 , \24741_25043 , \24742_25044 , \24743_25045 , \24744_25046 , \24745_25047 , \24746_25048 , \24747_25049 , \24748_25050 , \24749_25051 , \24750_25052 , \24751_25053 , \24752_25054 , \24753_25055 , \24754_25056 , \24755_25057 , \24756_25058 , \24757_25059 , \24758_25060 , \24759_25061 );
and \U$15943 ( \24761_25063 , RIfcb7968_7111, \9163_9462 );
and \U$15944 ( \24762_25064 , RIee2a3a0_4939, \9165_9464 );
and \U$15945 ( \24763_25065 , RIfc51050_5944, \9167_9466 );
and \U$15946 ( \24764_25066 , RIfcd3fa0_7434, \9169_9468 );
and \U$15947 ( \24765_25067 , RIdf2a3a0_1857, \9171_9470 );
and \U$15948 ( \24766_25068 , RIdf28078_1832, \9173_9472 );
and \U$15949 ( \24767_25069 , RIfe81198_7813, \9175_9474 );
and \U$15950 ( \24768_25070 , RIdf24838_1792, \9177_9476 );
and \U$15951 ( \24769_25071 , RIfc84428_6527, \9179_9478 );
and \U$15952 ( \24770_25072 , RIfce7ed8_7661, \9181_9480 );
and \U$15953 ( \24771_25073 , RIdf22d80_1773, \9183_9482 );
and \U$15954 ( \24772_25074 , RIfc515f0_5948, \9185_9484 );
and \U$15955 ( \24773_25075 , RIdf21868_1758, \9187_9486 );
and \U$15956 ( \24774_25076 , RIdf1f978_1736, \9189_9488 );
and \U$15957 ( \24775_25077 , RIdf1b058_1684, \9191_9490 );
and \U$15958 ( \24776_25078 , RIdf192d0_1663, \9193_9492 );
and \U$15959 ( \24777_25079 , RIdf17110_1639, \9195_9494 );
and \U$15960 ( \24778_25080 , RIdf14410_1607, \9197_9496 );
and \U$15961 ( \24779_25081 , RIdf11710_1575, \9199_9498 );
and \U$15962 ( \24780_25082 , RIdf0ea10_1543, \9201_9500 );
and \U$15963 ( \24781_25083 , RIdf0bd10_1511, \9203_9502 );
and \U$15964 ( \24782_25084 , RIdf09010_1479, \9205_9504 );
and \U$15965 ( \24783_25085 , RIdf06310_1447, \9207_9506 );
and \U$15966 ( \24784_25086 , RIdf03610_1415, \9209_9508 );
and \U$15967 ( \24785_25087 , RIdefdc10_1351, \9211_9510 );
and \U$15968 ( \24786_25088 , RIdefaf10_1319, \9213_9512 );
and \U$15969 ( \24787_25089 , RIdef8210_1287, \9215_9514 );
and \U$15970 ( \24788_25090 , RIdef5510_1255, \9217_9516 );
and \U$15971 ( \24789_25091 , RIdef2810_1223, \9219_9518 );
and \U$15972 ( \24790_25092 , RIdeefb10_1191, \9221_9520 );
and \U$15973 ( \24791_25093 , RIdeece10_1159, \9223_9522 );
and \U$15974 ( \24792_25094 , RIdeea110_1127, \9225_9524 );
and \U$15975 ( \24793_25095 , RIfc7e1b8_6457, \9227_9526 );
and \U$15976 ( \24794_25096 , RIfca19d8_6861, \9229_9528 );
and \U$15977 ( \24795_25097 , RIfc7dab0_6452, \9231_9530 );
and \U$15978 ( \24796_25098 , RIfc7e488_6459, \9233_9532 );
and \U$15979 ( \24797_25099 , RIdee49e0_1065, \9235_9534 );
and \U$15980 ( \24798_25100 , RIfe80d60_7810, \9237_9536 );
and \U$15981 ( \24799_25101 , RIfeabba0_8270, \9239_9538 );
and \U$15982 ( \24800_25102 , RIfe80bf8_7809, \9241_9540 );
and \U$15983 ( \24801_25103 , RIfcb3750_7064, \9243_9542 );
and \U$15984 ( \24802_25104 , RIfce9f30_7684, \9245_9544 );
and \U$15985 ( \24803_25105 , RIfc7e5f0_6460, \9247_9546 );
and \U$15986 ( \24804_25106 , RIfc56a50_6008, \9249_9548 );
and \U$15987 ( \24805_25107 , RIfe81030_7812, \9251_9550 );
and \U$15988 ( \24806_25108 , RIded7420_913, \9253_9552 );
and \U$15989 ( \24807_25109 , RIfe80ec8_7811, \9255_9554 );
and \U$15990 ( \24808_25110 , RIded2f38_864, \9257_9556 );
and \U$15991 ( \24809_25111 , RIded0940_837, \9259_9558 );
and \U$15992 ( \24810_25112 , RIdecdc40_805, \9261_9560 );
and \U$15993 ( \24811_25113 , RIdecaf40_773, \9263_9562 );
and \U$15994 ( \24812_25114 , RIdec8240_741, \9265_9564 );
and \U$15995 ( \24813_25115 , RIdeb4740_517, \9267_9566 );
and \U$15996 ( \24814_25116 , RIde96c68_325, \9269_9568 );
and \U$15997 ( \24815_25117 , RIe16e348_2631, \9271_9570 );
and \U$15998 ( \24816_25118 , RIe15a140_2402, \9273_9572 );
and \U$15999 ( \24817_25119 , RIe143940_2146, \9275_9574 );
and \U$16000 ( \24818_25120 , RIdf38338_2016, \9277_9576 );
and \U$16001 ( \24819_25121 , RIdf2c998_1884, \9279_9578 );
and \U$16002 ( \24820_25122 , RIdf1d218_1708, \9281_9580 );
and \U$16003 ( \24821_25123 , RIdf00910_1383, \9283_9582 );
and \U$16004 ( \24822_25124 , RIdee7410_1095, \9285_9584 );
and \U$16005 ( \24823_25125 , RIdedc178_968, \9287_9586 );
and \U$16006 ( \24824_25126 , RIde7cbb0_198, \9289_9588 );
or \U$16007 ( \24825_25127 , \24761_25063 , \24762_25064 , \24763_25065 , \24764_25066 , \24765_25067 , \24766_25068 , \24767_25069 , \24768_25070 , \24769_25071 , \24770_25072 , \24771_25073 , \24772_25074 , \24773_25075 , \24774_25076 , \24775_25077 , \24776_25078 , \24777_25079 , \24778_25080 , \24779_25081 , \24780_25082 , \24781_25083 , \24782_25084 , \24783_25085 , \24784_25086 , \24785_25087 , \24786_25088 , \24787_25089 , \24788_25090 , \24789_25091 , \24790_25092 , \24791_25093 , \24792_25094 , \24793_25095 , \24794_25096 , \24795_25097 , \24796_25098 , \24797_25099 , \24798_25100 , \24799_25101 , \24800_25102 , \24801_25103 , \24802_25104 , \24803_25105 , \24804_25106 , \24805_25107 , \24806_25108 , \24807_25109 , \24808_25110 , \24809_25111 , \24810_25112 , \24811_25113 , \24812_25114 , \24813_25115 , \24814_25116 , \24815_25117 , \24816_25118 , \24817_25119 , \24818_25120 , \24819_25121 , \24820_25122 , \24821_25123 , \24822_25124 , \24823_25125 , \24824_25126 );
or \U$16008 ( \24826_25128 , \24760_25062 , \24825_25127 );
_DC \g5ba0/U$1 ( \24827 , \24826_25128 , \9298_9597 );
and \U$16009 ( \24828_25130 , RIe19d7d8_3169, \8760_9059 );
and \U$16010 ( \24829_25131 , RIe19aad8_3137, \8762_9061 );
and \U$16011 ( \24830_25132 , RIfcc2d68_7239, \8764_9063 );
and \U$16012 ( \24831_25133 , RIe197dd8_3105, \8766_9065 );
and \U$16013 ( \24832_25134 , RIfc5c5b8_6073, \8768_9067 );
and \U$16014 ( \24833_25135 , RIe1950d8_3073, \8770_9069 );
and \U$16015 ( \24834_25136 , RIe1923d8_3041, \8772_9071 );
and \U$16016 ( \24835_25137 , RIe18f6d8_3009, \8774_9073 );
and \U$16017 ( \24836_25138 , RIe189cd8_2945, \8776_9075 );
and \U$16018 ( \24837_25139 , RIe186fd8_2913, \8778_9077 );
and \U$16019 ( \24838_25140 , RIf1438d0_5228, \8780_9079 );
and \U$16020 ( \24839_25141 , RIe1842d8_2881, \8782_9081 );
and \U$16021 ( \24840_25142 , RIfc5b370_6060, \8784_9083 );
and \U$16022 ( \24841_25143 , RIe1815d8_2849, \8786_9085 );
and \U$16023 ( \24842_25144 , RIe17e8d8_2817, \8788_9087 );
and \U$16024 ( \24843_25145 , RIe17bbd8_2785, \8790_9089 );
and \U$16025 ( \24844_25146 , RIfcbb748_7155, \8792_9091 );
and \U$16026 ( \24845_25147 , RIfc59480_6038, \8794_9093 );
and \U$16027 ( \24846_25148 , RIfcbbce8_7159, \8796_9095 );
and \U$16028 ( \24847_25149 , RIe175c38_2717, \8798_9097 );
and \U$16029 ( \24848_25150 , RIfcdb890_7520, \8800_9099 );
and \U$16030 ( \24849_25151 , RIfc59b88_6043, \8802_9101 );
and \U$16031 ( \24850_25152 , RIfc8ada0_6602, \8804_9103 );
and \U$16032 ( \24851_25153 , RIfcb5eb0_7092, \8806_9105 );
and \U$16033 ( \24852_25154 , RIfc57c98_6021, \8808_9107 );
and \U$16034 ( \24853_25155 , RIfc57158_6013, \8810_9109 );
and \U$16035 ( \24854_25156 , RIfc58aa8_6031, \8812_9111 );
and \U$16036 ( \24855_25157 , RIe173910_2692, \8814_9113 );
and \U$16037 ( \24856_25158 , RIfcc62d8_7277, \8816_9115 );
and \U$16038 ( \24857_25159 , RIfc8a968_6599, \8818_9117 );
and \U$16039 ( \24858_25160 , RIfc57428_6015, \8820_9119 );
and \U$16040 ( \24859_25161 , RIfc56d20_6010, \8822_9121 );
and \U$16041 ( \24860_25162 , RIfc408e0_5760, \8824_9123 );
and \U$16042 ( \24861_25163 , RIe223b30_4696, \8826_9125 );
and \U$16043 ( \24862_25164 , RIfc82970_6508, \8828_9127 );
and \U$16044 ( \24863_25165 , RIe220e30_4664, \8830_9129 );
and \U$16045 ( \24864_25166 , RIfcecc30_7716, \8832_9131 );
and \U$16046 ( \24865_25167 , RIe21e130_4632, \8834_9133 );
and \U$16047 ( \24866_25168 , RIe218730_4568, \8836_9135 );
and \U$16048 ( \24867_25169 , RIe215a30_4536, \8838_9137 );
and \U$16049 ( \24868_25170 , RIfc3fad0_5750, \8840_9139 );
and \U$16050 ( \24869_25171 , RIe212d30_4504, \8842_9141 );
and \U$16051 ( \24870_25172 , RIf169148_5655, \8844_9143 );
and \U$16052 ( \24871_25173 , RIe210030_4472, \8846_9145 );
and \U$16053 ( \24872_25174 , RIfc545c0_5982, \8848_9147 );
and \U$16054 ( \24873_25175 , RIe20d330_4440, \8850_9149 );
and \U$16055 ( \24874_25176 , RIe20a630_4408, \8852_9151 );
and \U$16056 ( \24875_25177 , RIe207930_4376, \8854_9153 );
and \U$16057 ( \24876_25178 , RIfc88d48_6579, \8856_9155 );
and \U$16058 ( \24877_25179 , RIfc4bec0_5886, \8858_9157 );
and \U$16059 ( \24878_25180 , RIe202638_4317, \8860_9159 );
and \U$16060 ( \24879_25181 , RIe200b80_4298, \8862_9161 );
and \U$16061 ( \24880_25182 , RIfc88910_6576, \8864_9163 );
and \U$16062 ( \24881_25183 , RIfc4c190_5888, \8866_9165 );
and \U$16063 ( \24882_25184 , RIfc4c2f8_5889, \8868_9167 );
and \U$16064 ( \24883_25185 , RIfcba398_7141, \8870_9169 );
and \U$16065 ( \24884_25186 , RIfcd4270_7436, \8872_9171 );
and \U$16066 ( \24885_25187 , RIfcba0c8_7139, \8874_9173 );
and \U$16067 ( \24886_25188 , RIe1fcda0_4254, \8876_9175 );
and \U$16068 ( \24887_25189 , RIe1fbb58_4241, \8878_9177 );
and \U$16069 ( \24888_25190 , RIfc53d50_5976, \8880_9179 );
and \U$16070 ( \24889_25191 , RIfc9b768_6791, \8882_9181 );
and \U$16071 ( \24890_25192 , RIfc537b0_5972, \8884_9183 );
and \U$16072 ( \24891_25193 , RIfc4c5c8_5891, \8886_9185 );
or \U$16073 ( \24892_25194 , \24828_25130 , \24829_25131 , \24830_25132 , \24831_25133 , \24832_25134 , \24833_25135 , \24834_25136 , \24835_25137 , \24836_25138 , \24837_25139 , \24838_25140 , \24839_25141 , \24840_25142 , \24841_25143 , \24842_25144 , \24843_25145 , \24844_25146 , \24845_25147 , \24846_25148 , \24847_25149 , \24848_25150 , \24849_25151 , \24850_25152 , \24851_25153 , \24852_25154 , \24853_25155 , \24854_25156 , \24855_25157 , \24856_25158 , \24857_25159 , \24858_25160 , \24859_25161 , \24860_25162 , \24861_25163 , \24862_25164 , \24863_25165 , \24864_25166 , \24865_25167 , \24866_25168 , \24867_25169 , \24868_25170 , \24869_25171 , \24870_25172 , \24871_25173 , \24872_25174 , \24873_25175 , \24874_25176 , \24875_25177 , \24876_25178 , \24877_25179 , \24878_25180 , \24879_25181 , \24880_25182 , \24881_25183 , \24882_25184 , \24883_25185 , \24884_25186 , \24885_25187 , \24886_25188 , \24887_25189 , \24888_25190 , \24889_25191 , \24890_25192 , \24891_25193 );
and \U$16074 ( \24893_25195 , RIfc9e468_6823, \8889_9188 );
and \U$16075 ( \24894_25196 , RIf157da8_5459, \8891_9190 );
and \U$16076 ( \24895_25197 , RIfcb9f60_7138, \8893_9192 );
and \U$16077 ( \24896_25198 , RIe1fa208_4223, \8895_9194 );
and \U$16078 ( \24897_25199 , RIfc849c8_6531, \8897_9196 );
and \U$16079 ( \24898_25200 , RIfc529a0_5962, \8899_9198 );
and \U$16080 ( \24899_25201 , RIfc9f6b0_6836, \8901_9200 );
and \U$16081 ( \24900_25202 , RIe1f5618_4169, \8903_9202 );
and \U$16082 ( \24901_25203 , RIf153320_5406, \8905_9204 );
and \U$16083 ( \24902_25204 , RIfcc4988_7259, \8907_9206 );
and \U$16084 ( \24903_25205 , RIf150d28_5379, \8909_9208 );
and \U$16085 ( \24904_25206 , RIfebe458_8285, \8911_9210 );
and \U$16086 ( \24905_25207 , RIfc87f38_6569, \8913_9212 );
and \U$16087 ( \24906_25208 , RIfcb7f08_7115, \8915_9214 );
and \U$16088 ( \24907_25209 , RIf14e190_5348, \8917_9216 );
and \U$16089 ( \24908_25210 , RIfe80658_7805, \8919_9218 );
and \U$16090 ( \24909_25211 , RIe1eb898_4057, \8921_9220 );
and \U$16091 ( \24910_25212 , RIe1e8b98_4025, \8923_9222 );
and \U$16092 ( \24911_25213 , RIe1e5e98_3993, \8925_9224 );
and \U$16093 ( \24912_25214 , RIe1e3198_3961, \8927_9226 );
and \U$16094 ( \24913_25215 , RIe1e0498_3929, \8929_9228 );
and \U$16095 ( \24914_25216 , RIe1dd798_3897, \8931_9230 );
and \U$16096 ( \24915_25217 , RIe1daa98_3865, \8933_9232 );
and \U$16097 ( \24916_25218 , RIe1d7d98_3833, \8935_9234 );
and \U$16098 ( \24917_25219 , RIe1d2398_3769, \8937_9236 );
and \U$16099 ( \24918_25220 , RIe1cf698_3737, \8939_9238 );
and \U$16100 ( \24919_25221 , RIe1cc998_3705, \8941_9240 );
and \U$16101 ( \24920_25222 , RIe1c9c98_3673, \8943_9242 );
and \U$16102 ( \24921_25223 , RIe1c6f98_3641, \8945_9244 );
and \U$16103 ( \24922_25224 , RIe1c4298_3609, \8947_9246 );
and \U$16104 ( \24923_25225 , RIe1c1598_3577, \8949_9248 );
and \U$16105 ( \24924_25226 , RIe1be898_3545, \8951_9250 );
and \U$16106 ( \24925_25227 , RIf14cc78_5333, \8953_9252 );
and \U$16107 ( \24926_25228 , RIf14ba30_5320, \8955_9254 );
and \U$16108 ( \24927_25229 , RIe1b92d0_3484, \8957_9256 );
and \U$16109 ( \24928_25230 , RIe1b7278_3461, \8959_9258 );
and \U$16110 ( \24929_25231 , RIf14a7e8_5307, \8961_9260 );
and \U$16111 ( \24930_25232 , RIf149ca8_5299, \8963_9262 );
and \U$16112 ( \24931_25233 , RIfebe5c0_8286, \8965_9264 );
and \U$16113 ( \24932_25234 , RIfe807c0_7806, \8967_9266 );
and \U$16114 ( \24933_25235 , RIfc50510_5936, \8969_9268 );
and \U$16115 ( \24934_25236 , RIfce4f08_7627, \8971_9270 );
and \U$16116 ( \24935_25237 , RIfe80a90_7808, \8973_9272 );
and \U$16117 ( \24936_25238 , RIfebe890_8288, \8975_9274 );
and \U$16118 ( \24937_25239 , RIfc9cde8_6807, \8977_9276 );
and \U$16119 ( \24938_25240 , RIfc87560_6562, \8979_9278 );
and \U$16120 ( \24939_25241 , RIfe80928_7807, \8981_9280 );
and \U$16121 ( \24940_25242 , RIfebe728_8287, \8983_9282 );
and \U$16122 ( \24941_25243 , RIe1a8bd8_3297, \8985_9284 );
and \U$16123 ( \24942_25244 , RIe1a5ed8_3265, \8987_9286 );
and \U$16124 ( \24943_25245 , RIe1a31d8_3233, \8989_9288 );
and \U$16125 ( \24944_25246 , RIe1a04d8_3201, \8991_9290 );
and \U$16126 ( \24945_25247 , RIe18c9d8_2977, \8993_9292 );
and \U$16127 ( \24946_25248 , RIe178ed8_2753, \8995_9294 );
and \U$16128 ( \24947_25249 , RIe226830_4728, \8997_9296 );
and \U$16129 ( \24948_25250 , RIe21b430_4600, \8999_9298 );
and \U$16130 ( \24949_25251 , RIe204c30_4344, \9001_9300 );
and \U$16131 ( \24950_25252 , RIe1fec90_4276, \9003_9302 );
and \U$16132 ( \24951_25253 , RIe1f8048_4199, \9005_9304 );
and \U$16133 ( \24952_25254 , RIe1f0b90_4116, \9007_9306 );
and \U$16134 ( \24953_25255 , RIe1d5098_3801, \9009_9308 );
and \U$16135 ( \24954_25256 , RIe1bbb98_3513, \9011_9310 );
and \U$16136 ( \24955_25257 , RIe1aea10_3364, \9013_9312 );
and \U$16137 ( \24956_25258 , RIe171048_2663, \9015_9314 );
or \U$16138 ( \24957_25259 , \24893_25195 , \24894_25196 , \24895_25197 , \24896_25198 , \24897_25199 , \24898_25200 , \24899_25201 , \24900_25202 , \24901_25203 , \24902_25204 , \24903_25205 , \24904_25206 , \24905_25207 , \24906_25208 , \24907_25209 , \24908_25210 , \24909_25211 , \24910_25212 , \24911_25213 , \24912_25214 , \24913_25215 , \24914_25216 , \24915_25217 , \24916_25218 , \24917_25219 , \24918_25220 , \24919_25221 , \24920_25222 , \24921_25223 , \24922_25224 , \24923_25225 , \24924_25226 , \24925_25227 , \24926_25228 , \24927_25229 , \24928_25230 , \24929_25231 , \24930_25232 , \24931_25233 , \24932_25234 , \24933_25235 , \24934_25236 , \24935_25237 , \24936_25238 , \24937_25239 , \24938_25240 , \24939_25241 , \24940_25242 , \24941_25243 , \24942_25244 , \24943_25245 , \24944_25246 , \24945_25247 , \24946_25248 , \24947_25249 , \24948_25250 , \24949_25251 , \24950_25252 , \24951_25253 , \24952_25254 , \24953_25255 , \24954_25256 , \24955_25257 , \24956_25258 );
or \U$16139 ( \24958_25260 , \24892_25194 , \24957_25259 );
_DC \g5c24/U$1 ( \24959 , \24958_25260 , \9024_9323 );
xor g5c25_GF_PartitionCandidate( \24960_25262_nG5c25 , \24827 , \24959 );
buf \U$16140 ( \24961_25263 , \24960_25262_nG5c25 );
xor \U$16141 ( \24962_25264 , \24961_25263 , \23836_24135 );
and \U$16142 ( \24963_25265 , \10385_10687 , \24962_25264 );
xor \U$16143 ( \24964_25266 , \24695_24997 , \24963_25265 );
xor \U$16144 ( \24965_25267 , \24686_24988 , \24964_25266 );
and \U$16145 ( \24966_25268 , \23900_24199 , \10681_10983 );
_DC \g65b9/U$1 ( \24967 , \24826_25128 , \9298_9597 );
_DC \g65ba/U$1 ( \24968 , \24958_25260 , \9024_9323 );
and g65bb_GF_PartitionCandidate( \24969_25271_nG65bb , \24967 , \24968 );
buf \U$16146 ( \24970_25272 , \24969_25271_nG65bb );
and \U$16147 ( \24971_25273 , \24970_25272 , \10389_10691 );
nor \U$16148 ( \24972_25274 , \24966_25268 , \24971_25273 );
xnor \U$16149 ( \24973_25275 , \24972_25274 , \10678_10980 );
and \U$16150 ( \24974_25276 , \11287_11586 , \22243_22542 );
and \U$16151 ( \24975_25277 , \12146_12448 , \21801_22103 );
nor \U$16152 ( \24976_25278 , \24974_25276 , \24975_25277 );
xnor \U$16153 ( \24977_25279 , \24976_25278 , \22249_22548 );
xor \U$16154 ( \24978_25280 , \24973_25275 , \24977_25279 );
and \U$16155 ( \24979_25281 , \10686_10988 , \23839_24138 );
and \U$16156 ( \24980_25282 , \10968_11270 , \23328_23630 );
nor \U$16157 ( \24981_25283 , \24979_25281 , \24980_25282 );
xnor \U$16158 ( \24982_25284 , \24981_25283 , \23845_24144 );
xor \U$16159 ( \24983_25285 , \24978_25280 , \24982_25284 );
xor \U$16160 ( \24984_25286 , \24965_25267 , \24983_25285 );
xor \U$16161 ( \24985_25287 , \24682_24984 , \24984_25286 );
xor \U$16162 ( \24986_25288 , \24643_24945 , \24985_25287 );
and \U$16163 ( \24987_25289 , \23548_23847 , \23552_23851 );
and \U$16164 ( \24988_25290 , \23552_23851 , \23916_24215 );
and \U$16165 ( \24989_25291 , \23548_23847 , \23916_24215 );
or \U$16166 ( \24990_25292 , \24987_25289 , \24988_25290 , \24989_25291 );
xor \U$16167 ( \24991_25293 , \24986_25288 , \24990_25292 );
and \U$16168 ( \24992_25294 , \23917_24216 , \23921_24220 );
and \U$16169 ( \24993_25295 , \23922_24221 , \23925_24224 );
or \U$16170 ( \24994_25296 , \24992_25294 , \24993_25295 );
xor \U$16171 ( \24995_25297 , \24991_25293 , \24994_25296 );
buf g9bcc_GF_PartitionCandidate( \24996_25298_nG9bcc , \24995_25297 );
and \U$16172 ( \24997_25299 , \10402_10704 , \24996_25298_nG9bcc );
or \U$16173 ( \24998_25300 , \24617_24919 , \24997_25299 );
xor \U$16174 ( \24999_25301 , \10399_10703 , \24998_25300 );
buf \U$16175 ( \25000_25302 , \24999_25301 );
buf \U$16177 ( \25001_25303 , \25000_25302 );
xor \U$16178 ( \25002_25304 , \24616_24918 , \25001_25303 );
buf \U$16179 ( \25003_25305 , \25002_25304 );
xor \U$16180 ( \25004_25306 , \24577_24879 , \25003_25305 );
and \U$16181 ( \25005_25307 , \23484_23786 , \23542_23841 );
and \U$16182 ( \25006_25308 , \23484_23786 , \23932_24231 );
and \U$16183 ( \25007_25309 , \23542_23841 , \23932_24231 );
or \U$16184 ( \25008_25310 , \25005_25307 , \25006_25308 , \25007_25309 );
buf \U$16185 ( \25009_25311 , \25008_25310 );
xor \U$16186 ( \25010_25312 , \25004_25306 , \25009_25311 );
buf \U$16187 ( \25011_25313 , \25010_25312 );
xor \U$16188 ( \25012_25314 , \24572_24874 , \25011_25313 );
and \U$16189 ( \25013_25315 , \24497_24799 , \25012_25314 );
and \U$16190 ( \25014_25316 , \23447_23749 , \23452_23754 );
and \U$16191 ( \25015_25317 , \23447_23749 , \23934_24233 );
and \U$16192 ( \25016_25318 , \23452_23754 , \23934_24233 );
or \U$16193 ( \25017_25319 , \25014_25316 , \25015_25317 , \25016_25318 );
and \U$16194 ( \25018_25320 , \24497_24799 , \25017_25319 );
and \U$16195 ( \25019_25321 , \25012_25314 , \25017_25319 );
or \U$16196 ( \25020_25322 , \25013_25315 , \25018_25320 , \25019_25321 );
and \U$16197 ( \25021_25323 , \23936_24235 , \23940_24239 );
and \U$16198 ( \25022_25324 , \23936_24235 , \24496_24798 );
and \U$16199 ( \25023_25325 , \23940_24239 , \24496_24798 );
or \U$16200 ( \25024_25326 , \25021_25323 , \25022_25324 , \25023_25325 );
xor \U$16201 ( \25025_25327 , \25020_25322 , \25024_25326 );
and \U$16202 ( \25026_25328 , \24579_24881 , \24585_24887 );
and \U$16203 ( \25027_25329 , \24579_24881 , \24592_24894 );
and \U$16204 ( \25028_25330 , \24585_24887 , \24592_24894 );
or \U$16205 ( \25029_25331 , \25026_25328 , \25027_25329 , \25028_25330 );
buf \U$16206 ( \25030_25332 , \25029_25331 );
and \U$16207 ( \25031_25333 , \24489_24788 , \24493_24795 );
buf \U$16208 ( \25032_25334 , \25031_25333 );
buf \U$16210 ( \25033_25335 , \25032_25334 );
and \U$16211 ( \25034_25336 , \23495_23201 , \10981_11283_nG9c08 );
and \U$16212 ( \25035_25337 , \22899_23198 , \11299_11598_nG9c05 );
or \U$16213 ( \25036_25338 , \25034_25336 , \25035_25337 );
xor \U$16214 ( \25037_25339 , \22898_23197 , \25036_25338 );
buf \U$16215 ( \25038_25340 , \25037_25339 );
buf \U$16217 ( \25039_25341 , \25038_25340 );
xor \U$16218 ( \25040_25342 , \25033_25335 , \25039_25341 );
buf \U$16219 ( \25041_25343 , \25040_25342 );
not \U$15659 ( \25042_24790 , \24490_24789 );
xor \U$15660 ( \25043_24791 , \24484_24783_nG4412 , \24487_24786_nG4415 );
and \U$15661 ( \25044_24792 , \25042_24790 , \25043_24791 );
and \U$16220 ( \25045_25344 , \25044_24792 , \10392_10694_nG9c0e );
and \U$16221 ( \25046_25345 , \24490_24789 , \10693_10995_nG9c0b );
or \U$16222 ( \25047_25346 , \25045_25344 , \25046_25345 );
xor \U$16223 ( \25048_25347 , \24489_24788 , \25047_25346 );
buf \U$16224 ( \25049_25348 , \25048_25347 );
buf \U$16226 ( \25050_25349 , \25049_25348 );
xor \U$16227 ( \25051_25350 , \25041_25343 , \25050_25349 );
and \U$16228 ( \25052_25351 , \21908_21658 , \12168_12470_nG9c02 );
and \U$16229 ( \25053_25352 , \21356_21655 , \12502_12801_nG9bff );
or \U$16230 ( \25054_25353 , \25052_25351 , \25053_25352 );
xor \U$16231 ( \25055_25354 , \21355_21654 , \25054_25353 );
buf \U$16232 ( \25056_25355 , \25055_25354 );
buf \U$16234 ( \25057_25356 , \25056_25355 );
xor \U$16235 ( \25058_25357 , \25051_25350 , \25057_25356 );
buf \U$16236 ( \25059_25358 , \25058_25357 );
xor \U$16237 ( \25060_25359 , \25030_25332 , \25059_25358 );
and \U$16238 ( \25061_25360 , \17437_17297 , \16013_16315_nG9bf0 );
and \U$16239 ( \25062_25361 , \16995_17294 , \16378_16680_nG9bed );
or \U$16240 ( \25063_25362 , \25061_25360 , \25062_25361 );
xor \U$16241 ( \25064_25363 , \16994_17293 , \25063_25362 );
buf \U$16242 ( \25065_25364 , \25064_25363 );
buf \U$16244 ( \25066_25365 , \25065_25364 );
xor \U$16245 ( \25067_25366 , \25060_25359 , \25066_25365 );
buf \U$16246 ( \25068_25367 , \25067_25366 );
and \U$16247 ( \25069_25368 , \14710_14631 , \18789_19091_nG9be4 );
and \U$16248 ( \25070_25369 , \14329_14628 , \19287_19586_nG9be1 );
or \U$16249 ( \25071_25370 , \25069_25368 , \25070_25369 );
xor \U$16250 ( \25072_25371 , \14328_14627 , \25071_25370 );
buf \U$16251 ( \25073_25372 , \25072_25371 );
buf \U$16253 ( \25074_25373 , \25073_25372 );
xor \U$16254 ( \25075_25374 , \25068_25367 , \25074_25373 );
and \U$16255 ( \25076_25375 , \13431_13370 , \20306_20608_nG9bde );
and \U$16256 ( \25077_25376 , \13068_13367 , \20787_21086_nG9bdb );
or \U$16257 ( \25078_25377 , \25076_25375 , \25077_25376 );
xor \U$16258 ( \25079_25378 , \13067_13366 , \25078_25377 );
buf \U$16259 ( \25080_25379 , \25079_25378 );
buf \U$16261 ( \25081_25380 , \25080_25379 );
xor \U$16262 ( \25082_25381 , \25075_25374 , \25081_25380 );
buf \U$16263 ( \25083_25382 , \25082_25381 );
and \U$16264 ( \25084_25383 , \24512_24814 , \24526_24828 );
and \U$16265 ( \25085_25384 , \24512_24814 , \24533_24835 );
and \U$16266 ( \25086_25385 , \24526_24828 , \24533_24835 );
or \U$16267 ( \25087_25386 , \25084_25383 , \25085_25384 , \25086_25385 );
buf \U$16268 ( \25088_25387 , \25087_25386 );
and \U$16269 ( \25089_25388 , \24518_24820 , \24524_24826 );
buf \U$16270 ( \25090_25389 , \25089_25388 );
and \U$16271 ( \25091_25390 , \20353_20155 , \13403_13705_nG9bfc );
and \U$16272 ( \25092_25391 , \19853_20152 , \13771_14070_nG9bf9 );
or \U$16273 ( \25093_25392 , \25091_25390 , \25092_25391 );
xor \U$16274 ( \25094_25393 , \19852_20151 , \25093_25392 );
buf \U$16275 ( \25095_25394 , \25094_25393 );
buf \U$16277 ( \25096_25395 , \25095_25394 );
xor \U$16278 ( \25097_25396 , \25090_25389 , \25096_25395 );
and \U$16279 ( \25098_25397 , \18908_18702 , \14682_14984_nG9bf6 );
and \U$16280 ( \25099_25398 , \18400_18699 , \15074_15373_nG9bf3 );
or \U$16281 ( \25100_25399 , \25098_25397 , \25099_25398 );
xor \U$16282 ( \25101_25400 , \18399_18698 , \25100_25399 );
buf \U$16283 ( \25102_25401 , \25101_25400 );
buf \U$16285 ( \25103_25402 , \25102_25401 );
xor \U$16286 ( \25104_25403 , \25097_25396 , \25103_25402 );
buf \U$16287 ( \25105_25404 , \25104_25403 );
xor \U$16288 ( \25106_25405 , \25088_25387 , \25105_25404 );
and \U$16289 ( \25107_25406 , \16405_15940 , \17363_17665_nG9bea );
and \U$16290 ( \25108_25407 , \15638_15937 , \17808_18107_nG9be7 );
or \U$16291 ( \25109_25408 , \25107_25406 , \25108_25407 );
xor \U$16292 ( \25110_25409 , \15637_15936 , \25109_25408 );
buf \U$16293 ( \25111_25410 , \25110_25409 );
buf \U$16295 ( \25112_25411 , \25111_25410 );
xor \U$16296 ( \25113_25412 , \25106_25405 , \25112_25411 );
buf \U$16297 ( \25114_25413 , \25113_25412 );
xor \U$16298 ( \25115_25414 , \25083_25382 , \25114_25413 );
and \U$16299 ( \25116_25415 , \10996_10421 , \23394_23696_nG9bd2 );
and \U$16300 ( \25117_25416 , \10119_10418 , \23927_24226_nG9bcf );
or \U$16301 ( \25118_25417 , \25116_25415 , \25117_25416 );
xor \U$16302 ( \25119_25418 , \10118_10417 , \25118_25417 );
buf \U$16303 ( \25120_25419 , \25119_25418 );
buf \U$16305 ( \25121_25420 , \25120_25419 );
xor \U$16306 ( \25122_25421 , \25115_25414 , \25121_25420 );
buf \U$16307 ( \25123_25422 , \25122_25421 );
and \U$16308 ( \25124_25423 , \24507_24809 , \24549_24851 );
and \U$16309 ( \25125_25424 , \24507_24809 , \24569_24871 );
and \U$16310 ( \25126_25425 , \24549_24851 , \24569_24871 );
or \U$16311 ( \25127_25426 , \25124_25423 , \25125_25424 , \25126_25425 );
buf \U$16312 ( \25128_25427 , \25127_25426 );
xor \U$16313 ( \25129_25428 , \25123_25422 , \25128_25427 );
and \U$16314 ( \25130_25429 , \24535_24837 , \24540_24842 );
and \U$16315 ( \25131_25430 , \24535_24837 , \24547_24849 );
and \U$16316 ( \25132_25431 , \24540_24842 , \24547_24849 );
or \U$16317 ( \25133_25432 , \25130_25429 , \25131_25430 , \25132_25431 );
buf \U$16318 ( \25134_25433 , \25133_25432 );
and \U$16319 ( \25135_25434 , \24594_24896 , \24600_24902 );
and \U$16320 ( \25136_25435 , \24594_24896 , \24607_24909 );
and \U$16321 ( \25137_25436 , \24600_24902 , \24607_24909 );
or \U$16322 ( \25138_25437 , \25135_25434 , \25136_25435 , \25137_25436 );
buf \U$16323 ( \25139_25438 , \25138_25437 );
xor \U$16324 ( \25140_25439 , \25134_25433 , \25139_25438 );
and \U$16325 ( \25141_25440 , \12183_12157 , \21827_22129_nG9bd8 );
and \U$16326 ( \25142_25441 , \11855_12154 , \22330_22629_nG9bd5 );
or \U$16327 ( \25143_25442 , \25141_25440 , \25142_25441 );
xor \U$16328 ( \25144_25443 , \11854_12153 , \25143_25442 );
buf \U$16329 ( \25145_25444 , \25144_25443 );
buf \U$16331 ( \25146_25445 , \25145_25444 );
xor \U$16332 ( \25147_25446 , \25140_25439 , \25146_25445 );
buf \U$16333 ( \25148_25447 , \25147_25446 );
xor \U$16334 ( \25149_25448 , \25129_25428 , \25148_25447 );
buf \U$16335 ( \25150_25449 , \25149_25448 );
and \U$16336 ( \25151_25450 , \24577_24879 , \25003_25305 );
and \U$16337 ( \25152_25451 , \24577_24879 , \25009_25311 );
and \U$16338 ( \25153_25452 , \25003_25305 , \25009_25311 );
or \U$16339 ( \25154_25453 , \25151_25450 , \25152_25451 , \25153_25452 );
buf \U$16340 ( \25155_25454 , \25154_25453 );
xor \U$16341 ( \25156_25455 , \25150_25449 , \25155_25454 );
and \U$16342 ( \25157_25456 , \24609_24911 , \24615_24917 );
and \U$16343 ( \25158_25457 , \24609_24911 , \25001_25303 );
and \U$16344 ( \25159_25458 , \24615_24917 , \25001_25303 );
or \U$16345 ( \25160_25459 , \25157_25456 , \25158_25457 , \25159_25458 );
buf \U$16346 ( \25161_25460 , \25160_25459 );
and \U$16347 ( \25162_25461 , \24555_24857 , \24560_24862 );
and \U$16348 ( \25163_25462 , \24555_24857 , \24567_24869 );
and \U$16349 ( \25164_25463 , \24560_24862 , \24567_24869 );
or \U$16350 ( \25165_25464 , \25162_25461 , \25163_25462 , \25164_25463 );
buf \U$16351 ( \25166_25465 , \25165_25464 );
xor \U$16352 ( \25167_25466 , \25161_25460 , \25166_25465 );
and \U$16353 ( \25168_25467 , \10411_10707 , \24996_25298_nG9bcc );
and \U$16354 ( \25169_25468 , \24625_24927 , \24629_24931 );
and \U$16355 ( \25170_25469 , \24629_24931 , \24641_24943 );
and \U$16356 ( \25171_25470 , \24625_24927 , \24641_24943 );
or \U$16357 ( \25172_25471 , \25169_25468 , \25170_25469 , \25171_25470 );
and \U$16358 ( \25173_25472 , \24647_24949 , \24681_24983 );
and \U$16359 ( \25174_25473 , \24681_24983 , \24984_25286 );
and \U$16360 ( \25175_25474 , \24647_24949 , \24984_25286 );
or \U$16361 ( \25176_25475 , \25173_25472 , \25174_25473 , \25175_25474 );
xor \U$16362 ( \25177_25476 , \25172_25471 , \25176_25475 );
and \U$16363 ( \25178_25477 , \24686_24988 , \24964_25266 );
and \U$16364 ( \25179_25478 , \24964_25266 , \24983_25285 );
and \U$16365 ( \25180_25479 , \24686_24988 , \24983_25285 );
or \U$16366 ( \25181_25480 , \25178_25477 , \25179_25478 , \25180_25479 );
and \U$16367 ( \25182_25481 , \24634_24936 , \24638_24940 );
and \U$16368 ( \25183_25482 , \24638_24940 , \24640_24942 );
and \U$16369 ( \25184_25483 , \24634_24936 , \24640_24942 );
or \U$16370 ( \25185_25484 , \25182_25481 , \25183_25482 , \25184_25483 );
and \U$16371 ( \25186_25485 , \20242_20544 , \13755_14054 );
and \U$16372 ( \25187_25486 , \20734_21033 , \13390_13692 );
nor \U$16373 ( \25188_25487 , \25186_25485 , \25187_25486 );
xnor \U$16374 ( \25189_25488 , \25188_25487 , \13736_14035 );
and \U$16375 ( \25190_25489 , \14648_14950 , \19235_19534 );
and \U$16376 ( \25191_25490 , \15022_15321 , \18743_19045 );
nor \U$16377 ( \25192_25491 , \25190_25489 , \25191_25490 );
xnor \U$16378 ( \25193_25492 , \25192_25491 , \19241_19540 );
xor \U$16379 ( \25194_25493 , \25189_25488 , \25193_25492 );
and \U$16380 ( \25195_25494 , \13377_13679 , \20706_21005 );
and \U$16381 ( \25196_25495 , \13725_14024 , \20255_20557 );
nor \U$16382 ( \25197_25496 , \25195_25494 , \25196_25495 );
xnor \U$16383 ( \25198_25497 , \25197_25496 , \20712_21011 );
xor \U$16384 ( \25199_25498 , \25194_25493 , \25198_25497 );
xor \U$16385 ( \25200_25499 , \25185_25484 , \25199_25498 );
and \U$16386 ( \25201_25500 , \23315_23617 , \11275_11574 );
and \U$16387 ( \25202_25501 , \23900_24199 , \10976_11278 );
nor \U$16388 ( \25203_25502 , \25201_25500 , \25202_25501 );
xnor \U$16389 ( \25204_25503 , \25203_25502 , \11281_11580 );
not \U$16390 ( \25205_25504 , \24963_25265 );
and \U$16391 ( \25206_25505 , RIdec56a8_710, \9034_9333 );
and \U$16392 ( \25207_25506 , RIdec29a8_678, \9036_9335 );
and \U$16393 ( \25208_25507 , RIfc54020_5978, \9038_9337 );
and \U$16394 ( \25209_25508 , RIdebfca8_646, \9040_9339 );
and \U$16395 ( \25210_25509 , RIee1f540_4815, \9042_9341 );
and \U$16396 ( \25211_25510 , RIdebcfa8_614, \9044_9343 );
and \U$16397 ( \25212_25511 , RIdeba2a8_582, \9046_9345 );
and \U$16398 ( \25213_25512 , RIdeb75a8_550, \9048_9347 );
and \U$16399 ( \25214_25513 , RIfc4fe08_5931, \9050_9349 );
and \U$16400 ( \25215_25514 , RIdeb1ba8_486, \9052_9351 );
and \U$16401 ( \25216_25515 , RIfc6b630_6244, \9054_9353 );
and \U$16402 ( \25217_25516 , RIdeaeea8_454, \9056_9355 );
and \U$16403 ( \25218_25517 , RIfc6a118_6229, \9058_9357 );
and \U$16404 ( \25219_25518 , RIdeaaab0_422, \9060_9359 );
and \U$16405 ( \25220_25519 , RIdea41b0_390, \9062_9361 );
and \U$16406 ( \25221_25520 , RIde9d8b0_358, \9064_9363 );
and \U$16407 ( \25222_25521 , RIfc69ce0_6226, \9066_9365 );
and \U$16408 ( \25223_25522 , RIee1be68_4776, \9068_9367 );
and \U$16409 ( \25224_25523 , RIfc653c0_6174, \9070_9369 );
and \U$16410 ( \25225_25524 , RIee1ac20_4763, \9072_9371 );
and \U$16411 ( \25226_25525 , RIde91718_299, \9074_9373 );
and \U$16412 ( \25227_25526 , RIde8df50_282, \9076_9375 );
and \U$16413 ( \25228_25527 , RIde89db0_262, \9078_9377 );
and \U$16414 ( \25229_25528 , RIde85c10_242, \9080_9379 );
and \U$16415 ( \25230_25529 , RIde81db8_223, \9082_9381 );
and \U$16416 ( \25231_25530 , RIfca76a8_6927, \9084_9383 );
and \U$16417 ( \25232_25531 , RIfcca4f0_7324, \9086_9385 );
and \U$16418 ( \25233_25532 , RIfc4ce38_5897, \9088_9387 );
and \U$16419 ( \25234_25533 , RIfc6b360_6242, \9090_9389 );
and \U$16420 ( \25235_25534 , RIe16b918_2601, \9092_9391 );
and \U$16421 ( \25236_25535 , RIe169cf8_2581, \9094_9393 );
and \U$16422 ( \25237_25536 , RIe167f70_2560, \9096_9395 );
and \U$16423 ( \25238_25537 , RIe1656a8_2531, \9098_9397 );
and \U$16424 ( \25239_25538 , RIe1629a8_2499, \9100_9399 );
and \U$16425 ( \25240_25539 , RIee37690_5089, \9102_9401 );
and \U$16426 ( \25241_25540 , RIe15fca8_2467, \9104_9403 );
and \U$16427 ( \25242_25541 , RIfce93f0_7676, \9106_9405 );
and \U$16428 ( \25243_25542 , RIe15cfa8_2435, \9108_9407 );
and \U$16429 ( \25244_25543 , RIe1575a8_2371, \9110_9409 );
and \U$16430 ( \25245_25544 , RIe1548a8_2339, \9112_9411 );
and \U$16431 ( \25246_25545 , RIee35908_5068, \9114_9413 );
and \U$16432 ( \25247_25546 , RIe151ba8_2307, \9116_9415 );
and \U$16433 ( \25248_25547 , RIee34f30_5061, \9118_9417 );
and \U$16434 ( \25249_25548 , RIe14eea8_2275, \9120_9419 );
and \U$16435 ( \25250_25549 , RIfce32e8_7607, \9122_9421 );
and \U$16436 ( \25251_25550 , RIe14c1a8_2243, \9124_9423 );
and \U$16437 ( \25252_25551 , RIe1494a8_2211, \9126_9425 );
and \U$16438 ( \25253_25552 , RIe1467a8_2179, \9128_9427 );
and \U$16439 ( \25254_25553 , RIfcde2c0_7550, \9130_9429 );
and \U$16440 ( \25255_25554 , RIfc687c8_6211, \9132_9431 );
and \U$16441 ( \25256_25555 , RIfca9160_6946, \9134_9433 );
and \U$16442 ( \25257_25556 , RIfcb1590_7040, \9136_9435 );
and \U$16443 ( \25258_25557 , RIe141078_2117, \9138_9437 );
and \U$16444 ( \25259_25558 , RIdf3ef80_2093, \9140_9439 );
and \U$16445 ( \25260_25559 , RIdf3cdc0_2069, \9142_9441 );
and \U$16446 ( \25261_25560 , RIfebeb60_8290, \9144_9443 );
and \U$16447 ( \25262_25561 , RIfc64448_6163, \9146_9445 );
and \U$16448 ( \25263_25562 , RIee2fad0_5001, \9148_9447 );
and \U$16449 ( \25264_25563 , RIfca7978_6929, \9150_9449 );
and \U$16450 ( \25265_25564 , RIfc676e8_6199, \9152_9451 );
and \U$16451 ( \25266_25565 , RIdf35a70_1987, \9154_9453 );
and \U$16452 ( \25267_25566 , RIdf335e0_1961, \9156_9455 );
and \U$16453 ( \25268_25567 , RIdf31420_1937, \9158_9457 );
and \U$16454 ( \25269_25568 , RIdf2f3c8_1914, \9160_9459 );
or \U$16455 ( \25270_25569 , \25206_25505 , \25207_25506 , \25208_25507 , \25209_25508 , \25210_25509 , \25211_25510 , \25212_25511 , \25213_25512 , \25214_25513 , \25215_25514 , \25216_25515 , \25217_25516 , \25218_25517 , \25219_25518 , \25220_25519 , \25221_25520 , \25222_25521 , \25223_25522 , \25224_25523 , \25225_25524 , \25226_25525 , \25227_25526 , \25228_25527 , \25229_25528 , \25230_25529 , \25231_25530 , \25232_25531 , \25233_25532 , \25234_25533 , \25235_25534 , \25236_25535 , \25237_25536 , \25238_25537 , \25239_25538 , \25240_25539 , \25241_25540 , \25242_25541 , \25243_25542 , \25244_25543 , \25245_25544 , \25246_25545 , \25247_25546 , \25248_25547 , \25249_25548 , \25250_25549 , \25251_25550 , \25252_25551 , \25253_25552 , \25254_25553 , \25255_25554 , \25256_25555 , \25257_25556 , \25258_25557 , \25259_25558 , \25260_25559 , \25261_25560 , \25262_25561 , \25263_25562 , \25264_25563 , \25265_25564 , \25266_25565 , \25267_25566 , \25268_25567 , \25269_25568 );
and \U$16456 ( \25271_25570 , RIfccef78_7377, \9163_9462 );
and \U$16457 ( \25272_25571 , RIfca6fa0_6922, \9165_9464 );
and \U$16458 ( \25273_25572 , RIfc62558_6141, \9167_9466 );
and \U$16459 ( \25274_25573 , RIfc61fb8_6137, \9169_9468 );
and \U$16460 ( \25275_25574 , RIfe81b70_7820, \9171_9470 );
and \U$16461 ( \25276_25575 , RIdf281e0_1833, \9173_9472 );
and \U$16462 ( \25277_25576 , RIfe81cd8_7821, \9175_9474 );
and \U$16463 ( \25278_25577 , RIdf249a0_1793, \9177_9476 );
and \U$16464 ( \25279_25578 , RIfc44300_5798, \9179_9478 );
and \U$16465 ( \25280_25579 , RIfcafc40_7022, \9181_9480 );
and \U$16466 ( \25281_25580 , RIdf22ee8_1774, \9183_9482 );
and \U$16467 ( \25282_25581 , RIfcaac18_6965, \9185_9484 );
and \U$16468 ( \25283_25582 , RIdf219d0_1759, \9187_9486 );
and \U$16469 ( \25284_25583 , RIdf1fae0_1737, \9189_9488 );
and \U$16470 ( \25285_25584 , RIdf1b1c0_1685, \9191_9490 );
and \U$16471 ( \25286_25585 , RIdf19438_1664, \9193_9492 );
and \U$16472 ( \25287_25586 , RIdf17278_1640, \9195_9494 );
and \U$16473 ( \25288_25587 , RIdf14578_1608, \9197_9496 );
and \U$16474 ( \25289_25588 , RIdf11878_1576, \9199_9498 );
and \U$16475 ( \25290_25589 , RIdf0eb78_1544, \9201_9500 );
and \U$16476 ( \25291_25590 , RIdf0be78_1512, \9203_9502 );
and \U$16477 ( \25292_25591 , RIdf09178_1480, \9205_9504 );
and \U$16478 ( \25293_25592 , RIdf06478_1448, \9207_9506 );
and \U$16479 ( \25294_25593 , RIdf03778_1416, \9209_9508 );
and \U$16480 ( \25295_25594 , RIdefdd78_1352, \9211_9510 );
and \U$16481 ( \25296_25595 , RIdefb078_1320, \9213_9512 );
and \U$16482 ( \25297_25596 , RIdef8378_1288, \9215_9514 );
and \U$16483 ( \25298_25597 , RIdef5678_1256, \9217_9516 );
and \U$16484 ( \25299_25598 , RIdef2978_1224, \9219_9518 );
and \U$16485 ( \25300_25599 , RIdeefc78_1192, \9221_9520 );
and \U$16486 ( \25301_25600 , RIdeecf78_1160, \9223_9522 );
and \U$16487 ( \25302_25601 , RIdeea278_1128, \9225_9524 );
and \U$16488 ( \25303_25602 , RIfc611a8_6127, \9227_9526 );
and \U$16489 ( \25304_25603 , RIfc61a18_6133, \9229_9528 );
and \U$16490 ( \25305_25604 , RIfca65c8_6915, \9231_9530 );
and \U$16491 ( \25306_25605 , RIfca6b68_6919, \9233_9532 );
and \U$16492 ( \25307_25606 , RIdee4b48_1066, \9235_9534 );
and \U$16493 ( \25308_25607 , RIdee2dc0_1045, \9237_9536 );
and \U$16494 ( \25309_25608 , RIdee0c00_1021, \9239_9538 );
and \U$16495 ( \25310_25609 , RIdedeba8_998, \9241_9540 );
and \U$16496 ( \25311_25610 , RIfc626c0_6142, \9243_9542 );
and \U$16497 ( \25312_25611 , RIfc738f8_6337, \9245_9544 );
and \U$16498 ( \25313_25612 , RIfcb31b0_7060, \9247_9546 );
and \U$16499 ( \25314_25613 , RIee21430_4837, \9249_9548 );
and \U$16500 ( \25315_25614 , RIded9a18_940, \9251_9550 );
and \U$16501 ( \25316_25615 , RIded7588_914, \9253_9552 );
and \U$16502 ( \25317_25616 , RIded5698_892, \9255_9554 );
and \U$16503 ( \25318_25617 , RIded30a0_865, \9257_9556 );
and \U$16504 ( \25319_25618 , RIded0aa8_838, \9259_9558 );
and \U$16505 ( \25320_25619 , RIdecdda8_806, \9261_9560 );
and \U$16506 ( \25321_25620 , RIdecb0a8_774, \9263_9562 );
and \U$16507 ( \25322_25621 , RIdec83a8_742, \9265_9564 );
and \U$16508 ( \25323_25622 , RIdeb48a8_518, \9267_9566 );
and \U$16509 ( \25324_25623 , RIde96fb0_326, \9269_9568 );
and \U$16510 ( \25325_25624 , RIe16e4b0_2632, \9271_9570 );
and \U$16511 ( \25326_25625 , RIe15a2a8_2403, \9273_9572 );
and \U$16512 ( \25327_25626 , RIe143aa8_2147, \9275_9574 );
and \U$16513 ( \25328_25627 , RIdf384a0_2017, \9277_9576 );
and \U$16514 ( \25329_25628 , RIdf2cb00_1885, \9279_9578 );
and \U$16515 ( \25330_25629 , RIdf1d380_1709, \9281_9580 );
and \U$16516 ( \25331_25630 , RIdf00a78_1384, \9283_9582 );
and \U$16517 ( \25332_25631 , RIdee7578_1096, \9285_9584 );
and \U$16518 ( \25333_25632 , RIdedc2e0_969, \9287_9586 );
and \U$16519 ( \25334_25633 , RIde7cef8_199, \9289_9588 );
or \U$16520 ( \25335_25634 , \25271_25570 , \25272_25571 , \25273_25572 , \25274_25573 , \25275_25574 , \25276_25575 , \25277_25576 , \25278_25577 , \25279_25578 , \25280_25579 , \25281_25580 , \25282_25581 , \25283_25582 , \25284_25583 , \25285_25584 , \25286_25585 , \25287_25586 , \25288_25587 , \25289_25588 , \25290_25589 , \25291_25590 , \25292_25591 , \25293_25592 , \25294_25593 , \25295_25594 , \25296_25595 , \25297_25596 , \25298_25597 , \25299_25598 , \25300_25599 , \25301_25600 , \25302_25601 , \25303_25602 , \25304_25603 , \25305_25604 , \25306_25605 , \25307_25606 , \25308_25607 , \25309_25608 , \25310_25609 , \25311_25610 , \25312_25611 , \25313_25612 , \25314_25613 , \25315_25614 , \25316_25615 , \25317_25616 , \25318_25617 , \25319_25618 , \25320_25619 , \25321_25620 , \25322_25621 , \25323_25622 , \25324_25623 , \25325_25624 , \25326_25625 , \25327_25626 , \25328_25627 , \25329_25628 , \25330_25629 , \25331_25630 , \25332_25631 , \25333_25632 , \25334_25633 );
or \U$16521 ( \25336_25635 , \25270_25569 , \25335_25634 );
_DC \g5ca9/U$1 ( \25337 , \25336_25635 , \9298_9597 );
and \U$16522 ( \25338_25637 , RIe19d940_3170, \8760_9059 );
and \U$16523 ( \25339_25638 , RIe19ac40_3138, \8762_9061 );
and \U$16524 ( \25340_25639 , RIfc64880_6166, \8764_9063 );
and \U$16525 ( \25341_25640 , RIe197f40_3106, \8766_9065 );
and \U$16526 ( \25342_25641 , RIf144848_5239, \8768_9067 );
and \U$16527 ( \25343_25642 , RIe195240_3074, \8770_9069 );
and \U$16528 ( \25344_25643 , RIe192540_3042, \8772_9071 );
and \U$16529 ( \25345_25644 , RIe18f840_3010, \8774_9073 );
and \U$16530 ( \25346_25645 , RIe189e40_2946, \8776_9075 );
and \U$16531 ( \25347_25646 , RIe187140_2914, \8778_9077 );
and \U$16532 ( \25348_25647 , RIf143a38_5229, \8780_9079 );
and \U$16533 ( \25349_25648 , RIe184440_2882, \8782_9081 );
and \U$16534 ( \25350_25649 , RIfc6f140_6286, \8784_9083 );
and \U$16535 ( \25351_25650 , RIe181740_2850, \8786_9085 );
and \U$16536 ( \25352_25651 , RIe17ea40_2818, \8788_9087 );
and \U$16537 ( \25353_25652 , RIe17bd40_2786, \8790_9089 );
and \U$16538 ( \25354_25653 , RIfc64f88_6171, \8792_9091 );
and \U$16539 ( \25355_25654 , RIf141008_5199, \8794_9093 );
and \U$16540 ( \25356_25655 , RIe177150_2732, \8796_9095 );
and \U$16541 ( \25357_25656 , RIfe81738_7817, \8798_9097 );
and \U$16542 ( \25358_25657 , RIfccabf8_7329, \8800_9099 );
and \U$16543 ( \25359_25658 , RIf13f3e8_5179, \8802_9101 );
and \U$16544 ( \25360_25659 , RIfca81e8_6935, \8804_9103 );
and \U$16545 ( \25361_25660 , RIee3d630_5157, \8806_9105 );
and \U$16546 ( \25362_25661 , RIfc66068_6183, \8808_9107 );
and \U$16547 ( \25363_25662 , RIfc6ed08_6283, \8810_9109 );
and \U$16548 ( \25364_25663 , RIfcdde88_7547, \8812_9111 );
and \U$16549 ( \25365_25664 , RIe173a78_2693, \8814_9113 );
and \U$16550 ( \25366_25665 , RIfc66338_6185, \8816_9115 );
and \U$16551 ( \25367_25666 , RIfc6eba0_6282, \8818_9117 );
and \U$16552 ( \25368_25667 , RIfc664a0_6186, \8820_9119 );
and \U$16553 ( \25369_25668 , RIfcacdd8_6989, \8822_9121 );
and \U$16554 ( \25370_25669 , RIfe81468_7815, \8824_9123 );
and \U$16555 ( \25371_25670 , RIe223c98_4697, \8826_9125 );
and \U$16556 ( \25372_25671 , RIfc66d10_6192, \8828_9127 );
and \U$16557 ( \25373_25672 , RIe220f98_4665, \8830_9129 );
and \U$16558 ( \25374_25673 , RIf16b038_5677, \8832_9131 );
and \U$16559 ( \25375_25674 , RIe21e298_4633, \8834_9133 );
and \U$16560 ( \25376_25675 , RIe218898_4569, \8836_9135 );
and \U$16561 ( \25377_25676 , RIe215b98_4537, \8838_9137 );
and \U$16562 ( \25378_25677 , RIfc3fc38_5751, \8840_9139 );
and \U$16563 ( \25379_25678 , RIe212e98_4505, \8842_9141 );
and \U$16564 ( \25380_25679 , RIfc67850_6200, \8844_9143 );
and \U$16565 ( \25381_25680 , RIe210198_4473, \8846_9145 );
and \U$16566 ( \25382_25681 , RIf167f00_5642, \8848_9147 );
and \U$16567 ( \25383_25682 , RIe20d498_4441, \8850_9149 );
and \U$16568 ( \25384_25683 , RIe20a798_4409, \8852_9151 );
and \U$16569 ( \25385_25684 , RIe207a98_4377, \8854_9153 );
and \U$16570 ( \25386_25685 , RIfcacb08_6987, \8856_9155 );
and \U$16571 ( \25387_25686 , RIfcac9a0_6986, \8858_9157 );
and \U$16572 ( \25388_25687 , RIfea8900_8234, \8860_9159 );
and \U$16573 ( \25389_25688 , RIfe818a0_7818, \8862_9161 );
and \U$16574 ( \25390_25689 , RIfca8a58_6941, \8864_9163 );
and \U$16575 ( \25391_25690 , RIfccad60_7330, \8866_9165 );
and \U$16576 ( \25392_25691 , RIfcac838_6985, \8868_9167 );
and \U$16577 ( \25393_25692 , RIfc67418_6197, \8870_9169 );
and \U$16578 ( \25394_25693 , RIf160340_5554, \8872_9171 );
and \U$16579 ( \25395_25694 , RIf15e450_5532, \8874_9173 );
and \U$16580 ( \25396_25695 , RIfe81a08_7819, \8876_9175 );
and \U$16581 ( \25397_25696 , RIfe81300_7814, \8878_9177 );
and \U$16582 ( \25398_25697 , RIfc6dac0_6270, \8880_9179 );
and \U$16583 ( \25399_25698 , RIf15ba20_5502, \8882_9181 );
and \U$16584 ( \25400_25699 , RIfc6d958_6269, \8884_9183 );
and \U$16585 ( \25401_25700 , RIfc6d7f0_6268, \8886_9185 );
or \U$16586 ( \25402_25701 , \25338_25637 , \25339_25638 , \25340_25639 , \25341_25640 , \25342_25641 , \25343_25642 , \25344_25643 , \25345_25644 , \25346_25645 , \25347_25646 , \25348_25647 , \25349_25648 , \25350_25649 , \25351_25650 , \25352_25651 , \25353_25652 , \25354_25653 , \25355_25654 , \25356_25655 , \25357_25656 , \25358_25657 , \25359_25658 , \25360_25659 , \25361_25660 , \25362_25661 , \25363_25662 , \25364_25663 , \25365_25664 , \25366_25665 , \25367_25666 , \25368_25667 , \25369_25668 , \25370_25669 , \25371_25670 , \25372_25671 , \25373_25672 , \25374_25673 , \25375_25674 , \25376_25675 , \25377_25676 , \25378_25677 , \25379_25678 , \25380_25679 , \25381_25680 , \25382_25681 , \25383_25682 , \25384_25683 , \25385_25684 , \25386_25685 , \25387_25686 , \25388_25687 , \25389_25688 , \25390_25689 , \25391_25690 , \25392_25691 , \25393_25692 , \25394_25693 , \25395_25694 , \25396_25695 , \25397_25696 , \25398_25697 , \25399_25698 , \25400_25699 , \25401_25700 );
and \U$16587 ( \25403_25702 , RIfc587d8_6029, \8889_9188 );
and \U$16588 ( \25404_25703 , RIfc6cf80_6262, \8891_9190 );
and \U$16589 ( \25405_25704 , RIfc6d3b8_6265, \8893_9192 );
and \U$16590 ( \25406_25705 , RIfe815d0_7816, \8895_9194 );
and \U$16591 ( \25407_25706 , RIfc6d520_6266, \8897_9196 );
and \U$16592 ( \25408_25707 , RIfcabe60_6978, \8899_9198 );
and \U$16593 ( \25409_25708 , RIfc6d0e8_6263, \8901_9200 );
and \U$16594 ( \25410_25709 , RIe1f5780_4170, \8903_9202 );
and \U$16595 ( \25411_25710 , RIfc6c5a8_6255, \8905_9204 );
and \U$16596 ( \25412_25711 , RIfc68d68_6215, \8907_9206 );
and \U$16597 ( \25413_25712 , RIfc68c00_6214, \8909_9208 );
and \U$16598 ( \25414_25713 , RIe1f3458_4145, \8911_9210 );
and \U$16599 ( \25415_25714 , RIfc68a98_6213, \8913_9212 );
and \U$16600 ( \25416_25715 , RIfccb8a0_7338, \8915_9214 );
and \U$16601 ( \25417_25716 , RIfca9b38_6953, \8917_9216 );
and \U$16602 ( \25418_25717 , RIe1ee160_4086, \8919_9218 );
and \U$16603 ( \25419_25718 , RIe1eba00_4058, \8921_9220 );
and \U$16604 ( \25420_25719 , RIe1e8d00_4026, \8923_9222 );
and \U$16605 ( \25421_25720 , RIe1e6000_3994, \8925_9224 );
and \U$16606 ( \25422_25721 , RIe1e3300_3962, \8927_9226 );
and \U$16607 ( \25423_25722 , RIe1e0600_3930, \8929_9228 );
and \U$16608 ( \25424_25723 , RIe1dd900_3898, \8931_9230 );
and \U$16609 ( \25425_25724 , RIe1dac00_3866, \8933_9232 );
and \U$16610 ( \25426_25725 , RIe1d7f00_3834, \8935_9234 );
and \U$16611 ( \25427_25726 , RIe1d2500_3770, \8937_9236 );
and \U$16612 ( \25428_25727 , RIe1cf800_3738, \8939_9238 );
and \U$16613 ( \25429_25728 , RIe1ccb00_3706, \8941_9240 );
and \U$16614 ( \25430_25729 , RIe1c9e00_3674, \8943_9242 );
and \U$16615 ( \25431_25730 , RIe1c7100_3642, \8945_9244 );
and \U$16616 ( \25432_25731 , RIe1c4400_3610, \8947_9246 );
and \U$16617 ( \25433_25732 , RIe1c1700_3578, \8949_9248 );
and \U$16618 ( \25434_25733 , RIe1bea00_3546, \8951_9250 );
and \U$16619 ( \25435_25734 , RIfc6bbd0_6248, \8953_9252 );
and \U$16620 ( \25436_25735 , RIfcdd348_7539, \8955_9254 );
and \U$16621 ( \25437_25736 , RIe1b9438_3485, \8957_9256 );
and \U$16622 ( \25438_25737 , RIe1b73e0_3462, \8959_9258 );
and \U$16623 ( \25439_25738 , RIfcab5f0_6972, \8961_9260 );
and \U$16624 ( \25440_25739 , RIfccbb70_7340, \8963_9262 );
and \U$16625 ( \25441_25740 , RIe1b5220_3438, \8965_9264 );
and \U$16626 ( \25442_25741 , RIe1b3e70_3424, \8967_9266 );
and \U$16627 ( \25443_25742 , RIfc6c9e0_6258, \8969_9268 );
and \U$16628 ( \25444_25743 , RIfcab488_6971, \8971_9270 );
and \U$16629 ( \25445_25744 , RIfea7dc0_8226, \8973_9272 );
and \U$16630 ( \25446_25745 , RIe1b0bd0_3388, \8975_9274 );
and \U$16631 ( \25447_25746 , RIfc6ce18_6261, \8977_9276 );
and \U$16632 ( \25448_25747 , RIfcabfc8_6979, \8979_9278 );
and \U$16633 ( \25449_25748 , RIe1ac580_3338, \8981_9280 );
and \U$16634 ( \25450_25749 , RIe1aaf00_3322, \8983_9282 );
and \U$16635 ( \25451_25750 , RIe1a8d40_3298, \8985_9284 );
and \U$16636 ( \25452_25751 , RIe1a6040_3266, \8987_9286 );
and \U$16637 ( \25453_25752 , RIe1a3340_3234, \8989_9288 );
and \U$16638 ( \25454_25753 , RIe1a0640_3202, \8991_9290 );
and \U$16639 ( \25455_25754 , RIe18cb40_2978, \8993_9292 );
and \U$16640 ( \25456_25755 , RIe179040_2754, \8995_9294 );
and \U$16641 ( \25457_25756 , RIe226998_4729, \8997_9296 );
and \U$16642 ( \25458_25757 , RIe21b598_4601, \8999_9298 );
and \U$16643 ( \25459_25758 , RIe204d98_4345, \9001_9300 );
and \U$16644 ( \25460_25759 , RIe1fedf8_4277, \9003_9302 );
and \U$16645 ( \25461_25760 , RIe1f81b0_4200, \9005_9304 );
and \U$16646 ( \25462_25761 , RIe1f0cf8_4117, \9007_9306 );
and \U$16647 ( \25463_25762 , RIe1d5200_3802, \9009_9308 );
and \U$16648 ( \25464_25763 , RIe1bbd00_3514, \9011_9310 );
and \U$16649 ( \25465_25764 , RIe1aeb78_3365, \9013_9312 );
and \U$16650 ( \25466_25765 , RIe1711b0_2664, \9015_9314 );
or \U$16651 ( \25467_25766 , \25403_25702 , \25404_25703 , \25405_25704 , \25406_25705 , \25407_25706 , \25408_25707 , \25409_25708 , \25410_25709 , \25411_25710 , \25412_25711 , \25413_25712 , \25414_25713 , \25415_25714 , \25416_25715 , \25417_25716 , \25418_25717 , \25419_25718 , \25420_25719 , \25421_25720 , \25422_25721 , \25423_25722 , \25424_25723 , \25425_25724 , \25426_25725 , \25427_25726 , \25428_25727 , \25429_25728 , \25430_25729 , \25431_25730 , \25432_25731 , \25433_25732 , \25434_25733 , \25435_25734 , \25436_25735 , \25437_25736 , \25438_25737 , \25439_25738 , \25440_25739 , \25441_25740 , \25442_25741 , \25443_25742 , \25444_25743 , \25445_25744 , \25446_25745 , \25447_25746 , \25448_25747 , \25449_25748 , \25450_25749 , \25451_25750 , \25452_25751 , \25453_25752 , \25454_25753 , \25455_25754 , \25456_25755 , \25457_25756 , \25458_25757 , \25459_25758 , \25460_25759 , \25461_25760 , \25462_25761 , \25463_25762 , \25464_25763 , \25465_25764 , \25466_25765 );
or \U$16652 ( \25468_25767 , \25402_25701 , \25467_25766 );
_DC \g5d2d/U$1 ( \25469 , \25468_25767 , \9024_9323 );
xor g5d2e_GF_PartitionCandidate( \25470_25769_nG5d2e , \25337 , \25469 );
buf \U$16653 ( \25471_25770 , \25470_25769_nG5d2e );
and \U$16654 ( \25472_25771 , \24961_25263 , \23836_24135 );
not \U$16655 ( \25473_25772 , \25472_25771 );
and \U$16656 ( \25474_25773 , \25471_25770 , \25473_25772 );
and \U$16657 ( \25475_25774 , \25205_25504 , \25474_25773 );
xor \U$16658 ( \25476_25775 , \25204_25503 , \25475_25774 );
and \U$16659 ( \25477_25776 , \17325_17627 , \16333_16635 );
and \U$16660 ( \25478_25777 , \17736_18035 , \15999_16301 );
nor \U$16661 ( \25479_25778 , \25477_25776 , \25478_25777 );
xnor \U$16662 ( \25480_25779 , \25479_25778 , \16323_16625 );
xor \U$16663 ( \25481_25780 , \25476_25775 , \25480_25779 );
and \U$16664 ( \25482_25781 , \15965_16267 , \17791_18090 );
and \U$16665 ( \25483_25782 , \16353_16655 , \17353_17655 );
nor \U$16666 ( \25484_25783 , \25482_25781 , \25483_25782 );
xnor \U$16667 ( \25485_25784 , \25484_25783 , \17747_18046 );
xor \U$16668 ( \25486_25785 , \25481_25780 , \25485_25784 );
xor \U$16669 ( \25487_25786 , \25200_25499 , \25486_25785 );
xor \U$16670 ( \25488_25787 , \25181_25480 , \25487_25786 );
and \U$16671 ( \25489_25788 , \24651_24953 , \24665_24967 );
and \U$16672 ( \25490_25789 , \24665_24967 , \24680_24982 );
and \U$16673 ( \25491_25790 , \24651_24953 , \24680_24982 );
or \U$16674 ( \25492_25791 , \25489_25788 , \25490_25789 , \25491_25790 );
and \U$16675 ( \25493_25792 , \24690_24992 , \24694_24996 );
and \U$16676 ( \25494_25793 , \24694_24996 , \24963_25265 );
and \U$16677 ( \25495_25794 , \24690_24992 , \24963_25265 );
or \U$16678 ( \25496_25795 , \25493_25792 , \25494_25793 , \25495_25794 );
and \U$16679 ( \25497_25796 , \24973_25275 , \24977_25279 );
and \U$16680 ( \25498_25797 , \24977_25279 , \24982_25284 );
and \U$16681 ( \25499_25798 , \24973_25275 , \24982_25284 );
or \U$16682 ( \25500_25799 , \25497_25796 , \25498_25797 , \25499_25798 );
xor \U$16683 ( \25501_25800 , \25496_25795 , \25500_25799 );
and \U$16684 ( \25502_25801 , \24670_24972 , \24674_24976 );
and \U$16685 ( \25503_25802 , \24674_24976 , \24679_24981 );
and \U$16686 ( \25504_25803 , \24670_24972 , \24679_24981 );
or \U$16687 ( \25505_25804 , \25502_25801 , \25503_25802 , \25504_25803 );
xor \U$16688 ( \25506_25805 , \25501_25800 , \25505_25804 );
xor \U$16689 ( \25507_25806 , \25492_25791 , \25506_25805 );
and \U$16690 ( \25508_25807 , \24655_24957 , \24659_24961 );
and \U$16691 ( \25509_25808 , \24659_24961 , \24664_24966 );
and \U$16692 ( \25510_25809 , \24655_24957 , \24664_24966 );
or \U$16693 ( \25511_25810 , \25508_25807 , \25509_25808 , \25510_25809 );
and \U$16694 ( \25512_25811 , \24970_25272 , \10681_10983 );
_DC \g65bc/U$1 ( \25513 , \25336_25635 , \9298_9597 );
_DC \g65bd/U$1 ( \25514 , \25468_25767 , \9024_9323 );
and g65be_GF_PartitionCandidate( \25515_25814_nG65be , \25513 , \25514 );
buf \U$16695 ( \25516_25815 , \25515_25814_nG65be );
and \U$16696 ( \25517_25816 , \25516_25815 , \10389_10691 );
nor \U$16697 ( \25518_25817 , \25512_25811 , \25517_25816 );
xnor \U$16698 ( \25519_25818 , \25518_25817 , \10678_10980 );
and \U$16699 ( \25520_25819 , \21788_22090 , \12491_12790 );
and \U$16700 ( \25521_25820 , \22257_22556 , \12159_12461 );
nor \U$16701 ( \25522_25821 , \25520_25819 , \25521_25820 );
xnor \U$16702 ( \25523_25822 , \25522_25821 , \12481_12780 );
xor \U$16703 ( \25524_25823 , \25519_25818 , \25523_25822 );
xor \U$16704 ( \25525_25824 , \25471_25770 , \24961_25263 );
not \U$16705 ( \25526_25825 , \24962_25264 );
and \U$16706 ( \25527_25826 , \25525_25824 , \25526_25825 );
and \U$16707 ( \25528_25827 , \10385_10687 , \25527_25826 );
and \U$16708 ( \25529_25828 , \10686_10988 , \24962_25264 );
nor \U$16709 ( \25530_25829 , \25528_25827 , \25529_25828 );
xnor \U$16710 ( \25531_25830 , \25530_25829 , \25474_25773 );
xor \U$16711 ( \25532_25831 , \25524_25823 , \25531_25830 );
xor \U$16712 ( \25533_25832 , \25511_25810 , \25532_25831 );
and \U$16713 ( \25534_25833 , \18730_19032 , \15037_15336 );
and \U$16714 ( \25535_25834 , \19259_19558 , \14661_14963 );
nor \U$16715 ( \25536_25835 , \25534_25833 , \25535_25834 );
xnor \U$16716 ( \25537_25836 , \25536_25835 , \15043_15342 );
and \U$16717 ( \25538_25837 , \12146_12448 , \22243_22542 );
and \U$16718 ( \25539_25838 , \12470_12769 , \21801_22103 );
nor \U$16719 ( \25540_25839 , \25538_25837 , \25539_25838 );
xnor \U$16720 ( \25541_25840 , \25540_25839 , \22249_22548 );
xor \U$16721 ( \25542_25841 , \25537_25836 , \25541_25840 );
and \U$16722 ( \25543_25842 , \10968_11270 , \23839_24138 );
and \U$16723 ( \25544_25843 , \11287_11586 , \23328_23630 );
nor \U$16724 ( \25545_25844 , \25543_25842 , \25544_25843 );
xnor \U$16725 ( \25546_25845 , \25545_25844 , \23845_24144 );
xor \U$16726 ( \25547_25846 , \25542_25841 , \25546_25845 );
xor \U$16727 ( \25548_25847 , \25533_25832 , \25547_25846 );
xor \U$16728 ( \25549_25848 , \25507_25806 , \25548_25847 );
xor \U$16729 ( \25550_25849 , \25488_25787 , \25549_25848 );
xor \U$16730 ( \25551_25850 , \25177_25476 , \25550_25849 );
and \U$16731 ( \25552_25851 , \24621_24923 , \24642_24944 );
and \U$16732 ( \25553_25852 , \24642_24944 , \24985_25287 );
and \U$16733 ( \25554_25853 , \24621_24923 , \24985_25287 );
or \U$16734 ( \25555_25854 , \25552_25851 , \25553_25852 , \25554_25853 );
xor \U$16735 ( \25556_25855 , \25551_25850 , \25555_25854 );
and \U$16736 ( \25557_25856 , \24986_25288 , \24990_25292 );
and \U$16737 ( \25558_25857 , \24991_25293 , \24994_25296 );
or \U$16738 ( \25559_25858 , \25557_25856 , \25558_25857 );
xor \U$16739 ( \25560_25859 , \25556_25855 , \25559_25858 );
buf g9bc9_GF_PartitionCandidate( \25561_25860_nG9bc9 , \25560_25859 );
and \U$16740 ( \25562_25861 , \10402_10704 , \25561_25860_nG9bc9 );
or \U$16741 ( \25563_25862 , \25168_25467 , \25562_25861 );
xor \U$16742 ( \25564_25863 , \10399_10703 , \25563_25862 );
buf \U$16743 ( \25565_25864 , \25564_25863 );
buf \U$16745 ( \25566_25865 , \25565_25864 );
xor \U$16746 ( \25567_25866 , \25167_25466 , \25566_25865 );
buf \U$16747 ( \25568_25867 , \25567_25866 );
xor \U$16748 ( \25569_25868 , \25156_25455 , \25568_25867 );
xor \U$16749 ( \25570_25869 , \25025_25327 , \25569_25868 );
and \U$16750 ( \25571_25870 , \24502_24804 , \24571_24873 );
and \U$16751 ( \25572_25871 , \24502_24804 , \25011_25313 );
and \U$16752 ( \25573_25872 , \24571_24873 , \25011_25313 );
or \U$16753 ( \25574_25873 , \25571_25870 , \25572_25871 , \25573_25872 );
and \U$16754 ( \25575_25874 , \25570_25869 , \25574_25873 );
and \U$16755 ( \25576_25875 , \25020_25322 , \25024_25326 );
and \U$16756 ( \25577_25876 , \25020_25322 , \25569_25868 );
and \U$16757 ( \25578_25877 , \25024_25326 , \25569_25868 );
or \U$16758 ( \25579_25878 , \25576_25875 , \25577_25876 , \25578_25877 );
xor \U$16759 ( \25580_25879 , \25575_25874 , \25579_25878 );
and \U$16760 ( \25581_25880 , RIdec5978_712, \8760_9059 );
and \U$16761 ( \25582_25881 , RIdec2c78_680, \8762_9061 );
and \U$16762 ( \25583_25882 , RIfc8aad0_6600, \8764_9063 );
and \U$16763 ( \25584_25883 , RIdebff78_648, \8766_9065 );
and \U$16764 ( \25585_25884 , RIfc8ac38_6601, \8768_9067 );
and \U$16765 ( \25586_25885 , RIdebd278_616, \8770_9069 );
and \U$16766 ( \25587_25886 , RIdeba578_584, \8772_9071 );
and \U$16767 ( \25588_25887 , RIdeb7878_552, \8774_9073 );
and \U$16768 ( \25589_25888 , RIfc40e80_5764, \8776_9075 );
and \U$16769 ( \25590_25889 , RIdeb1e78_488, \8778_9077 );
and \U$16770 ( \25591_25890 , RIfcdaeb8_7513, \8780_9079 );
and \U$16771 ( \25592_25891 , RIdeaf178_456, \8782_9081 );
and \U$16772 ( \25593_25892 , RIee1dbf0_4797, \8784_9083 );
and \U$16773 ( \25594_25893 , RIdeab140_424, \8786_9085 );
and \U$16774 ( \25595_25894 , RIdea4840_392, \8788_9087 );
and \U$16775 ( \25596_25895 , RIde9df40_360, \8790_9089 );
and \U$16776 ( \25597_25896 , RIfc8b070_6604, \8792_9091 );
and \U$16777 ( \25598_25897 , RIfcc38a8_7247, \8794_9093 );
and \U$16778 ( \25599_25898 , RIfc807b0_6484, \8796_9095 );
and \U$16779 ( \25600_25899 , RIfcbb8b0_7156, \8798_9097 );
and \U$16780 ( \25601_25900 , RIde91a60_300, \8800_9099 );
and \U$16781 ( \25602_25901 , RIde8e298_283, \8802_9101 );
and \U$16782 ( \25603_25902 , RIde8a440_264, \8804_9103 );
and \U$16783 ( \25604_25903 , RIde862a0_244, \8806_9105 );
and \U$16784 ( \25605_25904 , RIde82100_224, \8808_9107 );
and \U$16785 ( \25606_25905 , RIfcbbb80_7158, \8810_9109 );
and \U$16786 ( \25607_25906 , RIfc8c150_6616, \8812_9111 );
and \U$16787 ( \25608_25907 , RIfcbbfb8_7161, \8814_9113 );
and \U$16788 ( \25609_25908 , RIfc54458_5981, \8816_9115 );
and \U$16789 ( \25610_25909 , RIe16bbe8_2603, \8818_9117 );
and \U$16790 ( \25611_25910 , RIfc8c2b8_6617, \8820_9119 );
and \U$16791 ( \25612_25911 , RIe168240_2562, \8822_9121 );
and \U$16792 ( \25613_25912 , RIe165978_2533, \8824_9123 );
and \U$16793 ( \25614_25913 , RIe162c78_2501, \8826_9125 );
and \U$16794 ( \25615_25914 , RIee37960_5091, \8828_9127 );
and \U$16795 ( \25616_25915 , RIe15ff78_2469, \8830_9129 );
and \U$16796 ( \25617_25916 , RIfcd6b38_7465, \8832_9131 );
and \U$16797 ( \25618_25917 , RIe15d278_2437, \8834_9133 );
and \U$16798 ( \25619_25918 , RIe157878_2373, \8836_9135 );
and \U$16799 ( \25620_25919 , RIe154b78_2341, \8838_9137 );
and \U$16800 ( \25621_25920 , RIfc8e5e0_6642, \8840_9139 );
and \U$16801 ( \25622_25921 , RIe151e78_2309, \8842_9141 );
and \U$16802 ( \25623_25922 , RIfcb4290_7072, \8844_9143 );
and \U$16803 ( \25624_25923 , RIe14f178_2277, \8846_9145 );
and \U$16804 ( \25625_25924 , RIfc56ff0_6012, \8848_9147 );
and \U$16805 ( \25626_25925 , RIe14c478_2245, \8850_9149 );
and \U$16806 ( \25627_25926 , RIe149778_2213, \8852_9151 );
and \U$16807 ( \25628_25927 , RIe146a78_2181, \8854_9153 );
and \U$16808 ( \25629_25928 , RIee346c0_5055, \8856_9155 );
and \U$16809 ( \25630_25929 , RIee335e0_5043, \8858_9157 );
and \U$16810 ( \25631_25930 , RIee32398_5030, \8860_9159 );
and \U$16811 ( \25632_25931 , RIee31420_5019, \8862_9161 );
and \U$16812 ( \25633_25932 , RIe141348_2119, \8864_9163 );
and \U$16813 ( \25634_25933 , RIe13f020_2094, \8866_9165 );
and \U$16814 ( \25635_25934 , RIfec16f8_8321, \8868_9167 );
and \U$16815 ( \25636_25935 , RIdf3a930_2043, \8870_9169 );
and \U$16816 ( \25637_25936 , RIfce3e28_7615, \8872_9171 );
and \U$16817 ( \25638_25937 , RIfc56780_6006, \8874_9173 );
and \U$16818 ( \25639_25938 , RIfcb4128_7071, \8876_9175 );
and \U$16819 ( \25640_25939 , RIfce2eb0_7604, \8878_9177 );
and \U$16820 ( \25641_25940 , RIdf35d40_1989, \8880_9179 );
and \U$16821 ( \25642_25941 , RIfe88218_7893, \8882_9181 );
and \U$16822 ( \25643_25942 , RIdf316f0_1939, \8884_9183 );
and \U$16823 ( \25644_25943 , RIdf2f698_1916, \8886_9185 );
or \U$16824 ( \25645_25944 , \25581_25880 , \25582_25881 , \25583_25882 , \25584_25883 , \25585_25884 , \25586_25885 , \25587_25886 , \25588_25887 , \25589_25888 , \25590_25889 , \25591_25890 , \25592_25891 , \25593_25892 , \25594_25893 , \25595_25894 , \25596_25895 , \25597_25896 , \25598_25897 , \25599_25898 , \25600_25899 , \25601_25900 , \25602_25901 , \25603_25902 , \25604_25903 , \25605_25904 , \25606_25905 , \25607_25906 , \25608_25907 , \25609_25908 , \25610_25909 , \25611_25910 , \25612_25911 , \25613_25912 , \25614_25913 , \25615_25914 , \25616_25915 , \25617_25916 , \25618_25917 , \25619_25918 , \25620_25919 , \25621_25920 , \25622_25921 , \25623_25922 , \25624_25923 , \25625_25924 , \25626_25925 , \25627_25926 , \25628_25927 , \25629_25928 , \25630_25929 , \25631_25930 , \25632_25931 , \25633_25932 , \25634_25933 , \25635_25934 , \25636_25935 , \25637_25936 , \25638_25937 , \25639_25938 , \25640_25939 , \25641_25940 , \25642_25941 , \25643_25942 , \25644_25943 );
and \U$16825 ( \25646_25945 , RIfc7f9a0_6474, \8889_9188 );
and \U$16826 ( \25647_25946 , RIfce4260_7618, \8891_9190 );
and \U$16827 ( \25648_25947 , RIfcd62c8_7459, \8893_9192 );
and \U$16828 ( \25649_25948 , RIfce9990_7680, \8895_9194 );
and \U$16829 ( \25650_25949 , RIdf2a670_1859, \8897_9196 );
and \U$16830 ( \25651_25950 , RIdf284b0_1835, \8899_9198 );
and \U$16831 ( \25652_25951 , RIdf26728_1814, \8901_9200 );
and \U$16832 ( \25653_25952 , RIdf24c70_1795, \8903_9202 );
and \U$16833 ( \25654_25953 , RIfc7ecf8_6465, \8905_9204 );
and \U$16834 ( \25655_25954 , RIfcc31a0_7242, \8907_9206 );
and \U$16835 ( \25656_25955 , RIfc99008_6763, \8909_9208 );
and \U$16836 ( \25657_25956 , RIfc46e98_5829, \8911_9210 );
and \U$16837 ( \25658_25957 , RIfce2a78_7601, \8913_9212 );
and \U$16838 ( \25659_25958 , RIdf1fdb0_1739, \8915_9214 );
and \U$16839 ( \25660_25959 , RIfcc6e18_7285, \8917_9216 );
and \U$16840 ( \25661_25960 , RIdf19708_1666, \8919_9218 );
and \U$16841 ( \25662_25961 , RIdf17548_1642, \8921_9220 );
and \U$16842 ( \25663_25962 , RIdf14848_1610, \8923_9222 );
and \U$16843 ( \25664_25963 , RIdf11b48_1578, \8925_9224 );
and \U$16844 ( \25665_25964 , RIdf0ee48_1546, \8927_9226 );
and \U$16845 ( \25666_25965 , RIdf0c148_1514, \8929_9228 );
and \U$16846 ( \25667_25966 , RIdf09448_1482, \8931_9230 );
and \U$16847 ( \25668_25967 , RIdf06748_1450, \8933_9232 );
and \U$16848 ( \25669_25968 , RIdf03a48_1418, \8935_9234 );
and \U$16849 ( \25670_25969 , RIdefe048_1354, \8937_9236 );
and \U$16850 ( \25671_25970 , RIdefb348_1322, \8939_9238 );
and \U$16851 ( \25672_25971 , RIdef8648_1290, \8941_9240 );
and \U$16852 ( \25673_25972 , RIdef5948_1258, \8943_9242 );
and \U$16853 ( \25674_25973 , RIdef2c48_1226, \8945_9244 );
and \U$16854 ( \25675_25974 , RIdeeff48_1194, \8947_9246 );
and \U$16855 ( \25676_25975 , RIdeed248_1162, \8949_9248 );
and \U$16856 ( \25677_25976 , RIdeea548_1130, \8951_9250 );
and \U$16857 ( \25678_25977 , RIfcd9130_7492, \8953_9252 );
and \U$16858 ( \25679_25978 , RIfc7cb38_6441, \8955_9254 );
and \U$16859 ( \25680_25979 , RIfc97af0_6748, \8957_9256 );
and \U$16860 ( \25681_25980 , RIfcb3e58_7069, \8959_9258 );
and \U$16861 ( \25682_25981 , RIdee4e18_1068, \8961_9260 );
and \U$16862 ( \25683_25982 , RIdee3090_1047, \8963_9262 );
and \U$16863 ( \25684_25983 , RIdee0ed0_1023, \8965_9264 );
and \U$16864 ( \25685_25984 , RIfe88380_7894, \8967_9266 );
and \U$16865 ( \25686_25985 , RIfc97dc0_6750, \8969_9268 );
and \U$16866 ( \25687_25986 , RIfcc2930_7236, \8971_9270 );
and \U$16867 ( \25688_25987 , RIfcd9298_7493, \8973_9272 );
and \U$16868 ( \25689_25988 , RIfc7c868_6439, \8975_9274 );
and \U$16869 ( \25690_25989 , RIded9ce8_942, \8977_9276 );
and \U$16870 ( \25691_25990 , RIded76f0_915, \8979_9278 );
and \U$16871 ( \25692_25991 , RIded5968_894, \8981_9280 );
and \U$16872 ( \25693_25992 , RIded3370_867, \8983_9282 );
and \U$16873 ( \25694_25993 , RIded0d78_840, \8985_9284 );
and \U$16874 ( \25695_25994 , RIdece078_808, \8987_9286 );
and \U$16875 ( \25696_25995 , RIdecb378_776, \8989_9288 );
and \U$16876 ( \25697_25996 , RIdec8678_744, \8991_9290 );
and \U$16877 ( \25698_25997 , RIdeb4b78_520, \8993_9292 );
and \U$16878 ( \25699_25998 , RIde97640_328, \8995_9294 );
and \U$16879 ( \25700_25999 , RIe16e780_2634, \8997_9296 );
and \U$16880 ( \25701_26000 , RIe15a578_2405, \8999_9298 );
and \U$16881 ( \25702_26001 , RIe143d78_2149, \9001_9300 );
and \U$16882 ( \25703_26002 , RIdf38770_2019, \9003_9302 );
and \U$16883 ( \25704_26003 , RIdf2cdd0_1887, \9005_9304 );
and \U$16884 ( \25705_26004 , RIdf1d650_1711, \9007_9306 );
and \U$16885 ( \25706_26005 , RIdf00d48_1386, \9009_9308 );
and \U$16886 ( \25707_26006 , RIdee7848_1098, \9011_9310 );
and \U$16887 ( \25708_26007 , RIdedc5b0_971, \9013_9312 );
and \U$16888 ( \25709_26008 , RIde7d588_201, \9015_9314 );
or \U$16889 ( \25710_26009 , \25646_25945 , \25647_25946 , \25648_25947 , \25649_25948 , \25650_25949 , \25651_25950 , \25652_25951 , \25653_25952 , \25654_25953 , \25655_25954 , \25656_25955 , \25657_25956 , \25658_25957 , \25659_25958 , \25660_25959 , \25661_25960 , \25662_25961 , \25663_25962 , \25664_25963 , \25665_25964 , \25666_25965 , \25667_25966 , \25668_25967 , \25669_25968 , \25670_25969 , \25671_25970 , \25672_25971 , \25673_25972 , \25674_25973 , \25675_25974 , \25676_25975 , \25677_25976 , \25678_25977 , \25679_25978 , \25680_25979 , \25681_25980 , \25682_25981 , \25683_25982 , \25684_25983 , \25685_25984 , \25686_25985 , \25687_25986 , \25688_25987 , \25689_25988 , \25690_25989 , \25691_25990 , \25692_25991 , \25693_25992 , \25694_25993 , \25695_25994 , \25696_25995 , \25697_25996 , \25698_25997 , \25699_25998 , \25700_25999 , \25701_26000 , \25702_26001 , \25703_26002 , \25704_26003 , \25705_26004 , \25706_26005 , \25707_26006 , \25708_26007 , \25709_26008 );
or \U$16890 ( \25711_26010 , \25645_25944 , \25710_26009 );
_DC \g2553/U$1 ( \25712 , \25711_26010 , \9024_9323 );
buf \U$16891 ( \25713_26012 , \25712 );
and \U$16892 ( \25714_26013 , RIe19dc10_3172, \9034_9333 );
and \U$16893 ( \25715_26014 , RIe19af10_3140, \9036_9335 );
and \U$16894 ( \25716_26015 , RIfec1590_8320, \9038_9337 );
and \U$16895 ( \25717_26016 , RIe198210_3108, \9040_9339 );
and \U$16896 ( \25718_26017 , RIfec1428_8319, \9042_9341 );
and \U$16897 ( \25719_26018 , RIe195510_3076, \9044_9343 );
and \U$16898 ( \25720_26019 , RIe192810_3044, \9046_9345 );
and \U$16899 ( \25721_26020 , RIe18fb10_3012, \9048_9347 );
and \U$16900 ( \25722_26021 , RIe18a110_2948, \9050_9349 );
and \U$16901 ( \25723_26022 , RIe187410_2916, \9052_9351 );
and \U$16902 ( \25724_26023 , RIfec12c0_8318, \9054_9353 );
and \U$16903 ( \25725_26024 , RIe184710_2884, \9056_9355 );
and \U$16904 ( \25726_26025 , RIfc88370_6572, \9058_9357 );
and \U$16905 ( \25727_26026 , RIe181a10_2852, \9060_9359 );
and \U$16906 ( \25728_26027 , RIe17ed10_2820, \9062_9361 );
and \U$16907 ( \25729_26028 , RIe17c010_2788, \9064_9363 );
and \U$16908 ( \25730_26029 , RIfc6ccb0_6260, \9066_9365 );
and \U$16909 ( \25731_26030 , RIfc5f858_6109, \9068_9367 );
and \U$16910 ( \25732_26031 , RIfca88f0_6940, \9070_9369 );
and \U$16911 ( \25733_26032 , RIe175f08_2719, \9072_9371 );
and \U$16912 ( \25734_26033 , RIfc81020_6490, \9074_9373 );
and \U$16913 ( \25735_26034 , RIfcc6008_7275, \9076_9375 );
and \U$16914 ( \25736_26035 , RIfc4ea58_5917, \9078_9377 );
and \U$16915 ( \25737_26036 , RIfc42140_5774, \9080_9379 );
and \U$16916 ( \25738_26037 , RIfca3b98_6885, \9082_9381 );
and \U$16917 ( \25739_26038 , RIfc5ac68_6055, \9084_9383 );
and \U$16918 ( \25740_26039 , RIfc984c8_6755, \9086_9385 );
and \U$16919 ( \25741_26040 , RIe173d48_2695, \9088_9387 );
and \U$16920 ( \25742_26041 , RIfc9b330_6788, \9090_9389 );
and \U$16921 ( \25743_26042 , RIf16f688_5727, \9092_9391 );
and \U$16922 ( \25744_26043 , RIfc42410_5776, \9094_9393 );
and \U$16923 ( \25745_26044 , RIfc5f588_6107, \9096_9395 );
and \U$16924 ( \25746_26045 , RIfe880b0_7892, \9098_9397 );
and \U$16925 ( \25747_26046 , RIe223f68_4699, \9100_9399 );
and \U$16926 ( \25748_26047 , RIf16bfb0_5688, \9102_9401 );
and \U$16927 ( \25749_26048 , RIe221268_4667, \9104_9403 );
and \U$16928 ( \25750_26049 , RIfc86cf0_6556, \9106_9405 );
and \U$16929 ( \25751_26050 , RIe21e568_4635, \9108_9407 );
and \U$16930 ( \25752_26051 , RIe218b68_4571, \9110_9409 );
and \U$16931 ( \25753_26052 , RIe215e68_4539, \9112_9411 );
and \U$16932 ( \25754_26053 , RIfe87de0_7890, \9114_9413 );
and \U$16933 ( \25755_26054 , RIe213168_4507, \9116_9415 );
and \U$16934 ( \25756_26055 , RIf1692b0_5656, \9118_9417 );
and \U$16935 ( \25757_26056 , RIe210468_4475, \9120_9419 );
and \U$16936 ( \25758_26057 , RIfcdf670_7564, \9122_9421 );
and \U$16937 ( \25759_26058 , RIe20d768_4443, \9124_9423 );
and \U$16938 ( \25760_26059 , RIe20aa68_4411, \9126_9425 );
and \U$16939 ( \25761_26060 , RIe207d68_4379, \9128_9427 );
and \U$16940 ( \25762_26061 , RIfca6460_6914, \9130_9429 );
and \U$16941 ( \25763_26062 , RIf1662e0_5622, \9132_9431 );
and \U$16942 ( \25764_26063 , RIe202908_4319, \9134_9433 );
and \U$16943 ( \25765_26064 , RIfe87b10_7888, \9136_9435 );
and \U$16944 ( \25766_26065 , RIfc58c10_6032, \9138_9437 );
and \U$16945 ( \25767_26066 , RIfc50ab0_5940, \9140_9439 );
and \U$16946 ( \25768_26067 , RIfccd790_7360, \9142_9441 );
and \U$16947 ( \25769_26068 , RIfccd1f0_7356, \9144_9443 );
and \U$16948 ( \25770_26069 , RIf160610_5556, \9146_9445 );
and \U$16949 ( \25771_26070 , RIf15e720_5534, \9148_9447 );
and \U$16950 ( \25772_26071 , RIfe87c78_7889, \9150_9449 );
and \U$16951 ( \25773_26072 , RIfe87f48_7891, \9152_9451 );
and \U$16952 ( \25774_26073 , RIfce7668_7655, \9154_9453 );
and \U$16953 ( \25775_26074 , RIfc86480_6550, \9156_9455 );
and \U$16954 ( \25776_26075 , RIfcd2218_7413, \9158_9457 );
and \U$16955 ( \25777_26076 , RIfcb01e0_7026, \9160_9459 );
or \U$16956 ( \25778_26077 , \25714_26013 , \25715_26014 , \25716_26015 , \25717_26016 , \25718_26017 , \25719_26018 , \25720_26019 , \25721_26020 , \25722_26021 , \25723_26022 , \25724_26023 , \25725_26024 , \25726_26025 , \25727_26026 , \25728_26027 , \25729_26028 , \25730_26029 , \25731_26030 , \25732_26031 , \25733_26032 , \25734_26033 , \25735_26034 , \25736_26035 , \25737_26036 , \25738_26037 , \25739_26038 , \25740_26039 , \25741_26040 , \25742_26041 , \25743_26042 , \25744_26043 , \25745_26044 , \25746_26045 , \25747_26046 , \25748_26047 , \25749_26048 , \25750_26049 , \25751_26050 , \25752_26051 , \25753_26052 , \25754_26053 , \25755_26054 , \25756_26055 , \25757_26056 , \25758_26057 , \25759_26058 , \25760_26059 , \25761_26060 , \25762_26061 , \25763_26062 , \25764_26063 , \25765_26064 , \25766_26065 , \25767_26066 , \25768_26067 , \25769_26068 , \25770_26069 , \25771_26070 , \25772_26071 , \25773_26072 , \25774_26073 , \25775_26074 , \25776_26075 , \25777_26076 );
and \U$16957 ( \25779_26078 , RIfc47b40_5838, \9163_9462 );
and \U$16958 ( \25780_26079 , RIfc84158_6525, \9165_9464 );
and \U$16959 ( \25781_26080 , RIfc4b920_5882, \9167_9466 );
and \U$16960 ( \25782_26081 , RIe1fa4d8_4225, \9169_9468 );
and \U$16961 ( \25783_26082 , RIfc4ba88_5883, \9171_9470 );
and \U$16962 ( \25784_26083 , RIfcb7530_7108, \9173_9472 );
and \U$16963 ( \25785_26084 , RIfcd58f0_7452, \9175_9474 );
and \U$16964 ( \25786_26085 , RIe1f5a50_4172, \9177_9476 );
and \U$16965 ( \25787_26086 , RIf153488_5407, \9179_9478 );
and \U$16966 ( \25788_26087 , RIf151ca0_5390, \9181_9480 );
and \U$16967 ( \25789_26088 , RIfc51e60_5954, \9183_9482 );
and \U$16968 ( \25790_26089 , RIe1f3728_4147, \9185_9484 );
and \U$16969 ( \25791_26090 , RIfc9aef8_6785, \9187_9486 );
and \U$16970 ( \25792_26091 , RIfcbaaa0_7146, \9189_9488 );
and \U$16971 ( \25793_26092 , RIfc52130_5956, \9191_9490 );
and \U$16972 ( \25794_26093 , RIe1ee430_4088, \9193_9492 );
and \U$16973 ( \25795_26094 , RIe1ebcd0_4060, \9195_9494 );
and \U$16974 ( \25796_26095 , RIe1e8fd0_4028, \9197_9496 );
and \U$16975 ( \25797_26096 , RIe1e62d0_3996, \9199_9498 );
and \U$16976 ( \25798_26097 , RIe1e35d0_3964, \9201_9500 );
and \U$16977 ( \25799_26098 , RIe1e08d0_3932, \9203_9502 );
and \U$16978 ( \25800_26099 , RIe1ddbd0_3900, \9205_9504 );
and \U$16979 ( \25801_26100 , RIe1daed0_3868, \9207_9506 );
and \U$16980 ( \25802_26101 , RIe1d81d0_3836, \9209_9508 );
and \U$16981 ( \25803_26102 , RIe1d27d0_3772, \9211_9510 );
and \U$16982 ( \25804_26103 , RIe1cfad0_3740, \9213_9512 );
and \U$16983 ( \25805_26104 , RIe1ccdd0_3708, \9215_9514 );
and \U$16984 ( \25806_26105 , RIe1ca0d0_3676, \9217_9516 );
and \U$16985 ( \25807_26106 , RIe1c73d0_3644, \9219_9518 );
and \U$16986 ( \25808_26107 , RIe1c46d0_3612, \9221_9520 );
and \U$16987 ( \25809_26108 , RIe1c19d0_3580, \9223_9522 );
and \U$16988 ( \25810_26109 , RIe1becd0_3548, \9225_9524 );
and \U$16989 ( \25811_26110 , RIfce0b88_7579, \9227_9526 );
and \U$16990 ( \25812_26111 , RIfc82808_6507, \9229_9528 );
and \U$16991 ( \25813_26112 , RIe1b9708_3487, \9231_9530 );
and \U$16992 ( \25814_26113 , RIe1b76b0_3464, \9233_9532 );
and \U$16993 ( \25815_26114 , RIfcd5bc0_7454, \9235_9534 );
and \U$16994 ( \25816_26115 , RIfcb69f0_7100, \9237_9536 );
and \U$16995 ( \25817_26116 , RIe1b54f0_3440, \9239_9538 );
and \U$16996 ( \25818_26117 , RIe1b4140_3426, \9241_9540 );
and \U$16997 ( \25819_26118 , RIfc89f90_6592, \9243_9542 );
and \U$16998 ( \25820_26119 , RIfce9af8_7681, \9245_9544 );
and \U$16999 ( \25821_26120 , RIe1b2958_3409, \9247_9546 );
and \U$17000 ( \25822_26121 , RIe1b0ea0_3390, \9249_9548 );
and \U$17001 ( \25823_26122 , RIfc4a138_5865, \9251_9550 );
and \U$17002 ( \25824_26123 , RIfc8a260_6594, \9253_9552 );
and \U$17003 ( \25825_26124 , RIe1ac850_3340, \9255_9554 );
and \U$17004 ( \25826_26125 , RIe1ab1d0_3324, \9257_9556 );
and \U$17005 ( \25827_26126 , RIe1a9010_3300, \9259_9558 );
and \U$17006 ( \25828_26127 , RIe1a6310_3268, \9261_9560 );
and \U$17007 ( \25829_26128 , RIe1a3610_3236, \9263_9562 );
and \U$17008 ( \25830_26129 , RIe1a0910_3204, \9265_9564 );
and \U$17009 ( \25831_26130 , RIe18ce10_2980, \9267_9566 );
and \U$17010 ( \25832_26131 , RIe179310_2756, \9269_9568 );
and \U$17011 ( \25833_26132 , RIe226c68_4731, \9271_9570 );
and \U$17012 ( \25834_26133 , RIe21b868_4603, \9273_9572 );
and \U$17013 ( \25835_26134 , RIe205068_4347, \9275_9574 );
and \U$17014 ( \25836_26135 , RIe1ff0c8_4279, \9277_9576 );
and \U$17015 ( \25837_26136 , RIe1f8480_4202, \9279_9578 );
and \U$17016 ( \25838_26137 , RIe1f0fc8_4119, \9281_9580 );
and \U$17017 ( \25839_26138 , RIe1d54d0_3804, \9283_9582 );
and \U$17018 ( \25840_26139 , RIe1bbfd0_3516, \9285_9584 );
and \U$17019 ( \25841_26140 , RIe1aee48_3367, \9287_9586 );
and \U$17020 ( \25842_26141 , RIe171480_2666, \9289_9588 );
or \U$17021 ( \25843_26142 , \25779_26078 , \25780_26079 , \25781_26080 , \25782_26081 , \25783_26082 , \25784_26083 , \25785_26084 , \25786_26085 , \25787_26086 , \25788_26087 , \25789_26088 , \25790_26089 , \25791_26090 , \25792_26091 , \25793_26092 , \25794_26093 , \25795_26094 , \25796_26095 , \25797_26096 , \25798_26097 , \25799_26098 , \25800_26099 , \25801_26100 , \25802_26101 , \25803_26102 , \25804_26103 , \25805_26104 , \25806_26105 , \25807_26106 , \25808_26107 , \25809_26108 , \25810_26109 , \25811_26110 , \25812_26111 , \25813_26112 , \25814_26113 , \25815_26114 , \25816_26115 , \25817_26116 , \25818_26117 , \25819_26118 , \25820_26119 , \25821_26120 , \25822_26121 , \25823_26122 , \25824_26123 , \25825_26124 , \25826_26125 , \25827_26126 , \25828_26127 , \25829_26128 , \25830_26129 , \25831_26130 , \25832_26131 , \25833_26132 , \25834_26133 , \25835_26134 , \25836_26135 , \25837_26136 , \25838_26137 , \25839_26138 , \25840_26139 , \25841_26140 , \25842_26141 );
or \U$17022 ( \25844_26143 , \25778_26077 , \25843_26142 );
_DC \g3680/U$1 ( \25845 , \25844_26143 , \9298_9597 );
buf \U$17023 ( \25846_26145 , \25845 );
xor \U$17024 ( \25847_26146 , \25713_26012 , \25846_26145 );
and \U$17025 ( \25848_26147 , RIdec5810_711, \8760_9059 );
and \U$17026 ( \25849_26148 , RIdec2b10_679, \8762_9061 );
and \U$17027 ( \25850_26149 , RIfce6f60_7650, \8764_9063 );
and \U$17028 ( \25851_26150 , RIdebfe10_647, \8766_9065 );
and \U$17029 ( \25852_26151 , RIfc95228_6719, \8768_9067 );
and \U$17030 ( \25853_26152 , RIdebd110_615, \8770_9069 );
and \U$17031 ( \25854_26153 , RIdeba410_583, \8772_9071 );
and \U$17032 ( \25855_26154 , RIdeb7710_551, \8774_9073 );
and \U$17033 ( \25856_26155 , RIfe879a8_7887, \8776_9075 );
and \U$17034 ( \25857_26156 , RIdeb1d10_487, \8778_9077 );
and \U$17035 ( \25858_26157 , RIfcc16e8_7223, \8780_9079 );
and \U$17036 ( \25859_26158 , RIdeaf010_455, \8782_9081 );
and \U$17037 ( \25860_26159 , RIfca4f48_6899, \8784_9083 );
and \U$17038 ( \25861_26160 , RIdeaadf8_423, \8786_9085 );
and \U$17039 ( \25862_26161 , RIdea44f8_391, \8788_9087 );
and \U$17040 ( \25863_26162 , RIde9dbf8_359, \8790_9089 );
and \U$17041 ( \25864_26163 , RIee1cf48_4788, \8792_9091 );
and \U$17042 ( \25865_26164 , RIee1bfd0_4777, \8794_9093 );
and \U$17043 ( \25866_26165 , RIfc95660_6722, \8796_9095 );
and \U$17044 ( \25867_26166 , RIfcee148_7731, \8798_9097 );
and \U$17045 ( \25868_26167 , RIfe87840_7886, \8800_9099 );
and \U$17046 ( \25869_26168 , RIfe876d8_7885, \8802_9101 );
and \U$17047 ( \25870_26169 , RIde8a0f8_263, \8804_9103 );
and \U$17048 ( \25871_26170 , RIde85f58_243, \8806_9105 );
and \U$17049 ( \25872_26171 , RIfcb0780_7030, \8808_9107 );
and \U$17050 ( \25873_26172 , RIfcee9b8_7737, \8810_9109 );
and \U$17051 ( \25874_26173 , RIfc5f150_6104, \8812_9111 );
and \U$17052 ( \25875_26174 , RIfcdee00_7558, \8814_9113 );
and \U$17053 ( \25876_26175 , RIfcd8050_7480, \8816_9115 );
and \U$17054 ( \25877_26176 , RIe16ba80_2602, \8818_9117 );
and \U$17055 ( \25878_26177 , RIfca5380_6902, \8820_9119 );
and \U$17056 ( \25879_26178 , RIe1680d8_2561, \8822_9121 );
and \U$17057 ( \25880_26179 , RIe165810_2532, \8824_9123 );
and \U$17058 ( \25881_26180 , RIe162b10_2500, \8826_9125 );
and \U$17059 ( \25882_26181 , RIee377f8_5090, \8828_9127 );
and \U$17060 ( \25883_26182 , RIe15fe10_2468, \8830_9129 );
and \U$17061 ( \25884_26183 , RIee36448_5076, \8832_9131 );
and \U$17062 ( \25885_26184 , RIe15d110_2436, \8834_9133 );
and \U$17063 ( \25886_26185 , RIe157710_2372, \8836_9135 );
and \U$17064 ( \25887_26186 , RIe154a10_2340, \8838_9137 );
and \U$17065 ( \25888_26187 , RIfc3f3c8_5745, \8840_9139 );
and \U$17066 ( \25889_26188 , RIe151d10_2308, \8842_9141 );
and \U$17067 ( \25890_26189 , RIfcde9c8_7555, \8844_9143 );
and \U$17068 ( \25891_26190 , RIe14f010_2276, \8846_9145 );
and \U$17069 ( \25892_26191 , RIfc4a2a0_5866, \8848_9147 );
and \U$17070 ( \25893_26192 , RIe14c310_2244, \8850_9149 );
and \U$17071 ( \25894_26193 , RIe149610_2212, \8852_9151 );
and \U$17072 ( \25895_26194 , RIe146910_2180, \8854_9153 );
and \U$17073 ( \25896_26195 , RIfc62288_6139, \8856_9155 );
and \U$17074 ( \25897_26196 , RIee33478_5042, \8858_9157 );
and \U$17075 ( \25898_26197 , RIfc71b70_6316, \8860_9159 );
and \U$17076 ( \25899_26198 , RIee312b8_5018, \8862_9161 );
and \U$17077 ( \25900_26199 , RIe1411e0_2118, \8864_9163 );
and \U$17078 ( \25901_26200 , RIfe87570_7884, \8866_9165 );
and \U$17079 ( \25902_26201 , RIdf3cf28_2070, \8868_9167 );
and \U$17080 ( \25903_26202 , RIfe87408_7883, \8870_9169 );
and \U$17081 ( \25904_26203 , RIfcc99b0_7316, \8872_9171 );
and \U$17082 ( \25905_26204 , RIfccf0e0_7378, \8874_9173 );
and \U$17083 ( \25906_26205 , RIfcaeb60_7010, \8876_9175 );
and \U$17084 ( \25907_26206 , RIfcca220_7322, \8878_9177 );
and \U$17085 ( \25908_26207 , RIdf35bd8_1988, \8880_9179 );
and \U$17086 ( \25909_26208 , RIdf33748_1962, \8882_9181 );
and \U$17087 ( \25910_26209 , RIdf31588_1938, \8884_9183 );
and \U$17088 ( \25911_26210 , RIdf2f530_1915, \8886_9185 );
or \U$17089 ( \25912_26211 , \25848_26147 , \25849_26148 , \25850_26149 , \25851_26150 , \25852_26151 , \25853_26152 , \25854_26153 , \25855_26154 , \25856_26155 , \25857_26156 , \25858_26157 , \25859_26158 , \25860_26159 , \25861_26160 , \25862_26161 , \25863_26162 , \25864_26163 , \25865_26164 , \25866_26165 , \25867_26166 , \25868_26167 , \25869_26168 , \25870_26169 , \25871_26170 , \25872_26171 , \25873_26172 , \25874_26173 , \25875_26174 , \25876_26175 , \25877_26176 , \25878_26177 , \25879_26178 , \25880_26179 , \25881_26180 , \25882_26181 , \25883_26182 , \25884_26183 , \25885_26184 , \25886_26185 , \25887_26186 , \25888_26187 , \25889_26188 , \25890_26189 , \25891_26190 , \25892_26191 , \25893_26192 , \25894_26193 , \25895_26194 , \25896_26195 , \25897_26196 , \25898_26197 , \25899_26198 , \25900_26199 , \25901_26200 , \25902_26201 , \25903_26202 , \25904_26203 , \25905_26204 , \25906_26205 , \25907_26206 , \25908_26207 , \25909_26208 , \25910_26209 , \25911_26210 );
and \U$17090 ( \25913_26212 , RIee2be58_4958, \8889_9188 );
and \U$17091 ( \25914_26213 , RIee2a508_4940, \8891_9190 );
and \U$17092 ( \25915_26214 , RIee28ff0_4925, \8893_9192 );
and \U$17093 ( \25916_26215 , RIee27da8_4912, \8895_9194 );
and \U$17094 ( \25917_26216 , RIdf2a508_1858, \8897_9196 );
and \U$17095 ( \25918_26217 , RIdf28348_1834, \8899_9198 );
and \U$17096 ( \25919_26218 , RIdf265c0_1813, \8901_9200 );
and \U$17097 ( \25920_26219 , RIdf24b08_1794, \8903_9202 );
and \U$17098 ( \25921_26220 , RIfc74708_6347, \8905_9204 );
and \U$17099 ( \25922_26221 , RIfc42578_5777, \8907_9206 );
and \U$17100 ( \25923_26222 , RIfc43388_5787, \8909_9208 );
and \U$17101 ( \25924_26223 , RIfc745a0_6346, \8911_9210 );
and \U$17102 ( \25925_26224 , RIfcb0078_7025, \8913_9212 );
and \U$17103 ( \25926_26225 , RIdf1fc48_1738, \8915_9214 );
and \U$17104 ( \25927_26226 , RIfcaff10_7024, \8917_9216 );
and \U$17105 ( \25928_26227 , RIdf195a0_1665, \8919_9218 );
and \U$17106 ( \25929_26228 , RIdf173e0_1641, \8921_9220 );
and \U$17107 ( \25930_26229 , RIdf146e0_1609, \8923_9222 );
and \U$17108 ( \25931_26230 , RIdf119e0_1577, \8925_9224 );
and \U$17109 ( \25932_26231 , RIdf0ece0_1545, \8927_9226 );
and \U$17110 ( \25933_26232 , RIdf0bfe0_1513, \8929_9228 );
and \U$17111 ( \25934_26233 , RIdf092e0_1481, \8931_9230 );
and \U$17112 ( \25935_26234 , RIdf065e0_1449, \8933_9232 );
and \U$17113 ( \25936_26235 , RIdf038e0_1417, \8935_9234 );
and \U$17114 ( \25937_26236 , RIdefdee0_1353, \8937_9236 );
and \U$17115 ( \25938_26237 , RIdefb1e0_1321, \8939_9238 );
and \U$17116 ( \25939_26238 , RIdef84e0_1289, \8941_9240 );
and \U$17117 ( \25940_26239 , RIdef57e0_1257, \8943_9242 );
and \U$17118 ( \25941_26240 , RIdef2ae0_1225, \8945_9244 );
and \U$17119 ( \25942_26241 , RIdeefde0_1193, \8947_9246 );
and \U$17120 ( \25943_26242 , RIdeed0e0_1161, \8949_9248 );
and \U$17121 ( \25944_26243 , RIdeea3e0_1129, \8951_9250 );
and \U$17122 ( \25945_26244 , RIee257b0_4885, \8953_9252 );
and \U$17123 ( \25946_26245 , RIfca73d8_6925, \8955_9254 );
and \U$17124 ( \25947_26246 , RIee23e60_4867, \8957_9256 );
and \U$17125 ( \25948_26247 , RIfce66f0_7644, \8959_9258 );
and \U$17126 ( \25949_26248 , RIdee4cb0_1067, \8961_9260 );
and \U$17127 ( \25950_26249 , RIdee2f28_1046, \8963_9262 );
and \U$17128 ( \25951_26250 , RIdee0d68_1022, \8965_9264 );
and \U$17129 ( \25952_26251 , RIdeded10_999, \8967_9266 );
and \U$17130 ( \25953_26252 , RIfcca388_7323, \8969_9268 );
and \U$17131 ( \25954_26253 , RIfce6858_7645, \8971_9270 );
and \U$17132 ( \25955_26254 , RIfcceca8_7375, \8973_9272 );
and \U$17133 ( \25956_26255 , RIfcdc970_7532, \8975_9274 );
and \U$17134 ( \25957_26256 , RIded9b80_941, \8977_9276 );
and \U$17135 ( \25958_26257 , RIfeaaac0_8258, \8979_9278 );
and \U$17136 ( \25959_26258 , RIded5800_893, \8981_9280 );
and \U$17137 ( \25960_26259 , RIded3208_866, \8983_9282 );
and \U$17138 ( \25961_26260 , RIded0c10_839, \8985_9284 );
and \U$17139 ( \25962_26261 , RIdecdf10_807, \8987_9286 );
and \U$17140 ( \25963_26262 , RIdecb210_775, \8989_9288 );
and \U$17141 ( \25964_26263 , RIdec8510_743, \8991_9290 );
and \U$17142 ( \25965_26264 , RIdeb4a10_519, \8993_9292 );
and \U$17143 ( \25966_26265 , RIde972f8_327, \8995_9294 );
and \U$17144 ( \25967_26266 , RIe16e618_2633, \8997_9296 );
and \U$17145 ( \25968_26267 , RIe15a410_2404, \8999_9298 );
and \U$17146 ( \25969_26268 , RIe143c10_2148, \9001_9300 );
and \U$17147 ( \25970_26269 , RIdf38608_2018, \9003_9302 );
and \U$17148 ( \25971_26270 , RIdf2cc68_1886, \9005_9304 );
and \U$17149 ( \25972_26271 , RIdf1d4e8_1710, \9007_9306 );
and \U$17150 ( \25973_26272 , RIdf00be0_1385, \9009_9308 );
and \U$17151 ( \25974_26273 , RIdee76e0_1097, \9011_9310 );
and \U$17152 ( \25975_26274 , RIdedc448_970, \9013_9312 );
and \U$17153 ( \25976_26275 , RIde7d240_200, \9015_9314 );
or \U$17154 ( \25977_26276 , \25913_26212 , \25914_26213 , \25915_26214 , \25916_26215 , \25917_26216 , \25918_26217 , \25919_26218 , \25920_26219 , \25921_26220 , \25922_26221 , \25923_26222 , \25924_26223 , \25925_26224 , \25926_26225 , \25927_26226 , \25928_26227 , \25929_26228 , \25930_26229 , \25931_26230 , \25932_26231 , \25933_26232 , \25934_26233 , \25935_26234 , \25936_26235 , \25937_26236 , \25938_26237 , \25939_26238 , \25940_26239 , \25941_26240 , \25942_26241 , \25943_26242 , \25944_26243 , \25945_26244 , \25946_26245 , \25947_26246 , \25948_26247 , \25949_26248 , \25950_26249 , \25951_26250 , \25952_26251 , \25953_26252 , \25954_26253 , \25955_26254 , \25956_26255 , \25957_26256 , \25958_26257 , \25959_26258 , \25960_26259 , \25961_26260 , \25962_26261 , \25963_26262 , \25964_26263 , \25965_26264 , \25966_26265 , \25967_26266 , \25968_26267 , \25969_26268 , \25970_26269 , \25971_26270 , \25972_26271 , \25973_26272 , \25974_26273 , \25975_26274 , \25976_26275 );
or \U$17155 ( \25978_26277 , \25912_26211 , \25977_26276 );
_DC \g25d8/U$1 ( \25979 , \25978_26277 , \9024_9323 );
buf \U$17156 ( \25980_26279 , \25979 );
and \U$17157 ( \25981_26280 , RIe19daa8_3171, \9034_9333 );
and \U$17158 ( \25982_26281 , RIe19ada8_3139, \9036_9335 );
and \U$17159 ( \25983_26282 , RIf1457c0_5250, \9038_9337 );
and \U$17160 ( \25984_26283 , RIe1980a8_3107, \9040_9339 );
and \U$17161 ( \25985_26284 , RIf1449b0_5240, \9042_9341 );
and \U$17162 ( \25986_26285 , RIe1953a8_3075, \9044_9343 );
and \U$17163 ( \25987_26286 , RIe1926a8_3043, \9046_9345 );
and \U$17164 ( \25988_26287 , RIe18f9a8_3011, \9048_9347 );
and \U$17165 ( \25989_26288 , RIe189fa8_2947, \9050_9349 );
and \U$17166 ( \25990_26289 , RIe1872a8_2915, \9052_9351 );
and \U$17167 ( \25991_26290 , RIf143ba0_5230, \9054_9353 );
and \U$17168 ( \25992_26291 , RIe1845a8_2883, \9056_9355 );
and \U$17169 ( \25993_26292 , RIfc912e0_6674, \9058_9357 );
and \U$17170 ( \25994_26293 , RIe1818a8_2851, \9060_9359 );
and \U$17171 ( \25995_26294 , RIe17eba8_2819, \9062_9361 );
and \U$17172 ( \25996_26295 , RIe17bea8_2787, \9064_9363 );
and \U$17173 ( \25997_26296 , RIfc915b0_6676, \9066_9365 );
and \U$17174 ( \25998_26297 , RIfcbe5b0_7188, \9068_9367 );
and \U$17175 ( \25999_26298 , RIfce3b58_7613, \9070_9369 );
and \U$17176 ( \26000_26299 , RIe175da0_2718, \9072_9371 );
and \U$17177 ( \26001_26300 , RIfceb448_7699, \9074_9373 );
and \U$17178 ( \26002_26301 , RIfcc7958_7293, \9076_9375 );
and \U$17179 ( \26003_26302 , RIfc42de8_5783, \9078_9377 );
and \U$17180 ( \26004_26303 , RIfc96e48_6739, \9080_9379 );
and \U$17181 ( \26005_26304 , RIfc7a810_6416, \9082_9381 );
and \U$17182 ( \26006_26305 , RIfc96ce0_6738, \9084_9383 );
and \U$17183 ( \26007_26306 , RIfcc7ac0_7294, \9086_9385 );
and \U$17184 ( \26008_26307 , RIe173be0_2694, \9088_9387 );
and \U$17185 ( \26009_26308 , RIfce39f0_7612, \9090_9389 );
and \U$17186 ( \26010_26309 , RIfc7a540_6414, \9092_9391 );
and \U$17187 ( \26011_26310 , RIfc91b50_6680, \9094_9393 );
and \U$17188 ( \26012_26311 , RIfc429b0_5780, \9096_9395 );
and \U$17189 ( \26013_26312 , RIfea9710_8244, \9098_9397 );
and \U$17190 ( \26014_26313 , RIe223e00_4698, \9100_9399 );
and \U$17191 ( \26015_26314 , RIfcd8488_7483, \9102_9401 );
and \U$17192 ( \26016_26315 , RIe221100_4666, \9104_9403 );
and \U$17193 ( \26017_26316 , RIfc920f0_6684, \9106_9405 );
and \U$17194 ( \26018_26317 , RIe21e400_4634, \9108_9407 );
and \U$17195 ( \26019_26318 , RIe218a00_4570, \9110_9409 );
and \U$17196 ( \26020_26319 , RIe215d00_4538, \9112_9411 );
and \U$17197 ( \26021_26320 , RIfc79e38_6409, \9114_9413 );
and \U$17198 ( \26022_26321 , RIe213000_4506, \9116_9415 );
and \U$17199 ( \26023_26322 , RIfcbee20_7194, \9118_9417 );
and \U$17200 ( \26024_26323 , RIe210300_4474, \9120_9419 );
and \U$17201 ( \26025_26324 , RIf168068_5643, \9122_9421 );
and \U$17202 ( \26026_26325 , RIe20d600_4442, \9124_9423 );
and \U$17203 ( \26027_26326 , RIe20a900_4410, \9126_9425 );
and \U$17204 ( \26028_26327 , RIe207c00_4378, \9128_9427 );
and \U$17205 ( \26029_26328 , RIfc5af38_6057, \9130_9429 );
and \U$17206 ( \26030_26329 , RIfcd73a8_7471, \9132_9431 );
and \U$17207 ( \26031_26330 , RIe2027a0_4318, \9134_9433 );
and \U$17208 ( \26032_26331 , RIe200ce8_4299, \9136_9435 );
and \U$17209 ( \26033_26332 , RIfcb2670_7052, \9138_9437 );
and \U$17210 ( \26034_26333 , RIfcdf940_7566, \9140_9439 );
and \U$17211 ( \26035_26334 , RIfc5b208_6059, \9142_9441 );
and \U$17212 ( \26036_26335 , RIfcbf3c0_7198, \9144_9443 );
and \U$17213 ( \26037_26336 , RIf1604a8_5555, \9146_9445 );
and \U$17214 ( \26038_26337 , RIf15e5b8_5533, \9148_9447 );
and \U$17215 ( \26039_26338 , RIfe872a0_7882, \9150_9449 );
and \U$17216 ( \26040_26339 , RIfe87138_7881, \9152_9451 );
and \U$17217 ( \26041_26340 , RIfc78920_6394, \9154_9453 );
and \U$17218 ( \26042_26341 , RIfec1158_8317, \9156_9455 );
and \U$17219 ( \26043_26342 , RIfc93338_6697, \9158_9457 );
and \U$17220 ( \26044_26343 , RIfcea368_7687, \9160_9459 );
or \U$17221 ( \26045_26344 , \25981_26280 , \25982_26281 , \25983_26282 , \25984_26283 , \25985_26284 , \25986_26285 , \25987_26286 , \25988_26287 , \25989_26288 , \25990_26289 , \25991_26290 , \25992_26291 , \25993_26292 , \25994_26293 , \25995_26294 , \25996_26295 , \25997_26296 , \25998_26297 , \25999_26298 , \26000_26299 , \26001_26300 , \26002_26301 , \26003_26302 , \26004_26303 , \26005_26304 , \26006_26305 , \26007_26306 , \26008_26307 , \26009_26308 , \26010_26309 , \26011_26310 , \26012_26311 , \26013_26312 , \26014_26313 , \26015_26314 , \26016_26315 , \26017_26316 , \26018_26317 , \26019_26318 , \26020_26319 , \26021_26320 , \26022_26321 , \26023_26322 , \26024_26323 , \26025_26324 , \26026_26325 , \26027_26326 , \26028_26327 , \26029_26328 , \26030_26329 , \26031_26330 , \26032_26331 , \26033_26332 , \26034_26333 , \26035_26334 , \26036_26335 , \26037_26336 , \26038_26337 , \26039_26338 , \26040_26339 , \26041_26340 , \26042_26341 , \26043_26342 , \26044_26343 );
and \U$17222 ( \26046_26345 , RIfcb23a0_7050, \9163_9462 );
and \U$17223 ( \26047_26346 , RIfc5bbe0_6066, \9165_9464 );
and \U$17224 ( \26048_26347 , RIfcede78_7729, \9167_9466 );
and \U$17225 ( \26049_26348 , RIe1fa370_4224, \9169_9468 );
and \U$17226 ( \26050_26349 , RIfcd4c48_7443, \9171_9470 );
and \U$17227 ( \26051_26350 , RIfce1dd0_7592, \9173_9472 );
and \U$17228 ( \26052_26351 , RIfcbf960_7202, \9175_9474 );
and \U$17229 ( \26053_26352 , RIe1f58e8_4171, \9177_9476 );
and \U$17230 ( \26054_26353 , RIfcbfc30_7204, \9179_9478 );
and \U$17231 ( \26055_26354 , RIfc78380_6390, \9181_9480 );
and \U$17232 ( \26056_26355 , RIfc93770_6700, \9183_9482 );
and \U$17233 ( \26057_26356 , RIe1f35c0_4146, \9185_9484 );
and \U$17234 ( \26058_26357 , RIfcb1f68_7047, \9187_9486 );
and \U$17235 ( \26059_26358 , RIfce1b00_7590, \9189_9488 );
and \U$17236 ( \26060_26359 , RIfc93a40_6702, \9191_9490 );
and \U$17237 ( \26061_26360 , RIe1ee2c8_4087, \9193_9492 );
and \U$17238 ( \26062_26361 , RIe1ebb68_4059, \9195_9494 );
and \U$17239 ( \26063_26362 , RIe1e8e68_4027, \9197_9496 );
and \U$17240 ( \26064_26363 , RIe1e6168_3995, \9199_9498 );
and \U$17241 ( \26065_26364 , RIe1e3468_3963, \9201_9500 );
and \U$17242 ( \26066_26365 , RIe1e0768_3931, \9203_9502 );
and \U$17243 ( \26067_26366 , RIe1dda68_3899, \9205_9504 );
and \U$17244 ( \26068_26367 , RIe1dad68_3867, \9207_9506 );
and \U$17245 ( \26069_26368 , RIe1d8068_3835, \9209_9508 );
and \U$17246 ( \26070_26369 , RIe1d2668_3771, \9211_9510 );
and \U$17247 ( \26071_26370 , RIe1cf968_3739, \9213_9512 );
and \U$17248 ( \26072_26371 , RIe1ccc68_3707, \9215_9514 );
and \U$17249 ( \26073_26372 , RIe1c9f68_3675, \9217_9516 );
and \U$17250 ( \26074_26373 , RIe1c7268_3643, \9219_9518 );
and \U$17251 ( \26075_26374 , RIe1c4568_3611, \9221_9520 );
and \U$17252 ( \26076_26375 , RIe1c1868_3579, \9223_9522 );
and \U$17253 ( \26077_26376 , RIe1beb68_3547, \9225_9524 );
and \U$17254 ( \26078_26377 , RIfcdec98_7557, \9227_9526 );
and \U$17255 ( \26079_26378 , RIfc94148_6707, \9229_9528 );
and \U$17256 ( \26080_26379 , RIe1b95a0_3486, \9231_9530 );
and \U$17257 ( \26081_26380 , RIe1b7548_3463, \9233_9532 );
and \U$17258 ( \26082_26381 , RIfcd12a0_7402, \9235_9534 );
and \U$17259 ( \26083_26382 , RIfceabd8_7693, \9237_9536 );
and \U$17260 ( \26084_26383 , RIe1b5388_3439, \9239_9538 );
and \U$17261 ( \26085_26384 , RIe1b3fd8_3425, \9241_9540 );
and \U$17262 ( \26086_26385 , RIfc94850_6712, \9243_9542 );
and \U$17263 ( \26087_26386 , RIfcd7c18_7477, \9245_9544 );
and \U$17264 ( \26088_26387 , RIe1b27f0_3408, \9247_9546 );
and \U$17265 ( \26089_26388 , RIe1b0d38_3389, \9249_9548 );
and \U$17266 ( \26090_26389 , RIfc76a30_6372, \9251_9550 );
and \U$17267 ( \26091_26390 , RIfce2640_7598, \9253_9552 );
and \U$17268 ( \26092_26391 , RIe1ac6e8_3339, \9255_9554 );
and \U$17269 ( \26093_26392 , RIe1ab068_3323, \9257_9556 );
and \U$17270 ( \26094_26393 , RIe1a8ea8_3299, \9259_9558 );
and \U$17271 ( \26095_26394 , RIe1a61a8_3267, \9261_9560 );
and \U$17272 ( \26096_26395 , RIe1a34a8_3235, \9263_9562 );
and \U$17273 ( \26097_26396 , RIe1a07a8_3203, \9265_9564 );
and \U$17274 ( \26098_26397 , RIe18cca8_2979, \9267_9566 );
and \U$17275 ( \26099_26398 , RIe1791a8_2755, \9269_9568 );
and \U$17276 ( \26100_26399 , RIe226b00_4730, \9271_9570 );
and \U$17277 ( \26101_26400 , RIe21b700_4602, \9273_9572 );
and \U$17278 ( \26102_26401 , RIe204f00_4346, \9275_9574 );
and \U$17279 ( \26103_26402 , RIe1fef60_4278, \9277_9576 );
and \U$17280 ( \26104_26403 , RIe1f8318_4201, \9279_9578 );
and \U$17281 ( \26105_26404 , RIe1f0e60_4118, \9281_9580 );
and \U$17282 ( \26106_26405 , RIe1d5368_3803, \9283_9582 );
and \U$17283 ( \26107_26406 , RIe1bbe68_3515, \9285_9584 );
and \U$17284 ( \26108_26407 , RIe1aece0_3366, \9287_9586 );
and \U$17285 ( \26109_26408 , RIe171318_2665, \9289_9588 );
or \U$17286 ( \26110_26409 , \26046_26345 , \26047_26346 , \26048_26347 , \26049_26348 , \26050_26349 , \26051_26350 , \26052_26351 , \26053_26352 , \26054_26353 , \26055_26354 , \26056_26355 , \26057_26356 , \26058_26357 , \26059_26358 , \26060_26359 , \26061_26360 , \26062_26361 , \26063_26362 , \26064_26363 , \26065_26364 , \26066_26365 , \26067_26366 , \26068_26367 , \26069_26368 , \26070_26369 , \26071_26370 , \26072_26371 , \26073_26372 , \26074_26373 , \26075_26374 , \26076_26375 , \26077_26376 , \26078_26377 , \26079_26378 , \26080_26379 , \26081_26380 , \26082_26381 , \26083_26382 , \26084_26383 , \26085_26384 , \26086_26385 , \26087_26386 , \26088_26387 , \26089_26388 , \26090_26389 , \26091_26390 , \26092_26391 , \26093_26392 , \26094_26393 , \26095_26394 , \26096_26395 , \26097_26396 , \26098_26397 , \26099_26398 , \26100_26399 , \26101_26400 , \26102_26401 , \26103_26402 , \26104_26403 , \26105_26404 , \26106_26405 , \26107_26406 , \26108_26407 , \26109_26408 );
or \U$17287 ( \26111_26410 , \26045_26344 , \26110_26409 );
_DC \g3705/U$1 ( \26112 , \26111_26410 , \9298_9597 );
buf \U$17288 ( \26113_26412 , \26112 );
and \U$17289 ( \26114_26413 , \25980_26279 , \26113_26412 );
and \U$17290 ( \26115_26414 , \24074_24373 , \24207_24506 );
and \U$17291 ( \26116_26415 , \24207_24506 , \24482_24781 );
and \U$17292 ( \26117_26416 , \24074_24373 , \24482_24781 );
or \U$17293 ( \26118_26417 , \26115_26414 , \26116_26415 , \26117_26416 );
and \U$17294 ( \26119_26418 , \26113_26412 , \26118_26417 );
and \U$17295 ( \26120_26419 , \25980_26279 , \26118_26417 );
or \U$17296 ( \26121_26420 , \26114_26413 , \26119_26418 , \26120_26419 );
xor \U$17297 ( \26122_26421 , \25847_26146 , \26121_26420 );
buf g440c_GF_PartitionCandidate( \26123_26422_nG440c , \26122_26421 );
xor \U$17298 ( \26124_26423 , \25980_26279 , \26113_26412 );
xor \U$17299 ( \26125_26424 , \26124_26423 , \26118_26417 );
buf g440f_GF_PartitionCandidate( \26126_26425_nG440f , \26125_26424 );
nand \U$17300 ( \26127_26426 , \26126_26425_nG440f , \24484_24783_nG4412 );
and \U$17301 ( \26128_26427 , \26123_26422_nG440c , \26127_26426 );
xor \U$17302 ( \26129_26428 , \26126_26425_nG440f , \24484_24783_nG4412 );
and \U$17307 ( \26130_26432 , \26129_26428 , \10392_10694_nG9c0e );
or \U$17308 ( \26131_26433 , 1'b0 , \26130_26432 );
xor \U$17309 ( \26132_26434 , \26128_26427 , \26131_26433 );
xor \U$17310 ( \26133_26435 , \26128_26427 , \26132_26434 );
buf \U$17311 ( \26134_26436 , \26133_26435 );
buf \U$17312 ( \26135_26437 , \26134_26436 );
xor \U$17313 ( \26136_26438 , \25580_25879 , \26135_26437 );
and \U$17314 ( \26137_26439 , \25150_25449 , \25155_25454 );
and \U$17315 ( \26138_26440 , \25150_25449 , \25568_25867 );
and \U$17316 ( \26139_26441 , \25155_25454 , \25568_25867 );
or \U$17317 ( \26140_26442 , \26137_26439 , \26138_26440 , \26139_26441 );
and \U$17318 ( \26141_26443 , \26136_26438 , \26140_26442 );
and \U$17319 ( \26142_26444 , \25161_25460 , \25166_25465 );
and \U$17320 ( \26143_26445 , \25161_25460 , \25566_25865 );
and \U$17321 ( \26144_26446 , \25166_25465 , \25566_25865 );
or \U$17322 ( \26145_26447 , \26142_26444 , \26143_26445 , \26144_26446 );
buf \U$17323 ( \26146_26448 , \26145_26447 );
and \U$17324 ( \26147_26449 , \25041_25343 , \25050_25349 );
and \U$17325 ( \26148_26450 , \25041_25343 , \25057_25356 );
and \U$17326 ( \26149_26451 , \25050_25349 , \25057_25356 );
or \U$17327 ( \26150_26452 , \26147_26449 , \26148_26450 , \26149_26451 );
buf \U$17328 ( \26151_26453 , \26150_26452 );
and \U$17329 ( \26152_26454 , \25044_24792 , \10693_10995_nG9c0b );
and \U$17330 ( \26153_26455 , \24490_24789 , \10981_11283_nG9c08 );
or \U$17331 ( \26154_26456 , \26152_26454 , \26153_26455 );
xor \U$17332 ( \26155_26457 , \24489_24788 , \26154_26456 );
buf \U$17333 ( \26156_26458 , \26155_26457 );
buf \U$17335 ( \26157_26459 , \26156_26458 );
and \U$17336 ( \26158_26460 , \23495_23201 , \11299_11598_nG9c05 );
and \U$17337 ( \26159_26461 , \22899_23198 , \12168_12470_nG9c02 );
or \U$17338 ( \26160_26462 , \26158_26460 , \26159_26461 );
xor \U$17339 ( \26161_26463 , \22898_23197 , \26160_26462 );
buf \U$17340 ( \26162_26464 , \26161_26463 );
buf \U$17342 ( \26163_26465 , \26162_26464 );
xor \U$17343 ( \26164_26466 , \26157_26459 , \26163_26465 );
buf \U$17344 ( \26165_26467 , \26164_26466 );
xor \U$17345 ( \26166_26468 , \26151_26453 , \26165_26467 );
and \U$17346 ( \26167_26469 , \18908_18702 , \15074_15373_nG9bf3 );
and \U$17347 ( \26168_26470 , \18400_18699 , \16013_16315_nG9bf0 );
or \U$17348 ( \26169_26471 , \26167_26469 , \26168_26470 );
xor \U$17349 ( \26170_26472 , \18399_18698 , \26169_26471 );
buf \U$17350 ( \26171_26473 , \26170_26472 );
buf \U$17352 ( \26172_26474 , \26171_26473 );
xor \U$17353 ( \26173_26475 , \26166_26468 , \26172_26474 );
buf \U$17354 ( \26174_26476 , \26173_26475 );
and \U$17355 ( \26175_26477 , \16405_15940 , \17808_18107_nG9be7 );
and \U$17356 ( \26176_26478 , \15638_15937 , \18789_19091_nG9be4 );
or \U$17357 ( \26177_26479 , \26175_26477 , \26176_26478 );
xor \U$17358 ( \26178_26480 , \15637_15936 , \26177_26479 );
buf \U$17359 ( \26179_26481 , \26178_26480 );
buf \U$17361 ( \26180_26482 , \26179_26481 );
xor \U$17362 ( \26181_26483 , \26174_26476 , \26180_26482 );
and \U$17363 ( \26182_26484 , \14710_14631 , \19287_19586_nG9be1 );
and \U$17364 ( \26183_26485 , \14329_14628 , \20306_20608_nG9bde );
or \U$17365 ( \26184_26486 , \26182_26484 , \26183_26485 );
xor \U$17366 ( \26185_26487 , \14328_14627 , \26184_26486 );
buf \U$17367 ( \26186_26488 , \26185_26487 );
buf \U$17369 ( \26187_26489 , \26186_26488 );
xor \U$17370 ( \26188_26490 , \26181_26483 , \26187_26489 );
buf \U$17371 ( \26189_26491 , \26188_26490 );
and \U$17372 ( \26190_26492 , \25068_25367 , \25074_25373 );
and \U$17373 ( \26191_26493 , \25068_25367 , \25081_25380 );
and \U$17374 ( \26192_26494 , \25074_25373 , \25081_25380 );
or \U$17375 ( \26193_26495 , \26190_26492 , \26191_26493 , \26192_26494 );
buf \U$17376 ( \26194_26496 , \26193_26495 );
xor \U$17377 ( \26195_26497 , \26189_26491 , \26194_26496 );
and \U$17378 ( \26196_26498 , \10411_10707 , \25561_25860_nG9bc9 );
and \U$17379 ( \26197_26499 , \25181_25480 , \25487_25786 );
and \U$17380 ( \26198_26500 , \25487_25786 , \25549_25848 );
and \U$17381 ( \26199_26501 , \25181_25480 , \25549_25848 );
or \U$17382 ( \26200_26502 , \26197_26499 , \26198_26500 , \26199_26501 );
and \U$17383 ( \26201_26503 , \25511_25810 , \25532_25831 );
and \U$17384 ( \26202_26504 , \25532_25831 , \25547_25846 );
and \U$17385 ( \26203_26505 , \25511_25810 , \25547_25846 );
or \U$17386 ( \26204_26506 , \26201_26503 , \26202_26504 , \26203_26505 );
and \U$17387 ( \26205_26507 , \25189_25488 , \25193_25492 );
and \U$17388 ( \26206_26508 , \25193_25492 , \25198_25497 );
and \U$17389 ( \26207_26509 , \25189_25488 , \25198_25497 );
or \U$17390 ( \26208_26510 , \26205_26507 , \26206_26508 , \26207_26509 );
and \U$17391 ( \26209_26511 , \25519_25818 , \25523_25822 );
and \U$17392 ( \26210_26512 , \25523_25822 , \25531_25830 );
and \U$17393 ( \26211_26513 , \25519_25818 , \25531_25830 );
or \U$17394 ( \26212_26514 , \26209_26511 , \26210_26512 , \26211_26513 );
xor \U$17395 ( \26213_26515 , \26208_26510 , \26212_26514 );
and \U$17396 ( \26214_26516 , \22257_22556 , \12491_12790 );
and \U$17397 ( \26215_26517 , \23315_23617 , \12159_12461 );
nor \U$17398 ( \26216_26518 , \26214_26516 , \26215_26517 );
xnor \U$17399 ( \26217_26519 , \26216_26518 , \12481_12780 );
and \U$17400 ( \26218_26520 , \17736_18035 , \16333_16635 );
and \U$17401 ( \26219_26521 , \18730_19032 , \15999_16301 );
nor \U$17402 ( \26220_26522 , \26218_26520 , \26219_26521 );
xnor \U$17403 ( \26221_26523 , \26220_26522 , \16323_16625 );
xor \U$17404 ( \26222_26524 , \26217_26519 , \26221_26523 );
and \U$17405 ( \26223_26525 , \10686_10988 , \25527_25826 );
and \U$17406 ( \26224_26526 , \10968_11270 , \24962_25264 );
nor \U$17407 ( \26225_26527 , \26223_26525 , \26224_26526 );
xnor \U$17408 ( \26226_26528 , \26225_26527 , \25474_25773 );
xor \U$17409 ( \26227_26529 , \26222_26524 , \26226_26528 );
xor \U$17410 ( \26228_26530 , \26213_26515 , \26227_26529 );
xor \U$17411 ( \26229_26531 , \26204_26506 , \26228_26530 );
and \U$17412 ( \26230_26532 , \23900_24199 , \11275_11574 );
and \U$17413 ( \26231_26533 , \24970_25272 , \10976_11278 );
nor \U$17414 ( \26232_26534 , \26230_26532 , \26231_26533 );
xnor \U$17415 ( \26233_26535 , \26232_26534 , \11281_11580 );
and \U$17416 ( \26234_26536 , \20734_21033 , \13755_14054 );
and \U$17417 ( \26235_26537 , \21788_22090 , \13390_13692 );
nor \U$17418 ( \26236_26538 , \26234_26536 , \26235_26537 );
xnor \U$17419 ( \26237_26539 , \26236_26538 , \13736_14035 );
xor \U$17420 ( \26238_26540 , \26233_26535 , \26237_26539 );
and \U$17421 ( \26239_26541 , RIdec5810_711, \9034_9333 );
and \U$17422 ( \26240_26542 , RIdec2b10_679, \9036_9335 );
and \U$17423 ( \26241_26543 , RIfce6f60_7650, \9038_9337 );
and \U$17424 ( \26242_26544 , RIdebfe10_647, \9040_9339 );
and \U$17425 ( \26243_26545 , RIfc95228_6719, \9042_9341 );
and \U$17426 ( \26244_26546 , RIdebd110_615, \9044_9343 );
and \U$17427 ( \26245_26547 , RIdeba410_583, \9046_9345 );
and \U$17428 ( \26246_26548 , RIdeb7710_551, \9048_9347 );
and \U$17429 ( \26247_26549 , RIfe879a8_7887, \9050_9349 );
and \U$17430 ( \26248_26550 , RIdeb1d10_487, \9052_9351 );
and \U$17431 ( \26249_26551 , RIfcc16e8_7223, \9054_9353 );
and \U$17432 ( \26250_26552 , RIdeaf010_455, \9056_9355 );
and \U$17433 ( \26251_26553 , RIfca4f48_6899, \9058_9357 );
and \U$17434 ( \26252_26554 , RIdeaadf8_423, \9060_9359 );
and \U$17435 ( \26253_26555 , RIdea44f8_391, \9062_9361 );
and \U$17436 ( \26254_26556 , RIde9dbf8_359, \9064_9363 );
and \U$17437 ( \26255_26557 , RIee1cf48_4788, \9066_9365 );
and \U$17438 ( \26256_26558 , RIee1bfd0_4777, \9068_9367 );
and \U$17439 ( \26257_26559 , RIfc95660_6722, \9070_9369 );
and \U$17440 ( \26258_26560 , RIfcee148_7731, \9072_9371 );
and \U$17441 ( \26259_26561 , RIfe87840_7886, \9074_9373 );
and \U$17442 ( \26260_26562 , RIfe876d8_7885, \9076_9375 );
and \U$17443 ( \26261_26563 , RIde8a0f8_263, \9078_9377 );
and \U$17444 ( \26262_26564 , RIde85f58_243, \9080_9379 );
and \U$17445 ( \26263_26565 , RIfcb0780_7030, \9082_9381 );
and \U$17446 ( \26264_26566 , RIfcee9b8_7737, \9084_9383 );
and \U$17447 ( \26265_26567 , RIfc5f150_6104, \9086_9385 );
and \U$17448 ( \26266_26568 , RIfcdee00_7558, \9088_9387 );
and \U$17449 ( \26267_26569 , RIfcd8050_7480, \9090_9389 );
and \U$17450 ( \26268_26570 , RIe16ba80_2602, \9092_9391 );
and \U$17451 ( \26269_26571 , RIfca5380_6902, \9094_9393 );
and \U$17452 ( \26270_26572 , RIe1680d8_2561, \9096_9395 );
and \U$17453 ( \26271_26573 , RIe165810_2532, \9098_9397 );
and \U$17454 ( \26272_26574 , RIe162b10_2500, \9100_9399 );
and \U$17455 ( \26273_26575 , RIee377f8_5090, \9102_9401 );
and \U$17456 ( \26274_26576 , RIe15fe10_2468, \9104_9403 );
and \U$17457 ( \26275_26577 , RIee36448_5076, \9106_9405 );
and \U$17458 ( \26276_26578 , RIe15d110_2436, \9108_9407 );
and \U$17459 ( \26277_26579 , RIe157710_2372, \9110_9409 );
and \U$17460 ( \26278_26580 , RIe154a10_2340, \9112_9411 );
and \U$17461 ( \26279_26581 , RIfc3f3c8_5745, \9114_9413 );
and \U$17462 ( \26280_26582 , RIe151d10_2308, \9116_9415 );
and \U$17463 ( \26281_26583 , RIfcde9c8_7555, \9118_9417 );
and \U$17464 ( \26282_26584 , RIe14f010_2276, \9120_9419 );
and \U$17465 ( \26283_26585 , RIfc4a2a0_5866, \9122_9421 );
and \U$17466 ( \26284_26586 , RIe14c310_2244, \9124_9423 );
and \U$17467 ( \26285_26587 , RIe149610_2212, \9126_9425 );
and \U$17468 ( \26286_26588 , RIe146910_2180, \9128_9427 );
and \U$17469 ( \26287_26589 , RIfc62288_6139, \9130_9429 );
and \U$17470 ( \26288_26590 , RIee33478_5042, \9132_9431 );
and \U$17471 ( \26289_26591 , RIfc71b70_6316, \9134_9433 );
and \U$17472 ( \26290_26592 , RIee312b8_5018, \9136_9435 );
and \U$17473 ( \26291_26593 , RIe1411e0_2118, \9138_9437 );
and \U$17474 ( \26292_26594 , RIfe87570_7884, \9140_9439 );
and \U$17475 ( \26293_26595 , RIdf3cf28_2070, \9142_9441 );
and \U$17476 ( \26294_26596 , RIfe87408_7883, \9144_9443 );
and \U$17477 ( \26295_26597 , RIfcc99b0_7316, \9146_9445 );
and \U$17478 ( \26296_26598 , RIfccf0e0_7378, \9148_9447 );
and \U$17479 ( \26297_26599 , RIfcaeb60_7010, \9150_9449 );
and \U$17480 ( \26298_26600 , RIfcca220_7322, \9152_9451 );
and \U$17481 ( \26299_26601 , RIdf35bd8_1988, \9154_9453 );
and \U$17482 ( \26300_26602 , RIdf33748_1962, \9156_9455 );
and \U$17483 ( \26301_26603 , RIdf31588_1938, \9158_9457 );
and \U$17484 ( \26302_26604 , RIdf2f530_1915, \9160_9459 );
or \U$17485 ( \26303_26605 , \26239_26541 , \26240_26542 , \26241_26543 , \26242_26544 , \26243_26545 , \26244_26546 , \26245_26547 , \26246_26548 , \26247_26549 , \26248_26550 , \26249_26551 , \26250_26552 , \26251_26553 , \26252_26554 , \26253_26555 , \26254_26556 , \26255_26557 , \26256_26558 , \26257_26559 , \26258_26560 , \26259_26561 , \26260_26562 , \26261_26563 , \26262_26564 , \26263_26565 , \26264_26566 , \26265_26567 , \26266_26568 , \26267_26569 , \26268_26570 , \26269_26571 , \26270_26572 , \26271_26573 , \26272_26574 , \26273_26575 , \26274_26576 , \26275_26577 , \26276_26578 , \26277_26579 , \26278_26580 , \26279_26581 , \26280_26582 , \26281_26583 , \26282_26584 , \26283_26585 , \26284_26586 , \26285_26587 , \26286_26588 , \26287_26589 , \26288_26590 , \26289_26591 , \26290_26592 , \26291_26593 , \26292_26594 , \26293_26595 , \26294_26596 , \26295_26597 , \26296_26598 , \26297_26599 , \26298_26600 , \26299_26601 , \26300_26602 , \26301_26603 , \26302_26604 );
and \U$17486 ( \26304_26606 , RIee2be58_4958, \9163_9462 );
and \U$17487 ( \26305_26607 , RIee2a508_4940, \9165_9464 );
and \U$17488 ( \26306_26608 , RIee28ff0_4925, \9167_9466 );
and \U$17489 ( \26307_26609 , RIee27da8_4912, \9169_9468 );
and \U$17490 ( \26308_26610 , RIdf2a508_1858, \9171_9470 );
and \U$17491 ( \26309_26611 , RIdf28348_1834, \9173_9472 );
and \U$17492 ( \26310_26612 , RIdf265c0_1813, \9175_9474 );
and \U$17493 ( \26311_26613 , RIdf24b08_1794, \9177_9476 );
and \U$17494 ( \26312_26614 , RIfc74708_6347, \9179_9478 );
and \U$17495 ( \26313_26615 , RIfc42578_5777, \9181_9480 );
and \U$17496 ( \26314_26616 , RIfc43388_5787, \9183_9482 );
and \U$17497 ( \26315_26617 , RIfc745a0_6346, \9185_9484 );
and \U$17498 ( \26316_26618 , RIfcb0078_7025, \9187_9486 );
and \U$17499 ( \26317_26619 , RIdf1fc48_1738, \9189_9488 );
and \U$17500 ( \26318_26620 , RIfcaff10_7024, \9191_9490 );
and \U$17501 ( \26319_26621 , RIdf195a0_1665, \9193_9492 );
and \U$17502 ( \26320_26622 , RIdf173e0_1641, \9195_9494 );
and \U$17503 ( \26321_26623 , RIdf146e0_1609, \9197_9496 );
and \U$17504 ( \26322_26624 , RIdf119e0_1577, \9199_9498 );
and \U$17505 ( \26323_26625 , RIdf0ece0_1545, \9201_9500 );
and \U$17506 ( \26324_26626 , RIdf0bfe0_1513, \9203_9502 );
and \U$17507 ( \26325_26627 , RIdf092e0_1481, \9205_9504 );
and \U$17508 ( \26326_26628 , RIdf065e0_1449, \9207_9506 );
and \U$17509 ( \26327_26629 , RIdf038e0_1417, \9209_9508 );
and \U$17510 ( \26328_26630 , RIdefdee0_1353, \9211_9510 );
and \U$17511 ( \26329_26631 , RIdefb1e0_1321, \9213_9512 );
and \U$17512 ( \26330_26632 , RIdef84e0_1289, \9215_9514 );
and \U$17513 ( \26331_26633 , RIdef57e0_1257, \9217_9516 );
and \U$17514 ( \26332_26634 , RIdef2ae0_1225, \9219_9518 );
and \U$17515 ( \26333_26635 , RIdeefde0_1193, \9221_9520 );
and \U$17516 ( \26334_26636 , RIdeed0e0_1161, \9223_9522 );
and \U$17517 ( \26335_26637 , RIdeea3e0_1129, \9225_9524 );
and \U$17518 ( \26336_26638 , RIee257b0_4885, \9227_9526 );
and \U$17519 ( \26337_26639 , RIfca73d8_6925, \9229_9528 );
and \U$17520 ( \26338_26640 , RIee23e60_4867, \9231_9530 );
and \U$17521 ( \26339_26641 , RIfce66f0_7644, \9233_9532 );
and \U$17522 ( \26340_26642 , RIdee4cb0_1067, \9235_9534 );
and \U$17523 ( \26341_26643 , RIdee2f28_1046, \9237_9536 );
and \U$17524 ( \26342_26644 , RIdee0d68_1022, \9239_9538 );
and \U$17525 ( \26343_26645 , RIdeded10_999, \9241_9540 );
and \U$17526 ( \26344_26646 , RIfcca388_7323, \9243_9542 );
and \U$17527 ( \26345_26647 , RIfce6858_7645, \9245_9544 );
and \U$17528 ( \26346_26648 , RIfcceca8_7375, \9247_9546 );
and \U$17529 ( \26347_26649 , RIfcdc970_7532, \9249_9548 );
and \U$17530 ( \26348_26650 , RIded9b80_941, \9251_9550 );
and \U$17531 ( \26349_26651 , RIfeaaac0_8258, \9253_9552 );
and \U$17532 ( \26350_26652 , RIded5800_893, \9255_9554 );
and \U$17533 ( \26351_26653 , RIded3208_866, \9257_9556 );
and \U$17534 ( \26352_26654 , RIded0c10_839, \9259_9558 );
and \U$17535 ( \26353_26655 , RIdecdf10_807, \9261_9560 );
and \U$17536 ( \26354_26656 , RIdecb210_775, \9263_9562 );
and \U$17537 ( \26355_26657 , RIdec8510_743, \9265_9564 );
and \U$17538 ( \26356_26658 , RIdeb4a10_519, \9267_9566 );
and \U$17539 ( \26357_26659 , RIde972f8_327, \9269_9568 );
and \U$17540 ( \26358_26660 , RIe16e618_2633, \9271_9570 );
and \U$17541 ( \26359_26661 , RIe15a410_2404, \9273_9572 );
and \U$17542 ( \26360_26662 , RIe143c10_2148, \9275_9574 );
and \U$17543 ( \26361_26663 , RIdf38608_2018, \9277_9576 );
and \U$17544 ( \26362_26664 , RIdf2cc68_1886, \9279_9578 );
and \U$17545 ( \26363_26665 , RIdf1d4e8_1710, \9281_9580 );
and \U$17546 ( \26364_26666 , RIdf00be0_1385, \9283_9582 );
and \U$17547 ( \26365_26667 , RIdee76e0_1097, \9285_9584 );
and \U$17548 ( \26366_26668 , RIdedc448_970, \9287_9586 );
and \U$17549 ( \26367_26669 , RIde7d240_200, \9289_9588 );
or \U$17550 ( \26368_26670 , \26304_26606 , \26305_26607 , \26306_26608 , \26307_26609 , \26308_26610 , \26309_26611 , \26310_26612 , \26311_26613 , \26312_26614 , \26313_26615 , \26314_26616 , \26315_26617 , \26316_26618 , \26317_26619 , \26318_26620 , \26319_26621 , \26320_26622 , \26321_26623 , \26322_26624 , \26323_26625 , \26324_26626 , \26325_26627 , \26326_26628 , \26327_26629 , \26328_26630 , \26329_26631 , \26330_26632 , \26331_26633 , \26332_26634 , \26333_26635 , \26334_26636 , \26335_26637 , \26336_26638 , \26337_26639 , \26338_26640 , \26339_26641 , \26340_26642 , \26341_26643 , \26342_26644 , \26343_26645 , \26344_26646 , \26345_26647 , \26346_26648 , \26347_26649 , \26348_26650 , \26349_26651 , \26350_26652 , \26351_26653 , \26352_26654 , \26353_26655 , \26354_26656 , \26355_26657 , \26356_26658 , \26357_26659 , \26358_26660 , \26359_26661 , \26360_26662 , \26361_26663 , \26362_26664 , \26363_26665 , \26364_26666 , \26365_26667 , \26366_26668 , \26367_26669 );
or \U$17551 ( \26369_26671 , \26303_26605 , \26368_26670 );
_DC \g5db2/U$1 ( \26370 , \26369_26671 , \9298_9597 );
and \U$17552 ( \26371_26673 , RIe19daa8_3171, \8760_9059 );
and \U$17553 ( \26372_26674 , RIe19ada8_3139, \8762_9061 );
and \U$17554 ( \26373_26675 , RIf1457c0_5250, \8764_9063 );
and \U$17555 ( \26374_26676 , RIe1980a8_3107, \8766_9065 );
and \U$17556 ( \26375_26677 , RIf1449b0_5240, \8768_9067 );
and \U$17557 ( \26376_26678 , RIe1953a8_3075, \8770_9069 );
and \U$17558 ( \26377_26679 , RIe1926a8_3043, \8772_9071 );
and \U$17559 ( \26378_26680 , RIe18f9a8_3011, \8774_9073 );
and \U$17560 ( \26379_26681 , RIe189fa8_2947, \8776_9075 );
and \U$17561 ( \26380_26682 , RIe1872a8_2915, \8778_9077 );
and \U$17562 ( \26381_26683 , RIf143ba0_5230, \8780_9079 );
and \U$17563 ( \26382_26684 , RIe1845a8_2883, \8782_9081 );
and \U$17564 ( \26383_26685 , RIfc912e0_6674, \8784_9083 );
and \U$17565 ( \26384_26686 , RIe1818a8_2851, \8786_9085 );
and \U$17566 ( \26385_26687 , RIe17eba8_2819, \8788_9087 );
and \U$17567 ( \26386_26688 , RIe17bea8_2787, \8790_9089 );
and \U$17568 ( \26387_26689 , RIfc915b0_6676, \8792_9091 );
and \U$17569 ( \26388_26690 , RIfcbe5b0_7188, \8794_9093 );
and \U$17570 ( \26389_26691 , RIfce3b58_7613, \8796_9095 );
and \U$17571 ( \26390_26692 , RIe175da0_2718, \8798_9097 );
and \U$17572 ( \26391_26693 , RIfceb448_7699, \8800_9099 );
and \U$17573 ( \26392_26694 , RIfcc7958_7293, \8802_9101 );
and \U$17574 ( \26393_26695 , RIfc42de8_5783, \8804_9103 );
and \U$17575 ( \26394_26696 , RIfc96e48_6739, \8806_9105 );
and \U$17576 ( \26395_26697 , RIfc7a810_6416, \8808_9107 );
and \U$17577 ( \26396_26698 , RIfc96ce0_6738, \8810_9109 );
and \U$17578 ( \26397_26699 , RIfcc7ac0_7294, \8812_9111 );
and \U$17579 ( \26398_26700 , RIe173be0_2694, \8814_9113 );
and \U$17580 ( \26399_26701 , RIfce39f0_7612, \8816_9115 );
and \U$17581 ( \26400_26702 , RIfc7a540_6414, \8818_9117 );
and \U$17582 ( \26401_26703 , RIfc91b50_6680, \8820_9119 );
and \U$17583 ( \26402_26704 , RIfc429b0_5780, \8822_9121 );
and \U$17584 ( \26403_26705 , RIfea9710_8244, \8824_9123 );
and \U$17585 ( \26404_26706 , RIe223e00_4698, \8826_9125 );
and \U$17586 ( \26405_26707 , RIfcd8488_7483, \8828_9127 );
and \U$17587 ( \26406_26708 , RIe221100_4666, \8830_9129 );
and \U$17588 ( \26407_26709 , RIfc920f0_6684, \8832_9131 );
and \U$17589 ( \26408_26710 , RIe21e400_4634, \8834_9133 );
and \U$17590 ( \26409_26711 , RIe218a00_4570, \8836_9135 );
and \U$17591 ( \26410_26712 , RIe215d00_4538, \8838_9137 );
and \U$17592 ( \26411_26713 , RIfc79e38_6409, \8840_9139 );
and \U$17593 ( \26412_26714 , RIe213000_4506, \8842_9141 );
and \U$17594 ( \26413_26715 , RIfcbee20_7194, \8844_9143 );
and \U$17595 ( \26414_26716 , RIe210300_4474, \8846_9145 );
and \U$17596 ( \26415_26717 , RIf168068_5643, \8848_9147 );
and \U$17597 ( \26416_26718 , RIe20d600_4442, \8850_9149 );
and \U$17598 ( \26417_26719 , RIe20a900_4410, \8852_9151 );
and \U$17599 ( \26418_26720 , RIe207c00_4378, \8854_9153 );
and \U$17600 ( \26419_26721 , RIfc5af38_6057, \8856_9155 );
and \U$17601 ( \26420_26722 , RIfcd73a8_7471, \8858_9157 );
and \U$17602 ( \26421_26723 , RIe2027a0_4318, \8860_9159 );
and \U$17603 ( \26422_26724 , RIe200ce8_4299, \8862_9161 );
and \U$17604 ( \26423_26725 , RIfcb2670_7052, \8864_9163 );
and \U$17605 ( \26424_26726 , RIfcdf940_7566, \8866_9165 );
and \U$17606 ( \26425_26727 , RIfc5b208_6059, \8868_9167 );
and \U$17607 ( \26426_26728 , RIfcbf3c0_7198, \8870_9169 );
and \U$17608 ( \26427_26729 , RIf1604a8_5555, \8872_9171 );
and \U$17609 ( \26428_26730 , RIf15e5b8_5533, \8874_9173 );
and \U$17610 ( \26429_26731 , RIfe872a0_7882, \8876_9175 );
and \U$17611 ( \26430_26732 , RIfe87138_7881, \8878_9177 );
and \U$17612 ( \26431_26733 , RIfc78920_6394, \8880_9179 );
and \U$17613 ( \26432_26734 , RIfec1158_8317, \8882_9181 );
and \U$17614 ( \26433_26735 , RIfc93338_6697, \8884_9183 );
and \U$17615 ( \26434_26736 , RIfcea368_7687, \8886_9185 );
or \U$17616 ( \26435_26737 , \26371_26673 , \26372_26674 , \26373_26675 , \26374_26676 , \26375_26677 , \26376_26678 , \26377_26679 , \26378_26680 , \26379_26681 , \26380_26682 , \26381_26683 , \26382_26684 , \26383_26685 , \26384_26686 , \26385_26687 , \26386_26688 , \26387_26689 , \26388_26690 , \26389_26691 , \26390_26692 , \26391_26693 , \26392_26694 , \26393_26695 , \26394_26696 , \26395_26697 , \26396_26698 , \26397_26699 , \26398_26700 , \26399_26701 , \26400_26702 , \26401_26703 , \26402_26704 , \26403_26705 , \26404_26706 , \26405_26707 , \26406_26708 , \26407_26709 , \26408_26710 , \26409_26711 , \26410_26712 , \26411_26713 , \26412_26714 , \26413_26715 , \26414_26716 , \26415_26717 , \26416_26718 , \26417_26719 , \26418_26720 , \26419_26721 , \26420_26722 , \26421_26723 , \26422_26724 , \26423_26725 , \26424_26726 , \26425_26727 , \26426_26728 , \26427_26729 , \26428_26730 , \26429_26731 , \26430_26732 , \26431_26733 , \26432_26734 , \26433_26735 , \26434_26736 );
and \U$17617 ( \26436_26738 , RIfcb23a0_7050, \8889_9188 );
and \U$17618 ( \26437_26739 , RIfc5bbe0_6066, \8891_9190 );
and \U$17619 ( \26438_26740 , RIfcede78_7729, \8893_9192 );
and \U$17620 ( \26439_26741 , RIe1fa370_4224, \8895_9194 );
and \U$17621 ( \26440_26742 , RIfcd4c48_7443, \8897_9196 );
and \U$17622 ( \26441_26743 , RIfce1dd0_7592, \8899_9198 );
and \U$17623 ( \26442_26744 , RIfcbf960_7202, \8901_9200 );
and \U$17624 ( \26443_26745 , RIe1f58e8_4171, \8903_9202 );
and \U$17625 ( \26444_26746 , RIfcbfc30_7204, \8905_9204 );
and \U$17626 ( \26445_26747 , RIfc78380_6390, \8907_9206 );
and \U$17627 ( \26446_26748 , RIfc93770_6700, \8909_9208 );
and \U$17628 ( \26447_26749 , RIe1f35c0_4146, \8911_9210 );
and \U$17629 ( \26448_26750 , RIfcb1f68_7047, \8913_9212 );
and \U$17630 ( \26449_26751 , RIfce1b00_7590, \8915_9214 );
and \U$17631 ( \26450_26752 , RIfc93a40_6702, \8917_9216 );
and \U$17632 ( \26451_26753 , RIe1ee2c8_4087, \8919_9218 );
and \U$17633 ( \26452_26754 , RIe1ebb68_4059, \8921_9220 );
and \U$17634 ( \26453_26755 , RIe1e8e68_4027, \8923_9222 );
and \U$17635 ( \26454_26756 , RIe1e6168_3995, \8925_9224 );
and \U$17636 ( \26455_26757 , RIe1e3468_3963, \8927_9226 );
and \U$17637 ( \26456_26758 , RIe1e0768_3931, \8929_9228 );
and \U$17638 ( \26457_26759 , RIe1dda68_3899, \8931_9230 );
and \U$17639 ( \26458_26760 , RIe1dad68_3867, \8933_9232 );
and \U$17640 ( \26459_26761 , RIe1d8068_3835, \8935_9234 );
and \U$17641 ( \26460_26762 , RIe1d2668_3771, \8937_9236 );
and \U$17642 ( \26461_26763 , RIe1cf968_3739, \8939_9238 );
and \U$17643 ( \26462_26764 , RIe1ccc68_3707, \8941_9240 );
and \U$17644 ( \26463_26765 , RIe1c9f68_3675, \8943_9242 );
and \U$17645 ( \26464_26766 , RIe1c7268_3643, \8945_9244 );
and \U$17646 ( \26465_26767 , RIe1c4568_3611, \8947_9246 );
and \U$17647 ( \26466_26768 , RIe1c1868_3579, \8949_9248 );
and \U$17648 ( \26467_26769 , RIe1beb68_3547, \8951_9250 );
and \U$17649 ( \26468_26770 , RIfcdec98_7557, \8953_9252 );
and \U$17650 ( \26469_26771 , RIfc94148_6707, \8955_9254 );
and \U$17651 ( \26470_26772 , RIe1b95a0_3486, \8957_9256 );
and \U$17652 ( \26471_26773 , RIe1b7548_3463, \8959_9258 );
and \U$17653 ( \26472_26774 , RIfcd12a0_7402, \8961_9260 );
and \U$17654 ( \26473_26775 , RIfceabd8_7693, \8963_9262 );
and \U$17655 ( \26474_26776 , RIe1b5388_3439, \8965_9264 );
and \U$17656 ( \26475_26777 , RIe1b3fd8_3425, \8967_9266 );
and \U$17657 ( \26476_26778 , RIfc94850_6712, \8969_9268 );
and \U$17658 ( \26477_26779 , RIfcd7c18_7477, \8971_9270 );
and \U$17659 ( \26478_26780 , RIe1b27f0_3408, \8973_9272 );
and \U$17660 ( \26479_26781 , RIe1b0d38_3389, \8975_9274 );
and \U$17661 ( \26480_26782 , RIfc76a30_6372, \8977_9276 );
and \U$17662 ( \26481_26783 , RIfce2640_7598, \8979_9278 );
and \U$17663 ( \26482_26784 , RIe1ac6e8_3339, \8981_9280 );
and \U$17664 ( \26483_26785 , RIe1ab068_3323, \8983_9282 );
and \U$17665 ( \26484_26786 , RIe1a8ea8_3299, \8985_9284 );
and \U$17666 ( \26485_26787 , RIe1a61a8_3267, \8987_9286 );
and \U$17667 ( \26486_26788 , RIe1a34a8_3235, \8989_9288 );
and \U$17668 ( \26487_26789 , RIe1a07a8_3203, \8991_9290 );
and \U$17669 ( \26488_26790 , RIe18cca8_2979, \8993_9292 );
and \U$17670 ( \26489_26791 , RIe1791a8_2755, \8995_9294 );
and \U$17671 ( \26490_26792 , RIe226b00_4730, \8997_9296 );
and \U$17672 ( \26491_26793 , RIe21b700_4602, \8999_9298 );
and \U$17673 ( \26492_26794 , RIe204f00_4346, \9001_9300 );
and \U$17674 ( \26493_26795 , RIe1fef60_4278, \9003_9302 );
and \U$17675 ( \26494_26796 , RIe1f8318_4201, \9005_9304 );
and \U$17676 ( \26495_26797 , RIe1f0e60_4118, \9007_9306 );
and \U$17677 ( \26496_26798 , RIe1d5368_3803, \9009_9308 );
and \U$17678 ( \26497_26799 , RIe1bbe68_3515, \9011_9310 );
and \U$17679 ( \26498_26800 , RIe1aece0_3366, \9013_9312 );
and \U$17680 ( \26499_26801 , RIe171318_2665, \9015_9314 );
or \U$17681 ( \26500_26802 , \26436_26738 , \26437_26739 , \26438_26740 , \26439_26741 , \26440_26742 , \26441_26743 , \26442_26744 , \26443_26745 , \26444_26746 , \26445_26747 , \26446_26748 , \26447_26749 , \26448_26750 , \26449_26751 , \26450_26752 , \26451_26753 , \26452_26754 , \26453_26755 , \26454_26756 , \26455_26757 , \26456_26758 , \26457_26759 , \26458_26760 , \26459_26761 , \26460_26762 , \26461_26763 , \26462_26764 , \26463_26765 , \26464_26766 , \26465_26767 , \26466_26768 , \26467_26769 , \26468_26770 , \26469_26771 , \26470_26772 , \26471_26773 , \26472_26774 , \26473_26775 , \26474_26776 , \26475_26777 , \26476_26778 , \26477_26779 , \26478_26780 , \26479_26781 , \26480_26782 , \26481_26783 , \26482_26784 , \26483_26785 , \26484_26786 , \26485_26787 , \26486_26788 , \26487_26789 , \26488_26790 , \26489_26791 , \26490_26792 , \26491_26793 , \26492_26794 , \26493_26795 , \26494_26796 , \26495_26797 , \26496_26798 , \26497_26799 , \26498_26800 , \26499_26801 );
or \U$17682 ( \26501_26803 , \26435_26737 , \26500_26802 );
_DC \g5e36/U$1 ( \26502 , \26501_26803 , \9024_9323 );
xor g5e37_GF_PartitionCandidate( \26503_26805_nG5e37 , \26370 , \26502 );
buf \U$17683 ( \26504_26806 , \26503_26805_nG5e37 );
xor \U$17684 ( \26505_26807 , \26504_26806 , \25471_25770 );
and \U$17685 ( \26506_26808 , \10385_10687 , \26505_26807 );
xor \U$17686 ( \26507_26809 , \26238_26540 , \26506_26808 );
and \U$17687 ( \26508_26810 , \19259_19558 , \15037_15336 );
and \U$17688 ( \26509_26811 , \20242_20544 , \14661_14963 );
nor \U$17689 ( \26510_26812 , \26508_26810 , \26509_26811 );
xnor \U$17690 ( \26511_26813 , \26510_26812 , \15043_15342 );
and \U$17691 ( \26512_26814 , \15022_15321 , \19235_19534 );
and \U$17692 ( \26513_26815 , \15965_16267 , \18743_19045 );
nor \U$17693 ( \26514_26816 , \26512_26814 , \26513_26815 );
xnor \U$17694 ( \26515_26817 , \26514_26816 , \19241_19540 );
xor \U$17695 ( \26516_26818 , \26511_26813 , \26515_26817 );
and \U$17696 ( \26517_26819 , \13725_14024 , \20706_21005 );
and \U$17697 ( \26518_26820 , \14648_14950 , \20255_20557 );
nor \U$17698 ( \26519_26821 , \26517_26819 , \26518_26820 );
xnor \U$17699 ( \26520_26822 , \26519_26821 , \20712_21011 );
xor \U$17700 ( \26521_26823 , \26516_26818 , \26520_26822 );
xor \U$17701 ( \26522_26824 , \26507_26809 , \26521_26823 );
and \U$17702 ( \26523_26825 , \25516_25815 , \10681_10983 );
_DC \g65bf/U$1 ( \26524 , \26369_26671 , \9298_9597 );
_DC \g65c0/U$1 ( \26525 , \26501_26803 , \9024_9323 );
and g65c1_GF_PartitionCandidate( \26526_26828_nG65c1 , \26524 , \26525 );
buf \U$17703 ( \26527_26829 , \26526_26828_nG65c1 );
and \U$17704 ( \26528_26830 , \26527_26829 , \10389_10691 );
nor \U$17705 ( \26529_26831 , \26523_26825 , \26528_26830 );
xnor \U$17706 ( \26530_26832 , \26529_26831 , \10678_10980 );
and \U$17707 ( \26531_26833 , \12470_12769 , \22243_22542 );
and \U$17708 ( \26532_26834 , \13377_13679 , \21801_22103 );
nor \U$17709 ( \26533_26835 , \26531_26833 , \26532_26834 );
xnor \U$17710 ( \26534_26836 , \26533_26835 , \22249_22548 );
xor \U$17711 ( \26535_26837 , \26530_26832 , \26534_26836 );
and \U$17712 ( \26536_26838 , \11287_11586 , \23839_24138 );
and \U$17713 ( \26537_26839 , \12146_12448 , \23328_23630 );
nor \U$17714 ( \26538_26840 , \26536_26838 , \26537_26839 );
xnor \U$17715 ( \26539_26841 , \26538_26840 , \23845_24144 );
xor \U$17716 ( \26540_26842 , \26535_26837 , \26539_26841 );
xor \U$17717 ( \26541_26843 , \26522_26824 , \26540_26842 );
xor \U$17718 ( \26542_26844 , \26229_26531 , \26541_26843 );
xor \U$17719 ( \26543_26845 , \26200_26502 , \26542_26844 );
and \U$17720 ( \26544_26846 , \25185_25484 , \25199_25498 );
and \U$17721 ( \26545_26847 , \25199_25498 , \25486_25785 );
and \U$17722 ( \26546_26848 , \25185_25484 , \25486_25785 );
or \U$17723 ( \26547_26849 , \26544_26846 , \26545_26847 , \26546_26848 );
and \U$17724 ( \26548_26850 , \25492_25791 , \25506_25805 );
and \U$17725 ( \26549_26851 , \25506_25805 , \25548_25847 );
and \U$17726 ( \26550_26852 , \25492_25791 , \25548_25847 );
or \U$17727 ( \26551_26853 , \26548_26850 , \26549_26851 , \26550_26852 );
xor \U$17728 ( \26552_26854 , \26547_26849 , \26551_26853 );
and \U$17729 ( \26553_26855 , \25496_25795 , \25500_25799 );
and \U$17730 ( \26554_26856 , \25500_25799 , \25505_25804 );
and \U$17731 ( \26555_26857 , \25496_25795 , \25505_25804 );
or \U$17732 ( \26556_26858 , \26553_26855 , \26554_26856 , \26555_26857 );
and \U$17733 ( \26557_26859 , \25476_25775 , \25480_25779 );
and \U$17734 ( \26558_26860 , \25480_25779 , \25485_25784 );
and \U$17735 ( \26559_26861 , \25476_25775 , \25485_25784 );
or \U$17736 ( \26560_26862 , \26557_26859 , \26558_26860 , \26559_26861 );
xor \U$17737 ( \26561_26863 , \26556_26858 , \26560_26862 );
and \U$17738 ( \26562_26864 , \25537_25836 , \25541_25840 );
and \U$17739 ( \26563_26865 , \25541_25840 , \25546_25845 );
and \U$17740 ( \26564_26866 , \25537_25836 , \25546_25845 );
or \U$17741 ( \26565_26867 , \26562_26864 , \26563_26865 , \26564_26866 );
and \U$17742 ( \26566_26868 , \25204_25503 , \25475_25774 );
xor \U$17743 ( \26567_26869 , \26565_26867 , \26566_26868 );
and \U$17744 ( \26568_26870 , \16353_16655 , \17791_18090 );
and \U$17745 ( \26569_26871 , \17325_17627 , \17353_17655 );
nor \U$17746 ( \26570_26872 , \26568_26870 , \26569_26871 );
xnor \U$17747 ( \26571_26873 , \26570_26872 , \17747_18046 );
xor \U$17748 ( \26572_26874 , \26567_26869 , \26571_26873 );
xor \U$17749 ( \26573_26875 , \26561_26863 , \26572_26874 );
xor \U$17750 ( \26574_26876 , \26552_26854 , \26573_26875 );
xor \U$17751 ( \26575_26877 , \26543_26845 , \26574_26876 );
and \U$17752 ( \26576_26878 , \25172_25471 , \25176_25475 );
and \U$17753 ( \26577_26879 , \25176_25475 , \25550_25849 );
and \U$17754 ( \26578_26880 , \25172_25471 , \25550_25849 );
or \U$17755 ( \26579_26881 , \26576_26878 , \26577_26879 , \26578_26880 );
xor \U$17756 ( \26580_26882 , \26575_26877 , \26579_26881 );
and \U$17757 ( \26581_26883 , \25551_25850 , \25555_25854 );
and \U$17758 ( \26582_26884 , \25556_25855 , \25559_25858 );
or \U$17759 ( \26583_26885 , \26581_26883 , \26582_26884 );
xor \U$17760 ( \26584_26886 , \26580_26882 , \26583_26885 );
buf g9bc6_GF_PartitionCandidate( \26585_26887_nG9bc6 , \26584_26886 );
and \U$17761 ( \26586_26888 , \10402_10704 , \26585_26887_nG9bc6 );
or \U$17762 ( \26587_26889 , \26196_26498 , \26586_26888 );
xor \U$17763 ( \26588_26890 , \10399_10703 , \26587_26889 );
buf \U$17764 ( \26589_26891 , \26588_26890 );
buf \U$17766 ( \26590_26892 , \26589_26891 );
xor \U$17767 ( \26591_26893 , \26195_26497 , \26590_26892 );
buf \U$17768 ( \26592_26894 , \26591_26893 );
xor \U$17769 ( \26593_26895 , \26146_26448 , \26592_26894 );
and \U$17770 ( \26594_26896 , \25083_25382 , \25114_25413 );
and \U$17771 ( \26595_26897 , \25083_25382 , \25121_25420 );
and \U$17772 ( \26596_26898 , \25114_25413 , \25121_25420 );
or \U$17773 ( \26597_26899 , \26594_26896 , \26595_26897 , \26596_26898 );
buf \U$17774 ( \26598_26900 , \26597_26899 );
xor \U$17775 ( \26599_26901 , \26593_26895 , \26598_26900 );
buf \U$17776 ( \26600_26902 , \26599_26901 );
and \U$17777 ( \26601_26903 , \25134_25433 , \25139_25438 );
and \U$17778 ( \26602_26904 , \25134_25433 , \25146_25445 );
and \U$17779 ( \26603_26905 , \25139_25438 , \25146_25445 );
or \U$17780 ( \26604_26906 , \26601_26903 , \26602_26904 , \26603_26905 );
buf \U$17781 ( \26605_26907 , \26604_26906 );
and \U$17782 ( \26606_26908 , \25088_25387 , \25105_25404 );
and \U$17783 ( \26607_26909 , \25088_25387 , \25112_25411 );
and \U$17784 ( \26608_26910 , \25105_25404 , \25112_25411 );
or \U$17785 ( \26609_26911 , \26606_26908 , \26607_26909 , \26608_26910 );
buf \U$17786 ( \26610_26912 , \26609_26911 );
and \U$17787 ( \26611_26913 , \12183_12157 , \22330_22629_nG9bd5 );
and \U$17788 ( \26612_26914 , \11855_12154 , \23394_23696_nG9bd2 );
or \U$17789 ( \26613_26915 , \26611_26913 , \26612_26914 );
xor \U$17790 ( \26614_26916 , \11854_12153 , \26613_26915 );
buf \U$17791 ( \26615_26917 , \26614_26916 );
buf \U$17793 ( \26616_26918 , \26615_26917 );
xor \U$17794 ( \26617_26919 , \26610_26912 , \26616_26918 );
and \U$17795 ( \26618_26920 , \10996_10421 , \23927_24226_nG9bcf );
and \U$17796 ( \26619_26921 , \10119_10418 , \24996_25298_nG9bcc );
or \U$17797 ( \26620_26922 , \26618_26920 , \26619_26921 );
xor \U$17798 ( \26621_26923 , \10118_10417 , \26620_26922 );
buf \U$17799 ( \26622_26924 , \26621_26923 );
buf \U$17801 ( \26623_26925 , \26622_26924 );
xor \U$17802 ( \26624_26926 , \26617_26919 , \26623_26925 );
buf \U$17803 ( \26625_26927 , \26624_26926 );
xor \U$17804 ( \26626_26928 , \26605_26907 , \26625_26927 );
and \U$17805 ( \26627_26929 , \25090_25389 , \25096_25395 );
and \U$17806 ( \26628_26930 , \25090_25389 , \25103_25402 );
and \U$17807 ( \26629_26931 , \25096_25395 , \25103_25402 );
or \U$17808 ( \26630_26932 , \26627_26929 , \26628_26930 , \26629_26931 );
buf \U$17809 ( \26631_26933 , \26630_26932 );
and \U$17810 ( \26632_26934 , \25033_25335 , \25039_25341 );
buf \U$17811 ( \26633_26935 , \26632_26934 );
and \U$17812 ( \26634_26936 , \21908_21658 , \12502_12801_nG9bff );
and \U$17813 ( \26635_26937 , \21356_21655 , \13403_13705_nG9bfc );
or \U$17814 ( \26636_26938 , \26634_26936 , \26635_26937 );
xor \U$17815 ( \26637_26939 , \21355_21654 , \26636_26938 );
buf \U$17816 ( \26638_26940 , \26637_26939 );
buf \U$17818 ( \26639_26941 , \26638_26940 );
xor \U$17819 ( \26640_26942 , \26633_26935 , \26639_26941 );
and \U$17820 ( \26641_26943 , \20353_20155 , \13771_14070_nG9bf9 );
and \U$17821 ( \26642_26944 , \19853_20152 , \14682_14984_nG9bf6 );
or \U$17822 ( \26643_26945 , \26641_26943 , \26642_26944 );
xor \U$17823 ( \26644_26946 , \19852_20151 , \26643_26945 );
buf \U$17824 ( \26645_26947 , \26644_26946 );
buf \U$17826 ( \26646_26948 , \26645_26947 );
xor \U$17827 ( \26647_26949 , \26640_26942 , \26646_26948 );
buf \U$17828 ( \26648_26950 , \26647_26949 );
xor \U$17829 ( \26649_26951 , \26631_26933 , \26648_26950 );
and \U$17830 ( \26650_26952 , \17437_17297 , \16378_16680_nG9bed );
and \U$17831 ( \26651_26953 , \16995_17294 , \17363_17665_nG9bea );
or \U$17832 ( \26652_26954 , \26650_26952 , \26651_26953 );
xor \U$17833 ( \26653_26955 , \16994_17293 , \26652_26954 );
buf \U$17834 ( \26654_26956 , \26653_26955 );
buf \U$17836 ( \26655_26957 , \26654_26956 );
xor \U$17837 ( \26656_26958 , \26649_26951 , \26655_26957 );
buf \U$17838 ( \26657_26959 , \26656_26958 );
and \U$17839 ( \26658_26960 , \25030_25332 , \25059_25358 );
and \U$17840 ( \26659_26961 , \25030_25332 , \25066_25365 );
and \U$17841 ( \26660_26962 , \25059_25358 , \25066_25365 );
or \U$17842 ( \26661_26963 , \26658_26960 , \26659_26961 , \26660_26962 );
buf \U$17843 ( \26662_26964 , \26661_26963 );
xor \U$17844 ( \26663_26965 , \26657_26959 , \26662_26964 );
and \U$17845 ( \26664_26966 , \13431_13370 , \20787_21086_nG9bdb );
and \U$17846 ( \26665_26967 , \13068_13367 , \21827_22129_nG9bd8 );
or \U$17847 ( \26666_26968 , \26664_26966 , \26665_26967 );
xor \U$17848 ( \26667_26969 , \13067_13366 , \26666_26968 );
buf \U$17849 ( \26668_26970 , \26667_26969 );
buf \U$17851 ( \26669_26971 , \26668_26970 );
xor \U$17852 ( \26670_26972 , \26663_26965 , \26669_26971 );
buf \U$17853 ( \26671_26973 , \26670_26972 );
xor \U$17854 ( \26672_26974 , \26626_26928 , \26671_26973 );
buf \U$17855 ( \26673_26975 , \26672_26974 );
xor \U$17856 ( \26674_26976 , \26600_26902 , \26673_26975 );
and \U$17857 ( \26675_26977 , \25123_25422 , \25128_25427 );
and \U$17858 ( \26676_26978 , \25123_25422 , \25148_25447 );
and \U$17859 ( \26677_26979 , \25128_25427 , \25148_25447 );
or \U$17860 ( \26678_26980 , \26675_26977 , \26676_26978 , \26677_26979 );
buf \U$17861 ( \26679_26981 , \26678_26980 );
xor \U$17862 ( \26680_26982 , \26674_26976 , \26679_26981 );
and \U$17863 ( \26681_26983 , \26136_26438 , \26680_26982 );
and \U$17864 ( \26682_26984 , \26140_26442 , \26680_26982 );
or \U$17865 ( \26683_26985 , \26141_26443 , \26681_26983 , \26682_26984 );
and \U$17866 ( \26684_26986 , \25575_25874 , \25579_25878 );
and \U$17867 ( \26685_26987 , \25575_25874 , \26135_26437 );
and \U$17868 ( \26686_26988 , \25579_25878 , \26135_26437 );
or \U$17869 ( \26687_26989 , \26684_26986 , \26685_26987 , \26686_26988 );
xor \U$17870 ( \26688_26990 , \26683_26985 , \26687_26989 );
and \U$17871 ( \26689_26991 , \26600_26902 , \26673_26975 );
and \U$17872 ( \26690_26992 , \26600_26902 , \26679_26981 );
and \U$17873 ( \26691_26993 , \26673_26975 , \26679_26981 );
or \U$17874 ( \26692_26994 , \26689_26991 , \26690_26992 , \26691_26993 );
xor \U$17875 ( \26693_26995 , \26688_26990 , \26692_26994 );
and \U$17876 ( \26694_26996 , \26605_26907 , \26625_26927 );
and \U$17877 ( \26695_26997 , \26605_26907 , \26671_26973 );
and \U$17878 ( \26696_26998 , \26625_26927 , \26671_26973 );
or \U$17879 ( \26697_26999 , \26694_26996 , \26695_26997 , \26696_26998 );
buf \U$17880 ( \26698_27000 , \26697_26999 );
and \U$17881 ( \26699_27001 , \26657_26959 , \26662_26964 );
and \U$17882 ( \26700_27002 , \26657_26959 , \26669_26971 );
and \U$17883 ( \26701_27003 , \26662_26964 , \26669_26971 );
or \U$17884 ( \26702_27004 , \26699_27001 , \26700_27002 , \26701_27003 );
buf \U$17885 ( \26703_27005 , \26702_27004 );
and \U$17886 ( \26704_27006 , \10996_10421 , \24996_25298_nG9bcc );
and \U$17887 ( \26705_27007 , \10119_10418 , \25561_25860_nG9bc9 );
or \U$17888 ( \26706_27008 , \26704_27006 , \26705_27007 );
xor \U$17889 ( \26707_27009 , \10118_10417 , \26706_27008 );
buf \U$17890 ( \26708_27010 , \26707_27009 );
buf \U$17892 ( \26709_27011 , \26708_27010 );
xor \U$17893 ( \26710_27012 , \26703_27005 , \26709_27011 );
and \U$17894 ( \26711_27013 , \10411_10707 , \26585_26887_nG9bc6 );
and \U$17895 ( \26712_27014 , \26547_26849 , \26551_26853 );
and \U$17896 ( \26713_27015 , \26551_26853 , \26573_26875 );
and \U$17897 ( \26714_27016 , \26547_26849 , \26573_26875 );
or \U$17898 ( \26715_27017 , \26712_27014 , \26713_27015 , \26714_27016 );
and \U$17899 ( \26716_27018 , \26208_26510 , \26212_26514 );
and \U$17900 ( \26717_27019 , \26212_26514 , \26227_26529 );
and \U$17901 ( \26718_27020 , \26208_26510 , \26227_26529 );
or \U$17902 ( \26719_27021 , \26716_27018 , \26717_27019 , \26718_27020 );
and \U$17903 ( \26720_27022 , \24970_25272 , \11275_11574 );
and \U$17904 ( \26721_27023 , \25516_25815 , \10976_11278 );
nor \U$17905 ( \26722_27024 , \26720_27022 , \26721_27023 );
xnor \U$17906 ( \26723_27025 , \26722_27024 , \11281_11580 );
not \U$17907 ( \26724_27026 , \26506_26808 );
and \U$17908 ( \26725_27027 , RIdec5978_712, \9034_9333 );
and \U$17909 ( \26726_27028 , RIdec2c78_680, \9036_9335 );
and \U$17910 ( \26727_27029 , RIfc8aad0_6600, \9038_9337 );
and \U$17911 ( \26728_27030 , RIdebff78_648, \9040_9339 );
and \U$17912 ( \26729_27031 , RIfc8ac38_6601, \9042_9341 );
and \U$17913 ( \26730_27032 , RIdebd278_616, \9044_9343 );
and \U$17914 ( \26731_27033 , RIdeba578_584, \9046_9345 );
and \U$17915 ( \26732_27034 , RIdeb7878_552, \9048_9347 );
and \U$17916 ( \26733_27035 , RIfc40e80_5764, \9050_9349 );
and \U$17917 ( \26734_27036 , RIdeb1e78_488, \9052_9351 );
and \U$17918 ( \26735_27037 , RIfcdaeb8_7513, \9054_9353 );
and \U$17919 ( \26736_27038 , RIdeaf178_456, \9056_9355 );
and \U$17920 ( \26737_27039 , RIee1dbf0_4797, \9058_9357 );
and \U$17921 ( \26738_27040 , RIdeab140_424, \9060_9359 );
and \U$17922 ( \26739_27041 , RIdea4840_392, \9062_9361 );
and \U$17923 ( \26740_27042 , RIde9df40_360, \9064_9363 );
and \U$17924 ( \26741_27043 , RIfc8b070_6604, \9066_9365 );
and \U$17925 ( \26742_27044 , RIfcc38a8_7247, \9068_9367 );
and \U$17926 ( \26743_27045 , RIfc807b0_6484, \9070_9369 );
and \U$17927 ( \26744_27046 , RIfcbb8b0_7156, \9072_9371 );
and \U$17928 ( \26745_27047 , RIde91a60_300, \9074_9373 );
and \U$17929 ( \26746_27048 , RIde8e298_283, \9076_9375 );
and \U$17930 ( \26747_27049 , RIde8a440_264, \9078_9377 );
and \U$17931 ( \26748_27050 , RIde862a0_244, \9080_9379 );
and \U$17932 ( \26749_27051 , RIde82100_224, \9082_9381 );
and \U$17933 ( \26750_27052 , RIfcbbb80_7158, \9084_9383 );
and \U$17934 ( \26751_27053 , RIfc8c150_6616, \9086_9385 );
and \U$17935 ( \26752_27054 , RIfcbbfb8_7161, \9088_9387 );
and \U$17936 ( \26753_27055 , RIfc54458_5981, \9090_9389 );
and \U$17937 ( \26754_27056 , RIe16bbe8_2603, \9092_9391 );
and \U$17938 ( \26755_27057 , RIfc8c2b8_6617, \9094_9393 );
and \U$17939 ( \26756_27058 , RIe168240_2562, \9096_9395 );
and \U$17940 ( \26757_27059 , RIe165978_2533, \9098_9397 );
and \U$17941 ( \26758_27060 , RIe162c78_2501, \9100_9399 );
and \U$17942 ( \26759_27061 , RIee37960_5091, \9102_9401 );
and \U$17943 ( \26760_27062 , RIe15ff78_2469, \9104_9403 );
and \U$17944 ( \26761_27063 , RIfcd6b38_7465, \9106_9405 );
and \U$17945 ( \26762_27064 , RIe15d278_2437, \9108_9407 );
and \U$17946 ( \26763_27065 , RIe157878_2373, \9110_9409 );
and \U$17947 ( \26764_27066 , RIe154b78_2341, \9112_9411 );
and \U$17948 ( \26765_27067 , RIfc8e5e0_6642, \9114_9413 );
and \U$17949 ( \26766_27068 , RIe151e78_2309, \9116_9415 );
and \U$17950 ( \26767_27069 , RIfcb4290_7072, \9118_9417 );
and \U$17951 ( \26768_27070 , RIe14f178_2277, \9120_9419 );
and \U$17952 ( \26769_27071 , RIfc56ff0_6012, \9122_9421 );
and \U$17953 ( \26770_27072 , RIe14c478_2245, \9124_9423 );
and \U$17954 ( \26771_27073 , RIe149778_2213, \9126_9425 );
and \U$17955 ( \26772_27074 , RIe146a78_2181, \9128_9427 );
and \U$17956 ( \26773_27075 , RIee346c0_5055, \9130_9429 );
and \U$17957 ( \26774_27076 , RIee335e0_5043, \9132_9431 );
and \U$17958 ( \26775_27077 , RIee32398_5030, \9134_9433 );
and \U$17959 ( \26776_27078 , RIee31420_5019, \9136_9435 );
and \U$17960 ( \26777_27079 , RIe141348_2119, \9138_9437 );
and \U$17961 ( \26778_27080 , RIe13f020_2094, \9140_9439 );
and \U$17962 ( \26779_27081 , RIfec16f8_8321, \9142_9441 );
and \U$17963 ( \26780_27082 , RIdf3a930_2043, \9144_9443 );
and \U$17964 ( \26781_27083 , RIfce3e28_7615, \9146_9445 );
and \U$17965 ( \26782_27084 , RIfc56780_6006, \9148_9447 );
and \U$17966 ( \26783_27085 , RIfcb4128_7071, \9150_9449 );
and \U$17967 ( \26784_27086 , RIfce2eb0_7604, \9152_9451 );
and \U$17968 ( \26785_27087 , RIdf35d40_1989, \9154_9453 );
and \U$17969 ( \26786_27088 , RIfe88218_7893, \9156_9455 );
and \U$17970 ( \26787_27089 , RIdf316f0_1939, \9158_9457 );
and \U$17971 ( \26788_27090 , RIdf2f698_1916, \9160_9459 );
or \U$17972 ( \26789_27091 , \26725_27027 , \26726_27028 , \26727_27029 , \26728_27030 , \26729_27031 , \26730_27032 , \26731_27033 , \26732_27034 , \26733_27035 , \26734_27036 , \26735_27037 , \26736_27038 , \26737_27039 , \26738_27040 , \26739_27041 , \26740_27042 , \26741_27043 , \26742_27044 , \26743_27045 , \26744_27046 , \26745_27047 , \26746_27048 , \26747_27049 , \26748_27050 , \26749_27051 , \26750_27052 , \26751_27053 , \26752_27054 , \26753_27055 , \26754_27056 , \26755_27057 , \26756_27058 , \26757_27059 , \26758_27060 , \26759_27061 , \26760_27062 , \26761_27063 , \26762_27064 , \26763_27065 , \26764_27066 , \26765_27067 , \26766_27068 , \26767_27069 , \26768_27070 , \26769_27071 , \26770_27072 , \26771_27073 , \26772_27074 , \26773_27075 , \26774_27076 , \26775_27077 , \26776_27078 , \26777_27079 , \26778_27080 , \26779_27081 , \26780_27082 , \26781_27083 , \26782_27084 , \26783_27085 , \26784_27086 , \26785_27087 , \26786_27088 , \26787_27089 , \26788_27090 );
and \U$17973 ( \26790_27092 , RIfc7f9a0_6474, \9163_9462 );
and \U$17974 ( \26791_27093 , RIfce4260_7618, \9165_9464 );
and \U$17975 ( \26792_27094 , RIfcd62c8_7459, \9167_9466 );
and \U$17976 ( \26793_27095 , RIfce9990_7680, \9169_9468 );
and \U$17977 ( \26794_27096 , RIdf2a670_1859, \9171_9470 );
and \U$17978 ( \26795_27097 , RIdf284b0_1835, \9173_9472 );
and \U$17979 ( \26796_27098 , RIdf26728_1814, \9175_9474 );
and \U$17980 ( \26797_27099 , RIdf24c70_1795, \9177_9476 );
and \U$17981 ( \26798_27100 , RIfc7ecf8_6465, \9179_9478 );
and \U$17982 ( \26799_27101 , RIfcc31a0_7242, \9181_9480 );
and \U$17983 ( \26800_27102 , RIfc99008_6763, \9183_9482 );
and \U$17984 ( \26801_27103 , RIfc46e98_5829, \9185_9484 );
and \U$17985 ( \26802_27104 , RIfce2a78_7601, \9187_9486 );
and \U$17986 ( \26803_27105 , RIdf1fdb0_1739, \9189_9488 );
and \U$17987 ( \26804_27106 , RIfcc6e18_7285, \9191_9490 );
and \U$17988 ( \26805_27107 , RIdf19708_1666, \9193_9492 );
and \U$17989 ( \26806_27108 , RIdf17548_1642, \9195_9494 );
and \U$17990 ( \26807_27109 , RIdf14848_1610, \9197_9496 );
and \U$17991 ( \26808_27110 , RIdf11b48_1578, \9199_9498 );
and \U$17992 ( \26809_27111 , RIdf0ee48_1546, \9201_9500 );
and \U$17993 ( \26810_27112 , RIdf0c148_1514, \9203_9502 );
and \U$17994 ( \26811_27113 , RIdf09448_1482, \9205_9504 );
and \U$17995 ( \26812_27114 , RIdf06748_1450, \9207_9506 );
and \U$17996 ( \26813_27115 , RIdf03a48_1418, \9209_9508 );
and \U$17997 ( \26814_27116 , RIdefe048_1354, \9211_9510 );
and \U$17998 ( \26815_27117 , RIdefb348_1322, \9213_9512 );
and \U$17999 ( \26816_27118 , RIdef8648_1290, \9215_9514 );
and \U$18000 ( \26817_27119 , RIdef5948_1258, \9217_9516 );
and \U$18001 ( \26818_27120 , RIdef2c48_1226, \9219_9518 );
and \U$18002 ( \26819_27121 , RIdeeff48_1194, \9221_9520 );
and \U$18003 ( \26820_27122 , RIdeed248_1162, \9223_9522 );
and \U$18004 ( \26821_27123 , RIdeea548_1130, \9225_9524 );
and \U$18005 ( \26822_27124 , RIfcd9130_7492, \9227_9526 );
and \U$18006 ( \26823_27125 , RIfc7cb38_6441, \9229_9528 );
and \U$18007 ( \26824_27126 , RIfc97af0_6748, \9231_9530 );
and \U$18008 ( \26825_27127 , RIfcb3e58_7069, \9233_9532 );
and \U$18009 ( \26826_27128 , RIdee4e18_1068, \9235_9534 );
and \U$18010 ( \26827_27129 , RIdee3090_1047, \9237_9536 );
and \U$18011 ( \26828_27130 , RIdee0ed0_1023, \9239_9538 );
and \U$18012 ( \26829_27131 , RIfe88380_7894, \9241_9540 );
and \U$18013 ( \26830_27132 , RIfc97dc0_6750, \9243_9542 );
and \U$18014 ( \26831_27133 , RIfcc2930_7236, \9245_9544 );
and \U$18015 ( \26832_27134 , RIfcd9298_7493, \9247_9546 );
and \U$18016 ( \26833_27135 , RIfc7c868_6439, \9249_9548 );
and \U$18017 ( \26834_27136 , RIded9ce8_942, \9251_9550 );
and \U$18018 ( \26835_27137 , RIded76f0_915, \9253_9552 );
and \U$18019 ( \26836_27138 , RIded5968_894, \9255_9554 );
and \U$18020 ( \26837_27139 , RIded3370_867, \9257_9556 );
and \U$18021 ( \26838_27140 , RIded0d78_840, \9259_9558 );
and \U$18022 ( \26839_27141 , RIdece078_808, \9261_9560 );
and \U$18023 ( \26840_27142 , RIdecb378_776, \9263_9562 );
and \U$18024 ( \26841_27143 , RIdec8678_744, \9265_9564 );
and \U$18025 ( \26842_27144 , RIdeb4b78_520, \9267_9566 );
and \U$18026 ( \26843_27145 , RIde97640_328, \9269_9568 );
and \U$18027 ( \26844_27146 , RIe16e780_2634, \9271_9570 );
and \U$18028 ( \26845_27147 , RIe15a578_2405, \9273_9572 );
and \U$18029 ( \26846_27148 , RIe143d78_2149, \9275_9574 );
and \U$18030 ( \26847_27149 , RIdf38770_2019, \9277_9576 );
and \U$18031 ( \26848_27150 , RIdf2cdd0_1887, \9279_9578 );
and \U$18032 ( \26849_27151 , RIdf1d650_1711, \9281_9580 );
and \U$18033 ( \26850_27152 , RIdf00d48_1386, \9283_9582 );
and \U$18034 ( \26851_27153 , RIdee7848_1098, \9285_9584 );
and \U$18035 ( \26852_27154 , RIdedc5b0_971, \9287_9586 );
and \U$18036 ( \26853_27155 , RIde7d588_201, \9289_9588 );
or \U$18037 ( \26854_27156 , \26790_27092 , \26791_27093 , \26792_27094 , \26793_27095 , \26794_27096 , \26795_27097 , \26796_27098 , \26797_27099 , \26798_27100 , \26799_27101 , \26800_27102 , \26801_27103 , \26802_27104 , \26803_27105 , \26804_27106 , \26805_27107 , \26806_27108 , \26807_27109 , \26808_27110 , \26809_27111 , \26810_27112 , \26811_27113 , \26812_27114 , \26813_27115 , \26814_27116 , \26815_27117 , \26816_27118 , \26817_27119 , \26818_27120 , \26819_27121 , \26820_27122 , \26821_27123 , \26822_27124 , \26823_27125 , \26824_27126 , \26825_27127 , \26826_27128 , \26827_27129 , \26828_27130 , \26829_27131 , \26830_27132 , \26831_27133 , \26832_27134 , \26833_27135 , \26834_27136 , \26835_27137 , \26836_27138 , \26837_27139 , \26838_27140 , \26839_27141 , \26840_27142 , \26841_27143 , \26842_27144 , \26843_27145 , \26844_27146 , \26845_27147 , \26846_27148 , \26847_27149 , \26848_27150 , \26849_27151 , \26850_27152 , \26851_27153 , \26852_27154 , \26853_27155 );
or \U$18038 ( \26855_27157 , \26789_27091 , \26854_27156 );
_DC \g5ebb/U$1 ( \26856 , \26855_27157 , \9298_9597 );
and \U$18039 ( \26857_27159 , RIe19dc10_3172, \8760_9059 );
and \U$18040 ( \26858_27160 , RIe19af10_3140, \8762_9061 );
and \U$18041 ( \26859_27161 , RIfec1590_8320, \8764_9063 );
and \U$18042 ( \26860_27162 , RIe198210_3108, \8766_9065 );
and \U$18043 ( \26861_27163 , RIfec1428_8319, \8768_9067 );
and \U$18044 ( \26862_27164 , RIe195510_3076, \8770_9069 );
and \U$18045 ( \26863_27165 , RIe192810_3044, \8772_9071 );
and \U$18046 ( \26864_27166 , RIe18fb10_3012, \8774_9073 );
and \U$18047 ( \26865_27167 , RIe18a110_2948, \8776_9075 );
and \U$18048 ( \26866_27168 , RIe187410_2916, \8778_9077 );
and \U$18049 ( \26867_27169 , RIfec12c0_8318, \8780_9079 );
and \U$18050 ( \26868_27170 , RIe184710_2884, \8782_9081 );
and \U$18051 ( \26869_27171 , RIfc88370_6572, \8784_9083 );
and \U$18052 ( \26870_27172 , RIe181a10_2852, \8786_9085 );
and \U$18053 ( \26871_27173 , RIe17ed10_2820, \8788_9087 );
and \U$18054 ( \26872_27174 , RIe17c010_2788, \8790_9089 );
and \U$18055 ( \26873_27175 , RIfc6ccb0_6260, \8792_9091 );
and \U$18056 ( \26874_27176 , RIfc5f858_6109, \8794_9093 );
and \U$18057 ( \26875_27177 , RIfca88f0_6940, \8796_9095 );
and \U$18058 ( \26876_27178 , RIe175f08_2719, \8798_9097 );
and \U$18059 ( \26877_27179 , RIfc81020_6490, \8800_9099 );
and \U$18060 ( \26878_27180 , RIfcc6008_7275, \8802_9101 );
and \U$18061 ( \26879_27181 , RIfc4ea58_5917, \8804_9103 );
and \U$18062 ( \26880_27182 , RIfc42140_5774, \8806_9105 );
and \U$18063 ( \26881_27183 , RIfca3b98_6885, \8808_9107 );
and \U$18064 ( \26882_27184 , RIfc5ac68_6055, \8810_9109 );
and \U$18065 ( \26883_27185 , RIfc984c8_6755, \8812_9111 );
and \U$18066 ( \26884_27186 , RIe173d48_2695, \8814_9113 );
and \U$18067 ( \26885_27187 , RIfc9b330_6788, \8816_9115 );
and \U$18068 ( \26886_27188 , RIf16f688_5727, \8818_9117 );
and \U$18069 ( \26887_27189 , RIfc42410_5776, \8820_9119 );
and \U$18070 ( \26888_27190 , RIfc5f588_6107, \8822_9121 );
and \U$18071 ( \26889_27191 , RIfe880b0_7892, \8824_9123 );
and \U$18072 ( \26890_27192 , RIe223f68_4699, \8826_9125 );
and \U$18073 ( \26891_27193 , RIf16bfb0_5688, \8828_9127 );
and \U$18074 ( \26892_27194 , RIe221268_4667, \8830_9129 );
and \U$18075 ( \26893_27195 , RIfc86cf0_6556, \8832_9131 );
and \U$18076 ( \26894_27196 , RIe21e568_4635, \8834_9133 );
and \U$18077 ( \26895_27197 , RIe218b68_4571, \8836_9135 );
and \U$18078 ( \26896_27198 , RIe215e68_4539, \8838_9137 );
and \U$18079 ( \26897_27199 , RIfe87de0_7890, \8840_9139 );
and \U$18080 ( \26898_27200 , RIe213168_4507, \8842_9141 );
and \U$18081 ( \26899_27201 , RIf1692b0_5656, \8844_9143 );
and \U$18082 ( \26900_27202 , RIe210468_4475, \8846_9145 );
and \U$18083 ( \26901_27203 , RIfcdf670_7564, \8848_9147 );
and \U$18084 ( \26902_27204 , RIe20d768_4443, \8850_9149 );
and \U$18085 ( \26903_27205 , RIe20aa68_4411, \8852_9151 );
and \U$18086 ( \26904_27206 , RIe207d68_4379, \8854_9153 );
and \U$18087 ( \26905_27207 , RIfca6460_6914, \8856_9155 );
and \U$18088 ( \26906_27208 , RIf1662e0_5622, \8858_9157 );
and \U$18089 ( \26907_27209 , RIe202908_4319, \8860_9159 );
and \U$18090 ( \26908_27210 , RIfe87b10_7888, \8862_9161 );
and \U$18091 ( \26909_27211 , RIfc58c10_6032, \8864_9163 );
and \U$18092 ( \26910_27212 , RIfc50ab0_5940, \8866_9165 );
and \U$18093 ( \26911_27213 , RIfccd790_7360, \8868_9167 );
and \U$18094 ( \26912_27214 , RIfccd1f0_7356, \8870_9169 );
and \U$18095 ( \26913_27215 , RIf160610_5556, \8872_9171 );
and \U$18096 ( \26914_27216 , RIf15e720_5534, \8874_9173 );
and \U$18097 ( \26915_27217 , RIfe87c78_7889, \8876_9175 );
and \U$18098 ( \26916_27218 , RIfe87f48_7891, \8878_9177 );
and \U$18099 ( \26917_27219 , RIfce7668_7655, \8880_9179 );
and \U$18100 ( \26918_27220 , RIfc86480_6550, \8882_9181 );
and \U$18101 ( \26919_27221 , RIfcd2218_7413, \8884_9183 );
and \U$18102 ( \26920_27222 , RIfcb01e0_7026, \8886_9185 );
or \U$18103 ( \26921_27223 , \26857_27159 , \26858_27160 , \26859_27161 , \26860_27162 , \26861_27163 , \26862_27164 , \26863_27165 , \26864_27166 , \26865_27167 , \26866_27168 , \26867_27169 , \26868_27170 , \26869_27171 , \26870_27172 , \26871_27173 , \26872_27174 , \26873_27175 , \26874_27176 , \26875_27177 , \26876_27178 , \26877_27179 , \26878_27180 , \26879_27181 , \26880_27182 , \26881_27183 , \26882_27184 , \26883_27185 , \26884_27186 , \26885_27187 , \26886_27188 , \26887_27189 , \26888_27190 , \26889_27191 , \26890_27192 , \26891_27193 , \26892_27194 , \26893_27195 , \26894_27196 , \26895_27197 , \26896_27198 , \26897_27199 , \26898_27200 , \26899_27201 , \26900_27202 , \26901_27203 , \26902_27204 , \26903_27205 , \26904_27206 , \26905_27207 , \26906_27208 , \26907_27209 , \26908_27210 , \26909_27211 , \26910_27212 , \26911_27213 , \26912_27214 , \26913_27215 , \26914_27216 , \26915_27217 , \26916_27218 , \26917_27219 , \26918_27220 , \26919_27221 , \26920_27222 );
and \U$18104 ( \26922_27224 , RIfc47b40_5838, \8889_9188 );
and \U$18105 ( \26923_27225 , RIfc84158_6525, \8891_9190 );
and \U$18106 ( \26924_27226 , RIfc4b920_5882, \8893_9192 );
and \U$18107 ( \26925_27227 , RIe1fa4d8_4225, \8895_9194 );
and \U$18108 ( \26926_27228 , RIfc4ba88_5883, \8897_9196 );
and \U$18109 ( \26927_27229 , RIfcb7530_7108, \8899_9198 );
and \U$18110 ( \26928_27230 , RIfcd58f0_7452, \8901_9200 );
and \U$18111 ( \26929_27231 , RIe1f5a50_4172, \8903_9202 );
and \U$18112 ( \26930_27232 , RIf153488_5407, \8905_9204 );
and \U$18113 ( \26931_27233 , RIf151ca0_5390, \8907_9206 );
and \U$18114 ( \26932_27234 , RIfc51e60_5954, \8909_9208 );
and \U$18115 ( \26933_27235 , RIe1f3728_4147, \8911_9210 );
and \U$18116 ( \26934_27236 , RIfc9aef8_6785, \8913_9212 );
and \U$18117 ( \26935_27237 , RIfcbaaa0_7146, \8915_9214 );
and \U$18118 ( \26936_27238 , RIfc52130_5956, \8917_9216 );
and \U$18119 ( \26937_27239 , RIe1ee430_4088, \8919_9218 );
and \U$18120 ( \26938_27240 , RIe1ebcd0_4060, \8921_9220 );
and \U$18121 ( \26939_27241 , RIe1e8fd0_4028, \8923_9222 );
and \U$18122 ( \26940_27242 , RIe1e62d0_3996, \8925_9224 );
and \U$18123 ( \26941_27243 , RIe1e35d0_3964, \8927_9226 );
and \U$18124 ( \26942_27244 , RIe1e08d0_3932, \8929_9228 );
and \U$18125 ( \26943_27245 , RIe1ddbd0_3900, \8931_9230 );
and \U$18126 ( \26944_27246 , RIe1daed0_3868, \8933_9232 );
and \U$18127 ( \26945_27247 , RIe1d81d0_3836, \8935_9234 );
and \U$18128 ( \26946_27248 , RIe1d27d0_3772, \8937_9236 );
and \U$18129 ( \26947_27249 , RIe1cfad0_3740, \8939_9238 );
and \U$18130 ( \26948_27250 , RIe1ccdd0_3708, \8941_9240 );
and \U$18131 ( \26949_27251 , RIe1ca0d0_3676, \8943_9242 );
and \U$18132 ( \26950_27252 , RIe1c73d0_3644, \8945_9244 );
and \U$18133 ( \26951_27253 , RIe1c46d0_3612, \8947_9246 );
and \U$18134 ( \26952_27254 , RIe1c19d0_3580, \8949_9248 );
and \U$18135 ( \26953_27255 , RIe1becd0_3548, \8951_9250 );
and \U$18136 ( \26954_27256 , RIfce0b88_7579, \8953_9252 );
and \U$18137 ( \26955_27257 , RIfc82808_6507, \8955_9254 );
and \U$18138 ( \26956_27258 , RIe1b9708_3487, \8957_9256 );
and \U$18139 ( \26957_27259 , RIe1b76b0_3464, \8959_9258 );
and \U$18140 ( \26958_27260 , RIfcd5bc0_7454, \8961_9260 );
and \U$18141 ( \26959_27261 , RIfcb69f0_7100, \8963_9262 );
and \U$18142 ( \26960_27262 , RIe1b54f0_3440, \8965_9264 );
and \U$18143 ( \26961_27263 , RIe1b4140_3426, \8967_9266 );
and \U$18144 ( \26962_27264 , RIfc89f90_6592, \8969_9268 );
and \U$18145 ( \26963_27265 , RIfce9af8_7681, \8971_9270 );
and \U$18146 ( \26964_27266 , RIe1b2958_3409, \8973_9272 );
and \U$18147 ( \26965_27267 , RIe1b0ea0_3390, \8975_9274 );
and \U$18148 ( \26966_27268 , RIfc4a138_5865, \8977_9276 );
and \U$18149 ( \26967_27269 , RIfc8a260_6594, \8979_9278 );
and \U$18150 ( \26968_27270 , RIe1ac850_3340, \8981_9280 );
and \U$18151 ( \26969_27271 , RIe1ab1d0_3324, \8983_9282 );
and \U$18152 ( \26970_27272 , RIe1a9010_3300, \8985_9284 );
and \U$18153 ( \26971_27273 , RIe1a6310_3268, \8987_9286 );
and \U$18154 ( \26972_27274 , RIe1a3610_3236, \8989_9288 );
and \U$18155 ( \26973_27275 , RIe1a0910_3204, \8991_9290 );
and \U$18156 ( \26974_27276 , RIe18ce10_2980, \8993_9292 );
and \U$18157 ( \26975_27277 , RIe179310_2756, \8995_9294 );
and \U$18158 ( \26976_27278 , RIe226c68_4731, \8997_9296 );
and \U$18159 ( \26977_27279 , RIe21b868_4603, \8999_9298 );
and \U$18160 ( \26978_27280 , RIe205068_4347, \9001_9300 );
and \U$18161 ( \26979_27281 , RIe1ff0c8_4279, \9003_9302 );
and \U$18162 ( \26980_27282 , RIe1f8480_4202, \9005_9304 );
and \U$18163 ( \26981_27283 , RIe1f0fc8_4119, \9007_9306 );
and \U$18164 ( \26982_27284 , RIe1d54d0_3804, \9009_9308 );
and \U$18165 ( \26983_27285 , RIe1bbfd0_3516, \9011_9310 );
and \U$18166 ( \26984_27286 , RIe1aee48_3367, \9013_9312 );
and \U$18167 ( \26985_27287 , RIe171480_2666, \9015_9314 );
or \U$18168 ( \26986_27288 , \26922_27224 , \26923_27225 , \26924_27226 , \26925_27227 , \26926_27228 , \26927_27229 , \26928_27230 , \26929_27231 , \26930_27232 , \26931_27233 , \26932_27234 , \26933_27235 , \26934_27236 , \26935_27237 , \26936_27238 , \26937_27239 , \26938_27240 , \26939_27241 , \26940_27242 , \26941_27243 , \26942_27244 , \26943_27245 , \26944_27246 , \26945_27247 , \26946_27248 , \26947_27249 , \26948_27250 , \26949_27251 , \26950_27252 , \26951_27253 , \26952_27254 , \26953_27255 , \26954_27256 , \26955_27257 , \26956_27258 , \26957_27259 , \26958_27260 , \26959_27261 , \26960_27262 , \26961_27263 , \26962_27264 , \26963_27265 , \26964_27266 , \26965_27267 , \26966_27268 , \26967_27269 , \26968_27270 , \26969_27271 , \26970_27272 , \26971_27273 , \26972_27274 , \26973_27275 , \26974_27276 , \26975_27277 , \26976_27278 , \26977_27279 , \26978_27280 , \26979_27281 , \26980_27282 , \26981_27283 , \26982_27284 , \26983_27285 , \26984_27286 , \26985_27287 );
or \U$18169 ( \26987_27289 , \26921_27223 , \26986_27288 );
_DC \g5f3f/U$1 ( \26988 , \26987_27289 , \9024_9323 );
xor g5f40_GF_PartitionCandidate( \26989_27291_nG5f40 , \26856 , \26988 );
buf \U$18170 ( \26990_27292 , \26989_27291_nG5f40 );
and \U$18171 ( \26991_27293 , \26504_26806 , \25471_25770 );
not \U$18172 ( \26992_27294 , \26991_27293 );
and \U$18173 ( \26993_27295 , \26990_27292 , \26992_27294 );
and \U$18174 ( \26994_27296 , \26724_27026 , \26993_27295 );
xor \U$18175 ( \26995_27297 , \26723_27025 , \26994_27296 );
and \U$18176 ( \26996_27298 , \26511_26813 , \26515_26817 );
and \U$18177 ( \26997_27299 , \26515_26817 , \26520_26822 );
and \U$18178 ( \26998_27300 , \26511_26813 , \26520_26822 );
or \U$18179 ( \26999_27301 , \26996_27298 , \26997_27299 , \26998_27300 );
xor \U$18180 ( \27000_27302 , \26995_27297 , \26999_27301 );
and \U$18181 ( \27001_27303 , \26530_26832 , \26534_26836 );
and \U$18182 ( \27002_27304 , \26534_26836 , \26539_26841 );
and \U$18183 ( \27003_27305 , \26530_26832 , \26539_26841 );
or \U$18184 ( \27004_27306 , \27001_27303 , \27002_27304 , \27003_27305 );
xor \U$18185 ( \27005_27307 , \27000_27302 , \27004_27306 );
xor \U$18186 ( \27006_27308 , \26719_27021 , \27005_27307 );
and \U$18187 ( \27007_27309 , \26527_26829 , \10681_10983 );
_DC \g65c2/U$1 ( \27008 , \26855_27157 , \9298_9597 );
_DC \g65c3/U$1 ( \27009 , \26987_27289 , \9024_9323 );
and g65c4_GF_PartitionCandidate( \27010_27312_nG65c4 , \27008 , \27009 );
buf \U$18188 ( \27011_27313 , \27010_27312_nG65c4 );
and \U$18189 ( \27012_27314 , \27011_27313 , \10389_10691 );
nor \U$18190 ( \27013_27315 , \27007_27309 , \27012_27314 );
xnor \U$18191 ( \27014_27316 , \27013_27315 , \10678_10980 );
and \U$18192 ( \27015_27317 , \18730_19032 , \16333_16635 );
and \U$18193 ( \27016_27318 , \19259_19558 , \15999_16301 );
nor \U$18194 ( \27017_27319 , \27015_27317 , \27016_27318 );
xnor \U$18195 ( \27018_27320 , \27017_27319 , \16323_16625 );
xor \U$18196 ( \27019_27321 , \27014_27316 , \27018_27320 );
and \U$18197 ( \27020_27322 , \10968_11270 , \25527_25826 );
and \U$18198 ( \27021_27323 , \11287_11586 , \24962_25264 );
nor \U$18199 ( \27022_27324 , \27020_27322 , \27021_27323 );
xnor \U$18200 ( \27023_27325 , \27022_27324 , \25474_25773 );
xor \U$18201 ( \27024_27326 , \27019_27321 , \27023_27325 );
and \U$18202 ( \27025_27327 , \20242_20544 , \15037_15336 );
and \U$18203 ( \27026_27328 , \20734_21033 , \14661_14963 );
nor \U$18204 ( \27027_27329 , \27025_27327 , \27026_27328 );
xnor \U$18205 ( \27028_27330 , \27027_27329 , \15043_15342 );
and \U$18206 ( \27029_27331 , \13377_13679 , \22243_22542 );
and \U$18207 ( \27030_27332 , \13725_14024 , \21801_22103 );
nor \U$18208 ( \27031_27333 , \27029_27331 , \27030_27332 );
xnor \U$18209 ( \27032_27334 , \27031_27333 , \22249_22548 );
xor \U$18210 ( \27033_27335 , \27028_27330 , \27032_27334 );
and \U$18211 ( \27034_27336 , \12146_12448 , \23839_24138 );
and \U$18212 ( \27035_27337 , \12470_12769 , \23328_23630 );
nor \U$18213 ( \27036_27338 , \27034_27336 , \27035_27337 );
xnor \U$18214 ( \27037_27339 , \27036_27338 , \23845_24144 );
xor \U$18215 ( \27038_27340 , \27033_27335 , \27037_27339 );
xor \U$18216 ( \27039_27341 , \27024_27326 , \27038_27340 );
and \U$18217 ( \27040_27342 , \21788_22090 , \13755_14054 );
and \U$18218 ( \27041_27343 , \22257_22556 , \13390_13692 );
nor \U$18219 ( \27042_27344 , \27040_27342 , \27041_27343 );
xnor \U$18220 ( \27043_27345 , \27042_27344 , \13736_14035 );
and \U$18221 ( \27044_27346 , \15965_16267 , \19235_19534 );
and \U$18222 ( \27045_27347 , \16353_16655 , \18743_19045 );
nor \U$18223 ( \27046_27348 , \27044_27346 , \27045_27347 );
xnor \U$18224 ( \27047_27349 , \27046_27348 , \19241_19540 );
xor \U$18225 ( \27048_27350 , \27043_27345 , \27047_27349 );
and \U$18226 ( \27049_27351 , \14648_14950 , \20706_21005 );
and \U$18227 ( \27050_27352 , \15022_15321 , \20255_20557 );
nor \U$18228 ( \27051_27353 , \27049_27351 , \27050_27352 );
xnor \U$18229 ( \27052_27354 , \27051_27353 , \20712_21011 );
xor \U$18230 ( \27053_27355 , \27048_27350 , \27052_27354 );
xor \U$18231 ( \27054_27356 , \27039_27341 , \27053_27355 );
xor \U$18232 ( \27055_27357 , \27006_27308 , \27054_27356 );
xor \U$18233 ( \27056_27358 , \26715_27017 , \27055_27357 );
and \U$18234 ( \27057_27359 , \26556_26858 , \26560_26862 );
and \U$18235 ( \27058_27360 , \26560_26862 , \26572_26874 );
and \U$18236 ( \27059_27361 , \26556_26858 , \26572_26874 );
or \U$18237 ( \27060_27362 , \27057_27359 , \27058_27360 , \27059_27361 );
and \U$18238 ( \27061_27363 , \26204_26506 , \26228_26530 );
and \U$18239 ( \27062_27364 , \26228_26530 , \26541_26843 );
and \U$18240 ( \27063_27365 , \26204_26506 , \26541_26843 );
or \U$18241 ( \27064_27366 , \27061_27363 , \27062_27364 , \27063_27365 );
xor \U$18242 ( \27065_27367 , \27060_27362 , \27064_27366 );
and \U$18243 ( \27066_27368 , \26565_26867 , \26566_26868 );
and \U$18244 ( \27067_27369 , \26566_26868 , \26571_26873 );
and \U$18245 ( \27068_27370 , \26565_26867 , \26571_26873 );
or \U$18246 ( \27069_27371 , \27066_27368 , \27067_27369 , \27068_27370 );
and \U$18247 ( \27070_27372 , \26507_26809 , \26521_26823 );
and \U$18248 ( \27071_27373 , \26521_26823 , \26540_26842 );
and \U$18249 ( \27072_27374 , \26507_26809 , \26540_26842 );
or \U$18250 ( \27073_27375 , \27070_27372 , \27071_27373 , \27072_27374 );
xor \U$18251 ( \27074_27376 , \27069_27371 , \27073_27375 );
and \U$18252 ( \27075_27377 , \26233_26535 , \26237_26539 );
and \U$18253 ( \27076_27378 , \26237_26539 , \26506_26808 );
and \U$18254 ( \27077_27379 , \26233_26535 , \26506_26808 );
or \U$18255 ( \27078_27380 , \27075_27377 , \27076_27378 , \27077_27379 );
and \U$18256 ( \27079_27381 , \26217_26519 , \26221_26523 );
and \U$18257 ( \27080_27382 , \26221_26523 , \26226_26528 );
and \U$18258 ( \27081_27383 , \26217_26519 , \26226_26528 );
or \U$18259 ( \27082_27384 , \27079_27381 , \27080_27382 , \27081_27383 );
xor \U$18260 ( \27083_27385 , \27078_27380 , \27082_27384 );
and \U$18261 ( \27084_27386 , \23315_23617 , \12491_12790 );
and \U$18262 ( \27085_27387 , \23900_24199 , \12159_12461 );
nor \U$18263 ( \27086_27388 , \27084_27386 , \27085_27387 );
xnor \U$18264 ( \27087_27389 , \27086_27388 , \12481_12780 );
and \U$18265 ( \27088_27390 , \17325_17627 , \17791_18090 );
and \U$18266 ( \27089_27391 , \17736_18035 , \17353_17655 );
nor \U$18267 ( \27090_27392 , \27088_27390 , \27089_27391 );
xnor \U$18268 ( \27091_27393 , \27090_27392 , \17747_18046 );
xor \U$18269 ( \27092_27394 , \27087_27389 , \27091_27393 );
xor \U$18270 ( \27093_27395 , \26990_27292 , \26504_26806 );
not \U$18271 ( \27094_27396 , \26505_26807 );
and \U$18272 ( \27095_27397 , \27093_27395 , \27094_27396 );
and \U$18273 ( \27096_27398 , \10385_10687 , \27095_27397 );
and \U$18274 ( \27097_27399 , \10686_10988 , \26505_26807 );
nor \U$18275 ( \27098_27400 , \27096_27398 , \27097_27399 );
xnor \U$18276 ( \27099_27401 , \27098_27400 , \26993_27295 );
xor \U$18277 ( \27100_27402 , \27092_27394 , \27099_27401 );
xor \U$18278 ( \27101_27403 , \27083_27385 , \27100_27402 );
xor \U$18279 ( \27102_27404 , \27074_27376 , \27101_27403 );
xor \U$18280 ( \27103_27405 , \27065_27367 , \27102_27404 );
xor \U$18281 ( \27104_27406 , \27056_27358 , \27103_27405 );
and \U$18282 ( \27105_27407 , \26200_26502 , \26542_26844 );
and \U$18283 ( \27106_27408 , \26542_26844 , \26574_26876 );
and \U$18284 ( \27107_27409 , \26200_26502 , \26574_26876 );
or \U$18285 ( \27108_27410 , \27105_27407 , \27106_27408 , \27107_27409 );
xor \U$18286 ( \27109_27411 , \27104_27406 , \27108_27410 );
and \U$18287 ( \27110_27412 , \26575_26877 , \26579_26881 );
and \U$18288 ( \27111_27413 , \26580_26882 , \26583_26885 );
or \U$18289 ( \27112_27414 , \27110_27412 , \27111_27413 );
xor \U$18290 ( \27113_27415 , \27109_27411 , \27112_27414 );
buf g9bc3_GF_PartitionCandidate( \27114_27416_nG9bc3 , \27113_27415 );
and \U$18291 ( \27115_27417 , \10402_10704 , \27114_27416_nG9bc3 );
or \U$18292 ( \27116_27418 , \26711_27013 , \27115_27417 );
xor \U$18293 ( \27117_27419 , \10399_10703 , \27116_27418 );
buf \U$18294 ( \27118_27420 , \27117_27419 );
buf \U$18296 ( \27119_27421 , \27118_27420 );
xor \U$18297 ( \27120_27422 , \26710_27012 , \27119_27421 );
buf \U$18298 ( \27121_27423 , \27120_27422 );
xor \U$18299 ( \27122_27424 , \26698_27000 , \27121_27423 );
and \U$18300 ( \27123_27425 , \26633_26935 , \26639_26941 );
and \U$18301 ( \27124_27426 , \26633_26935 , \26646_26948 );
and \U$18302 ( \27125_27427 , \26639_26941 , \26646_26948 );
or \U$18303 ( \27126_27428 , \27123_27425 , \27124_27426 , \27125_27427 );
buf \U$18304 ( \27127_27429 , \27126_27428 );
and \U$18305 ( \27128_27430 , \26128_26427 , \26132_26434 );
buf \U$18306 ( \27129_27431 , \27128_27430 );
buf \U$18308 ( \27130_27432 , \27129_27431 );
and \U$18309 ( \27131_27433 , \25044_24792 , \10981_11283_nG9c08 );
and \U$18310 ( \27132_27434 , \24490_24789 , \11299_11598_nG9c05 );
or \U$18311 ( \27133_27435 , \27131_27433 , \27132_27434 );
xor \U$18312 ( \27134_27436 , \24489_24788 , \27133_27435 );
buf \U$18313 ( \27135_27437 , \27134_27436 );
buf \U$18315 ( \27136_27438 , \27135_27437 );
xor \U$18316 ( \27137_27439 , \27130_27432 , \27136_27438 );
buf \U$18317 ( \27138_27440 , \27137_27439 );
not \U$17303 ( \27139_26429 , \26129_26428 );
xor \U$17304 ( \27140_26430 , \26123_26422_nG440c , \26126_26425_nG440f );
and \U$17305 ( \27141_26431 , \27139_26429 , \27140_26430 );
and \U$18318 ( \27142_27441 , \27141_26431 , \10392_10694_nG9c0e );
and \U$18319 ( \27143_27442 , \26129_26428 , \10693_10995_nG9c0b );
or \U$18320 ( \27144_27443 , \27142_27441 , \27143_27442 );
xor \U$18321 ( \27145_27444 , \26128_26427 , \27144_27443 );
buf \U$18322 ( \27146_27445 , \27145_27444 );
buf \U$18324 ( \27147_27446 , \27146_27445 );
xor \U$18325 ( \27148_27447 , \27138_27440 , \27147_27446 );
and \U$18326 ( \27149_27448 , \23495_23201 , \12168_12470_nG9c02 );
and \U$18327 ( \27150_27449 , \22899_23198 , \12502_12801_nG9bff );
or \U$18328 ( \27151_27450 , \27149_27448 , \27150_27449 );
xor \U$18329 ( \27152_27451 , \22898_23197 , \27151_27450 );
buf \U$18330 ( \27153_27452 , \27152_27451 );
buf \U$18332 ( \27154_27453 , \27153_27452 );
xor \U$18333 ( \27155_27454 , \27148_27447 , \27154_27453 );
buf \U$18334 ( \27156_27455 , \27155_27454 );
xor \U$18335 ( \27157_27456 , \27127_27429 , \27156_27455 );
and \U$18336 ( \27158_27457 , \18908_18702 , \16013_16315_nG9bf0 );
and \U$18337 ( \27159_27458 , \18400_18699 , \16378_16680_nG9bed );
or \U$18338 ( \27160_27459 , \27158_27457 , \27159_27458 );
xor \U$18339 ( \27161_27460 , \18399_18698 , \27160_27459 );
buf \U$18340 ( \27162_27461 , \27161_27460 );
buf \U$18342 ( \27163_27462 , \27162_27461 );
xor \U$18343 ( \27164_27463 , \27157_27456 , \27163_27462 );
buf \U$18344 ( \27165_27464 , \27164_27463 );
and \U$18345 ( \27166_27465 , \16405_15940 , \18789_19091_nG9be4 );
and \U$18346 ( \27167_27466 , \15638_15937 , \19287_19586_nG9be1 );
or \U$18347 ( \27168_27467 , \27166_27465 , \27167_27466 );
xor \U$18348 ( \27169_27468 , \15637_15936 , \27168_27467 );
buf \U$18349 ( \27170_27469 , \27169_27468 );
buf \U$18351 ( \27171_27470 , \27170_27469 );
xor \U$18352 ( \27172_27471 , \27165_27464 , \27171_27470 );
and \U$18353 ( \27173_27472 , \14710_14631 , \20306_20608_nG9bde );
and \U$18354 ( \27174_27473 , \14329_14628 , \20787_21086_nG9bdb );
or \U$18355 ( \27175_27474 , \27173_27472 , \27174_27473 );
xor \U$18356 ( \27176_27475 , \14328_14627 , \27175_27474 );
buf \U$18357 ( \27177_27476 , \27176_27475 );
buf \U$18359 ( \27178_27477 , \27177_27476 );
xor \U$18360 ( \27179_27478 , \27172_27471 , \27178_27477 );
buf \U$18361 ( \27180_27479 , \27179_27478 );
and \U$18362 ( \27181_27480 , \26157_26459 , \26163_26465 );
buf \U$18363 ( \27182_27481 , \27181_27480 );
and \U$18364 ( \27183_27482 , \21908_21658 , \13403_13705_nG9bfc );
and \U$18365 ( \27184_27483 , \21356_21655 , \13771_14070_nG9bf9 );
or \U$18366 ( \27185_27484 , \27183_27482 , \27184_27483 );
xor \U$18367 ( \27186_27485 , \21355_21654 , \27185_27484 );
buf \U$18368 ( \27187_27486 , \27186_27485 );
buf \U$18370 ( \27188_27487 , \27187_27486 );
xor \U$18371 ( \27189_27488 , \27182_27481 , \27188_27487 );
and \U$18372 ( \27190_27489 , \20353_20155 , \14682_14984_nG9bf6 );
and \U$18373 ( \27191_27490 , \19853_20152 , \15074_15373_nG9bf3 );
or \U$18374 ( \27192_27491 , \27190_27489 , \27191_27490 );
xor \U$18375 ( \27193_27492 , \19852_20151 , \27192_27491 );
buf \U$18376 ( \27194_27493 , \27193_27492 );
buf \U$18378 ( \27195_27494 , \27194_27493 );
xor \U$18379 ( \27196_27495 , \27189_27488 , \27195_27494 );
buf \U$18380 ( \27197_27496 , \27196_27495 );
and \U$18381 ( \27198_27497 , \26151_26453 , \26165_26467 );
and \U$18382 ( \27199_27498 , \26151_26453 , \26172_26474 );
and \U$18383 ( \27200_27499 , \26165_26467 , \26172_26474 );
or \U$18384 ( \27201_27500 , \27198_27497 , \27199_27498 , \27200_27499 );
buf \U$18385 ( \27202_27501 , \27201_27500 );
xor \U$18386 ( \27203_27502 , \27197_27496 , \27202_27501 );
and \U$18387 ( \27204_27503 , \17437_17297 , \17363_17665_nG9bea );
and \U$18388 ( \27205_27504 , \16995_17294 , \17808_18107_nG9be7 );
or \U$18389 ( \27206_27505 , \27204_27503 , \27205_27504 );
xor \U$18390 ( \27207_27506 , \16994_17293 , \27206_27505 );
buf \U$18391 ( \27208_27507 , \27207_27506 );
buf \U$18393 ( \27209_27508 , \27208_27507 );
xor \U$18394 ( \27210_27509 , \27203_27502 , \27209_27508 );
buf \U$18395 ( \27211_27510 , \27210_27509 );
xor \U$18396 ( \27212_27511 , \27180_27479 , \27211_27510 );
and \U$18397 ( \27213_27512 , \12183_12157 , \23394_23696_nG9bd2 );
and \U$18398 ( \27214_27513 , \11855_12154 , \23927_24226_nG9bcf );
or \U$18399 ( \27215_27514 , \27213_27512 , \27214_27513 );
xor \U$18400 ( \27216_27515 , \11854_12153 , \27215_27514 );
buf \U$18401 ( \27217_27516 , \27216_27515 );
buf \U$18403 ( \27218_27517 , \27217_27516 );
xor \U$18404 ( \27219_27518 , \27212_27511 , \27218_27517 );
buf \U$18405 ( \27220_27519 , \27219_27518 );
xor \U$18406 ( \27221_27520 , \27122_27424 , \27220_27519 );
buf \U$18407 ( \27222_27521 , \27221_27520 );
and \U$18408 ( \27223_27522 , \26146_26448 , \26592_26894 );
and \U$18409 ( \27224_27523 , \26146_26448 , \26598_26900 );
and \U$18410 ( \27225_27524 , \26592_26894 , \26598_26900 );
or \U$18411 ( \27226_27525 , \27223_27522 , \27224_27523 , \27225_27524 );
buf \U$18412 ( \27227_27526 , \27226_27525 );
xor \U$18413 ( \27228_27527 , \27222_27521 , \27227_27526 );
and \U$18414 ( \27229_27528 , \26610_26912 , \26616_26918 );
and \U$18415 ( \27230_27529 , \26610_26912 , \26623_26925 );
and \U$18416 ( \27231_27530 , \26616_26918 , \26623_26925 );
or \U$18417 ( \27232_27531 , \27229_27528 , \27230_27529 , \27231_27530 );
buf \U$18418 ( \27233_27532 , \27232_27531 );
and \U$18419 ( \27234_27533 , \26174_26476 , \26180_26482 );
and \U$18420 ( \27235_27534 , \26174_26476 , \26187_26489 );
and \U$18421 ( \27236_27535 , \26180_26482 , \26187_26489 );
or \U$18422 ( \27237_27536 , \27234_27533 , \27235_27534 , \27236_27535 );
buf \U$18423 ( \27238_27537 , \27237_27536 );
and \U$18424 ( \27239_27538 , \26631_26933 , \26648_26950 );
and \U$18425 ( \27240_27539 , \26631_26933 , \26655_26957 );
and \U$18426 ( \27241_27540 , \26648_26950 , \26655_26957 );
or \U$18427 ( \27242_27541 , \27239_27538 , \27240_27539 , \27241_27540 );
buf \U$18428 ( \27243_27542 , \27242_27541 );
xor \U$18429 ( \27244_27543 , \27238_27537 , \27243_27542 );
and \U$18430 ( \27245_27544 , \13431_13370 , \21827_22129_nG9bd8 );
and \U$18431 ( \27246_27545 , \13068_13367 , \22330_22629_nG9bd5 );
or \U$18432 ( \27247_27546 , \27245_27544 , \27246_27545 );
xor \U$18433 ( \27248_27547 , \13067_13366 , \27247_27546 );
buf \U$18434 ( \27249_27548 , \27248_27547 );
buf \U$18436 ( \27250_27549 , \27249_27548 );
xor \U$18437 ( \27251_27550 , \27244_27543 , \27250_27549 );
buf \U$18438 ( \27252_27551 , \27251_27550 );
xor \U$18439 ( \27253_27552 , \27233_27532 , \27252_27551 );
and \U$18440 ( \27254_27553 , \26189_26491 , \26194_26496 );
and \U$18441 ( \27255_27554 , \26189_26491 , \26590_26892 );
and \U$18442 ( \27256_27555 , \26194_26496 , \26590_26892 );
or \U$18443 ( \27257_27556 , \27254_27553 , \27255_27554 , \27256_27555 );
buf \U$18444 ( \27258_27557 , \27257_27556 );
xor \U$18445 ( \27259_27558 , \27253_27552 , \27258_27557 );
buf \U$18446 ( \27260_27559 , \27259_27558 );
xor \U$18447 ( \27261_27560 , \27228_27527 , \27260_27559 );
and \U$18448 ( \27262_27561 , \26693_26995 , \27261_27560 );
and \U$18449 ( \27263_27562 , \26683_26985 , \26687_26989 );
and \U$18450 ( \27264_27563 , \26683_26985 , \26692_26994 );
and \U$18451 ( \27265_27564 , \26687_26989 , \26692_26994 );
or \U$18452 ( \27266_27565 , \27263_27562 , \27264_27563 , \27265_27564 );
xor \U$18453 ( \27267_27566 , \27262_27561 , \27266_27565 );
and \U$18454 ( \27268_27567 , RIdec5c48_714, \8760_9059 );
and \U$18455 ( \27269_27568 , RIdec2f48_682, \8762_9061 );
and \U$18456 ( \27270_27569 , RIfc7c160_6434, \8764_9063 );
and \U$18457 ( \27271_27570 , RIdec0248_650, \8766_9065 );
and \U$18458 ( \27272_27571 , RIfcb38b8_7065, \8768_9067 );
and \U$18459 ( \27273_27572 , RIdebd548_618, \8770_9069 );
and \U$18460 ( \27274_27573 , RIdeba848_586, \8772_9071 );
and \U$18461 ( \27275_27574 , RIdeb7b48_554, \8774_9073 );
and \U$18462 ( \27276_27575 , RIfce7c08_7659, \8776_9075 );
and \U$18463 ( \27277_27576 , RIdeb2148_490, \8778_9077 );
and \U$18464 ( \27278_27577 , RIfce7aa0_7658, \8780_9079 );
and \U$18465 ( \27279_27578 , RIdeaf448_458, \8782_9081 );
and \U$18466 ( \27280_27579 , RIfca38c8_6883, \8784_9083 );
and \U$18467 ( \27281_27580 , RIdeab7d0_426, \8786_9085 );
and \U$18468 ( \27282_27581 , RIdea4ed0_394, \8788_9087 );
and \U$18469 ( \27283_27582 , RIde9e5d0_362, \8790_9089 );
and \U$18470 ( \27284_27583 , RIfc41e70_5772, \8792_9091 );
and \U$18471 ( \27285_27584 , RIfc5b0a0_6058, \8794_9093 );
and \U$18472 ( \27286_27585 , RIfcdbb60_7522, \8796_9095 );
and \U$18473 ( \27287_27586 , RIfc78650_6392, \8798_9097 );
and \U$18474 ( \27288_27587 , RIfea92d8_8241, \8800_9099 );
and \U$18475 ( \27289_27588 , RIde8e5e0_284, \8802_9101 );
and \U$18476 ( \27290_27589 , RIfea0d40_8174, \8804_9103 );
and \U$18477 ( \27291_27590 , RIfea0bd8_8173, \8806_9105 );
and \U$18478 ( \27292_27591 , RIfcdf508_7563, \8808_9107 );
and \U$18479 ( \27293_27592 , RIfcb1b30_7044, \8810_9109 );
and \U$18480 ( \27294_27593 , RIfc5ccc0_6078, \8812_9111 );
and \U$18481 ( \27295_27594 , RIfcb16f8_7041, \8814_9113 );
and \U$18482 ( \27296_27595 , RIfc77b10_6384, \8816_9115 );
and \U$18483 ( \27297_27596 , RIe16beb8_2605, \8818_9117 );
and \U$18484 ( \27298_27597 , RIe169e60_2582, \8820_9119 );
and \U$18485 ( \27299_27598 , RIe168510_2564, \8822_9121 );
and \U$18486 ( \27300_27599 , RIe165c48_2535, \8824_9123 );
and \U$18487 ( \27301_27600 , RIe162f48_2503, \8826_9125 );
and \U$18488 ( \27302_27601 , RIfc4f9d0_5928, \8828_9127 );
and \U$18489 ( \27303_27602 , RIe160248_2471, \8830_9129 );
and \U$18490 ( \27304_27603 , RIfc4e8f0_5916, \8832_9131 );
and \U$18491 ( \27305_27604 , RIe15d548_2439, \8834_9133 );
and \U$18492 ( \27306_27605 , RIe157b48_2375, \8836_9135 );
and \U$18493 ( \27307_27606 , RIe154e48_2343, \8838_9137 );
and \U$18494 ( \27308_27607 , RIfc4e1e8_5911, \8840_9139 );
and \U$18495 ( \27309_27608 , RIe152148_2311, \8842_9141 );
and \U$18496 ( \27310_27609 , RIfc868b8_6553, \8844_9143 );
and \U$18497 ( \27311_27610 , RIe14f448_2279, \8846_9145 );
and \U$18498 ( \27312_27611 , RIfc865e8_6551, \8848_9147 );
and \U$18499 ( \27313_27612 , RIe14c748_2247, \8850_9149 );
and \U$18500 ( \27314_27613 , RIe149a48_2215, \8852_9151 );
and \U$18501 ( \27315_27614 , RIe146d48_2183, \8854_9153 );
and \U$18502 ( \27316_27615 , RIfc9eb70_6828, \8856_9155 );
and \U$18503 ( \27317_27616 , RIfc9ecd8_6829, \8858_9157 );
and \U$18504 ( \27318_27617 , RIfcc5630_7268, \8860_9159 );
and \U$18505 ( \27319_27618 , RIfc83bb8_6521, \8862_9161 );
and \U$18506 ( \27320_27619 , RIe141618_2121, \8864_9163 );
and \U$18507 ( \27321_27620 , RIfea0ea8_8175, \8866_9165 );
and \U$18508 ( \27322_27621 , RIdf3d1f8_2072, \8868_9167 );
and \U$18509 ( \27323_27622 , RIdf3ac00_2045, \8870_9169 );
and \U$18510 ( \27324_27623 , RIee308e0_5011, \8872_9171 );
and \U$18511 ( \27325_27624 , RIfcd3cd0_7432, \8874_9173 );
and \U$18512 ( \27326_27625 , RIfc84e00_6534, \8876_9175 );
and \U$18513 ( \27327_27626 , RIfc834b0_6516, \8878_9177 );
and \U$18514 ( \27328_27627 , RIdf36010_1991, \8880_9179 );
and \U$18515 ( \27329_27628 , RIdf33a18_1964, \8882_9181 );
and \U$18516 ( \27330_27629 , RIdf31858_1940, \8884_9183 );
and \U$18517 ( \27331_27630 , RIdf2f968_1918, \8886_9185 );
or \U$18518 ( \27332_27631 , \27268_27567 , \27269_27568 , \27270_27569 , \27271_27570 , \27272_27571 , \27273_27572 , \27274_27573 , \27275_27574 , \27276_27575 , \27277_27576 , \27278_27577 , \27279_27578 , \27280_27579 , \27281_27580 , \27282_27581 , \27283_27582 , \27284_27583 , \27285_27584 , \27286_27585 , \27287_27586 , \27288_27587 , \27289_27588 , \27290_27589 , \27291_27590 , \27292_27591 , \27293_27592 , \27294_27593 , \27295_27594 , \27296_27595 , \27297_27596 , \27298_27597 , \27299_27598 , \27300_27599 , \27301_27600 , \27302_27601 , \27303_27602 , \27304_27603 , \27305_27604 , \27306_27605 , \27307_27606 , \27308_27607 , \27309_27608 , \27310_27609 , \27311_27610 , \27312_27611 , \27313_27612 , \27314_27613 , \27315_27614 , \27316_27615 , \27317_27616 , \27318_27617 , \27319_27618 , \27320_27619 , \27321_27620 , \27322_27621 , \27323_27622 , \27324_27623 , \27325_27624 , \27326_27625 , \27327_27626 , \27328_27627 , \27329_27628 , \27330_27629 , \27331_27630 );
and \U$18519 ( \27333_27632 , RIee2c128_4960, \8889_9188 );
and \U$18520 ( \27334_27633 , RIee2a7d8_4942, \8891_9190 );
and \U$18521 ( \27335_27634 , RIee292c0_4927, \8893_9192 );
and \U$18522 ( \27336_27635 , RIee28078_4914, \8895_9194 );
and \U$18523 ( \27337_27636 , RIdf2a940_1861, \8897_9196 );
and \U$18524 ( \27338_27637 , RIdf28780_1837, \8899_9198 );
and \U$18525 ( \27339_27638 , RIfea0a70_8172, \8901_9200 );
and \U$18526 ( \27340_27639 , RIfea0908_8171, \8903_9202 );
and \U$18527 ( \27341_27640 , RIfcd4f18_7445, \8905_9204 );
and \U$18528 ( \27342_27641 , RIfca0628_6847, \8907_9206 );
and \U$18529 ( \27343_27642 , RIdf23050_1775, \8909_9208 );
and \U$18530 ( \27344_27643 , RIfcd3190_7424, \8911_9210 );
and \U$18531 ( \27345_27644 , RIdf21b38_1760, \8913_9212 );
and \U$18532 ( \27346_27645 , RIdf20080_1741, \8915_9214 );
and \U$18533 ( \27347_27646 , RIdf1b328_1686, \8917_9216 );
and \U$18534 ( \27348_27647 , RIdf199d8_1668, \8919_9218 );
and \U$18535 ( \27349_27648 , RIdf17818_1644, \8921_9220 );
and \U$18536 ( \27350_27649 , RIdf14b18_1612, \8923_9222 );
and \U$18537 ( \27351_27650 , RIdf11e18_1580, \8925_9224 );
and \U$18538 ( \27352_27651 , RIdf0f118_1548, \8927_9226 );
and \U$18539 ( \27353_27652 , RIdf0c418_1516, \8929_9228 );
and \U$18540 ( \27354_27653 , RIdf09718_1484, \8931_9230 );
and \U$18541 ( \27355_27654 , RIdf06a18_1452, \8933_9232 );
and \U$18542 ( \27356_27655 , RIdf03d18_1420, \8935_9234 );
and \U$18543 ( \27357_27656 , RIdefe318_1356, \8937_9236 );
and \U$18544 ( \27358_27657 , RIdefb618_1324, \8939_9238 );
and \U$18545 ( \27359_27658 , RIdef8918_1292, \8941_9240 );
and \U$18546 ( \27360_27659 , RIdef5c18_1260, \8943_9242 );
and \U$18547 ( \27361_27660 , RIdef2f18_1228, \8945_9244 );
and \U$18548 ( \27362_27661 , RIdef0218_1196, \8947_9246 );
and \U$18549 ( \27363_27662 , RIdeed518_1164, \8949_9248 );
and \U$18550 ( \27364_27663 , RIdeea818_1132, \8951_9250 );
and \U$18551 ( \27365_27664 , RIfcdf3a0_7562, \8953_9252 );
and \U$18552 ( \27366_27665 , RIfca5218_6901, \8955_9254 );
and \U$18553 ( \27367_27666 , RIfcdc538_7529, \8957_9256 );
and \U$18554 ( \27368_27667 , RIfcdc6a0_7530, \8959_9258 );
and \U$18555 ( \27369_27668 , RIdee50e8_1070, \8961_9260 );
and \U$18556 ( \27370_27669 , RIdee3360_1049, \8963_9262 );
and \U$18557 ( \27371_27670 , RIfea07a0_8170, \8965_9264 );
and \U$18558 ( \27372_27671 , RIdedefe0_1001, \8967_9266 );
and \U$18559 ( \27373_27672 , RIfcb0d20_7034, \8969_9268 );
and \U$18560 ( \27374_27673 , RIfcd4978_7441, \8971_9270 );
and \U$18561 ( \27375_27674 , RIfca49a8_6895, \8973_9272 );
and \U$18562 ( \27376_27675 , RIfca1708_6859, \8975_9274 );
and \U$18563 ( \27377_27676 , RIded9fb8_944, \8977_9276 );
and \U$18564 ( \27378_27677 , RIded79c0_917, \8979_9278 );
and \U$18565 ( \27379_27678 , RIded5ad0_895, \8981_9280 );
and \U$18566 ( \27380_27679 , RIfeab498_8265, \8983_9282 );
and \U$18567 ( \27381_27680 , RIded1048_842, \8985_9284 );
and \U$18568 ( \27382_27681 , RIdece348_810, \8987_9286 );
and \U$18569 ( \27383_27682 , RIdecb648_778, \8989_9288 );
and \U$18570 ( \27384_27683 , RIdec8948_746, \8991_9290 );
and \U$18571 ( \27385_27684 , RIdeb4e48_522, \8993_9292 );
and \U$18572 ( \27386_27685 , RIde97cd0_330, \8995_9294 );
and \U$18573 ( \27387_27686 , RIe16ea50_2636, \8997_9296 );
and \U$18574 ( \27388_27687 , RIe15a848_2407, \8999_9298 );
and \U$18575 ( \27389_27688 , RIe144048_2151, \9001_9300 );
and \U$18576 ( \27390_27689 , RIdf38a40_2021, \9003_9302 );
and \U$18577 ( \27391_27690 , RIdf2d0a0_1889, \9005_9304 );
and \U$18578 ( \27392_27691 , RIdf1d920_1713, \9007_9306 );
and \U$18579 ( \27393_27692 , RIdf01018_1388, \9009_9308 );
and \U$18580 ( \27394_27693 , RIdee7b18_1100, \9011_9310 );
and \U$18581 ( \27395_27694 , RIdedc880_973, \9013_9312 );
and \U$18582 ( \27396_27695 , RIde7dc18_203, \9015_9314 );
or \U$18583 ( \27397_27696 , \27333_27632 , \27334_27633 , \27335_27634 , \27336_27635 , \27337_27636 , \27338_27637 , \27339_27638 , \27340_27639 , \27341_27640 , \27342_27641 , \27343_27642 , \27344_27643 , \27345_27644 , \27346_27645 , \27347_27646 , \27348_27647 , \27349_27648 , \27350_27649 , \27351_27650 , \27352_27651 , \27353_27652 , \27354_27653 , \27355_27654 , \27356_27655 , \27357_27656 , \27358_27657 , \27359_27658 , \27360_27659 , \27361_27660 , \27362_27661 , \27363_27662 , \27364_27663 , \27365_27664 , \27366_27665 , \27367_27666 , \27368_27667 , \27369_27668 , \27370_27669 , \27371_27670 , \27372_27671 , \27373_27672 , \27374_27673 , \27375_27674 , \27376_27675 , \27377_27676 , \27378_27677 , \27379_27678 , \27380_27679 , \27381_27680 , \27382_27681 , \27383_27682 , \27384_27683 , \27385_27684 , \27386_27685 , \27387_27686 , \27388_27687 , \27389_27688 , \27390_27689 , \27391_27690 , \27392_27691 , \27393_27692 , \27394_27693 , \27395_27694 , \27396_27695 );
or \U$18584 ( \27398_27697 , \27332_27631 , \27397_27696 );
_DC \g2449/U$1 ( \27399 , \27398_27697 , \9024_9323 );
buf \U$18585 ( \27400_27699 , \27399 );
and \U$18586 ( \27401_27700 , RIe19dee0_3174, \9034_9333 );
and \U$18587 ( \27402_27701 , RIe19b1e0_3142, \9036_9335 );
and \U$18588 ( \27403_27702 , RIfc67580_6198, \9038_9337 );
and \U$18589 ( \27404_27703 , RIe1984e0_3110, \9040_9339 );
and \U$18590 ( \27405_27704 , RIfccb030_7332, \9042_9341 );
and \U$18591 ( \27406_27705 , RIe1957e0_3078, \9044_9343 );
and \U$18592 ( \27407_27706 , RIe192ae0_3046, \9046_9345 );
and \U$18593 ( \27408_27707 , RIe18fde0_3014, \9048_9347 );
and \U$18594 ( \27409_27708 , RIe18a3e0_2950, \9050_9349 );
and \U$18595 ( \27410_27709 , RIe1876e0_2918, \9052_9351 );
and \U$18596 ( \27411_27710 , RIfc6a550_6232, \9054_9353 );
and \U$18597 ( \27412_27711 , RIe1849e0_2886, \9056_9355 );
and \U$18598 ( \27413_27712 , RIfcaa7e0_6962, \9058_9357 );
and \U$18599 ( \27414_27713 , RIe181ce0_2854, \9060_9359 );
and \U$18600 ( \27415_27714 , RIe17efe0_2822, \9062_9361 );
and \U$18601 ( \27416_27715 , RIe17c2e0_2790, \9064_9363 );
and \U$18602 ( \27417_27716 , RIfc65d98_6181, \9066_9365 );
and \U$18603 ( \27418_27717 , RIfc65690_6176, \9068_9367 );
and \U$18604 ( \27419_27718 , RIe1772b8_2733, \9070_9369 );
and \U$18605 ( \27420_27719 , RIfea0638_8169, \9072_9371 );
and \U$18606 ( \27421_27720 , RIfcca928_7327, \9074_9373 );
and \U$18607 ( \27422_27721 , RIfc607d0_6120, \9076_9375 );
and \U$18608 ( \27423_27722 , RIfc65258_6173, \9078_9377 );
and \U$18609 ( \27424_27723 , RIee3d798_5158, \9080_9379 );
and \U$18610 ( \27425_27724 , RIee3c3e8_5144, \9082_9381 );
and \U$18611 ( \27426_27725 , RIfca9430_6948, \9084_9383 );
and \U$18612 ( \27427_27726 , RIee39f58_5118, \9086_9385 );
and \U$18613 ( \27428_27727 , RIe174018_2697, \9088_9387 );
and \U$18614 ( \27429_27728 , RIfcecf00_7718, \9090_9389 );
and \U$18615 ( \27430_27729 , RIfc650f0_6172, \9092_9391 );
and \U$18616 ( \27431_27730 , RIf16e5a8_5715, \9094_9393 );
and \U$18617 ( \27432_27731 , RIfc43a90_5792, \9096_9395 );
and \U$18618 ( \27433_27732 , RIfc65528_6175, \9098_9397 );
and \U$18619 ( \27434_27733 , RIe224238_4701, \9100_9399 );
and \U$18620 ( \27435_27734 , RIfca9f70_6956, \9102_9401 );
and \U$18621 ( \27436_27735 , RIe221538_4669, \9104_9403 );
and \U$18622 ( \27437_27736 , RIfc6b4c8_6243, \9106_9405 );
and \U$18623 ( \27438_27737 , RIe21e838_4637, \9108_9407 );
and \U$18624 ( \27439_27738 , RIe218e38_4573, \9110_9409 );
and \U$18625 ( \27440_27739 , RIe216138_4541, \9112_9411 );
and \U$18626 ( \27441_27740 , RIfc3fda0_5752, \9114_9413 );
and \U$18627 ( \27442_27741 , RIe213438_4509, \9116_9415 );
and \U$18628 ( \27443_27742 , RIfc61310_6128, \9118_9417 );
and \U$18629 ( \27444_27743 , RIe210738_4477, \9120_9419 );
and \U$18630 ( \27445_27744 , RIfc60c08_6123, \9122_9421 );
and \U$18631 ( \27446_27745 , RIe20da38_4445, \9124_9423 );
and \U$18632 ( \27447_27746 , RIe20ad38_4413, \9126_9425 );
and \U$18633 ( \27448_27747 , RIe208038_4381, \9128_9427 );
and \U$18634 ( \27449_27748 , RIfc66ba8_6191, \9130_9429 );
and \U$18635 ( \27450_27749 , RIfccbcd8_7341, \9132_9431 );
and \U$18636 ( \27451_27750 , RIe202bd8_4321, \9134_9433 );
and \U$18637 ( \27452_27751 , RIe200fb8_4301, \9136_9435 );
and \U$18638 ( \27453_27752 , RIfcadbe8_6999, \9138_9437 );
and \U$18639 ( \27454_27753 , RIfccbe40_7342, \9140_9439 );
and \U$18640 ( \27455_27754 , RIfca7540_6926, \9142_9441 );
and \U$18641 ( \27456_27755 , RIfc6a3e8_6231, \9144_9443 );
and \U$18642 ( \27457_27756 , RIfca6898_6917, \9146_9445 );
and \U$18643 ( \27458_27757 , RIfc73358_6333, \9148_9447 );
and \U$18644 ( \27459_27758 , RIe1fd070_4256, \9150_9449 );
and \U$18645 ( \27460_27759 , RIe1fbe28_4243, \9152_9451 );
and \U$18646 ( \27461_27760 , RIfcc2660_7234, \9154_9453 );
and \U$18647 ( \27462_27761 , RIfc44468_5799, \9156_9455 );
and \U$18648 ( \27463_27762 , RIf15a940_5490, \9158_9457 );
and \U$18649 ( \27464_27763 , RIfca7270_6924, \9160_9459 );
or \U$18650 ( \27465_27764 , \27401_27700 , \27402_27701 , \27403_27702 , \27404_27703 , \27405_27704 , \27406_27705 , \27407_27706 , \27408_27707 , \27409_27708 , \27410_27709 , \27411_27710 , \27412_27711 , \27413_27712 , \27414_27713 , \27415_27714 , \27416_27715 , \27417_27716 , \27418_27717 , \27419_27718 , \27420_27719 , \27421_27720 , \27422_27721 , \27423_27722 , \27424_27723 , \27425_27724 , \27426_27725 , \27427_27726 , \27428_27727 , \27429_27728 , \27430_27729 , \27431_27730 , \27432_27731 , \27433_27732 , \27434_27733 , \27435_27734 , \27436_27735 , \27437_27736 , \27438_27737 , \27439_27738 , \27440_27739 , \27441_27740 , \27442_27741 , \27443_27742 , \27444_27743 , \27445_27744 , \27446_27745 , \27447_27746 , \27448_27747 , \27449_27748 , \27450_27749 , \27451_27750 , \27452_27751 , \27453_27752 , \27454_27753 , \27455_27754 , \27456_27755 , \27457_27756 , \27458_27757 , \27459_27758 , \27460_27759 , \27461_27760 , \27462_27761 , \27463_27762 , \27464_27763 );
and \U$18651 ( \27466_27765 , RIfc5e070_6092, \9163_9462 );
and \U$18652 ( \27467_27766 , RIfc5dda0_6090, \9165_9464 );
and \U$18653 ( \27468_27767 , RIfc7e050_6456, \9167_9466 );
and \U$18654 ( \27469_27768 , RIe1fa7a8_4227, \9169_9468 );
and \U$18655 ( \27470_27769 , RIfc5d968_6087, \9171_9470 );
and \U$18656 ( \27471_27770 , RIfcd9568_7495, \9173_9472 );
and \U$18657 ( \27472_27771 , RIfc8d668_6631, \9175_9474 );
and \U$18658 ( \27473_27772 , RIe1f5d20_4174, \9177_9476 );
and \U$18659 ( \27474_27773 , RIfca4138_6889, \9179_9478 );
and \U$18660 ( \27475_27774 , RIfc8cdf8_6625, \9181_9480 );
and \U$18661 ( \27476_27775 , RIfcc7c28_7295, \9183_9482 );
and \U$18662 ( \27477_27776 , RIe1f39f8_4149, \9185_9484 );
and \U$18663 ( \27478_27777 , RIfc99440_6766, \9187_9486 );
and \U$18664 ( \27479_27778 , RIfcbc3f0_7164, \9189_9488 );
and \U$18665 ( \27480_27779 , RIfc5a128_6047, \9191_9490 );
and \U$18666 ( \27481_27780 , RIe1ee700_4090, \9193_9492 );
and \U$18667 ( \27482_27781 , RIe1ebfa0_4062, \9195_9494 );
and \U$18668 ( \27483_27782 , RIe1e92a0_4030, \9197_9496 );
and \U$18669 ( \27484_27783 , RIe1e65a0_3998, \9199_9498 );
and \U$18670 ( \27485_27784 , RIe1e38a0_3966, \9201_9500 );
and \U$18671 ( \27486_27785 , RIe1e0ba0_3934, \9203_9502 );
and \U$18672 ( \27487_27786 , RIe1ddea0_3902, \9205_9504 );
and \U$18673 ( \27488_27787 , RIe1db1a0_3870, \9207_9506 );
and \U$18674 ( \27489_27788 , RIe1d84a0_3838, \9209_9508 );
and \U$18675 ( \27490_27789 , RIe1d2aa0_3774, \9211_9510 );
and \U$18676 ( \27491_27790 , RIe1cfda0_3742, \9213_9512 );
and \U$18677 ( \27492_27791 , RIe1cd0a0_3710, \9215_9514 );
and \U$18678 ( \27493_27792 , RIe1ca3a0_3678, \9217_9516 );
and \U$18679 ( \27494_27793 , RIe1c76a0_3646, \9219_9518 );
and \U$18680 ( \27495_27794 , RIe1c49a0_3614, \9221_9520 );
and \U$18681 ( \27496_27795 , RIe1c1ca0_3582, \9223_9522 );
and \U$18682 ( \27497_27796 , RIe1befa0_3550, \9225_9524 );
and \U$18683 ( \27498_27797 , RIf14cde0_5334, \9227_9526 );
and \U$18684 ( \27499_27798 , RIf14bb98_5321, \9229_9528 );
and \U$18685 ( \27500_27799 , RIe1b99d8_3489, \9231_9530 );
and \U$18686 ( \27501_27800 , RIe1b7980_3466, \9233_9532 );
and \U$18687 ( \27502_27801 , RIfc4c460_5890, \9235_9534 );
and \U$18688 ( \27503_27802 , RIfc9e738_6825, \9237_9536 );
and \U$18689 ( \27504_27803 , RIe1b5658_3441, \9239_9538 );
and \U$18690 ( \27505_27804 , RIfec54d8_8365, \9241_9540 );
and \U$18691 ( \27506_27805 , RIf149168_5291, \9243_9542 );
and \U$18692 ( \27507_27806 , RIf147f20_5278, \9245_9544 );
and \U$18693 ( \27508_27807 , RIe1b2ac0_3410, \9247_9546 );
and \U$18694 ( \27509_27808 , RIe1b1170_3392, \9249_9548 );
and \U$18695 ( \27510_27809 , RIf1473e0_5270, \9251_9550 );
and \U$18696 ( \27511_27810 , RIf1468a0_5262, \9253_9552 );
and \U$18697 ( \27512_27811 , RIe1acb20_3342, \9255_9554 );
and \U$18698 ( \27513_27812 , RIe1ab338_3325, \9257_9556 );
and \U$18699 ( \27514_27813 , RIe1a92e0_3302, \9259_9558 );
and \U$18700 ( \27515_27814 , RIe1a65e0_3270, \9261_9560 );
and \U$18701 ( \27516_27815 , RIe1a38e0_3238, \9263_9562 );
and \U$18702 ( \27517_27816 , RIe1a0be0_3206, \9265_9564 );
and \U$18703 ( \27518_27817 , RIe18d0e0_2982, \9267_9566 );
and \U$18704 ( \27519_27818 , RIe1795e0_2758, \9269_9568 );
and \U$18705 ( \27520_27819 , RIe226f38_4733, \9271_9570 );
and \U$18706 ( \27521_27820 , RIe21bb38_4605, \9273_9572 );
and \U$18707 ( \27522_27821 , RIe205338_4349, \9275_9574 );
and \U$18708 ( \27523_27822 , RIe1ff398_4281, \9277_9576 );
and \U$18709 ( \27524_27823 , RIe1f8750_4204, \9279_9578 );
and \U$18710 ( \27525_27824 , RIe1f1298_4121, \9281_9580 );
and \U$18711 ( \27526_27825 , RIe1d57a0_3806, \9283_9582 );
and \U$18712 ( \27527_27826 , RIe1bc2a0_3518, \9285_9584 );
and \U$18713 ( \27528_27827 , RIe1af118_3369, \9287_9586 );
and \U$18714 ( \27529_27828 , RIe171750_2668, \9289_9588 );
or \U$18715 ( \27530_27829 , \27466_27765 , \27467_27766 , \27468_27767 , \27469_27768 , \27470_27769 , \27471_27770 , \27472_27771 , \27473_27772 , \27474_27773 , \27475_27774 , \27476_27775 , \27477_27776 , \27478_27777 , \27479_27778 , \27480_27779 , \27481_27780 , \27482_27781 , \27483_27782 , \27484_27783 , \27485_27784 , \27486_27785 , \27487_27786 , \27488_27787 , \27489_27788 , \27490_27789 , \27491_27790 , \27492_27791 , \27493_27792 , \27494_27793 , \27495_27794 , \27496_27795 , \27497_27796 , \27498_27797 , \27499_27798 , \27500_27799 , \27501_27800 , \27502_27801 , \27503_27802 , \27504_27803 , \27505_27804 , \27506_27805 , \27507_27806 , \27508_27807 , \27509_27808 , \27510_27809 , \27511_27810 , \27512_27811 , \27513_27812 , \27514_27813 , \27515_27814 , \27516_27815 , \27517_27816 , \27518_27817 , \27519_27818 , \27520_27819 , \27521_27820 , \27522_27821 , \27523_27822 , \27524_27823 , \27525_27824 , \27526_27825 , \27527_27826 , \27528_27827 , \27529_27828 );
or \U$18716 ( \27531_27830 , \27465_27764 , \27530_27829 );
_DC \g3576/U$1 ( \27532 , \27531_27830 , \9298_9597 );
buf \U$18717 ( \27533_27832 , \27532 );
xor \U$18718 ( \27534_27833 , \27400_27699 , \27533_27832 );
and \U$18719 ( \27535_27834 , RIdec5ae0_713, \8760_9059 );
and \U$18720 ( \27536_27835 , RIdec2de0_681, \8762_9061 );
and \U$18721 ( \27537_27836 , RIfc82268_6503, \8764_9063 );
and \U$18722 ( \27538_27837 , RIdec00e0_649, \8766_9065 );
and \U$18723 ( \27539_27838 , RIfcb8d18_7125, \8768_9067 );
and \U$18724 ( \27540_27839 , RIdebd3e0_617, \8770_9069 );
and \U$18725 ( \27541_27840 , RIdeba6e0_585, \8772_9071 );
and \U$18726 ( \27542_27841 , RIdeb79e0_553, \8774_9073 );
and \U$18727 ( \27543_27842 , RIfcb9858_7133, \8776_9075 );
and \U$18728 ( \27544_27843 , RIdeb1fe0_489, \8778_9077 );
and \U$18729 ( \27545_27844 , RIfc9efa8_6831, \8780_9079 );
and \U$18730 ( \27546_27845 , RIdeaf2e0_457, \8782_9081 );
and \U$18731 ( \27547_27846 , RIfce0750_7576, \8784_9083 );
and \U$18732 ( \27548_27847 , RIdeab488_425, \8786_9085 );
and \U$18733 ( \27549_27848 , RIdea4b88_393, \8788_9087 );
and \U$18734 ( \27550_27849 , RIde9e288_361, \8790_9089 );
and \U$18735 ( \27551_27850 , RIee1d0b0_4789, \8792_9091 );
and \U$18736 ( \27552_27851 , RIee1c138_4778, \8794_9093 );
and \U$18737 ( \27553_27852 , RIfcd0e68_7399, \8796_9095 );
and \U$18738 ( \27554_27853 , RIfc76d00_6374, \8798_9097 );
and \U$18739 ( \27555_27854 , RIfe89028_7903, \8800_9099 );
and \U$18740 ( \27556_27855 , RIfe88d58_7901, \8802_9101 );
and \U$18741 ( \27557_27856 , RIfe88ec0_7902, \8804_9103 );
and \U$18742 ( \27558_27857 , RIfe88bf0_7900, \8806_9105 );
and \U$18743 ( \27559_27858 , RIfcda7b0_7508, \8808_9107 );
and \U$18744 ( \27560_27859 , RIfc4d810_5904, \8810_9109 );
and \U$18745 ( \27561_27860 , RIfc52dd8_5965, \8812_9111 );
and \U$18746 ( \27562_27861 , RIfcde590_7552, \8814_9113 );
and \U$18747 ( \27563_27862 , RIfc4f868_5927, \8816_9115 );
and \U$18748 ( \27564_27863 , RIe16bd50_2604, \8818_9117 );
and \U$18749 ( \27565_27864 , RIfc68930_6212, \8820_9119 );
and \U$18750 ( \27566_27865 , RIe1683a8_2563, \8822_9121 );
and \U$18751 ( \27567_27866 , RIe165ae0_2534, \8824_9123 );
and \U$18752 ( \27568_27867 , RIe162de0_2502, \8826_9125 );
and \U$18753 ( \27569_27868 , RIfe88a88_7899, \8828_9127 );
and \U$18754 ( \27570_27869 , RIe1600e0_2470, \8830_9129 );
and \U$18755 ( \27571_27870 , RIfcc9140_7310, \8832_9131 );
and \U$18756 ( \27572_27871 , RIe15d3e0_2438, \8834_9133 );
and \U$18757 ( \27573_27872 , RIe1579e0_2374, \8836_9135 );
and \U$18758 ( \27574_27873 , RIe154ce0_2342, \8838_9137 );
and \U$18759 ( \27575_27874 , RIfc698a8_6223, \8840_9139 );
and \U$18760 ( \27576_27875 , RIe151fe0_2310, \8842_9141 );
and \U$18761 ( \27577_27876 , RIee35098_5062, \8844_9143 );
and \U$18762 ( \27578_27877 , RIe14f2e0_2278, \8846_9145 );
and \U$18763 ( \27579_27878 , RIfcc0338_7209, \8848_9147 );
and \U$18764 ( \27580_27879 , RIe14c5e0_2246, \8850_9149 );
and \U$18765 ( \27581_27880 , RIe1498e0_2214, \8852_9151 );
and \U$18766 ( \27582_27881 , RIe146be0_2182, \8854_9153 );
and \U$18767 ( \27583_27882 , RIfc88208_6571, \8856_9155 );
and \U$18768 ( \27584_27883 , RIfc85670_6540, \8858_9157 );
and \U$18769 ( \27585_27884 , RIfc81f98_6501, \8860_9159 );
and \U$18770 ( \27586_27885 , RIfcc4f28_7263, \8862_9161 );
and \U$18771 ( \27587_27886 , RIe1414b0_2120, \8864_9163 );
and \U$18772 ( \27588_27887 , RIe13f188_2095, \8866_9165 );
and \U$18773 ( \27589_27888 , RIdf3d090_2071, \8868_9167 );
and \U$18774 ( \27590_27889 , RIdf3aa98_2044, \8870_9169 );
and \U$18775 ( \27591_27890 , RIfcd2920_7418, \8872_9171 );
and \U$18776 ( \27592_27891 , RIfc7d7e0_6450, \8874_9173 );
and \U$18777 ( \27593_27892 , RIfc49760_5858, \8876_9175 );
and \U$18778 ( \27594_27893 , RIfce5a48_7635, \8878_9177 );
and \U$18779 ( \27595_27894 , RIdf35ea8_1990, \8880_9179 );
and \U$18780 ( \27596_27895 , RIdf338b0_1963, \8882_9181 );
and \U$18781 ( \27597_27896 , RIfe88920_7898, \8884_9183 );
and \U$18782 ( \27598_27897 , RIdf2f800_1917, \8886_9185 );
or \U$18783 ( \27599_27898 , \27535_27834 , \27536_27835 , \27537_27836 , \27538_27837 , \27539_27838 , \27540_27839 , \27541_27840 , \27542_27841 , \27543_27842 , \27544_27843 , \27545_27844 , \27546_27845 , \27547_27846 , \27548_27847 , \27549_27848 , \27550_27849 , \27551_27850 , \27552_27851 , \27553_27852 , \27554_27853 , \27555_27854 , \27556_27855 , \27557_27856 , \27558_27857 , \27559_27858 , \27560_27859 , \27561_27860 , \27562_27861 , \27563_27862 , \27564_27863 , \27565_27864 , \27566_27865 , \27567_27866 , \27568_27867 , \27569_27868 , \27570_27869 , \27571_27870 , \27572_27871 , \27573_27872 , \27574_27873 , \27575_27874 , \27576_27875 , \27577_27876 , \27578_27877 , \27579_27878 , \27580_27879 , \27581_27880 , \27582_27881 , \27583_27882 , \27584_27883 , \27585_27884 , \27586_27885 , \27587_27886 , \27588_27887 , \27589_27888 , \27590_27889 , \27591_27890 , \27592_27891 , \27593_27892 , \27594_27893 , \27595_27894 , \27596_27895 , \27597_27896 , \27598_27897 );
and \U$18784 ( \27600_27899 , RIee2bfc0_4959, \8889_9188 );
and \U$18785 ( \27601_27900 , RIee2a670_4941, \8891_9190 );
and \U$18786 ( \27602_27901 , RIee29158_4926, \8893_9192 );
and \U$18787 ( \27603_27902 , RIee27f10_4913, \8895_9194 );
and \U$18788 ( \27604_27903 , RIdf2a7d8_1860, \8897_9196 );
and \U$18789 ( \27605_27904 , RIdf28618_1836, \8899_9198 );
and \U$18790 ( \27606_27905 , RIdf26890_1815, \8901_9200 );
and \U$18791 ( \27607_27906 , RIdf24dd8_1796, \8903_9202 );
and \U$18792 ( \27608_27907 , RIfcad918_6997, \8905_9204 );
and \U$18793 ( \27609_27908 , RIfc69fb0_6228, \8907_9206 );
and \U$18794 ( \27610_27909 , RIfc63368_6151, \8909_9208 );
and \U$18795 ( \27611_27910 , RIfc623f0_6140, \8911_9210 );
and \U$18796 ( \27612_27911 , RIfc60938_6121, \8913_9212 );
and \U$18797 ( \27613_27912 , RIdf1ff18_1740, \8915_9214 );
and \U$18798 ( \27614_27913 , RIfcba500_7142, \8917_9216 );
and \U$18799 ( \27615_27914 , RIdf19870_1667, \8919_9218 );
and \U$18800 ( \27616_27915 , RIdf176b0_1643, \8921_9220 );
and \U$18801 ( \27617_27916 , RIdf149b0_1611, \8923_9222 );
and \U$18802 ( \27618_27917 , RIdf11cb0_1579, \8925_9224 );
and \U$18803 ( \27619_27918 , RIdf0efb0_1547, \8927_9226 );
and \U$18804 ( \27620_27919 , RIdf0c2b0_1515, \8929_9228 );
and \U$18805 ( \27621_27920 , RIdf095b0_1483, \8931_9230 );
and \U$18806 ( \27622_27921 , RIdf068b0_1451, \8933_9232 );
and \U$18807 ( \27623_27922 , RIdf03bb0_1419, \8935_9234 );
and \U$18808 ( \27624_27923 , RIdefe1b0_1355, \8937_9236 );
and \U$18809 ( \27625_27924 , RIdefb4b0_1323, \8939_9238 );
and \U$18810 ( \27626_27925 , RIdef87b0_1291, \8941_9240 );
and \U$18811 ( \27627_27926 , RIdef5ab0_1259, \8943_9242 );
and \U$18812 ( \27628_27927 , RIdef2db0_1227, \8945_9244 );
and \U$18813 ( \27629_27928 , RIdef00b0_1195, \8947_9246 );
and \U$18814 ( \27630_27929 , RIdeed3b0_1163, \8949_9248 );
and \U$18815 ( \27631_27930 , RIdeea6b0_1131, \8951_9250 );
and \U$18816 ( \27632_27931 , RIfcc9848_7315, \8953_9252 );
and \U$18817 ( \27633_27932 , RIfc69a10_6224, \8955_9254 );
and \U$18818 ( \27634_27933 , RIfcacc70_6988, \8957_9256 );
and \U$18819 ( \27635_27934 , RIfccbfa8_7343, \8959_9258 );
and \U$18820 ( \27636_27935 , RIdee4f80_1069, \8961_9260 );
and \U$18821 ( \27637_27936 , RIdee31f8_1048, \8963_9262 );
and \U$18822 ( \27638_27937 , RIdee1038_1024, \8965_9264 );
and \U$18823 ( \27639_27938 , RIdedee78_1000, \8967_9266 );
and \U$18824 ( \27640_27939 , RIfc84590_6528, \8969_9268 );
and \U$18825 ( \27641_27940 , RIfc9bba0_6794, \8971_9270 );
and \U$18826 ( \27642_27941 , RIee21b38_4842, \8973_9272 );
and \U$18827 ( \27643_27942 , RIfc47168_5831, \8975_9274 );
and \U$18828 ( \27644_27943 , RIded9e50_943, \8977_9276 );
and \U$18829 ( \27645_27944 , RIded7858_916, \8979_9278 );
and \U$18830 ( \27646_27945 , RIfe887b8_7897, \8981_9280 );
and \U$18831 ( \27647_27946 , RIded34d8_868, \8983_9282 );
and \U$18832 ( \27648_27947 , RIded0ee0_841, \8985_9284 );
and \U$18833 ( \27649_27948 , RIdece1e0_809, \8987_9286 );
and \U$18834 ( \27650_27949 , RIdecb4e0_777, \8989_9288 );
and \U$18835 ( \27651_27950 , RIdec87e0_745, \8991_9290 );
and \U$18836 ( \27652_27951 , RIdeb4ce0_521, \8993_9292 );
and \U$18837 ( \27653_27952 , RIde97988_329, \8995_9294 );
and \U$18838 ( \27654_27953 , RIe16e8e8_2635, \8997_9296 );
and \U$18839 ( \27655_27954 , RIe15a6e0_2406, \8999_9298 );
and \U$18840 ( \27656_27955 , RIe143ee0_2150, \9001_9300 );
and \U$18841 ( \27657_27956 , RIdf388d8_2020, \9003_9302 );
and \U$18842 ( \27658_27957 , RIdf2cf38_1888, \9005_9304 );
and \U$18843 ( \27659_27958 , RIdf1d7b8_1712, \9007_9306 );
and \U$18844 ( \27660_27959 , RIdf00eb0_1387, \9009_9308 );
and \U$18845 ( \27661_27960 , RIdee79b0_1099, \9011_9310 );
and \U$18846 ( \27662_27961 , RIdedc718_972, \9013_9312 );
and \U$18847 ( \27663_27962 , RIde7d8d0_202, \9015_9314 );
or \U$18848 ( \27664_27963 , \27600_27899 , \27601_27900 , \27602_27901 , \27603_27902 , \27604_27903 , \27605_27904 , \27606_27905 , \27607_27906 , \27608_27907 , \27609_27908 , \27610_27909 , \27611_27910 , \27612_27911 , \27613_27912 , \27614_27913 , \27615_27914 , \27616_27915 , \27617_27916 , \27618_27917 , \27619_27918 , \27620_27919 , \27621_27920 , \27622_27921 , \27623_27922 , \27624_27923 , \27625_27924 , \27626_27925 , \27627_27926 , \27628_27927 , \27629_27928 , \27630_27929 , \27631_27930 , \27632_27931 , \27633_27932 , \27634_27933 , \27635_27934 , \27636_27935 , \27637_27936 , \27638_27937 , \27639_27938 , \27640_27939 , \27641_27940 , \27642_27941 , \27643_27942 , \27644_27943 , \27645_27944 , \27646_27945 , \27647_27946 , \27648_27947 , \27649_27948 , \27650_27949 , \27651_27950 , \27652_27951 , \27653_27952 , \27654_27953 , \27655_27954 , \27656_27955 , \27657_27956 , \27658_27957 , \27659_27958 , \27660_27959 , \27661_27960 , \27662_27961 , \27663_27962 );
or \U$18849 ( \27665_27964 , \27599_27898 , \27664_27963 );
_DC \g24ce/U$1 ( \27666 , \27665_27964 , \9024_9323 );
buf \U$18850 ( \27667_27966 , \27666 );
and \U$18851 ( \27668_27967 , RIe19dd78_3173, \9034_9333 );
and \U$18852 ( \27669_27968 , RIe19b078_3141, \9036_9335 );
and \U$18853 ( \27670_27969 , RIfca1438_6857, \9038_9337 );
and \U$18854 ( \27671_27970 , RIe198378_3109, \9040_9339 );
and \U$18855 ( \27672_27971 , RIfca35f8_6881, \9042_9341 );
and \U$18856 ( \27673_27972 , RIe195678_3077, \9044_9343 );
and \U$18857 ( \27674_27973 , RIe192978_3045, \9046_9345 );
and \U$18858 ( \27675_27974 , RIe18fc78_3013, \9048_9347 );
and \U$18859 ( \27676_27975 , RIe18a278_2949, \9050_9349 );
and \U$18860 ( \27677_27976 , RIe187578_2917, \9052_9351 );
and \U$18861 ( \27678_27977 , RIfcba230_7140, \9054_9353 );
and \U$18862 ( \27679_27978 , RIe184878_2885, \9056_9355 );
and \U$18863 ( \27680_27979 , RIf142d90_5220, \9058_9357 );
and \U$18864 ( \27681_27980 , RIe181b78_2853, \9060_9359 );
and \U$18865 ( \27682_27981 , RIe17ee78_2821, \9062_9361 );
and \U$18866 ( \27683_27982 , RIe17c178_2789, \9064_9363 );
and \U$18867 ( \27684_27983 , RIfc9be70_6796, \9066_9365 );
and \U$18868 ( \27685_27984 , RIfc9bd08_6795, \9068_9367 );
and \U$18869 ( \27686_27985 , RIfc4ccd0_5896, \9070_9369 );
and \U$18870 ( \27687_27986 , RIe176070_2720, \9072_9371 );
and \U$18871 ( \27688_27987 , RIfc87c68_6567, \9074_9373 );
and \U$18872 ( \27689_27988 , RIfc87b00_6566, \9076_9375 );
and \U$18873 ( \27690_27989 , RIfcc4c58_7261, \9078_9377 );
and \U$18874 ( \27691_27990 , RIfc4fca0_5930, \9080_9379 );
and \U$18875 ( \27692_27991 , RIfc4f598_5925, \9082_9381 );
and \U$18876 ( \27693_27992 , RIfc876c8_6563, \9084_9383 );
and \U$18877 ( \27694_27993 , RIfc4dae0_5906, \9086_9385 );
and \U$18878 ( \27695_27994 , RIe173eb0_2696, \9088_9387 );
and \U$18879 ( \27696_27995 , RIfcb9420_7130, \9090_9389 );
and \U$18880 ( \27697_27996 , RIfc4e080_5910, \9092_9391 );
and \U$18881 ( \27698_27997 , RIfc4e350_5912, \9094_9393 );
and \U$18882 ( \27699_27998 , RIfc9d388_6811, \9096_9395 );
and \U$18883 ( \27700_27999 , RIfc40a48_5761, \9098_9397 );
and \U$18884 ( \27701_28000 , RIe2240d0_4700, \9100_9399 );
and \U$18885 ( \27702_28001 , RIfc85508_6539, \9102_9401 );
and \U$18886 ( \27703_28002 , RIe2213d0_4668, \9104_9403 );
and \U$18887 ( \27704_28003 , RIfc9ba38_6793, \9106_9405 );
and \U$18888 ( \27705_28004 , RIe21e6d0_4636, \9108_9407 );
and \U$18889 ( \27706_28005 , RIe218cd0_4572, \9110_9409 );
and \U$18890 ( \27707_28006 , RIe215fd0_4540, \9112_9411 );
and \U$18891 ( \27708_28007 , RIfc52c70_5964, \9114_9413 );
and \U$18892 ( \27709_28008 , RIe2132d0_4508, \9116_9415 );
and \U$18893 ( \27710_28009 , RIfca3760_6882, \9118_9417 );
and \U$18894 ( \27711_28010 , RIe2105d0_4476, \9120_9419 );
and \U$18895 ( \27712_28011 , RIfc97988_6747, \9122_9421 );
and \U$18896 ( \27713_28012 , RIe20d8d0_4444, \9124_9423 );
and \U$18897 ( \27714_28013 , RIe20abd0_4412, \9126_9425 );
and \U$18898 ( \27715_28014 , RIe207ed0_4380, \9128_9427 );
and \U$18899 ( \27716_28015 , RIfceb5b0_7700, \9130_9429 );
and \U$18900 ( \27717_28016 , RIfcddbb8_7545, \9132_9431 );
and \U$18901 ( \27718_28017 , RIe202a70_4320, \9134_9433 );
and \U$18902 ( \27719_28018 , RIe200e50_4300, \9136_9435 );
and \U$18903 ( \27720_28019 , RIfc73d30_6340, \9138_9437 );
and \U$18904 ( \27721_28020 , RIfcaf100_7014, \9140_9439 );
and \U$18905 ( \27722_28021 , RIfc71468_6311, \9142_9441 );
and \U$18906 ( \27723_28022 , RIfcdcad8_7533, \9144_9443 );
and \U$18907 ( \27724_28023 , RIfcdda50_7544, \9146_9445 );
and \U$18908 ( \27725_28024 , RIfca8620_6938, \9148_9447 );
and \U$18909 ( \27726_28025 , RIe1fcf08_4255, \9150_9449 );
and \U$18910 ( \27727_28026 , RIe1fbcc0_4242, \9152_9451 );
and \U$18911 ( \27728_28027 , RIfc6c008_6251, \9154_9453 );
and \U$18912 ( \27729_28028 , RIfcdd1e0_7538, \9156_9455 );
and \U$18913 ( \27730_28029 , RIfca9700_6950, \9158_9457 );
and \U$18914 ( \27731_28030 , RIfca92c8_6947, \9160_9459 );
or \U$18915 ( \27732_28031 , \27668_27967 , \27669_27968 , \27670_27969 , \27671_27970 , \27672_27971 , \27673_27972 , \27674_27973 , \27675_27974 , \27676_27975 , \27677_27976 , \27678_27977 , \27679_27978 , \27680_27979 , \27681_27980 , \27682_27981 , \27683_27982 , \27684_27983 , \27685_27984 , \27686_27985 , \27687_27986 , \27688_27987 , \27689_27988 , \27690_27989 , \27691_27990 , \27692_27991 , \27693_27992 , \27694_27993 , \27695_27994 , \27696_27995 , \27697_27996 , \27698_27997 , \27699_27998 , \27700_27999 , \27701_28000 , \27702_28001 , \27703_28002 , \27704_28003 , \27705_28004 , \27706_28005 , \27707_28006 , \27708_28007 , \27709_28008 , \27710_28009 , \27711_28010 , \27712_28011 , \27713_28012 , \27714_28013 , \27715_28014 , \27716_28015 , \27717_28016 , \27718_28017 , \27719_28018 , \27720_28019 , \27721_28020 , \27722_28021 , \27723_28022 , \27724_28023 , \27725_28024 , \27726_28025 , \27727_28026 , \27728_28027 , \27729_28028 , \27730_28029 , \27731_28030 );
and \U$18916 ( \27733_28032 , RIfcce5a0_7370, \9163_9462 );
and \U$18917 ( \27734_28033 , RIfc6ba68_6247, \9165_9464 );
and \U$18918 ( \27735_28034 , RIfc6f410_6288, \9167_9466 );
and \U$18919 ( \27736_28035 , RIe1fa640_4226, \9169_9468 );
and \U$18920 ( \27737_28036 , RIfcce000_7366, \9171_9470 );
and \U$18921 ( \27738_28037 , RIfc53918_5973, \9173_9472 );
and \U$18922 ( \27739_28038 , RIfcce708_7371, \9175_9474 );
and \U$18923 ( \27740_28039 , RIe1f5bb8_4173, \9177_9476 );
and \U$18924 ( \27741_28040 , RIf1535f0_5408, \9179_9478 );
and \U$18925 ( \27742_28041 , RIf151e08_5391, \9181_9480 );
and \U$18926 ( \27743_28042 , RIfc72db8_6329, \9183_9482 );
and \U$18927 ( \27744_28043 , RIe1f3890_4148, \9185_9484 );
and \U$18928 ( \27745_28044 , RIf14fc48_5367, \9187_9486 );
and \U$18929 ( \27746_28045 , RIfc72c50_6328, \9189_9488 );
and \U$18930 ( \27747_28046 , RIfc73e98_6341, \9191_9490 );
and \U$18931 ( \27748_28047 , RIe1ee598_4089, \9193_9492 );
and \U$18932 ( \27749_28048 , RIe1ebe38_4061, \9195_9494 );
and \U$18933 ( \27750_28049 , RIe1e9138_4029, \9197_9496 );
and \U$18934 ( \27751_28050 , RIe1e6438_3997, \9199_9498 );
and \U$18935 ( \27752_28051 , RIe1e3738_3965, \9201_9500 );
and \U$18936 ( \27753_28052 , RIe1e0a38_3933, \9203_9502 );
and \U$18937 ( \27754_28053 , RIe1ddd38_3901, \9205_9504 );
and \U$18938 ( \27755_28054 , RIe1db038_3869, \9207_9506 );
and \U$18939 ( \27756_28055 , RIe1d8338_3837, \9209_9508 );
and \U$18940 ( \27757_28056 , RIe1d2938_3773, \9211_9510 );
and \U$18941 ( \27758_28057 , RIe1cfc38_3741, \9213_9512 );
and \U$18942 ( \27759_28058 , RIe1ccf38_3709, \9215_9514 );
and \U$18943 ( \27760_28059 , RIe1ca238_3677, \9217_9516 );
and \U$18944 ( \27761_28060 , RIe1c7538_3645, \9219_9518 );
and \U$18945 ( \27762_28061 , RIe1c4838_3613, \9221_9520 );
and \U$18946 ( \27763_28062 , RIe1c1b38_3581, \9223_9522 );
and \U$18947 ( \27764_28063 , RIe1bee38_3549, \9225_9524 );
and \U$18948 ( \27765_28064 , RIfcb8a48_7123, \9227_9526 );
and \U$18949 ( \27766_28065 , RIfcb84a8_7119, \9229_9528 );
and \U$18950 ( \27767_28066 , RIe1b9870_3488, \9231_9530 );
and \U$18951 ( \27768_28067 , RIe1b7818_3465, \9233_9532 );
and \U$18952 ( \27769_28068 , RIfc85940_6542, \9235_9534 );
and \U$18953 ( \27770_28069 , RIfc9e198_6821, \9237_9536 );
and \U$18954 ( \27771_28070 , RIfeac140_8274, \9239_9538 );
and \U$18955 ( \27772_28071 , RIe1b42a8_3427, \9241_9540 );
and \U$18956 ( \27773_28072 , RIfc518c0_5950, \9243_9542 );
and \U$18957 ( \27774_28073 , RIfc838e8_6519, \9245_9544 );
and \U$18958 ( \27775_28074 , RIfe884e8_7895, \9247_9546 );
and \U$18959 ( \27776_28075 , RIe1b1008_3391, \9249_9548 );
and \U$18960 ( \27777_28076 , RIfcc5900_7270, \9251_9550 );
and \U$18961 ( \27778_28077 , RIfc82ad8_6509, \9253_9552 );
and \U$18962 ( \27779_28078 , RIe1ac9b8_3341, \9255_9554 );
and \U$18963 ( \27780_28079 , RIfe88650_7896, \9257_9556 );
and \U$18964 ( \27781_28080 , RIe1a9178_3301, \9259_9558 );
and \U$18965 ( \27782_28081 , RIe1a6478_3269, \9261_9560 );
and \U$18966 ( \27783_28082 , RIe1a3778_3237, \9263_9562 );
and \U$18967 ( \27784_28083 , RIe1a0a78_3205, \9265_9564 );
and \U$18968 ( \27785_28084 , RIe18cf78_2981, \9267_9566 );
and \U$18969 ( \27786_28085 , RIe179478_2757, \9269_9568 );
and \U$18970 ( \27787_28086 , RIe226dd0_4732, \9271_9570 );
and \U$18971 ( \27788_28087 , RIe21b9d0_4604, \9273_9572 );
and \U$18972 ( \27789_28088 , RIe2051d0_4348, \9275_9574 );
and \U$18973 ( \27790_28089 , RIe1ff230_4280, \9277_9576 );
and \U$18974 ( \27791_28090 , RIe1f85e8_4203, \9279_9578 );
and \U$18975 ( \27792_28091 , RIe1f1130_4120, \9281_9580 );
and \U$18976 ( \27793_28092 , RIe1d5638_3805, \9283_9582 );
and \U$18977 ( \27794_28093 , RIe1bc138_3517, \9285_9584 );
and \U$18978 ( \27795_28094 , RIe1aefb0_3368, \9287_9586 );
and \U$18979 ( \27796_28095 , RIe1715e8_2667, \9289_9588 );
or \U$18980 ( \27797_28096 , \27733_28032 , \27734_28033 , \27735_28034 , \27736_28035 , \27737_28036 , \27738_28037 , \27739_28038 , \27740_28039 , \27741_28040 , \27742_28041 , \27743_28042 , \27744_28043 , \27745_28044 , \27746_28045 , \27747_28046 , \27748_28047 , \27749_28048 , \27750_28049 , \27751_28050 , \27752_28051 , \27753_28052 , \27754_28053 , \27755_28054 , \27756_28055 , \27757_28056 , \27758_28057 , \27759_28058 , \27760_28059 , \27761_28060 , \27762_28061 , \27763_28062 , \27764_28063 , \27765_28064 , \27766_28065 , \27767_28066 , \27768_28067 , \27769_28068 , \27770_28069 , \27771_28070 , \27772_28071 , \27773_28072 , \27774_28073 , \27775_28074 , \27776_28075 , \27777_28076 , \27778_28077 , \27779_28078 , \27780_28079 , \27781_28080 , \27782_28081 , \27783_28082 , \27784_28083 , \27785_28084 , \27786_28085 , \27787_28086 , \27788_28087 , \27789_28088 , \27790_28089 , \27791_28090 , \27792_28091 , \27793_28092 , \27794_28093 , \27795_28094 , \27796_28095 );
or \U$18981 ( \27798_28097 , \27732_28031 , \27797_28096 );
_DC \g35fb/U$1 ( \27799 , \27798_28097 , \9298_9597 );
buf \U$18982 ( \27800_28099 , \27799 );
and \U$18983 ( \27801_28100 , \27667_27966 , \27800_28099 );
and \U$18984 ( \27802_28101 , \25713_26012 , \25846_26145 );
and \U$18985 ( \27803_28102 , \25846_26145 , \26121_26420 );
and \U$18986 ( \27804_28103 , \25713_26012 , \26121_26420 );
or \U$18987 ( \27805_28104 , \27802_28101 , \27803_28102 , \27804_28103 );
and \U$18988 ( \27806_28105 , \27800_28099 , \27805_28104 );
and \U$18989 ( \27807_28106 , \27667_27966 , \27805_28104 );
or \U$18990 ( \27808_28107 , \27801_28100 , \27806_28105 , \27807_28106 );
xor \U$18991 ( \27809_28108 , \27534_27833 , \27808_28107 );
buf g4406_GF_PartitionCandidate( \27810_28109_nG4406 , \27809_28108 );
xor \U$18992 ( \27811_28110 , \27667_27966 , \27800_28099 );
xor \U$18993 ( \27812_28111 , \27811_28110 , \27805_28104 );
buf g4409_GF_PartitionCandidate( \27813_28112_nG4409 , \27812_28111 );
nand \U$18994 ( \27814_28113 , \27813_28112_nG4409 , \26123_26422_nG440c );
and \U$18995 ( \27815_28114 , \27810_28109_nG4406 , \27814_28113 );
xor \U$18996 ( \27816_28115 , \27813_28112_nG4409 , \26123_26422_nG440c );
and \U$19001 ( \27817_28119 , \27816_28115 , \10392_10694_nG9c0e );
or \U$19002 ( \27818_28120 , 1'b0 , \27817_28119 );
xor \U$19003 ( \27819_28121 , \27815_28114 , \27818_28120 );
xor \U$19004 ( \27820_28122 , \27815_28114 , \27819_28121 );
buf \U$19005 ( \27821_28123 , \27820_28122 );
buf \U$19006 ( \27822_28124 , \27821_28123 );
xor \U$19007 ( \27823_28125 , \27267_27566 , \27822_28124 );
and \U$19008 ( \27824_28126 , \27222_27521 , \27227_27526 );
and \U$19009 ( \27825_28127 , \27222_27521 , \27260_27559 );
and \U$19010 ( \27826_28128 , \27227_27526 , \27260_27559 );
or \U$19011 ( \27827_28129 , \27824_28126 , \27825_28127 , \27826_28128 );
and \U$19012 ( \27828_28130 , \27823_28125 , \27827_28129 );
and \U$19013 ( \27829_28131 , \27233_27532 , \27252_27551 );
and \U$19014 ( \27830_28132 , \27233_27532 , \27258_27557 );
and \U$19015 ( \27831_28133 , \27252_27551 , \27258_27557 );
or \U$19016 ( \27832_28134 , \27829_28131 , \27830_28132 , \27831_28133 );
buf \U$19017 ( \27833_28135 , \27832_28134 );
and \U$19018 ( \27834_28136 , \27197_27496 , \27202_27501 );
and \U$19019 ( \27835_28137 , \27197_27496 , \27209_27508 );
and \U$19020 ( \27836_28138 , \27202_27501 , \27209_27508 );
or \U$19021 ( \27837_28139 , \27834_28136 , \27835_28137 , \27836_28138 );
buf \U$19022 ( \27838_28140 , \27837_28139 );
and \U$19023 ( \27839_28141 , \13431_13370 , \22330_22629_nG9bd5 );
and \U$19024 ( \27840_28142 , \13068_13367 , \23394_23696_nG9bd2 );
or \U$19025 ( \27841_28143 , \27839_28141 , \27840_28142 );
xor \U$19026 ( \27842_28144 , \13067_13366 , \27841_28143 );
buf \U$19027 ( \27843_28145 , \27842_28144 );
buf \U$19029 ( \27844_28146 , \27843_28145 );
xor \U$19030 ( \27845_28147 , \27838_28140 , \27844_28146 );
and \U$19031 ( \27846_28148 , \12183_12157 , \23927_24226_nG9bcf );
and \U$19032 ( \27847_28149 , \11855_12154 , \24996_25298_nG9bcc );
or \U$19033 ( \27848_28150 , \27846_28148 , \27847_28149 );
xor \U$19034 ( \27849_28151 , \11854_12153 , \27848_28150 );
buf \U$19035 ( \27850_28152 , \27849_28151 );
buf \U$19037 ( \27851_28153 , \27850_28152 );
xor \U$19038 ( \27852_28154 , \27845_28147 , \27851_28153 );
buf \U$19039 ( \27853_28155 , \27852_28154 );
and \U$19040 ( \27854_28156 , \27130_27432 , \27136_27438 );
buf \U$19041 ( \27855_28157 , \27854_28156 );
and \U$19042 ( \27856_28158 , \23495_23201 , \12502_12801_nG9bff );
and \U$19043 ( \27857_28159 , \22899_23198 , \13403_13705_nG9bfc );
or \U$19044 ( \27858_28160 , \27856_28158 , \27857_28159 );
xor \U$19045 ( \27859_28161 , \22898_23197 , \27858_28160 );
buf \U$19046 ( \27860_28162 , \27859_28161 );
buf \U$19048 ( \27861_28163 , \27860_28162 );
xor \U$19049 ( \27862_28164 , \27855_28157 , \27861_28163 );
and \U$19050 ( \27863_28165 , \21908_21658 , \13771_14070_nG9bf9 );
and \U$19051 ( \27864_28166 , \21356_21655 , \14682_14984_nG9bf6 );
or \U$19052 ( \27865_28167 , \27863_28165 , \27864_28166 );
xor \U$19053 ( \27866_28168 , \21355_21654 , \27865_28167 );
buf \U$19054 ( \27867_28169 , \27866_28168 );
buf \U$19056 ( \27868_28170 , \27867_28169 );
xor \U$19057 ( \27869_28171 , \27862_28164 , \27868_28170 );
buf \U$19058 ( \27870_28172 , \27869_28171 );
and \U$19059 ( \27871_28173 , \18908_18702 , \16378_16680_nG9bed );
and \U$19060 ( \27872_28174 , \18400_18699 , \17363_17665_nG9bea );
or \U$19061 ( \27873_28175 , \27871_28173 , \27872_28174 );
xor \U$19062 ( \27874_28176 , \18399_18698 , \27873_28175 );
buf \U$19063 ( \27875_28177 , \27874_28176 );
buf \U$19065 ( \27876_28178 , \27875_28177 );
xor \U$19066 ( \27877_28179 , \27870_28172 , \27876_28178 );
and \U$19067 ( \27878_28180 , \17437_17297 , \17808_18107_nG9be7 );
and \U$19068 ( \27879_28181 , \16995_17294 , \18789_19091_nG9be4 );
or \U$19069 ( \27880_28182 , \27878_28180 , \27879_28181 );
xor \U$19070 ( \27881_28183 , \16994_17293 , \27880_28182 );
buf \U$19071 ( \27882_28184 , \27881_28183 );
buf \U$19073 ( \27883_28185 , \27882_28184 );
xor \U$19074 ( \27884_28186 , \27877_28179 , \27883_28185 );
buf \U$19075 ( \27885_28187 , \27884_28186 );
and \U$19076 ( \27886_28188 , \27127_27429 , \27156_27455 );
and \U$19077 ( \27887_28189 , \27127_27429 , \27163_27462 );
and \U$19078 ( \27888_28190 , \27156_27455 , \27163_27462 );
or \U$19079 ( \27889_28191 , \27886_28188 , \27887_28189 , \27888_28190 );
buf \U$19080 ( \27890_28192 , \27889_28191 );
xor \U$19081 ( \27891_28193 , \27885_28187 , \27890_28192 );
and \U$19082 ( \27892_28194 , \16405_15940 , \19287_19586_nG9be1 );
and \U$19083 ( \27893_28195 , \15638_15937 , \20306_20608_nG9bde );
or \U$19084 ( \27894_28196 , \27892_28194 , \27893_28195 );
xor \U$19085 ( \27895_28197 , \15637_15936 , \27894_28196 );
buf \U$19086 ( \27896_28198 , \27895_28197 );
buf \U$19088 ( \27897_28199 , \27896_28198 );
xor \U$19089 ( \27898_28200 , \27891_28193 , \27897_28199 );
buf \U$19090 ( \27899_28201 , \27898_28200 );
xor \U$19091 ( \27900_28202 , \27853_28155 , \27899_28201 );
and \U$19092 ( \27901_28203 , \10411_10707 , \27114_27416_nG9bc3 );
and \U$19093 ( \27902_28204 , \27060_27362 , \27064_27366 );
and \U$19094 ( \27903_28205 , \27064_27366 , \27102_27404 );
and \U$19095 ( \27904_28206 , \27060_27362 , \27102_27404 );
or \U$19096 ( \27905_28207 , \27902_28204 , \27903_28205 , \27904_28206 );
and \U$19097 ( \27906_28208 , \27069_27371 , \27073_27375 );
and \U$19098 ( \27907_28209 , \27073_27375 , \27101_27403 );
and \U$19099 ( \27908_28210 , \27069_27371 , \27101_27403 );
or \U$19100 ( \27909_28211 , \27906_28208 , \27907_28209 , \27908_28210 );
and \U$19101 ( \27910_28212 , \26719_27021 , \27005_27307 );
and \U$19102 ( \27911_28213 , \27005_27307 , \27054_27356 );
and \U$19103 ( \27912_28214 , \26719_27021 , \27054_27356 );
or \U$19104 ( \27913_28215 , \27910_28212 , \27911_28213 , \27912_28214 );
xor \U$19105 ( \27914_28216 , \27909_28211 , \27913_28215 );
and \U$19106 ( \27915_28217 , \26995_27297 , \26999_27301 );
and \U$19107 ( \27916_28218 , \26999_27301 , \27004_27306 );
and \U$19108 ( \27917_28219 , \26995_27297 , \27004_27306 );
or \U$19109 ( \27918_28220 , \27915_28217 , \27916_28218 , \27917_28219 );
and \U$19110 ( \27919_28221 , \27078_27380 , \27082_27384 );
and \U$19111 ( \27920_28222 , \27082_27384 , \27100_27402 );
and \U$19112 ( \27921_28223 , \27078_27380 , \27100_27402 );
or \U$19113 ( \27922_28224 , \27919_28221 , \27920_28222 , \27921_28223 );
xor \U$19114 ( \27923_28225 , \27918_28220 , \27922_28224 );
and \U$19115 ( \27924_28226 , \27024_27326 , \27038_27340 );
and \U$19116 ( \27925_28227 , \27038_27340 , \27053_27355 );
and \U$19117 ( \27926_28228 , \27024_27326 , \27053_27355 );
or \U$19118 ( \27927_28229 , \27924_28226 , \27925_28227 , \27926_28228 );
xor \U$19119 ( \27928_28230 , \27923_28225 , \27927_28229 );
xor \U$19120 ( \27929_28231 , \27914_28216 , \27928_28230 );
xor \U$19121 ( \27930_28232 , \27905_28207 , \27929_28231 );
and \U$19122 ( \27931_28233 , \27014_27316 , \27018_27320 );
and \U$19123 ( \27932_28234 , \27018_27320 , \27023_27325 );
and \U$19124 ( \27933_28235 , \27014_27316 , \27023_27325 );
or \U$19125 ( \27934_28236 , \27931_28233 , \27932_28234 , \27933_28235 );
and \U$19126 ( \27935_28237 , \27028_27330 , \27032_27334 );
and \U$19127 ( \27936_28238 , \27032_27334 , \27037_27339 );
and \U$19128 ( \27937_28239 , \27028_27330 , \27037_27339 );
or \U$19129 ( \27938_28240 , \27935_28237 , \27936_28238 , \27937_28239 );
xor \U$19130 ( \27939_28241 , \27934_28236 , \27938_28240 );
and \U$19131 ( \27940_28242 , \27043_27345 , \27047_27349 );
and \U$19132 ( \27941_28243 , \27047_27349 , \27052_27354 );
and \U$19133 ( \27942_28244 , \27043_27345 , \27052_27354 );
or \U$19134 ( \27943_28245 , \27940_28242 , \27941_28243 , \27942_28244 );
xor \U$19135 ( \27944_28246 , \27939_28241 , \27943_28245 );
and \U$19136 ( \27945_28247 , \27087_27389 , \27091_27393 );
and \U$19137 ( \27946_28248 , \27091_27393 , \27099_27401 );
and \U$19138 ( \27947_28249 , \27087_27389 , \27099_27401 );
or \U$19139 ( \27948_28250 , \27945_28247 , \27946_28248 , \27947_28249 );
and \U$19140 ( \27949_28251 , \25516_25815 , \11275_11574 );
and \U$19141 ( \27950_28252 , \26527_26829 , \10976_11278 );
nor \U$19142 ( \27951_28253 , \27949_28251 , \27950_28252 );
xnor \U$19143 ( \27952_28254 , \27951_28253 , \11281_11580 );
and \U$19144 ( \27953_28255 , \22257_22556 , \13755_14054 );
and \U$19145 ( \27954_28256 , \23315_23617 , \13390_13692 );
nor \U$19146 ( \27955_28257 , \27953_28255 , \27954_28256 );
xnor \U$19147 ( \27956_28258 , \27955_28257 , \13736_14035 );
xor \U$19148 ( \27957_28259 , \27952_28254 , \27956_28258 );
and \U$19149 ( \27958_28260 , RIdec5ae0_713, \9034_9333 );
and \U$19150 ( \27959_28261 , RIdec2de0_681, \9036_9335 );
and \U$19151 ( \27960_28262 , RIfc82268_6503, \9038_9337 );
and \U$19152 ( \27961_28263 , RIdec00e0_649, \9040_9339 );
and \U$19153 ( \27962_28264 , RIfcb8d18_7125, \9042_9341 );
and \U$19154 ( \27963_28265 , RIdebd3e0_617, \9044_9343 );
and \U$19155 ( \27964_28266 , RIdeba6e0_585, \9046_9345 );
and \U$19156 ( \27965_28267 , RIdeb79e0_553, \9048_9347 );
and \U$19157 ( \27966_28268 , RIfcb9858_7133, \9050_9349 );
and \U$19158 ( \27967_28269 , RIdeb1fe0_489, \9052_9351 );
and \U$19159 ( \27968_28270 , RIfc9efa8_6831, \9054_9353 );
and \U$19160 ( \27969_28271 , RIdeaf2e0_457, \9056_9355 );
and \U$19161 ( \27970_28272 , RIfce0750_7576, \9058_9357 );
and \U$19162 ( \27971_28273 , RIdeab488_425, \9060_9359 );
and \U$19163 ( \27972_28274 , RIdea4b88_393, \9062_9361 );
and \U$19164 ( \27973_28275 , RIde9e288_361, \9064_9363 );
and \U$19165 ( \27974_28276 , RIee1d0b0_4789, \9066_9365 );
and \U$19166 ( \27975_28277 , RIee1c138_4778, \9068_9367 );
and \U$19167 ( \27976_28278 , RIfcd0e68_7399, \9070_9369 );
and \U$19168 ( \27977_28279 , RIfc76d00_6374, \9072_9371 );
and \U$19169 ( \27978_28280 , RIfe89028_7903, \9074_9373 );
and \U$19170 ( \27979_28281 , RIfe88d58_7901, \9076_9375 );
and \U$19171 ( \27980_28282 , RIfe88ec0_7902, \9078_9377 );
and \U$19172 ( \27981_28283 , RIfe88bf0_7900, \9080_9379 );
and \U$19173 ( \27982_28284 , RIfcda7b0_7508, \9082_9381 );
and \U$19174 ( \27983_28285 , RIfc4d810_5904, \9084_9383 );
and \U$19175 ( \27984_28286 , RIfc52dd8_5965, \9086_9385 );
and \U$19176 ( \27985_28287 , RIfcde590_7552, \9088_9387 );
and \U$19177 ( \27986_28288 , RIfc4f868_5927, \9090_9389 );
and \U$19178 ( \27987_28289 , RIe16bd50_2604, \9092_9391 );
and \U$19179 ( \27988_28290 , RIfc68930_6212, \9094_9393 );
and \U$19180 ( \27989_28291 , RIe1683a8_2563, \9096_9395 );
and \U$19181 ( \27990_28292 , RIe165ae0_2534, \9098_9397 );
and \U$19182 ( \27991_28293 , RIe162de0_2502, \9100_9399 );
and \U$19183 ( \27992_28294 , RIfe88a88_7899, \9102_9401 );
and \U$19184 ( \27993_28295 , RIe1600e0_2470, \9104_9403 );
and \U$19185 ( \27994_28296 , RIfcc9140_7310, \9106_9405 );
and \U$19186 ( \27995_28297 , RIe15d3e0_2438, \9108_9407 );
and \U$19187 ( \27996_28298 , RIe1579e0_2374, \9110_9409 );
and \U$19188 ( \27997_28299 , RIe154ce0_2342, \9112_9411 );
and \U$19189 ( \27998_28300 , RIfc698a8_6223, \9114_9413 );
and \U$19190 ( \27999_28301 , RIe151fe0_2310, \9116_9415 );
and \U$19191 ( \28000_28302 , RIee35098_5062, \9118_9417 );
and \U$19192 ( \28001_28303 , RIe14f2e0_2278, \9120_9419 );
and \U$19193 ( \28002_28304 , RIfcc0338_7209, \9122_9421 );
and \U$19194 ( \28003_28305 , RIe14c5e0_2246, \9124_9423 );
and \U$19195 ( \28004_28306 , RIe1498e0_2214, \9126_9425 );
and \U$19196 ( \28005_28307 , RIe146be0_2182, \9128_9427 );
and \U$19197 ( \28006_28308 , RIfc88208_6571, \9130_9429 );
and \U$19198 ( \28007_28309 , RIfc85670_6540, \9132_9431 );
and \U$19199 ( \28008_28310 , RIfc81f98_6501, \9134_9433 );
and \U$19200 ( \28009_28311 , RIfcc4f28_7263, \9136_9435 );
and \U$19201 ( \28010_28312 , RIe1414b0_2120, \9138_9437 );
and \U$19202 ( \28011_28313 , RIe13f188_2095, \9140_9439 );
and \U$19203 ( \28012_28314 , RIdf3d090_2071, \9142_9441 );
and \U$19204 ( \28013_28315 , RIdf3aa98_2044, \9144_9443 );
and \U$19205 ( \28014_28316 , RIfcd2920_7418, \9146_9445 );
and \U$19206 ( \28015_28317 , RIfc7d7e0_6450, \9148_9447 );
and \U$19207 ( \28016_28318 , RIfc49760_5858, \9150_9449 );
and \U$19208 ( \28017_28319 , RIfce5a48_7635, \9152_9451 );
and \U$19209 ( \28018_28320 , RIdf35ea8_1990, \9154_9453 );
and \U$19210 ( \28019_28321 , RIdf338b0_1963, \9156_9455 );
and \U$19211 ( \28020_28322 , RIfe88920_7898, \9158_9457 );
and \U$19212 ( \28021_28323 , RIdf2f800_1917, \9160_9459 );
or \U$19213 ( \28022_28324 , \27958_28260 , \27959_28261 , \27960_28262 , \27961_28263 , \27962_28264 , \27963_28265 , \27964_28266 , \27965_28267 , \27966_28268 , \27967_28269 , \27968_28270 , \27969_28271 , \27970_28272 , \27971_28273 , \27972_28274 , \27973_28275 , \27974_28276 , \27975_28277 , \27976_28278 , \27977_28279 , \27978_28280 , \27979_28281 , \27980_28282 , \27981_28283 , \27982_28284 , \27983_28285 , \27984_28286 , \27985_28287 , \27986_28288 , \27987_28289 , \27988_28290 , \27989_28291 , \27990_28292 , \27991_28293 , \27992_28294 , \27993_28295 , \27994_28296 , \27995_28297 , \27996_28298 , \27997_28299 , \27998_28300 , \27999_28301 , \28000_28302 , \28001_28303 , \28002_28304 , \28003_28305 , \28004_28306 , \28005_28307 , \28006_28308 , \28007_28309 , \28008_28310 , \28009_28311 , \28010_28312 , \28011_28313 , \28012_28314 , \28013_28315 , \28014_28316 , \28015_28317 , \28016_28318 , \28017_28319 , \28018_28320 , \28019_28321 , \28020_28322 , \28021_28323 );
and \U$19214 ( \28023_28325 , RIee2bfc0_4959, \9163_9462 );
and \U$19215 ( \28024_28326 , RIee2a670_4941, \9165_9464 );
and \U$19216 ( \28025_28327 , RIee29158_4926, \9167_9466 );
and \U$19217 ( \28026_28328 , RIee27f10_4913, \9169_9468 );
and \U$19218 ( \28027_28329 , RIdf2a7d8_1860, \9171_9470 );
and \U$19219 ( \28028_28330 , RIdf28618_1836, \9173_9472 );
and \U$19220 ( \28029_28331 , RIdf26890_1815, \9175_9474 );
and \U$19221 ( \28030_28332 , RIdf24dd8_1796, \9177_9476 );
and \U$19222 ( \28031_28333 , RIfcad918_6997, \9179_9478 );
and \U$19223 ( \28032_28334 , RIfc69fb0_6228, \9181_9480 );
and \U$19224 ( \28033_28335 , RIfc63368_6151, \9183_9482 );
and \U$19225 ( \28034_28336 , RIfc623f0_6140, \9185_9484 );
and \U$19226 ( \28035_28337 , RIfc60938_6121, \9187_9486 );
and \U$19227 ( \28036_28338 , RIdf1ff18_1740, \9189_9488 );
and \U$19228 ( \28037_28339 , RIfcba500_7142, \9191_9490 );
and \U$19229 ( \28038_28340 , RIdf19870_1667, \9193_9492 );
and \U$19230 ( \28039_28341 , RIdf176b0_1643, \9195_9494 );
and \U$19231 ( \28040_28342 , RIdf149b0_1611, \9197_9496 );
and \U$19232 ( \28041_28343 , RIdf11cb0_1579, \9199_9498 );
and \U$19233 ( \28042_28344 , RIdf0efb0_1547, \9201_9500 );
and \U$19234 ( \28043_28345 , RIdf0c2b0_1515, \9203_9502 );
and \U$19235 ( \28044_28346 , RIdf095b0_1483, \9205_9504 );
and \U$19236 ( \28045_28347 , RIdf068b0_1451, \9207_9506 );
and \U$19237 ( \28046_28348 , RIdf03bb0_1419, \9209_9508 );
and \U$19238 ( \28047_28349 , RIdefe1b0_1355, \9211_9510 );
and \U$19239 ( \28048_28350 , RIdefb4b0_1323, \9213_9512 );
and \U$19240 ( \28049_28351 , RIdef87b0_1291, \9215_9514 );
and \U$19241 ( \28050_28352 , RIdef5ab0_1259, \9217_9516 );
and \U$19242 ( \28051_28353 , RIdef2db0_1227, \9219_9518 );
and \U$19243 ( \28052_28354 , RIdef00b0_1195, \9221_9520 );
and \U$19244 ( \28053_28355 , RIdeed3b0_1163, \9223_9522 );
and \U$19245 ( \28054_28356 , RIdeea6b0_1131, \9225_9524 );
and \U$19246 ( \28055_28357 , RIfcc9848_7315, \9227_9526 );
and \U$19247 ( \28056_28358 , RIfc69a10_6224, \9229_9528 );
and \U$19248 ( \28057_28359 , RIfcacc70_6988, \9231_9530 );
and \U$19249 ( \28058_28360 , RIfccbfa8_7343, \9233_9532 );
and \U$19250 ( \28059_28361 , RIdee4f80_1069, \9235_9534 );
and \U$19251 ( \28060_28362 , RIdee31f8_1048, \9237_9536 );
and \U$19252 ( \28061_28363 , RIdee1038_1024, \9239_9538 );
and \U$19253 ( \28062_28364 , RIdedee78_1000, \9241_9540 );
and \U$19254 ( \28063_28365 , RIfc84590_6528, \9243_9542 );
and \U$19255 ( \28064_28366 , RIfc9bba0_6794, \9245_9544 );
and \U$19256 ( \28065_28367 , RIee21b38_4842, \9247_9546 );
and \U$19257 ( \28066_28368 , RIfc47168_5831, \9249_9548 );
and \U$19258 ( \28067_28369 , RIded9e50_943, \9251_9550 );
and \U$19259 ( \28068_28370 , RIded7858_916, \9253_9552 );
and \U$19260 ( \28069_28371 , RIfe887b8_7897, \9255_9554 );
and \U$19261 ( \28070_28372 , RIded34d8_868, \9257_9556 );
and \U$19262 ( \28071_28373 , RIded0ee0_841, \9259_9558 );
and \U$19263 ( \28072_28374 , RIdece1e0_809, \9261_9560 );
and \U$19264 ( \28073_28375 , RIdecb4e0_777, \9263_9562 );
and \U$19265 ( \28074_28376 , RIdec87e0_745, \9265_9564 );
and \U$19266 ( \28075_28377 , RIdeb4ce0_521, \9267_9566 );
and \U$19267 ( \28076_28378 , RIde97988_329, \9269_9568 );
and \U$19268 ( \28077_28379 , RIe16e8e8_2635, \9271_9570 );
and \U$19269 ( \28078_28380 , RIe15a6e0_2406, \9273_9572 );
and \U$19270 ( \28079_28381 , RIe143ee0_2150, \9275_9574 );
and \U$19271 ( \28080_28382 , RIdf388d8_2020, \9277_9576 );
and \U$19272 ( \28081_28383 , RIdf2cf38_1888, \9279_9578 );
and \U$19273 ( \28082_28384 , RIdf1d7b8_1712, \9281_9580 );
and \U$19274 ( \28083_28385 , RIdf00eb0_1387, \9283_9582 );
and \U$19275 ( \28084_28386 , RIdee79b0_1099, \9285_9584 );
and \U$19276 ( \28085_28387 , RIdedc718_972, \9287_9586 );
and \U$19277 ( \28086_28388 , RIde7d8d0_202, \9289_9588 );
or \U$19278 ( \28087_28389 , \28023_28325 , \28024_28326 , \28025_28327 , \28026_28328 , \28027_28329 , \28028_28330 , \28029_28331 , \28030_28332 , \28031_28333 , \28032_28334 , \28033_28335 , \28034_28336 , \28035_28337 , \28036_28338 , \28037_28339 , \28038_28340 , \28039_28341 , \28040_28342 , \28041_28343 , \28042_28344 , \28043_28345 , \28044_28346 , \28045_28347 , \28046_28348 , \28047_28349 , \28048_28350 , \28049_28351 , \28050_28352 , \28051_28353 , \28052_28354 , \28053_28355 , \28054_28356 , \28055_28357 , \28056_28358 , \28057_28359 , \28058_28360 , \28059_28361 , \28060_28362 , \28061_28363 , \28062_28364 , \28063_28365 , \28064_28366 , \28065_28367 , \28066_28368 , \28067_28369 , \28068_28370 , \28069_28371 , \28070_28372 , \28071_28373 , \28072_28374 , \28073_28375 , \28074_28376 , \28075_28377 , \28076_28378 , \28077_28379 , \28078_28380 , \28079_28381 , \28080_28382 , \28081_28383 , \28082_28384 , \28083_28385 , \28084_28386 , \28085_28387 , \28086_28388 );
or \U$19279 ( \28088_28390 , \28022_28324 , \28087_28389 );
_DC \g5fc4/U$1 ( \28089 , \28088_28390 , \9298_9597 );
and \U$19280 ( \28090_28392 , RIe19dd78_3173, \8760_9059 );
and \U$19281 ( \28091_28393 , RIe19b078_3141, \8762_9061 );
and \U$19282 ( \28092_28394 , RIfca1438_6857, \8764_9063 );
and \U$19283 ( \28093_28395 , RIe198378_3109, \8766_9065 );
and \U$19284 ( \28094_28396 , RIfca35f8_6881, \8768_9067 );
and \U$19285 ( \28095_28397 , RIe195678_3077, \8770_9069 );
and \U$19286 ( \28096_28398 , RIe192978_3045, \8772_9071 );
and \U$19287 ( \28097_28399 , RIe18fc78_3013, \8774_9073 );
and \U$19288 ( \28098_28400 , RIe18a278_2949, \8776_9075 );
and \U$19289 ( \28099_28401 , RIe187578_2917, \8778_9077 );
and \U$19290 ( \28100_28402 , RIfcba230_7140, \8780_9079 );
and \U$19291 ( \28101_28403 , RIe184878_2885, \8782_9081 );
and \U$19292 ( \28102_28404 , RIf142d90_5220, \8784_9083 );
and \U$19293 ( \28103_28405 , RIe181b78_2853, \8786_9085 );
and \U$19294 ( \28104_28406 , RIe17ee78_2821, \8788_9087 );
and \U$19295 ( \28105_28407 , RIe17c178_2789, \8790_9089 );
and \U$19296 ( \28106_28408 , RIfc9be70_6796, \8792_9091 );
and \U$19297 ( \28107_28409 , RIfc9bd08_6795, \8794_9093 );
and \U$19298 ( \28108_28410 , RIfc4ccd0_5896, \8796_9095 );
and \U$19299 ( \28109_28411 , RIe176070_2720, \8798_9097 );
and \U$19300 ( \28110_28412 , RIfc87c68_6567, \8800_9099 );
and \U$19301 ( \28111_28413 , RIfc87b00_6566, \8802_9101 );
and \U$19302 ( \28112_28414 , RIfcc4c58_7261, \8804_9103 );
and \U$19303 ( \28113_28415 , RIfc4fca0_5930, \8806_9105 );
and \U$19304 ( \28114_28416 , RIfc4f598_5925, \8808_9107 );
and \U$19305 ( \28115_28417 , RIfc876c8_6563, \8810_9109 );
and \U$19306 ( \28116_28418 , RIfc4dae0_5906, \8812_9111 );
and \U$19307 ( \28117_28419 , RIe173eb0_2696, \8814_9113 );
and \U$19308 ( \28118_28420 , RIfcb9420_7130, \8816_9115 );
and \U$19309 ( \28119_28421 , RIfc4e080_5910, \8818_9117 );
and \U$19310 ( \28120_28422 , RIfc4e350_5912, \8820_9119 );
and \U$19311 ( \28121_28423 , RIfc9d388_6811, \8822_9121 );
and \U$19312 ( \28122_28424 , RIfc40a48_5761, \8824_9123 );
and \U$19313 ( \28123_28425 , RIe2240d0_4700, \8826_9125 );
and \U$19314 ( \28124_28426 , RIfc85508_6539, \8828_9127 );
and \U$19315 ( \28125_28427 , RIe2213d0_4668, \8830_9129 );
and \U$19316 ( \28126_28428 , RIfc9ba38_6793, \8832_9131 );
and \U$19317 ( \28127_28429 , RIe21e6d0_4636, \8834_9133 );
and \U$19318 ( \28128_28430 , RIe218cd0_4572, \8836_9135 );
and \U$19319 ( \28129_28431 , RIe215fd0_4540, \8838_9137 );
and \U$19320 ( \28130_28432 , RIfc52c70_5964, \8840_9139 );
and \U$19321 ( \28131_28433 , RIe2132d0_4508, \8842_9141 );
and \U$19322 ( \28132_28434 , RIfca3760_6882, \8844_9143 );
and \U$19323 ( \28133_28435 , RIe2105d0_4476, \8846_9145 );
and \U$19324 ( \28134_28436 , RIfc97988_6747, \8848_9147 );
and \U$19325 ( \28135_28437 , RIe20d8d0_4444, \8850_9149 );
and \U$19326 ( \28136_28438 , RIe20abd0_4412, \8852_9151 );
and \U$19327 ( \28137_28439 , RIe207ed0_4380, \8854_9153 );
and \U$19328 ( \28138_28440 , RIfceb5b0_7700, \8856_9155 );
and \U$19329 ( \28139_28441 , RIfcddbb8_7545, \8858_9157 );
and \U$19330 ( \28140_28442 , RIe202a70_4320, \8860_9159 );
and \U$19331 ( \28141_28443 , RIe200e50_4300, \8862_9161 );
and \U$19332 ( \28142_28444 , RIfc73d30_6340, \8864_9163 );
and \U$19333 ( \28143_28445 , RIfcaf100_7014, \8866_9165 );
and \U$19334 ( \28144_28446 , RIfc71468_6311, \8868_9167 );
and \U$19335 ( \28145_28447 , RIfcdcad8_7533, \8870_9169 );
and \U$19336 ( \28146_28448 , RIfcdda50_7544, \8872_9171 );
and \U$19337 ( \28147_28449 , RIfca8620_6938, \8874_9173 );
and \U$19338 ( \28148_28450 , RIe1fcf08_4255, \8876_9175 );
and \U$19339 ( \28149_28451 , RIe1fbcc0_4242, \8878_9177 );
and \U$19340 ( \28150_28452 , RIfc6c008_6251, \8880_9179 );
and \U$19341 ( \28151_28453 , RIfcdd1e0_7538, \8882_9181 );
and \U$19342 ( \28152_28454 , RIfca9700_6950, \8884_9183 );
and \U$19343 ( \28153_28455 , RIfca92c8_6947, \8886_9185 );
or \U$19344 ( \28154_28456 , \28090_28392 , \28091_28393 , \28092_28394 , \28093_28395 , \28094_28396 , \28095_28397 , \28096_28398 , \28097_28399 , \28098_28400 , \28099_28401 , \28100_28402 , \28101_28403 , \28102_28404 , \28103_28405 , \28104_28406 , \28105_28407 , \28106_28408 , \28107_28409 , \28108_28410 , \28109_28411 , \28110_28412 , \28111_28413 , \28112_28414 , \28113_28415 , \28114_28416 , \28115_28417 , \28116_28418 , \28117_28419 , \28118_28420 , \28119_28421 , \28120_28422 , \28121_28423 , \28122_28424 , \28123_28425 , \28124_28426 , \28125_28427 , \28126_28428 , \28127_28429 , \28128_28430 , \28129_28431 , \28130_28432 , \28131_28433 , \28132_28434 , \28133_28435 , \28134_28436 , \28135_28437 , \28136_28438 , \28137_28439 , \28138_28440 , \28139_28441 , \28140_28442 , \28141_28443 , \28142_28444 , \28143_28445 , \28144_28446 , \28145_28447 , \28146_28448 , \28147_28449 , \28148_28450 , \28149_28451 , \28150_28452 , \28151_28453 , \28152_28454 , \28153_28455 );
and \U$19345 ( \28155_28457 , RIfcce5a0_7370, \8889_9188 );
and \U$19346 ( \28156_28458 , RIfc6ba68_6247, \8891_9190 );
and \U$19347 ( \28157_28459 , RIfc6f410_6288, \8893_9192 );
and \U$19348 ( \28158_28460 , RIe1fa640_4226, \8895_9194 );
and \U$19349 ( \28159_28461 , RIfcce000_7366, \8897_9196 );
and \U$19350 ( \28160_28462 , RIfc53918_5973, \8899_9198 );
and \U$19351 ( \28161_28463 , RIfcce708_7371, \8901_9200 );
and \U$19352 ( \28162_28464 , RIe1f5bb8_4173, \8903_9202 );
and \U$19353 ( \28163_28465 , RIf1535f0_5408, \8905_9204 );
and \U$19354 ( \28164_28466 , RIf151e08_5391, \8907_9206 );
and \U$19355 ( \28165_28467 , RIfc72db8_6329, \8909_9208 );
and \U$19356 ( \28166_28468 , RIe1f3890_4148, \8911_9210 );
and \U$19357 ( \28167_28469 , RIf14fc48_5367, \8913_9212 );
and \U$19358 ( \28168_28470 , RIfc72c50_6328, \8915_9214 );
and \U$19359 ( \28169_28471 , RIfc73e98_6341, \8917_9216 );
and \U$19360 ( \28170_28472 , RIe1ee598_4089, \8919_9218 );
and \U$19361 ( \28171_28473 , RIe1ebe38_4061, \8921_9220 );
and \U$19362 ( \28172_28474 , RIe1e9138_4029, \8923_9222 );
and \U$19363 ( \28173_28475 , RIe1e6438_3997, \8925_9224 );
and \U$19364 ( \28174_28476 , RIe1e3738_3965, \8927_9226 );
and \U$19365 ( \28175_28477 , RIe1e0a38_3933, \8929_9228 );
and \U$19366 ( \28176_28478 , RIe1ddd38_3901, \8931_9230 );
and \U$19367 ( \28177_28479 , RIe1db038_3869, \8933_9232 );
and \U$19368 ( \28178_28480 , RIe1d8338_3837, \8935_9234 );
and \U$19369 ( \28179_28481 , RIe1d2938_3773, \8937_9236 );
and \U$19370 ( \28180_28482 , RIe1cfc38_3741, \8939_9238 );
and \U$19371 ( \28181_28483 , RIe1ccf38_3709, \8941_9240 );
and \U$19372 ( \28182_28484 , RIe1ca238_3677, \8943_9242 );
and \U$19373 ( \28183_28485 , RIe1c7538_3645, \8945_9244 );
and \U$19374 ( \28184_28486 , RIe1c4838_3613, \8947_9246 );
and \U$19375 ( \28185_28487 , RIe1c1b38_3581, \8949_9248 );
and \U$19376 ( \28186_28488 , RIe1bee38_3549, \8951_9250 );
and \U$19377 ( \28187_28489 , RIfcb8a48_7123, \8953_9252 );
and \U$19378 ( \28188_28490 , RIfcb84a8_7119, \8955_9254 );
and \U$19379 ( \28189_28491 , RIe1b9870_3488, \8957_9256 );
and \U$19380 ( \28190_28492 , RIe1b7818_3465, \8959_9258 );
and \U$19381 ( \28191_28493 , RIfc85940_6542, \8961_9260 );
and \U$19382 ( \28192_28494 , RIfc9e198_6821, \8963_9262 );
and \U$19383 ( \28193_28495 , RIfeac140_8274, \8965_9264 );
and \U$19384 ( \28194_28496 , RIe1b42a8_3427, \8967_9266 );
and \U$19385 ( \28195_28497 , RIfc518c0_5950, \8969_9268 );
and \U$19386 ( \28196_28498 , RIfc838e8_6519, \8971_9270 );
and \U$19387 ( \28197_28499 , RIfe884e8_7895, \8973_9272 );
and \U$19388 ( \28198_28500 , RIe1b1008_3391, \8975_9274 );
and \U$19389 ( \28199_28501 , RIfcc5900_7270, \8977_9276 );
and \U$19390 ( \28200_28502 , RIfc82ad8_6509, \8979_9278 );
and \U$19391 ( \28201_28503 , RIe1ac9b8_3341, \8981_9280 );
and \U$19392 ( \28202_28504 , RIfe88650_7896, \8983_9282 );
and \U$19393 ( \28203_28505 , RIe1a9178_3301, \8985_9284 );
and \U$19394 ( \28204_28506 , RIe1a6478_3269, \8987_9286 );
and \U$19395 ( \28205_28507 , RIe1a3778_3237, \8989_9288 );
and \U$19396 ( \28206_28508 , RIe1a0a78_3205, \8991_9290 );
and \U$19397 ( \28207_28509 , RIe18cf78_2981, \8993_9292 );
and \U$19398 ( \28208_28510 , RIe179478_2757, \8995_9294 );
and \U$19399 ( \28209_28511 , RIe226dd0_4732, \8997_9296 );
and \U$19400 ( \28210_28512 , RIe21b9d0_4604, \8999_9298 );
and \U$19401 ( \28211_28513 , RIe2051d0_4348, \9001_9300 );
and \U$19402 ( \28212_28514 , RIe1ff230_4280, \9003_9302 );
and \U$19403 ( \28213_28515 , RIe1f85e8_4203, \9005_9304 );
and \U$19404 ( \28214_28516 , RIe1f1130_4120, \9007_9306 );
and \U$19405 ( \28215_28517 , RIe1d5638_3805, \9009_9308 );
and \U$19406 ( \28216_28518 , RIe1bc138_3517, \9011_9310 );
and \U$19407 ( \28217_28519 , RIe1aefb0_3368, \9013_9312 );
and \U$19408 ( \28218_28520 , RIe1715e8_2667, \9015_9314 );
or \U$19409 ( \28219_28521 , \28155_28457 , \28156_28458 , \28157_28459 , \28158_28460 , \28159_28461 , \28160_28462 , \28161_28463 , \28162_28464 , \28163_28465 , \28164_28466 , \28165_28467 , \28166_28468 , \28167_28469 , \28168_28470 , \28169_28471 , \28170_28472 , \28171_28473 , \28172_28474 , \28173_28475 , \28174_28476 , \28175_28477 , \28176_28478 , \28177_28479 , \28178_28480 , \28179_28481 , \28180_28482 , \28181_28483 , \28182_28484 , \28183_28485 , \28184_28486 , \28185_28487 , \28186_28488 , \28187_28489 , \28188_28490 , \28189_28491 , \28190_28492 , \28191_28493 , \28192_28494 , \28193_28495 , \28194_28496 , \28195_28497 , \28196_28498 , \28197_28499 , \28198_28500 , \28199_28501 , \28200_28502 , \28201_28503 , \28202_28504 , \28203_28505 , \28204_28506 , \28205_28507 , \28206_28508 , \28207_28509 , \28208_28510 , \28209_28511 , \28210_28512 , \28211_28513 , \28212_28514 , \28213_28515 , \28214_28516 , \28215_28517 , \28216_28518 , \28217_28519 , \28218_28520 );
or \U$19410 ( \28220_28522 , \28154_28456 , \28219_28521 );
_DC \g6048/U$1 ( \28221 , \28220_28522 , \9024_9323 );
xor g6049_GF_PartitionCandidate( \28222_28524_nG6049 , \28089 , \28221 );
buf \U$19411 ( \28223_28525 , \28222_28524_nG6049 );
xor \U$19412 ( \28224_28526 , \28223_28525 , \26990_27292 );
and \U$19413 ( \28225_28527 , \10385_10687 , \28224_28526 );
xor \U$19414 ( \28226_28528 , \27957_28259 , \28225_28527 );
xor \U$19415 ( \28227_28529 , \27948_28250 , \28226_28528 );
and \U$19416 ( \28228_28530 , \27011_27313 , \10681_10983 );
_DC \g65c5/U$1 ( \28229 , \28088_28390 , \9298_9597 );
_DC \g65c6/U$1 ( \28230 , \28220_28522 , \9024_9323 );
and g65c7_GF_PartitionCandidate( \28231_28533_nG65c7 , \28229 , \28230 );
buf \U$19417 ( \28232_28534 , \28231_28533_nG65c7 );
and \U$19418 ( \28233_28535 , \28232_28534 , \10389_10691 );
nor \U$19419 ( \28234_28536 , \28228_28530 , \28233_28535 );
xnor \U$19420 ( \28235_28537 , \28234_28536 , \10678_10980 );
and \U$19421 ( \28236_28538 , \13725_14024 , \22243_22542 );
and \U$19422 ( \28237_28539 , \14648_14950 , \21801_22103 );
nor \U$19423 ( \28238_28540 , \28236_28538 , \28237_28539 );
xnor \U$19424 ( \28239_28541 , \28238_28540 , \22249_22548 );
xor \U$19425 ( \28240_28542 , \28235_28537 , \28239_28541 );
and \U$19426 ( \28241_28543 , \12470_12769 , \23839_24138 );
and \U$19427 ( \28242_28544 , \13377_13679 , \23328_23630 );
nor \U$19428 ( \28243_28545 , \28241_28543 , \28242_28544 );
xnor \U$19429 ( \28244_28546 , \28243_28545 , \23845_24144 );
xor \U$19430 ( \28245_28547 , \28240_28542 , \28244_28546 );
xor \U$19431 ( \28246_28548 , \28227_28529 , \28245_28547 );
xor \U$19432 ( \28247_28549 , \27944_28246 , \28246_28548 );
and \U$19433 ( \28248_28550 , \19259_19558 , \16333_16635 );
and \U$19434 ( \28249_28551 , \20242_20544 , \15999_16301 );
nor \U$19435 ( \28250_28552 , \28248_28550 , \28249_28551 );
xnor \U$19436 ( \28251_28553 , \28250_28552 , \16323_16625 );
and \U$19437 ( \28252_28554 , \11287_11586 , \25527_25826 );
and \U$19438 ( \28253_28555 , \12146_12448 , \24962_25264 );
nor \U$19439 ( \28254_28556 , \28252_28554 , \28253_28555 );
xnor \U$19440 ( \28255_28557 , \28254_28556 , \25474_25773 );
xor \U$19441 ( \28256_28558 , \28251_28553 , \28255_28557 );
and \U$19442 ( \28257_28559 , \10686_10988 , \27095_27397 );
and \U$19443 ( \28258_28560 , \10968_11270 , \26505_26807 );
nor \U$19444 ( \28259_28561 , \28257_28559 , \28258_28560 );
xnor \U$19445 ( \28260_28562 , \28259_28561 , \26993_27295 );
xor \U$19446 ( \28261_28563 , \28256_28558 , \28260_28562 );
and \U$19447 ( \28262_28564 , \20734_21033 , \15037_15336 );
and \U$19448 ( \28263_28565 , \21788_22090 , \14661_14963 );
nor \U$19449 ( \28264_28566 , \28262_28564 , \28263_28565 );
xnor \U$19450 ( \28265_28567 , \28264_28566 , \15043_15342 );
and \U$19451 ( \28266_28568 , \16353_16655 , \19235_19534 );
and \U$19452 ( \28267_28569 , \17325_17627 , \18743_19045 );
nor \U$19453 ( \28268_28570 , \28266_28568 , \28267_28569 );
xnor \U$19454 ( \28269_28571 , \28268_28570 , \19241_19540 );
xor \U$19455 ( \28270_28572 , \28265_28567 , \28269_28571 );
and \U$19456 ( \28271_28573 , \15022_15321 , \20706_21005 );
and \U$19457 ( \28272_28574 , \15965_16267 , \20255_20557 );
nor \U$19458 ( \28273_28575 , \28271_28573 , \28272_28574 );
xnor \U$19459 ( \28274_28576 , \28273_28575 , \20712_21011 );
xor \U$19460 ( \28275_28577 , \28270_28572 , \28274_28576 );
xor \U$19461 ( \28276_28578 , \28261_28563 , \28275_28577 );
and \U$19462 ( \28277_28579 , \26723_27025 , \26994_27296 );
and \U$19463 ( \28278_28580 , \23900_24199 , \12491_12790 );
and \U$19464 ( \28279_28581 , \24970_25272 , \12159_12461 );
nor \U$19465 ( \28280_28582 , \28278_28580 , \28279_28581 );
xnor \U$19466 ( \28281_28583 , \28280_28582 , \12481_12780 );
xor \U$19467 ( \28282_28584 , \28277_28579 , \28281_28583 );
and \U$19468 ( \28283_28585 , \17736_18035 , \17791_18090 );
and \U$19469 ( \28284_28586 , \18730_19032 , \17353_17655 );
nor \U$19470 ( \28285_28587 , \28283_28585 , \28284_28586 );
xnor \U$19471 ( \28286_28588 , \28285_28587 , \17747_18046 );
xor \U$19472 ( \28287_28589 , \28282_28584 , \28286_28588 );
xor \U$19473 ( \28288_28590 , \28276_28578 , \28287_28589 );
xor \U$19474 ( \28289_28591 , \28247_28549 , \28288_28590 );
xor \U$19475 ( \28290_28592 , \27930_28232 , \28289_28591 );
and \U$19476 ( \28291_28593 , \26715_27017 , \27055_27357 );
and \U$19477 ( \28292_28594 , \27055_27357 , \27103_27405 );
and \U$19478 ( \28293_28595 , \26715_27017 , \27103_27405 );
or \U$19479 ( \28294_28596 , \28291_28593 , \28292_28594 , \28293_28595 );
xor \U$19480 ( \28295_28597 , \28290_28592 , \28294_28596 );
and \U$19481 ( \28296_28598 , \27104_27406 , \27108_27410 );
and \U$19482 ( \28297_28599 , \27109_27411 , \27112_27414 );
or \U$19483 ( \28298_28600 , \28296_28598 , \28297_28599 );
xor \U$19484 ( \28299_28601 , \28295_28597 , \28298_28600 );
buf g9bc0_GF_PartitionCandidate( \28300_28602_nG9bc0 , \28299_28601 );
and \U$19485 ( \28301_28603 , \10402_10704 , \28300_28602_nG9bc0 );
or \U$19486 ( \28302_28604 , \27901_28203 , \28301_28603 );
xor \U$19487 ( \28303_28605 , \10399_10703 , \28302_28604 );
buf \U$19488 ( \28304_28606 , \28303_28605 );
buf \U$19490 ( \28305_28607 , \28304_28606 );
xor \U$19491 ( \28306_28608 , \27900_28202 , \28305_28607 );
buf \U$19492 ( \28307_28609 , \28306_28608 );
xor \U$19493 ( \28308_28610 , \27833_28135 , \28307_28609 );
and \U$19494 ( \28309_28611 , \26703_27005 , \26709_27011 );
and \U$19495 ( \28310_28612 , \26703_27005 , \27119_27421 );
and \U$19496 ( \28311_28613 , \26709_27011 , \27119_27421 );
or \U$19497 ( \28312_28614 , \28309_28611 , \28310_28612 , \28311_28613 );
buf \U$19498 ( \28313_28615 , \28312_28614 );
xor \U$19499 ( \28314_28616 , \28308_28610 , \28313_28615 );
buf \U$19500 ( \28315_28617 , \28314_28616 );
and \U$19501 ( \28316_28618 , \27165_27464 , \27171_27470 );
and \U$19502 ( \28317_28619 , \27165_27464 , \27178_27477 );
and \U$19503 ( \28318_28620 , \27171_27470 , \27178_27477 );
or \U$19504 ( \28319_28621 , \28316_28618 , \28317_28619 , \28318_28620 );
buf \U$19505 ( \28320_28622 , \28319_28621 );
and \U$19506 ( \28321_28623 , \27138_27440 , \27147_27446 );
and \U$19507 ( \28322_28624 , \27138_27440 , \27154_27453 );
and \U$19508 ( \28323_28625 , \27147_27446 , \27154_27453 );
or \U$19509 ( \28324_28626 , \28321_28623 , \28322_28624 , \28323_28625 );
buf \U$19510 ( \28325_28627 , \28324_28626 );
and \U$19511 ( \28326_28628 , \27141_26431 , \10693_10995_nG9c0b );
and \U$19512 ( \28327_28629 , \26129_26428 , \10981_11283_nG9c08 );
or \U$19513 ( \28328_28630 , \28326_28628 , \28327_28629 );
xor \U$19514 ( \28329_28631 , \26128_26427 , \28328_28630 );
buf \U$19515 ( \28330_28632 , \28329_28631 );
buf \U$19517 ( \28331_28633 , \28330_28632 );
and \U$19518 ( \28332_28634 , \25044_24792 , \11299_11598_nG9c05 );
and \U$19519 ( \28333_28635 , \24490_24789 , \12168_12470_nG9c02 );
or \U$19520 ( \28334_28636 , \28332_28634 , \28333_28635 );
xor \U$19521 ( \28335_28637 , \24489_24788 , \28334_28636 );
buf \U$19522 ( \28336_28638 , \28335_28637 );
buf \U$19524 ( \28337_28639 , \28336_28638 );
xor \U$19525 ( \28338_28640 , \28331_28633 , \28337_28639 );
buf \U$19526 ( \28339_28641 , \28338_28640 );
xor \U$19527 ( \28340_28642 , \28325_28627 , \28339_28641 );
and \U$19528 ( \28341_28643 , \20353_20155 , \15074_15373_nG9bf3 );
and \U$19529 ( \28342_28644 , \19853_20152 , \16013_16315_nG9bf0 );
or \U$19530 ( \28343_28645 , \28341_28643 , \28342_28644 );
xor \U$19531 ( \28344_28646 , \19852_20151 , \28343_28645 );
buf \U$19532 ( \28345_28647 , \28344_28646 );
buf \U$19534 ( \28346_28648 , \28345_28647 );
xor \U$19535 ( \28347_28649 , \28340_28642 , \28346_28648 );
buf \U$19536 ( \28348_28650 , \28347_28649 );
and \U$19537 ( \28349_28651 , \27182_27481 , \27188_27487 );
and \U$19538 ( \28350_28652 , \27182_27481 , \27195_27494 );
and \U$19539 ( \28351_28653 , \27188_27487 , \27195_27494 );
or \U$19540 ( \28352_28654 , \28349_28651 , \28350_28652 , \28351_28653 );
buf \U$19541 ( \28353_28655 , \28352_28654 );
xor \U$19542 ( \28354_28656 , \28348_28650 , \28353_28655 );
and \U$19543 ( \28355_28657 , \14710_14631 , \20787_21086_nG9bdb );
and \U$19544 ( \28356_28658 , \14329_14628 , \21827_22129_nG9bd8 );
or \U$19545 ( \28357_28659 , \28355_28657 , \28356_28658 );
xor \U$19546 ( \28358_28660 , \14328_14627 , \28357_28659 );
buf \U$19547 ( \28359_28661 , \28358_28660 );
buf \U$19549 ( \28360_28662 , \28359_28661 );
xor \U$19550 ( \28361_28663 , \28354_28656 , \28360_28662 );
buf \U$19551 ( \28362_28664 , \28361_28663 );
xor \U$19552 ( \28363_28665 , \28320_28622 , \28362_28664 );
and \U$19553 ( \28364_28666 , \10996_10421 , \25561_25860_nG9bc9 );
and \U$19554 ( \28365_28667 , \10119_10418 , \26585_26887_nG9bc6 );
or \U$19555 ( \28366_28668 , \28364_28666 , \28365_28667 );
xor \U$19556 ( \28367_28669 , \10118_10417 , \28366_28668 );
buf \U$19557 ( \28368_28670 , \28367_28669 );
buf \U$19559 ( \28369_28671 , \28368_28670 );
xor \U$19560 ( \28370_28672 , \28363_28665 , \28369_28671 );
buf \U$19561 ( \28371_28673 , \28370_28672 );
and \U$19562 ( \28372_28674 , \27180_27479 , \27211_27510 );
and \U$19563 ( \28373_28675 , \27180_27479 , \27218_27517 );
and \U$19564 ( \28374_28676 , \27211_27510 , \27218_27517 );
or \U$19565 ( \28375_28677 , \28372_28674 , \28373_28675 , \28374_28676 );
buf \U$19566 ( \28376_28678 , \28375_28677 );
xor \U$19567 ( \28377_28679 , \28371_28673 , \28376_28678 );
and \U$19568 ( \28378_28680 , \27238_27537 , \27243_27542 );
and \U$19569 ( \28379_28681 , \27238_27537 , \27250_27549 );
and \U$19570 ( \28380_28682 , \27243_27542 , \27250_27549 );
or \U$19571 ( \28381_28683 , \28378_28680 , \28379_28681 , \28380_28682 );
buf \U$19572 ( \28382_28684 , \28381_28683 );
xor \U$19573 ( \28383_28685 , \28377_28679 , \28382_28684 );
buf \U$19574 ( \28384_28686 , \28383_28685 );
xor \U$19575 ( \28385_28687 , \28315_28617 , \28384_28686 );
and \U$19576 ( \28386_28688 , \26698_27000 , \27121_27423 );
and \U$19577 ( \28387_28689 , \26698_27000 , \27220_27519 );
and \U$19578 ( \28388_28690 , \27121_27423 , \27220_27519 );
or \U$19579 ( \28389_28691 , \28386_28688 , \28387_28689 , \28388_28690 );
buf \U$19580 ( \28390_28692 , \28389_28691 );
xor \U$19581 ( \28391_28693 , \28385_28687 , \28390_28692 );
and \U$19582 ( \28392_28694 , \27823_28125 , \28391_28693 );
and \U$19583 ( \28393_28695 , \27827_28129 , \28391_28693 );
or \U$19584 ( \28394_28696 , \27828_28130 , \28392_28694 , \28393_28695 );
and \U$19585 ( \28395_28697 , \27262_27561 , \27266_27565 );
and \U$19586 ( \28396_28698 , \27262_27561 , \27822_28124 );
and \U$19587 ( \28397_28699 , \27266_27565 , \27822_28124 );
or \U$19588 ( \28398_28700 , \28395_28697 , \28396_28698 , \28397_28699 );
xor \U$19589 ( \28399_28701 , \28394_28696 , \28398_28700 );
and \U$19590 ( \28400_28702 , \28315_28617 , \28384_28686 );
and \U$19591 ( \28401_28703 , \28315_28617 , \28390_28692 );
and \U$19592 ( \28402_28704 , \28384_28686 , \28390_28692 );
or \U$19593 ( \28403_28705 , \28400_28702 , \28401_28703 , \28402_28704 );
xor \U$19594 ( \28404_28706 , \28399_28701 , \28403_28705 );
and \U$19595 ( \28405_28707 , \28371_28673 , \28376_28678 );
and \U$19596 ( \28406_28708 , \28371_28673 , \28382_28684 );
and \U$19597 ( \28407_28709 , \28376_28678 , \28382_28684 );
or \U$19598 ( \28408_28710 , \28405_28707 , \28406_28708 , \28407_28709 );
buf \U$19599 ( \28409_28711 , \28408_28710 );
and \U$19600 ( \28410_28712 , \27885_28187 , \27890_28192 );
and \U$19601 ( \28411_28713 , \27885_28187 , \27897_28199 );
and \U$19602 ( \28412_28714 , \27890_28192 , \27897_28199 );
or \U$19603 ( \28413_28715 , \28410_28712 , \28411_28713 , \28412_28714 );
buf \U$19604 ( \28414_28716 , \28413_28715 );
and \U$19605 ( \28415_28717 , \27870_28172 , \27876_28178 );
and \U$19606 ( \28416_28718 , \27870_28172 , \27883_28185 );
and \U$19607 ( \28417_28719 , \27876_28178 , \27883_28185 );
or \U$19608 ( \28418_28720 , \28415_28717 , \28416_28718 , \28417_28719 );
buf \U$19609 ( \28419_28721 , \28418_28720 );
and \U$19610 ( \28420_28722 , \14710_14631 , \21827_22129_nG9bd8 );
and \U$19611 ( \28421_28723 , \14329_14628 , \22330_22629_nG9bd5 );
or \U$19612 ( \28422_28724 , \28420_28722 , \28421_28723 );
xor \U$19613 ( \28423_28725 , \14328_14627 , \28422_28724 );
buf \U$19614 ( \28424_28726 , \28423_28725 );
buf \U$19616 ( \28425_28727 , \28424_28726 );
xor \U$19617 ( \28426_28728 , \28419_28721 , \28425_28727 );
and \U$19618 ( \28427_28729 , \13431_13370 , \23394_23696_nG9bd2 );
and \U$19619 ( \28428_28730 , \13068_13367 , \23927_24226_nG9bcf );
or \U$19620 ( \28429_28731 , \28427_28729 , \28428_28730 );
xor \U$19621 ( \28430_28732 , \13067_13366 , \28429_28731 );
buf \U$19622 ( \28431_28733 , \28430_28732 );
buf \U$19624 ( \28432_28734 , \28431_28733 );
xor \U$19625 ( \28433_28735 , \28426_28728 , \28432_28734 );
buf \U$19626 ( \28434_28736 , \28433_28735 );
xor \U$19627 ( \28435_28737 , \28414_28716 , \28434_28736 );
and \U$19628 ( \28436_28738 , \27838_28140 , \27844_28146 );
and \U$19629 ( \28437_28739 , \27838_28140 , \27851_28153 );
and \U$19630 ( \28438_28740 , \27844_28146 , \27851_28153 );
or \U$19631 ( \28439_28741 , \28436_28738 , \28437_28739 , \28438_28740 );
buf \U$19632 ( \28440_28742 , \28439_28741 );
xor \U$19633 ( \28441_28743 , \28435_28737 , \28440_28742 );
buf \U$19634 ( \28442_28744 , \28441_28743 );
xor \U$19635 ( \28443_28745 , \28409_28711 , \28442_28744 );
and \U$19636 ( \28444_28746 , \27853_28155 , \27899_28201 );
and \U$19637 ( \28445_28747 , \27853_28155 , \28305_28607 );
and \U$19638 ( \28446_28748 , \27899_28201 , \28305_28607 );
or \U$19639 ( \28447_28749 , \28444_28746 , \28445_28747 , \28446_28748 );
buf \U$19640 ( \28448_28750 , \28447_28749 );
xor \U$19641 ( \28449_28751 , \28443_28745 , \28448_28750 );
buf \U$19642 ( \28450_28752 , \28449_28751 );
and \U$19643 ( \28451_28753 , \12183_12157 , \24996_25298_nG9bcc );
and \U$19644 ( \28452_28754 , \11855_12154 , \25561_25860_nG9bc9 );
or \U$19645 ( \28453_28755 , \28451_28753 , \28452_28754 );
xor \U$19646 ( \28454_28756 , \11854_12153 , \28453_28755 );
buf \U$19647 ( \28455_28757 , \28454_28756 );
buf \U$19649 ( \28456_28758 , \28455_28757 );
and \U$19650 ( \28457_28759 , \10996_10421 , \26585_26887_nG9bc6 );
and \U$19651 ( \28458_28760 , \10119_10418 , \27114_27416_nG9bc3 );
or \U$19652 ( \28459_28761 , \28457_28759 , \28458_28760 );
xor \U$19653 ( \28460_28762 , \10118_10417 , \28459_28761 );
buf \U$19654 ( \28461_28763 , \28460_28762 );
buf \U$19656 ( \28462_28764 , \28461_28763 );
xor \U$19657 ( \28463_28765 , \28456_28758 , \28462_28764 );
and \U$19658 ( \28464_28766 , \10411_10707 , \28300_28602_nG9bc0 );
and \U$19659 ( \28465_28767 , \27905_28207 , \27929_28231 );
and \U$19660 ( \28466_28768 , \27929_28231 , \28289_28591 );
and \U$19661 ( \28467_28769 , \27905_28207 , \28289_28591 );
or \U$19662 ( \28468_28770 , \28465_28767 , \28466_28768 , \28467_28769 );
and \U$19663 ( \28469_28771 , \27909_28211 , \27913_28215 );
and \U$19664 ( \28470_28772 , \27913_28215 , \27928_28230 );
and \U$19665 ( \28471_28773 , \27909_28211 , \27928_28230 );
or \U$19666 ( \28472_28774 , \28469_28771 , \28470_28772 , \28471_28773 );
and \U$19667 ( \28473_28775 , \28261_28563 , \28275_28577 );
and \U$19668 ( \28474_28776 , \28275_28577 , \28287_28589 );
and \U$19669 ( \28475_28777 , \28261_28563 , \28287_28589 );
or \U$19670 ( \28476_28778 , \28473_28775 , \28474_28776 , \28475_28777 );
and \U$19671 ( \28477_28779 , \23315_23617 , \13755_14054 );
and \U$19672 ( \28478_28780 , \23900_24199 , \13390_13692 );
nor \U$19673 ( \28479_28781 , \28477_28779 , \28478_28780 );
xnor \U$19674 ( \28480_28782 , \28479_28781 , \13736_14035 );
and \U$19675 ( \28481_28783 , \17325_17627 , \19235_19534 );
and \U$19676 ( \28482_28784 , \17736_18035 , \18743_19045 );
nor \U$19677 ( \28483_28785 , \28481_28783 , \28482_28784 );
xnor \U$19678 ( \28484_28786 , \28483_28785 , \19241_19540 );
xor \U$19679 ( \28485_28787 , \28480_28782 , \28484_28786 );
and \U$19680 ( \28486_28788 , \15965_16267 , \20706_21005 );
and \U$19681 ( \28487_28789 , \16353_16655 , \20255_20557 );
nor \U$19682 ( \28488_28790 , \28486_28788 , \28487_28789 );
xnor \U$19683 ( \28489_28791 , \28488_28790 , \20712_21011 );
xor \U$19684 ( \28490_28792 , \28485_28787 , \28489_28791 );
and \U$19685 ( \28491_28793 , \24970_25272 , \12491_12790 );
and \U$19686 ( \28492_28794 , \25516_25815 , \12159_12461 );
nor \U$19687 ( \28493_28795 , \28491_28793 , \28492_28794 );
xnor \U$19688 ( \28494_28796 , \28493_28795 , \12481_12780 );
and \U$19689 ( \28495_28797 , \10968_11270 , \27095_27397 );
and \U$19690 ( \28496_28798 , \11287_11586 , \26505_26807 );
nor \U$19691 ( \28497_28799 , \28495_28797 , \28496_28798 );
xnor \U$19692 ( \28498_28800 , \28497_28799 , \26993_27295 );
xor \U$19693 ( \28499_28801 , \28494_28796 , \28498_28800 );
and \U$19694 ( \28500_28802 , RIdec5c48_714, \9034_9333 );
and \U$19695 ( \28501_28803 , RIdec2f48_682, \9036_9335 );
and \U$19696 ( \28502_28804 , RIfc7c160_6434, \9038_9337 );
and \U$19697 ( \28503_28805 , RIdec0248_650, \9040_9339 );
and \U$19698 ( \28504_28806 , RIfcb38b8_7065, \9042_9341 );
and \U$19699 ( \28505_28807 , RIdebd548_618, \9044_9343 );
and \U$19700 ( \28506_28808 , RIdeba848_586, \9046_9345 );
and \U$19701 ( \28507_28809 , RIdeb7b48_554, \9048_9347 );
and \U$19702 ( \28508_28810 , RIfce7c08_7659, \9050_9349 );
and \U$19703 ( \28509_28811 , RIdeb2148_490, \9052_9351 );
and \U$19704 ( \28510_28812 , RIfce7aa0_7658, \9054_9353 );
and \U$19705 ( \28511_28813 , RIdeaf448_458, \9056_9355 );
and \U$19706 ( \28512_28814 , RIfca38c8_6883, \9058_9357 );
and \U$19707 ( \28513_28815 , RIdeab7d0_426, \9060_9359 );
and \U$19708 ( \28514_28816 , RIdea4ed0_394, \9062_9361 );
and \U$19709 ( \28515_28817 , RIde9e5d0_362, \9064_9363 );
and \U$19710 ( \28516_28818 , RIfc41e70_5772, \9066_9365 );
and \U$19711 ( \28517_28819 , RIfc5b0a0_6058, \9068_9367 );
and \U$19712 ( \28518_28820 , RIfcdbb60_7522, \9070_9369 );
and \U$19713 ( \28519_28821 , RIfc78650_6392, \9072_9371 );
and \U$19714 ( \28520_28822 , RIfea92d8_8241, \9074_9373 );
and \U$19715 ( \28521_28823 , RIde8e5e0_284, \9076_9375 );
and \U$19716 ( \28522_28824 , RIfea0d40_8174, \9078_9377 );
and \U$19717 ( \28523_28825 , RIfea0bd8_8173, \9080_9379 );
and \U$19718 ( \28524_28826 , RIfcdf508_7563, \9082_9381 );
and \U$19719 ( \28525_28827 , RIfcb1b30_7044, \9084_9383 );
and \U$19720 ( \28526_28828 , RIfc5ccc0_6078, \9086_9385 );
and \U$19721 ( \28527_28829 , RIfcb16f8_7041, \9088_9387 );
and \U$19722 ( \28528_28830 , RIfc77b10_6384, \9090_9389 );
and \U$19723 ( \28529_28831 , RIe16beb8_2605, \9092_9391 );
and \U$19724 ( \28530_28832 , RIe169e60_2582, \9094_9393 );
and \U$19725 ( \28531_28833 , RIe168510_2564, \9096_9395 );
and \U$19726 ( \28532_28834 , RIe165c48_2535, \9098_9397 );
and \U$19727 ( \28533_28835 , RIe162f48_2503, \9100_9399 );
and \U$19728 ( \28534_28836 , RIfc4f9d0_5928, \9102_9401 );
and \U$19729 ( \28535_28837 , RIe160248_2471, \9104_9403 );
and \U$19730 ( \28536_28838 , RIfc4e8f0_5916, \9106_9405 );
and \U$19731 ( \28537_28839 , RIe15d548_2439, \9108_9407 );
and \U$19732 ( \28538_28840 , RIe157b48_2375, \9110_9409 );
and \U$19733 ( \28539_28841 , RIe154e48_2343, \9112_9411 );
and \U$19734 ( \28540_28842 , RIfc4e1e8_5911, \9114_9413 );
and \U$19735 ( \28541_28843 , RIe152148_2311, \9116_9415 );
and \U$19736 ( \28542_28844 , RIfc868b8_6553, \9118_9417 );
and \U$19737 ( \28543_28845 , RIe14f448_2279, \9120_9419 );
and \U$19738 ( \28544_28846 , RIfc865e8_6551, \9122_9421 );
and \U$19739 ( \28545_28847 , RIe14c748_2247, \9124_9423 );
and \U$19740 ( \28546_28848 , RIe149a48_2215, \9126_9425 );
and \U$19741 ( \28547_28849 , RIe146d48_2183, \9128_9427 );
and \U$19742 ( \28548_28850 , RIfc9eb70_6828, \9130_9429 );
and \U$19743 ( \28549_28851 , RIfc9ecd8_6829, \9132_9431 );
and \U$19744 ( \28550_28852 , RIfcc5630_7268, \9134_9433 );
and \U$19745 ( \28551_28853 , RIfc83bb8_6521, \9136_9435 );
and \U$19746 ( \28552_28854 , RIe141618_2121, \9138_9437 );
and \U$19747 ( \28553_28855 , RIfea0ea8_8175, \9140_9439 );
and \U$19748 ( \28554_28856 , RIdf3d1f8_2072, \9142_9441 );
and \U$19749 ( \28555_28857 , RIdf3ac00_2045, \9144_9443 );
and \U$19750 ( \28556_28858 , RIee308e0_5011, \9146_9445 );
and \U$19751 ( \28557_28859 , RIfcd3cd0_7432, \9148_9447 );
and \U$19752 ( \28558_28860 , RIfc84e00_6534, \9150_9449 );
and \U$19753 ( \28559_28861 , RIfc834b0_6516, \9152_9451 );
and \U$19754 ( \28560_28862 , RIdf36010_1991, \9154_9453 );
and \U$19755 ( \28561_28863 , RIdf33a18_1964, \9156_9455 );
and \U$19756 ( \28562_28864 , RIdf31858_1940, \9158_9457 );
and \U$19757 ( \28563_28865 , RIdf2f968_1918, \9160_9459 );
or \U$19758 ( \28564_28866 , \28500_28802 , \28501_28803 , \28502_28804 , \28503_28805 , \28504_28806 , \28505_28807 , \28506_28808 , \28507_28809 , \28508_28810 , \28509_28811 , \28510_28812 , \28511_28813 , \28512_28814 , \28513_28815 , \28514_28816 , \28515_28817 , \28516_28818 , \28517_28819 , \28518_28820 , \28519_28821 , \28520_28822 , \28521_28823 , \28522_28824 , \28523_28825 , \28524_28826 , \28525_28827 , \28526_28828 , \28527_28829 , \28528_28830 , \28529_28831 , \28530_28832 , \28531_28833 , \28532_28834 , \28533_28835 , \28534_28836 , \28535_28837 , \28536_28838 , \28537_28839 , \28538_28840 , \28539_28841 , \28540_28842 , \28541_28843 , \28542_28844 , \28543_28845 , \28544_28846 , \28545_28847 , \28546_28848 , \28547_28849 , \28548_28850 , \28549_28851 , \28550_28852 , \28551_28853 , \28552_28854 , \28553_28855 , \28554_28856 , \28555_28857 , \28556_28858 , \28557_28859 , \28558_28860 , \28559_28861 , \28560_28862 , \28561_28863 , \28562_28864 , \28563_28865 );
and \U$19759 ( \28565_28867 , RIee2c128_4960, \9163_9462 );
and \U$19760 ( \28566_28868 , RIee2a7d8_4942, \9165_9464 );
and \U$19761 ( \28567_28869 , RIee292c0_4927, \9167_9466 );
and \U$19762 ( \28568_28870 , RIee28078_4914, \9169_9468 );
and \U$19763 ( \28569_28871 , RIdf2a940_1861, \9171_9470 );
and \U$19764 ( \28570_28872 , RIdf28780_1837, \9173_9472 );
and \U$19765 ( \28571_28873 , RIfea0a70_8172, \9175_9474 );
and \U$19766 ( \28572_28874 , RIfea0908_8171, \9177_9476 );
and \U$19767 ( \28573_28875 , RIfcd4f18_7445, \9179_9478 );
and \U$19768 ( \28574_28876 , RIfca0628_6847, \9181_9480 );
and \U$19769 ( \28575_28877 , RIdf23050_1775, \9183_9482 );
and \U$19770 ( \28576_28878 , RIfcd3190_7424, \9185_9484 );
and \U$19771 ( \28577_28879 , RIdf21b38_1760, \9187_9486 );
and \U$19772 ( \28578_28880 , RIdf20080_1741, \9189_9488 );
and \U$19773 ( \28579_28881 , RIdf1b328_1686, \9191_9490 );
and \U$19774 ( \28580_28882 , RIdf199d8_1668, \9193_9492 );
and \U$19775 ( \28581_28883 , RIdf17818_1644, \9195_9494 );
and \U$19776 ( \28582_28884 , RIdf14b18_1612, \9197_9496 );
and \U$19777 ( \28583_28885 , RIdf11e18_1580, \9199_9498 );
and \U$19778 ( \28584_28886 , RIdf0f118_1548, \9201_9500 );
and \U$19779 ( \28585_28887 , RIdf0c418_1516, \9203_9502 );
and \U$19780 ( \28586_28888 , RIdf09718_1484, \9205_9504 );
and \U$19781 ( \28587_28889 , RIdf06a18_1452, \9207_9506 );
and \U$19782 ( \28588_28890 , RIdf03d18_1420, \9209_9508 );
and \U$19783 ( \28589_28891 , RIdefe318_1356, \9211_9510 );
and \U$19784 ( \28590_28892 , RIdefb618_1324, \9213_9512 );
and \U$19785 ( \28591_28893 , RIdef8918_1292, \9215_9514 );
and \U$19786 ( \28592_28894 , RIdef5c18_1260, \9217_9516 );
and \U$19787 ( \28593_28895 , RIdef2f18_1228, \9219_9518 );
and \U$19788 ( \28594_28896 , RIdef0218_1196, \9221_9520 );
and \U$19789 ( \28595_28897 , RIdeed518_1164, \9223_9522 );
and \U$19790 ( \28596_28898 , RIdeea818_1132, \9225_9524 );
and \U$19791 ( \28597_28899 , RIfcdf3a0_7562, \9227_9526 );
and \U$19792 ( \28598_28900 , RIfca5218_6901, \9229_9528 );
and \U$19793 ( \28599_28901 , RIfcdc538_7529, \9231_9530 );
and \U$19794 ( \28600_28902 , RIfcdc6a0_7530, \9233_9532 );
and \U$19795 ( \28601_28903 , RIdee50e8_1070, \9235_9534 );
and \U$19796 ( \28602_28904 , RIdee3360_1049, \9237_9536 );
and \U$19797 ( \28603_28905 , RIfea07a0_8170, \9239_9538 );
and \U$19798 ( \28604_28906 , RIdedefe0_1001, \9241_9540 );
and \U$19799 ( \28605_28907 , RIfcb0d20_7034, \9243_9542 );
and \U$19800 ( \28606_28908 , RIfcd4978_7441, \9245_9544 );
and \U$19801 ( \28607_28909 , RIfca49a8_6895, \9247_9546 );
and \U$19802 ( \28608_28910 , RIfca1708_6859, \9249_9548 );
and \U$19803 ( \28609_28911 , RIded9fb8_944, \9251_9550 );
and \U$19804 ( \28610_28912 , RIded79c0_917, \9253_9552 );
and \U$19805 ( \28611_28913 , RIded5ad0_895, \9255_9554 );
and \U$19806 ( \28612_28914 , RIfeab498_8265, \9257_9556 );
and \U$19807 ( \28613_28915 , RIded1048_842, \9259_9558 );
and \U$19808 ( \28614_28916 , RIdece348_810, \9261_9560 );
and \U$19809 ( \28615_28917 , RIdecb648_778, \9263_9562 );
and \U$19810 ( \28616_28918 , RIdec8948_746, \9265_9564 );
and \U$19811 ( \28617_28919 , RIdeb4e48_522, \9267_9566 );
and \U$19812 ( \28618_28920 , RIde97cd0_330, \9269_9568 );
and \U$19813 ( \28619_28921 , RIe16ea50_2636, \9271_9570 );
and \U$19814 ( \28620_28922 , RIe15a848_2407, \9273_9572 );
and \U$19815 ( \28621_28923 , RIe144048_2151, \9275_9574 );
and \U$19816 ( \28622_28924 , RIdf38a40_2021, \9277_9576 );
and \U$19817 ( \28623_28925 , RIdf2d0a0_1889, \9279_9578 );
and \U$19818 ( \28624_28926 , RIdf1d920_1713, \9281_9580 );
and \U$19819 ( \28625_28927 , RIdf01018_1388, \9283_9582 );
and \U$19820 ( \28626_28928 , RIdee7b18_1100, \9285_9584 );
and \U$19821 ( \28627_28929 , RIdedc880_973, \9287_9586 );
and \U$19822 ( \28628_28930 , RIde7dc18_203, \9289_9588 );
or \U$19823 ( \28629_28931 , \28565_28867 , \28566_28868 , \28567_28869 , \28568_28870 , \28569_28871 , \28570_28872 , \28571_28873 , \28572_28874 , \28573_28875 , \28574_28876 , \28575_28877 , \28576_28878 , \28577_28879 , \28578_28880 , \28579_28881 , \28580_28882 , \28581_28883 , \28582_28884 , \28583_28885 , \28584_28886 , \28585_28887 , \28586_28888 , \28587_28889 , \28588_28890 , \28589_28891 , \28590_28892 , \28591_28893 , \28592_28894 , \28593_28895 , \28594_28896 , \28595_28897 , \28596_28898 , \28597_28899 , \28598_28900 , \28599_28901 , \28600_28902 , \28601_28903 , \28602_28904 , \28603_28905 , \28604_28906 , \28605_28907 , \28606_28908 , \28607_28909 , \28608_28910 , \28609_28911 , \28610_28912 , \28611_28913 , \28612_28914 , \28613_28915 , \28614_28916 , \28615_28917 , \28616_28918 , \28617_28919 , \28618_28920 , \28619_28921 , \28620_28922 , \28621_28923 , \28622_28924 , \28623_28925 , \28624_28926 , \28625_28927 , \28626_28928 , \28627_28929 , \28628_28930 );
or \U$19824 ( \28630_28932 , \28564_28866 , \28629_28931 );
_DC \g60cd/U$1 ( \28631 , \28630_28932 , \9298_9597 );
and \U$19825 ( \28632_28934 , RIe19dee0_3174, \8760_9059 );
and \U$19826 ( \28633_28935 , RIe19b1e0_3142, \8762_9061 );
and \U$19827 ( \28634_28936 , RIfc67580_6198, \8764_9063 );
and \U$19828 ( \28635_28937 , RIe1984e0_3110, \8766_9065 );
and \U$19829 ( \28636_28938 , RIfccb030_7332, \8768_9067 );
and \U$19830 ( \28637_28939 , RIe1957e0_3078, \8770_9069 );
and \U$19831 ( \28638_28940 , RIe192ae0_3046, \8772_9071 );
and \U$19832 ( \28639_28941 , RIe18fde0_3014, \8774_9073 );
and \U$19833 ( \28640_28942 , RIe18a3e0_2950, \8776_9075 );
and \U$19834 ( \28641_28943 , RIe1876e0_2918, \8778_9077 );
and \U$19835 ( \28642_28944 , RIfc6a550_6232, \8780_9079 );
and \U$19836 ( \28643_28945 , RIe1849e0_2886, \8782_9081 );
and \U$19837 ( \28644_28946 , RIfcaa7e0_6962, \8784_9083 );
and \U$19838 ( \28645_28947 , RIe181ce0_2854, \8786_9085 );
and \U$19839 ( \28646_28948 , RIe17efe0_2822, \8788_9087 );
and \U$19840 ( \28647_28949 , RIe17c2e0_2790, \8790_9089 );
and \U$19841 ( \28648_28950 , RIfc65d98_6181, \8792_9091 );
and \U$19842 ( \28649_28951 , RIfc65690_6176, \8794_9093 );
and \U$19843 ( \28650_28952 , RIe1772b8_2733, \8796_9095 );
and \U$19844 ( \28651_28953 , RIfea0638_8169, \8798_9097 );
and \U$19845 ( \28652_28954 , RIfcca928_7327, \8800_9099 );
and \U$19846 ( \28653_28955 , RIfc607d0_6120, \8802_9101 );
and \U$19847 ( \28654_28956 , RIfc65258_6173, \8804_9103 );
and \U$19848 ( \28655_28957 , RIee3d798_5158, \8806_9105 );
and \U$19849 ( \28656_28958 , RIee3c3e8_5144, \8808_9107 );
and \U$19850 ( \28657_28959 , RIfca9430_6948, \8810_9109 );
and \U$19851 ( \28658_28960 , RIee39f58_5118, \8812_9111 );
and \U$19852 ( \28659_28961 , RIe174018_2697, \8814_9113 );
and \U$19853 ( \28660_28962 , RIfcecf00_7718, \8816_9115 );
and \U$19854 ( \28661_28963 , RIfc650f0_6172, \8818_9117 );
and \U$19855 ( \28662_28964 , RIf16e5a8_5715, \8820_9119 );
and \U$19856 ( \28663_28965 , RIfc43a90_5792, \8822_9121 );
and \U$19857 ( \28664_28966 , RIfc65528_6175, \8824_9123 );
and \U$19858 ( \28665_28967 , RIe224238_4701, \8826_9125 );
and \U$19859 ( \28666_28968 , RIfca9f70_6956, \8828_9127 );
and \U$19860 ( \28667_28969 , RIe221538_4669, \8830_9129 );
and \U$19861 ( \28668_28970 , RIfc6b4c8_6243, \8832_9131 );
and \U$19862 ( \28669_28971 , RIe21e838_4637, \8834_9133 );
and \U$19863 ( \28670_28972 , RIe218e38_4573, \8836_9135 );
and \U$19864 ( \28671_28973 , RIe216138_4541, \8838_9137 );
and \U$19865 ( \28672_28974 , RIfc3fda0_5752, \8840_9139 );
and \U$19866 ( \28673_28975 , RIe213438_4509, \8842_9141 );
and \U$19867 ( \28674_28976 , RIfc61310_6128, \8844_9143 );
and \U$19868 ( \28675_28977 , RIe210738_4477, \8846_9145 );
and \U$19869 ( \28676_28978 , RIfc60c08_6123, \8848_9147 );
and \U$19870 ( \28677_28979 , RIe20da38_4445, \8850_9149 );
and \U$19871 ( \28678_28980 , RIe20ad38_4413, \8852_9151 );
and \U$19872 ( \28679_28981 , RIe208038_4381, \8854_9153 );
and \U$19873 ( \28680_28982 , RIfc66ba8_6191, \8856_9155 );
and \U$19874 ( \28681_28983 , RIfccbcd8_7341, \8858_9157 );
and \U$19875 ( \28682_28984 , RIe202bd8_4321, \8860_9159 );
and \U$19876 ( \28683_28985 , RIe200fb8_4301, \8862_9161 );
and \U$19877 ( \28684_28986 , RIfcadbe8_6999, \8864_9163 );
and \U$19878 ( \28685_28987 , RIfccbe40_7342, \8866_9165 );
and \U$19879 ( \28686_28988 , RIfca7540_6926, \8868_9167 );
and \U$19880 ( \28687_28989 , RIfc6a3e8_6231, \8870_9169 );
and \U$19881 ( \28688_28990 , RIfca6898_6917, \8872_9171 );
and \U$19882 ( \28689_28991 , RIfc73358_6333, \8874_9173 );
and \U$19883 ( \28690_28992 , RIe1fd070_4256, \8876_9175 );
and \U$19884 ( \28691_28993 , RIe1fbe28_4243, \8878_9177 );
and \U$19885 ( \28692_28994 , RIfcc2660_7234, \8880_9179 );
and \U$19886 ( \28693_28995 , RIfc44468_5799, \8882_9181 );
and \U$19887 ( \28694_28996 , RIf15a940_5490, \8884_9183 );
and \U$19888 ( \28695_28997 , RIfca7270_6924, \8886_9185 );
or \U$19889 ( \28696_28998 , \28632_28934 , \28633_28935 , \28634_28936 , \28635_28937 , \28636_28938 , \28637_28939 , \28638_28940 , \28639_28941 , \28640_28942 , \28641_28943 , \28642_28944 , \28643_28945 , \28644_28946 , \28645_28947 , \28646_28948 , \28647_28949 , \28648_28950 , \28649_28951 , \28650_28952 , \28651_28953 , \28652_28954 , \28653_28955 , \28654_28956 , \28655_28957 , \28656_28958 , \28657_28959 , \28658_28960 , \28659_28961 , \28660_28962 , \28661_28963 , \28662_28964 , \28663_28965 , \28664_28966 , \28665_28967 , \28666_28968 , \28667_28969 , \28668_28970 , \28669_28971 , \28670_28972 , \28671_28973 , \28672_28974 , \28673_28975 , \28674_28976 , \28675_28977 , \28676_28978 , \28677_28979 , \28678_28980 , \28679_28981 , \28680_28982 , \28681_28983 , \28682_28984 , \28683_28985 , \28684_28986 , \28685_28987 , \28686_28988 , \28687_28989 , \28688_28990 , \28689_28991 , \28690_28992 , \28691_28993 , \28692_28994 , \28693_28995 , \28694_28996 , \28695_28997 );
and \U$19890 ( \28697_28999 , RIfc5e070_6092, \8889_9188 );
and \U$19891 ( \28698_29000 , RIfc5dda0_6090, \8891_9190 );
and \U$19892 ( \28699_29001 , RIfc7e050_6456, \8893_9192 );
and \U$19893 ( \28700_29002 , RIe1fa7a8_4227, \8895_9194 );
and \U$19894 ( \28701_29003 , RIfc5d968_6087, \8897_9196 );
and \U$19895 ( \28702_29004 , RIfcd9568_7495, \8899_9198 );
and \U$19896 ( \28703_29005 , RIfc8d668_6631, \8901_9200 );
and \U$19897 ( \28704_29006 , RIe1f5d20_4174, \8903_9202 );
and \U$19898 ( \28705_29007 , RIfca4138_6889, \8905_9204 );
and \U$19899 ( \28706_29008 , RIfc8cdf8_6625, \8907_9206 );
and \U$19900 ( \28707_29009 , RIfcc7c28_7295, \8909_9208 );
and \U$19901 ( \28708_29010 , RIe1f39f8_4149, \8911_9210 );
and \U$19902 ( \28709_29011 , RIfc99440_6766, \8913_9212 );
and \U$19903 ( \28710_29012 , RIfcbc3f0_7164, \8915_9214 );
and \U$19904 ( \28711_29013 , RIfc5a128_6047, \8917_9216 );
and \U$19905 ( \28712_29014 , RIe1ee700_4090, \8919_9218 );
and \U$19906 ( \28713_29015 , RIe1ebfa0_4062, \8921_9220 );
and \U$19907 ( \28714_29016 , RIe1e92a0_4030, \8923_9222 );
and \U$19908 ( \28715_29017 , RIe1e65a0_3998, \8925_9224 );
and \U$19909 ( \28716_29018 , RIe1e38a0_3966, \8927_9226 );
and \U$19910 ( \28717_29019 , RIe1e0ba0_3934, \8929_9228 );
and \U$19911 ( \28718_29020 , RIe1ddea0_3902, \8931_9230 );
and \U$19912 ( \28719_29021 , RIe1db1a0_3870, \8933_9232 );
and \U$19913 ( \28720_29022 , RIe1d84a0_3838, \8935_9234 );
and \U$19914 ( \28721_29023 , RIe1d2aa0_3774, \8937_9236 );
and \U$19915 ( \28722_29024 , RIe1cfda0_3742, \8939_9238 );
and \U$19916 ( \28723_29025 , RIe1cd0a0_3710, \8941_9240 );
and \U$19917 ( \28724_29026 , RIe1ca3a0_3678, \8943_9242 );
and \U$19918 ( \28725_29027 , RIe1c76a0_3646, \8945_9244 );
and \U$19919 ( \28726_29028 , RIe1c49a0_3614, \8947_9246 );
and \U$19920 ( \28727_29029 , RIe1c1ca0_3582, \8949_9248 );
and \U$19921 ( \28728_29030 , RIe1befa0_3550, \8951_9250 );
and \U$19922 ( \28729_29031 , RIf14cde0_5334, \8953_9252 );
and \U$19923 ( \28730_29032 , RIf14bb98_5321, \8955_9254 );
and \U$19924 ( \28731_29033 , RIe1b99d8_3489, \8957_9256 );
and \U$19925 ( \28732_29034 , RIe1b7980_3466, \8959_9258 );
and \U$19926 ( \28733_29035 , RIfc4c460_5890, \8961_9260 );
and \U$19927 ( \28734_29036 , RIfc9e738_6825, \8963_9262 );
and \U$19928 ( \28735_29037 , RIe1b5658_3441, \8965_9264 );
and \U$19929 ( \28736_29038 , RIfec54d8_8365, \8967_9266 );
and \U$19930 ( \28737_29039 , RIf149168_5291, \8969_9268 );
and \U$19931 ( \28738_29040 , RIf147f20_5278, \8971_9270 );
and \U$19932 ( \28739_29041 , RIe1b2ac0_3410, \8973_9272 );
and \U$19933 ( \28740_29042 , RIe1b1170_3392, \8975_9274 );
and \U$19934 ( \28741_29043 , RIf1473e0_5270, \8977_9276 );
and \U$19935 ( \28742_29044 , RIf1468a0_5262, \8979_9278 );
and \U$19936 ( \28743_29045 , RIe1acb20_3342, \8981_9280 );
and \U$19937 ( \28744_29046 , RIe1ab338_3325, \8983_9282 );
and \U$19938 ( \28745_29047 , RIe1a92e0_3302, \8985_9284 );
and \U$19939 ( \28746_29048 , RIe1a65e0_3270, \8987_9286 );
and \U$19940 ( \28747_29049 , RIe1a38e0_3238, \8989_9288 );
and \U$19941 ( \28748_29050 , RIe1a0be0_3206, \8991_9290 );
and \U$19942 ( \28749_29051 , RIe18d0e0_2982, \8993_9292 );
and \U$19943 ( \28750_29052 , RIe1795e0_2758, \8995_9294 );
and \U$19944 ( \28751_29053 , RIe226f38_4733, \8997_9296 );
and \U$19945 ( \28752_29054 , RIe21bb38_4605, \8999_9298 );
and \U$19946 ( \28753_29055 , RIe205338_4349, \9001_9300 );
and \U$19947 ( \28754_29056 , RIe1ff398_4281, \9003_9302 );
and \U$19948 ( \28755_29057 , RIe1f8750_4204, \9005_9304 );
and \U$19949 ( \28756_29058 , RIe1f1298_4121, \9007_9306 );
and \U$19950 ( \28757_29059 , RIe1d57a0_3806, \9009_9308 );
and \U$19951 ( \28758_29060 , RIe1bc2a0_3518, \9011_9310 );
and \U$19952 ( \28759_29061 , RIe1af118_3369, \9013_9312 );
and \U$19953 ( \28760_29062 , RIe171750_2668, \9015_9314 );
or \U$19954 ( \28761_29063 , \28697_28999 , \28698_29000 , \28699_29001 , \28700_29002 , \28701_29003 , \28702_29004 , \28703_29005 , \28704_29006 , \28705_29007 , \28706_29008 , \28707_29009 , \28708_29010 , \28709_29011 , \28710_29012 , \28711_29013 , \28712_29014 , \28713_29015 , \28714_29016 , \28715_29017 , \28716_29018 , \28717_29019 , \28718_29020 , \28719_29021 , \28720_29022 , \28721_29023 , \28722_29024 , \28723_29025 , \28724_29026 , \28725_29027 , \28726_29028 , \28727_29029 , \28728_29030 , \28729_29031 , \28730_29032 , \28731_29033 , \28732_29034 , \28733_29035 , \28734_29036 , \28735_29037 , \28736_29038 , \28737_29039 , \28738_29040 , \28739_29041 , \28740_29042 , \28741_29043 , \28742_29044 , \28743_29045 , \28744_29046 , \28745_29047 , \28746_29048 , \28747_29049 , \28748_29050 , \28749_29051 , \28750_29052 , \28751_29053 , \28752_29054 , \28753_29055 , \28754_29056 , \28755_29057 , \28756_29058 , \28757_29059 , \28758_29060 , \28759_29061 , \28760_29062 );
or \U$19955 ( \28762_29064 , \28696_28998 , \28761_29063 );
_DC \g6151/U$1 ( \28763 , \28762_29064 , \9024_9323 );
xor g6152_GF_PartitionCandidate( \28764_29066_nG6152 , \28631 , \28763 );
buf \U$19956 ( \28765_29067 , \28764_29066_nG6152 );
xor \U$19957 ( \28766_29068 , \28765_29067 , \28223_28525 );
not \U$19958 ( \28767_29069 , \28224_28526 );
and \U$19959 ( \28768_29070 , \28766_29068 , \28767_29069 );
and \U$19960 ( \28769_29071 , \10385_10687 , \28768_29070 );
and \U$19961 ( \28770_29072 , \10686_10988 , \28224_28526 );
nor \U$19962 ( \28771_29073 , \28769_29071 , \28770_29072 );
and \U$19963 ( \28772_29074 , \28223_28525 , \26990_27292 );
not \U$19964 ( \28773_29075 , \28772_29074 );
and \U$19965 ( \28774_29076 , \28765_29067 , \28773_29075 );
xnor \U$19966 ( \28775_29077 , \28771_29073 , \28774_29076 );
xor \U$19967 ( \28776_29078 , \28499_28801 , \28775_29077 );
xor \U$19968 ( \28777_29079 , \28490_28792 , \28776_29078 );
and \U$19969 ( \28778_29080 , \28232_28534 , \10681_10983 );
_DC \g65c8/U$1 ( \28779 , \28630_28932 , \9298_9597 );
_DC \g65c9/U$1 ( \28780 , \28762_29064 , \9024_9323 );
and g65ca_GF_PartitionCandidate( \28781_29083_nG65ca , \28779 , \28780 );
buf \U$19970 ( \28782_29084 , \28781_29083_nG65ca );
and \U$19971 ( \28783_29085 , \28782_29084 , \10389_10691 );
nor \U$19972 ( \28784_29086 , \28778_29080 , \28783_29085 );
xnor \U$19973 ( \28785_29087 , \28784_29086 , \10678_10980 );
and \U$19974 ( \28786_29088 , \20242_20544 , \16333_16635 );
and \U$19975 ( \28787_29089 , \20734_21033 , \15999_16301 );
nor \U$19976 ( \28788_29090 , \28786_29088 , \28787_29089 );
xnor \U$19977 ( \28789_29091 , \28788_29090 , \16323_16625 );
xor \U$19978 ( \28790_29092 , \28785_29087 , \28789_29091 );
and \U$19979 ( \28791_29093 , \12146_12448 , \25527_25826 );
and \U$19980 ( \28792_29094 , \12470_12769 , \24962_25264 );
nor \U$19981 ( \28793_29095 , \28791_29093 , \28792_29094 );
xnor \U$19982 ( \28794_29096 , \28793_29095 , \25474_25773 );
xor \U$19983 ( \28795_29097 , \28790_29092 , \28794_29096 );
xor \U$19984 ( \28796_29098 , \28777_29079 , \28795_29097 );
xor \U$19985 ( \28797_29099 , \28476_28778 , \28796_29098 );
and \U$19986 ( \28798_29100 , \28277_28579 , \28281_28583 );
and \U$19987 ( \28799_29101 , \28281_28583 , \28286_28588 );
and \U$19988 ( \28800_29102 , \28277_28579 , \28286_28588 );
or \U$19989 ( \28801_29103 , \28798_29100 , \28799_29101 , \28800_29102 );
and \U$19990 ( \28802_29104 , \21788_22090 , \15037_15336 );
and \U$19991 ( \28803_29105 , \22257_22556 , \14661_14963 );
nor \U$19992 ( \28804_29106 , \28802_29104 , \28803_29105 );
xnor \U$19993 ( \28805_29107 , \28804_29106 , \15043_15342 );
and \U$19994 ( \28806_29108 , \14648_14950 , \22243_22542 );
and \U$19995 ( \28807_29109 , \15022_15321 , \21801_22103 );
nor \U$19996 ( \28808_29110 , \28806_29108 , \28807_29109 );
xnor \U$19997 ( \28809_29111 , \28808_29110 , \22249_22548 );
xor \U$19998 ( \28810_29112 , \28805_29107 , \28809_29111 );
and \U$19999 ( \28811_29113 , \13377_13679 , \23839_24138 );
and \U$20000 ( \28812_29114 , \13725_14024 , \23328_23630 );
nor \U$20001 ( \28813_29115 , \28811_29113 , \28812_29114 );
xnor \U$20002 ( \28814_29116 , \28813_29115 , \23845_24144 );
xor \U$20003 ( \28815_29117 , \28810_29112 , \28814_29116 );
xor \U$20004 ( \28816_29118 , \28801_29103 , \28815_29117 );
and \U$20005 ( \28817_29119 , \26527_26829 , \11275_11574 );
and \U$20006 ( \28818_29120 , \27011_27313 , \10976_11278 );
nor \U$20007 ( \28819_29121 , \28817_29119 , \28818_29120 );
xnor \U$20008 ( \28820_29122 , \28819_29121 , \11281_11580 );
not \U$20009 ( \28821_29123 , \28225_28527 );
and \U$20010 ( \28822_29124 , \28821_29123 , \28774_29076 );
xor \U$20011 ( \28823_29125 , \28820_29122 , \28822_29124 );
and \U$20012 ( \28824_29126 , \27952_28254 , \27956_28258 );
and \U$20013 ( \28825_29127 , \27956_28258 , \28225_28527 );
and \U$20014 ( \28826_29128 , \27952_28254 , \28225_28527 );
or \U$20015 ( \28827_29129 , \28824_29126 , \28825_29127 , \28826_29128 );
xor \U$20016 ( \28828_29130 , \28823_29125 , \28827_29129 );
and \U$20017 ( \28829_29131 , \18730_19032 , \17791_18090 );
and \U$20018 ( \28830_29132 , \19259_19558 , \17353_17655 );
nor \U$20019 ( \28831_29133 , \28829_29131 , \28830_29132 );
xnor \U$20020 ( \28832_29134 , \28831_29133 , \17747_18046 );
xor \U$20021 ( \28833_29135 , \28828_29130 , \28832_29134 );
xor \U$20022 ( \28834_29136 , \28816_29118 , \28833_29135 );
xor \U$20023 ( \28835_29137 , \28797_29099 , \28834_29136 );
xor \U$20024 ( \28836_29138 , \28472_28774 , \28835_29137 );
and \U$20025 ( \28837_29139 , \27918_28220 , \27922_28224 );
and \U$20026 ( \28838_29140 , \27922_28224 , \27927_28229 );
and \U$20027 ( \28839_29141 , \27918_28220 , \27927_28229 );
or \U$20028 ( \28840_29142 , \28837_29139 , \28838_29140 , \28839_29141 );
and \U$20029 ( \28841_29143 , \27944_28246 , \28246_28548 );
and \U$20030 ( \28842_29144 , \28246_28548 , \28288_28590 );
and \U$20031 ( \28843_29145 , \27944_28246 , \28288_28590 );
or \U$20032 ( \28844_29146 , \28841_29143 , \28842_29144 , \28843_29145 );
xor \U$20033 ( \28845_29147 , \28840_29142 , \28844_29146 );
and \U$20034 ( \28846_29148 , \27934_28236 , \27938_28240 );
and \U$20035 ( \28847_29149 , \27938_28240 , \27943_28245 );
and \U$20036 ( \28848_29150 , \27934_28236 , \27943_28245 );
or \U$20037 ( \28849_29151 , \28846_29148 , \28847_29149 , \28848_29150 );
and \U$20038 ( \28850_29152 , \27948_28250 , \28226_28528 );
and \U$20039 ( \28851_29153 , \28226_28528 , \28245_28547 );
and \U$20040 ( \28852_29154 , \27948_28250 , \28245_28547 );
or \U$20041 ( \28853_29155 , \28850_29152 , \28851_29153 , \28852_29154 );
xor \U$20042 ( \28854_29156 , \28849_29151 , \28853_29155 );
and \U$20043 ( \28855_29157 , \28235_28537 , \28239_28541 );
and \U$20044 ( \28856_29158 , \28239_28541 , \28244_28546 );
and \U$20045 ( \28857_29159 , \28235_28537 , \28244_28546 );
or \U$20046 ( \28858_29160 , \28855_29157 , \28856_29158 , \28857_29159 );
and \U$20047 ( \28859_29161 , \28251_28553 , \28255_28557 );
and \U$20048 ( \28860_29162 , \28255_28557 , \28260_28562 );
and \U$20049 ( \28861_29163 , \28251_28553 , \28260_28562 );
or \U$20050 ( \28862_29164 , \28859_29161 , \28860_29162 , \28861_29163 );
xor \U$20051 ( \28863_29165 , \28858_29160 , \28862_29164 );
and \U$20052 ( \28864_29166 , \28265_28567 , \28269_28571 );
and \U$20053 ( \28865_29167 , \28269_28571 , \28274_28576 );
and \U$20054 ( \28866_29168 , \28265_28567 , \28274_28576 );
or \U$20055 ( \28867_29169 , \28864_29166 , \28865_29167 , \28866_29168 );
xor \U$20056 ( \28868_29170 , \28863_29165 , \28867_29169 );
xor \U$20057 ( \28869_29171 , \28854_29156 , \28868_29170 );
xor \U$20058 ( \28870_29172 , \28845_29147 , \28869_29171 );
xor \U$20059 ( \28871_29173 , \28836_29138 , \28870_29172 );
xor \U$20060 ( \28872_29174 , \28468_28770 , \28871_29173 );
and \U$20061 ( \28873_29175 , \28290_28592 , \28294_28596 );
and \U$20062 ( \28874_29176 , \28295_28597 , \28298_28600 );
or \U$20063 ( \28875_29177 , \28873_29175 , \28874_29176 );
xor \U$20064 ( \28876_29178 , \28872_29174 , \28875_29177 );
buf g9bbd_GF_PartitionCandidate( \28877_29179_nG9bbd , \28876_29178 );
and \U$20065 ( \28878_29180 , \10402_10704 , \28877_29179_nG9bbd );
or \U$20066 ( \28879_29181 , \28464_28766 , \28878_29180 );
xor \U$20067 ( \28880_29182 , \10399_10703 , \28879_29181 );
buf \U$20068 ( \28881_29183 , \28880_29182 );
buf \U$20070 ( \28882_29184 , \28881_29183 );
xor \U$20071 ( \28883_29185 , \28463_28765 , \28882_29184 );
buf \U$20072 ( \28884_29186 , \28883_29185 );
and \U$20073 ( \28885_29187 , \28320_28622 , \28362_28664 );
and \U$20074 ( \28886_29188 , \28320_28622 , \28369_28671 );
and \U$20075 ( \28887_29189 , \28362_28664 , \28369_28671 );
or \U$20076 ( \28888_29190 , \28885_29187 , \28886_29188 , \28887_29189 );
buf \U$20077 ( \28889_29191 , \28888_29190 );
xor \U$20078 ( \28890_29192 , \28884_29186 , \28889_29191 );
and \U$20079 ( \28891_29193 , \28348_28650 , \28353_28655 );
and \U$20080 ( \28892_29194 , \28348_28650 , \28360_28662 );
and \U$20081 ( \28893_29195 , \28353_28655 , \28360_28662 );
or \U$20082 ( \28894_29196 , \28891_29193 , \28892_29194 , \28893_29195 );
buf \U$20083 ( \28895_29197 , \28894_29196 );
and \U$20084 ( \28896_29198 , \28325_28627 , \28339_28641 );
and \U$20085 ( \28897_29199 , \28325_28627 , \28346_28648 );
and \U$20086 ( \28898_29200 , \28339_28641 , \28346_28648 );
or \U$20087 ( \28899_29201 , \28896_29198 , \28897_29199 , \28898_29200 );
buf \U$20088 ( \28900_29202 , \28899_29201 );
and \U$20089 ( \28901_29203 , \28331_28633 , \28337_28639 );
buf \U$20090 ( \28902_29204 , \28901_29203 );
and \U$20091 ( \28903_29205 , \23495_23201 , \13403_13705_nG9bfc );
and \U$20092 ( \28904_29206 , \22899_23198 , \13771_14070_nG9bf9 );
or \U$20093 ( \28905_29207 , \28903_29205 , \28904_29206 );
xor \U$20094 ( \28906_29208 , \22898_23197 , \28905_29207 );
buf \U$20095 ( \28907_29209 , \28906_29208 );
buf \U$20097 ( \28908_29210 , \28907_29209 );
xor \U$20098 ( \28909_29211 , \28902_29204 , \28908_29210 );
and \U$20099 ( \28910_29212 , \21908_21658 , \14682_14984_nG9bf6 );
and \U$20100 ( \28911_29213 , \21356_21655 , \15074_15373_nG9bf3 );
or \U$20101 ( \28912_29214 , \28910_29212 , \28911_29213 );
xor \U$20102 ( \28913_29215 , \21355_21654 , \28912_29214 );
buf \U$20103 ( \28914_29216 , \28913_29215 );
buf \U$20105 ( \28915_29217 , \28914_29216 );
xor \U$20106 ( \28916_29218 , \28909_29211 , \28915_29217 );
buf \U$20107 ( \28917_29219 , \28916_29218 );
xor \U$20108 ( \28918_29220 , \28900_29202 , \28917_29219 );
and \U$20109 ( \28919_29221 , \18908_18702 , \17363_17665_nG9bea );
and \U$20110 ( \28920_29222 , \18400_18699 , \17808_18107_nG9be7 );
or \U$20111 ( \28921_29223 , \28919_29221 , \28920_29222 );
xor \U$20112 ( \28922_29224 , \18399_18698 , \28921_29223 );
buf \U$20113 ( \28923_29225 , \28922_29224 );
buf \U$20115 ( \28924_29226 , \28923_29225 );
xor \U$20116 ( \28925_29227 , \28918_29220 , \28924_29226 );
buf \U$20117 ( \28926_29228 , \28925_29227 );
xor \U$20118 ( \28927_29229 , \28895_29197 , \28926_29228 );
and \U$20119 ( \28928_29230 , \27855_28157 , \27861_28163 );
and \U$20120 ( \28929_29231 , \27855_28157 , \27868_28170 );
and \U$20121 ( \28930_29232 , \27861_28163 , \27868_28170 );
or \U$20122 ( \28931_29233 , \28928_29230 , \28929_29231 , \28930_29232 );
buf \U$20123 ( \28932_29234 , \28931_29233 );
and \U$20124 ( \28933_29235 , \27815_28114 , \27819_28121 );
buf \U$20125 ( \28934_29236 , \28933_29235 );
buf \U$20127 ( \28935_29237 , \28934_29236 );
and \U$20128 ( \28936_29238 , \27141_26431 , \10981_11283_nG9c08 );
and \U$20129 ( \28937_29239 , \26129_26428 , \11299_11598_nG9c05 );
or \U$20130 ( \28938_29240 , \28936_29238 , \28937_29239 );
xor \U$20131 ( \28939_29241 , \26128_26427 , \28938_29240 );
buf \U$20132 ( \28940_29242 , \28939_29241 );
buf \U$20134 ( \28941_29243 , \28940_29242 );
xor \U$20135 ( \28942_29244 , \28935_29237 , \28941_29243 );
buf \U$20136 ( \28943_29245 , \28942_29244 );
not \U$18997 ( \28944_28116 , \27816_28115 );
xor \U$18998 ( \28945_28117 , \27810_28109_nG4406 , \27813_28112_nG4409 );
and \U$18999 ( \28946_28118 , \28944_28116 , \28945_28117 );
and \U$20137 ( \28947_29246 , \28946_28118 , \10392_10694_nG9c0e );
and \U$20138 ( \28948_29247 , \27816_28115 , \10693_10995_nG9c0b );
or \U$20139 ( \28949_29248 , \28947_29246 , \28948_29247 );
xor \U$20140 ( \28950_29249 , \27815_28114 , \28949_29248 );
buf \U$20141 ( \28951_29250 , \28950_29249 );
buf \U$20143 ( \28952_29251 , \28951_29250 );
xor \U$20144 ( \28953_29252 , \28943_29245 , \28952_29251 );
and \U$20145 ( \28954_29253 , \25044_24792 , \12168_12470_nG9c02 );
and \U$20146 ( \28955_29254 , \24490_24789 , \12502_12801_nG9bff );
or \U$20147 ( \28956_29255 , \28954_29253 , \28955_29254 );
xor \U$20148 ( \28957_29256 , \24489_24788 , \28956_29255 );
buf \U$20149 ( \28958_29257 , \28957_29256 );
buf \U$20151 ( \28959_29258 , \28958_29257 );
xor \U$20152 ( \28960_29259 , \28953_29252 , \28959_29258 );
buf \U$20153 ( \28961_29260 , \28960_29259 );
xor \U$20154 ( \28962_29261 , \28932_29234 , \28961_29260 );
and \U$20155 ( \28963_29262 , \20353_20155 , \16013_16315_nG9bf0 );
and \U$20156 ( \28964_29263 , \19853_20152 , \16378_16680_nG9bed );
or \U$20157 ( \28965_29264 , \28963_29262 , \28964_29263 );
xor \U$20158 ( \28966_29265 , \19852_20151 , \28965_29264 );
buf \U$20159 ( \28967_29266 , \28966_29265 );
buf \U$20161 ( \28968_29267 , \28967_29266 );
xor \U$20162 ( \28969_29268 , \28962_29261 , \28968_29267 );
buf \U$20163 ( \28970_29269 , \28969_29268 );
and \U$20164 ( \28971_29270 , \17437_17297 , \18789_19091_nG9be4 );
and \U$20165 ( \28972_29271 , \16995_17294 , \19287_19586_nG9be1 );
or \U$20166 ( \28973_29272 , \28971_29270 , \28972_29271 );
xor \U$20167 ( \28974_29273 , \16994_17293 , \28973_29272 );
buf \U$20168 ( \28975_29274 , \28974_29273 );
buf \U$20170 ( \28976_29275 , \28975_29274 );
xor \U$20171 ( \28977_29276 , \28970_29269 , \28976_29275 );
and \U$20172 ( \28978_29277 , \16405_15940 , \20306_20608_nG9bde );
and \U$20173 ( \28979_29278 , \15638_15937 , \20787_21086_nG9bdb );
or \U$20174 ( \28980_29279 , \28978_29277 , \28979_29278 );
xor \U$20175 ( \28981_29280 , \15637_15936 , \28980_29279 );
buf \U$20176 ( \28982_29281 , \28981_29280 );
buf \U$20178 ( \28983_29282 , \28982_29281 );
xor \U$20179 ( \28984_29283 , \28977_29276 , \28983_29282 );
buf \U$20180 ( \28985_29284 , \28984_29283 );
xor \U$20181 ( \28986_29285 , \28927_29229 , \28985_29284 );
buf \U$20182 ( \28987_29286 , \28986_29285 );
xor \U$20183 ( \28988_29287 , \28890_29192 , \28987_29286 );
buf \U$20184 ( \28989_29288 , \28988_29287 );
xor \U$20185 ( \28990_29289 , \28450_28752 , \28989_29288 );
and \U$20186 ( \28991_29290 , \27833_28135 , \28307_28609 );
and \U$20187 ( \28992_29291 , \27833_28135 , \28313_28615 );
and \U$20188 ( \28993_29292 , \28307_28609 , \28313_28615 );
or \U$20189 ( \28994_29293 , \28991_29290 , \28992_29291 , \28993_29292 );
buf \U$20190 ( \28995_29294 , \28994_29293 );
xor \U$20191 ( \28996_29295 , \28990_29289 , \28995_29294 );
and \U$20192 ( \28997_29296 , \28404_28706 , \28996_29295 );
and \U$20193 ( \28998_29297 , \28394_28696 , \28398_28700 );
and \U$20194 ( \28999_29298 , \28394_28696 , \28403_28705 );
and \U$20195 ( \29000_29299 , \28398_28700 , \28403_28705 );
or \U$20196 ( \29001_29300 , \28998_29297 , \28999_29298 , \29000_29299 );
xor \U$20197 ( \29002_29301 , \28997_29296 , \29001_29300 );
and \U$20198 ( \29003_29302 , RIdec5f18_716, \8760_9059 );
and \U$20199 ( \29004_29303 , RIdec3218_684, \8762_9061 );
and \U$20200 ( \29005_29304 , RIee20350_4825, \8764_9063 );
and \U$20201 ( \29006_29305 , RIdec0518_652, \8766_9065 );
and \U$20202 ( \29007_29306 , RIee1f6a8_4816, \8768_9067 );
and \U$20203 ( \29008_29307 , RIdebd818_620, \8770_9069 );
and \U$20204 ( \29009_29308 , RIdebab18_588, \8772_9071 );
and \U$20205 ( \29010_29309 , RIdeb7e18_556, \8774_9073 );
and \U$20206 ( \29011_29310 , RIfce4da0_7626, \8776_9075 );
and \U$20207 ( \29012_29311 , RIdeb2418_492, \8778_9077 );
and \U$20208 ( \29013_29312 , RIfcea908_7691, \8780_9079 );
and \U$20209 ( \29014_29313 , RIdeaf718_460, \8782_9081 );
and \U$20210 ( \29015_29314 , RIfce20a0_7594, \8784_9083 );
and \U$20211 ( \29016_29315 , RIdeabe60_428, \8786_9085 );
and \U$20212 ( \29017_29316 , RIdea5560_396, \8788_9087 );
and \U$20213 ( \29018_29317 , RIde9ec60_364, \8790_9089 );
and \U$20214 ( \29019_29318 , RIfce6420_7642, \8792_9091 );
and \U$20215 ( \29020_29319 , RIee1c2a0_4779, \8794_9093 );
and \U$20216 ( \29021_29320 , RIfc75950_6360, \8796_9095 );
and \U$20217 ( \29022_29321 , RIee1ad88_4764, \8798_9097 );
and \U$20218 ( \29023_29322 , RIde920f0_302, \8800_9099 );
and \U$20219 ( \29024_29323 , RIfea4148_8211, \8802_9101 );
and \U$20220 ( \29025_29324 , RIfeaa688_8255, \8804_9103 );
and \U$20221 ( \29026_29325 , RIfea3fe0_8210, \8806_9105 );
and \U$20222 ( \29027_29326 , RIde82790_226, \8808_9107 );
and \U$20223 ( \29028_29327 , RIfc6f848_6291, \8810_9109 );
and \U$20224 ( \29029_29328 , RIfc5dc38_6089, \8812_9111 );
and \U$20225 ( \29030_29329 , RIfc76b98_6373, \8814_9113 );
and \U$20226 ( \29031_29330 , RIfcae2f0_7004, \8816_9115 );
and \U$20227 ( \29032_29331 , RIe16c020_2606, \8818_9117 );
and \U$20228 ( \29033_29332 , RIe16a130_2584, \8820_9119 );
and \U$20229 ( \29034_29333 , RIe1687e0_2566, \8822_9121 );
and \U$20230 ( \29035_29334 , RIe165f18_2537, \8824_9123 );
and \U$20231 ( \29036_29335 , RIe163218_2505, \8826_9125 );
and \U$20232 ( \29037_29336 , RIfcadd50_7000, \8828_9127 );
and \U$20233 ( \29038_29337 , RIe160518_2473, \8830_9129 );
and \U$20234 ( \29039_29338 , RIfc55268_5991, \8832_9131 );
and \U$20235 ( \29040_29339 , RIe15d818_2441, \8834_9133 );
and \U$20236 ( \29041_29340 , RIe157e18_2377, \8836_9135 );
and \U$20237 ( \29042_29341 , RIe155118_2345, \8838_9137 );
and \U$20238 ( \29043_29342 , RIfc45548_5811, \8840_9139 );
and \U$20239 ( \29044_29343 , RIe152418_2313, \8842_9141 );
and \U$20240 ( \29045_29344 , RIfc498c8_5859, \8844_9143 );
and \U$20241 ( \29046_29345 , RIe14f718_2281, \8846_9145 );
and \U$20242 ( \29047_29346 , RIfcbda70_7180, \8848_9147 );
and \U$20243 ( \29048_29347 , RIe14ca18_2249, \8850_9149 );
and \U$20244 ( \29049_29348 , RIe149d18_2217, \8852_9151 );
and \U$20245 ( \29050_29349 , RIe147018_2185, \8854_9153 );
and \U$20246 ( \29051_29350 , RIee34828_5056, \8856_9155 );
and \U$20247 ( \29052_29351 , RIee33748_5044, \8858_9157 );
and \U$20248 ( \29053_29352 , RIee32668_5032, \8860_9159 );
and \U$20249 ( \29054_29353 , RIee31588_5020, \8862_9161 );
and \U$20250 ( \29055_29354 , RIe1418e8_2123, \8864_9163 );
and \U$20251 ( \29056_29355 , RIe13f458_2097, \8866_9165 );
and \U$20252 ( \29057_29356 , RIdf3d360_2073, \8868_9167 );
and \U$20253 ( \29058_29357 , RIdf3aed0_2047, \8870_9169 );
and \U$20254 ( \29059_29358 , RIfc526d0_5960, \8872_9171 );
and \U$20255 ( \29060_29359 , RIfc42848_5779, \8874_9173 );
and \U$20256 ( \29061_29360 , RIfcae9f8_7009, \8876_9175 );
and \U$20257 ( \29062_29361 , RIfcb7260_7106, \8878_9177 );
and \U$20258 ( \29063_29362 , RIfea42b0_8212, \8880_9179 );
and \U$20259 ( \29064_29363 , RIdf33ce8_1966, \8882_9181 );
and \U$20260 ( \29065_29364 , RIdf31b28_1942, \8884_9183 );
and \U$20261 ( \29066_29365 , RIdf2fc38_1920, \8886_9185 );
or \U$20262 ( \29067_29366 , \29003_29302 , \29004_29303 , \29005_29304 , \29006_29305 , \29007_29306 , \29008_29307 , \29009_29308 , \29010_29309 , \29011_29310 , \29012_29311 , \29013_29312 , \29014_29313 , \29015_29314 , \29016_29315 , \29017_29316 , \29018_29317 , \29019_29318 , \29020_29319 , \29021_29320 , \29022_29321 , \29023_29322 , \29024_29323 , \29025_29324 , \29026_29325 , \29027_29326 , \29028_29327 , \29029_29328 , \29030_29329 , \29031_29330 , \29032_29331 , \29033_29332 , \29034_29333 , \29035_29334 , \29036_29335 , \29037_29336 , \29038_29337 , \29039_29338 , \29040_29339 , \29041_29340 , \29042_29341 , \29043_29342 , \29044_29343 , \29045_29344 , \29046_29345 , \29047_29346 , \29048_29347 , \29049_29348 , \29050_29349 , \29051_29350 , \29052_29351 , \29053_29352 , \29054_29353 , \29055_29354 , \29056_29355 , \29057_29356 , \29058_29357 , \29059_29358 , \29060_29359 , \29061_29360 , \29062_29361 , \29063_29362 , \29064_29363 , \29065_29364 , \29066_29365 );
and \U$20263 ( \29068_29367 , RIee2c3f8_4962, \8889_9188 );
and \U$20264 ( \29069_29368 , RIfc4cfa0_5898, \8891_9190 );
and \U$20265 ( \29070_29369 , RIfc572c0_6014, \8893_9192 );
and \U$20266 ( \29071_29370 , RIfc4f430_5924, \8895_9194 );
and \U$20267 ( \29072_29371 , RIfea3e78_8209, \8897_9196 );
and \U$20268 ( \29073_29372 , RIdf28a50_1839, \8899_9198 );
and \U$20269 ( \29074_29373 , RIdf26b60_1817, \8901_9200 );
and \U$20270 ( \29075_29374 , RIdf250a8_1798, \8903_9202 );
and \U$20271 ( \29076_29375 , RIfc9b600_6790, \8905_9204 );
and \U$20272 ( \29077_29376 , RIfcb9df8_7137, \8907_9206 );
and \U$20273 ( \29078_29377 , RIdf23320_1777, \8909_9208 );
and \U$20274 ( \29079_29378 , RIfc86318_6549, \8911_9210 );
and \U$20275 ( \29080_29379 , RIfeabfd8_8273, \8913_9212 );
and \U$20276 ( \29081_29380 , RIdf201e8_1742, \8915_9214 );
and \U$20277 ( \29082_29381 , RIdf1b5f8_1688, \8917_9216 );
and \U$20278 ( \29083_29382 , RIdf19ca8_1670, \8919_9218 );
and \U$20279 ( \29084_29383 , RIdf17ae8_1646, \8921_9220 );
and \U$20280 ( \29085_29384 , RIdf14de8_1614, \8923_9222 );
and \U$20281 ( \29086_29385 , RIdf120e8_1582, \8925_9224 );
and \U$20282 ( \29087_29386 , RIdf0f3e8_1550, \8927_9226 );
and \U$20283 ( \29088_29387 , RIdf0c6e8_1518, \8929_9228 );
and \U$20284 ( \29089_29388 , RIdf099e8_1486, \8931_9230 );
and \U$20285 ( \29090_29389 , RIdf06ce8_1454, \8933_9232 );
and \U$20286 ( \29091_29390 , RIdf03fe8_1422, \8935_9234 );
and \U$20287 ( \29092_29391 , RIdefe5e8_1358, \8937_9236 );
and \U$20288 ( \29093_29392 , RIdefb8e8_1326, \8939_9238 );
and \U$20289 ( \29094_29393 , RIdef8be8_1294, \8941_9240 );
and \U$20290 ( \29095_29394 , RIdef5ee8_1262, \8943_9242 );
and \U$20291 ( \29096_29395 , RIdef31e8_1230, \8945_9244 );
and \U$20292 ( \29097_29396 , RIdef04e8_1198, \8947_9246 );
and \U$20293 ( \29098_29397 , RIdeed7e8_1166, \8949_9248 );
and \U$20294 ( \29099_29398 , RIdeeaae8_1134, \8951_9250 );
and \U$20295 ( \29100_29399 , RIfc89018_6581, \8953_9252 );
and \U$20296 ( \29101_29400 , RIfcc54c8_7267, \8955_9254 );
and \U$20297 ( \29102_29401 , RIfc89180_6582, \8957_9256 );
and \U$20298 ( \29103_29402 , RIfc4b380_5878, \8959_9258 );
and \U$20299 ( \29104_29403 , RIdee53b8_1072, \8961_9260 );
and \U$20300 ( \29105_29404 , RIdee34c8_1050, \8963_9262 );
and \U$20301 ( \29106_29405 , RIfea3d10_8208, \8965_9264 );
and \U$20302 ( \29107_29406 , RIdedf148_1002, \8967_9266 );
and \U$20303 ( \29108_29407 , RIfcae188_7003, \8969_9268 );
and \U$20304 ( \29109_29408 , RIfc4b0b0_5876, \8971_9270 );
and \U$20305 ( \29110_29409 , RIfc74870_6348, \8973_9272 );
and \U$20306 ( \29111_29410 , RIfce4968_7623, \8975_9274 );
and \U$20307 ( \29112_29411 , RIdeda288_946, \8977_9276 );
and \U$20308 ( \29113_29412 , RIded7c90_919, \8979_9278 );
and \U$20309 ( \29114_29413 , RIded5da0_897, \8981_9280 );
and \U$20310 ( \29115_29414 , RIded3640_869, \8983_9282 );
and \U$20311 ( \29116_29415 , RIded1318_844, \8985_9284 );
and \U$20312 ( \29117_29416 , RIdece618_812, \8987_9286 );
and \U$20313 ( \29118_29417 , RIdecb918_780, \8989_9288 );
and \U$20314 ( \29119_29418 , RIdec8c18_748, \8991_9290 );
and \U$20315 ( \29120_29419 , RIdeb5118_524, \8993_9292 );
and \U$20316 ( \29121_29420 , RIde98360_332, \8995_9294 );
and \U$20317 ( \29122_29421 , RIe16ed20_2638, \8997_9296 );
and \U$20318 ( \29123_29422 , RIe15ab18_2409, \8999_9298 );
and \U$20319 ( \29124_29423 , RIe144318_2153, \9001_9300 );
and \U$20320 ( \29125_29424 , RIdf38d10_2023, \9003_9302 );
and \U$20321 ( \29126_29425 , RIdf2d370_1891, \9005_9304 );
and \U$20322 ( \29127_29426 , RIdf1dbf0_1715, \9007_9306 );
and \U$20323 ( \29128_29427 , RIdf012e8_1390, \9009_9308 );
and \U$20324 ( \29129_29428 , RIdee7de8_1102, \9011_9310 );
and \U$20325 ( \29130_29429 , RIdedcb50_975, \9013_9312 );
and \U$20326 ( \29131_29430 , RIde7e2a8_205, \9015_9314 );
or \U$20327 ( \29132_29431 , \29068_29367 , \29069_29368 , \29070_29369 , \29071_29370 , \29072_29371 , \29073_29372 , \29074_29373 , \29075_29374 , \29076_29375 , \29077_29376 , \29078_29377 , \29079_29378 , \29080_29379 , \29081_29380 , \29082_29381 , \29083_29382 , \29084_29383 , \29085_29384 , \29086_29385 , \29087_29386 , \29088_29387 , \29089_29388 , \29090_29389 , \29091_29390 , \29092_29391 , \29093_29392 , \29094_29393 , \29095_29394 , \29096_29395 , \29097_29396 , \29098_29397 , \29099_29398 , \29100_29399 , \29101_29400 , \29102_29401 , \29103_29402 , \29104_29403 , \29105_29404 , \29106_29405 , \29107_29406 , \29108_29407 , \29109_29408 , \29110_29409 , \29111_29410 , \29112_29411 , \29113_29412 , \29114_29413 , \29115_29414 , \29116_29415 , \29117_29416 , \29118_29417 , \29119_29418 , \29120_29419 , \29121_29420 , \29122_29421 , \29123_29422 , \29124_29423 , \29125_29424 , \29126_29425 , \29127_29426 , \29128_29427 , \29129_29428 , \29130_29429 , \29131_29430 );
or \U$20328 ( \29133_29432 , \29067_29366 , \29132_29431 );
_DC \g233f/U$1 ( \29134 , \29133_29432 , \9024_9323 );
buf \U$20329 ( \29135_29434 , \29134 );
and \U$20330 ( \29136_29435 , RIe19e1b0_3176, \9034_9333 );
and \U$20331 ( \29137_29436 , RIe19b4b0_3144, \9036_9335 );
and \U$20332 ( \29138_29437 , RIfc9cf50_6808, \9038_9337 );
and \U$20333 ( \29139_29438 , RIe1987b0_3112, \9040_9339 );
and \U$20334 ( \29140_29439 , RIfc87290_6560, \9042_9341 );
and \U$20335 ( \29141_29440 , RIe195ab0_3080, \9044_9343 );
and \U$20336 ( \29142_29441 , RIe192db0_3048, \9046_9345 );
and \U$20337 ( \29143_29442 , RIe1900b0_3016, \9048_9347 );
and \U$20338 ( \29144_29443 , RIe18a6b0_2952, \9050_9349 );
and \U$20339 ( \29145_29444 , RIe1879b0_2920, \9052_9351 );
and \U$20340 ( \29146_29445 , RIfc842c0_6526, \9054_9353 );
and \U$20341 ( \29147_29446 , RIe184cb0_2888, \9056_9355 );
and \U$20342 ( \29148_29447 , RIfc83a50_6520, \9058_9357 );
and \U$20343 ( \29149_29448 , RIe181fb0_2856, \9060_9359 );
and \U$20344 ( \29150_29449 , RIe17f2b0_2824, \9062_9361 );
and \U$20345 ( \29151_29450 , RIe17c5b0_2792, \9064_9363 );
and \U$20346 ( \29152_29451 , RIfc9d0b8_6809, \9066_9365 );
and \U$20347 ( \29153_29452 , RIfc9e030_6820, \9068_9367 );
and \U$20348 ( \29154_29453 , RIe177420_2734, \9070_9369 );
and \U$20349 ( \29155_29454 , RIe176340_2722, \9072_9371 );
and \U$20350 ( \29156_29455 , RIfc4f700_5926, \9074_9373 );
and \U$20351 ( \29157_29456 , RIfcc4820_7258, \9076_9375 );
and \U$20352 ( \29158_29457 , RIfc4fb38_5929, \9078_9377 );
and \U$20353 ( \29159_29458 , RIfce8040_7662, \9080_9379 );
and \U$20354 ( \29160_29459 , RIee3c6b8_5146, \9082_9381 );
and \U$20355 ( \29161_29460 , RIee3b308_5132, \9084_9383 );
and \U$20356 ( \29162_29461 , RIfc812f0_6492, \9086_9385 );
and \U$20357 ( \29163_29462 , RIe174180_2698, \9088_9387 );
and \U$20358 ( \29164_29463 , RIfcd3028_7423, \9090_9389 );
and \U$20359 ( \29165_29464 , RIfc7f400_6470, \9092_9391 );
and \U$20360 ( \29166_29465 , RIfc46a60_5826, \9094_9393 );
and \U$20361 ( \29167_29466 , RIfc472d0_5832, \9096_9395 );
and \U$20362 ( \29168_29467 , RIf16cc58_5697, \9098_9397 );
and \U$20363 ( \29169_29468 , RIe224508_4703, \9100_9399 );
and \U$20364 ( \29170_29469 , RIfc7d3a8_6447, \9102_9401 );
and \U$20365 ( \29171_29470 , RIe221808_4671, \9104_9403 );
and \U$20366 ( \29172_29471 , RIfc97c58_6749, \9106_9405 );
and \U$20367 ( \29173_29472 , RIe21eb08_4639, \9108_9407 );
and \U$20368 ( \29174_29473 , RIe219108_4575, \9110_9409 );
and \U$20369 ( \29175_29474 , RIe216408_4543, \9112_9411 );
and \U$20370 ( \29176_29475 , RIfcdbe30_7524, \9114_9413 );
and \U$20371 ( \29177_29476 , RIe213708_4511, \9116_9415 );
and \U$20372 ( \29178_29477 , RIf169580_5658, \9118_9417 );
and \U$20373 ( \29179_29478 , RIe210a08_4479, \9120_9419 );
and \U$20374 ( \29180_29479 , RIfca4570_6892, \9122_9421 );
and \U$20375 ( \29181_29480 , RIe20dd08_4447, \9124_9423 );
and \U$20376 ( \29182_29481 , RIe20b008_4415, \9126_9425 );
and \U$20377 ( \29183_29482 , RIe208308_4383, \9128_9427 );
and \U$20378 ( \29184_29483 , RIfc7b080_6422, \9130_9429 );
and \U$20379 ( \29185_29484 , RIfc59cf0_6044, \9132_9431 );
and \U$20380 ( \29186_29485 , RIfea9b48_8247, \9134_9433 );
and \U$20381 ( \29187_29486 , RIfea4418_8213, \9136_9435 );
and \U$20382 ( \29188_29487 , RIfc79cd0_6408, \9138_9437 );
and \U$20383 ( \29189_29488 , RIfcd19a8_7407, \9140_9439 );
and \U$20384 ( \29190_29489 , RIfcc81c8_7299, \9142_9441 );
and \U$20385 ( \29191_29490 , RIf162230_5576, \9144_9443 );
and \U$20386 ( \29192_29491 , RIf160778_5557, \9146_9445 );
and \U$20387 ( \29193_29492 , RIf15e888_5535, \9148_9447 );
and \U$20388 ( \29194_29493 , RIfea4580_8214, \9150_9449 );
and \U$20389 ( \29195_29494 , RIfea46e8_8215, \9152_9451 );
and \U$20390 ( \29196_29495 , RIfc77f48_6387, \9154_9453 );
and \U$20391 ( \29197_29496 , RIfc41fd8_5773, \9156_9455 );
and \U$20392 ( \29198_29497 , RIf15aaa8_5491, \9158_9457 );
and \U$20393 ( \29199_29498 , RIfc7c430_6436, \9160_9459 );
or \U$20394 ( \29200_29499 , \29136_29435 , \29137_29436 , \29138_29437 , \29139_29438 , \29140_29439 , \29141_29440 , \29142_29441 , \29143_29442 , \29144_29443 , \29145_29444 , \29146_29445 , \29147_29446 , \29148_29447 , \29149_29448 , \29150_29449 , \29151_29450 , \29152_29451 , \29153_29452 , \29154_29453 , \29155_29454 , \29156_29455 , \29157_29456 , \29158_29457 , \29159_29458 , \29160_29459 , \29161_29460 , \29162_29461 , \29163_29462 , \29164_29463 , \29165_29464 , \29166_29465 , \29167_29466 , \29168_29467 , \29169_29468 , \29170_29469 , \29171_29470 , \29172_29471 , \29173_29472 , \29174_29473 , \29175_29474 , \29176_29475 , \29177_29476 , \29178_29477 , \29179_29478 , \29180_29479 , \29181_29480 , \29182_29481 , \29183_29482 , \29184_29483 , \29185_29484 , \29186_29485 , \29187_29486 , \29188_29487 , \29189_29488 , \29190_29489 , \29191_29490 , \29192_29491 , \29193_29492 , \29194_29493 , \29195_29494 , \29196_29495 , \29197_29496 , \29198_29497 , \29199_29498 );
and \U$20395 ( \29201_29500 , RIf159158_5473, \9163_9462 );
and \U$20396 ( \29202_29501 , RIf157f10_5460, \9165_9464 );
and \U$20397 ( \29203_29502 , RIfcae890_7008, \9167_9466 );
and \U$20398 ( \29204_29503 , RIe1faa78_4229, \9169_9468 );
and \U$20399 ( \29205_29504 , RIfc4a840_5870, \9171_9470 );
and \U$20400 ( \29206_29505 , RIfc4ed28_5919, \9173_9472 );
and \U$20401 ( \29207_29506 , RIfce0e58_7581, \9175_9474 );
and \U$20402 ( \29208_29507 , RIe1f5ff0_4176, \9177_9476 );
and \U$20403 ( \29209_29508 , RIf153758_5409, \9179_9478 );
and \U$20404 ( \29210_29509 , RIf151f70_5392, \9181_9480 );
and \U$20405 ( \29211_29510 , RIfccb468_7335, \9183_9482 );
and \U$20406 ( \29212_29511 , RIe1f3cc8_4151, \9185_9484 );
and \U$20407 ( \29213_29512 , RIfc68ed0_6216, \9187_9486 );
and \U$20408 ( \29214_29513 , RIfc6d250_6264, \9189_9488 );
and \U$20409 ( \29215_29514 , RIfca9ca0_6954, \9191_9490 );
and \U$20410 ( \29216_29515 , RIe1ee9d0_4092, \9193_9492 );
and \U$20411 ( \29217_29516 , RIe1ec270_4064, \9195_9494 );
and \U$20412 ( \29218_29517 , RIe1e9570_4032, \9197_9496 );
and \U$20413 ( \29219_29518 , RIe1e6870_4000, \9199_9498 );
and \U$20414 ( \29220_29519 , RIe1e3b70_3968, \9201_9500 );
and \U$20415 ( \29221_29520 , RIe1e0e70_3936, \9203_9502 );
and \U$20416 ( \29222_29521 , RIe1de170_3904, \9205_9504 );
and \U$20417 ( \29223_29522 , RIe1db470_3872, \9207_9506 );
and \U$20418 ( \29224_29523 , RIe1d8770_3840, \9209_9508 );
and \U$20419 ( \29225_29524 , RIe1d2d70_3776, \9211_9510 );
and \U$20420 ( \29226_29525 , RIe1d0070_3744, \9213_9512 );
and \U$20421 ( \29227_29526 , RIe1cd370_3712, \9215_9514 );
and \U$20422 ( \29228_29527 , RIe1ca670_3680, \9217_9516 );
and \U$20423 ( \29229_29528 , RIe1c7970_3648, \9219_9518 );
and \U$20424 ( \29230_29529 , RIe1c4c70_3616, \9221_9520 );
and \U$20425 ( \29231_29530 , RIe1c1f70_3584, \9223_9522 );
and \U$20426 ( \29232_29531 , RIe1bf270_3552, \9225_9524 );
and \U$20427 ( \29233_29532 , RIfc784e8_6391, \9227_9526 );
and \U$20428 ( \29234_29533 , RIfcbef88_7195, \9229_9528 );
and \U$20429 ( \29235_29534 , RIe1b9ca8_3491, \9231_9530 );
and \U$20430 ( \29236_29535 , RIe1b7ae8_3467, \9233_9532 );
and \U$20431 ( \29237_29536 , RIfcc20c0_7230, \9235_9534 );
and \U$20432 ( \29238_29537 , RIfca6190_6912, \9237_9536 );
and \U$20433 ( \29239_29538 , RIe1b5928_3443, \9239_9538 );
and \U$20434 ( \29240_29539 , RIe1b4410_3428, \9241_9540 );
and \U$20435 ( \29241_29540 , RIfcb81d8_7117, \9243_9542 );
and \U$20436 ( \29242_29541 , RIfcc5090_7264, \9245_9544 );
and \U$20437 ( \29243_29542 , RIe1b2d90_3412, \9247_9546 );
and \U$20438 ( \29244_29543 , RIe1b1440_3394, \9249_9548 );
and \U$20439 ( \29245_29544 , RIfcd5350_7448, \9251_9550 );
and \U$20440 ( \29246_29545 , RIfcb9588_7131, \9253_9552 );
and \U$20441 ( \29247_29546 , RIe1acc88_3343, \9255_9554 );
and \U$20442 ( \29248_29547 , RIe1ab4a0_3326, \9257_9556 );
and \U$20443 ( \29249_29548 , RIe1a95b0_3304, \9259_9558 );
and \U$20444 ( \29250_29549 , RIe1a68b0_3272, \9261_9560 );
and \U$20445 ( \29251_29550 , RIe1a3bb0_3240, \9263_9562 );
and \U$20446 ( \29252_29551 , RIe1a0eb0_3208, \9265_9564 );
and \U$20447 ( \29253_29552 , RIe18d3b0_2984, \9267_9566 );
and \U$20448 ( \29254_29553 , RIe1798b0_2760, \9269_9568 );
and \U$20449 ( \29255_29554 , RIe227208_4735, \9271_9570 );
and \U$20450 ( \29256_29555 , RIe21be08_4607, \9273_9572 );
and \U$20451 ( \29257_29556 , RIe205608_4351, \9275_9574 );
and \U$20452 ( \29258_29557 , RIe1ff668_4283, \9277_9576 );
and \U$20453 ( \29259_29558 , RIe1f8a20_4206, \9279_9578 );
and \U$20454 ( \29260_29559 , RIe1f1568_4123, \9281_9580 );
and \U$20455 ( \29261_29560 , RIe1d5a70_3808, \9283_9582 );
and \U$20456 ( \29262_29561 , RIe1bc570_3520, \9285_9584 );
and \U$20457 ( \29263_29562 , RIe1af3e8_3371, \9287_9586 );
and \U$20458 ( \29264_29563 , RIe171a20_2670, \9289_9588 );
or \U$20459 ( \29265_29564 , \29201_29500 , \29202_29501 , \29203_29502 , \29204_29503 , \29205_29504 , \29206_29505 , \29207_29506 , \29208_29507 , \29209_29508 , \29210_29509 , \29211_29510 , \29212_29511 , \29213_29512 , \29214_29513 , \29215_29514 , \29216_29515 , \29217_29516 , \29218_29517 , \29219_29518 , \29220_29519 , \29221_29520 , \29222_29521 , \29223_29522 , \29224_29523 , \29225_29524 , \29226_29525 , \29227_29526 , \29228_29527 , \29229_29528 , \29230_29529 , \29231_29530 , \29232_29531 , \29233_29532 , \29234_29533 , \29235_29534 , \29236_29535 , \29237_29536 , \29238_29537 , \29239_29538 , \29240_29539 , \29241_29540 , \29242_29541 , \29243_29542 , \29244_29543 , \29245_29544 , \29246_29545 , \29247_29546 , \29248_29547 , \29249_29548 , \29250_29549 , \29251_29550 , \29252_29551 , \29253_29552 , \29254_29553 , \29255_29554 , \29256_29555 , \29257_29556 , \29258_29557 , \29259_29558 , \29260_29559 , \29261_29560 , \29262_29561 , \29263_29562 , \29264_29563 );
or \U$20460 ( \29266_29565 , \29200_29499 , \29265_29564 );
_DC \g346c/U$1 ( \29267 , \29266_29565 , \9298_9597 );
buf \U$20461 ( \29268_29567 , \29267 );
xor \U$20462 ( \29269_29568 , \29135_29434 , \29268_29567 );
and \U$20463 ( \29270_29569 , RIdec5db0_715, \8760_9059 );
and \U$20464 ( \29271_29570 , RIdec30b0_683, \8762_9061 );
and \U$20465 ( \29272_29571 , RIee201e8_4824, \8764_9063 );
and \U$20466 ( \29273_29572 , RIdec03b0_651, \8766_9065 );
and \U$20467 ( \29274_29573 , RIfcaf538_7017, \8768_9067 );
and \U$20468 ( \29275_29574 , RIdebd6b0_619, \8770_9069 );
and \U$20469 ( \29276_29575 , RIdeba9b0_587, \8772_9071 );
and \U$20470 ( \29277_29576 , RIdeb7cb0_555, \8774_9073 );
and \U$20471 ( \29278_29577 , RIfc40fe8_5765, \8776_9075 );
and \U$20472 ( \29279_29578 , RIdeb22b0_491, \8778_9077 );
and \U$20473 ( \29280_29579 , RIfcd08c8_7395, \8780_9079 );
and \U$20474 ( \29281_29580 , RIdeaf5b0_459, \8782_9081 );
and \U$20475 ( \29282_29581 , RIee1dd58_4798, \8784_9083 );
and \U$20476 ( \29283_29582 , RIdeabb18_427, \8786_9085 );
and \U$20477 ( \29284_29583 , RIdea5218_395, \8788_9087 );
and \U$20478 ( \29285_29584 , RIde9e918_363, \8790_9089 );
and \U$20479 ( \29286_29585 , RIee1d218_4790, \8792_9091 );
and \U$20480 ( \29287_29586 , RIfcedd10_7728, \8794_9093 );
and \U$20481 ( \29288_29587 , RIfce62b8_7641, \8796_9095 );
and \U$20482 ( \29289_29588 , RIfcc92a8_7311, \8798_9097 );
and \U$20483 ( \29290_29589 , RIde91da8_301, \8800_9099 );
and \U$20484 ( \29291_29590 , RIde8e928_285, \8802_9101 );
and \U$20485 ( \29292_29591 , RIde8a788_265, \8804_9103 );
and \U$20486 ( \29293_29592 , RIde865e8_245, \8806_9105 );
and \U$20487 ( \29294_29593 , RIde82448_225, \8808_9107 );
and \U$20488 ( \29295_29594 , RIfea1448_8179, \8810_9109 );
and \U$20489 ( \29296_29595 , RIfc750e0_6354, \8812_9111 );
and \U$20490 ( \29297_29596 , RIfcc19b8_7225, \8814_9113 );
and \U$20491 ( \29298_29597 , RIfced8d8_7725, \8816_9115 );
and \U$20492 ( \29299_29598 , RIfec5eb0_8372, \8818_9117 );
and \U$20493 ( \29300_29599 , RIe169fc8_2583, \8820_9119 );
and \U$20494 ( \29301_29600 , RIe168678_2565, \8822_9121 );
and \U$20495 ( \29302_29601 , RIe165db0_2536, \8824_9123 );
and \U$20496 ( \29303_29602 , RIe1630b0_2504, \8826_9125 );
and \U$20497 ( \29304_29603 , RIfccfc20_7386, \8828_9127 );
and \U$20498 ( \29305_29604 , RIe1603b0_2472, \8830_9129 );
and \U$20499 ( \29306_29605 , RIee365b0_5077, \8832_9131 );
and \U$20500 ( \29307_29606 , RIe15d6b0_2440, \8834_9133 );
and \U$20501 ( \29308_29607 , RIe157cb0_2376, \8836_9135 );
and \U$20502 ( \29309_29608 , RIe154fb0_2344, \8838_9137 );
and \U$20503 ( \29310_29609 , RIfea1718_8181, \8840_9139 );
and \U$20504 ( \29311_29610 , RIe1522b0_2312, \8842_9141 );
and \U$20505 ( \29312_29611 , RIee35200_5063, \8844_9143 );
and \U$20506 ( \29313_29612 , RIe14f5b0_2280, \8846_9145 );
and \U$20507 ( \29314_29613 , RIfcb0348_7027, \8848_9147 );
and \U$20508 ( \29315_29614 , RIe14c8b0_2248, \8850_9149 );
and \U$20509 ( \29316_29615 , RIe149bb0_2216, \8852_9151 );
and \U$20510 ( \29317_29616 , RIe146eb0_2184, \8854_9153 );
and \U$20511 ( \29318_29617 , RIfc73790_6336, \8856_9155 );
and \U$20512 ( \29319_29618 , RIfcdf238_7561, \8858_9157 );
and \U$20513 ( \29320_29619 , RIee32500_5031, \8860_9159 );
and \U$20514 ( \29321_29620 , RIfc94f58_6717, \8862_9161 );
and \U$20515 ( \29322_29621 , RIe141780_2122, \8864_9163 );
and \U$20516 ( \29323_29622 , RIe13f2f0_2096, \8866_9165 );
and \U$20517 ( \29324_29623 , RIfec5be0_8370, \8868_9167 );
and \U$20518 ( \29325_29624 , RIdf3ad68_2046, \8870_9169 );
and \U$20519 ( \29326_29625 , RIfea15b0_8180, \8872_9171 );
and \U$20520 ( \29327_29626 , RIfc5fb28_6111, \8874_9173 );
and \U$20521 ( \29328_29627 , RIfcae728_7007, \8876_9175 );
and \U$20522 ( \29329_29628 , RIfc74438_6345, \8878_9177 );
and \U$20523 ( \29330_29629 , RIdf36178_1992, \8880_9179 );
and \U$20524 ( \29331_29630 , RIdf33b80_1965, \8882_9181 );
and \U$20525 ( \29332_29631 , RIdf319c0_1941, \8884_9183 );
and \U$20526 ( \29333_29632 , RIdf2fad0_1919, \8886_9185 );
or \U$20527 ( \29334_29633 , \29270_29569 , \29271_29570 , \29272_29571 , \29273_29572 , \29274_29573 , \29275_29574 , \29276_29575 , \29277_29576 , \29278_29577 , \29279_29578 , \29280_29579 , \29281_29580 , \29282_29581 , \29283_29582 , \29284_29583 , \29285_29584 , \29286_29585 , \29287_29586 , \29288_29587 , \29289_29588 , \29290_29589 , \29291_29590 , \29292_29591 , \29293_29592 , \29294_29593 , \29295_29594 , \29296_29595 , \29297_29596 , \29298_29597 , \29299_29598 , \29300_29599 , \29301_29600 , \29302_29601 , \29303_29602 , \29304_29603 , \29305_29604 , \29306_29605 , \29307_29606 , \29308_29607 , \29309_29608 , \29310_29609 , \29311_29610 , \29312_29611 , \29313_29612 , \29314_29613 , \29315_29614 , \29316_29615 , \29317_29616 , \29318_29617 , \29319_29618 , \29320_29619 , \29321_29620 , \29322_29621 , \29323_29622 , \29324_29623 , \29325_29624 , \29326_29625 , \29327_29626 , \29328_29627 , \29329_29628 , \29330_29629 , \29331_29630 , \29332_29631 , \29333_29632 );
and \U$20528 ( \29335_29634 , RIee2c290_4961, \8889_9188 );
and \U$20529 ( \29336_29635 , RIee2a940_4943, \8891_9190 );
and \U$20530 ( \29337_29636 , RIfc70658_6301, \8893_9192 );
and \U$20531 ( \29338_29637 , RIfc704f0_6300, \8895_9194 );
and \U$20532 ( \29339_29638 , RIdf2aaa8_1862, \8897_9196 );
and \U$20533 ( \29340_29639 , RIdf288e8_1838, \8899_9198 );
and \U$20534 ( \29341_29640 , RIdf269f8_1816, \8901_9200 );
and \U$20535 ( \29342_29641 , RIdf24f40_1797, \8903_9202 );
and \U$20536 ( \29343_29642 , RIfc64b50_6168, \8905_9204 );
and \U$20537 ( \29344_29643 , RIfccaa90_7328, \8907_9206 );
and \U$20538 ( \29345_29644 , RIdf231b8_1776, \8909_9208 );
and \U$20539 ( \29346_29645 , RIfcad4e0_6994, \8911_9210 );
and \U$20540 ( \29347_29646 , RIdf21ca0_1761, \8913_9212 );
and \U$20541 ( \29348_29647 , RIfeaad90_8260, \8915_9214 );
and \U$20542 ( \29349_29648 , RIdf1b490_1687, \8917_9216 );
and \U$20543 ( \29350_29649 , RIdf19b40_1669, \8919_9218 );
and \U$20544 ( \29351_29650 , RIdf17980_1645, \8921_9220 );
and \U$20545 ( \29352_29651 , RIdf14c80_1613, \8923_9222 );
and \U$20546 ( \29353_29652 , RIdf11f80_1581, \8925_9224 );
and \U$20547 ( \29354_29653 , RIdf0f280_1549, \8927_9226 );
and \U$20548 ( \29355_29654 , RIdf0c580_1517, \8929_9228 );
and \U$20549 ( \29356_29655 , RIdf09880_1485, \8931_9230 );
and \U$20550 ( \29357_29656 , RIdf06b80_1453, \8933_9232 );
and \U$20551 ( \29358_29657 , RIdf03e80_1421, \8935_9234 );
and \U$20552 ( \29359_29658 , RIdefe480_1357, \8937_9236 );
and \U$20553 ( \29360_29659 , RIdefb780_1325, \8939_9238 );
and \U$20554 ( \29361_29660 , RIdef8a80_1293, \8941_9240 );
and \U$20555 ( \29362_29661 , RIdef5d80_1261, \8943_9242 );
and \U$20556 ( \29363_29662 , RIdef3080_1229, \8945_9244 );
and \U$20557 ( \29364_29663 , RIdef0380_1197, \8947_9246 );
and \U$20558 ( \29365_29664 , RIdeed680_1165, \8949_9248 );
and \U$20559 ( \29366_29665 , RIdeea980_1133, \8951_9250 );
and \U$20560 ( \29367_29666 , RIfc595e8_6039, \8953_9252 );
and \U$20561 ( \29368_29667 , RIfcac568_6983, \8955_9254 );
and \U$20562 ( \29369_29668 , RIfcccf20_7354, \8957_9256 );
and \U$20563 ( \29370_29669 , RIfccd358_7357, \8959_9258 );
and \U$20564 ( \29371_29670 , RIdee5250_1071, \8961_9260 );
and \U$20565 ( \29372_29671 , RIfea7f28_8227, \8963_9262 );
and \U$20566 ( \29373_29672 , RIdee11a0_1025, \8965_9264 );
and \U$20567 ( \29374_29673 , RIfea12e0_8178, \8967_9266 );
and \U$20568 ( \29375_29674 , RIfc679b8_6201, \8969_9268 );
and \U$20569 ( \29376_29675 , RIee22510_4849, \8971_9270 );
and \U$20570 ( \29377_29676 , RIfc6dd90_6272, \8973_9272 );
and \U$20571 ( \29378_29677 , RIfc6cb48_6259, \8975_9274 );
and \U$20572 ( \29379_29678 , RIdeda120_945, \8977_9276 );
and \U$20573 ( \29380_29679 , RIded7b28_918, \8979_9278 );
and \U$20574 ( \29381_29680 , RIded5c38_896, \8981_9280 );
and \U$20575 ( \29382_29681 , RIfec5d48_8371, \8983_9282 );
and \U$20576 ( \29383_29682 , RIded11b0_843, \8985_9284 );
and \U$20577 ( \29384_29683 , RIdece4b0_811, \8987_9286 );
and \U$20578 ( \29385_29684 , RIdecb7b0_779, \8989_9288 );
and \U$20579 ( \29386_29685 , RIdec8ab0_747, \8991_9290 );
and \U$20580 ( \29387_29686 , RIdeb4fb0_523, \8993_9292 );
and \U$20581 ( \29388_29687 , RIde98018_331, \8995_9294 );
and \U$20582 ( \29389_29688 , RIe16ebb8_2637, \8997_9296 );
and \U$20583 ( \29390_29689 , RIe15a9b0_2408, \8999_9298 );
and \U$20584 ( \29391_29690 , RIe1441b0_2152, \9001_9300 );
and \U$20585 ( \29392_29691 , RIdf38ba8_2022, \9003_9302 );
and \U$20586 ( \29393_29692 , RIdf2d208_1890, \9005_9304 );
and \U$20587 ( \29394_29693 , RIdf1da88_1714, \9007_9306 );
and \U$20588 ( \29395_29694 , RIdf01180_1389, \9009_9308 );
and \U$20589 ( \29396_29695 , RIdee7c80_1101, \9011_9310 );
and \U$20590 ( \29397_29696 , RIdedc9e8_974, \9013_9312 );
and \U$20591 ( \29398_29697 , RIde7df60_204, \9015_9314 );
or \U$20592 ( \29399_29698 , \29335_29634 , \29336_29635 , \29337_29636 , \29338_29637 , \29339_29638 , \29340_29639 , \29341_29640 , \29342_29641 , \29343_29642 , \29344_29643 , \29345_29644 , \29346_29645 , \29347_29646 , \29348_29647 , \29349_29648 , \29350_29649 , \29351_29650 , \29352_29651 , \29353_29652 , \29354_29653 , \29355_29654 , \29356_29655 , \29357_29656 , \29358_29657 , \29359_29658 , \29360_29659 , \29361_29660 , \29362_29661 , \29363_29662 , \29364_29663 , \29365_29664 , \29366_29665 , \29367_29666 , \29368_29667 , \29369_29668 , \29370_29669 , \29371_29670 , \29372_29671 , \29373_29672 , \29374_29673 , \29375_29674 , \29376_29675 , \29377_29676 , \29378_29677 , \29379_29678 , \29380_29679 , \29381_29680 , \29382_29681 , \29383_29682 , \29384_29683 , \29385_29684 , \29386_29685 , \29387_29686 , \29388_29687 , \29389_29688 , \29390_29689 , \29391_29690 , \29392_29691 , \29393_29692 , \29394_29693 , \29395_29694 , \29396_29695 , \29397_29696 , \29398_29697 );
or \U$20593 ( \29400_29699 , \29334_29633 , \29399_29698 );
_DC \g23c4/U$1 ( \29401 , \29400_29699 , \9024_9323 );
buf \U$20594 ( \29402_29701 , \29401 );
and \U$20595 ( \29403_29702 , RIe19e048_3175, \9034_9333 );
and \U$20596 ( \29404_29703 , RIe19b348_3143, \9036_9335 );
and \U$20597 ( \29405_29704 , RIfcc3ce0_7250, \9038_9337 );
and \U$20598 ( \29406_29705 , RIe198648_3111, \9040_9339 );
and \U$20599 ( \29407_29706 , RIfc7efc8_6467, \9042_9341 );
and \U$20600 ( \29408_29707 , RIe195948_3079, \9044_9343 );
and \U$20601 ( \29409_29708 , RIe192c48_3047, \9046_9345 );
and \U$20602 ( \29410_29709 , RIe18ff48_3015, \9048_9347 );
and \U$20603 ( \29411_29710 , RIe18a548_2951, \9050_9349 );
and \U$20604 ( \29412_29711 , RIe187848_2919, \9052_9351 );
and \U$20605 ( \29413_29712 , RIfc46790_5824, \9054_9353 );
and \U$20606 ( \29414_29713 , RIe184b48_2887, \9056_9355 );
and \U$20607 ( \29415_29714 , RIfc98d38_6761, \9058_9357 );
and \U$20608 ( \29416_29715 , RIe181e48_2855, \9060_9359 );
and \U$20609 ( \29417_29716 , RIe17f148_2823, \9062_9361 );
and \U$20610 ( \29418_29717 , RIe17c448_2791, \9064_9363 );
and \U$20611 ( \29419_29718 , RIfcb5d48_7091, \9066_9365 );
and \U$20612 ( \29420_29719 , RIfc995a8_6767, \9068_9367 );
and \U$20613 ( \29421_29720 , RIfc9a3b8_6777, \9070_9369 );
and \U$20614 ( \29422_29721 , RIe1761d8_2721, \9072_9371 );
and \U$20615 ( \29423_29722 , RIfc54188_5979, \9074_9373 );
and \U$20616 ( \29424_29723 , RIfcd2bf0_7420, \9076_9375 );
and \U$20617 ( \29425_29724 , RIfc8b778_6609, \9078_9377 );
and \U$20618 ( \29426_29725 , RIfc7dee8_6455, \9080_9379 );
and \U$20619 ( \29427_29726 , RIee3c550_5145, \9082_9381 );
and \U$20620 ( \29428_29727 , RIfc8c420_6618, \9084_9383 );
and \U$20621 ( \29429_29728 , RIee3a0c0_5119, \9086_9385 );
and \U$20622 ( \29430_29729 , RIfeaba38_8269, \9088_9387 );
and \U$20623 ( \29431_29730 , RIfc46628_5823, \9090_9389 );
and \U$20624 ( \29432_29731 , RIfcbc288_7163, \9092_9391 );
and \U$20625 ( \29433_29732 , RIf16e710_5716, \9094_9393 );
and \U$20626 ( \29434_29733 , RIfc8fdc8_6659, \9096_9395 );
and \U$20627 ( \29435_29734 , RIfc48c20_5850, \9098_9397 );
and \U$20628 ( \29436_29735 , RIe2243a0_4702, \9100_9399 );
and \U$20629 ( \29437_29736 , RIfca0358_6845, \9102_9401 );
and \U$20630 ( \29438_29737 , RIe2216a0_4670, \9104_9403 );
and \U$20631 ( \29439_29738 , RIfc9a688_6779, \9106_9405 );
and \U$20632 ( \29440_29739 , RIe21e9a0_4638, \9108_9407 );
and \U$20633 ( \29441_29740 , RIe218fa0_4574, \9110_9409 );
and \U$20634 ( \29442_29741 , RIe2162a0_4542, \9112_9411 );
and \U$20635 ( \29443_29742 , RIfc456b0_5812, \9114_9413 );
and \U$20636 ( \29444_29743 , RIe2135a0_4510, \9116_9415 );
and \U$20637 ( \29445_29744 , RIf169418_5657, \9118_9417 );
and \U$20638 ( \29446_29745 , RIe2108a0_4478, \9120_9419 );
and \U$20639 ( \29447_29746 , RIfc8bfe8_6615, \9122_9421 );
and \U$20640 ( \29448_29747 , RIe20dba0_4446, \9124_9423 );
and \U$20641 ( \29449_29748 , RIe20aea0_4414, \9126_9425 );
and \U$20642 ( \29450_29749 , RIe2081a0_4382, \9128_9427 );
and \U$20643 ( \29451_29750 , RIfc8c9c0_6622, \9130_9429 );
and \U$20644 ( \29452_29751 , RIfc7f568_6471, \9132_9431 );
and \U$20645 ( \29453_29752 , RIe202d40_4322, \9134_9433 );
and \U$20646 ( \29454_29753 , RIe201120_4302, \9136_9435 );
and \U$20647 ( \29455_29754 , RIfce2910_7600, \9138_9437 );
and \U$20648 ( \29456_29755 , RIfc487e8_5847, \9140_9439 );
and \U$20649 ( \29457_29756 , RIfc46d30_5828, \9142_9441 );
and \U$20650 ( \29458_29757 , RIfc992d8_6765, \9144_9443 );
and \U$20651 ( \29459_29758 , RIfca2680_6870, \9146_9445 );
and \U$20652 ( \29460_29759 , RIfc44a08_5803, \9148_9447 );
and \U$20653 ( \29461_29760 , RIe1fd1d8_4257, \9150_9449 );
and \U$20654 ( \29462_29761 , RIe1fbf90_4244, \9152_9451 );
and \U$20655 ( \29463_29762 , RIfc580d0_6024, \9154_9453 );
and \U$20656 ( \29464_29763 , RIfcbdbd8_7181, \9156_9455 );
and \U$20657 ( \29465_29764 , RIfc8dd70_6636, \9158_9457 );
and \U$20658 ( \29466_29765 , RIfce01b0_7572, \9160_9459 );
or \U$20659 ( \29467_29766 , \29403_29702 , \29404_29703 , \29405_29704 , \29406_29705 , \29407_29706 , \29408_29707 , \29409_29708 , \29410_29709 , \29411_29710 , \29412_29711 , \29413_29712 , \29414_29713 , \29415_29714 , \29416_29715 , \29417_29716 , \29418_29717 , \29419_29718 , \29420_29719 , \29421_29720 , \29422_29721 , \29423_29722 , \29424_29723 , \29425_29724 , \29426_29725 , \29427_29726 , \29428_29727 , \29429_29728 , \29430_29729 , \29431_29730 , \29432_29731 , \29433_29732 , \29434_29733 , \29435_29734 , \29436_29735 , \29437_29736 , \29438_29737 , \29439_29738 , \29440_29739 , \29441_29740 , \29442_29741 , \29443_29742 , \29444_29743 , \29445_29744 , \29446_29745 , \29447_29746 , \29448_29747 , \29449_29748 , \29450_29749 , \29451_29750 , \29452_29751 , \29453_29752 , \29454_29753 , \29455_29754 , \29456_29755 , \29457_29756 , \29458_29757 , \29459_29758 , \29460_29759 , \29461_29760 , \29462_29761 , \29463_29762 , \29464_29763 , \29465_29764 , \29466_29765 );
and \U$20660 ( \29468_29767 , RIfc7bbc0_6430, \9163_9462 );
and \U$20661 ( \29469_29768 , RIfc90368_6663, \9165_9464 );
and \U$20662 ( \29470_29769 , RIfc7b8f0_6428, \9167_9466 );
and \U$20663 ( \29471_29770 , RIe1fa910_4228, \9169_9468 );
and \U$20664 ( \29472_29771 , RIfcd8b90_7488, \9171_9470 );
and \U$20665 ( \29473_29772 , RIfc43ec8_5795, \9173_9472 );
and \U$20666 ( \29474_29773 , RIfc7b788_6427, \9175_9474 );
and \U$20667 ( \29475_29774 , RIe1f5e88_4175, \9177_9476 );
and \U$20668 ( \29476_29775 , RIfc7b350_6424, \9179_9478 );
and \U$20669 ( \29477_29776 , RIfc90d40_6670, \9181_9480 );
and \U$20670 ( \29478_29777 , RIfca3490_6880, \9183_9482 );
and \U$20671 ( \29479_29778 , RIe1f3b60_4150, \9185_9484 );
and \U$20672 ( \29480_29779 , RIfc91010_6672, \9187_9486 );
and \U$20673 ( \29481_29780 , RIfcdb728_7519, \9189_9488 );
and \U$20674 ( \29482_29781 , RIfcd8758_7485, \9191_9490 );
and \U$20675 ( \29483_29782 , RIe1ee868_4091, \9193_9492 );
and \U$20676 ( \29484_29783 , RIe1ec108_4063, \9195_9494 );
and \U$20677 ( \29485_29784 , RIe1e9408_4031, \9197_9496 );
and \U$20678 ( \29486_29785 , RIe1e6708_3999, \9199_9498 );
and \U$20679 ( \29487_29786 , RIe1e3a08_3967, \9201_9500 );
and \U$20680 ( \29488_29787 , RIe1e0d08_3935, \9203_9502 );
and \U$20681 ( \29489_29788 , RIe1de008_3903, \9205_9504 );
and \U$20682 ( \29490_29789 , RIe1db308_3871, \9207_9506 );
and \U$20683 ( \29491_29790 , RIe1d8608_3839, \9209_9508 );
and \U$20684 ( \29492_29791 , RIe1d2c08_3775, \9211_9510 );
and \U$20685 ( \29493_29792 , RIe1cff08_3743, \9213_9512 );
and \U$20686 ( \29494_29793 , RIe1cd208_3711, \9215_9514 );
and \U$20687 ( \29495_29794 , RIe1ca508_3679, \9217_9516 );
and \U$20688 ( \29496_29795 , RIe1c7808_3647, \9219_9518 );
and \U$20689 ( \29497_29796 , RIe1c4b08_3615, \9221_9520 );
and \U$20690 ( \29498_29797 , RIe1c1e08_3583, \9223_9522 );
and \U$20691 ( \29499_29798 , RIe1bf108_3551, \9225_9524 );
and \U$20692 ( \29500_29799 , RIf14cf48_5335, \9227_9526 );
and \U$20693 ( \29501_29800 , RIfc78d58_6397, \9229_9528 );
and \U$20694 ( \29502_29801 , RIe1b9b40_3490, \9231_9530 );
and \U$20695 ( \29503_29802 , RIfec5910_8368, \9233_9532 );
and \U$20696 ( \29504_29803 , RIfc78a88_6395, \9235_9534 );
and \U$20697 ( \29505_29804 , RIfcd51e8_7447, \9237_9536 );
and \U$20698 ( \29506_29805 , RIe1b57c0_3442, \9239_9538 );
and \U$20699 ( \29507_29806 , RIfea1010_8176, \9241_9540 );
and \U$20700 ( \29508_29807 , RIf1492d0_5292, \9243_9542 );
and \U$20701 ( \29509_29808 , RIfec5a78_8369, \9245_9544 );
and \U$20702 ( \29510_29809 , RIe1b2c28_3411, \9247_9546 );
and \U$20703 ( \29511_29810 , RIe1b12d8_3393, \9249_9548 );
and \U$20704 ( \29512_29811 , RIfec5640_8366, \9251_9550 );
and \U$20705 ( \29513_29812 , RIf146a08_5263, \9253_9552 );
and \U$20706 ( \29514_29813 , RIfec57a8_8367, \9255_9554 );
and \U$20707 ( \29515_29814 , RIfea1178_8177, \9257_9556 );
and \U$20708 ( \29516_29815 , RIe1a9448_3303, \9259_9558 );
and \U$20709 ( \29517_29816 , RIe1a6748_3271, \9261_9560 );
and \U$20710 ( \29518_29817 , RIe1a3a48_3239, \9263_9562 );
and \U$20711 ( \29519_29818 , RIe1a0d48_3207, \9265_9564 );
and \U$20712 ( \29520_29819 , RIe18d248_2983, \9267_9566 );
and \U$20713 ( \29521_29820 , RIe179748_2759, \9269_9568 );
and \U$20714 ( \29522_29821 , RIe2270a0_4734, \9271_9570 );
and \U$20715 ( \29523_29822 , RIe21bca0_4606, \9273_9572 );
and \U$20716 ( \29524_29823 , RIe2054a0_4350, \9275_9574 );
and \U$20717 ( \29525_29824 , RIe1ff500_4282, \9277_9576 );
and \U$20718 ( \29526_29825 , RIe1f88b8_4205, \9279_9578 );
and \U$20719 ( \29527_29826 , RIe1f1400_4122, \9281_9580 );
and \U$20720 ( \29528_29827 , RIe1d5908_3807, \9283_9582 );
and \U$20721 ( \29529_29828 , RIe1bc408_3519, \9285_9584 );
and \U$20722 ( \29530_29829 , RIe1af280_3370, \9287_9586 );
and \U$20723 ( \29531_29830 , RIe1718b8_2669, \9289_9588 );
or \U$20724 ( \29532_29831 , \29468_29767 , \29469_29768 , \29470_29769 , \29471_29770 , \29472_29771 , \29473_29772 , \29474_29773 , \29475_29774 , \29476_29775 , \29477_29776 , \29478_29777 , \29479_29778 , \29480_29779 , \29481_29780 , \29482_29781 , \29483_29782 , \29484_29783 , \29485_29784 , \29486_29785 , \29487_29786 , \29488_29787 , \29489_29788 , \29490_29789 , \29491_29790 , \29492_29791 , \29493_29792 , \29494_29793 , \29495_29794 , \29496_29795 , \29497_29796 , \29498_29797 , \29499_29798 , \29500_29799 , \29501_29800 , \29502_29801 , \29503_29802 , \29504_29803 , \29505_29804 , \29506_29805 , \29507_29806 , \29508_29807 , \29509_29808 , \29510_29809 , \29511_29810 , \29512_29811 , \29513_29812 , \29514_29813 , \29515_29814 , \29516_29815 , \29517_29816 , \29518_29817 , \29519_29818 , \29520_29819 , \29521_29820 , \29522_29821 , \29523_29822 , \29524_29823 , \29525_29824 , \29526_29825 , \29527_29826 , \29528_29827 , \29529_29828 , \29530_29829 , \29531_29830 );
or \U$20725 ( \29533_29832 , \29467_29766 , \29532_29831 );
_DC \g34f1/U$1 ( \29534 , \29533_29832 , \9298_9597 );
buf \U$20726 ( \29535_29834 , \29534 );
and \U$20727 ( \29536_29835 , \29402_29701 , \29535_29834 );
and \U$20728 ( \29537_29836 , \27400_27699 , \27533_27832 );
and \U$20729 ( \29538_29837 , \27533_27832 , \27808_28107 );
and \U$20730 ( \29539_29838 , \27400_27699 , \27808_28107 );
or \U$20731 ( \29540_29839 , \29537_29836 , \29538_29837 , \29539_29838 );
and \U$20732 ( \29541_29840 , \29535_29834 , \29540_29839 );
and \U$20733 ( \29542_29841 , \29402_29701 , \29540_29839 );
or \U$20734 ( \29543_29842 , \29536_29835 , \29541_29840 , \29542_29841 );
xor \U$20735 ( \29544_29843 , \29269_29568 , \29543_29842 );
buf g4400_GF_PartitionCandidate( \29545_29844_nG4400 , \29544_29843 );
xor \U$20736 ( \29546_29845 , \29402_29701 , \29535_29834 );
xor \U$20737 ( \29547_29846 , \29546_29845 , \29540_29839 );
buf g4403_GF_PartitionCandidate( \29548_29847_nG4403 , \29547_29846 );
nand \U$20738 ( \29549_29848 , \29548_29847_nG4403 , \27810_28109_nG4406 );
and \U$20739 ( \29550_29849 , \29545_29844_nG4400 , \29549_29848 );
xor \U$20740 ( \29551_29850 , \29548_29847_nG4403 , \27810_28109_nG4406 );
and \U$20745 ( \29552_29854 , \29551_29850 , \10392_10694_nG9c0e );
or \U$20746 ( \29553_29855 , 1'b0 , \29552_29854 );
xor \U$20747 ( \29554_29856 , \29550_29849 , \29553_29855 );
xor \U$20748 ( \29555_29857 , \29550_29849 , \29554_29856 );
buf \U$20749 ( \29556_29858 , \29555_29857 );
buf \U$20750 ( \29557_29859 , \29556_29858 );
xor \U$20751 ( \29558_29860 , \29002_29301 , \29557_29859 );
and \U$20752 ( \29559_29861 , \28450_28752 , \28989_29288 );
and \U$20753 ( \29560_29862 , \28450_28752 , \28995_29294 );
and \U$20754 ( \29561_29863 , \28989_29288 , \28995_29294 );
or \U$20755 ( \29562_29864 , \29559_29861 , \29560_29862 , \29561_29863 );
and \U$20756 ( \29563_29865 , \29558_29860 , \29562_29864 );
and \U$20757 ( \29564_29866 , \28884_29186 , \28889_29191 );
and \U$20758 ( \29565_29867 , \28884_29186 , \28987_29286 );
and \U$20759 ( \29566_29868 , \28889_29191 , \28987_29286 );
or \U$20760 ( \29567_29869 , \29564_29866 , \29565_29867 , \29566_29868 );
buf \U$20761 ( \29568_29870 , \29567_29869 );
and \U$20762 ( \29569_29871 , \28895_29197 , \28926_29228 );
and \U$20763 ( \29570_29872 , \28895_29197 , \28985_29284 );
and \U$20764 ( \29571_29873 , \28926_29228 , \28985_29284 );
or \U$20765 ( \29572_29874 , \29569_29871 , \29570_29872 , \29571_29873 );
buf \U$20766 ( \29573_29875 , \29572_29874 );
and \U$20767 ( \29574_29876 , \28900_29202 , \28917_29219 );
and \U$20768 ( \29575_29877 , \28900_29202 , \28924_29226 );
and \U$20769 ( \29576_29878 , \28917_29219 , \28924_29226 );
or \U$20770 ( \29577_29879 , \29574_29876 , \29575_29877 , \29576_29878 );
buf \U$20771 ( \29578_29880 , \29577_29879 );
and \U$20772 ( \29579_29881 , \14710_14631 , \22330_22629_nG9bd5 );
and \U$20773 ( \29580_29882 , \14329_14628 , \23394_23696_nG9bd2 );
or \U$20774 ( \29581_29883 , \29579_29881 , \29580_29882 );
xor \U$20775 ( \29582_29884 , \14328_14627 , \29581_29883 );
buf \U$20776 ( \29583_29885 , \29582_29884 );
buf \U$20778 ( \29584_29886 , \29583_29885 );
xor \U$20779 ( \29585_29887 , \29578_29880 , \29584_29886 );
and \U$20780 ( \29586_29888 , \13431_13370 , \23927_24226_nG9bcf );
and \U$20781 ( \29587_29889 , \13068_13367 , \24996_25298_nG9bcc );
or \U$20782 ( \29588_29890 , \29586_29888 , \29587_29889 );
xor \U$20783 ( \29589_29891 , \13067_13366 , \29588_29890 );
buf \U$20784 ( \29590_29892 , \29589_29891 );
buf \U$20786 ( \29591_29893 , \29590_29892 );
xor \U$20787 ( \29592_29894 , \29585_29887 , \29591_29893 );
buf \U$20788 ( \29593_29895 , \29592_29894 );
xor \U$20789 ( \29594_29896 , \29573_29875 , \29593_29895 );
and \U$20790 ( \29595_29897 , \28419_28721 , \28425_28727 );
and \U$20791 ( \29596_29898 , \28419_28721 , \28432_28734 );
and \U$20792 ( \29597_29899 , \28425_28727 , \28432_28734 );
or \U$20793 ( \29598_29900 , \29595_29897 , \29596_29898 , \29597_29899 );
buf \U$20794 ( \29599_29901 , \29598_29900 );
xor \U$20795 ( \29600_29902 , \29594_29896 , \29599_29901 );
buf \U$20796 ( \29601_29903 , \29600_29902 );
xor \U$20797 ( \29602_29904 , \29568_29870 , \29601_29903 );
and \U$20798 ( \29603_29905 , \28932_29234 , \28961_29260 );
and \U$20799 ( \29604_29906 , \28932_29234 , \28968_29267 );
and \U$20800 ( \29605_29907 , \28961_29260 , \28968_29267 );
or \U$20801 ( \29606_29908 , \29603_29905 , \29604_29906 , \29605_29907 );
buf \U$20802 ( \29607_29909 , \29606_29908 );
and \U$20803 ( \29608_29910 , \28902_29204 , \28908_29210 );
and \U$20804 ( \29609_29911 , \28902_29204 , \28915_29217 );
and \U$20805 ( \29610_29912 , \28908_29210 , \28915_29217 );
or \U$20806 ( \29611_29913 , \29608_29910 , \29609_29911 , \29610_29912 );
buf \U$20807 ( \29612_29914 , \29611_29913 );
and \U$20808 ( \29613_29915 , \28935_29237 , \28941_29243 );
buf \U$20809 ( \29614_29916 , \29613_29915 );
and \U$20810 ( \29615_29917 , \25044_24792 , \12502_12801_nG9bff );
and \U$20811 ( \29616_29918 , \24490_24789 , \13403_13705_nG9bfc );
or \U$20812 ( \29617_29919 , \29615_29917 , \29616_29918 );
xor \U$20813 ( \29618_29920 , \24489_24788 , \29617_29919 );
buf \U$20814 ( \29619_29921 , \29618_29920 );
buf \U$20816 ( \29620_29922 , \29619_29921 );
xor \U$20817 ( \29621_29923 , \29614_29916 , \29620_29922 );
and \U$20818 ( \29622_29924 , \23495_23201 , \13771_14070_nG9bf9 );
and \U$20819 ( \29623_29925 , \22899_23198 , \14682_14984_nG9bf6 );
or \U$20820 ( \29624_29926 , \29622_29924 , \29623_29925 );
xor \U$20821 ( \29625_29927 , \22898_23197 , \29624_29926 );
buf \U$20822 ( \29626_29928 , \29625_29927 );
buf \U$20824 ( \29627_29929 , \29626_29928 );
xor \U$20825 ( \29628_29930 , \29621_29923 , \29627_29929 );
buf \U$20826 ( \29629_29931 , \29628_29930 );
xor \U$20827 ( \29630_29932 , \29612_29914 , \29629_29931 );
and \U$20828 ( \29631_29933 , \20353_20155 , \16378_16680_nG9bed );
and \U$20829 ( \29632_29934 , \19853_20152 , \17363_17665_nG9bea );
or \U$20830 ( \29633_29935 , \29631_29933 , \29632_29934 );
xor \U$20831 ( \29634_29936 , \19852_20151 , \29633_29935 );
buf \U$20832 ( \29635_29937 , \29634_29936 );
buf \U$20834 ( \29636_29938 , \29635_29937 );
xor \U$20835 ( \29637_29939 , \29630_29932 , \29636_29938 );
buf \U$20836 ( \29638_29940 , \29637_29939 );
xor \U$20837 ( \29639_29941 , \29607_29909 , \29638_29940 );
and \U$20838 ( \29640_29942 , \17437_17297 , \19287_19586_nG9be1 );
and \U$20839 ( \29641_29943 , \16995_17294 , \20306_20608_nG9bde );
or \U$20840 ( \29642_29944 , \29640_29942 , \29641_29943 );
xor \U$20841 ( \29643_29945 , \16994_17293 , \29642_29944 );
buf \U$20842 ( \29644_29946 , \29643_29945 );
buf \U$20844 ( \29645_29947 , \29644_29946 );
xor \U$20845 ( \29646_29948 , \29639_29941 , \29645_29947 );
buf \U$20846 ( \29647_29949 , \29646_29948 );
and \U$20847 ( \29648_29950 , \12183_12157 , \25561_25860_nG9bc9 );
and \U$20848 ( \29649_29951 , \11855_12154 , \26585_26887_nG9bc6 );
or \U$20849 ( \29650_29952 , \29648_29950 , \29649_29951 );
xor \U$20850 ( \29651_29953 , \11854_12153 , \29650_29952 );
buf \U$20851 ( \29652_29954 , \29651_29953 );
buf \U$20853 ( \29653_29955 , \29652_29954 );
xor \U$20854 ( \29654_29956 , \29647_29949 , \29653_29955 );
and \U$20855 ( \29655_29957 , \10411_10707 , \28877_29179_nG9bbd );
and \U$20856 ( \29656_29958 , \28840_29142 , \28844_29146 );
and \U$20857 ( \29657_29959 , \28844_29146 , \28869_29171 );
and \U$20858 ( \29658_29960 , \28840_29142 , \28869_29171 );
or \U$20859 ( \29659_29961 , \29656_29958 , \29657_29959 , \29658_29960 );
and \U$20860 ( \29660_29962 , \28801_29103 , \28815_29117 );
and \U$20861 ( \29661_29963 , \28815_29117 , \28833_29135 );
and \U$20862 ( \29662_29964 , \28801_29103 , \28833_29135 );
or \U$20863 ( \29663_29965 , \29660_29962 , \29661_29963 , \29662_29964 );
and \U$20864 ( \29664_29966 , \28849_29151 , \28853_29155 );
and \U$20865 ( \29665_29967 , \28853_29155 , \28868_29170 );
and \U$20866 ( \29666_29968 , \28849_29151 , \28868_29170 );
or \U$20867 ( \29667_29969 , \29664_29966 , \29665_29967 , \29666_29968 );
xor \U$20868 ( \29668_29970 , \29663_29965 , \29667_29969 );
and \U$20869 ( \29669_29971 , \27011_27313 , \11275_11574 );
and \U$20870 ( \29670_29972 , \28232_28534 , \10976_11278 );
nor \U$20871 ( \29671_29973 , \29669_29971 , \29670_29972 );
xnor \U$20872 ( \29672_29974 , \29671_29973 , \11281_11580 );
and \U$20873 ( \29673_29975 , \23900_24199 , \13755_14054 );
and \U$20874 ( \29674_29976 , \24970_25272 , \13390_13692 );
nor \U$20875 ( \29675_29977 , \29673_29975 , \29674_29976 );
xnor \U$20876 ( \29676_29978 , \29675_29977 , \13736_14035 );
xor \U$20877 ( \29677_29979 , \29672_29974 , \29676_29978 );
and \U$20878 ( \29678_29980 , RIdec5db0_715, \9034_9333 );
and \U$20879 ( \29679_29981 , RIdec30b0_683, \9036_9335 );
and \U$20880 ( \29680_29982 , RIee201e8_4824, \9038_9337 );
and \U$20881 ( \29681_29983 , RIdec03b0_651, \9040_9339 );
and \U$20882 ( \29682_29984 , RIfcaf538_7017, \9042_9341 );
and \U$20883 ( \29683_29985 , RIdebd6b0_619, \9044_9343 );
and \U$20884 ( \29684_29986 , RIdeba9b0_587, \9046_9345 );
and \U$20885 ( \29685_29987 , RIdeb7cb0_555, \9048_9347 );
and \U$20886 ( \29686_29988 , RIfc40fe8_5765, \9050_9349 );
and \U$20887 ( \29687_29989 , RIdeb22b0_491, \9052_9351 );
and \U$20888 ( \29688_29990 , RIfcd08c8_7395, \9054_9353 );
and \U$20889 ( \29689_29991 , RIdeaf5b0_459, \9056_9355 );
and \U$20890 ( \29690_29992 , RIee1dd58_4798, \9058_9357 );
and \U$20891 ( \29691_29993 , RIdeabb18_427, \9060_9359 );
and \U$20892 ( \29692_29994 , RIdea5218_395, \9062_9361 );
and \U$20893 ( \29693_29995 , RIde9e918_363, \9064_9363 );
and \U$20894 ( \29694_29996 , RIee1d218_4790, \9066_9365 );
and \U$20895 ( \29695_29997 , RIfcedd10_7728, \9068_9367 );
and \U$20896 ( \29696_29998 , RIfce62b8_7641, \9070_9369 );
and \U$20897 ( \29697_29999 , RIfcc92a8_7311, \9072_9371 );
and \U$20898 ( \29698_30000 , RIde91da8_301, \9074_9373 );
and \U$20899 ( \29699_30001 , RIde8e928_285, \9076_9375 );
and \U$20900 ( \29700_30002 , RIde8a788_265, \9078_9377 );
and \U$20901 ( \29701_30003 , RIde865e8_245, \9080_9379 );
and \U$20902 ( \29702_30004 , RIde82448_225, \9082_9381 );
and \U$20903 ( \29703_30005 , RIfea1448_8179, \9084_9383 );
and \U$20904 ( \29704_30006 , RIfc750e0_6354, \9086_9385 );
and \U$20905 ( \29705_30007 , RIfcc19b8_7225, \9088_9387 );
and \U$20906 ( \29706_30008 , RIfced8d8_7725, \9090_9389 );
and \U$20907 ( \29707_30009 , RIfec5eb0_8372, \9092_9391 );
and \U$20908 ( \29708_30010 , RIe169fc8_2583, \9094_9393 );
and \U$20909 ( \29709_30011 , RIe168678_2565, \9096_9395 );
and \U$20910 ( \29710_30012 , RIe165db0_2536, \9098_9397 );
and \U$20911 ( \29711_30013 , RIe1630b0_2504, \9100_9399 );
and \U$20912 ( \29712_30014 , RIfccfc20_7386, \9102_9401 );
and \U$20913 ( \29713_30015 , RIe1603b0_2472, \9104_9403 );
and \U$20914 ( \29714_30016 , RIee365b0_5077, \9106_9405 );
and \U$20915 ( \29715_30017 , RIe15d6b0_2440, \9108_9407 );
and \U$20916 ( \29716_30018 , RIe157cb0_2376, \9110_9409 );
and \U$20917 ( \29717_30019 , RIe154fb0_2344, \9112_9411 );
and \U$20918 ( \29718_30020 , RIfea1718_8181, \9114_9413 );
and \U$20919 ( \29719_30021 , RIe1522b0_2312, \9116_9415 );
and \U$20920 ( \29720_30022 , RIee35200_5063, \9118_9417 );
and \U$20921 ( \29721_30023 , RIe14f5b0_2280, \9120_9419 );
and \U$20922 ( \29722_30024 , RIfcb0348_7027, \9122_9421 );
and \U$20923 ( \29723_30025 , RIe14c8b0_2248, \9124_9423 );
and \U$20924 ( \29724_30026 , RIe149bb0_2216, \9126_9425 );
and \U$20925 ( \29725_30027 , RIe146eb0_2184, \9128_9427 );
and \U$20926 ( \29726_30028 , RIfc73790_6336, \9130_9429 );
and \U$20927 ( \29727_30029 , RIfcdf238_7561, \9132_9431 );
and \U$20928 ( \29728_30030 , RIee32500_5031, \9134_9433 );
and \U$20929 ( \29729_30031 , RIfc94f58_6717, \9136_9435 );
and \U$20930 ( \29730_30032 , RIe141780_2122, \9138_9437 );
and \U$20931 ( \29731_30033 , RIe13f2f0_2096, \9140_9439 );
and \U$20932 ( \29732_30034 , RIfec5be0_8370, \9142_9441 );
and \U$20933 ( \29733_30035 , RIdf3ad68_2046, \9144_9443 );
and \U$20934 ( \29734_30036 , RIfea15b0_8180, \9146_9445 );
and \U$20935 ( \29735_30037 , RIfc5fb28_6111, \9148_9447 );
and \U$20936 ( \29736_30038 , RIfcae728_7007, \9150_9449 );
and \U$20937 ( \29737_30039 , RIfc74438_6345, \9152_9451 );
and \U$20938 ( \29738_30040 , RIdf36178_1992, \9154_9453 );
and \U$20939 ( \29739_30041 , RIdf33b80_1965, \9156_9455 );
and \U$20940 ( \29740_30042 , RIdf319c0_1941, \9158_9457 );
and \U$20941 ( \29741_30043 , RIdf2fad0_1919, \9160_9459 );
or \U$20942 ( \29742_30044 , \29678_29980 , \29679_29981 , \29680_29982 , \29681_29983 , \29682_29984 , \29683_29985 , \29684_29986 , \29685_29987 , \29686_29988 , \29687_29989 , \29688_29990 , \29689_29991 , \29690_29992 , \29691_29993 , \29692_29994 , \29693_29995 , \29694_29996 , \29695_29997 , \29696_29998 , \29697_29999 , \29698_30000 , \29699_30001 , \29700_30002 , \29701_30003 , \29702_30004 , \29703_30005 , \29704_30006 , \29705_30007 , \29706_30008 , \29707_30009 , \29708_30010 , \29709_30011 , \29710_30012 , \29711_30013 , \29712_30014 , \29713_30015 , \29714_30016 , \29715_30017 , \29716_30018 , \29717_30019 , \29718_30020 , \29719_30021 , \29720_30022 , \29721_30023 , \29722_30024 , \29723_30025 , \29724_30026 , \29725_30027 , \29726_30028 , \29727_30029 , \29728_30030 , \29729_30031 , \29730_30032 , \29731_30033 , \29732_30034 , \29733_30035 , \29734_30036 , \29735_30037 , \29736_30038 , \29737_30039 , \29738_30040 , \29739_30041 , \29740_30042 , \29741_30043 );
and \U$20943 ( \29743_30045 , RIee2c290_4961, \9163_9462 );
and \U$20944 ( \29744_30046 , RIee2a940_4943, \9165_9464 );
and \U$20945 ( \29745_30047 , RIfc70658_6301, \9167_9466 );
and \U$20946 ( \29746_30048 , RIfc704f0_6300, \9169_9468 );
and \U$20947 ( \29747_30049 , RIdf2aaa8_1862, \9171_9470 );
and \U$20948 ( \29748_30050 , RIdf288e8_1838, \9173_9472 );
and \U$20949 ( \29749_30051 , RIdf269f8_1816, \9175_9474 );
and \U$20950 ( \29750_30052 , RIdf24f40_1797, \9177_9476 );
and \U$20951 ( \29751_30053 , RIfc64b50_6168, \9179_9478 );
and \U$20952 ( \29752_30054 , RIfccaa90_7328, \9181_9480 );
and \U$20953 ( \29753_30055 , RIdf231b8_1776, \9183_9482 );
and \U$20954 ( \29754_30056 , RIfcad4e0_6994, \9185_9484 );
and \U$20955 ( \29755_30057 , RIdf21ca0_1761, \9187_9486 );
and \U$20956 ( \29756_30058 , RIfeaad90_8260, \9189_9488 );
and \U$20957 ( \29757_30059 , RIdf1b490_1687, \9191_9490 );
and \U$20958 ( \29758_30060 , RIdf19b40_1669, \9193_9492 );
and \U$20959 ( \29759_30061 , RIdf17980_1645, \9195_9494 );
and \U$20960 ( \29760_30062 , RIdf14c80_1613, \9197_9496 );
and \U$20961 ( \29761_30063 , RIdf11f80_1581, \9199_9498 );
and \U$20962 ( \29762_30064 , RIdf0f280_1549, \9201_9500 );
and \U$20963 ( \29763_30065 , RIdf0c580_1517, \9203_9502 );
and \U$20964 ( \29764_30066 , RIdf09880_1485, \9205_9504 );
and \U$20965 ( \29765_30067 , RIdf06b80_1453, \9207_9506 );
and \U$20966 ( \29766_30068 , RIdf03e80_1421, \9209_9508 );
and \U$20967 ( \29767_30069 , RIdefe480_1357, \9211_9510 );
and \U$20968 ( \29768_30070 , RIdefb780_1325, \9213_9512 );
and \U$20969 ( \29769_30071 , RIdef8a80_1293, \9215_9514 );
and \U$20970 ( \29770_30072 , RIdef5d80_1261, \9217_9516 );
and \U$20971 ( \29771_30073 , RIdef3080_1229, \9219_9518 );
and \U$20972 ( \29772_30074 , RIdef0380_1197, \9221_9520 );
and \U$20973 ( \29773_30075 , RIdeed680_1165, \9223_9522 );
and \U$20974 ( \29774_30076 , RIdeea980_1133, \9225_9524 );
and \U$20975 ( \29775_30077 , RIfc595e8_6039, \9227_9526 );
and \U$20976 ( \29776_30078 , RIfcac568_6983, \9229_9528 );
and \U$20977 ( \29777_30079 , RIfcccf20_7354, \9231_9530 );
and \U$20978 ( \29778_30080 , RIfccd358_7357, \9233_9532 );
and \U$20979 ( \29779_30081 , RIdee5250_1071, \9235_9534 );
and \U$20980 ( \29780_30082 , RIfea7f28_8227, \9237_9536 );
and \U$20981 ( \29781_30083 , RIdee11a0_1025, \9239_9538 );
and \U$20982 ( \29782_30084 , RIfea12e0_8178, \9241_9540 );
and \U$20983 ( \29783_30085 , RIfc679b8_6201, \9243_9542 );
and \U$20984 ( \29784_30086 , RIee22510_4849, \9245_9544 );
and \U$20985 ( \29785_30087 , RIfc6dd90_6272, \9247_9546 );
and \U$20986 ( \29786_30088 , RIfc6cb48_6259, \9249_9548 );
and \U$20987 ( \29787_30089 , RIdeda120_945, \9251_9550 );
and \U$20988 ( \29788_30090 , RIded7b28_918, \9253_9552 );
and \U$20989 ( \29789_30091 , RIded5c38_896, \9255_9554 );
and \U$20990 ( \29790_30092 , RIfec5d48_8371, \9257_9556 );
and \U$20991 ( \29791_30093 , RIded11b0_843, \9259_9558 );
and \U$20992 ( \29792_30094 , RIdece4b0_811, \9261_9560 );
and \U$20993 ( \29793_30095 , RIdecb7b0_779, \9263_9562 );
and \U$20994 ( \29794_30096 , RIdec8ab0_747, \9265_9564 );
and \U$20995 ( \29795_30097 , RIdeb4fb0_523, \9267_9566 );
and \U$20996 ( \29796_30098 , RIde98018_331, \9269_9568 );
and \U$20997 ( \29797_30099 , RIe16ebb8_2637, \9271_9570 );
and \U$20998 ( \29798_30100 , RIe15a9b0_2408, \9273_9572 );
and \U$20999 ( \29799_30101 , RIe1441b0_2152, \9275_9574 );
and \U$21000 ( \29800_30102 , RIdf38ba8_2022, \9277_9576 );
and \U$21001 ( \29801_30103 , RIdf2d208_1890, \9279_9578 );
and \U$21002 ( \29802_30104 , RIdf1da88_1714, \9281_9580 );
and \U$21003 ( \29803_30105 , RIdf01180_1389, \9283_9582 );
and \U$21004 ( \29804_30106 , RIdee7c80_1101, \9285_9584 );
and \U$21005 ( \29805_30107 , RIdedc9e8_974, \9287_9586 );
and \U$21006 ( \29806_30108 , RIde7df60_204, \9289_9588 );
or \U$21007 ( \29807_30109 , \29743_30045 , \29744_30046 , \29745_30047 , \29746_30048 , \29747_30049 , \29748_30050 , \29749_30051 , \29750_30052 , \29751_30053 , \29752_30054 , \29753_30055 , \29754_30056 , \29755_30057 , \29756_30058 , \29757_30059 , \29758_30060 , \29759_30061 , \29760_30062 , \29761_30063 , \29762_30064 , \29763_30065 , \29764_30066 , \29765_30067 , \29766_30068 , \29767_30069 , \29768_30070 , \29769_30071 , \29770_30072 , \29771_30073 , \29772_30074 , \29773_30075 , \29774_30076 , \29775_30077 , \29776_30078 , \29777_30079 , \29778_30080 , \29779_30081 , \29780_30082 , \29781_30083 , \29782_30084 , \29783_30085 , \29784_30086 , \29785_30087 , \29786_30088 , \29787_30089 , \29788_30090 , \29789_30091 , \29790_30092 , \29791_30093 , \29792_30094 , \29793_30095 , \29794_30096 , \29795_30097 , \29796_30098 , \29797_30099 , \29798_30100 , \29799_30101 , \29800_30102 , \29801_30103 , \29802_30104 , \29803_30105 , \29804_30106 , \29805_30107 , \29806_30108 );
or \U$21008 ( \29808_30110 , \29742_30044 , \29807_30109 );
_DC \g61d6/U$1 ( \29809 , \29808_30110 , \9298_9597 );
and \U$21009 ( \29810_30112 , RIe19e048_3175, \8760_9059 );
and \U$21010 ( \29811_30113 , RIe19b348_3143, \8762_9061 );
and \U$21011 ( \29812_30114 , RIfcc3ce0_7250, \8764_9063 );
and \U$21012 ( \29813_30115 , RIe198648_3111, \8766_9065 );
and \U$21013 ( \29814_30116 , RIfc7efc8_6467, \8768_9067 );
and \U$21014 ( \29815_30117 , RIe195948_3079, \8770_9069 );
and \U$21015 ( \29816_30118 , RIe192c48_3047, \8772_9071 );
and \U$21016 ( \29817_30119 , RIe18ff48_3015, \8774_9073 );
and \U$21017 ( \29818_30120 , RIe18a548_2951, \8776_9075 );
and \U$21018 ( \29819_30121 , RIe187848_2919, \8778_9077 );
and \U$21019 ( \29820_30122 , RIfc46790_5824, \8780_9079 );
and \U$21020 ( \29821_30123 , RIe184b48_2887, \8782_9081 );
and \U$21021 ( \29822_30124 , RIfc98d38_6761, \8784_9083 );
and \U$21022 ( \29823_30125 , RIe181e48_2855, \8786_9085 );
and \U$21023 ( \29824_30126 , RIe17f148_2823, \8788_9087 );
and \U$21024 ( \29825_30127 , RIe17c448_2791, \8790_9089 );
and \U$21025 ( \29826_30128 , RIfcb5d48_7091, \8792_9091 );
and \U$21026 ( \29827_30129 , RIfc995a8_6767, \8794_9093 );
and \U$21027 ( \29828_30130 , RIfc9a3b8_6777, \8796_9095 );
and \U$21028 ( \29829_30131 , RIe1761d8_2721, \8798_9097 );
and \U$21029 ( \29830_30132 , RIfc54188_5979, \8800_9099 );
and \U$21030 ( \29831_30133 , RIfcd2bf0_7420, \8802_9101 );
and \U$21031 ( \29832_30134 , RIfc8b778_6609, \8804_9103 );
and \U$21032 ( \29833_30135 , RIfc7dee8_6455, \8806_9105 );
and \U$21033 ( \29834_30136 , RIee3c550_5145, \8808_9107 );
and \U$21034 ( \29835_30137 , RIfc8c420_6618, \8810_9109 );
and \U$21035 ( \29836_30138 , RIee3a0c0_5119, \8812_9111 );
and \U$21036 ( \29837_30139 , RIfeaba38_8269, \8814_9113 );
and \U$21037 ( \29838_30140 , RIfc46628_5823, \8816_9115 );
and \U$21038 ( \29839_30141 , RIfcbc288_7163, \8818_9117 );
and \U$21039 ( \29840_30142 , RIf16e710_5716, \8820_9119 );
and \U$21040 ( \29841_30143 , RIfc8fdc8_6659, \8822_9121 );
and \U$21041 ( \29842_30144 , RIfc48c20_5850, \8824_9123 );
and \U$21042 ( \29843_30145 , RIe2243a0_4702, \8826_9125 );
and \U$21043 ( \29844_30146 , RIfca0358_6845, \8828_9127 );
and \U$21044 ( \29845_30147 , RIe2216a0_4670, \8830_9129 );
and \U$21045 ( \29846_30148 , RIfc9a688_6779, \8832_9131 );
and \U$21046 ( \29847_30149 , RIe21e9a0_4638, \8834_9133 );
and \U$21047 ( \29848_30150 , RIe218fa0_4574, \8836_9135 );
and \U$21048 ( \29849_30151 , RIe2162a0_4542, \8838_9137 );
and \U$21049 ( \29850_30152 , RIfc456b0_5812, \8840_9139 );
and \U$21050 ( \29851_30153 , RIe2135a0_4510, \8842_9141 );
and \U$21051 ( \29852_30154 , RIf169418_5657, \8844_9143 );
and \U$21052 ( \29853_30155 , RIe2108a0_4478, \8846_9145 );
and \U$21053 ( \29854_30156 , RIfc8bfe8_6615, \8848_9147 );
and \U$21054 ( \29855_30157 , RIe20dba0_4446, \8850_9149 );
and \U$21055 ( \29856_30158 , RIe20aea0_4414, \8852_9151 );
and \U$21056 ( \29857_30159 , RIe2081a0_4382, \8854_9153 );
and \U$21057 ( \29858_30160 , RIfc8c9c0_6622, \8856_9155 );
and \U$21058 ( \29859_30161 , RIfc7f568_6471, \8858_9157 );
and \U$21059 ( \29860_30162 , RIe202d40_4322, \8860_9159 );
and \U$21060 ( \29861_30163 , RIe201120_4302, \8862_9161 );
and \U$21061 ( \29862_30164 , RIfce2910_7600, \8864_9163 );
and \U$21062 ( \29863_30165 , RIfc487e8_5847, \8866_9165 );
and \U$21063 ( \29864_30166 , RIfc46d30_5828, \8868_9167 );
and \U$21064 ( \29865_30167 , RIfc992d8_6765, \8870_9169 );
and \U$21065 ( \29866_30168 , RIfca2680_6870, \8872_9171 );
and \U$21066 ( \29867_30169 , RIfc44a08_5803, \8874_9173 );
and \U$21067 ( \29868_30170 , RIe1fd1d8_4257, \8876_9175 );
and \U$21068 ( \29869_30171 , RIe1fbf90_4244, \8878_9177 );
and \U$21069 ( \29870_30172 , RIfc580d0_6024, \8880_9179 );
and \U$21070 ( \29871_30173 , RIfcbdbd8_7181, \8882_9181 );
and \U$21071 ( \29872_30174 , RIfc8dd70_6636, \8884_9183 );
and \U$21072 ( \29873_30175 , RIfce01b0_7572, \8886_9185 );
or \U$21073 ( \29874_30176 , \29810_30112 , \29811_30113 , \29812_30114 , \29813_30115 , \29814_30116 , \29815_30117 , \29816_30118 , \29817_30119 , \29818_30120 , \29819_30121 , \29820_30122 , \29821_30123 , \29822_30124 , \29823_30125 , \29824_30126 , \29825_30127 , \29826_30128 , \29827_30129 , \29828_30130 , \29829_30131 , \29830_30132 , \29831_30133 , \29832_30134 , \29833_30135 , \29834_30136 , \29835_30137 , \29836_30138 , \29837_30139 , \29838_30140 , \29839_30141 , \29840_30142 , \29841_30143 , \29842_30144 , \29843_30145 , \29844_30146 , \29845_30147 , \29846_30148 , \29847_30149 , \29848_30150 , \29849_30151 , \29850_30152 , \29851_30153 , \29852_30154 , \29853_30155 , \29854_30156 , \29855_30157 , \29856_30158 , \29857_30159 , \29858_30160 , \29859_30161 , \29860_30162 , \29861_30163 , \29862_30164 , \29863_30165 , \29864_30166 , \29865_30167 , \29866_30168 , \29867_30169 , \29868_30170 , \29869_30171 , \29870_30172 , \29871_30173 , \29872_30174 , \29873_30175 );
and \U$21074 ( \29875_30177 , RIfc7bbc0_6430, \8889_9188 );
and \U$21075 ( \29876_30178 , RIfc90368_6663, \8891_9190 );
and \U$21076 ( \29877_30179 , RIfc7b8f0_6428, \8893_9192 );
and \U$21077 ( \29878_30180 , RIe1fa910_4228, \8895_9194 );
and \U$21078 ( \29879_30181 , RIfcd8b90_7488, \8897_9196 );
and \U$21079 ( \29880_30182 , RIfc43ec8_5795, \8899_9198 );
and \U$21080 ( \29881_30183 , RIfc7b788_6427, \8901_9200 );
and \U$21081 ( \29882_30184 , RIe1f5e88_4175, \8903_9202 );
and \U$21082 ( \29883_30185 , RIfc7b350_6424, \8905_9204 );
and \U$21083 ( \29884_30186 , RIfc90d40_6670, \8907_9206 );
and \U$21084 ( \29885_30187 , RIfca3490_6880, \8909_9208 );
and \U$21085 ( \29886_30188 , RIe1f3b60_4150, \8911_9210 );
and \U$21086 ( \29887_30189 , RIfc91010_6672, \8913_9212 );
and \U$21087 ( \29888_30190 , RIfcdb728_7519, \8915_9214 );
and \U$21088 ( \29889_30191 , RIfcd8758_7485, \8917_9216 );
and \U$21089 ( \29890_30192 , RIe1ee868_4091, \8919_9218 );
and \U$21090 ( \29891_30193 , RIe1ec108_4063, \8921_9220 );
and \U$21091 ( \29892_30194 , RIe1e9408_4031, \8923_9222 );
and \U$21092 ( \29893_30195 , RIe1e6708_3999, \8925_9224 );
and \U$21093 ( \29894_30196 , RIe1e3a08_3967, \8927_9226 );
and \U$21094 ( \29895_30197 , RIe1e0d08_3935, \8929_9228 );
and \U$21095 ( \29896_30198 , RIe1de008_3903, \8931_9230 );
and \U$21096 ( \29897_30199 , RIe1db308_3871, \8933_9232 );
and \U$21097 ( \29898_30200 , RIe1d8608_3839, \8935_9234 );
and \U$21098 ( \29899_30201 , RIe1d2c08_3775, \8937_9236 );
and \U$21099 ( \29900_30202 , RIe1cff08_3743, \8939_9238 );
and \U$21100 ( \29901_30203 , RIe1cd208_3711, \8941_9240 );
and \U$21101 ( \29902_30204 , RIe1ca508_3679, \8943_9242 );
and \U$21102 ( \29903_30205 , RIe1c7808_3647, \8945_9244 );
and \U$21103 ( \29904_30206 , RIe1c4b08_3615, \8947_9246 );
and \U$21104 ( \29905_30207 , RIe1c1e08_3583, \8949_9248 );
and \U$21105 ( \29906_30208 , RIe1bf108_3551, \8951_9250 );
and \U$21106 ( \29907_30209 , RIf14cf48_5335, \8953_9252 );
and \U$21107 ( \29908_30210 , RIfc78d58_6397, \8955_9254 );
and \U$21108 ( \29909_30211 , RIe1b9b40_3490, \8957_9256 );
and \U$21109 ( \29910_30212 , RIfec5910_8368, \8959_9258 );
and \U$21110 ( \29911_30213 , RIfc78a88_6395, \8961_9260 );
and \U$21111 ( \29912_30214 , RIfcd51e8_7447, \8963_9262 );
and \U$21112 ( \29913_30215 , RIe1b57c0_3442, \8965_9264 );
and \U$21113 ( \29914_30216 , RIfea1010_8176, \8967_9266 );
and \U$21114 ( \29915_30217 , RIf1492d0_5292, \8969_9268 );
and \U$21115 ( \29916_30218 , RIfec5a78_8369, \8971_9270 );
and \U$21116 ( \29917_30219 , RIe1b2c28_3411, \8973_9272 );
and \U$21117 ( \29918_30220 , RIe1b12d8_3393, \8975_9274 );
and \U$21118 ( \29919_30221 , RIfec5640_8366, \8977_9276 );
and \U$21119 ( \29920_30222 , RIf146a08_5263, \8979_9278 );
and \U$21120 ( \29921_30223 , RIfec57a8_8367, \8981_9280 );
and \U$21121 ( \29922_30224 , RIfea1178_8177, \8983_9282 );
and \U$21122 ( \29923_30225 , RIe1a9448_3303, \8985_9284 );
and \U$21123 ( \29924_30226 , RIe1a6748_3271, \8987_9286 );
and \U$21124 ( \29925_30227 , RIe1a3a48_3239, \8989_9288 );
and \U$21125 ( \29926_30228 , RIe1a0d48_3207, \8991_9290 );
and \U$21126 ( \29927_30229 , RIe18d248_2983, \8993_9292 );
and \U$21127 ( \29928_30230 , RIe179748_2759, \8995_9294 );
and \U$21128 ( \29929_30231 , RIe2270a0_4734, \8997_9296 );
and \U$21129 ( \29930_30232 , RIe21bca0_4606, \8999_9298 );
and \U$21130 ( \29931_30233 , RIe2054a0_4350, \9001_9300 );
and \U$21131 ( \29932_30234 , RIe1ff500_4282, \9003_9302 );
and \U$21132 ( \29933_30235 , RIe1f88b8_4205, \9005_9304 );
and \U$21133 ( \29934_30236 , RIe1f1400_4122, \9007_9306 );
and \U$21134 ( \29935_30237 , RIe1d5908_3807, \9009_9308 );
and \U$21135 ( \29936_30238 , RIe1bc408_3519, \9011_9310 );
and \U$21136 ( \29937_30239 , RIe1af280_3370, \9013_9312 );
and \U$21137 ( \29938_30240 , RIe1718b8_2669, \9015_9314 );
or \U$21138 ( \29939_30241 , \29875_30177 , \29876_30178 , \29877_30179 , \29878_30180 , \29879_30181 , \29880_30182 , \29881_30183 , \29882_30184 , \29883_30185 , \29884_30186 , \29885_30187 , \29886_30188 , \29887_30189 , \29888_30190 , \29889_30191 , \29890_30192 , \29891_30193 , \29892_30194 , \29893_30195 , \29894_30196 , \29895_30197 , \29896_30198 , \29897_30199 , \29898_30200 , \29899_30201 , \29900_30202 , \29901_30203 , \29902_30204 , \29903_30205 , \29904_30206 , \29905_30207 , \29906_30208 , \29907_30209 , \29908_30210 , \29909_30211 , \29910_30212 , \29911_30213 , \29912_30214 , \29913_30215 , \29914_30216 , \29915_30217 , \29916_30218 , \29917_30219 , \29918_30220 , \29919_30221 , \29920_30222 , \29921_30223 , \29922_30224 , \29923_30225 , \29924_30226 , \29925_30227 , \29926_30228 , \29927_30229 , \29928_30230 , \29929_30231 , \29930_30232 , \29931_30233 , \29932_30234 , \29933_30235 , \29934_30236 , \29935_30237 , \29936_30238 , \29937_30239 , \29938_30240 );
or \U$21139 ( \29940_30242 , \29874_30176 , \29939_30241 );
_DC \g625a/U$1 ( \29941 , \29940_30242 , \9024_9323 );
xor g625b_GF_PartitionCandidate( \29942_30244_nG625b , \29809 , \29941 );
buf \U$21140 ( \29943_30245 , \29942_30244_nG625b );
xor \U$21141 ( \29944_30246 , \29943_30245 , \28765_29067 );
and \U$21142 ( \29945_30247 , \10385_10687 , \29944_30246 );
xor \U$21143 ( \29946_30248 , \29677_29979 , \29945_30247 );
and \U$21144 ( \29947_30249 , \25516_25815 , \12491_12790 );
and \U$21145 ( \29948_30250 , \26527_26829 , \12159_12461 );
nor \U$21146 ( \29949_30251 , \29947_30249 , \29948_30250 );
xnor \U$21147 ( \29950_30252 , \29949_30251 , \12481_12780 );
and \U$21148 ( \29951_30253 , \19259_19558 , \17791_18090 );
and \U$21149 ( \29952_30254 , \20242_20544 , \17353_17655 );
nor \U$21150 ( \29953_30255 , \29951_30253 , \29952_30254 );
xnor \U$21151 ( \29954_30256 , \29953_30255 , \17747_18046 );
xor \U$21152 ( \29955_30257 , \29950_30252 , \29954_30256 );
and \U$21153 ( \29956_30258 , \10686_10988 , \28768_29070 );
and \U$21154 ( \29957_30259 , \10968_11270 , \28224_28526 );
nor \U$21155 ( \29958_30260 , \29956_30258 , \29957_30259 );
xnor \U$21156 ( \29959_30261 , \29958_30260 , \28774_29076 );
xor \U$21157 ( \29960_30262 , \29955_30257 , \29959_30261 );
xor \U$21158 ( \29961_30263 , \29946_30248 , \29960_30262 );
and \U$21159 ( \29962_30264 , \28782_29084 , \10681_10983 );
_DC \g65cb/U$1 ( \29963 , \29808_30110 , \9298_9597 );
_DC \g65cc/U$1 ( \29964 , \29940_30242 , \9024_9323 );
and g65cd_GF_PartitionCandidate( \29965_30267_nG65cd , \29963 , \29964 );
buf \U$21160 ( \29966_30268 , \29965_30267_nG65cd );
and \U$21161 ( \29967_30269 , \29966_30268 , \10389_10691 );
nor \U$21162 ( \29968_30270 , \29962_30264 , \29967_30269 );
xnor \U$21163 ( \29969_30271 , \29968_30270 , \10678_10980 );
and \U$21164 ( \29970_30272 , \15022_15321 , \22243_22542 );
and \U$21165 ( \29971_30273 , \15965_16267 , \21801_22103 );
nor \U$21166 ( \29972_30274 , \29970_30272 , \29971_30273 );
xnor \U$21167 ( \29973_30275 , \29972_30274 , \22249_22548 );
xor \U$21168 ( \29974_30276 , \29969_30271 , \29973_30275 );
and \U$21169 ( \29975_30277 , \13725_14024 , \23839_24138 );
and \U$21170 ( \29976_30278 , \14648_14950 , \23328_23630 );
nor \U$21171 ( \29977_30279 , \29975_30277 , \29976_30278 );
xnor \U$21172 ( \29978_30280 , \29977_30279 , \23845_24144 );
xor \U$21173 ( \29979_30281 , \29974_30276 , \29978_30280 );
xor \U$21174 ( \29980_30282 , \29961_30263 , \29979_30281 );
xor \U$21175 ( \29981_30283 , \29668_29970 , \29980_30282 );
xor \U$21176 ( \29982_30284 , \29659_29961 , \29981_30283 );
and \U$21177 ( \29983_30285 , \28476_28778 , \28796_29098 );
and \U$21178 ( \29984_30286 , \28796_29098 , \28834_29136 );
and \U$21179 ( \29985_30287 , \28476_28778 , \28834_29136 );
or \U$21180 ( \29986_30288 , \29983_30285 , \29984_30286 , \29985_30287 );
and \U$21181 ( \29987_30289 , \28858_29160 , \28862_29164 );
and \U$21182 ( \29988_30290 , \28862_29164 , \28867_29169 );
and \U$21183 ( \29989_30291 , \28858_29160 , \28867_29169 );
or \U$21184 ( \29990_30292 , \29987_30289 , \29988_30290 , \29989_30291 );
and \U$21185 ( \29991_30293 , \28823_29125 , \28827_29129 );
and \U$21186 ( \29992_30294 , \28827_29129 , \28832_29134 );
and \U$21187 ( \29993_30295 , \28823_29125 , \28832_29134 );
or \U$21188 ( \29994_30296 , \29991_30293 , \29992_30294 , \29993_30295 );
xor \U$21189 ( \29995_30297 , \29990_30292 , \29994_30296 );
and \U$21190 ( \29996_30298 , \20734_21033 , \16333_16635 );
and \U$21191 ( \29997_30299 , \21788_22090 , \15999_16301 );
nor \U$21192 ( \29998_30300 , \29996_30298 , \29997_30299 );
xnor \U$21193 ( \29999_30301 , \29998_30300 , \16323_16625 );
and \U$21194 ( \30000_30302 , \12470_12769 , \25527_25826 );
and \U$21195 ( \30001_30303 , \13377_13679 , \24962_25264 );
nor \U$21196 ( \30002_30304 , \30000_30302 , \30001_30303 );
xnor \U$21197 ( \30003_30305 , \30002_30304 , \25474_25773 );
xor \U$21198 ( \30004_30306 , \29999_30301 , \30003_30305 );
and \U$21199 ( \30005_30307 , \11287_11586 , \27095_27397 );
and \U$21200 ( \30006_30308 , \12146_12448 , \26505_26807 );
nor \U$21201 ( \30007_30309 , \30005_30307 , \30006_30308 );
xnor \U$21202 ( \30008_30310 , \30007_30309 , \26993_27295 );
xor \U$21203 ( \30009_30311 , \30004_30306 , \30008_30310 );
xor \U$21204 ( \30010_30312 , \29995_30297 , \30009_30311 );
xor \U$21205 ( \30011_30313 , \29986_30288 , \30010_30312 );
and \U$21206 ( \30012_30314 , \28490_28792 , \28776_29078 );
and \U$21207 ( \30013_30315 , \28776_29078 , \28795_29097 );
and \U$21208 ( \30014_30316 , \28490_28792 , \28795_29097 );
or \U$21209 ( \30015_30317 , \30012_30314 , \30013_30315 , \30014_30316 );
and \U$21210 ( \30016_30318 , \28480_28782 , \28484_28786 );
and \U$21211 ( \30017_30319 , \28484_28786 , \28489_28791 );
and \U$21212 ( \30018_30320 , \28480_28782 , \28489_28791 );
or \U$21213 ( \30019_30321 , \30016_30318 , \30017_30319 , \30018_30320 );
and \U$21214 ( \30020_30322 , \28805_29107 , \28809_29111 );
and \U$21215 ( \30021_30323 , \28809_29111 , \28814_29116 );
and \U$21216 ( \30022_30324 , \28805_29107 , \28814_29116 );
or \U$21217 ( \30023_30325 , \30020_30322 , \30021_30323 , \30022_30324 );
xor \U$21218 ( \30024_30326 , \30019_30321 , \30023_30325 );
and \U$21219 ( \30025_30327 , \28820_29122 , \28822_29124 );
xor \U$21220 ( \30026_30328 , \30024_30326 , \30025_30327 );
xor \U$21221 ( \30027_30329 , \30015_30317 , \30026_30328 );
and \U$21222 ( \30028_30330 , \28494_28796 , \28498_28800 );
and \U$21223 ( \30029_30331 , \28498_28800 , \28775_29077 );
and \U$21224 ( \30030_30332 , \28494_28796 , \28775_29077 );
or \U$21225 ( \30031_30333 , \30028_30330 , \30029_30331 , \30030_30332 );
and \U$21226 ( \30032_30334 , \28785_29087 , \28789_29091 );
and \U$21227 ( \30033_30335 , \28789_29091 , \28794_29096 );
and \U$21228 ( \30034_30336 , \28785_29087 , \28794_29096 );
or \U$21229 ( \30035_30337 , \30032_30334 , \30033_30335 , \30034_30336 );
xor \U$21230 ( \30036_30338 , \30031_30333 , \30035_30337 );
and \U$21231 ( \30037_30339 , \22257_22556 , \15037_15336 );
and \U$21232 ( \30038_30340 , \23315_23617 , \14661_14963 );
nor \U$21233 ( \30039_30341 , \30037_30339 , \30038_30340 );
xnor \U$21234 ( \30040_30342 , \30039_30341 , \15043_15342 );
and \U$21235 ( \30041_30343 , \17736_18035 , \19235_19534 );
and \U$21236 ( \30042_30344 , \18730_19032 , \18743_19045 );
nor \U$21237 ( \30043_30345 , \30041_30343 , \30042_30344 );
xnor \U$21238 ( \30044_30346 , \30043_30345 , \19241_19540 );
xor \U$21239 ( \30045_30347 , \30040_30342 , \30044_30346 );
and \U$21240 ( \30046_30348 , \16353_16655 , \20706_21005 );
and \U$21241 ( \30047_30349 , \17325_17627 , \20255_20557 );
nor \U$21242 ( \30048_30350 , \30046_30348 , \30047_30349 );
xnor \U$21243 ( \30049_30351 , \30048_30350 , \20712_21011 );
xor \U$21244 ( \30050_30352 , \30045_30347 , \30049_30351 );
xor \U$21245 ( \30051_30353 , \30036_30338 , \30050_30352 );
xor \U$21246 ( \30052_30354 , \30027_30329 , \30051_30353 );
xor \U$21247 ( \30053_30355 , \30011_30313 , \30052_30354 );
xor \U$21248 ( \30054_30356 , \29982_30284 , \30053_30355 );
and \U$21249 ( \30055_30357 , \28472_28774 , \28835_29137 );
and \U$21250 ( \30056_30358 , \28835_29137 , \28870_29172 );
and \U$21251 ( \30057_30359 , \28472_28774 , \28870_29172 );
or \U$21252 ( \30058_30360 , \30055_30357 , \30056_30358 , \30057_30359 );
xor \U$21253 ( \30059_30361 , \30054_30356 , \30058_30360 );
and \U$21254 ( \30060_30362 , \28468_28770 , \28871_29173 );
and \U$21255 ( \30061_30363 , \28872_29174 , \28875_29177 );
or \U$21256 ( \30062_30364 , \30060_30362 , \30061_30363 );
xor \U$21257 ( \30063_30365 , \30059_30361 , \30062_30364 );
buf g9bba_GF_PartitionCandidate( \30064_30366_nG9bba , \30063_30365 );
and \U$21258 ( \30065_30367 , \10402_10704 , \30064_30366_nG9bba );
or \U$21259 ( \30066_30368 , \29655_29957 , \30065_30367 );
xor \U$21260 ( \30067_30369 , \10399_10703 , \30066_30368 );
buf \U$21261 ( \30068_30370 , \30067_30369 );
buf \U$21263 ( \30069_30371 , \30068_30370 );
xor \U$21264 ( \30070_30372 , \29654_29956 , \30069_30371 );
buf \U$21265 ( \30071_30373 , \30070_30372 );
xor \U$21266 ( \30072_30374 , \29602_29904 , \30071_30373 );
buf \U$21267 ( \30073_30375 , \30072_30374 );
and \U$21268 ( \30074_30376 , \28409_28711 , \28442_28744 );
and \U$21269 ( \30075_30377 , \28409_28711 , \28448_28750 );
and \U$21270 ( \30076_30378 , \28442_28744 , \28448_28750 );
or \U$21271 ( \30077_30379 , \30074_30376 , \30075_30377 , \30076_30378 );
buf \U$21272 ( \30078_30380 , \30077_30379 );
xor \U$21273 ( \30079_30381 , \30073_30375 , \30078_30380 );
and \U$21274 ( \30080_30382 , \28414_28716 , \28434_28736 );
and \U$21275 ( \30081_30383 , \28414_28716 , \28440_28742 );
and \U$21276 ( \30082_30384 , \28434_28736 , \28440_28742 );
or \U$21277 ( \30083_30385 , \30080_30382 , \30081_30383 , \30082_30384 );
buf \U$21278 ( \30084_30386 , \30083_30385 );
and \U$21279 ( \30085_30387 , \28970_29269 , \28976_29275 );
and \U$21280 ( \30086_30388 , \28970_29269 , \28983_29282 );
and \U$21281 ( \30087_30389 , \28976_29275 , \28983_29282 );
or \U$21282 ( \30088_30390 , \30085_30387 , \30086_30388 , \30087_30389 );
buf \U$21283 ( \30089_30391 , \30088_30390 );
and \U$21284 ( \30090_30392 , \28943_29245 , \28952_29251 );
and \U$21285 ( \30091_30393 , \28943_29245 , \28959_29258 );
and \U$21286 ( \30092_30394 , \28952_29251 , \28959_29258 );
or \U$21287 ( \30093_30395 , \30090_30392 , \30091_30393 , \30092_30394 );
buf \U$21288 ( \30094_30396 , \30093_30395 );
and \U$21289 ( \30095_30397 , \28946_28118 , \10693_10995_nG9c0b );
and \U$21290 ( \30096_30398 , \27816_28115 , \10981_11283_nG9c08 );
or \U$21291 ( \30097_30399 , \30095_30397 , \30096_30398 );
xor \U$21292 ( \30098_30400 , \27815_28114 , \30097_30399 );
buf \U$21293 ( \30099_30401 , \30098_30400 );
buf \U$21295 ( \30100_30402 , \30099_30401 );
and \U$21296 ( \30101_30403 , \27141_26431 , \11299_11598_nG9c05 );
and \U$21297 ( \30102_30404 , \26129_26428 , \12168_12470_nG9c02 );
or \U$21298 ( \30103_30405 , \30101_30403 , \30102_30404 );
xor \U$21299 ( \30104_30406 , \26128_26427 , \30103_30405 );
buf \U$21300 ( \30105_30407 , \30104_30406 );
buf \U$21302 ( \30106_30408 , \30105_30407 );
xor \U$21303 ( \30107_30409 , \30100_30402 , \30106_30408 );
buf \U$21304 ( \30108_30410 , \30107_30409 );
xor \U$21305 ( \30109_30411 , \30094_30396 , \30108_30410 );
and \U$21306 ( \30110_30412 , \21908_21658 , \15074_15373_nG9bf3 );
and \U$21307 ( \30111_30413 , \21356_21655 , \16013_16315_nG9bf0 );
or \U$21308 ( \30112_30414 , \30110_30412 , \30111_30413 );
xor \U$21309 ( \30113_30415 , \21355_21654 , \30112_30414 );
buf \U$21310 ( \30114_30416 , \30113_30415 );
buf \U$21312 ( \30115_30417 , \30114_30416 );
xor \U$21313 ( \30116_30418 , \30109_30411 , \30115_30417 );
buf \U$21314 ( \30117_30419 , \30116_30418 );
and \U$21315 ( \30118_30420 , \18908_18702 , \17808_18107_nG9be7 );
and \U$21316 ( \30119_30421 , \18400_18699 , \18789_19091_nG9be4 );
or \U$21317 ( \30120_30422 , \30118_30420 , \30119_30421 );
xor \U$21318 ( \30121_30423 , \18399_18698 , \30120_30422 );
buf \U$21319 ( \30122_30424 , \30121_30423 );
buf \U$21321 ( \30123_30425 , \30122_30424 );
xor \U$21322 ( \30124_30426 , \30117_30419 , \30123_30425 );
and \U$21323 ( \30125_30427 , \16405_15940 , \20787_21086_nG9bdb );
and \U$21324 ( \30126_30428 , \15638_15937 , \21827_22129_nG9bd8 );
or \U$21325 ( \30127_30429 , \30125_30427 , \30126_30428 );
xor \U$21326 ( \30128_30430 , \15637_15936 , \30127_30429 );
buf \U$21327 ( \30129_30431 , \30128_30430 );
buf \U$21329 ( \30130_30432 , \30129_30431 );
xor \U$21330 ( \30131_30433 , \30124_30426 , \30130_30432 );
buf \U$21331 ( \30132_30434 , \30131_30433 );
xor \U$21332 ( \30133_30435 , \30089_30391 , \30132_30434 );
and \U$21333 ( \30134_30436 , \10996_10421 , \27114_27416_nG9bc3 );
and \U$21334 ( \30135_30437 , \10119_10418 , \28300_28602_nG9bc0 );
or \U$21335 ( \30136_30438 , \30134_30436 , \30135_30437 );
xor \U$21336 ( \30137_30439 , \10118_10417 , \30136_30438 );
buf \U$21337 ( \30138_30440 , \30137_30439 );
buf \U$21339 ( \30139_30441 , \30138_30440 );
xor \U$21340 ( \30140_30442 , \30133_30435 , \30139_30441 );
buf \U$21341 ( \30141_30443 , \30140_30442 );
xor \U$21342 ( \30142_30444 , \30084_30386 , \30141_30443 );
and \U$21343 ( \30143_30445 , \28456_28758 , \28462_28764 );
and \U$21344 ( \30144_30446 , \28456_28758 , \28882_29184 );
and \U$21345 ( \30145_30447 , \28462_28764 , \28882_29184 );
or \U$21346 ( \30146_30448 , \30143_30445 , \30144_30446 , \30145_30447 );
buf \U$21347 ( \30147_30449 , \30146_30448 );
xor \U$21348 ( \30148_30450 , \30142_30444 , \30147_30449 );
buf \U$21349 ( \30149_30451 , \30148_30450 );
xor \U$21350 ( \30150_30452 , \30079_30381 , \30149_30451 );
and \U$21351 ( \30151_30453 , \29558_29860 , \30150_30452 );
and \U$21352 ( \30152_30454 , \29562_29864 , \30150_30452 );
or \U$21353 ( \30153_30455 , \29563_29865 , \30151_30453 , \30152_30454 );
and \U$21354 ( \30154_30456 , \28997_29296 , \29001_29300 );
and \U$21355 ( \30155_30457 , \28997_29296 , \29557_29859 );
and \U$21356 ( \30156_30458 , \29001_29300 , \29557_29859 );
or \U$21357 ( \30157_30459 , \30154_30456 , \30155_30457 , \30156_30458 );
xor \U$21358 ( \30158_30460 , \30153_30455 , \30157_30459 );
and \U$21359 ( \30159_30461 , \30073_30375 , \30078_30380 );
and \U$21360 ( \30160_30462 , \30073_30375 , \30149_30451 );
and \U$21361 ( \30161_30463 , \30078_30380 , \30149_30451 );
or \U$21362 ( \30162_30464 , \30159_30461 , \30160_30462 , \30161_30463 );
xor \U$21363 ( \30163_30465 , \30158_30460 , \30162_30464 );
and \U$21364 ( \30164_30466 , \30094_30396 , \30108_30410 );
and \U$21365 ( \30165_30467 , \30094_30396 , \30115_30417 );
and \U$21366 ( \30166_30468 , \30108_30410 , \30115_30417 );
or \U$21367 ( \30167_30469 , \30164_30466 , \30165_30467 , \30166_30468 );
buf \U$21368 ( \30168_30470 , \30167_30469 );
and \U$21369 ( \30169_30471 , \30100_30402 , \30106_30408 );
buf \U$21370 ( \30170_30472 , \30169_30471 );
and \U$21371 ( \30171_30473 , \25044_24792 , \13403_13705_nG9bfc );
and \U$21372 ( \30172_30474 , \24490_24789 , \13771_14070_nG9bf9 );
or \U$21373 ( \30173_30475 , \30171_30473 , \30172_30474 );
xor \U$21374 ( \30174_30476 , \24489_24788 , \30173_30475 );
buf \U$21375 ( \30175_30477 , \30174_30476 );
buf \U$21377 ( \30176_30478 , \30175_30477 );
xor \U$21378 ( \30177_30479 , \30170_30472 , \30176_30478 );
and \U$21379 ( \30178_30480 , \23495_23201 , \14682_14984_nG9bf6 );
and \U$21380 ( \30179_30481 , \22899_23198 , \15074_15373_nG9bf3 );
or \U$21381 ( \30180_30482 , \30178_30480 , \30179_30481 );
xor \U$21382 ( \30181_30483 , \22898_23197 , \30180_30482 );
buf \U$21383 ( \30182_30484 , \30181_30483 );
buf \U$21385 ( \30183_30485 , \30182_30484 );
xor \U$21386 ( \30184_30486 , \30177_30479 , \30183_30485 );
buf \U$21387 ( \30185_30487 , \30184_30486 );
xor \U$21388 ( \30186_30488 , \30168_30470 , \30185_30487 );
and \U$21389 ( \30187_30489 , \20353_20155 , \17363_17665_nG9bea );
and \U$21390 ( \30188_30490 , \19853_20152 , \17808_18107_nG9be7 );
or \U$21391 ( \30189_30491 , \30187_30489 , \30188_30490 );
xor \U$21392 ( \30190_30492 , \19852_20151 , \30189_30491 );
buf \U$21393 ( \30191_30493 , \30190_30492 );
buf \U$21395 ( \30192_30494 , \30191_30493 );
xor \U$21396 ( \30193_30495 , \30186_30488 , \30192_30494 );
buf \U$21397 ( \30194_30496 , \30193_30495 );
and \U$21398 ( \30195_30497 , \29612_29914 , \29629_29931 );
and \U$21399 ( \30196_30498 , \29612_29914 , \29636_29938 );
and \U$21400 ( \30197_30499 , \29629_29931 , \29636_29938 );
or \U$21401 ( \30198_30500 , \30195_30497 , \30196_30498 , \30197_30499 );
buf \U$21402 ( \30199_30501 , \30198_30500 );
xor \U$21403 ( \30200_30502 , \30194_30496 , \30199_30501 );
and \U$21404 ( \30201_30503 , \16405_15940 , \21827_22129_nG9bd8 );
and \U$21405 ( \30202_30504 , \15638_15937 , \22330_22629_nG9bd5 );
or \U$21406 ( \30203_30505 , \30201_30503 , \30202_30504 );
xor \U$21407 ( \30204_30506 , \15637_15936 , \30203_30505 );
buf \U$21408 ( \30205_30507 , \30204_30506 );
buf \U$21410 ( \30206_30508 , \30205_30507 );
xor \U$21411 ( \30207_30509 , \30200_30502 , \30206_30508 );
buf \U$21412 ( \30208_30510 , \30207_30509 );
and \U$21413 ( \30209_30511 , \29607_29909 , \29638_29940 );
and \U$21414 ( \30210_30512 , \29607_29909 , \29645_29947 );
and \U$21415 ( \30211_30513 , \29638_29940 , \29645_29947 );
or \U$21416 ( \30212_30514 , \30209_30511 , \30210_30512 , \30211_30513 );
buf \U$21417 ( \30213_30515 , \30212_30514 );
xor \U$21418 ( \30214_30516 , \30208_30510 , \30213_30515 );
and \U$21419 ( \30215_30517 , \10411_10707 , \30064_30366_nG9bba );
and \U$21420 ( \30216_30518 , \29663_29965 , \29667_29969 );
and \U$21421 ( \30217_30519 , \29667_29969 , \29980_30282 );
and \U$21422 ( \30218_30520 , \29663_29965 , \29980_30282 );
or \U$21423 ( \30219_30521 , \30216_30518 , \30217_30519 , \30218_30520 );
and \U$21424 ( \30220_30522 , \29986_30288 , \30010_30312 );
and \U$21425 ( \30221_30523 , \30010_30312 , \30052_30354 );
and \U$21426 ( \30222_30524 , \29986_30288 , \30052_30354 );
or \U$21427 ( \30223_30525 , \30220_30522 , \30221_30523 , \30222_30524 );
xor \U$21428 ( \30224_30526 , \30219_30521 , \30223_30525 );
and \U$21429 ( \30225_30527 , \30019_30321 , \30023_30325 );
and \U$21430 ( \30226_30528 , \30023_30325 , \30025_30327 );
and \U$21431 ( \30227_30529 , \30019_30321 , \30025_30327 );
or \U$21432 ( \30228_30530 , \30225_30527 , \30226_30528 , \30227_30529 );
and \U$21433 ( \30229_30531 , \29946_30248 , \29960_30262 );
and \U$21434 ( \30230_30532 , \29960_30262 , \29979_30281 );
and \U$21435 ( \30231_30533 , \29946_30248 , \29979_30281 );
or \U$21436 ( \30232_30534 , \30229_30531 , \30230_30532 , \30231_30533 );
xor \U$21437 ( \30233_30535 , \30228_30530 , \30232_30534 );
and \U$21438 ( \30234_30536 , \29966_30268 , \10681_10983 );
and \U$21439 ( \30235_30537 , RIdec5f18_716, \9034_9333 );
and \U$21440 ( \30236_30538 , RIdec3218_684, \9036_9335 );
and \U$21441 ( \30237_30539 , RIee20350_4825, \9038_9337 );
and \U$21442 ( \30238_30540 , RIdec0518_652, \9040_9339 );
and \U$21443 ( \30239_30541 , RIee1f6a8_4816, \9042_9341 );
and \U$21444 ( \30240_30542 , RIdebd818_620, \9044_9343 );
and \U$21445 ( \30241_30543 , RIdebab18_588, \9046_9345 );
and \U$21446 ( \30242_30544 , RIdeb7e18_556, \9048_9347 );
and \U$21447 ( \30243_30545 , RIfce4da0_7626, \9050_9349 );
and \U$21448 ( \30244_30546 , RIdeb2418_492, \9052_9351 );
and \U$21449 ( \30245_30547 , RIfcea908_7691, \9054_9353 );
and \U$21450 ( \30246_30548 , RIdeaf718_460, \9056_9355 );
and \U$21451 ( \30247_30549 , RIfce20a0_7594, \9058_9357 );
and \U$21452 ( \30248_30550 , RIdeabe60_428, \9060_9359 );
and \U$21453 ( \30249_30551 , RIdea5560_396, \9062_9361 );
and \U$21454 ( \30250_30552 , RIde9ec60_364, \9064_9363 );
and \U$21455 ( \30251_30553 , RIfce6420_7642, \9066_9365 );
and \U$21456 ( \30252_30554 , RIee1c2a0_4779, \9068_9367 );
and \U$21457 ( \30253_30555 , RIfc75950_6360, \9070_9369 );
and \U$21458 ( \30254_30556 , RIee1ad88_4764, \9072_9371 );
and \U$21459 ( \30255_30557 , RIde920f0_302, \9074_9373 );
and \U$21460 ( \30256_30558 , RIfea4148_8211, \9076_9375 );
and \U$21461 ( \30257_30559 , RIfeaa688_8255, \9078_9377 );
and \U$21462 ( \30258_30560 , RIfea3fe0_8210, \9080_9379 );
and \U$21463 ( \30259_30561 , RIde82790_226, \9082_9381 );
and \U$21464 ( \30260_30562 , RIfc6f848_6291, \9084_9383 );
and \U$21465 ( \30261_30563 , RIfc5dc38_6089, \9086_9385 );
and \U$21466 ( \30262_30564 , RIfc76b98_6373, \9088_9387 );
and \U$21467 ( \30263_30565 , RIfcae2f0_7004, \9090_9389 );
and \U$21468 ( \30264_30566 , RIe16c020_2606, \9092_9391 );
and \U$21469 ( \30265_30567 , RIe16a130_2584, \9094_9393 );
and \U$21470 ( \30266_30568 , RIe1687e0_2566, \9096_9395 );
and \U$21471 ( \30267_30569 , RIe165f18_2537, \9098_9397 );
and \U$21472 ( \30268_30570 , RIe163218_2505, \9100_9399 );
and \U$21473 ( \30269_30571 , RIfcadd50_7000, \9102_9401 );
and \U$21474 ( \30270_30572 , RIe160518_2473, \9104_9403 );
and \U$21475 ( \30271_30573 , RIfc55268_5991, \9106_9405 );
and \U$21476 ( \30272_30574 , RIe15d818_2441, \9108_9407 );
and \U$21477 ( \30273_30575 , RIe157e18_2377, \9110_9409 );
and \U$21478 ( \30274_30576 , RIe155118_2345, \9112_9411 );
and \U$21479 ( \30275_30577 , RIfc45548_5811, \9114_9413 );
and \U$21480 ( \30276_30578 , RIe152418_2313, \9116_9415 );
and \U$21481 ( \30277_30579 , RIfc498c8_5859, \9118_9417 );
and \U$21482 ( \30278_30580 , RIe14f718_2281, \9120_9419 );
and \U$21483 ( \30279_30581 , RIfcbda70_7180, \9122_9421 );
and \U$21484 ( \30280_30582 , RIe14ca18_2249, \9124_9423 );
and \U$21485 ( \30281_30583 , RIe149d18_2217, \9126_9425 );
and \U$21486 ( \30282_30584 , RIe147018_2185, \9128_9427 );
and \U$21487 ( \30283_30585 , RIee34828_5056, \9130_9429 );
and \U$21488 ( \30284_30586 , RIee33748_5044, \9132_9431 );
and \U$21489 ( \30285_30587 , RIee32668_5032, \9134_9433 );
and \U$21490 ( \30286_30588 , RIee31588_5020, \9136_9435 );
and \U$21491 ( \30287_30589 , RIe1418e8_2123, \9138_9437 );
and \U$21492 ( \30288_30590 , RIe13f458_2097, \9140_9439 );
and \U$21493 ( \30289_30591 , RIdf3d360_2073, \9142_9441 );
and \U$21494 ( \30290_30592 , RIdf3aed0_2047, \9144_9443 );
and \U$21495 ( \30291_30593 , RIfc526d0_5960, \9146_9445 );
and \U$21496 ( \30292_30594 , RIfc42848_5779, \9148_9447 );
and \U$21497 ( \30293_30595 , RIfcae9f8_7009, \9150_9449 );
and \U$21498 ( \30294_30596 , RIfcb7260_7106, \9152_9451 );
and \U$21499 ( \30295_30597 , RIfea42b0_8212, \9154_9453 );
and \U$21500 ( \30296_30598 , RIdf33ce8_1966, \9156_9455 );
and \U$21501 ( \30297_30599 , RIdf31b28_1942, \9158_9457 );
and \U$21502 ( \30298_30600 , RIdf2fc38_1920, \9160_9459 );
or \U$21503 ( \30299_30601 , \30235_30537 , \30236_30538 , \30237_30539 , \30238_30540 , \30239_30541 , \30240_30542 , \30241_30543 , \30242_30544 , \30243_30545 , \30244_30546 , \30245_30547 , \30246_30548 , \30247_30549 , \30248_30550 , \30249_30551 , \30250_30552 , \30251_30553 , \30252_30554 , \30253_30555 , \30254_30556 , \30255_30557 , \30256_30558 , \30257_30559 , \30258_30560 , \30259_30561 , \30260_30562 , \30261_30563 , \30262_30564 , \30263_30565 , \30264_30566 , \30265_30567 , \30266_30568 , \30267_30569 , \30268_30570 , \30269_30571 , \30270_30572 , \30271_30573 , \30272_30574 , \30273_30575 , \30274_30576 , \30275_30577 , \30276_30578 , \30277_30579 , \30278_30580 , \30279_30581 , \30280_30582 , \30281_30583 , \30282_30584 , \30283_30585 , \30284_30586 , \30285_30587 , \30286_30588 , \30287_30589 , \30288_30590 , \30289_30591 , \30290_30592 , \30291_30593 , \30292_30594 , \30293_30595 , \30294_30596 , \30295_30597 , \30296_30598 , \30297_30599 , \30298_30600 );
and \U$21504 ( \30300_30602 , RIee2c3f8_4962, \9163_9462 );
and \U$21505 ( \30301_30603 , RIfc4cfa0_5898, \9165_9464 );
and \U$21506 ( \30302_30604 , RIfc572c0_6014, \9167_9466 );
and \U$21507 ( \30303_30605 , RIfc4f430_5924, \9169_9468 );
and \U$21508 ( \30304_30606 , RIfea3e78_8209, \9171_9470 );
and \U$21509 ( \30305_30607 , RIdf28a50_1839, \9173_9472 );
and \U$21510 ( \30306_30608 , RIdf26b60_1817, \9175_9474 );
and \U$21511 ( \30307_30609 , RIdf250a8_1798, \9177_9476 );
and \U$21512 ( \30308_30610 , RIfc9b600_6790, \9179_9478 );
and \U$21513 ( \30309_30611 , RIfcb9df8_7137, \9181_9480 );
and \U$21514 ( \30310_30612 , RIdf23320_1777, \9183_9482 );
and \U$21515 ( \30311_30613 , RIfc86318_6549, \9185_9484 );
and \U$21516 ( \30312_30614 , RIfeabfd8_8273, \9187_9486 );
and \U$21517 ( \30313_30615 , RIdf201e8_1742, \9189_9488 );
and \U$21518 ( \30314_30616 , RIdf1b5f8_1688, \9191_9490 );
and \U$21519 ( \30315_30617 , RIdf19ca8_1670, \9193_9492 );
and \U$21520 ( \30316_30618 , RIdf17ae8_1646, \9195_9494 );
and \U$21521 ( \30317_30619 , RIdf14de8_1614, \9197_9496 );
and \U$21522 ( \30318_30620 , RIdf120e8_1582, \9199_9498 );
and \U$21523 ( \30319_30621 , RIdf0f3e8_1550, \9201_9500 );
and \U$21524 ( \30320_30622 , RIdf0c6e8_1518, \9203_9502 );
and \U$21525 ( \30321_30623 , RIdf099e8_1486, \9205_9504 );
and \U$21526 ( \30322_30624 , RIdf06ce8_1454, \9207_9506 );
and \U$21527 ( \30323_30625 , RIdf03fe8_1422, \9209_9508 );
and \U$21528 ( \30324_30626 , RIdefe5e8_1358, \9211_9510 );
and \U$21529 ( \30325_30627 , RIdefb8e8_1326, \9213_9512 );
and \U$21530 ( \30326_30628 , RIdef8be8_1294, \9215_9514 );
and \U$21531 ( \30327_30629 , RIdef5ee8_1262, \9217_9516 );
and \U$21532 ( \30328_30630 , RIdef31e8_1230, \9219_9518 );
and \U$21533 ( \30329_30631 , RIdef04e8_1198, \9221_9520 );
and \U$21534 ( \30330_30632 , RIdeed7e8_1166, \9223_9522 );
and \U$21535 ( \30331_30633 , RIdeeaae8_1134, \9225_9524 );
and \U$21536 ( \30332_30634 , RIfc89018_6581, \9227_9526 );
and \U$21537 ( \30333_30635 , RIfcc54c8_7267, \9229_9528 );
and \U$21538 ( \30334_30636 , RIfc89180_6582, \9231_9530 );
and \U$21539 ( \30335_30637 , RIfc4b380_5878, \9233_9532 );
and \U$21540 ( \30336_30638 , RIdee53b8_1072, \9235_9534 );
and \U$21541 ( \30337_30639 , RIdee34c8_1050, \9237_9536 );
and \U$21542 ( \30338_30640 , RIfea3d10_8208, \9239_9538 );
and \U$21543 ( \30339_30641 , RIdedf148_1002, \9241_9540 );
and \U$21544 ( \30340_30642 , RIfcae188_7003, \9243_9542 );
and \U$21545 ( \30341_30643 , RIfc4b0b0_5876, \9245_9544 );
and \U$21546 ( \30342_30644 , RIfc74870_6348, \9247_9546 );
and \U$21547 ( \30343_30645 , RIfce4968_7623, \9249_9548 );
and \U$21548 ( \30344_30646 , RIdeda288_946, \9251_9550 );
and \U$21549 ( \30345_30647 , RIded7c90_919, \9253_9552 );
and \U$21550 ( \30346_30648 , RIded5da0_897, \9255_9554 );
and \U$21551 ( \30347_30649 , RIded3640_869, \9257_9556 );
and \U$21552 ( \30348_30650 , RIded1318_844, \9259_9558 );
and \U$21553 ( \30349_30651 , RIdece618_812, \9261_9560 );
and \U$21554 ( \30350_30652 , RIdecb918_780, \9263_9562 );
and \U$21555 ( \30351_30653 , RIdec8c18_748, \9265_9564 );
and \U$21556 ( \30352_30654 , RIdeb5118_524, \9267_9566 );
and \U$21557 ( \30353_30655 , RIde98360_332, \9269_9568 );
and \U$21558 ( \30354_30656 , RIe16ed20_2638, \9271_9570 );
and \U$21559 ( \30355_30657 , RIe15ab18_2409, \9273_9572 );
and \U$21560 ( \30356_30658 , RIe144318_2153, \9275_9574 );
and \U$21561 ( \30357_30659 , RIdf38d10_2023, \9277_9576 );
and \U$21562 ( \30358_30660 , RIdf2d370_1891, \9279_9578 );
and \U$21563 ( \30359_30661 , RIdf1dbf0_1715, \9281_9580 );
and \U$21564 ( \30360_30662 , RIdf012e8_1390, \9283_9582 );
and \U$21565 ( \30361_30663 , RIdee7de8_1102, \9285_9584 );
and \U$21566 ( \30362_30664 , RIdedcb50_975, \9287_9586 );
and \U$21567 ( \30363_30665 , RIde7e2a8_205, \9289_9588 );
or \U$21568 ( \30364_30666 , \30300_30602 , \30301_30603 , \30302_30604 , \30303_30605 , \30304_30606 , \30305_30607 , \30306_30608 , \30307_30609 , \30308_30610 , \30309_30611 , \30310_30612 , \30311_30613 , \30312_30614 , \30313_30615 , \30314_30616 , \30315_30617 , \30316_30618 , \30317_30619 , \30318_30620 , \30319_30621 , \30320_30622 , \30321_30623 , \30322_30624 , \30323_30625 , \30324_30626 , \30325_30627 , \30326_30628 , \30327_30629 , \30328_30630 , \30329_30631 , \30330_30632 , \30331_30633 , \30332_30634 , \30333_30635 , \30334_30636 , \30335_30637 , \30336_30638 , \30337_30639 , \30338_30640 , \30339_30641 , \30340_30642 , \30341_30643 , \30342_30644 , \30343_30645 , \30344_30646 , \30345_30647 , \30346_30648 , \30347_30649 , \30348_30650 , \30349_30651 , \30350_30652 , \30351_30653 , \30352_30654 , \30353_30655 , \30354_30656 , \30355_30657 , \30356_30658 , \30357_30659 , \30358_30660 , \30359_30661 , \30360_30662 , \30361_30663 , \30362_30664 , \30363_30665 );
or \U$21569 ( \30365_30667 , \30299_30601 , \30364_30666 );
_DC \g65ce/U$1 ( \30366 , \30365_30667 , \9298_9597 );
and \U$21570 ( \30367_30669 , RIe19e1b0_3176, \8760_9059 );
and \U$21571 ( \30368_30670 , RIe19b4b0_3144, \8762_9061 );
and \U$21572 ( \30369_30671 , RIfc9cf50_6808, \8764_9063 );
and \U$21573 ( \30370_30672 , RIe1987b0_3112, \8766_9065 );
and \U$21574 ( \30371_30673 , RIfc87290_6560, \8768_9067 );
and \U$21575 ( \30372_30674 , RIe195ab0_3080, \8770_9069 );
and \U$21576 ( \30373_30675 , RIe192db0_3048, \8772_9071 );
and \U$21577 ( \30374_30676 , RIe1900b0_3016, \8774_9073 );
and \U$21578 ( \30375_30677 , RIe18a6b0_2952, \8776_9075 );
and \U$21579 ( \30376_30678 , RIe1879b0_2920, \8778_9077 );
and \U$21580 ( \30377_30679 , RIfc842c0_6526, \8780_9079 );
and \U$21581 ( \30378_30680 , RIe184cb0_2888, \8782_9081 );
and \U$21582 ( \30379_30681 , RIfc83a50_6520, \8784_9083 );
and \U$21583 ( \30380_30682 , RIe181fb0_2856, \8786_9085 );
and \U$21584 ( \30381_30683 , RIe17f2b0_2824, \8788_9087 );
and \U$21585 ( \30382_30684 , RIe17c5b0_2792, \8790_9089 );
and \U$21586 ( \30383_30685 , RIfc9d0b8_6809, \8792_9091 );
and \U$21587 ( \30384_30686 , RIfc9e030_6820, \8794_9093 );
and \U$21588 ( \30385_30687 , RIe177420_2734, \8796_9095 );
and \U$21589 ( \30386_30688 , RIe176340_2722, \8798_9097 );
and \U$21590 ( \30387_30689 , RIfc4f700_5926, \8800_9099 );
and \U$21591 ( \30388_30690 , RIfcc4820_7258, \8802_9101 );
and \U$21592 ( \30389_30691 , RIfc4fb38_5929, \8804_9103 );
and \U$21593 ( \30390_30692 , RIfce8040_7662, \8806_9105 );
and \U$21594 ( \30391_30693 , RIee3c6b8_5146, \8808_9107 );
and \U$21595 ( \30392_30694 , RIee3b308_5132, \8810_9109 );
and \U$21596 ( \30393_30695 , RIfc812f0_6492, \8812_9111 );
and \U$21597 ( \30394_30696 , RIe174180_2698, \8814_9113 );
and \U$21598 ( \30395_30697 , RIfcd3028_7423, \8816_9115 );
and \U$21599 ( \30396_30698 , RIfc7f400_6470, \8818_9117 );
and \U$21600 ( \30397_30699 , RIfc46a60_5826, \8820_9119 );
and \U$21601 ( \30398_30700 , RIfc472d0_5832, \8822_9121 );
and \U$21602 ( \30399_30701 , RIf16cc58_5697, \8824_9123 );
and \U$21603 ( \30400_30702 , RIe224508_4703, \8826_9125 );
and \U$21604 ( \30401_30703 , RIfc7d3a8_6447, \8828_9127 );
and \U$21605 ( \30402_30704 , RIe221808_4671, \8830_9129 );
and \U$21606 ( \30403_30705 , RIfc97c58_6749, \8832_9131 );
and \U$21607 ( \30404_30706 , RIe21eb08_4639, \8834_9133 );
and \U$21608 ( \30405_30707 , RIe219108_4575, \8836_9135 );
and \U$21609 ( \30406_30708 , RIe216408_4543, \8838_9137 );
and \U$21610 ( \30407_30709 , RIfcdbe30_7524, \8840_9139 );
and \U$21611 ( \30408_30710 , RIe213708_4511, \8842_9141 );
and \U$21612 ( \30409_30711 , RIf169580_5658, \8844_9143 );
and \U$21613 ( \30410_30712 , RIe210a08_4479, \8846_9145 );
and \U$21614 ( \30411_30713 , RIfca4570_6892, \8848_9147 );
and \U$21615 ( \30412_30714 , RIe20dd08_4447, \8850_9149 );
and \U$21616 ( \30413_30715 , RIe20b008_4415, \8852_9151 );
and \U$21617 ( \30414_30716 , RIe208308_4383, \8854_9153 );
and \U$21618 ( \30415_30717 , RIfc7b080_6422, \8856_9155 );
and \U$21619 ( \30416_30718 , RIfc59cf0_6044, \8858_9157 );
and \U$21620 ( \30417_30719 , RIfea9b48_8247, \8860_9159 );
and \U$21621 ( \30418_30720 , RIfea4418_8213, \8862_9161 );
and \U$21622 ( \30419_30721 , RIfc79cd0_6408, \8864_9163 );
and \U$21623 ( \30420_30722 , RIfcd19a8_7407, \8866_9165 );
and \U$21624 ( \30421_30723 , RIfcc81c8_7299, \8868_9167 );
and \U$21625 ( \30422_30724 , RIf162230_5576, \8870_9169 );
and \U$21626 ( \30423_30725 , RIf160778_5557, \8872_9171 );
and \U$21627 ( \30424_30726 , RIf15e888_5535, \8874_9173 );
and \U$21628 ( \30425_30727 , RIfea4580_8214, \8876_9175 );
and \U$21629 ( \30426_30728 , RIfea46e8_8215, \8878_9177 );
and \U$21630 ( \30427_30729 , RIfc77f48_6387, \8880_9179 );
and \U$21631 ( \30428_30730 , RIfc41fd8_5773, \8882_9181 );
and \U$21632 ( \30429_30731 , RIf15aaa8_5491, \8884_9183 );
and \U$21633 ( \30430_30732 , RIfc7c430_6436, \8886_9185 );
or \U$21634 ( \30431_30733 , \30367_30669 , \30368_30670 , \30369_30671 , \30370_30672 , \30371_30673 , \30372_30674 , \30373_30675 , \30374_30676 , \30375_30677 , \30376_30678 , \30377_30679 , \30378_30680 , \30379_30681 , \30380_30682 , \30381_30683 , \30382_30684 , \30383_30685 , \30384_30686 , \30385_30687 , \30386_30688 , \30387_30689 , \30388_30690 , \30389_30691 , \30390_30692 , \30391_30693 , \30392_30694 , \30393_30695 , \30394_30696 , \30395_30697 , \30396_30698 , \30397_30699 , \30398_30700 , \30399_30701 , \30400_30702 , \30401_30703 , \30402_30704 , \30403_30705 , \30404_30706 , \30405_30707 , \30406_30708 , \30407_30709 , \30408_30710 , \30409_30711 , \30410_30712 , \30411_30713 , \30412_30714 , \30413_30715 , \30414_30716 , \30415_30717 , \30416_30718 , \30417_30719 , \30418_30720 , \30419_30721 , \30420_30722 , \30421_30723 , \30422_30724 , \30423_30725 , \30424_30726 , \30425_30727 , \30426_30728 , \30427_30729 , \30428_30730 , \30429_30731 , \30430_30732 );
and \U$21635 ( \30432_30734 , RIf159158_5473, \8889_9188 );
and \U$21636 ( \30433_30735 , RIf157f10_5460, \8891_9190 );
and \U$21637 ( \30434_30736 , RIfcae890_7008, \8893_9192 );
and \U$21638 ( \30435_30737 , RIe1faa78_4229, \8895_9194 );
and \U$21639 ( \30436_30738 , RIfc4a840_5870, \8897_9196 );
and \U$21640 ( \30437_30739 , RIfc4ed28_5919, \8899_9198 );
and \U$21641 ( \30438_30740 , RIfce0e58_7581, \8901_9200 );
and \U$21642 ( \30439_30741 , RIe1f5ff0_4176, \8903_9202 );
and \U$21643 ( \30440_30742 , RIf153758_5409, \8905_9204 );
and \U$21644 ( \30441_30743 , RIf151f70_5392, \8907_9206 );
and \U$21645 ( \30442_30744 , RIfccb468_7335, \8909_9208 );
and \U$21646 ( \30443_30745 , RIe1f3cc8_4151, \8911_9210 );
and \U$21647 ( \30444_30746 , RIfc68ed0_6216, \8913_9212 );
and \U$21648 ( \30445_30747 , RIfc6d250_6264, \8915_9214 );
and \U$21649 ( \30446_30748 , RIfca9ca0_6954, \8917_9216 );
and \U$21650 ( \30447_30749 , RIe1ee9d0_4092, \8919_9218 );
and \U$21651 ( \30448_30750 , RIe1ec270_4064, \8921_9220 );
and \U$21652 ( \30449_30751 , RIe1e9570_4032, \8923_9222 );
and \U$21653 ( \30450_30752 , RIe1e6870_4000, \8925_9224 );
and \U$21654 ( \30451_30753 , RIe1e3b70_3968, \8927_9226 );
and \U$21655 ( \30452_30754 , RIe1e0e70_3936, \8929_9228 );
and \U$21656 ( \30453_30755 , RIe1de170_3904, \8931_9230 );
and \U$21657 ( \30454_30756 , RIe1db470_3872, \8933_9232 );
and \U$21658 ( \30455_30757 , RIe1d8770_3840, \8935_9234 );
and \U$21659 ( \30456_30758 , RIe1d2d70_3776, \8937_9236 );
and \U$21660 ( \30457_30759 , RIe1d0070_3744, \8939_9238 );
and \U$21661 ( \30458_30760 , RIe1cd370_3712, \8941_9240 );
and \U$21662 ( \30459_30761 , RIe1ca670_3680, \8943_9242 );
and \U$21663 ( \30460_30762 , RIe1c7970_3648, \8945_9244 );
and \U$21664 ( \30461_30763 , RIe1c4c70_3616, \8947_9246 );
and \U$21665 ( \30462_30764 , RIe1c1f70_3584, \8949_9248 );
and \U$21666 ( \30463_30765 , RIe1bf270_3552, \8951_9250 );
and \U$21667 ( \30464_30766 , RIfc784e8_6391, \8953_9252 );
and \U$21668 ( \30465_30767 , RIfcbef88_7195, \8955_9254 );
and \U$21669 ( \30466_30768 , RIe1b9ca8_3491, \8957_9256 );
and \U$21670 ( \30467_30769 , RIe1b7ae8_3467, \8959_9258 );
and \U$21671 ( \30468_30770 , RIfcc20c0_7230, \8961_9260 );
and \U$21672 ( \30469_30771 , RIfca6190_6912, \8963_9262 );
and \U$21673 ( \30470_30772 , RIe1b5928_3443, \8965_9264 );
and \U$21674 ( \30471_30773 , RIe1b4410_3428, \8967_9266 );
and \U$21675 ( \30472_30774 , RIfcb81d8_7117, \8969_9268 );
and \U$21676 ( \30473_30775 , RIfcc5090_7264, \8971_9270 );
and \U$21677 ( \30474_30776 , RIe1b2d90_3412, \8973_9272 );
and \U$21678 ( \30475_30777 , RIe1b1440_3394, \8975_9274 );
and \U$21679 ( \30476_30778 , RIfcd5350_7448, \8977_9276 );
and \U$21680 ( \30477_30779 , RIfcb9588_7131, \8979_9278 );
and \U$21681 ( \30478_30780 , RIe1acc88_3343, \8981_9280 );
and \U$21682 ( \30479_30781 , RIe1ab4a0_3326, \8983_9282 );
and \U$21683 ( \30480_30782 , RIe1a95b0_3304, \8985_9284 );
and \U$21684 ( \30481_30783 , RIe1a68b0_3272, \8987_9286 );
and \U$21685 ( \30482_30784 , RIe1a3bb0_3240, \8989_9288 );
and \U$21686 ( \30483_30785 , RIe1a0eb0_3208, \8991_9290 );
and \U$21687 ( \30484_30786 , RIe18d3b0_2984, \8993_9292 );
and \U$21688 ( \30485_30787 , RIe1798b0_2760, \8995_9294 );
and \U$21689 ( \30486_30788 , RIe227208_4735, \8997_9296 );
and \U$21690 ( \30487_30789 , RIe21be08_4607, \8999_9298 );
and \U$21691 ( \30488_30790 , RIe205608_4351, \9001_9300 );
and \U$21692 ( \30489_30791 , RIe1ff668_4283, \9003_9302 );
and \U$21693 ( \30490_30792 , RIe1f8a20_4206, \9005_9304 );
and \U$21694 ( \30491_30793 , RIe1f1568_4123, \9007_9306 );
and \U$21695 ( \30492_30794 , RIe1d5a70_3808, \9009_9308 );
and \U$21696 ( \30493_30795 , RIe1bc570_3520, \9011_9310 );
and \U$21697 ( \30494_30796 , RIe1af3e8_3371, \9013_9312 );
and \U$21698 ( \30495_30797 , RIe171a20_2670, \9015_9314 );
or \U$21699 ( \30496_30798 , \30432_30734 , \30433_30735 , \30434_30736 , \30435_30737 , \30436_30738 , \30437_30739 , \30438_30740 , \30439_30741 , \30440_30742 , \30441_30743 , \30442_30744 , \30443_30745 , \30444_30746 , \30445_30747 , \30446_30748 , \30447_30749 , \30448_30750 , \30449_30751 , \30450_30752 , \30451_30753 , \30452_30754 , \30453_30755 , \30454_30756 , \30455_30757 , \30456_30758 , \30457_30759 , \30458_30760 , \30459_30761 , \30460_30762 , \30461_30763 , \30462_30764 , \30463_30765 , \30464_30766 , \30465_30767 , \30466_30768 , \30467_30769 , \30468_30770 , \30469_30771 , \30470_30772 , \30471_30773 , \30472_30774 , \30473_30775 , \30474_30776 , \30475_30777 , \30476_30778 , \30477_30779 , \30478_30780 , \30479_30781 , \30480_30782 , \30481_30783 , \30482_30784 , \30483_30785 , \30484_30786 , \30485_30787 , \30486_30788 , \30487_30789 , \30488_30790 , \30489_30791 , \30490_30792 , \30491_30793 , \30492_30794 , \30493_30795 , \30494_30796 , \30495_30797 );
or \U$21700 ( \30497_30799 , \30431_30733 , \30496_30798 );
_DC \g65cf/U$1 ( \30498 , \30497_30799 , \9024_9323 );
and g65d0_GF_PartitionCandidate( \30499_30801_nG65d0 , \30366 , \30498 );
buf \U$21701 ( \30500_30802 , \30499_30801_nG65d0 );
and \U$21702 ( \30501_30803 , \30500_30802 , \10389_10691 );
nor \U$21703 ( \30502_30804 , \30234_30536 , \30501_30803 );
xnor \U$21704 ( \30503_30805 , \30502_30804 , \10678_10980 );
not \U$21705 ( \30504_30806 , \29945_30247 );
_DC \g62df/U$1 ( \30505 , \30365_30667 , \9298_9597 );
_DC \g6363/U$1 ( \30506 , \30497_30799 , \9024_9323 );
xor g6364_GF_PartitionCandidate( \30507_30809_nG6364 , \30505 , \30506 );
buf \U$21706 ( \30508_30810 , \30507_30809_nG6364 );
and \U$21707 ( \30509_30811 , \29943_30245 , \28765_29067 );
not \U$21708 ( \30510_30812 , \30509_30811 );
and \U$21709 ( \30511_30813 , \30508_30810 , \30510_30812 );
and \U$21710 ( \30512_30814 , \30504_30806 , \30511_30813 );
xor \U$21711 ( \30513_30815 , \30503_30805 , \30512_30814 );
and \U$21712 ( \30514_30816 , \10968_11270 , \28768_29070 );
and \U$21713 ( \30515_30817 , \11287_11586 , \28224_28526 );
nor \U$21714 ( \30516_30818 , \30514_30816 , \30515_30817 );
xnor \U$21715 ( \30517_30819 , \30516_30818 , \28774_29076 );
xor \U$21716 ( \30518_30820 , \30513_30815 , \30517_30819 );
xor \U$21717 ( \30519_30821 , \30508_30810 , \29943_30245 );
not \U$21718 ( \30520_30822 , \29944_30246 );
and \U$21719 ( \30521_30823 , \30519_30821 , \30520_30822 );
and \U$21720 ( \30522_30824 , \10385_10687 , \30521_30823 );
and \U$21721 ( \30523_30825 , \10686_10988 , \29944_30246 );
nor \U$21722 ( \30524_30826 , \30522_30824 , \30523_30825 );
xnor \U$21723 ( \30525_30827 , \30524_30826 , \30511_30813 );
xor \U$21724 ( \30526_30828 , \30518_30820 , \30525_30827 );
xor \U$21725 ( \30527_30829 , \30233_30535 , \30526_30828 );
and \U$21726 ( \30528_30830 , \30031_30333 , \30035_30337 );
and \U$21727 ( \30529_30831 , \30035_30337 , \30050_30352 );
and \U$21728 ( \30530_30832 , \30031_30333 , \30050_30352 );
or \U$21729 ( \30531_30833 , \30528_30830 , \30529_30831 , \30530_30832 );
and \U$21730 ( \30532_30834 , \29672_29974 , \29676_29978 );
and \U$21731 ( \30533_30835 , \29676_29978 , \29945_30247 );
and \U$21732 ( \30534_30836 , \29672_29974 , \29945_30247 );
or \U$21733 ( \30535_30837 , \30532_30834 , \30533_30835 , \30534_30836 );
and \U$21734 ( \30536_30838 , \29969_30271 , \29973_30275 );
and \U$21735 ( \30537_30839 , \29973_30275 , \29978_30280 );
and \U$21736 ( \30538_30840 , \29969_30271 , \29978_30280 );
or \U$21737 ( \30539_30841 , \30536_30838 , \30537_30839 , \30538_30840 );
xor \U$21738 ( \30540_30842 , \30535_30837 , \30539_30841 );
and \U$21739 ( \30541_30843 , \30040_30342 , \30044_30346 );
and \U$21740 ( \30542_30844 , \30044_30346 , \30049_30351 );
and \U$21741 ( \30543_30845 , \30040_30342 , \30049_30351 );
or \U$21742 ( \30544_30846 , \30541_30843 , \30542_30844 , \30543_30845 );
xor \U$21743 ( \30545_30847 , \30540_30842 , \30544_30846 );
xor \U$21744 ( \30546_30848 , \30531_30833 , \30545_30847 );
and \U$21745 ( \30547_30849 , \29950_30252 , \29954_30256 );
and \U$21746 ( \30548_30850 , \29954_30256 , \29959_30261 );
and \U$21747 ( \30549_30851 , \29950_30252 , \29959_30261 );
or \U$21748 ( \30550_30852 , \30547_30849 , \30548_30850 , \30549_30851 );
and \U$21749 ( \30551_30853 , \29999_30301 , \30003_30305 );
and \U$21750 ( \30552_30854 , \30003_30305 , \30008_30310 );
and \U$21751 ( \30553_30855 , \29999_30301 , \30008_30310 );
or \U$21752 ( \30554_30856 , \30551_30853 , \30552_30854 , \30553_30855 );
xor \U$21753 ( \30555_30857 , \30550_30852 , \30554_30856 );
and \U$21754 ( \30556_30858 , \28232_28534 , \11275_11574 );
and \U$21755 ( \30557_30859 , \28782_29084 , \10976_11278 );
nor \U$21756 ( \30558_30860 , \30556_30858 , \30557_30859 );
xnor \U$21757 ( \30559_30861 , \30558_30860 , \11281_11580 );
and \U$21758 ( \30560_30862 , \24970_25272 , \13755_14054 );
and \U$21759 ( \30561_30863 , \25516_25815 , \13390_13692 );
nor \U$21760 ( \30562_30864 , \30560_30862 , \30561_30863 );
xnor \U$21761 ( \30563_30865 , \30562_30864 , \13736_14035 );
xor \U$21762 ( \30564_30866 , \30559_30861 , \30563_30865 );
and \U$21763 ( \30565_30867 , \18730_19032 , \19235_19534 );
and \U$21764 ( \30566_30868 , \19259_19558 , \18743_19045 );
nor \U$21765 ( \30567_30869 , \30565_30867 , \30566_30868 );
xnor \U$21766 ( \30568_30870 , \30567_30869 , \19241_19540 );
xor \U$21767 ( \30569_30871 , \30564_30866 , \30568_30870 );
xor \U$21768 ( \30570_30872 , \30555_30857 , \30569_30871 );
xor \U$21769 ( \30571_30873 , \30546_30848 , \30570_30872 );
xor \U$21770 ( \30572_30874 , \30527_30829 , \30571_30873 );
and \U$21771 ( \30573_30875 , \29990_30292 , \29994_30296 );
and \U$21772 ( \30574_30876 , \29994_30296 , \30009_30311 );
and \U$21773 ( \30575_30877 , \29990_30292 , \30009_30311 );
or \U$21774 ( \30576_30878 , \30573_30875 , \30574_30876 , \30575_30877 );
and \U$21775 ( \30577_30879 , \30015_30317 , \30026_30328 );
and \U$21776 ( \30578_30880 , \30026_30328 , \30051_30353 );
and \U$21777 ( \30579_30881 , \30015_30317 , \30051_30353 );
or \U$21778 ( \30580_30882 , \30577_30879 , \30578_30880 , \30579_30881 );
xor \U$21779 ( \30581_30883 , \30576_30878 , \30580_30882 );
and \U$21780 ( \30582_30884 , \23315_23617 , \15037_15336 );
and \U$21781 ( \30583_30885 , \23900_24199 , \14661_14963 );
nor \U$21782 ( \30584_30886 , \30582_30884 , \30583_30885 );
xnor \U$21783 ( \30585_30887 , \30584_30886 , \15043_15342 );
and \U$21784 ( \30586_30888 , \17325_17627 , \20706_21005 );
and \U$21785 ( \30587_30889 , \17736_18035 , \20255_20557 );
nor \U$21786 ( \30588_30890 , \30586_30888 , \30587_30889 );
xnor \U$21787 ( \30589_30891 , \30588_30890 , \20712_21011 );
xor \U$21788 ( \30590_30892 , \30585_30887 , \30589_30891 );
and \U$21789 ( \30591_30893 , \15965_16267 , \22243_22542 );
and \U$21790 ( \30592_30894 , \16353_16655 , \21801_22103 );
nor \U$21791 ( \30593_30895 , \30591_30893 , \30592_30894 );
xnor \U$21792 ( \30594_30896 , \30593_30895 , \22249_22548 );
xor \U$21793 ( \30595_30897 , \30590_30892 , \30594_30896 );
and \U$21794 ( \30596_30898 , \26527_26829 , \12491_12790 );
and \U$21795 ( \30597_30899 , \27011_27313 , \12159_12461 );
nor \U$21796 ( \30598_30900 , \30596_30898 , \30597_30899 );
xnor \U$21797 ( \30599_30901 , \30598_30900 , \12481_12780 );
and \U$21798 ( \30600_30902 , \21788_22090 , \16333_16635 );
and \U$21799 ( \30601_30903 , \22257_22556 , \15999_16301 );
nor \U$21800 ( \30602_30904 , \30600_30902 , \30601_30903 );
xnor \U$21801 ( \30603_30905 , \30602_30904 , \16323_16625 );
xor \U$21802 ( \30604_30906 , \30599_30901 , \30603_30905 );
and \U$21803 ( \30605_30907 , \14648_14950 , \23839_24138 );
and \U$21804 ( \30606_30908 , \15022_15321 , \23328_23630 );
nor \U$21805 ( \30607_30909 , \30605_30907 , \30606_30908 );
xnor \U$21806 ( \30608_30910 , \30607_30909 , \23845_24144 );
xor \U$21807 ( \30609_30911 , \30604_30906 , \30608_30910 );
xor \U$21808 ( \30610_30912 , \30595_30897 , \30609_30911 );
and \U$21809 ( \30611_30913 , \20242_20544 , \17791_18090 );
and \U$21810 ( \30612_30914 , \20734_21033 , \17353_17655 );
nor \U$21811 ( \30613_30915 , \30611_30913 , \30612_30914 );
xnor \U$21812 ( \30614_30916 , \30613_30915 , \17747_18046 );
and \U$21813 ( \30615_30917 , \13377_13679 , \25527_25826 );
and \U$21814 ( \30616_30918 , \13725_14024 , \24962_25264 );
nor \U$21815 ( \30617_30919 , \30615_30917 , \30616_30918 );
xnor \U$21816 ( \30618_30920 , \30617_30919 , \25474_25773 );
xor \U$21817 ( \30619_30921 , \30614_30916 , \30618_30920 );
and \U$21818 ( \30620_30922 , \12146_12448 , \27095_27397 );
and \U$21819 ( \30621_30923 , \12470_12769 , \26505_26807 );
nor \U$21820 ( \30622_30924 , \30620_30922 , \30621_30923 );
xnor \U$21821 ( \30623_30925 , \30622_30924 , \26993_27295 );
xor \U$21822 ( \30624_30926 , \30619_30921 , \30623_30925 );
xor \U$21823 ( \30625_30927 , \30610_30912 , \30624_30926 );
xor \U$21824 ( \30626_30928 , \30581_30883 , \30625_30927 );
xor \U$21825 ( \30627_30929 , \30572_30874 , \30626_30928 );
xor \U$21826 ( \30628_30930 , \30224_30526 , \30627_30929 );
and \U$21827 ( \30629_30931 , \29659_29961 , \29981_30283 );
and \U$21828 ( \30630_30932 , \29981_30283 , \30053_30355 );
and \U$21829 ( \30631_30933 , \29659_29961 , \30053_30355 );
or \U$21830 ( \30632_30934 , \30629_30931 , \30630_30932 , \30631_30933 );
xor \U$21831 ( \30633_30935 , \30628_30930 , \30632_30934 );
and \U$21832 ( \30634_30936 , \30054_30356 , \30058_30360 );
and \U$21833 ( \30635_30937 , \30059_30361 , \30062_30364 );
or \U$21834 ( \30636_30938 , \30634_30936 , \30635_30937 );
xor \U$21835 ( \30637_30939 , \30633_30935 , \30636_30938 );
buf g9bb7_GF_PartitionCandidate( \30638_30940_nG9bb7 , \30637_30939 );
and \U$21836 ( \30639_30941 , \10402_10704 , \30638_30940_nG9bb7 );
or \U$21837 ( \30640_30942 , \30215_30517 , \30639_30941 );
xor \U$21838 ( \30641_30943 , \10399_10703 , \30640_30942 );
buf \U$21839 ( \30642_30944 , \30641_30943 );
buf \U$21841 ( \30643_30945 , \30642_30944 );
xor \U$21842 ( \30644_30946 , \30214_30516 , \30643_30945 );
buf \U$21843 ( \30645_30947 , \30644_30946 );
and \U$21844 ( \30646_30948 , \29647_29949 , \29653_29955 );
and \U$21845 ( \30647_30949 , \29647_29949 , \30069_30371 );
and \U$21846 ( \30648_30950 , \29653_29955 , \30069_30371 );
or \U$21847 ( \30649_30951 , \30646_30948 , \30647_30949 , \30648_30950 );
buf \U$21848 ( \30650_30952 , \30649_30951 );
xor \U$21849 ( \30651_30953 , \30645_30947 , \30650_30952 );
and \U$21850 ( \30652_30954 , \29614_29916 , \29620_29922 );
and \U$21851 ( \30653_30955 , \29614_29916 , \29627_29929 );
and \U$21852 ( \30654_30956 , \29620_29922 , \29627_29929 );
or \U$21853 ( \30655_30957 , \30652_30954 , \30653_30955 , \30654_30956 );
buf \U$21854 ( \30656_30958 , \30655_30957 );
and \U$21855 ( \30657_30959 , \29550_29849 , \29554_29856 );
buf \U$21856 ( \30658_30960 , \30657_30959 );
buf \U$21858 ( \30659_30961 , \30658_30960 );
and \U$21859 ( \30660_30962 , \28946_28118 , \10981_11283_nG9c08 );
and \U$21860 ( \30661_30963 , \27816_28115 , \11299_11598_nG9c05 );
or \U$21861 ( \30662_30964 , \30660_30962 , \30661_30963 );
xor \U$21862 ( \30663_30965 , \27815_28114 , \30662_30964 );
buf \U$21863 ( \30664_30966 , \30663_30965 );
buf \U$21865 ( \30665_30967 , \30664_30966 );
xor \U$21866 ( \30666_30968 , \30659_30961 , \30665_30967 );
buf \U$21867 ( \30667_30969 , \30666_30968 );
not \U$20741 ( \30668_29851 , \29551_29850 );
xor \U$20742 ( \30669_29852 , \29545_29844_nG4400 , \29548_29847_nG4403 );
and \U$20743 ( \30670_29853 , \30668_29851 , \30669_29852 );
and \U$21868 ( \30671_30970 , \30670_29853 , \10392_10694_nG9c0e );
and \U$21869 ( \30672_30971 , \29551_29850 , \10693_10995_nG9c0b );
or \U$21870 ( \30673_30972 , \30671_30970 , \30672_30971 );
xor \U$21871 ( \30674_30973 , \29550_29849 , \30673_30972 );
buf \U$21872 ( \30675_30974 , \30674_30973 );
buf \U$21874 ( \30676_30975 , \30675_30974 );
xor \U$21875 ( \30677_30976 , \30667_30969 , \30676_30975 );
and \U$21876 ( \30678_30977 , \27141_26431 , \12168_12470_nG9c02 );
and \U$21877 ( \30679_30978 , \26129_26428 , \12502_12801_nG9bff );
or \U$21878 ( \30680_30979 , \30678_30977 , \30679_30978 );
xor \U$21879 ( \30681_30980 , \26128_26427 , \30680_30979 );
buf \U$21880 ( \30682_30981 , \30681_30980 );
buf \U$21882 ( \30683_30982 , \30682_30981 );
xor \U$21883 ( \30684_30983 , \30677_30976 , \30683_30982 );
buf \U$21884 ( \30685_30984 , \30684_30983 );
xor \U$21885 ( \30686_30985 , \30656_30958 , \30685_30984 );
and \U$21886 ( \30687_30986 , \21908_21658 , \16013_16315_nG9bf0 );
and \U$21887 ( \30688_30987 , \21356_21655 , \16378_16680_nG9bed );
or \U$21888 ( \30689_30988 , \30687_30986 , \30688_30987 );
xor \U$21889 ( \30690_30989 , \21355_21654 , \30689_30988 );
buf \U$21890 ( \30691_30990 , \30690_30989 );
buf \U$21892 ( \30692_30991 , \30691_30990 );
xor \U$21893 ( \30693_30992 , \30686_30985 , \30692_30991 );
buf \U$21894 ( \30694_30993 , \30693_30992 );
and \U$21895 ( \30695_30994 , \18908_18702 , \18789_19091_nG9be4 );
and \U$21896 ( \30696_30995 , \18400_18699 , \19287_19586_nG9be1 );
or \U$21897 ( \30697_30996 , \30695_30994 , \30696_30995 );
xor \U$21898 ( \30698_30997 , \18399_18698 , \30697_30996 );
buf \U$21899 ( \30699_30998 , \30698_30997 );
buf \U$21901 ( \30700_30999 , \30699_30998 );
xor \U$21902 ( \30701_31000 , \30694_30993 , \30700_30999 );
and \U$21903 ( \30702_31001 , \17437_17297 , \20306_20608_nG9bde );
and \U$21904 ( \30703_31002 , \16995_17294 , \20787_21086_nG9bdb );
or \U$21905 ( \30704_31003 , \30702_31001 , \30703_31002 );
xor \U$21906 ( \30705_31004 , \16994_17293 , \30704_31003 );
buf \U$21907 ( \30706_31005 , \30705_31004 );
buf \U$21909 ( \30707_31006 , \30706_31005 );
xor \U$21910 ( \30708_31007 , \30701_31000 , \30707_31006 );
buf \U$21911 ( \30709_31008 , \30708_31007 );
and \U$21912 ( \30710_31009 , \13431_13370 , \24996_25298_nG9bcc );
and \U$21913 ( \30711_31010 , \13068_13367 , \25561_25860_nG9bc9 );
or \U$21914 ( \30712_31011 , \30710_31009 , \30711_31010 );
xor \U$21915 ( \30713_31012 , \13067_13366 , \30712_31011 );
buf \U$21916 ( \30714_31013 , \30713_31012 );
buf \U$21918 ( \30715_31014 , \30714_31013 );
xor \U$21919 ( \30716_31015 , \30709_31008 , \30715_31014 );
and \U$21920 ( \30717_31016 , \10996_10421 , \28300_28602_nG9bc0 );
and \U$21921 ( \30718_31017 , \10119_10418 , \28877_29179_nG9bbd );
or \U$21922 ( \30719_31018 , \30717_31016 , \30718_31017 );
xor \U$21923 ( \30720_31019 , \10118_10417 , \30719_31018 );
buf \U$21924 ( \30721_31020 , \30720_31019 );
buf \U$21926 ( \30722_31021 , \30721_31020 );
xor \U$21927 ( \30723_31022 , \30716_31015 , \30722_31021 );
buf \U$21928 ( \30724_31023 , \30723_31022 );
xor \U$21929 ( \30725_31024 , \30651_30953 , \30724_31023 );
buf \U$21930 ( \30726_31025 , \30725_31024 );
and \U$21931 ( \30727_31026 , \29568_29870 , \29601_29903 );
and \U$21932 ( \30728_31027 , \29568_29870 , \30071_30373 );
and \U$21933 ( \30729_31028 , \29601_29903 , \30071_30373 );
or \U$21934 ( \30730_31029 , \30727_31026 , \30728_31027 , \30729_31028 );
buf \U$21935 ( \30731_31030 , \30730_31029 );
xor \U$21936 ( \30732_31031 , \30726_31025 , \30731_31030 );
and \U$21937 ( \30733_31032 , \30117_30419 , \30123_30425 );
and \U$21938 ( \30734_31033 , \30117_30419 , \30130_30432 );
and \U$21939 ( \30735_31034 , \30123_30425 , \30130_30432 );
or \U$21940 ( \30736_31035 , \30733_31032 , \30734_31033 , \30735_31034 );
buf \U$21941 ( \30737_31036 , \30736_31035 );
and \U$21942 ( \30738_31037 , \14710_14631 , \23394_23696_nG9bd2 );
and \U$21943 ( \30739_31038 , \14329_14628 , \23927_24226_nG9bcf );
or \U$21944 ( \30740_31039 , \30738_31037 , \30739_31038 );
xor \U$21945 ( \30741_31040 , \14328_14627 , \30740_31039 );
buf \U$21946 ( \30742_31041 , \30741_31040 );
buf \U$21948 ( \30743_31042 , \30742_31041 );
xor \U$21949 ( \30744_31043 , \30737_31036 , \30743_31042 );
and \U$21950 ( \30745_31044 , \12183_12157 , \26585_26887_nG9bc6 );
and \U$21951 ( \30746_31045 , \11855_12154 , \27114_27416_nG9bc3 );
or \U$21952 ( \30747_31046 , \30745_31044 , \30746_31045 );
xor \U$21953 ( \30748_31047 , \11854_12153 , \30747_31046 );
buf \U$21954 ( \30749_31048 , \30748_31047 );
buf \U$21956 ( \30750_31049 , \30749_31048 );
xor \U$21957 ( \30751_31050 , \30744_31043 , \30750_31049 );
buf \U$21958 ( \30752_31051 , \30751_31050 );
and \U$21959 ( \30753_31052 , \30089_30391 , \30132_30434 );
and \U$21960 ( \30754_31053 , \30089_30391 , \30139_30441 );
and \U$21961 ( \30755_31054 , \30132_30434 , \30139_30441 );
or \U$21962 ( \30756_31055 , \30753_31052 , \30754_31053 , \30755_31054 );
buf \U$21963 ( \30757_31056 , \30756_31055 );
xor \U$21964 ( \30758_31057 , \30752_31051 , \30757_31056 );
and \U$21965 ( \30759_31058 , \29578_29880 , \29584_29886 );
and \U$21966 ( \30760_31059 , \29578_29880 , \29591_29893 );
and \U$21967 ( \30761_31060 , \29584_29886 , \29591_29893 );
or \U$21968 ( \30762_31061 , \30759_31058 , \30760_31059 , \30761_31060 );
buf \U$21969 ( \30763_31062 , \30762_31061 );
xor \U$21970 ( \30764_31063 , \30758_31057 , \30763_31062 );
buf \U$21971 ( \30765_31064 , \30764_31063 );
and \U$21972 ( \30766_31065 , \30084_30386 , \30141_30443 );
and \U$21973 ( \30767_31066 , \30084_30386 , \30147_30449 );
and \U$21974 ( \30768_31067 , \30141_30443 , \30147_30449 );
or \U$21975 ( \30769_31068 , \30766_31065 , \30767_31066 , \30768_31067 );
buf \U$21976 ( \30770_31069 , \30769_31068 );
xor \U$21977 ( \30771_31070 , \30765_31064 , \30770_31069 );
and \U$21978 ( \30772_31071 , \29573_29875 , \29593_29895 );
and \U$21979 ( \30773_31072 , \29573_29875 , \29599_29901 );
and \U$21980 ( \30774_31073 , \29593_29895 , \29599_29901 );
or \U$21981 ( \30775_31074 , \30772_31071 , \30773_31072 , \30774_31073 );
buf \U$21982 ( \30776_31075 , \30775_31074 );
xor \U$21983 ( \30777_31076 , \30771_31070 , \30776_31075 );
buf \U$21984 ( \30778_31077 , \30777_31076 );
xor \U$21985 ( \30779_31078 , \30732_31031 , \30778_31077 );
and \U$21986 ( \30780_31079 , \30163_30465 , \30779_31078 );
and \U$21987 ( \30781_31080 , \30153_30455 , \30157_30459 );
and \U$21988 ( \30782_31081 , \30153_30455 , \30162_30464 );
and \U$21989 ( \30783_31082 , \30157_30459 , \30162_30464 );
or \U$21990 ( \30784_31083 , \30781_31080 , \30782_31081 , \30783_31082 );
xor \U$21991 ( \30785_31084 , \30780_31079 , \30784_31083 );
and \U$21992 ( \30786_31085 , RIdec6350_719, \8760_9059 );
and \U$21993 ( \30787_31086 , RIdec3650_687, \8762_9061 );
and \U$21994 ( \30788_31087 , RIfcaf3d0_7016, \8764_9063 );
and \U$21995 ( \30789_31088 , RIdec0950_655, \8766_9065 );
and \U$21996 ( \30790_31089 , RIfc6a280_6230, \8768_9067 );
and \U$21997 ( \30791_31090 , RIdebdc50_623, \8770_9069 );
and \U$21998 ( \30792_31091 , RIdebaf50_591, \8772_9071 );
and \U$21999 ( \30793_31092 , RIdeb8250_559, \8774_9073 );
and \U$22000 ( \30794_31093 , RIfc42f50_5784, \8776_9075 );
and \U$22001 ( \30795_31094 , RIdeb2850_495, \8778_9077 );
and \U$22002 ( \30796_31095 , RIfc981f8_6753, \8780_9079 );
and \U$22003 ( \30797_31096 , RIdeafb50_463, \8782_9081 );
and \U$22004 ( \30798_31097 , RIfc8c6f0_6620, \8784_9083 );
and \U$22005 ( \30799_31098 , RIdeac838_431, \8786_9085 );
and \U$22006 ( \30800_31099 , RIdea5f38_399, \8788_9087 );
and \U$22007 ( \30801_31100 , RIde9f638_367, \8790_9089 );
and \U$22008 ( \30802_31101 , RIee1d4e8_4792, \8792_9091 );
and \U$22009 ( \30803_31102 , RIfcda648_7507, \8794_9093 );
and \U$22010 ( \30804_31103 , RIfcc6440_7278, \8796_9095 );
and \U$22011 ( \30805_31104 , RIfcd5620_7450, \8798_9097 );
and \U$22012 ( \30806_31105 , RIde92ac8_305, \8800_9099 );
and \U$22013 ( \30807_31106 , RIfea34a0_8202, \8802_9101 );
and \U$22014 ( \30808_31107 , RIfea31d0_8200, \8804_9103 );
and \U$22015 ( \30809_31108 , RIfea3338_8201, \8806_9105 );
and \U$22016 ( \30810_31109 , RIfcb6b58_7101, \8808_9107 );
and \U$22017 ( \30811_31110 , RIfcb6888_7099, \8810_9109 );
and \U$22018 ( \30812_31111 , RIfc9dd60_6818, \8812_9111 );
and \U$22019 ( \30813_31112 , RIee19708_4748, \8814_9113 );
and \U$22020 ( \30814_31113 , RIfc50c18_5941, \8816_9115 );
and \U$22021 ( \30815_31114 , RIe16c458_2609, \8818_9117 );
and \U$22022 ( \30816_31115 , RIfc80a80_6486, \8820_9119 );
and \U$22023 ( \30817_31116 , RIfec62e8_8375, \8822_9121 );
and \U$22024 ( \30818_31117 , RIe166350_2540, \8824_9123 );
and \U$22025 ( \30819_31118 , RIe163650_2508, \8826_9125 );
and \U$22026 ( \30820_31119 , RIee37d98_5094, \8828_9127 );
and \U$22027 ( \30821_31120 , RIe160950_2476, \8830_9129 );
and \U$22028 ( \30822_31121 , RIfcaa678_6961, \8832_9131 );
and \U$22029 ( \30823_31122 , RIe15dc50_2444, \8834_9133 );
and \U$22030 ( \30824_31123 , RIe158250_2380, \8836_9135 );
and \U$22031 ( \30825_31124 , RIe155550_2348, \8838_9137 );
and \U$22032 ( \30826_31125 , RIfea3ba8_8207, \8840_9139 );
and \U$22033 ( \30827_31126 , RIe152850_2316, \8842_9141 );
and \U$22034 ( \30828_31127 , RIee35638_5066, \8844_9143 );
and \U$22035 ( \30829_31128 , RIe14fb50_2284, \8846_9145 );
and \U$22036 ( \30830_31129 , RIfc62f30_6148, \8848_9147 );
and \U$22037 ( \30831_31130 , RIe14ce50_2252, \8850_9149 );
and \U$22038 ( \30832_31131 , RIe14a150_2220, \8852_9151 );
and \U$22039 ( \30833_31132 , RIe147450_2188, \8854_9153 );
and \U$22040 ( \30834_31133 , RIfc97f28_6751, \8856_9155 );
and \U$22041 ( \30835_31134 , RIfc89888_6587, \8858_9157 );
and \U$22042 ( \30836_31135 , RIfc8f558_6653, \8860_9159 );
and \U$22043 ( \30837_31136 , RIfc52838_5961, \8862_9161 );
and \U$22044 ( \30838_31137 , RIe141bb8_2125, \8864_9163 );
and \U$22045 ( \30839_31138 , RIe13f890_2100, \8866_9165 );
and \U$22046 ( \30840_31139 , RIdf3d798_2076, \8868_9167 );
and \U$22047 ( \30841_31140 , RIdf3b308_2050, \8870_9169 );
and \U$22048 ( \30842_31141 , RIee30a48_5012, \8872_9171 );
and \U$22049 ( \30843_31142 , RIfc568e8_6007, \8874_9173 );
and \U$22050 ( \30844_31143 , RIee2e9f0_4989, \8876_9175 );
and \U$22051 ( \30845_31144 , RIee2dbe0_4979, \8878_9177 );
and \U$22052 ( \30846_31145 , RIdf365b0_1995, \8880_9179 );
and \U$22053 ( \30847_31146 , RIfea38d8_8205, \8882_9181 );
and \U$22054 ( \30848_31147 , RIfea3a40_8206, \8884_9183 );
and \U$22055 ( \30849_31148 , RIdf2ff08_1922, \8886_9185 );
or \U$22056 ( \30850_31149 , \30786_31085 , \30787_31086 , \30788_31087 , \30789_31088 , \30790_31089 , \30791_31090 , \30792_31091 , \30793_31092 , \30794_31093 , \30795_31094 , \30796_31095 , \30797_31096 , \30798_31097 , \30799_31098 , \30800_31099 , \30801_31100 , \30802_31101 , \30803_31102 , \30804_31103 , \30805_31104 , \30806_31105 , \30807_31106 , \30808_31107 , \30809_31108 , \30810_31109 , \30811_31110 , \30812_31111 , \30813_31112 , \30814_31113 , \30815_31114 , \30816_31115 , \30817_31116 , \30818_31117 , \30819_31118 , \30820_31119 , \30821_31120 , \30822_31121 , \30823_31122 , \30824_31123 , \30825_31124 , \30826_31125 , \30827_31126 , \30828_31127 , \30829_31128 , \30830_31129 , \30831_31130 , \30832_31131 , \30833_31132 , \30834_31133 , \30835_31134 , \30836_31135 , \30837_31136 , \30838_31137 , \30839_31138 , \30840_31139 , \30841_31140 , \30842_31141 , \30843_31142 , \30844_31143 , \30845_31144 , \30846_31145 , \30847_31146 , \30848_31147 , \30849_31148 );
and \U$22057 ( \30851_31150 , RIee2c6c8_4964, \8889_9188 );
and \U$22058 ( \30852_31151 , RIee2ac10_4945, \8891_9190 );
and \U$22059 ( \30853_31152 , RIee29590_4929, \8893_9192 );
and \U$22060 ( \30854_31153 , RIee28348_4916, \8895_9194 );
and \U$22061 ( \30855_31154 , RIdf2ad78_1864, \8897_9196 );
and \U$22062 ( \30856_31155 , RIdf28e88_1842, \8899_9198 );
and \U$22063 ( \30857_31156 , RIfea3608_8203, \8901_9200 );
and \U$22064 ( \30858_31157 , RIfea3770_8204, \8903_9202 );
and \U$22065 ( \30859_31158 , RIfcc0d10_7216, \8905_9204 );
and \U$22066 ( \30860_31159 , RIfc75c20_6362, \8907_9206 );
and \U$22067 ( \30861_31160 , RIfca50b0_6900, \8909_9208 );
and \U$22068 ( \30862_31161 , RIfc74e10_6352, \8911_9210 );
and \U$22069 ( \30863_31162 , RIfcc9410_7312, \8913_9212 );
and \U$22070 ( \30864_31163 , RIdf20620_1745, \8915_9214 );
and \U$22071 ( \30865_31164 , RIfc73628_6335, \8917_9216 );
and \U$22072 ( \30866_31165 , RIdf1a0e0_1673, \8919_9218 );
and \U$22073 ( \30867_31166 , RIdf17f20_1649, \8921_9220 );
and \U$22074 ( \30868_31167 , RIdf15220_1617, \8923_9222 );
and \U$22075 ( \30869_31168 , RIdf12520_1585, \8925_9224 );
and \U$22076 ( \30870_31169 , RIdf0f820_1553, \8927_9226 );
and \U$22077 ( \30871_31170 , RIdf0cb20_1521, \8929_9228 );
and \U$22078 ( \30872_31171 , RIdf09e20_1489, \8931_9230 );
and \U$22079 ( \30873_31172 , RIdf07120_1457, \8933_9232 );
and \U$22080 ( \30874_31173 , RIdf04420_1425, \8935_9234 );
and \U$22081 ( \30875_31174 , RIdefea20_1361, \8937_9236 );
and \U$22082 ( \30876_31175 , RIdefbd20_1329, \8939_9238 );
and \U$22083 ( \30877_31176 , RIdef9020_1297, \8941_9240 );
and \U$22084 ( \30878_31177 , RIdef6320_1265, \8943_9242 );
and \U$22085 ( \30879_31178 , RIdef3620_1233, \8945_9244 );
and \U$22086 ( \30880_31179 , RIdef0920_1201, \8947_9246 );
and \U$22087 ( \30881_31180 , RIdeedc20_1169, \8949_9248 );
and \U$22088 ( \30882_31181 , RIdeeaf20_1137, \8951_9250 );
and \U$22089 ( \30883_31182 , RIfcab8c0_6974, \8953_9252 );
and \U$22090 ( \30884_31183 , RIfc7c598_6437, \8955_9254 );
and \U$22091 ( \30885_31184 , RIfc5beb0_6068, \8957_9256 );
and \U$22092 ( \30886_31185 , RIfc58ee0_6034, \8959_9258 );
and \U$22093 ( \30887_31186 , RIdee5688_1074, \8961_9260 );
and \U$22094 ( \30888_31187 , RIdee3798_1052, \8963_9262 );
and \U$22095 ( \30889_31188 , RIdee15d8_1028, \8965_9264 );
and \U$22096 ( \30890_31189 , RIdedf580_1005, \8967_9266 );
and \U$22097 ( \30891_31190 , RIfcb3048_7059, \8969_9268 );
and \U$22098 ( \30892_31191 , RIfc72ae8_6327, \8971_9270 );
and \U$22099 ( \30893_31192 , RIfca3d00_6886, \8973_9272 );
and \U$22100 ( \30894_31193 , RIfcb6450_7096, \8975_9274 );
and \U$22101 ( \30895_31194 , RIdeda558_948, \8977_9276 );
and \U$22102 ( \30896_31195 , RIded7f60_921, \8979_9278 );
and \U$22103 ( \30897_31196 , RIfea3068_8199, \8981_9280 );
and \U$22104 ( \30898_31197 , RIded3a78_872, \8983_9282 );
and \U$22105 ( \30899_31198 , RIded1750_847, \8985_9284 );
and \U$22106 ( \30900_31199 , RIdecea50_815, \8987_9286 );
and \U$22107 ( \30901_31200 , RIdecbd50_783, \8989_9288 );
and \U$22108 ( \30902_31201 , RIdec9050_751, \8991_9290 );
and \U$22109 ( \30903_31202 , RIdeb5550_527, \8993_9292 );
and \U$22110 ( \30904_31203 , RIde98d38_335, \8995_9294 );
and \U$22111 ( \30905_31204 , RIe16f158_2641, \8997_9296 );
and \U$22112 ( \30906_31205 , RIe15af50_2412, \8999_9298 );
and \U$22113 ( \30907_31206 , RIe144750_2156, \9001_9300 );
and \U$22114 ( \30908_31207 , RIdf39148_2026, \9003_9302 );
and \U$22115 ( \30909_31208 , RIdf2d7a8_1894, \9005_9304 );
and \U$22116 ( \30910_31209 , RIdf1e028_1718, \9007_9306 );
and \U$22117 ( \30911_31210 , RIdf01720_1393, \9009_9308 );
and \U$22118 ( \30912_31211 , RIdee8220_1105, \9011_9310 );
and \U$22119 ( \30913_31212 , RIdedcf88_978, \9013_9312 );
and \U$22120 ( \30914_31213 , RIde7ec80_208, \9015_9314 );
or \U$22121 ( \30915_31214 , \30851_31150 , \30852_31151 , \30853_31152 , \30854_31153 , \30855_31154 , \30856_31155 , \30857_31156 , \30858_31157 , \30859_31158 , \30860_31159 , \30861_31160 , \30862_31161 , \30863_31162 , \30864_31163 , \30865_31164 , \30866_31165 , \30867_31166 , \30868_31167 , \30869_31168 , \30870_31169 , \30871_31170 , \30872_31171 , \30873_31172 , \30874_31173 , \30875_31174 , \30876_31175 , \30877_31176 , \30878_31177 , \30879_31178 , \30880_31179 , \30881_31180 , \30882_31181 , \30883_31182 , \30884_31183 , \30885_31184 , \30886_31185 , \30887_31186 , \30888_31187 , \30889_31188 , \30890_31189 , \30891_31190 , \30892_31191 , \30893_31192 , \30894_31193 , \30895_31194 , \30896_31195 , \30897_31196 , \30898_31197 , \30899_31198 , \30900_31199 , \30901_31200 , \30902_31201 , \30903_31202 , \30904_31203 , \30905_31204 , \30906_31205 , \30907_31206 , \30908_31207 , \30909_31208 , \30910_31209 , \30911_31210 , \30912_31211 , \30913_31212 , \30914_31213 );
or \U$22122 ( \30916_31215 , \30850_31149 , \30915_31214 );
_DC \g2235/U$1 ( \30917 , \30916_31215 , \9024_9323 );
buf \U$22123 ( \30918_31217 , \30917 );
and \U$22124 ( \30919_31218 , RIe19e5e8_3179, \9034_9333 );
and \U$22125 ( \30920_31219 , RIe19b8e8_3147, \9036_9335 );
and \U$22126 ( \30921_31220 , RIfca84b8_6937, \9038_9337 );
and \U$22127 ( \30922_31221 , RIe198be8_3115, \9040_9339 );
and \U$22128 ( \30923_31222 , RIfc846f8_6529, \9042_9341 );
and \U$22129 ( \30924_31223 , RIe195ee8_3083, \9044_9343 );
and \U$22130 ( \30925_31224 , RIe1931e8_3051, \9046_9345 );
and \U$22131 ( \30926_31225 , RIe1904e8_3019, \9048_9347 );
and \U$22132 ( \30927_31226 , RIe18aae8_2955, \9050_9349 );
and \U$22133 ( \30928_31227 , RIe187de8_2923, \9052_9351 );
and \U$22134 ( \30929_31228 , RIfce2be0_7602, \9054_9353 );
and \U$22135 ( \30930_31229 , RIe1850e8_2891, \9056_9355 );
and \U$22136 ( \30931_31230 , RIfc8e310_6640, \9058_9357 );
and \U$22137 ( \30932_31231 , RIe1823e8_2859, \9060_9359 );
and \U$22138 ( \30933_31232 , RIe17f6e8_2827, \9062_9361 );
and \U$22139 ( \30934_31233 , RIe17c9e8_2795, \9064_9363 );
and \U$22140 ( \30935_31234 , RIfcd1570_7404, \9066_9365 );
and \U$22141 ( \30936_31235 , RIfccc278_7345, \9068_9367 );
and \U$22142 ( \30937_31236 , RIf1404c8_5191, \9070_9369 );
and \U$22143 ( \30938_31237 , RIfea2d98_8197, \9072_9371 );
and \U$22144 ( \30939_31238 , RIfcc1b20_7226, \9074_9373 );
and \U$22145 ( \30940_31239 , RIfc60398_6117, \9076_9375 );
and \U$22146 ( \30941_31240 , RIee3e5a8_5168, \9078_9377 );
and \U$22147 ( \30942_31241 , RIee3da68_5160, \9080_9379 );
and \U$22148 ( \30943_31242 , RIfc642e0_6162, \9082_9381 );
and \U$22149 ( \30944_31243 , RIfca7f18_6933, \9084_9383 );
and \U$22150 ( \30945_31244 , RIee3a228_5120, \9086_9385 );
and \U$22151 ( \30946_31245 , RIfec6180_8374, \9088_9387 );
and \U$22152 ( \30947_31246 , RIfca9598_6949, \9090_9389 );
and \U$22153 ( \30948_31247 , RIfc5c720_6074, \9092_9391 );
and \U$22154 ( \30949_31248 , RIfc6bea0_6250, \9094_9393 );
and \U$22155 ( \30950_31249 , RIfccaec8_7331, \9096_9395 );
and \U$22156 ( \30951_31250 , RIfc44cd8_5805, \9098_9397 );
and \U$22157 ( \30952_31251 , RIe224940_4706, \9100_9399 );
and \U$22158 ( \30953_31252 , RIfcb6180_7094, \9102_9401 );
and \U$22159 ( \30954_31253 , RIe221c40_4674, \9104_9403 );
and \U$22160 ( \30955_31254 , RIfc55ad8_5997, \9106_9405 );
and \U$22161 ( \30956_31255 , RIe21ef40_4642, \9108_9407 );
and \U$22162 ( \30957_31256 , RIe219540_4578, \9110_9409 );
and \U$22163 ( \30958_31257 , RIe216840_4546, \9112_9411 );
and \U$22164 ( \30959_31258 , RIfc4dc48_5907, \9114_9413 );
and \U$22165 ( \30960_31259 , RIe213b40_4514, \9116_9415 );
and \U$22166 ( \30961_31260 , RIfcdcf10_7536, \9118_9417 );
and \U$22167 ( \30962_31261 , RIe210e40_4482, \9120_9419 );
and \U$22168 ( \30963_31262 , RIfcab1b8_6969, \9122_9421 );
and \U$22169 ( \30964_31263 , RIe20e140_4450, \9124_9423 );
and \U$22170 ( \30965_31264 , RIe20b440_4418, \9126_9425 );
and \U$22171 ( \30966_31265 , RIe208740_4386, \9128_9427 );
and \U$22172 ( \30967_31266 , RIfce3720_7610, \9130_9429 );
and \U$22173 ( \30968_31267 , RIfc64178_6161, \9132_9431 );
and \U$22174 ( \30969_31268 , RIe203178_4325, \9134_9433 );
and \U$22175 ( \30970_31269 , RIe201558_4305, \9136_9435 );
and \U$22176 ( \30971_31270 , RIfcd2ec0_7422, \9138_9437 );
and \U$22177 ( \30972_31271 , RIf164828_5603, \9140_9439 );
and \U$22178 ( \30973_31272 , RIfc7f838_6473, \9142_9441 );
and \U$22179 ( \30974_31273 , RIf162398_5577, \9144_9443 );
and \U$22180 ( \30975_31274 , RIfcc9c80_7318, \9146_9445 );
and \U$22181 ( \30976_31275 , RIfca8bc0_6942, \9148_9447 );
and \U$22182 ( \30977_31276 , RIfea2ac8_8195, \9150_9449 );
and \U$22183 ( \30978_31277 , RIfea2c30_8196, \9152_9451 );
and \U$22184 ( \30979_31278 , RIfc59318_6037, \9154_9453 );
and \U$22185 ( \30980_31279 , RIfc4f160_5922, \9156_9455 );
and \U$22186 ( \30981_31280 , RIf15ac10_5492, \9158_9457 );
and \U$22187 ( \30982_31281 , RIfcebf88_7707, \9160_9459 );
or \U$22188 ( \30983_31282 , \30919_31218 , \30920_31219 , \30921_31220 , \30922_31221 , \30923_31222 , \30924_31223 , \30925_31224 , \30926_31225 , \30927_31226 , \30928_31227 , \30929_31228 , \30930_31229 , \30931_31230 , \30932_31231 , \30933_31232 , \30934_31233 , \30935_31234 , \30936_31235 , \30937_31236 , \30938_31237 , \30939_31238 , \30940_31239 , \30941_31240 , \30942_31241 , \30943_31242 , \30944_31243 , \30945_31244 , \30946_31245 , \30947_31246 , \30948_31247 , \30949_31248 , \30950_31249 , \30951_31250 , \30952_31251 , \30953_31252 , \30954_31253 , \30955_31254 , \30956_31255 , \30957_31256 , \30958_31257 , \30959_31258 , \30960_31259 , \30961_31260 , \30962_31261 , \30963_31262 , \30964_31263 , \30965_31264 , \30966_31265 , \30967_31266 , \30968_31267 , \30969_31268 , \30970_31269 , \30971_31270 , \30972_31271 , \30973_31272 , \30974_31273 , \30975_31274 , \30976_31275 , \30977_31276 , \30978_31277 , \30979_31278 , \30980_31279 , \30981_31280 , \30982_31281 );
and \U$22189 ( \30984_31283 , RIfcbb040_7150, \9163_9462 );
and \U$22190 ( \30985_31284 , RIfca1870_6860, \9165_9464 );
and \U$22191 ( \30986_31285 , RIfc93d10_6704, \9167_9466 );
and \U$22192 ( \30987_31286 , RIe1faeb0_4232, \9169_9468 );
and \U$22193 ( \30988_31287 , RIf1565c0_5442, \9171_9470 );
and \U$22194 ( \30989_31288 , RIf155a80_5434, \9173_9472 );
and \U$22195 ( \30990_31289 , RIfc45c50_5816, \9175_9474 );
and \U$22196 ( \30991_31290 , RIe1f6428_4179, \9177_9476 );
and \U$22197 ( \30992_31291 , RIfccdbc8_7363, \9179_9478 );
and \U$22198 ( \30993_31292 , RIfcccae8_7351, \9181_9480 );
and \U$22199 ( \30994_31293 , RIfca6cd0_6920, \9183_9482 );
and \U$22200 ( \30995_31294 , RIfec6018_8373, \9185_9484 );
and \U$22201 ( \30996_31295 , RIfc64010_6160, \9187_9486 );
and \U$22202 ( \30997_31296 , RIfc434f0_5788, \9189_9488 );
and \U$22203 ( \30998_31297 , RIfc4c028_5887, \9191_9490 );
and \U$22204 ( \30999_31298 , RIe1eee08_4095, \9193_9492 );
and \U$22205 ( \31000_31299 , RIe1ec6a8_4067, \9195_9494 );
and \U$22206 ( \31001_31300 , RIe1e99a8_4035, \9197_9496 );
and \U$22207 ( \31002_31301 , RIe1e6ca8_4003, \9199_9498 );
and \U$22208 ( \31003_31302 , RIe1e3fa8_3971, \9201_9500 );
and \U$22209 ( \31004_31303 , RIe1e12a8_3939, \9203_9502 );
and \U$22210 ( \31005_31304 , RIe1de5a8_3907, \9205_9504 );
and \U$22211 ( \31006_31305 , RIe1db8a8_3875, \9207_9506 );
and \U$22212 ( \31007_31306 , RIe1d8ba8_3843, \9209_9508 );
and \U$22213 ( \31008_31307 , RIe1d31a8_3779, \9211_9510 );
and \U$22214 ( \31009_31308 , RIe1d04a8_3747, \9213_9512 );
and \U$22215 ( \31010_31309 , RIe1cd7a8_3715, \9215_9514 );
and \U$22216 ( \31011_31310 , RIe1caaa8_3683, \9217_9516 );
and \U$22217 ( \31012_31311 , RIe1c7da8_3651, \9219_9518 );
and \U$22218 ( \31013_31312 , RIe1c50a8_3619, \9221_9520 );
and \U$22219 ( \31014_31313 , RIe1c23a8_3587, \9223_9522 );
and \U$22220 ( \31015_31314 , RIe1bf6a8_3555, \9225_9524 );
and \U$22221 ( \31016_31315 , RIfc63908_6155, \9227_9526 );
and \U$22222 ( \31017_31316 , RIfc6bd38_6249, \9229_9528 );
and \U$22223 ( \31018_31317 , RIe1ba0e0_3494, \9231_9530 );
and \U$22224 ( \31019_31318 , RIe1b7f20_3470, \9233_9532 );
and \U$22225 ( \31020_31319 , RIfc66fe0_6194, \9235_9534 );
and \U$22226 ( \31021_31320 , RIfc92ac8_6691, \9237_9536 );
and \U$22227 ( \31022_31321 , RIe1b5d60_3446, \9239_9538 );
and \U$22228 ( \31023_31322 , RIfea2f00_8198, \9241_9540 );
and \U$22229 ( \31024_31323 , RIfc9bfd8_6797, \9243_9542 );
and \U$22230 ( \31025_31324 , RIfc50d80_5942, \9245_9544 );
and \U$22231 ( \31026_31325 , RIe1b31c8_3415, \9247_9546 );
and \U$22232 ( \31027_31326 , RIe1b1878_3397, \9249_9548 );
and \U$22233 ( \31028_31327 , RIfc4df18_5909, \9251_9550 );
and \U$22234 ( \31029_31328 , RIfc9d658_6813, \9253_9552 );
and \U$22235 ( \31030_31329 , RIe1ad0c0_3346, \9255_9554 );
and \U$22236 ( \31031_31330 , RIe1ab8d8_3329, \9257_9556 );
and \U$22237 ( \31032_31331 , RIe1a99e8_3307, \9259_9558 );
and \U$22238 ( \31033_31332 , RIe1a6ce8_3275, \9261_9560 );
and \U$22239 ( \31034_31333 , RIe1a3fe8_3243, \9263_9562 );
and \U$22240 ( \31035_31334 , RIe1a12e8_3211, \9265_9564 );
and \U$22241 ( \31036_31335 , RIe18d7e8_2987, \9267_9566 );
and \U$22242 ( \31037_31336 , RIe179ce8_2763, \9269_9568 );
and \U$22243 ( \31038_31337 , RIe227640_4738, \9271_9570 );
and \U$22244 ( \31039_31338 , RIe21c240_4610, \9273_9572 );
and \U$22245 ( \31040_31339 , RIe205a40_4354, \9275_9574 );
and \U$22246 ( \31041_31340 , RIe1ffaa0_4286, \9277_9576 );
and \U$22247 ( \31042_31341 , RIe1f8e58_4209, \9279_9578 );
and \U$22248 ( \31043_31342 , RIe1f19a0_4126, \9281_9580 );
and \U$22249 ( \31044_31343 , RIe1d5ea8_3811, \9283_9582 );
and \U$22250 ( \31045_31344 , RIe1bc9a8_3523, \9285_9584 );
and \U$22251 ( \31046_31345 , RIe1af820_3374, \9287_9586 );
and \U$22252 ( \31047_31346 , RIe171e58_2673, \9289_9588 );
or \U$22253 ( \31048_31347 , \30984_31283 , \30985_31284 , \30986_31285 , \30987_31286 , \30988_31287 , \30989_31288 , \30990_31289 , \30991_31290 , \30992_31291 , \30993_31292 , \30994_31293 , \30995_31294 , \30996_31295 , \30997_31296 , \30998_31297 , \30999_31298 , \31000_31299 , \31001_31300 , \31002_31301 , \31003_31302 , \31004_31303 , \31005_31304 , \31006_31305 , \31007_31306 , \31008_31307 , \31009_31308 , \31010_31309 , \31011_31310 , \31012_31311 , \31013_31312 , \31014_31313 , \31015_31314 , \31016_31315 , \31017_31316 , \31018_31317 , \31019_31318 , \31020_31319 , \31021_31320 , \31022_31321 , \31023_31322 , \31024_31323 , \31025_31324 , \31026_31325 , \31027_31326 , \31028_31327 , \31029_31328 , \31030_31329 , \31031_31330 , \31032_31331 , \31033_31332 , \31034_31333 , \31035_31334 , \31036_31335 , \31037_31336 , \31038_31337 , \31039_31338 , \31040_31339 , \31041_31340 , \31042_31341 , \31043_31342 , \31044_31343 , \31045_31344 , \31046_31345 , \31047_31346 );
or \U$22254 ( \31049_31348 , \30983_31282 , \31048_31347 );
_DC \g3362/U$1 ( \31050 , \31049_31348 , \9298_9597 );
buf \U$22255 ( \31051_31350 , \31050 );
xor \U$22256 ( \31052_31351 , \30918_31217 , \31051_31350 );
and \U$22257 ( \31053_31352 , RIdec61e8_718, \8760_9059 );
and \U$22258 ( \31054_31353 , RIdec34e8_686, \8762_9061 );
and \U$22259 ( \31055_31354 , RIee20620_4827, \8764_9063 );
and \U$22260 ( \31056_31355 , RIdec07e8_654, \8766_9065 );
and \U$22261 ( \31057_31356 , RIfc4b7b8_5881, \8768_9067 );
and \U$22262 ( \31058_31357 , RIdebdae8_622, \8770_9069 );
and \U$22263 ( \31059_31358 , RIdebade8_590, \8772_9071 );
and \U$22264 ( \31060_31359 , RIdeb80e8_558, \8774_9073 );
and \U$22265 ( \31061_31360 , RIfc41150_5766, \8776_9075 );
and \U$22266 ( \31062_31361 , RIdeb26e8_494, \8778_9077 );
and \U$22267 ( \31063_31362 , RIfc87830_6564, \8780_9079 );
and \U$22268 ( \31064_31363 , RIdeaf9e8_462, \8782_9081 );
and \U$22269 ( \31065_31364 , RIee1dec0_4799, \8784_9083 );
and \U$22270 ( \31066_31365 , RIdeac4f0_430, \8786_9085 );
and \U$22271 ( \31067_31366 , RIdea5bf0_398, \8788_9087 );
and \U$22272 ( \31068_31367 , RIde9f2f0_366, \8790_9089 );
and \U$22273 ( \31069_31368 , RIee1d380_4791, \8792_9091 );
and \U$22274 ( \31070_31369 , RIfc77c78_6385, \8794_9093 );
and \U$22275 ( \31071_31370 , RIfc84f68_6535, \8796_9095 );
and \U$22276 ( \31072_31371 , RIfc6ff50_6296, \8798_9097 );
and \U$22277 ( \31073_31372 , RIde92780_304, \8800_9099 );
and \U$22278 ( \31074_31373 , RIde8efb8_287, \8802_9101 );
and \U$22279 ( \31075_31374 , RIde8ae18_267, \8804_9103 );
and \U$22280 ( \31076_31375 , RIde86c78_247, \8806_9105 );
and \U$22281 ( \31077_31376 , RIee1a680_4759, \8808_9107 );
and \U$22282 ( \31078_31377 , RIee19f78_4754, \8810_9109 );
and \U$22283 ( \31079_31378 , RIfcd7240_7470, \8812_9111 );
and \U$22284 ( \31080_31379 , RIfcbeb50_7192, \8814_9113 );
and \U$22285 ( \31081_31380 , RIfc76328_6367, \8816_9115 );
and \U$22286 ( \31082_31381 , RIe16c2f0_2608, \8818_9117 );
and \U$22287 ( \31083_31382 , RIee388d8_5102, \8820_9119 );
and \U$22288 ( \31084_31383 , RIfea20f0_8188, \8822_9121 );
and \U$22289 ( \31085_31384 , RIe1661e8_2539, \8824_9123 );
and \U$22290 ( \31086_31385 , RIe1634e8_2507, \8826_9125 );
and \U$22291 ( \31087_31386 , RIee37c30_5093, \8828_9127 );
and \U$22292 ( \31088_31387 , RIe1607e8_2475, \8830_9129 );
and \U$22293 ( \31089_31388 , RIfce7500_7654, \8832_9131 );
and \U$22294 ( \31090_31389 , RIe15dae8_2443, \8834_9133 );
and \U$22295 ( \31091_31390 , RIe1580e8_2379, \8836_9135 );
and \U$22296 ( \31092_31391 , RIe1553e8_2347, \8838_9137 );
and \U$22297 ( \31093_31392 , RIfc3f698_5747, \8840_9139 );
and \U$22298 ( \31094_31393 , RIe1526e8_2315, \8842_9141 );
and \U$22299 ( \31095_31394 , RIee354d0_5065, \8844_9143 );
and \U$22300 ( \31096_31395 , RIe14f9e8_2283, \8846_9145 );
and \U$22301 ( \31097_31396 , RIfc83e88_6523, \8848_9147 );
and \U$22302 ( \31098_31397 , RIe14cce8_2251, \8850_9149 );
and \U$22303 ( \31099_31398 , RIe149fe8_2219, \8852_9151 );
and \U$22304 ( \31100_31399 , RIe1472e8_2187, \8854_9153 );
and \U$22305 ( \31101_31400 , RIfcea4d0_7688, \8856_9155 );
and \U$22306 ( \31102_31401 , RIfcb7ad0_7112, \8858_9157 );
and \U$22307 ( \31103_31402 , RIfc695d8_6221, \8860_9159 );
and \U$22308 ( \31104_31403 , RIfc51a28_5951, \8862_9161 );
and \U$22309 ( \31105_31404 , RIe141a50_2124, \8864_9163 );
and \U$22310 ( \31106_31405 , RIe13f728_2099, \8866_9165 );
and \U$22311 ( \31107_31406 , RIdf3d630_2075, \8868_9167 );
and \U$22312 ( \31108_31407 , RIdf3b1a0_2049, \8870_9169 );
and \U$22313 ( \31109_31408 , RIfca9e08_6955, \8872_9171 );
and \U$22314 ( \31110_31409 , RIee2fda0_5003, \8874_9173 );
and \U$22315 ( \31111_31410 , RIfc88a78_6577, \8876_9175 );
and \U$22316 ( \31112_31411 , RIee2da78_4978, \8878_9177 );
and \U$22317 ( \31113_31412 , RIdf36448_1994, \8880_9179 );
and \U$22318 ( \31114_31413 , RIdf33fb8_1968, \8882_9181 );
and \U$22319 ( \31115_31414 , RIdf31df8_1944, \8884_9183 );
and \U$22320 ( \31116_31415 , RIfea2258_8189, \8886_9185 );
or \U$22321 ( \31117_31416 , \31053_31352 , \31054_31353 , \31055_31354 , \31056_31355 , \31057_31356 , \31058_31357 , \31059_31358 , \31060_31359 , \31061_31360 , \31062_31361 , \31063_31362 , \31064_31363 , \31065_31364 , \31066_31365 , \31067_31366 , \31068_31367 , \31069_31368 , \31070_31369 , \31071_31370 , \31072_31371 , \31073_31372 , \31074_31373 , \31075_31374 , \31076_31375 , \31077_31376 , \31078_31377 , \31079_31378 , \31080_31379 , \31081_31380 , \31082_31381 , \31083_31382 , \31084_31383 , \31085_31384 , \31086_31385 , \31087_31386 , \31088_31387 , \31089_31388 , \31090_31389 , \31091_31390 , \31092_31391 , \31093_31392 , \31094_31393 , \31095_31394 , \31096_31395 , \31097_31396 , \31098_31397 , \31099_31398 , \31100_31399 , \31101_31400 , \31102_31401 , \31103_31402 , \31104_31403 , \31105_31404 , \31106_31405 , \31107_31406 , \31108_31407 , \31109_31408 , \31110_31409 , \31111_31410 , \31112_31411 , \31113_31412 , \31114_31413 , \31115_31414 , \31116_31415 );
and \U$22322 ( \31118_31417 , RIee2c560_4963, \8889_9188 );
and \U$22323 ( \31119_31418 , RIee2aaa8_4944, \8891_9190 );
and \U$22324 ( \31120_31419 , RIee29428_4928, \8893_9192 );
and \U$22325 ( \31121_31420 , RIee281e0_4915, \8895_9194 );
and \U$22326 ( \31122_31421 , RIdf2ac10_1863, \8897_9196 );
and \U$22327 ( \31123_31422 , RIdf28d20_1841, \8899_9198 );
and \U$22328 ( \31124_31423 , RIfea27f8_8193, \8901_9200 );
and \U$22329 ( \31125_31424 , RIfea2960_8194, \8903_9202 );
and \U$22330 ( \31126_31425 , RIfcdabe8_7511, \8905_9204 );
and \U$22331 ( \31127_31426 , RIfca08f8_6849, \8907_9206 );
and \U$22332 ( \31128_31427 , RIfc8b1d8_6605, \8909_9208 );
and \U$22333 ( \31129_31428 , RIfc49058_5853, \8911_9210 );
and \U$22334 ( \31130_31429 , RIfca0a60_6850, \8913_9212 );
and \U$22335 ( \31131_31430 , RIdf204b8_1744, \8915_9214 );
and \U$22336 ( \31132_31431 , RIfc99cb0_6772, \8917_9216 );
and \U$22337 ( \31133_31432 , RIdf19f78_1672, \8919_9218 );
and \U$22338 ( \31134_31433 , RIdf17db8_1648, \8921_9220 );
and \U$22339 ( \31135_31434 , RIdf150b8_1616, \8923_9222 );
and \U$22340 ( \31136_31435 , RIdf123b8_1584, \8925_9224 );
and \U$22341 ( \31137_31436 , RIdf0f6b8_1552, \8927_9226 );
and \U$22342 ( \31138_31437 , RIdf0c9b8_1520, \8929_9228 );
and \U$22343 ( \31139_31438 , RIdf09cb8_1488, \8931_9230 );
and \U$22344 ( \31140_31439 , RIdf06fb8_1456, \8933_9232 );
and \U$22345 ( \31141_31440 , RIdf042b8_1424, \8935_9234 );
and \U$22346 ( \31142_31441 , RIdefe8b8_1360, \8937_9236 );
and \U$22347 ( \31143_31442 , RIdefbbb8_1328, \8939_9238 );
and \U$22348 ( \31144_31443 , RIdef8eb8_1296, \8941_9240 );
and \U$22349 ( \31145_31444 , RIdef61b8_1264, \8943_9242 );
and \U$22350 ( \31146_31445 , RIdef34b8_1232, \8945_9244 );
and \U$22351 ( \31147_31446 , RIdef07b8_1200, \8947_9246 );
and \U$22352 ( \31148_31447 , RIdeedab8_1168, \8949_9248 );
and \U$22353 ( \31149_31448 , RIdeeadb8_1136, \8951_9250 );
and \U$22354 ( \31150_31449 , RIfcd1f48_7411, \8953_9252 );
and \U$22355 ( \31151_31450 , RIfc57f68_6023, \8955_9254 );
and \U$22356 ( \31152_31451 , RIfcbe2e0_7186, \8957_9256 );
and \U$22357 ( \31153_31452 , RIfcd8fc8_7491, \8959_9258 );
and \U$22358 ( \31154_31453 , RIdee5520_1073, \8961_9260 );
and \U$22359 ( \31155_31454 , RIfea2690_8192, \8963_9262 );
and \U$22360 ( \31156_31455 , RIdee1470_1027, \8965_9264 );
and \U$22361 ( \31157_31456 , RIdedf418_1004, \8967_9266 );
and \U$22362 ( \31158_31457 , RIfc57b30_6020, \8969_9268 );
and \U$22363 ( \31159_31458 , RIfcb35e8_7063, \8971_9270 );
and \U$22364 ( \31160_31459 , RIfcbd7a0_7178, \8973_9272 );
and \U$22365 ( \31161_31460 , RIfc91178_6673, \8975_9274 );
and \U$22366 ( \31162_31461 , RIfea2528_8191, \8977_9276 );
and \U$22367 ( \31163_31462 , RIded7df8_920, \8979_9278 );
and \U$22368 ( \31164_31463 , RIfea23c0_8190, \8981_9280 );
and \U$22369 ( \31165_31464 , RIded3910_871, \8983_9282 );
and \U$22370 ( \31166_31465 , RIded15e8_846, \8985_9284 );
and \U$22371 ( \31167_31466 , RIdece8e8_814, \8987_9286 );
and \U$22372 ( \31168_31467 , RIdecbbe8_782, \8989_9288 );
and \U$22373 ( \31169_31468 , RIdec8ee8_750, \8991_9290 );
and \U$22374 ( \31170_31469 , RIdeb53e8_526, \8993_9292 );
and \U$22375 ( \31171_31470 , RIde989f0_334, \8995_9294 );
and \U$22376 ( \31172_31471 , RIe16eff0_2640, \8997_9296 );
and \U$22377 ( \31173_31472 , RIe15ade8_2411, \8999_9298 );
and \U$22378 ( \31174_31473 , RIe1445e8_2155, \9001_9300 );
and \U$22379 ( \31175_31474 , RIdf38fe0_2025, \9003_9302 );
and \U$22380 ( \31176_31475 , RIdf2d640_1893, \9005_9304 );
and \U$22381 ( \31177_31476 , RIdf1dec0_1717, \9007_9306 );
and \U$22382 ( \31178_31477 , RIdf015b8_1392, \9009_9308 );
and \U$22383 ( \31179_31478 , RIdee80b8_1104, \9011_9310 );
and \U$22384 ( \31180_31479 , RIdedce20_977, \9013_9312 );
and \U$22385 ( \31181_31480 , RIde7e938_207, \9015_9314 );
or \U$22386 ( \31182_31481 , \31118_31417 , \31119_31418 , \31120_31419 , \31121_31420 , \31122_31421 , \31123_31422 , \31124_31423 , \31125_31424 , \31126_31425 , \31127_31426 , \31128_31427 , \31129_31428 , \31130_31429 , \31131_31430 , \31132_31431 , \31133_31432 , \31134_31433 , \31135_31434 , \31136_31435 , \31137_31436 , \31138_31437 , \31139_31438 , \31140_31439 , \31141_31440 , \31142_31441 , \31143_31442 , \31144_31443 , \31145_31444 , \31146_31445 , \31147_31446 , \31148_31447 , \31149_31448 , \31150_31449 , \31151_31450 , \31152_31451 , \31153_31452 , \31154_31453 , \31155_31454 , \31156_31455 , \31157_31456 , \31158_31457 , \31159_31458 , \31160_31459 , \31161_31460 , \31162_31461 , \31163_31462 , \31164_31463 , \31165_31464 , \31166_31465 , \31167_31466 , \31168_31467 , \31169_31468 , \31170_31469 , \31171_31470 , \31172_31471 , \31173_31472 , \31174_31473 , \31175_31474 , \31176_31475 , \31177_31476 , \31178_31477 , \31179_31478 , \31180_31479 , \31181_31480 );
or \U$22387 ( \31183_31482 , \31117_31416 , \31182_31481 );
_DC \g22ba/U$1 ( \31184 , \31183_31482 , \9024_9323 );
buf \U$22388 ( \31185_31484 , \31184 );
and \U$22389 ( \31186_31485 , RIe19e480_3178, \9034_9333 );
and \U$22390 ( \31187_31486 , RIe19b780_3146, \9036_9335 );
and \U$22391 ( \31188_31487 , RIfccc980_7350, \9038_9337 );
and \U$22392 ( \31189_31488 , RIe198a80_3114, \9040_9339 );
and \U$22393 ( \31190_31489 , RIfcc1148_7219, \9042_9341 );
and \U$22394 ( \31191_31490 , RIe195d80_3082, \9044_9343 );
and \U$22395 ( \31192_31491 , RIe193080_3050, \9046_9345 );
and \U$22396 ( \31193_31492 , RIe190380_3018, \9048_9347 );
and \U$22397 ( \31194_31493 , RIe18a980_2954, \9050_9349 );
and \U$22398 ( \31195_31494 , RIe187c80_2922, \9052_9351 );
and \U$22399 ( \31196_31495 , RIfcb2ee0_7058, \9054_9353 );
and \U$22400 ( \31197_31496 , RIe184f80_2890, \9056_9355 );
and \U$22401 ( \31198_31497 , RIfc615e0_6130, \9058_9357 );
and \U$22402 ( \31199_31498 , RIe182280_2858, \9060_9359 );
and \U$22403 ( \31200_31499 , RIe17f580_2826, \9062_9361 );
and \U$22404 ( \31201_31500 , RIe17c880_2794, \9064_9363 );
and \U$22405 ( \31202_31501 , RIfc69038_6217, \9066_9365 );
and \U$22406 ( \31203_31502 , RIfc4c898_5893, \9068_9367 );
and \U$22407 ( \31204_31503 , RIfc6f2a8_6287, \9070_9369 );
and \U$22408 ( \31205_31504 , RIe1764a8_2723, \9072_9371 );
and \U$22409 ( \31206_31505 , RIfcad0a8_6991, \9074_9373 );
and \U$22410 ( \31207_31506 , RIfc6adc0_6238, \9076_9375 );
and \U$22411 ( \31208_31507 , RIfc70388_6299, \9078_9377 );
and \U$22412 ( \31209_31508 , RIfea1b50_8184, \9080_9379 );
and \U$22413 ( \31210_31509 , RIfea1f88_8187, \9082_9381 );
and \U$22414 ( \31211_31510 , RIfc56e88_6011, \9084_9383 );
and \U$22415 ( \31212_31511 , RIfea1cb8_8185, \9086_9385 );
and \U$22416 ( \31213_31512 , RIe174450_2700, \9088_9387 );
and \U$22417 ( \31214_31513 , RIfc60d70_6124, \9090_9389 );
and \U$22418 ( \31215_31514 , RIfc6a820_6234, \9092_9391 );
and \U$22419 ( \31216_31515 , RIfea1e20_8186, \9094_9393 );
and \U$22420 ( \31217_31516 , RIf16d798_5705, \9096_9395 );
and \U$22421 ( \31218_31517 , RIfc40bb0_5762, \9098_9397 );
and \U$22422 ( \31219_31518 , RIe2247d8_4705, \9100_9399 );
and \U$22423 ( \31220_31519 , RIfc77138_6377, \9102_9401 );
and \U$22424 ( \31221_31520 , RIe221ad8_4673, \9104_9403 );
and \U$22425 ( \31222_31521 , RIfcd7d80_7478, \9106_9405 );
and \U$22426 ( \31223_31522 , RIe21edd8_4641, \9108_9407 );
and \U$22427 ( \31224_31523 , RIe2193d8_4577, \9110_9409 );
and \U$22428 ( \31225_31524 , RIe2166d8_4545, \9112_9411 );
and \U$22429 ( \31226_31525 , RIfc40070_5754, \9114_9413 );
and \U$22430 ( \31227_31526 , RIe2139d8_4513, \9116_9415 );
and \U$22431 ( \31228_31527 , RIf169850_5660, \9118_9417 );
and \U$22432 ( \31229_31528 , RIe210cd8_4481, \9120_9419 );
and \U$22433 ( \31230_31529 , RIfcc1580_7222, \9122_9421 );
and \U$22434 ( \31231_31530 , RIe20dfd8_4449, \9124_9423 );
and \U$22435 ( \31232_31531 , RIe20b2d8_4417, \9126_9425 );
and \U$22436 ( \31233_31532 , RIe2085d8_4385, \9128_9427 );
and \U$22437 ( \31234_31533 , RIfcd0058_7389, \9130_9429 );
and \U$22438 ( \31235_31534 , RIfc749d8_6349, \9132_9431 );
and \U$22439 ( \31236_31535 , RIe203010_4324, \9134_9433 );
and \U$22440 ( \31237_31536 , RIe2013f0_4304, \9136_9435 );
and \U$22441 ( \31238_31537 , RIfc60230_6116, \9138_9437 );
and \U$22442 ( \31239_31538 , RIfc60668_6119, \9140_9439 );
and \U$22443 ( \31240_31539 , RIfcaf970_7020, \9142_9441 );
and \U$22444 ( \31241_31540 , RIfc45818_5813, \9144_9443 );
and \U$22445 ( \31242_31541 , RIf160a48_5559, \9146_9445 );
and \U$22446 ( \31243_31542 , RIf15eb58_5537, \9148_9447 );
and \U$22447 ( \31244_31543 , RIfea1880_8182, \9150_9449 );
and \U$22448 ( \31245_31544 , RIfea19e8_8183, \9152_9451 );
and \U$22449 ( \31246_31545 , RIfc72110_6320, \9154_9453 );
and \U$22450 ( \31247_31546 , RIfc49b98_5861, \9156_9455 );
and \U$22451 ( \31248_31547 , RIfcca0b8_7321, \9158_9457 );
and \U$22452 ( \31249_31548 , RIfc71738_6313, \9160_9459 );
or \U$22453 ( \31250_31549 , \31186_31485 , \31187_31486 , \31188_31487 , \31189_31488 , \31190_31489 , \31191_31490 , \31192_31491 , \31193_31492 , \31194_31493 , \31195_31494 , \31196_31495 , \31197_31496 , \31198_31497 , \31199_31498 , \31200_31499 , \31201_31500 , \31202_31501 , \31203_31502 , \31204_31503 , \31205_31504 , \31206_31505 , \31207_31506 , \31208_31507 , \31209_31508 , \31210_31509 , \31211_31510 , \31212_31511 , \31213_31512 , \31214_31513 , \31215_31514 , \31216_31515 , \31217_31516 , \31218_31517 , \31219_31518 , \31220_31519 , \31221_31520 , \31222_31521 , \31223_31522 , \31224_31523 , \31225_31524 , \31226_31525 , \31227_31526 , \31228_31527 , \31229_31528 , \31230_31529 , \31231_31530 , \31232_31531 , \31233_31532 , \31234_31533 , \31235_31534 , \31236_31535 , \31237_31536 , \31238_31537 , \31239_31538 , \31240_31539 , \31241_31540 , \31242_31541 , \31243_31542 , \31244_31543 , \31245_31544 , \31246_31545 , \31247_31546 , \31248_31547 , \31249_31548 );
and \U$22454 ( \31251_31550 , RIfc4ca00_5894, \9163_9462 );
and \U$22455 ( \31252_31551 , RIfc71030_6308, \9165_9464 );
and \U$22456 ( \31253_31552 , RIfcde428_7551, \9167_9466 );
and \U$22457 ( \31254_31553 , RIe1fad48_4231, \9169_9468 );
and \U$22458 ( \31255_31554 , RIfc70bf8_6305, \9171_9470 );
and \U$22459 ( \31256_31555 , RIfc63a70_6156, \9173_9472 );
and \U$22460 ( \31257_31556 , RIfca7db0_6932, \9175_9474 );
and \U$22461 ( \31258_31557 , RIe1f62c0_4178, \9177_9476 );
and \U$22462 ( \31259_31558 , RIfcada80_6998, \9179_9478 );
and \U$22463 ( \31260_31559 , RIfc6fde8_6295, \9181_9480 );
and \U$22464 ( \31261_31560 , RIfc6f578_6289, \9183_9482 );
and \U$22465 ( \31262_31561 , RIe1f3f98_4153, \9185_9484 );
and \U$22466 ( \31263_31562 , RIfcde158_7549, \9187_9486 );
and \U$22467 ( \31264_31563 , RIfcad378_6993, \9189_9488 );
and \U$22468 ( \31265_31564 , RIfc65f00_6182, \9191_9490 );
and \U$22469 ( \31266_31565 , RIe1eeca0_4094, \9193_9492 );
and \U$22470 ( \31267_31566 , RIe1ec540_4066, \9195_9494 );
and \U$22471 ( \31268_31567 , RIe1e9840_4034, \9197_9496 );
and \U$22472 ( \31269_31568 , RIe1e6b40_4002, \9199_9498 );
and \U$22473 ( \31270_31569 , RIe1e3e40_3970, \9201_9500 );
and \U$22474 ( \31271_31570 , RIe1e1140_3938, \9203_9502 );
and \U$22475 ( \31272_31571 , RIe1de440_3906, \9205_9504 );
and \U$22476 ( \31273_31572 , RIe1db740_3874, \9207_9506 );
and \U$22477 ( \31274_31573 , RIe1d8a40_3842, \9209_9508 );
and \U$22478 ( \31275_31574 , RIe1d3040_3778, \9211_9510 );
and \U$22479 ( \31276_31575 , RIe1d0340_3746, \9213_9512 );
and \U$22480 ( \31277_31576 , RIe1cd640_3714, \9215_9514 );
and \U$22481 ( \31278_31577 , RIe1ca940_3682, \9217_9516 );
and \U$22482 ( \31279_31578 , RIe1c7c40_3650, \9219_9518 );
and \U$22483 ( \31280_31579 , RIe1c4f40_3618, \9221_9520 );
and \U$22484 ( \31281_31580 , RIe1c2240_3586, \9223_9522 );
and \U$22485 ( \31282_31581 , RIe1bf540_3554, \9225_9524 );
and \U$22486 ( \31283_31582 , RIfc69308_6219, \9227_9526 );
and \U$22487 ( \31284_31583 , RIfccba08_7339, \9229_9528 );
and \U$22488 ( \31285_31584 , RIe1b9f78_3493, \9231_9530 );
and \U$22489 ( \31286_31585 , RIe1b7db8_3469, \9233_9532 );
and \U$22490 ( \31287_31586 , RIfccd628_7359, \9235_9534 );
and \U$22491 ( \31288_31587 , RIfc69740_6222, \9237_9536 );
and \U$22492 ( \31289_31588 , RIe1b5bf8_3445, \9239_9538 );
and \U$22493 ( \31290_31589 , RIe1b4578_3429, \9241_9540 );
and \U$22494 ( \31291_31590 , RIfccf950_7384, \9243_9542 );
and \U$22495 ( \31292_31591 , RIf148088_5279, \9245_9544 );
and \U$22496 ( \31293_31592 , RIe1b3060_3414, \9247_9546 );
and \U$22497 ( \31294_31593 , RIe1b1710_3396, \9249_9548 );
and \U$22498 ( \31295_31594 , RIfc9f818_6837, \9251_9550 );
and \U$22499 ( \31296_31595 , RIfcb9c90_7136, \9253_9552 );
and \U$22500 ( \31297_31596 , RIe1acf58_3345, \9255_9554 );
and \U$22501 ( \31298_31597 , RIe1ab770_3328, \9257_9556 );
and \U$22502 ( \31299_31598 , RIe1a9880_3306, \9259_9558 );
and \U$22503 ( \31300_31599 , RIe1a6b80_3274, \9261_9560 );
and \U$22504 ( \31301_31600 , RIe1a3e80_3242, \9263_9562 );
and \U$22505 ( \31302_31601 , RIe1a1180_3210, \9265_9564 );
and \U$22506 ( \31303_31602 , RIe18d680_2986, \9267_9566 );
and \U$22507 ( \31304_31603 , RIe179b80_2762, \9269_9568 );
and \U$22508 ( \31305_31604 , RIe2274d8_4737, \9271_9570 );
and \U$22509 ( \31306_31605 , RIe21c0d8_4609, \9273_9572 );
and \U$22510 ( \31307_31606 , RIe2058d8_4353, \9275_9574 );
and \U$22511 ( \31308_31607 , RIe1ff938_4285, \9277_9576 );
and \U$22512 ( \31309_31608 , RIe1f8cf0_4208, \9279_9578 );
and \U$22513 ( \31310_31609 , RIe1f1838_4125, \9281_9580 );
and \U$22514 ( \31311_31610 , RIe1d5d40_3810, \9283_9582 );
and \U$22515 ( \31312_31611 , RIe1bc840_3522, \9285_9584 );
and \U$22516 ( \31313_31612 , RIe1af6b8_3373, \9287_9586 );
and \U$22517 ( \31314_31613 , RIe171cf0_2672, \9289_9588 );
or \U$22518 ( \31315_31614 , \31251_31550 , \31252_31551 , \31253_31552 , \31254_31553 , \31255_31554 , \31256_31555 , \31257_31556 , \31258_31557 , \31259_31558 , \31260_31559 , \31261_31560 , \31262_31561 , \31263_31562 , \31264_31563 , \31265_31564 , \31266_31565 , \31267_31566 , \31268_31567 , \31269_31568 , \31270_31569 , \31271_31570 , \31272_31571 , \31273_31572 , \31274_31573 , \31275_31574 , \31276_31575 , \31277_31576 , \31278_31577 , \31279_31578 , \31280_31579 , \31281_31580 , \31282_31581 , \31283_31582 , \31284_31583 , \31285_31584 , \31286_31585 , \31287_31586 , \31288_31587 , \31289_31588 , \31290_31589 , \31291_31590 , \31292_31591 , \31293_31592 , \31294_31593 , \31295_31594 , \31296_31595 , \31297_31596 , \31298_31597 , \31299_31598 , \31300_31599 , \31301_31600 , \31302_31601 , \31303_31602 , \31304_31603 , \31305_31604 , \31306_31605 , \31307_31606 , \31308_31607 , \31309_31608 , \31310_31609 , \31311_31610 , \31312_31611 , \31313_31612 , \31314_31613 );
or \U$22519 ( \31316_31615 , \31250_31549 , \31315_31614 );
_DC \g33e7/U$1 ( \31317 , \31316_31615 , \9298_9597 );
buf \U$22520 ( \31318_31617 , \31317 );
and \U$22521 ( \31319_31618 , \31185_31484 , \31318_31617 );
and \U$22522 ( \31320_31619 , \29135_29434 , \29268_29567 );
and \U$22523 ( \31321_31620 , \29268_29567 , \29543_29842 );
and \U$22524 ( \31322_31621 , \29135_29434 , \29543_29842 );
or \U$22525 ( \31323_31622 , \31320_31619 , \31321_31620 , \31322_31621 );
and \U$22526 ( \31324_31623 , \31318_31617 , \31323_31622 );
and \U$22527 ( \31325_31624 , \31185_31484 , \31323_31622 );
or \U$22528 ( \31326_31625 , \31319_31618 , \31324_31623 , \31325_31624 );
xor \U$22529 ( \31327_31626 , \31052_31351 , \31326_31625 );
buf g43fa_GF_PartitionCandidate( \31328_31627_nG43fa , \31327_31626 );
xor \U$22530 ( \31329_31628 , \31185_31484 , \31318_31617 );
xor \U$22531 ( \31330_31629 , \31329_31628 , \31323_31622 );
buf g43fd_GF_PartitionCandidate( \31331_31630_nG43fd , \31330_31629 );
nand \U$22532 ( \31332_31631 , \31331_31630_nG43fd , \29545_29844_nG4400 );
and \U$22533 ( \31333_31632 , \31328_31627_nG43fa , \31332_31631 );
xor \U$22534 ( \31334_31633 , \31331_31630_nG43fd , \29545_29844_nG4400 );
and \U$22539 ( \31335_31637 , \31334_31633 , \10392_10694_nG9c0e );
or \U$22540 ( \31336_31638 , 1'b0 , \31335_31637 );
xor \U$22541 ( \31337_31639 , \31333_31632 , \31336_31638 );
xor \U$22542 ( \31338_31640 , \31333_31632 , \31337_31639 );
buf \U$22543 ( \31339_31641 , \31338_31640 );
buf \U$22544 ( \31340_31642 , \31339_31641 );
xor \U$22545 ( \31341_31643 , \30785_31084 , \31340_31642 );
and \U$22546 ( \31342_31644 , \30726_31025 , \30731_31030 );
and \U$22547 ( \31343_31645 , \30726_31025 , \30778_31077 );
and \U$22548 ( \31344_31646 , \30731_31030 , \30778_31077 );
or \U$22549 ( \31345_31647 , \31342_31644 , \31343_31645 , \31344_31646 );
and \U$22550 ( \31346_31648 , \31341_31643 , \31345_31647 );
and \U$22551 ( \31347_31649 , \30765_31064 , \30770_31069 );
and \U$22552 ( \31348_31650 , \30765_31064 , \30776_31075 );
and \U$22553 ( \31349_31651 , \30770_31069 , \30776_31075 );
or \U$22554 ( \31350_31652 , \31347_31649 , \31348_31650 , \31349_31651 );
buf \U$22555 ( \31351_31653 , \31350_31652 );
and \U$22556 ( \31352_31654 , \30645_30947 , \30650_30952 );
and \U$22557 ( \31353_31655 , \30645_30947 , \30724_31023 );
and \U$22558 ( \31354_31656 , \30650_30952 , \30724_31023 );
or \U$22559 ( \31355_31657 , \31352_31654 , \31353_31655 , \31354_31656 );
buf \U$22560 ( \31356_31658 , \31355_31657 );
and \U$22561 ( \31357_31659 , \30709_31008 , \30715_31014 );
and \U$22562 ( \31358_31660 , \30709_31008 , \30722_31021 );
and \U$22563 ( \31359_31661 , \30715_31014 , \30722_31021 );
or \U$22564 ( \31360_31662 , \31357_31659 , \31358_31660 , \31359_31661 );
buf \U$22565 ( \31361_31663 , \31360_31662 );
and \U$22566 ( \31362_31664 , \30694_30993 , \30700_30999 );
and \U$22567 ( \31363_31665 , \30694_30993 , \30707_31006 );
and \U$22568 ( \31364_31666 , \30700_30999 , \30707_31006 );
or \U$22569 ( \31365_31667 , \31362_31664 , \31363_31665 , \31364_31666 );
buf \U$22570 ( \31366_31668 , \31365_31667 );
and \U$22571 ( \31367_31669 , \20353_20155 , \17808_18107_nG9be7 );
and \U$22572 ( \31368_31670 , \19853_20152 , \18789_19091_nG9be4 );
or \U$22573 ( \31369_31671 , \31367_31669 , \31368_31670 );
xor \U$22574 ( \31370_31672 , \19852_20151 , \31369_31671 );
buf \U$22575 ( \31371_31673 , \31370_31672 );
buf \U$22577 ( \31372_31674 , \31371_31673 );
and \U$22578 ( \31373_31675 , \18908_18702 , \19287_19586_nG9be1 );
and \U$22579 ( \31374_31676 , \18400_18699 , \20306_20608_nG9bde );
or \U$22580 ( \31375_31677 , \31373_31675 , \31374_31676 );
xor \U$22581 ( \31376_31678 , \18399_18698 , \31375_31677 );
buf \U$22582 ( \31377_31679 , \31376_31678 );
buf \U$22584 ( \31378_31680 , \31377_31679 );
xor \U$22585 ( \31379_31681 , \31372_31674 , \31378_31680 );
and \U$22586 ( \31380_31682 , \17437_17297 , \20787_21086_nG9bdb );
and \U$22587 ( \31381_31683 , \16995_17294 , \21827_22129_nG9bd8 );
or \U$22588 ( \31382_31684 , \31380_31682 , \31381_31683 );
xor \U$22589 ( \31383_31685 , \16994_17293 , \31382_31684 );
buf \U$22590 ( \31384_31686 , \31383_31685 );
buf \U$22592 ( \31385_31687 , \31384_31686 );
xor \U$22593 ( \31386_31688 , \31379_31681 , \31385_31687 );
buf \U$22594 ( \31387_31689 , \31386_31688 );
xor \U$22595 ( \31388_31690 , \31366_31668 , \31387_31689 );
and \U$22596 ( \31389_31691 , \12183_12157 , \27114_27416_nG9bc3 );
and \U$22597 ( \31390_31692 , \11855_12154 , \28300_28602_nG9bc0 );
or \U$22598 ( \31391_31693 , \31389_31691 , \31390_31692 );
xor \U$22599 ( \31392_31694 , \11854_12153 , \31391_31693 );
buf \U$22600 ( \31393_31695 , \31392_31694 );
buf \U$22602 ( \31394_31696 , \31393_31695 );
xor \U$22603 ( \31395_31697 , \31388_31690 , \31394_31696 );
buf \U$22604 ( \31396_31698 , \31395_31697 );
xor \U$22605 ( \31397_31699 , \31361_31663 , \31396_31698 );
and \U$22606 ( \31398_31700 , \30737_31036 , \30743_31042 );
and \U$22607 ( \31399_31701 , \30737_31036 , \30750_31049 );
and \U$22608 ( \31400_31702 , \30743_31042 , \30750_31049 );
or \U$22609 ( \31401_31703 , \31398_31700 , \31399_31701 , \31400_31702 );
buf \U$22610 ( \31402_31704 , \31401_31703 );
xor \U$22611 ( \31403_31705 , \31397_31699 , \31402_31704 );
buf \U$22612 ( \31404_31706 , \31403_31705 );
xor \U$22613 ( \31405_31707 , \31356_31658 , \31404_31706 );
and \U$22614 ( \31406_31708 , \30194_30496 , \30199_30501 );
and \U$22615 ( \31407_31709 , \30194_30496 , \30206_30508 );
and \U$22616 ( \31408_31710 , \30199_30501 , \30206_30508 );
or \U$22617 ( \31409_31711 , \31406_31708 , \31407_31709 , \31408_31710 );
buf \U$22618 ( \31410_31712 , \31409_31711 );
and \U$22619 ( \31411_31713 , \30170_30472 , \30176_30478 );
and \U$22620 ( \31412_31714 , \30170_30472 , \30183_30485 );
and \U$22621 ( \31413_31715 , \30176_30478 , \30183_30485 );
or \U$22622 ( \31414_31716 , \31411_31713 , \31412_31714 , \31413_31715 );
buf \U$22623 ( \31415_31717 , \31414_31716 );
and \U$22624 ( \31416_31718 , \30659_30961 , \30665_30967 );
buf \U$22625 ( \31417_31719 , \31416_31718 );
and \U$22626 ( \31418_31720 , \27141_26431 , \12502_12801_nG9bff );
and \U$22627 ( \31419_31721 , \26129_26428 , \13403_13705_nG9bfc );
or \U$22628 ( \31420_31722 , \31418_31720 , \31419_31721 );
xor \U$22629 ( \31421_31723 , \26128_26427 , \31420_31722 );
buf \U$22630 ( \31422_31724 , \31421_31723 );
buf \U$22632 ( \31423_31725 , \31422_31724 );
xor \U$22633 ( \31424_31726 , \31417_31719 , \31423_31725 );
and \U$22634 ( \31425_31727 , \25044_24792 , \13771_14070_nG9bf9 );
and \U$22635 ( \31426_31728 , \24490_24789 , \14682_14984_nG9bf6 );
or \U$22636 ( \31427_31729 , \31425_31727 , \31426_31728 );
xor \U$22637 ( \31428_31730 , \24489_24788 , \31427_31729 );
buf \U$22638 ( \31429_31731 , \31428_31730 );
buf \U$22640 ( \31430_31732 , \31429_31731 );
xor \U$22641 ( \31431_31733 , \31424_31726 , \31430_31732 );
buf \U$22642 ( \31432_31734 , \31431_31733 );
xor \U$22643 ( \31433_31735 , \31415_31717 , \31432_31734 );
and \U$22644 ( \31434_31736 , \21908_21658 , \16378_16680_nG9bed );
and \U$22645 ( \31435_31737 , \21356_21655 , \17363_17665_nG9bea );
or \U$22646 ( \31436_31738 , \31434_31736 , \31435_31737 );
xor \U$22647 ( \31437_31739 , \21355_21654 , \31436_31738 );
buf \U$22648 ( \31438_31740 , \31437_31739 );
buf \U$22650 ( \31439_31741 , \31438_31740 );
xor \U$22651 ( \31440_31742 , \31433_31735 , \31439_31741 );
buf \U$22652 ( \31441_31743 , \31440_31742 );
and \U$22653 ( \31442_31744 , \16405_15940 , \22330_22629_nG9bd5 );
and \U$22654 ( \31443_31745 , \15638_15937 , \23394_23696_nG9bd2 );
or \U$22655 ( \31444_31746 , \31442_31744 , \31443_31745 );
xor \U$22656 ( \31445_31747 , \15637_15936 , \31444_31746 );
buf \U$22657 ( \31446_31748 , \31445_31747 );
buf \U$22659 ( \31447_31749 , \31446_31748 );
xor \U$22660 ( \31448_31750 , \31441_31743 , \31447_31749 );
and \U$22661 ( \31449_31751 , \14710_14631 , \23927_24226_nG9bcf );
and \U$22662 ( \31450_31752 , \14329_14628 , \24996_25298_nG9bcc );
or \U$22663 ( \31451_31753 , \31449_31751 , \31450_31752 );
xor \U$22664 ( \31452_31754 , \14328_14627 , \31451_31753 );
buf \U$22665 ( \31453_31755 , \31452_31754 );
buf \U$22667 ( \31454_31756 , \31453_31755 );
xor \U$22668 ( \31455_31757 , \31448_31750 , \31454_31756 );
buf \U$22669 ( \31456_31758 , \31455_31757 );
xor \U$22670 ( \31457_31759 , \31410_31712 , \31456_31758 );
and \U$22671 ( \31458_31760 , \10411_10707 , \30638_30940_nG9bb7 );
and \U$22672 ( \31459_31761 , \30527_30829 , \30571_30873 );
and \U$22673 ( \31460_31762 , \30571_30873 , \30626_30928 );
and \U$22674 ( \31461_31763 , \30527_30829 , \30626_30928 );
or \U$22675 ( \31462_31764 , \31459_31761 , \31460_31762 , \31461_31763 );
and \U$22676 ( \31463_31765 , \30228_30530 , \30232_30534 );
and \U$22677 ( \31464_31766 , \30232_30534 , \30526_30828 );
and \U$22678 ( \31465_31767 , \30228_30530 , \30526_30828 );
or \U$22679 ( \31466_31768 , \31463_31765 , \31464_31766 , \31465_31767 );
and \U$22680 ( \31467_31769 , \30531_30833 , \30545_30847 );
and \U$22681 ( \31468_31770 , \30545_30847 , \30570_30872 );
and \U$22682 ( \31469_31771 , \30531_30833 , \30570_30872 );
or \U$22683 ( \31470_31772 , \31467_31769 , \31468_31770 , \31469_31771 );
xor \U$22684 ( \31471_31773 , \31466_31768 , \31470_31772 );
and \U$22685 ( \31472_31774 , \20734_21033 , \17791_18090 );
and \U$22686 ( \31473_31775 , \21788_22090 , \17353_17655 );
nor \U$22687 ( \31474_31776 , \31472_31774 , \31473_31775 );
xnor \U$22688 ( \31475_31777 , \31474_31776 , \17747_18046 );
and \U$22689 ( \31476_31778 , \12470_12769 , \27095_27397 );
and \U$22690 ( \31477_31779 , \13377_13679 , \26505_26807 );
nor \U$22691 ( \31478_31780 , \31476_31778 , \31477_31779 );
xnor \U$22692 ( \31479_31781 , \31478_31780 , \26993_27295 );
xor \U$22693 ( \31480_31782 , \31475_31777 , \31479_31781 );
and \U$22694 ( \31481_31783 , \11287_11586 , \28768_29070 );
and \U$22695 ( \31482_31784 , \12146_12448 , \28224_28526 );
nor \U$22696 ( \31483_31785 , \31481_31783 , \31482_31784 );
xnor \U$22697 ( \31484_31786 , \31483_31785 , \28774_29076 );
xor \U$22698 ( \31485_31787 , \31480_31782 , \31484_31786 );
and \U$22699 ( \31486_31788 , \30500_30802 , \10681_10983 );
and \U$22700 ( \31487_31789 , RIdec61e8_718, \9034_9333 );
and \U$22701 ( \31488_31790 , RIdec34e8_686, \9036_9335 );
and \U$22702 ( \31489_31791 , RIee20620_4827, \9038_9337 );
and \U$22703 ( \31490_31792 , RIdec07e8_654, \9040_9339 );
and \U$22704 ( \31491_31793 , RIfc4b7b8_5881, \9042_9341 );
and \U$22705 ( \31492_31794 , RIdebdae8_622, \9044_9343 );
and \U$22706 ( \31493_31795 , RIdebade8_590, \9046_9345 );
and \U$22707 ( \31494_31796 , RIdeb80e8_558, \9048_9347 );
and \U$22708 ( \31495_31797 , RIfc41150_5766, \9050_9349 );
and \U$22709 ( \31496_31798 , RIdeb26e8_494, \9052_9351 );
and \U$22710 ( \31497_31799 , RIfc87830_6564, \9054_9353 );
and \U$22711 ( \31498_31800 , RIdeaf9e8_462, \9056_9355 );
and \U$22712 ( \31499_31801 , RIee1dec0_4799, \9058_9357 );
and \U$22713 ( \31500_31802 , RIdeac4f0_430, \9060_9359 );
and \U$22714 ( \31501_31803 , RIdea5bf0_398, \9062_9361 );
and \U$22715 ( \31502_31804 , RIde9f2f0_366, \9064_9363 );
and \U$22716 ( \31503_31805 , RIee1d380_4791, \9066_9365 );
and \U$22717 ( \31504_31806 , RIfc77c78_6385, \9068_9367 );
and \U$22718 ( \31505_31807 , RIfc84f68_6535, \9070_9369 );
and \U$22719 ( \31506_31808 , RIfc6ff50_6296, \9072_9371 );
and \U$22720 ( \31507_31809 , RIde92780_304, \9074_9373 );
and \U$22721 ( \31508_31810 , RIde8efb8_287, \9076_9375 );
and \U$22722 ( \31509_31811 , RIde8ae18_267, \9078_9377 );
and \U$22723 ( \31510_31812 , RIde86c78_247, \9080_9379 );
and \U$22724 ( \31511_31813 , RIee1a680_4759, \9082_9381 );
and \U$22725 ( \31512_31814 , RIee19f78_4754, \9084_9383 );
and \U$22726 ( \31513_31815 , RIfcd7240_7470, \9086_9385 );
and \U$22727 ( \31514_31816 , RIfcbeb50_7192, \9088_9387 );
and \U$22728 ( \31515_31817 , RIfc76328_6367, \9090_9389 );
and \U$22729 ( \31516_31818 , RIe16c2f0_2608, \9092_9391 );
and \U$22730 ( \31517_31819 , RIee388d8_5102, \9094_9393 );
and \U$22731 ( \31518_31820 , RIfea20f0_8188, \9096_9395 );
and \U$22732 ( \31519_31821 , RIe1661e8_2539, \9098_9397 );
and \U$22733 ( \31520_31822 , RIe1634e8_2507, \9100_9399 );
and \U$22734 ( \31521_31823 , RIee37c30_5093, \9102_9401 );
and \U$22735 ( \31522_31824 , RIe1607e8_2475, \9104_9403 );
and \U$22736 ( \31523_31825 , RIfce7500_7654, \9106_9405 );
and \U$22737 ( \31524_31826 , RIe15dae8_2443, \9108_9407 );
and \U$22738 ( \31525_31827 , RIe1580e8_2379, \9110_9409 );
and \U$22739 ( \31526_31828 , RIe1553e8_2347, \9112_9411 );
and \U$22740 ( \31527_31829 , RIfc3f698_5747, \9114_9413 );
and \U$22741 ( \31528_31830 , RIe1526e8_2315, \9116_9415 );
and \U$22742 ( \31529_31831 , RIee354d0_5065, \9118_9417 );
and \U$22743 ( \31530_31832 , RIe14f9e8_2283, \9120_9419 );
and \U$22744 ( \31531_31833 , RIfc83e88_6523, \9122_9421 );
and \U$22745 ( \31532_31834 , RIe14cce8_2251, \9124_9423 );
and \U$22746 ( \31533_31835 , RIe149fe8_2219, \9126_9425 );
and \U$22747 ( \31534_31836 , RIe1472e8_2187, \9128_9427 );
and \U$22748 ( \31535_31837 , RIfcea4d0_7688, \9130_9429 );
and \U$22749 ( \31536_31838 , RIfcb7ad0_7112, \9132_9431 );
and \U$22750 ( \31537_31839 , RIfc695d8_6221, \9134_9433 );
and \U$22751 ( \31538_31840 , RIfc51a28_5951, \9136_9435 );
and \U$22752 ( \31539_31841 , RIe141a50_2124, \9138_9437 );
and \U$22753 ( \31540_31842 , RIe13f728_2099, \9140_9439 );
and \U$22754 ( \31541_31843 , RIdf3d630_2075, \9142_9441 );
and \U$22755 ( \31542_31844 , RIdf3b1a0_2049, \9144_9443 );
and \U$22756 ( \31543_31845 , RIfca9e08_6955, \9146_9445 );
and \U$22757 ( \31544_31846 , RIee2fda0_5003, \9148_9447 );
and \U$22758 ( \31545_31847 , RIfc88a78_6577, \9150_9449 );
and \U$22759 ( \31546_31848 , RIee2da78_4978, \9152_9451 );
and \U$22760 ( \31547_31849 , RIdf36448_1994, \9154_9453 );
and \U$22761 ( \31548_31850 , RIdf33fb8_1968, \9156_9455 );
and \U$22762 ( \31549_31851 , RIdf31df8_1944, \9158_9457 );
and \U$22763 ( \31550_31852 , RIfea2258_8189, \9160_9459 );
or \U$22764 ( \31551_31853 , \31487_31789 , \31488_31790 , \31489_31791 , \31490_31792 , \31491_31793 , \31492_31794 , \31493_31795 , \31494_31796 , \31495_31797 , \31496_31798 , \31497_31799 , \31498_31800 , \31499_31801 , \31500_31802 , \31501_31803 , \31502_31804 , \31503_31805 , \31504_31806 , \31505_31807 , \31506_31808 , \31507_31809 , \31508_31810 , \31509_31811 , \31510_31812 , \31511_31813 , \31512_31814 , \31513_31815 , \31514_31816 , \31515_31817 , \31516_31818 , \31517_31819 , \31518_31820 , \31519_31821 , \31520_31822 , \31521_31823 , \31522_31824 , \31523_31825 , \31524_31826 , \31525_31827 , \31526_31828 , \31527_31829 , \31528_31830 , \31529_31831 , \31530_31832 , \31531_31833 , \31532_31834 , \31533_31835 , \31534_31836 , \31535_31837 , \31536_31838 , \31537_31839 , \31538_31840 , \31539_31841 , \31540_31842 , \31541_31843 , \31542_31844 , \31543_31845 , \31544_31846 , \31545_31847 , \31546_31848 , \31547_31849 , \31548_31850 , \31549_31851 , \31550_31852 );
and \U$22765 ( \31552_31854 , RIee2c560_4963, \9163_9462 );
and \U$22766 ( \31553_31855 , RIee2aaa8_4944, \9165_9464 );
and \U$22767 ( \31554_31856 , RIee29428_4928, \9167_9466 );
and \U$22768 ( \31555_31857 , RIee281e0_4915, \9169_9468 );
and \U$22769 ( \31556_31858 , RIdf2ac10_1863, \9171_9470 );
and \U$22770 ( \31557_31859 , RIdf28d20_1841, \9173_9472 );
and \U$22771 ( \31558_31860 , RIfea27f8_8193, \9175_9474 );
and \U$22772 ( \31559_31861 , RIfea2960_8194, \9177_9476 );
and \U$22773 ( \31560_31862 , RIfcdabe8_7511, \9179_9478 );
and \U$22774 ( \31561_31863 , RIfca08f8_6849, \9181_9480 );
and \U$22775 ( \31562_31864 , RIfc8b1d8_6605, \9183_9482 );
and \U$22776 ( \31563_31865 , RIfc49058_5853, \9185_9484 );
and \U$22777 ( \31564_31866 , RIfca0a60_6850, \9187_9486 );
and \U$22778 ( \31565_31867 , RIdf204b8_1744, \9189_9488 );
and \U$22779 ( \31566_31868 , RIfc99cb0_6772, \9191_9490 );
and \U$22780 ( \31567_31869 , RIdf19f78_1672, \9193_9492 );
and \U$22781 ( \31568_31870 , RIdf17db8_1648, \9195_9494 );
and \U$22782 ( \31569_31871 , RIdf150b8_1616, \9197_9496 );
and \U$22783 ( \31570_31872 , RIdf123b8_1584, \9199_9498 );
and \U$22784 ( \31571_31873 , RIdf0f6b8_1552, \9201_9500 );
and \U$22785 ( \31572_31874 , RIdf0c9b8_1520, \9203_9502 );
and \U$22786 ( \31573_31875 , RIdf09cb8_1488, \9205_9504 );
and \U$22787 ( \31574_31876 , RIdf06fb8_1456, \9207_9506 );
and \U$22788 ( \31575_31877 , RIdf042b8_1424, \9209_9508 );
and \U$22789 ( \31576_31878 , RIdefe8b8_1360, \9211_9510 );
and \U$22790 ( \31577_31879 , RIdefbbb8_1328, \9213_9512 );
and \U$22791 ( \31578_31880 , RIdef8eb8_1296, \9215_9514 );
and \U$22792 ( \31579_31881 , RIdef61b8_1264, \9217_9516 );
and \U$22793 ( \31580_31882 , RIdef34b8_1232, \9219_9518 );
and \U$22794 ( \31581_31883 , RIdef07b8_1200, \9221_9520 );
and \U$22795 ( \31582_31884 , RIdeedab8_1168, \9223_9522 );
and \U$22796 ( \31583_31885 , RIdeeadb8_1136, \9225_9524 );
and \U$22797 ( \31584_31886 , RIfcd1f48_7411, \9227_9526 );
and \U$22798 ( \31585_31887 , RIfc57f68_6023, \9229_9528 );
and \U$22799 ( \31586_31888 , RIfcbe2e0_7186, \9231_9530 );
and \U$22800 ( \31587_31889 , RIfcd8fc8_7491, \9233_9532 );
and \U$22801 ( \31588_31890 , RIdee5520_1073, \9235_9534 );
and \U$22802 ( \31589_31891 , RIfea2690_8192, \9237_9536 );
and \U$22803 ( \31590_31892 , RIdee1470_1027, \9239_9538 );
and \U$22804 ( \31591_31893 , RIdedf418_1004, \9241_9540 );
and \U$22805 ( \31592_31894 , RIfc57b30_6020, \9243_9542 );
and \U$22806 ( \31593_31895 , RIfcb35e8_7063, \9245_9544 );
and \U$22807 ( \31594_31896 , RIfcbd7a0_7178, \9247_9546 );
and \U$22808 ( \31595_31897 , RIfc91178_6673, \9249_9548 );
and \U$22809 ( \31596_31898 , RIfea2528_8191, \9251_9550 );
and \U$22810 ( \31597_31899 , RIded7df8_920, \9253_9552 );
and \U$22811 ( \31598_31900 , RIfea23c0_8190, \9255_9554 );
and \U$22812 ( \31599_31901 , RIded3910_871, \9257_9556 );
and \U$22813 ( \31600_31902 , RIded15e8_846, \9259_9558 );
and \U$22814 ( \31601_31903 , RIdece8e8_814, \9261_9560 );
and \U$22815 ( \31602_31904 , RIdecbbe8_782, \9263_9562 );
and \U$22816 ( \31603_31905 , RIdec8ee8_750, \9265_9564 );
and \U$22817 ( \31604_31906 , RIdeb53e8_526, \9267_9566 );
and \U$22818 ( \31605_31907 , RIde989f0_334, \9269_9568 );
and \U$22819 ( \31606_31908 , RIe16eff0_2640, \9271_9570 );
and \U$22820 ( \31607_31909 , RIe15ade8_2411, \9273_9572 );
and \U$22821 ( \31608_31910 , RIe1445e8_2155, \9275_9574 );
and \U$22822 ( \31609_31911 , RIdf38fe0_2025, \9277_9576 );
and \U$22823 ( \31610_31912 , RIdf2d640_1893, \9279_9578 );
and \U$22824 ( \31611_31913 , RIdf1dec0_1717, \9281_9580 );
and \U$22825 ( \31612_31914 , RIdf015b8_1392, \9283_9582 );
and \U$22826 ( \31613_31915 , RIdee80b8_1104, \9285_9584 );
and \U$22827 ( \31614_31916 , RIdedce20_977, \9287_9586 );
and \U$22828 ( \31615_31917 , RIde7e938_207, \9289_9588 );
or \U$22829 ( \31616_31918 , \31552_31854 , \31553_31855 , \31554_31856 , \31555_31857 , \31556_31858 , \31557_31859 , \31558_31860 , \31559_31861 , \31560_31862 , \31561_31863 , \31562_31864 , \31563_31865 , \31564_31866 , \31565_31867 , \31566_31868 , \31567_31869 , \31568_31870 , \31569_31871 , \31570_31872 , \31571_31873 , \31572_31874 , \31573_31875 , \31574_31876 , \31575_31877 , \31576_31878 , \31577_31879 , \31578_31880 , \31579_31881 , \31580_31882 , \31581_31883 , \31582_31884 , \31583_31885 , \31584_31886 , \31585_31887 , \31586_31888 , \31587_31889 , \31588_31890 , \31589_31891 , \31590_31892 , \31591_31893 , \31592_31894 , \31593_31895 , \31594_31896 , \31595_31897 , \31596_31898 , \31597_31899 , \31598_31900 , \31599_31901 , \31600_31902 , \31601_31903 , \31602_31904 , \31603_31905 , \31604_31906 , \31605_31907 , \31606_31908 , \31607_31909 , \31608_31910 , \31609_31911 , \31610_31912 , \31611_31913 , \31612_31914 , \31613_31915 , \31614_31916 , \31615_31917 );
or \U$22830 ( \31617_31919 , \31551_31853 , \31616_31918 );
_DC \g65d1/U$1 ( \31618 , \31617_31919 , \9298_9597 );
and \U$22831 ( \31619_31921 , RIe19e480_3178, \8760_9059 );
and \U$22832 ( \31620_31922 , RIe19b780_3146, \8762_9061 );
and \U$22833 ( \31621_31923 , RIfccc980_7350, \8764_9063 );
and \U$22834 ( \31622_31924 , RIe198a80_3114, \8766_9065 );
and \U$22835 ( \31623_31925 , RIfcc1148_7219, \8768_9067 );
and \U$22836 ( \31624_31926 , RIe195d80_3082, \8770_9069 );
and \U$22837 ( \31625_31927 , RIe193080_3050, \8772_9071 );
and \U$22838 ( \31626_31928 , RIe190380_3018, \8774_9073 );
and \U$22839 ( \31627_31929 , RIe18a980_2954, \8776_9075 );
and \U$22840 ( \31628_31930 , RIe187c80_2922, \8778_9077 );
and \U$22841 ( \31629_31931 , RIfcb2ee0_7058, \8780_9079 );
and \U$22842 ( \31630_31932 , RIe184f80_2890, \8782_9081 );
and \U$22843 ( \31631_31933 , RIfc615e0_6130, \8784_9083 );
and \U$22844 ( \31632_31934 , RIe182280_2858, \8786_9085 );
and \U$22845 ( \31633_31935 , RIe17f580_2826, \8788_9087 );
and \U$22846 ( \31634_31936 , RIe17c880_2794, \8790_9089 );
and \U$22847 ( \31635_31937 , RIfc69038_6217, \8792_9091 );
and \U$22848 ( \31636_31938 , RIfc4c898_5893, \8794_9093 );
and \U$22849 ( \31637_31939 , RIfc6f2a8_6287, \8796_9095 );
and \U$22850 ( \31638_31940 , RIe1764a8_2723, \8798_9097 );
and \U$22851 ( \31639_31941 , RIfcad0a8_6991, \8800_9099 );
and \U$22852 ( \31640_31942 , RIfc6adc0_6238, \8802_9101 );
and \U$22853 ( \31641_31943 , RIfc70388_6299, \8804_9103 );
and \U$22854 ( \31642_31944 , RIfea1b50_8184, \8806_9105 );
and \U$22855 ( \31643_31945 , RIfea1f88_8187, \8808_9107 );
and \U$22856 ( \31644_31946 , RIfc56e88_6011, \8810_9109 );
and \U$22857 ( \31645_31947 , RIfea1cb8_8185, \8812_9111 );
and \U$22858 ( \31646_31948 , RIe174450_2700, \8814_9113 );
and \U$22859 ( \31647_31949 , RIfc60d70_6124, \8816_9115 );
and \U$22860 ( \31648_31950 , RIfc6a820_6234, \8818_9117 );
and \U$22861 ( \31649_31951 , RIfea1e20_8186, \8820_9119 );
and \U$22862 ( \31650_31952 , RIf16d798_5705, \8822_9121 );
and \U$22863 ( \31651_31953 , RIfc40bb0_5762, \8824_9123 );
and \U$22864 ( \31652_31954 , RIe2247d8_4705, \8826_9125 );
and \U$22865 ( \31653_31955 , RIfc77138_6377, \8828_9127 );
and \U$22866 ( \31654_31956 , RIe221ad8_4673, \8830_9129 );
and \U$22867 ( \31655_31957 , RIfcd7d80_7478, \8832_9131 );
and \U$22868 ( \31656_31958 , RIe21edd8_4641, \8834_9133 );
and \U$22869 ( \31657_31959 , RIe2193d8_4577, \8836_9135 );
and \U$22870 ( \31658_31960 , RIe2166d8_4545, \8838_9137 );
and \U$22871 ( \31659_31961 , RIfc40070_5754, \8840_9139 );
and \U$22872 ( \31660_31962 , RIe2139d8_4513, \8842_9141 );
and \U$22873 ( \31661_31963 , RIf169850_5660, \8844_9143 );
and \U$22874 ( \31662_31964 , RIe210cd8_4481, \8846_9145 );
and \U$22875 ( \31663_31965 , RIfcc1580_7222, \8848_9147 );
and \U$22876 ( \31664_31966 , RIe20dfd8_4449, \8850_9149 );
and \U$22877 ( \31665_31967 , RIe20b2d8_4417, \8852_9151 );
and \U$22878 ( \31666_31968 , RIe2085d8_4385, \8854_9153 );
and \U$22879 ( \31667_31969 , RIfcd0058_7389, \8856_9155 );
and \U$22880 ( \31668_31970 , RIfc749d8_6349, \8858_9157 );
and \U$22881 ( \31669_31971 , RIe203010_4324, \8860_9159 );
and \U$22882 ( \31670_31972 , RIe2013f0_4304, \8862_9161 );
and \U$22883 ( \31671_31973 , RIfc60230_6116, \8864_9163 );
and \U$22884 ( \31672_31974 , RIfc60668_6119, \8866_9165 );
and \U$22885 ( \31673_31975 , RIfcaf970_7020, \8868_9167 );
and \U$22886 ( \31674_31976 , RIfc45818_5813, \8870_9169 );
and \U$22887 ( \31675_31977 , RIf160a48_5559, \8872_9171 );
and \U$22888 ( \31676_31978 , RIf15eb58_5537, \8874_9173 );
and \U$22889 ( \31677_31979 , RIfea1880_8182, \8876_9175 );
and \U$22890 ( \31678_31980 , RIfea19e8_8183, \8878_9177 );
and \U$22891 ( \31679_31981 , RIfc72110_6320, \8880_9179 );
and \U$22892 ( \31680_31982 , RIfc49b98_5861, \8882_9181 );
and \U$22893 ( \31681_31983 , RIfcca0b8_7321, \8884_9183 );
and \U$22894 ( \31682_31984 , RIfc71738_6313, \8886_9185 );
or \U$22895 ( \31683_31985 , \31619_31921 , \31620_31922 , \31621_31923 , \31622_31924 , \31623_31925 , \31624_31926 , \31625_31927 , \31626_31928 , \31627_31929 , \31628_31930 , \31629_31931 , \31630_31932 , \31631_31933 , \31632_31934 , \31633_31935 , \31634_31936 , \31635_31937 , \31636_31938 , \31637_31939 , \31638_31940 , \31639_31941 , \31640_31942 , \31641_31943 , \31642_31944 , \31643_31945 , \31644_31946 , \31645_31947 , \31646_31948 , \31647_31949 , \31648_31950 , \31649_31951 , \31650_31952 , \31651_31953 , \31652_31954 , \31653_31955 , \31654_31956 , \31655_31957 , \31656_31958 , \31657_31959 , \31658_31960 , \31659_31961 , \31660_31962 , \31661_31963 , \31662_31964 , \31663_31965 , \31664_31966 , \31665_31967 , \31666_31968 , \31667_31969 , \31668_31970 , \31669_31971 , \31670_31972 , \31671_31973 , \31672_31974 , \31673_31975 , \31674_31976 , \31675_31977 , \31676_31978 , \31677_31979 , \31678_31980 , \31679_31981 , \31680_31982 , \31681_31983 , \31682_31984 );
and \U$22896 ( \31684_31986 , RIfc4ca00_5894, \8889_9188 );
and \U$22897 ( \31685_31987 , RIfc71030_6308, \8891_9190 );
and \U$22898 ( \31686_31988 , RIfcde428_7551, \8893_9192 );
and \U$22899 ( \31687_31989 , RIe1fad48_4231, \8895_9194 );
and \U$22900 ( \31688_31990 , RIfc70bf8_6305, \8897_9196 );
and \U$22901 ( \31689_31991 , RIfc63a70_6156, \8899_9198 );
and \U$22902 ( \31690_31992 , RIfca7db0_6932, \8901_9200 );
and \U$22903 ( \31691_31993 , RIe1f62c0_4178, \8903_9202 );
and \U$22904 ( \31692_31994 , RIfcada80_6998, \8905_9204 );
and \U$22905 ( \31693_31995 , RIfc6fde8_6295, \8907_9206 );
and \U$22906 ( \31694_31996 , RIfc6f578_6289, \8909_9208 );
and \U$22907 ( \31695_31997 , RIe1f3f98_4153, \8911_9210 );
and \U$22908 ( \31696_31998 , RIfcde158_7549, \8913_9212 );
and \U$22909 ( \31697_31999 , RIfcad378_6993, \8915_9214 );
and \U$22910 ( \31698_32000 , RIfc65f00_6182, \8917_9216 );
and \U$22911 ( \31699_32001 , RIe1eeca0_4094, \8919_9218 );
and \U$22912 ( \31700_32002 , RIe1ec540_4066, \8921_9220 );
and \U$22913 ( \31701_32003 , RIe1e9840_4034, \8923_9222 );
and \U$22914 ( \31702_32004 , RIe1e6b40_4002, \8925_9224 );
and \U$22915 ( \31703_32005 , RIe1e3e40_3970, \8927_9226 );
and \U$22916 ( \31704_32006 , RIe1e1140_3938, \8929_9228 );
and \U$22917 ( \31705_32007 , RIe1de440_3906, \8931_9230 );
and \U$22918 ( \31706_32008 , RIe1db740_3874, \8933_9232 );
and \U$22919 ( \31707_32009 , RIe1d8a40_3842, \8935_9234 );
and \U$22920 ( \31708_32010 , RIe1d3040_3778, \8937_9236 );
and \U$22921 ( \31709_32011 , RIe1d0340_3746, \8939_9238 );
and \U$22922 ( \31710_32012 , RIe1cd640_3714, \8941_9240 );
and \U$22923 ( \31711_32013 , RIe1ca940_3682, \8943_9242 );
and \U$22924 ( \31712_32014 , RIe1c7c40_3650, \8945_9244 );
and \U$22925 ( \31713_32015 , RIe1c4f40_3618, \8947_9246 );
and \U$22926 ( \31714_32016 , RIe1c2240_3586, \8949_9248 );
and \U$22927 ( \31715_32017 , RIe1bf540_3554, \8951_9250 );
and \U$22928 ( \31716_32018 , RIfc69308_6219, \8953_9252 );
and \U$22929 ( \31717_32019 , RIfccba08_7339, \8955_9254 );
and \U$22930 ( \31718_32020 , RIe1b9f78_3493, \8957_9256 );
and \U$22931 ( \31719_32021 , RIe1b7db8_3469, \8959_9258 );
and \U$22932 ( \31720_32022 , RIfccd628_7359, \8961_9260 );
and \U$22933 ( \31721_32023 , RIfc69740_6222, \8963_9262 );
and \U$22934 ( \31722_32024 , RIe1b5bf8_3445, \8965_9264 );
and \U$22935 ( \31723_32025 , RIe1b4578_3429, \8967_9266 );
and \U$22936 ( \31724_32026 , RIfccf950_7384, \8969_9268 );
and \U$22937 ( \31725_32027 , RIf148088_5279, \8971_9270 );
and \U$22938 ( \31726_32028 , RIe1b3060_3414, \8973_9272 );
and \U$22939 ( \31727_32029 , RIe1b1710_3396, \8975_9274 );
and \U$22940 ( \31728_32030 , RIfc9f818_6837, \8977_9276 );
and \U$22941 ( \31729_32031 , RIfcb9c90_7136, \8979_9278 );
and \U$22942 ( \31730_32032 , RIe1acf58_3345, \8981_9280 );
and \U$22943 ( \31731_32033 , RIe1ab770_3328, \8983_9282 );
and \U$22944 ( \31732_32034 , RIe1a9880_3306, \8985_9284 );
and \U$22945 ( \31733_32035 , RIe1a6b80_3274, \8987_9286 );
and \U$22946 ( \31734_32036 , RIe1a3e80_3242, \8989_9288 );
and \U$22947 ( \31735_32037 , RIe1a1180_3210, \8991_9290 );
and \U$22948 ( \31736_32038 , RIe18d680_2986, \8993_9292 );
and \U$22949 ( \31737_32039 , RIe179b80_2762, \8995_9294 );
and \U$22950 ( \31738_32040 , RIe2274d8_4737, \8997_9296 );
and \U$22951 ( \31739_32041 , RIe21c0d8_4609, \8999_9298 );
and \U$22952 ( \31740_32042 , RIe2058d8_4353, \9001_9300 );
and \U$22953 ( \31741_32043 , RIe1ff938_4285, \9003_9302 );
and \U$22954 ( \31742_32044 , RIe1f8cf0_4208, \9005_9304 );
and \U$22955 ( \31743_32045 , RIe1f1838_4125, \9007_9306 );
and \U$22956 ( \31744_32046 , RIe1d5d40_3810, \9009_9308 );
and \U$22957 ( \31745_32047 , RIe1bc840_3522, \9011_9310 );
and \U$22958 ( \31746_32048 , RIe1af6b8_3373, \9013_9312 );
and \U$22959 ( \31747_32049 , RIe171cf0_2672, \9015_9314 );
or \U$22960 ( \31748_32050 , \31684_31986 , \31685_31987 , \31686_31988 , \31687_31989 , \31688_31990 , \31689_31991 , \31690_31992 , \31691_31993 , \31692_31994 , \31693_31995 , \31694_31996 , \31695_31997 , \31696_31998 , \31697_31999 , \31698_32000 , \31699_32001 , \31700_32002 , \31701_32003 , \31702_32004 , \31703_32005 , \31704_32006 , \31705_32007 , \31706_32008 , \31707_32009 , \31708_32010 , \31709_32011 , \31710_32012 , \31711_32013 , \31712_32014 , \31713_32015 , \31714_32016 , \31715_32017 , \31716_32018 , \31717_32019 , \31718_32020 , \31719_32021 , \31720_32022 , \31721_32023 , \31722_32024 , \31723_32025 , \31724_32026 , \31725_32027 , \31726_32028 , \31727_32029 , \31728_32030 , \31729_32031 , \31730_32032 , \31731_32033 , \31732_32034 , \31733_32035 , \31734_32036 , \31735_32037 , \31736_32038 , \31737_32039 , \31738_32040 , \31739_32041 , \31740_32042 , \31741_32043 , \31742_32044 , \31743_32045 , \31744_32046 , \31745_32047 , \31746_32048 , \31747_32049 );
or \U$22961 ( \31749_32051 , \31683_31985 , \31748_32050 );
_DC \g65d2/U$1 ( \31750 , \31749_32051 , \9024_9323 );
and g65d3_GF_PartitionCandidate( \31751_32053_nG65d3 , \31618 , \31750 );
buf \U$22962 ( \31752_32054 , \31751_32053_nG65d3 );
and \U$22963 ( \31753_32055 , \31752_32054 , \10389_10691 );
nor \U$22964 ( \31754_32056 , \31486_31788 , \31753_32055 );
xnor \U$22965 ( \31755_32057 , \31754_32056 , \10678_10980 );
and \U$22966 ( \31756_32058 , \28782_29084 , \11275_11574 );
and \U$22967 ( \31757_32059 , \29966_30268 , \10976_11278 );
nor \U$22968 ( \31758_32060 , \31756_32058 , \31757_32059 );
xnor \U$22969 ( \31759_32061 , \31758_32060 , \11281_11580 );
xor \U$22970 ( \31760_32062 , \31755_32057 , \31759_32061 );
_DC \g63e8/U$1 ( \31761 , \31617_31919 , \9298_9597 );
_DC \g646c/U$1 ( \31762 , \31749_32051 , \9024_9323 );
xor g646d_GF_PartitionCandidate( \31763_32065_nG646d , \31761 , \31762 );
buf \U$22971 ( \31764_32066 , \31763_32065_nG646d );
xor \U$22972 ( \31765_32067 , \31764_32066 , \30508_30810 );
and \U$22973 ( \31766_32068 , \10385_10687 , \31765_32067 );
xor \U$22974 ( \31767_32069 , \31760_32062 , \31766_32068 );
xor \U$22975 ( \31768_32070 , \31485_31787 , \31767_32069 );
and \U$22976 ( \31769_32071 , \27011_27313 , \12491_12790 );
and \U$22977 ( \31770_32072 , \28232_28534 , \12159_12461 );
nor \U$22978 ( \31771_32073 , \31769_32071 , \31770_32072 );
xnor \U$22979 ( \31772_32074 , \31771_32073 , \12481_12780 );
and \U$22980 ( \31773_32075 , \22257_22556 , \16333_16635 );
and \U$22981 ( \31774_32076 , \23315_23617 , \15999_16301 );
nor \U$22982 ( \31775_32077 , \31773_32075 , \31774_32076 );
xnor \U$22983 ( \31776_32078 , \31775_32077 , \16323_16625 );
xor \U$22984 ( \31777_32079 , \31772_32074 , \31776_32078 );
and \U$22985 ( \31778_32080 , \13725_14024 , \25527_25826 );
and \U$22986 ( \31779_32081 , \14648_14950 , \24962_25264 );
nor \U$22987 ( \31780_32082 , \31778_32080 , \31779_32081 );
xnor \U$22988 ( \31781_32083 , \31780_32082 , \25474_25773 );
xor \U$22989 ( \31782_32084 , \31777_32079 , \31781_32083 );
xor \U$22990 ( \31783_32085 , \31768_32070 , \31782_32084 );
xor \U$22991 ( \31784_32086 , \31471_31773 , \31783_32085 );
xor \U$22992 ( \31785_32087 , \31462_31764 , \31784_32086 );
and \U$22993 ( \31786_32088 , \30576_30878 , \30580_30882 );
and \U$22994 ( \31787_32089 , \30580_30882 , \30625_30927 );
and \U$22995 ( \31788_32090 , \30576_30878 , \30625_30927 );
or \U$22996 ( \31789_32091 , \31786_32088 , \31787_32089 , \31788_32090 );
and \U$22997 ( \31790_32092 , \30535_30837 , \30539_30841 );
and \U$22998 ( \31791_32093 , \30539_30841 , \30544_30846 );
and \U$22999 ( \31792_32094 , \30535_30837 , \30544_30846 );
or \U$23000 ( \31793_32095 , \31790_32092 , \31791_32093 , \31792_32094 );
and \U$23001 ( \31794_32096 , \30595_30897 , \30609_30911 );
and \U$23002 ( \31795_32097 , \30609_30911 , \30624_30926 );
and \U$23003 ( \31796_32098 , \30595_30897 , \30624_30926 );
or \U$23004 ( \31797_32099 , \31794_32096 , \31795_32097 , \31796_32098 );
xor \U$23005 ( \31798_32100 , \31793_32095 , \31797_32099 );
and \U$23006 ( \31799_32101 , \30559_30861 , \30563_30865 );
and \U$23007 ( \31800_32102 , \30563_30865 , \30568_30870 );
and \U$23008 ( \31801_32103 , \30559_30861 , \30568_30870 );
or \U$23009 ( \31802_32104 , \31799_32101 , \31800_32102 , \31801_32103 );
and \U$23010 ( \31803_32105 , \30503_30805 , \30512_30814 );
xor \U$23011 ( \31804_32106 , \31802_32104 , \31803_32105 );
and \U$23012 ( \31805_32107 , \10686_10988 , \30521_30823 );
and \U$23013 ( \31806_32108 , \10968_11270 , \29944_30246 );
nor \U$23014 ( \31807_32109 , \31805_32107 , \31806_32108 );
xnor \U$23015 ( \31808_32110 , \31807_32109 , \30511_30813 );
xor \U$23016 ( \31809_32111 , \31804_32106 , \31808_32110 );
xor \U$23017 ( \31810_32112 , \31798_32100 , \31809_32111 );
xor \U$23018 ( \31811_32113 , \31789_32091 , \31810_32112 );
and \U$23019 ( \31812_32114 , \30550_30852 , \30554_30856 );
and \U$23020 ( \31813_32115 , \30554_30856 , \30569_30871 );
and \U$23021 ( \31814_32116 , \30550_30852 , \30569_30871 );
or \U$23022 ( \31815_32117 , \31812_32114 , \31813_32115 , \31814_32116 );
and \U$23023 ( \31816_32118 , \30585_30887 , \30589_30891 );
and \U$23024 ( \31817_32119 , \30589_30891 , \30594_30896 );
and \U$23025 ( \31818_32120 , \30585_30887 , \30594_30896 );
or \U$23026 ( \31819_32121 , \31816_32118 , \31817_32119 , \31818_32120 );
and \U$23027 ( \31820_32122 , \30599_30901 , \30603_30905 );
and \U$23028 ( \31821_32123 , \30603_30905 , \30608_30910 );
and \U$23029 ( \31822_32124 , \30599_30901 , \30608_30910 );
or \U$23030 ( \31823_32125 , \31820_32122 , \31821_32123 , \31822_32124 );
xor \U$23031 ( \31824_32126 , \31819_32121 , \31823_32125 );
and \U$23032 ( \31825_32127 , \30614_30916 , \30618_30920 );
and \U$23033 ( \31826_32128 , \30618_30920 , \30623_30925 );
and \U$23034 ( \31827_32129 , \30614_30916 , \30623_30925 );
or \U$23035 ( \31828_32130 , \31825_32127 , \31826_32128 , \31827_32129 );
xor \U$23036 ( \31829_32131 , \31824_32126 , \31828_32130 );
xor \U$23037 ( \31830_32132 , \31815_32117 , \31829_32131 );
and \U$23038 ( \31831_32133 , \30513_30815 , \30517_30819 );
and \U$23039 ( \31832_32134 , \30517_30819 , \30525_30827 );
and \U$23040 ( \31833_32135 , \30513_30815 , \30525_30827 );
or \U$23041 ( \31834_32136 , \31831_32133 , \31832_32134 , \31833_32135 );
and \U$23042 ( \31835_32137 , \23900_24199 , \15037_15336 );
and \U$23043 ( \31836_32138 , \24970_25272 , \14661_14963 );
nor \U$23044 ( \31837_32139 , \31835_32137 , \31836_32138 );
xnor \U$23045 ( \31838_32140 , \31837_32139 , \15043_15342 );
and \U$23046 ( \31839_32141 , \16353_16655 , \22243_22542 );
and \U$23047 ( \31840_32142 , \17325_17627 , \21801_22103 );
nor \U$23048 ( \31841_32143 , \31839_32141 , \31840_32142 );
xnor \U$23049 ( \31842_32144 , \31841_32143 , \22249_22548 );
xor \U$23050 ( \31843_32145 , \31838_32140 , \31842_32144 );
and \U$23051 ( \31844_32146 , \15022_15321 , \23839_24138 );
and \U$23052 ( \31845_32147 , \15965_16267 , \23328_23630 );
nor \U$23053 ( \31846_32148 , \31844_32146 , \31845_32147 );
xnor \U$23054 ( \31847_32149 , \31846_32148 , \23845_24144 );
xor \U$23055 ( \31848_32150 , \31843_32145 , \31847_32149 );
xor \U$23056 ( \31849_32151 , \31834_32136 , \31848_32150 );
and \U$23057 ( \31850_32152 , \25516_25815 , \13755_14054 );
and \U$23058 ( \31851_32153 , \26527_26829 , \13390_13692 );
nor \U$23059 ( \31852_32154 , \31850_32152 , \31851_32153 );
xnor \U$23060 ( \31853_32155 , \31852_32154 , \13736_14035 );
and \U$23061 ( \31854_32156 , \19259_19558 , \19235_19534 );
and \U$23062 ( \31855_32157 , \20242_20544 , \18743_19045 );
nor \U$23063 ( \31856_32158 , \31854_32156 , \31855_32157 );
xnor \U$23064 ( \31857_32159 , \31856_32158 , \19241_19540 );
xor \U$23065 ( \31858_32160 , \31853_32155 , \31857_32159 );
and \U$23066 ( \31859_32161 , \17736_18035 , \20706_21005 );
and \U$23067 ( \31860_32162 , \18730_19032 , \20255_20557 );
nor \U$23068 ( \31861_32163 , \31859_32161 , \31860_32162 );
xnor \U$23069 ( \31862_32164 , \31861_32163 , \20712_21011 );
xor \U$23070 ( \31863_32165 , \31858_32160 , \31862_32164 );
xor \U$23071 ( \31864_32166 , \31849_32151 , \31863_32165 );
xor \U$23072 ( \31865_32167 , \31830_32132 , \31864_32166 );
xor \U$23073 ( \31866_32168 , \31811_32113 , \31865_32167 );
xor \U$23074 ( \31867_32169 , \31785_32087 , \31866_32168 );
and \U$23075 ( \31868_32170 , \30219_30521 , \30223_30525 );
and \U$23076 ( \31869_32171 , \30223_30525 , \30627_30929 );
and \U$23077 ( \31870_32172 , \30219_30521 , \30627_30929 );
or \U$23078 ( \31871_32173 , \31868_32170 , \31869_32171 , \31870_32172 );
xor \U$23079 ( \31872_32174 , \31867_32169 , \31871_32173 );
and \U$23080 ( \31873_32175 , \30628_30930 , \30632_30934 );
and \U$23081 ( \31874_32176 , \30633_30935 , \30636_30938 );
or \U$23082 ( \31875_32177 , \31873_32175 , \31874_32176 );
xor \U$23083 ( \31876_32178 , \31872_32174 , \31875_32177 );
buf g9bb4_GF_PartitionCandidate( \31877_32179_nG9bb4 , \31876_32178 );
and \U$23084 ( \31878_32180 , \10402_10704 , \31877_32179_nG9bb4 );
or \U$23085 ( \31879_32181 , \31458_31760 , \31878_32180 );
xor \U$23086 ( \31880_32182 , \10399_10703 , \31879_32181 );
buf \U$23087 ( \31881_32183 , \31880_32182 );
buf \U$23089 ( \31882_32184 , \31881_32183 );
xor \U$23090 ( \31883_32185 , \31457_31759 , \31882_32184 );
buf \U$23091 ( \31884_32186 , \31883_32185 );
xor \U$23092 ( \31885_32187 , \31405_31707 , \31884_32186 );
buf \U$23093 ( \31886_32188 , \31885_32187 );
xor \U$23094 ( \31887_32189 , \31351_31653 , \31886_32188 );
and \U$23095 ( \31888_32190 , \30752_31051 , \30757_31056 );
and \U$23096 ( \31889_32191 , \30752_31051 , \30763_31062 );
and \U$23097 ( \31890_32192 , \30757_31056 , \30763_31062 );
or \U$23098 ( \31891_32193 , \31888_32190 , \31889_32191 , \31890_32192 );
buf \U$23099 ( \31892_32194 , \31891_32193 );
and \U$23100 ( \31893_32195 , \30208_30510 , \30213_30515 );
and \U$23101 ( \31894_32196 , \30208_30510 , \30643_30945 );
and \U$23102 ( \31895_32197 , \30213_30515 , \30643_30945 );
or \U$23103 ( \31896_32198 , \31893_32195 , \31894_32196 , \31895_32197 );
buf \U$23104 ( \31897_32199 , \31896_32198 );
xor \U$23105 ( \31898_32200 , \31892_32194 , \31897_32199 );
and \U$23106 ( \31899_32201 , \30168_30470 , \30185_30487 );
and \U$23107 ( \31900_32202 , \30168_30470 , \30192_30494 );
and \U$23108 ( \31901_32203 , \30185_30487 , \30192_30494 );
or \U$23109 ( \31902_32204 , \31899_32201 , \31900_32202 , \31901_32203 );
buf \U$23110 ( \31903_32205 , \31902_32204 );
and \U$23111 ( \31904_32206 , \30656_30958 , \30685_30984 );
and \U$23112 ( \31905_32207 , \30656_30958 , \30692_30991 );
and \U$23113 ( \31906_32208 , \30685_30984 , \30692_30991 );
or \U$23114 ( \31907_32209 , \31904_32206 , \31905_32207 , \31906_32208 );
buf \U$23115 ( \31908_32210 , \31907_32209 );
xor \U$23116 ( \31909_32211 , \31903_32205 , \31908_32210 );
and \U$23117 ( \31910_32212 , \30667_30969 , \30676_30975 );
and \U$23118 ( \31911_32213 , \30667_30969 , \30683_30982 );
and \U$23119 ( \31912_32214 , \30676_30975 , \30683_30982 );
or \U$23120 ( \31913_32215 , \31910_32212 , \31911_32213 , \31912_32214 );
buf \U$23121 ( \31914_32216 , \31913_32215 );
and \U$23122 ( \31915_32217 , \30670_29853 , \10693_10995_nG9c0b );
and \U$23123 ( \31916_32218 , \29551_29850 , \10981_11283_nG9c08 );
or \U$23124 ( \31917_32219 , \31915_32217 , \31916_32218 );
xor \U$23125 ( \31918_32220 , \29550_29849 , \31917_32219 );
buf \U$23126 ( \31919_32221 , \31918_32220 );
buf \U$23128 ( \31920_32222 , \31919_32221 );
and \U$23129 ( \31921_32223 , \28946_28118 , \11299_11598_nG9c05 );
and \U$23130 ( \31922_32224 , \27816_28115 , \12168_12470_nG9c02 );
or \U$23131 ( \31923_32225 , \31921_32223 , \31922_32224 );
xor \U$23132 ( \31924_32226 , \27815_28114 , \31923_32225 );
buf \U$23133 ( \31925_32227 , \31924_32226 );
buf \U$23135 ( \31926_32228 , \31925_32227 );
xor \U$23136 ( \31927_32229 , \31920_32222 , \31926_32228 );
buf \U$23137 ( \31928_32230 , \31927_32229 );
xor \U$23138 ( \31929_32231 , \31914_32216 , \31928_32230 );
and \U$23139 ( \31930_32232 , \23495_23201 , \15074_15373_nG9bf3 );
and \U$23140 ( \31931_32233 , \22899_23198 , \16013_16315_nG9bf0 );
or \U$23141 ( \31932_32234 , \31930_32232 , \31931_32233 );
xor \U$23142 ( \31933_32235 , \22898_23197 , \31932_32234 );
buf \U$23143 ( \31934_32236 , \31933_32235 );
buf \U$23145 ( \31935_32237 , \31934_32236 );
xor \U$23146 ( \31936_32238 , \31929_32231 , \31935_32237 );
buf \U$23147 ( \31937_32239 , \31936_32238 );
xor \U$23148 ( \31938_32240 , \31909_32211 , \31937_32239 );
buf \U$23149 ( \31939_32241 , \31938_32240 );
and \U$23150 ( \31940_32242 , \13431_13370 , \25561_25860_nG9bc9 );
and \U$23151 ( \31941_32243 , \13068_13367 , \26585_26887_nG9bc6 );
or \U$23152 ( \31942_32244 , \31940_32242 , \31941_32243 );
xor \U$23153 ( \31943_32245 , \13067_13366 , \31942_32244 );
buf \U$23154 ( \31944_32246 , \31943_32245 );
buf \U$23156 ( \31945_32247 , \31944_32246 );
xor \U$23157 ( \31946_32248 , \31939_32241 , \31945_32247 );
and \U$23158 ( \31947_32249 , \10996_10421 , \28877_29179_nG9bbd );
and \U$23159 ( \31948_32250 , \10119_10418 , \30064_30366_nG9bba );
or \U$23160 ( \31949_32251 , \31947_32249 , \31948_32250 );
xor \U$23161 ( \31950_32252 , \10118_10417 , \31949_32251 );
buf \U$23162 ( \31951_32253 , \31950_32252 );
buf \U$23164 ( \31952_32254 , \31951_32253 );
xor \U$23165 ( \31953_32255 , \31946_32248 , \31952_32254 );
buf \U$23166 ( \31954_32256 , \31953_32255 );
xor \U$23167 ( \31955_32257 , \31898_32200 , \31954_32256 );
buf \U$23168 ( \31956_32258 , \31955_32257 );
xor \U$23169 ( \31957_32259 , \31887_32189 , \31956_32258 );
and \U$23170 ( \31958_32260 , \31341_31643 , \31957_32259 );
and \U$23171 ( \31959_32261 , \31345_31647 , \31957_32259 );
or \U$23172 ( \31960_32262 , \31346_31648 , \31958_32260 , \31959_32261 );
and \U$23173 ( \31961_32263 , \30780_31079 , \30784_31083 );
and \U$23174 ( \31962_32264 , \30780_31079 , \31340_31642 );
and \U$23175 ( \31963_32265 , \30784_31083 , \31340_31642 );
or \U$23176 ( \31964_32266 , \31961_32263 , \31962_32264 , \31963_32265 );
xor \U$23177 ( \31965_32267 , \31960_32262 , \31964_32266 );
and \U$23178 ( \31966_32268 , \31892_32194 , \31897_32199 );
and \U$23179 ( \31967_32269 , \31892_32194 , \31954_32256 );
and \U$23180 ( \31968_32270 , \31897_32199 , \31954_32256 );
or \U$23181 ( \31969_32271 , \31966_32268 , \31967_32269 , \31968_32270 );
buf \U$23182 ( \31970_32272 , \31969_32271 );
and \U$23183 ( \31971_32273 , \31417_31719 , \31423_31725 );
and \U$23184 ( \31972_32274 , \31417_31719 , \31430_31732 );
and \U$23185 ( \31973_32275 , \31423_31725 , \31430_31732 );
or \U$23186 ( \31974_32276 , \31971_32273 , \31972_32274 , \31973_32275 );
buf \U$23187 ( \31975_32277 , \31974_32276 );
and \U$23188 ( \31976_32278 , \31333_31632 , \31337_31639 );
buf \U$23189 ( \31977_32279 , \31976_32278 );
buf \U$23191 ( \31978_32280 , \31977_32279 );
and \U$23192 ( \31979_32281 , \30670_29853 , \10981_11283_nG9c08 );
and \U$23193 ( \31980_32282 , \29551_29850 , \11299_11598_nG9c05 );
or \U$23194 ( \31981_32283 , \31979_32281 , \31980_32282 );
xor \U$23195 ( \31982_32284 , \29550_29849 , \31981_32283 );
buf \U$23196 ( \31983_32285 , \31982_32284 );
buf \U$23198 ( \31984_32286 , \31983_32285 );
xor \U$23199 ( \31985_32287 , \31978_32280 , \31984_32286 );
buf \U$23200 ( \31986_32288 , \31985_32287 );
not \U$22535 ( \31987_31634 , \31334_31633 );
xor \U$22536 ( \31988_31635 , \31328_31627_nG43fa , \31331_31630_nG43fd );
and \U$22537 ( \31989_31636 , \31987_31634 , \31988_31635 );
and \U$23201 ( \31990_32289 , \31989_31636 , \10392_10694_nG9c0e );
and \U$23202 ( \31991_32290 , \31334_31633 , \10693_10995_nG9c0b );
or \U$23203 ( \31992_32291 , \31990_32289 , \31991_32290 );
xor \U$23204 ( \31993_32292 , \31333_31632 , \31992_32291 );
buf \U$23205 ( \31994_32293 , \31993_32292 );
buf \U$23207 ( \31995_32294 , \31994_32293 );
xor \U$23208 ( \31996_32295 , \31986_32288 , \31995_32294 );
and \U$23209 ( \31997_32296 , \28946_28118 , \12168_12470_nG9c02 );
and \U$23210 ( \31998_32297 , \27816_28115 , \12502_12801_nG9bff );
or \U$23211 ( \31999_32298 , \31997_32296 , \31998_32297 );
xor \U$23212 ( \32000_32299 , \27815_28114 , \31999_32298 );
buf \U$23213 ( \32001_32300 , \32000_32299 );
buf \U$23215 ( \32002_32301 , \32001_32300 );
xor \U$23216 ( \32003_32302 , \31996_32295 , \32002_32301 );
buf \U$23217 ( \32004_32303 , \32003_32302 );
xor \U$23218 ( \32005_32304 , \31975_32277 , \32004_32303 );
and \U$23219 ( \32006_32305 , \23495_23201 , \16013_16315_nG9bf0 );
and \U$23220 ( \32007_32306 , \22899_23198 , \16378_16680_nG9bed );
or \U$23221 ( \32008_32307 , \32006_32305 , \32007_32306 );
xor \U$23222 ( \32009_32308 , \22898_23197 , \32008_32307 );
buf \U$23223 ( \32010_32309 , \32009_32308 );
buf \U$23225 ( \32011_32310 , \32010_32309 );
xor \U$23226 ( \32012_32311 , \32005_32304 , \32011_32310 );
buf \U$23227 ( \32013_32312 , \32012_32311 );
and \U$23228 ( \32014_32313 , \20353_20155 , \18789_19091_nG9be4 );
and \U$23229 ( \32015_32314 , \19853_20152 , \19287_19586_nG9be1 );
or \U$23230 ( \32016_32315 , \32014_32313 , \32015_32314 );
xor \U$23231 ( \32017_32316 , \19852_20151 , \32016_32315 );
buf \U$23232 ( \32018_32317 , \32017_32316 );
buf \U$23234 ( \32019_32318 , \32018_32317 );
xor \U$23235 ( \32020_32319 , \32013_32312 , \32019_32318 );
and \U$23236 ( \32021_32320 , \18908_18702 , \20306_20608_nG9bde );
and \U$23237 ( \32022_32321 , \18400_18699 , \20787_21086_nG9bdb );
or \U$23238 ( \32023_32322 , \32021_32320 , \32022_32321 );
xor \U$23239 ( \32024_32323 , \18399_18698 , \32023_32322 );
buf \U$23240 ( \32025_32324 , \32024_32323 );
buf \U$23242 ( \32026_32325 , \32025_32324 );
xor \U$23243 ( \32027_32326 , \32020_32319 , \32026_32325 );
buf \U$23244 ( \32028_32327 , \32027_32326 );
and \U$23245 ( \32029_32328 , \13431_13370 , \26585_26887_nG9bc6 );
and \U$23246 ( \32030_32329 , \13068_13367 , \27114_27416_nG9bc3 );
or \U$23247 ( \32031_32330 , \32029_32328 , \32030_32329 );
xor \U$23248 ( \32032_32331 , \13067_13366 , \32031_32330 );
buf \U$23249 ( \32033_32332 , \32032_32331 );
buf \U$23251 ( \32034_32333 , \32033_32332 );
xor \U$23252 ( \32035_32334 , \32028_32327 , \32034_32333 );
and \U$23253 ( \32036_32335 , \12183_12157 , \28300_28602_nG9bc0 );
and \U$23254 ( \32037_32336 , \11855_12154 , \28877_29179_nG9bbd );
or \U$23255 ( \32038_32337 , \32036_32335 , \32037_32336 );
xor \U$23256 ( \32039_32338 , \11854_12153 , \32038_32337 );
buf \U$23257 ( \32040_32339 , \32039_32338 );
buf \U$23259 ( \32041_32340 , \32040_32339 );
xor \U$23260 ( \32042_32341 , \32035_32334 , \32041_32340 );
buf \U$23261 ( \32043_32342 , \32042_32341 );
and \U$23262 ( \32044_32343 , \31372_31674 , \31378_31680 );
and \U$23263 ( \32045_32344 , \31372_31674 , \31385_31687 );
and \U$23264 ( \32046_32345 , \31378_31680 , \31385_31687 );
or \U$23265 ( \32047_32346 , \32044_32343 , \32045_32344 , \32046_32345 );
buf \U$23266 ( \32048_32347 , \32047_32346 );
and \U$23267 ( \32049_32348 , \16405_15940 , \23394_23696_nG9bd2 );
and \U$23268 ( \32050_32349 , \15638_15937 , \23927_24226_nG9bcf );
or \U$23269 ( \32051_32350 , \32049_32348 , \32050_32349 );
xor \U$23270 ( \32052_32351 , \15637_15936 , \32051_32350 );
buf \U$23271 ( \32053_32352 , \32052_32351 );
buf \U$23273 ( \32054_32353 , \32053_32352 );
xor \U$23274 ( \32055_32354 , \32048_32347 , \32054_32353 );
and \U$23275 ( \32056_32355 , \14710_14631 , \24996_25298_nG9bcc );
and \U$23276 ( \32057_32356 , \14329_14628 , \25561_25860_nG9bc9 );
or \U$23277 ( \32058_32357 , \32056_32355 , \32057_32356 );
xor \U$23278 ( \32059_32358 , \14328_14627 , \32058_32357 );
buf \U$23279 ( \32060_32359 , \32059_32358 );
buf \U$23281 ( \32061_32360 , \32060_32359 );
xor \U$23282 ( \32062_32361 , \32055_32354 , \32061_32360 );
buf \U$23283 ( \32063_32362 , \32062_32361 );
xor \U$23284 ( \32064_32363 , \32043_32342 , \32063_32362 );
and \U$23285 ( \32065_32364 , \31939_32241 , \31945_32247 );
and \U$23286 ( \32066_32365 , \31939_32241 , \31952_32254 );
and \U$23287 ( \32067_32366 , \31945_32247 , \31952_32254 );
or \U$23288 ( \32068_32367 , \32065_32364 , \32066_32365 , \32067_32366 );
buf \U$23289 ( \32069_32368 , \32068_32367 );
xor \U$23290 ( \32070_32369 , \32064_32363 , \32069_32368 );
buf \U$23291 ( \32071_32370 , \32070_32369 );
xor \U$23292 ( \32072_32371 , \31970_32272 , \32071_32370 );
and \U$23293 ( \32073_32372 , \31361_31663 , \31396_31698 );
and \U$23294 ( \32074_32373 , \31361_31663 , \31402_31704 );
and \U$23295 ( \32075_32374 , \31396_31698 , \31402_31704 );
or \U$23296 ( \32076_32375 , \32073_32372 , \32074_32373 , \32075_32374 );
buf \U$23297 ( \32077_32376 , \32076_32375 );
xor \U$23298 ( \32078_32377 , \32072_32371 , \32077_32376 );
buf \U$23299 ( \32079_32378 , \32078_32377 );
and \U$23300 ( \32080_32379 , \31356_31658 , \31404_31706 );
and \U$23301 ( \32081_32380 , \31356_31658 , \31884_32186 );
and \U$23302 ( \32082_32381 , \31404_31706 , \31884_32186 );
or \U$23303 ( \32083_32382 , \32080_32379 , \32081_32380 , \32082_32381 );
buf \U$23304 ( \32084_32383 , \32083_32382 );
xor \U$23305 ( \32085_32384 , \32079_32378 , \32084_32383 );
and \U$23306 ( \32086_32385 , \31914_32216 , \31928_32230 );
and \U$23307 ( \32087_32386 , \31914_32216 , \31935_32237 );
and \U$23308 ( \32088_32387 , \31928_32230 , \31935_32237 );
or \U$23309 ( \32089_32388 , \32086_32385 , \32087_32386 , \32088_32387 );
buf \U$23310 ( \32090_32389 , \32089_32388 );
and \U$23311 ( \32091_32390 , \31920_32222 , \31926_32228 );
buf \U$23312 ( \32092_32391 , \32091_32390 );
and \U$23313 ( \32093_32392 , \27141_26431 , \13403_13705_nG9bfc );
and \U$23314 ( \32094_32393 , \26129_26428 , \13771_14070_nG9bf9 );
or \U$23315 ( \32095_32394 , \32093_32392 , \32094_32393 );
xor \U$23316 ( \32096_32395 , \26128_26427 , \32095_32394 );
buf \U$23317 ( \32097_32396 , \32096_32395 );
buf \U$23319 ( \32098_32397 , \32097_32396 );
xor \U$23320 ( \32099_32398 , \32092_32391 , \32098_32397 );
and \U$23321 ( \32100_32399 , \25044_24792 , \14682_14984_nG9bf6 );
and \U$23322 ( \32101_32400 , \24490_24789 , \15074_15373_nG9bf3 );
or \U$23323 ( \32102_32401 , \32100_32399 , \32101_32400 );
xor \U$23324 ( \32103_32402 , \24489_24788 , \32102_32401 );
buf \U$23325 ( \32104_32403 , \32103_32402 );
buf \U$23327 ( \32105_32404 , \32104_32403 );
xor \U$23328 ( \32106_32405 , \32099_32398 , \32105_32404 );
buf \U$23329 ( \32107_32406 , \32106_32405 );
xor \U$23330 ( \32108_32407 , \32090_32389 , \32107_32406 );
and \U$23331 ( \32109_32408 , \21908_21658 , \17363_17665_nG9bea );
and \U$23332 ( \32110_32409 , \21356_21655 , \17808_18107_nG9be7 );
or \U$23333 ( \32111_32410 , \32109_32408 , \32110_32409 );
xor \U$23334 ( \32112_32411 , \21355_21654 , \32111_32410 );
buf \U$23335 ( \32113_32412 , \32112_32411 );
buf \U$23337 ( \32114_32413 , \32113_32412 );
xor \U$23338 ( \32115_32414 , \32108_32407 , \32114_32413 );
buf \U$23339 ( \32116_32415 , \32115_32414 );
and \U$23340 ( \32117_32416 , \31415_31717 , \31432_31734 );
and \U$23341 ( \32118_32417 , \31415_31717 , \31439_31741 );
and \U$23342 ( \32119_32418 , \31432_31734 , \31439_31741 );
or \U$23343 ( \32120_32419 , \32117_32416 , \32118_32417 , \32119_32418 );
buf \U$23344 ( \32121_32420 , \32120_32419 );
xor \U$23345 ( \32122_32421 , \32116_32415 , \32121_32420 );
and \U$23346 ( \32123_32422 , \17437_17297 , \21827_22129_nG9bd8 );
and \U$23347 ( \32124_32423 , \16995_17294 , \22330_22629_nG9bd5 );
or \U$23348 ( \32125_32424 , \32123_32422 , \32124_32423 );
xor \U$23349 ( \32126_32425 , \16994_17293 , \32125_32424 );
buf \U$23350 ( \32127_32426 , \32126_32425 );
buf \U$23352 ( \32128_32427 , \32127_32426 );
xor \U$23353 ( \32129_32428 , \32122_32421 , \32128_32427 );
buf \U$23354 ( \32130_32429 , \32129_32428 );
and \U$23355 ( \32131_32430 , \31441_31743 , \31447_31749 );
and \U$23356 ( \32132_32431 , \31441_31743 , \31454_31756 );
and \U$23357 ( \32133_32432 , \31447_31749 , \31454_31756 );
or \U$23358 ( \32134_32433 , \32131_32430 , \32132_32431 , \32133_32432 );
buf \U$23359 ( \32135_32434 , \32134_32433 );
xor \U$23360 ( \32136_32435 , \32130_32429 , \32135_32434 );
and \U$23361 ( \32137_32436 , \31366_31668 , \31387_31689 );
and \U$23362 ( \32138_32437 , \31366_31668 , \31394_31696 );
and \U$23363 ( \32139_32438 , \31387_31689 , \31394_31696 );
or \U$23364 ( \32140_32439 , \32137_32436 , \32138_32437 , \32139_32438 );
buf \U$23365 ( \32141_32440 , \32140_32439 );
xor \U$23366 ( \32142_32441 , \32136_32435 , \32141_32440 );
buf \U$23367 ( \32143_32442 , \32142_32441 );
and \U$23368 ( \32144_32443 , \31903_32205 , \31908_32210 );
and \U$23369 ( \32145_32444 , \31903_32205 , \31937_32239 );
and \U$23370 ( \32146_32445 , \31908_32210 , \31937_32239 );
or \U$23371 ( \32147_32446 , \32144_32443 , \32145_32444 , \32146_32445 );
buf \U$23372 ( \32148_32447 , \32147_32446 );
and \U$23373 ( \32149_32448 , \10996_10421 , \30064_30366_nG9bba );
and \U$23374 ( \32150_32449 , \10119_10418 , \30638_30940_nG9bb7 );
or \U$23375 ( \32151_32450 , \32149_32448 , \32150_32449 );
xor \U$23376 ( \32152_32451 , \10118_10417 , \32151_32450 );
buf \U$23377 ( \32153_32452 , \32152_32451 );
buf \U$23379 ( \32154_32453 , \32153_32452 );
xor \U$23380 ( \32155_32454 , \32148_32447 , \32154_32453 );
and \U$23381 ( \32156_32455 , \10411_10707 , \31877_32179_nG9bb4 );
and \U$23382 ( \32157_32456 , \31789_32091 , \31810_32112 );
and \U$23383 ( \32158_32457 , \31810_32112 , \31865_32167 );
and \U$23384 ( \32159_32458 , \31789_32091 , \31865_32167 );
or \U$23385 ( \32160_32459 , \32157_32456 , \32158_32457 , \32159_32458 );
and \U$23386 ( \32161_32460 , \31793_32095 , \31797_32099 );
and \U$23387 ( \32162_32461 , \31797_32099 , \31809_32111 );
and \U$23388 ( \32163_32462 , \31793_32095 , \31809_32111 );
or \U$23389 ( \32164_32463 , \32161_32460 , \32162_32461 , \32163_32462 );
and \U$23390 ( \32165_32464 , \31815_32117 , \31829_32131 );
and \U$23391 ( \32166_32465 , \31829_32131 , \31864_32166 );
and \U$23392 ( \32167_32466 , \31815_32117 , \31864_32166 );
or \U$23393 ( \32168_32467 , \32165_32464 , \32166_32465 , \32167_32466 );
xor \U$23394 ( \32169_32468 , \32164_32463 , \32168_32467 );
and \U$23395 ( \32170_32469 , \31819_32121 , \31823_32125 );
and \U$23396 ( \32171_32470 , \31823_32125 , \31828_32130 );
and \U$23397 ( \32172_32471 , \31819_32121 , \31828_32130 );
or \U$23398 ( \32173_32472 , \32170_32469 , \32171_32470 , \32172_32471 );
and \U$23399 ( \32174_32473 , \23315_23617 , \16333_16635 );
and \U$23400 ( \32175_32474 , \23900_24199 , \15999_16301 );
nor \U$23401 ( \32176_32475 , \32174_32473 , \32175_32474 );
xnor \U$23402 ( \32177_32476 , \32176_32475 , \16323_16625 );
and \U$23403 ( \32178_32477 , \14648_14950 , \25527_25826 );
and \U$23404 ( \32179_32478 , \15022_15321 , \24962_25264 );
nor \U$23405 ( \32180_32479 , \32178_32477 , \32179_32478 );
xnor \U$23406 ( \32181_32480 , \32180_32479 , \25474_25773 );
xor \U$23407 ( \32182_32481 , \32177_32476 , \32181_32480 );
and \U$23408 ( \32183_32482 , \13377_13679 , \27095_27397 );
and \U$23409 ( \32184_32483 , \13725_14024 , \26505_26807 );
nor \U$23410 ( \32185_32484 , \32183_32482 , \32184_32483 );
xnor \U$23411 ( \32186_32485 , \32185_32484 , \26993_27295 );
xor \U$23412 ( \32187_32486 , \32182_32481 , \32186_32485 );
xor \U$23413 ( \32188_32487 , \32173_32472 , \32187_32486 );
and \U$23414 ( \32189_32488 , \28232_28534 , \12491_12790 );
and \U$23415 ( \32190_32489 , \28782_29084 , \12159_12461 );
nor \U$23416 ( \32191_32490 , \32189_32488 , \32190_32489 );
xnor \U$23417 ( \32192_32491 , \32191_32490 , \12481_12780 );
and \U$23418 ( \32193_32492 , \17325_17627 , \22243_22542 );
and \U$23419 ( \32194_32493 , \17736_18035 , \21801_22103 );
nor \U$23420 ( \32195_32494 , \32193_32492 , \32194_32493 );
xnor \U$23421 ( \32196_32495 , \32195_32494 , \22249_22548 );
xor \U$23422 ( \32197_32496 , \32192_32491 , \32196_32495 );
and \U$23423 ( \32198_32497 , \15965_16267 , \23839_24138 );
and \U$23424 ( \32199_32498 , \16353_16655 , \23328_23630 );
nor \U$23425 ( \32200_32499 , \32198_32497 , \32199_32498 );
xnor \U$23426 ( \32201_32500 , \32200_32499 , \23845_24144 );
xor \U$23427 ( \32202_32501 , \32197_32496 , \32201_32500 );
xor \U$23428 ( \32203_32502 , \32188_32487 , \32202_32501 );
xor \U$23429 ( \32204_32503 , \32169_32468 , \32203_32502 );
xor \U$23430 ( \32205_32504 , \32160_32459 , \32204_32503 );
and \U$23431 ( \32206_32505 , \31466_31768 , \31470_31772 );
and \U$23432 ( \32207_32506 , \31470_31772 , \31783_32085 );
and \U$23433 ( \32208_32507 , \31466_31768 , \31783_32085 );
or \U$23434 ( \32209_32508 , \32206_32505 , \32207_32506 , \32208_32507 );
and \U$23435 ( \32210_32509 , \31802_32104 , \31803_32105 );
and \U$23436 ( \32211_32510 , \31803_32105 , \31808_32110 );
and \U$23437 ( \32212_32511 , \31802_32104 , \31808_32110 );
or \U$23438 ( \32213_32512 , \32210_32509 , \32211_32510 , \32212_32511 );
and \U$23439 ( \32214_32513 , \31475_31777 , \31479_31781 );
and \U$23440 ( \32215_32514 , \31479_31781 , \31484_31786 );
and \U$23441 ( \32216_32515 , \31475_31777 , \31484_31786 );
or \U$23442 ( \32217_32516 , \32214_32513 , \32215_32514 , \32216_32515 );
and \U$23443 ( \32218_32517 , \31772_32074 , \31776_32078 );
and \U$23444 ( \32219_32518 , \31776_32078 , \31781_32083 );
and \U$23445 ( \32220_32519 , \31772_32074 , \31781_32083 );
or \U$23446 ( \32221_32520 , \32218_32517 , \32219_32518 , \32220_32519 );
xor \U$23447 ( \32222_32521 , \32217_32516 , \32221_32520 );
and \U$23448 ( \32223_32522 , \31838_32140 , \31842_32144 );
and \U$23449 ( \32224_32523 , \31842_32144 , \31847_32149 );
and \U$23450 ( \32225_32524 , \31838_32140 , \31847_32149 );
or \U$23451 ( \32226_32525 , \32223_32522 , \32224_32523 , \32225_32524 );
xor \U$23452 ( \32227_32526 , \32222_32521 , \32226_32525 );
xor \U$23453 ( \32228_32527 , \32213_32512 , \32227_32526 );
and \U$23454 ( \32229_32528 , \31752_32054 , \10681_10983 );
and \U$23455 ( \32230_32529 , RIdec6350_719, \9034_9333 );
and \U$23456 ( \32231_32530 , RIdec3650_687, \9036_9335 );
and \U$23457 ( \32232_32531 , RIfcaf3d0_7016, \9038_9337 );
and \U$23458 ( \32233_32532 , RIdec0950_655, \9040_9339 );
and \U$23459 ( \32234_32533 , RIfc6a280_6230, \9042_9341 );
and \U$23460 ( \32235_32534 , RIdebdc50_623, \9044_9343 );
and \U$23461 ( \32236_32535 , RIdebaf50_591, \9046_9345 );
and \U$23462 ( \32237_32536 , RIdeb8250_559, \9048_9347 );
and \U$23463 ( \32238_32537 , RIfc42f50_5784, \9050_9349 );
and \U$23464 ( \32239_32538 , RIdeb2850_495, \9052_9351 );
and \U$23465 ( \32240_32539 , RIfc981f8_6753, \9054_9353 );
and \U$23466 ( \32241_32540 , RIdeafb50_463, \9056_9355 );
and \U$23467 ( \32242_32541 , RIfc8c6f0_6620, \9058_9357 );
and \U$23468 ( \32243_32542 , RIdeac838_431, \9060_9359 );
and \U$23469 ( \32244_32543 , RIdea5f38_399, \9062_9361 );
and \U$23470 ( \32245_32544 , RIde9f638_367, \9064_9363 );
and \U$23471 ( \32246_32545 , RIee1d4e8_4792, \9066_9365 );
and \U$23472 ( \32247_32546 , RIfcda648_7507, \9068_9367 );
and \U$23473 ( \32248_32547 , RIfcc6440_7278, \9070_9369 );
and \U$23474 ( \32249_32548 , RIfcd5620_7450, \9072_9371 );
and \U$23475 ( \32250_32549 , RIde92ac8_305, \9074_9373 );
and \U$23476 ( \32251_32550 , RIfea34a0_8202, \9076_9375 );
and \U$23477 ( \32252_32551 , RIfea31d0_8200, \9078_9377 );
and \U$23478 ( \32253_32552 , RIfea3338_8201, \9080_9379 );
and \U$23479 ( \32254_32553 , RIfcb6b58_7101, \9082_9381 );
and \U$23480 ( \32255_32554 , RIfcb6888_7099, \9084_9383 );
and \U$23481 ( \32256_32555 , RIfc9dd60_6818, \9086_9385 );
and \U$23482 ( \32257_32556 , RIee19708_4748, \9088_9387 );
and \U$23483 ( \32258_32557 , RIfc50c18_5941, \9090_9389 );
and \U$23484 ( \32259_32558 , RIe16c458_2609, \9092_9391 );
and \U$23485 ( \32260_32559 , RIfc80a80_6486, \9094_9393 );
and \U$23486 ( \32261_32560 , RIfec62e8_8375, \9096_9395 );
and \U$23487 ( \32262_32561 , RIe166350_2540, \9098_9397 );
and \U$23488 ( \32263_32562 , RIe163650_2508, \9100_9399 );
and \U$23489 ( \32264_32563 , RIee37d98_5094, \9102_9401 );
and \U$23490 ( \32265_32564 , RIe160950_2476, \9104_9403 );
and \U$23491 ( \32266_32565 , RIfcaa678_6961, \9106_9405 );
and \U$23492 ( \32267_32566 , RIe15dc50_2444, \9108_9407 );
and \U$23493 ( \32268_32567 , RIe158250_2380, \9110_9409 );
and \U$23494 ( \32269_32568 , RIe155550_2348, \9112_9411 );
and \U$23495 ( \32270_32569 , RIfea3ba8_8207, \9114_9413 );
and \U$23496 ( \32271_32570 , RIe152850_2316, \9116_9415 );
and \U$23497 ( \32272_32571 , RIee35638_5066, \9118_9417 );
and \U$23498 ( \32273_32572 , RIe14fb50_2284, \9120_9419 );
and \U$23499 ( \32274_32573 , RIfc62f30_6148, \9122_9421 );
and \U$23500 ( \32275_32574 , RIe14ce50_2252, \9124_9423 );
and \U$23501 ( \32276_32575 , RIe14a150_2220, \9126_9425 );
and \U$23502 ( \32277_32576 , RIe147450_2188, \9128_9427 );
and \U$23503 ( \32278_32577 , RIfc97f28_6751, \9130_9429 );
and \U$23504 ( \32279_32578 , RIfc89888_6587, \9132_9431 );
and \U$23505 ( \32280_32579 , RIfc8f558_6653, \9134_9433 );
and \U$23506 ( \32281_32580 , RIfc52838_5961, \9136_9435 );
and \U$23507 ( \32282_32581 , RIe141bb8_2125, \9138_9437 );
and \U$23508 ( \32283_32582 , RIe13f890_2100, \9140_9439 );
and \U$23509 ( \32284_32583 , RIdf3d798_2076, \9142_9441 );
and \U$23510 ( \32285_32584 , RIdf3b308_2050, \9144_9443 );
and \U$23511 ( \32286_32585 , RIee30a48_5012, \9146_9445 );
and \U$23512 ( \32287_32586 , RIfc568e8_6007, \9148_9447 );
and \U$23513 ( \32288_32587 , RIee2e9f0_4989, \9150_9449 );
and \U$23514 ( \32289_32588 , RIee2dbe0_4979, \9152_9451 );
and \U$23515 ( \32290_32589 , RIdf365b0_1995, \9154_9453 );
and \U$23516 ( \32291_32590 , RIfea38d8_8205, \9156_9455 );
and \U$23517 ( \32292_32591 , RIfea3a40_8206, \9158_9457 );
and \U$23518 ( \32293_32592 , RIdf2ff08_1922, \9160_9459 );
or \U$23519 ( \32294_32593 , \32230_32529 , \32231_32530 , \32232_32531 , \32233_32532 , \32234_32533 , \32235_32534 , \32236_32535 , \32237_32536 , \32238_32537 , \32239_32538 , \32240_32539 , \32241_32540 , \32242_32541 , \32243_32542 , \32244_32543 , \32245_32544 , \32246_32545 , \32247_32546 , \32248_32547 , \32249_32548 , \32250_32549 , \32251_32550 , \32252_32551 , \32253_32552 , \32254_32553 , \32255_32554 , \32256_32555 , \32257_32556 , \32258_32557 , \32259_32558 , \32260_32559 , \32261_32560 , \32262_32561 , \32263_32562 , \32264_32563 , \32265_32564 , \32266_32565 , \32267_32566 , \32268_32567 , \32269_32568 , \32270_32569 , \32271_32570 , \32272_32571 , \32273_32572 , \32274_32573 , \32275_32574 , \32276_32575 , \32277_32576 , \32278_32577 , \32279_32578 , \32280_32579 , \32281_32580 , \32282_32581 , \32283_32582 , \32284_32583 , \32285_32584 , \32286_32585 , \32287_32586 , \32288_32587 , \32289_32588 , \32290_32589 , \32291_32590 , \32292_32591 , \32293_32592 );
and \U$23520 ( \32295_32594 , RIee2c6c8_4964, \9163_9462 );
and \U$23521 ( \32296_32595 , RIee2ac10_4945, \9165_9464 );
and \U$23522 ( \32297_32596 , RIee29590_4929, \9167_9466 );
and \U$23523 ( \32298_32597 , RIee28348_4916, \9169_9468 );
and \U$23524 ( \32299_32598 , RIdf2ad78_1864, \9171_9470 );
and \U$23525 ( \32300_32599 , RIdf28e88_1842, \9173_9472 );
and \U$23526 ( \32301_32600 , RIfea3608_8203, \9175_9474 );
and \U$23527 ( \32302_32601 , RIfea3770_8204, \9177_9476 );
and \U$23528 ( \32303_32602 , RIfcc0d10_7216, \9179_9478 );
and \U$23529 ( \32304_32603 , RIfc75c20_6362, \9181_9480 );
and \U$23530 ( \32305_32604 , RIfca50b0_6900, \9183_9482 );
and \U$23531 ( \32306_32605 , RIfc74e10_6352, \9185_9484 );
and \U$23532 ( \32307_32606 , RIfcc9410_7312, \9187_9486 );
and \U$23533 ( \32308_32607 , RIdf20620_1745, \9189_9488 );
and \U$23534 ( \32309_32608 , RIfc73628_6335, \9191_9490 );
and \U$23535 ( \32310_32609 , RIdf1a0e0_1673, \9193_9492 );
and \U$23536 ( \32311_32610 , RIdf17f20_1649, \9195_9494 );
and \U$23537 ( \32312_32611 , RIdf15220_1617, \9197_9496 );
and \U$23538 ( \32313_32612 , RIdf12520_1585, \9199_9498 );
and \U$23539 ( \32314_32613 , RIdf0f820_1553, \9201_9500 );
and \U$23540 ( \32315_32614 , RIdf0cb20_1521, \9203_9502 );
and \U$23541 ( \32316_32615 , RIdf09e20_1489, \9205_9504 );
and \U$23542 ( \32317_32616 , RIdf07120_1457, \9207_9506 );
and \U$23543 ( \32318_32617 , RIdf04420_1425, \9209_9508 );
and \U$23544 ( \32319_32618 , RIdefea20_1361, \9211_9510 );
and \U$23545 ( \32320_32619 , RIdefbd20_1329, \9213_9512 );
and \U$23546 ( \32321_32620 , RIdef9020_1297, \9215_9514 );
and \U$23547 ( \32322_32621 , RIdef6320_1265, \9217_9516 );
and \U$23548 ( \32323_32622 , RIdef3620_1233, \9219_9518 );
and \U$23549 ( \32324_32623 , RIdef0920_1201, \9221_9520 );
and \U$23550 ( \32325_32624 , RIdeedc20_1169, \9223_9522 );
and \U$23551 ( \32326_32625 , RIdeeaf20_1137, \9225_9524 );
and \U$23552 ( \32327_32626 , RIfcab8c0_6974, \9227_9526 );
and \U$23553 ( \32328_32627 , RIfc7c598_6437, \9229_9528 );
and \U$23554 ( \32329_32628 , RIfc5beb0_6068, \9231_9530 );
and \U$23555 ( \32330_32629 , RIfc58ee0_6034, \9233_9532 );
and \U$23556 ( \32331_32630 , RIdee5688_1074, \9235_9534 );
and \U$23557 ( \32332_32631 , RIdee3798_1052, \9237_9536 );
and \U$23558 ( \32333_32632 , RIdee15d8_1028, \9239_9538 );
and \U$23559 ( \32334_32633 , RIdedf580_1005, \9241_9540 );
and \U$23560 ( \32335_32634 , RIfcb3048_7059, \9243_9542 );
and \U$23561 ( \32336_32635 , RIfc72ae8_6327, \9245_9544 );
and \U$23562 ( \32337_32636 , RIfca3d00_6886, \9247_9546 );
and \U$23563 ( \32338_32637 , RIfcb6450_7096, \9249_9548 );
and \U$23564 ( \32339_32638 , RIdeda558_948, \9251_9550 );
and \U$23565 ( \32340_32639 , RIded7f60_921, \9253_9552 );
and \U$23566 ( \32341_32640 , RIfea3068_8199, \9255_9554 );
and \U$23567 ( \32342_32641 , RIded3a78_872, \9257_9556 );
and \U$23568 ( \32343_32642 , RIded1750_847, \9259_9558 );
and \U$23569 ( \32344_32643 , RIdecea50_815, \9261_9560 );
and \U$23570 ( \32345_32644 , RIdecbd50_783, \9263_9562 );
and \U$23571 ( \32346_32645 , RIdec9050_751, \9265_9564 );
and \U$23572 ( \32347_32646 , RIdeb5550_527, \9267_9566 );
and \U$23573 ( \32348_32647 , RIde98d38_335, \9269_9568 );
and \U$23574 ( \32349_32648 , RIe16f158_2641, \9271_9570 );
and \U$23575 ( \32350_32649 , RIe15af50_2412, \9273_9572 );
and \U$23576 ( \32351_32650 , RIe144750_2156, \9275_9574 );
and \U$23577 ( \32352_32651 , RIdf39148_2026, \9277_9576 );
and \U$23578 ( \32353_32652 , RIdf2d7a8_1894, \9279_9578 );
and \U$23579 ( \32354_32653 , RIdf1e028_1718, \9281_9580 );
and \U$23580 ( \32355_32654 , RIdf01720_1393, \9283_9582 );
and \U$23581 ( \32356_32655 , RIdee8220_1105, \9285_9584 );
and \U$23582 ( \32357_32656 , RIdedcf88_978, \9287_9586 );
and \U$23583 ( \32358_32657 , RIde7ec80_208, \9289_9588 );
or \U$23584 ( \32359_32658 , \32295_32594 , \32296_32595 , \32297_32596 , \32298_32597 , \32299_32598 , \32300_32599 , \32301_32600 , \32302_32601 , \32303_32602 , \32304_32603 , \32305_32604 , \32306_32605 , \32307_32606 , \32308_32607 , \32309_32608 , \32310_32609 , \32311_32610 , \32312_32611 , \32313_32612 , \32314_32613 , \32315_32614 , \32316_32615 , \32317_32616 , \32318_32617 , \32319_32618 , \32320_32619 , \32321_32620 , \32322_32621 , \32323_32622 , \32324_32623 , \32325_32624 , \32326_32625 , \32327_32626 , \32328_32627 , \32329_32628 , \32330_32629 , \32331_32630 , \32332_32631 , \32333_32632 , \32334_32633 , \32335_32634 , \32336_32635 , \32337_32636 , \32338_32637 , \32339_32638 , \32340_32639 , \32341_32640 , \32342_32641 , \32343_32642 , \32344_32643 , \32345_32644 , \32346_32645 , \32347_32646 , \32348_32647 , \32349_32648 , \32350_32649 , \32351_32650 , \32352_32651 , \32353_32652 , \32354_32653 , \32355_32654 , \32356_32655 , \32357_32656 , \32358_32657 );
or \U$23585 ( \32360_32659 , \32294_32593 , \32359_32658 );
_DC \g65d4/U$1 ( \32361 , \32360_32659 , \9298_9597 );
and \U$23586 ( \32362_32661 , RIe19e5e8_3179, \8760_9059 );
and \U$23587 ( \32363_32662 , RIe19b8e8_3147, \8762_9061 );
and \U$23588 ( \32364_32663 , RIfca84b8_6937, \8764_9063 );
and \U$23589 ( \32365_32664 , RIe198be8_3115, \8766_9065 );
and \U$23590 ( \32366_32665 , RIfc846f8_6529, \8768_9067 );
and \U$23591 ( \32367_32666 , RIe195ee8_3083, \8770_9069 );
and \U$23592 ( \32368_32667 , RIe1931e8_3051, \8772_9071 );
and \U$23593 ( \32369_32668 , RIe1904e8_3019, \8774_9073 );
and \U$23594 ( \32370_32669 , RIe18aae8_2955, \8776_9075 );
and \U$23595 ( \32371_32670 , RIe187de8_2923, \8778_9077 );
and \U$23596 ( \32372_32671 , RIfce2be0_7602, \8780_9079 );
and \U$23597 ( \32373_32672 , RIe1850e8_2891, \8782_9081 );
and \U$23598 ( \32374_32673 , RIfc8e310_6640, \8784_9083 );
and \U$23599 ( \32375_32674 , RIe1823e8_2859, \8786_9085 );
and \U$23600 ( \32376_32675 , RIe17f6e8_2827, \8788_9087 );
and \U$23601 ( \32377_32676 , RIe17c9e8_2795, \8790_9089 );
and \U$23602 ( \32378_32677 , RIfcd1570_7404, \8792_9091 );
and \U$23603 ( \32379_32678 , RIfccc278_7345, \8794_9093 );
and \U$23604 ( \32380_32679 , RIf1404c8_5191, \8796_9095 );
and \U$23605 ( \32381_32680 , RIfea2d98_8197, \8798_9097 );
and \U$23606 ( \32382_32681 , RIfcc1b20_7226, \8800_9099 );
and \U$23607 ( \32383_32682 , RIfc60398_6117, \8802_9101 );
and \U$23608 ( \32384_32683 , RIee3e5a8_5168, \8804_9103 );
and \U$23609 ( \32385_32684 , RIee3da68_5160, \8806_9105 );
and \U$23610 ( \32386_32685 , RIfc642e0_6162, \8808_9107 );
and \U$23611 ( \32387_32686 , RIfca7f18_6933, \8810_9109 );
and \U$23612 ( \32388_32687 , RIee3a228_5120, \8812_9111 );
and \U$23613 ( \32389_32688 , RIfec6180_8374, \8814_9113 );
and \U$23614 ( \32390_32689 , RIfca9598_6949, \8816_9115 );
and \U$23615 ( \32391_32690 , RIfc5c720_6074, \8818_9117 );
and \U$23616 ( \32392_32691 , RIfc6bea0_6250, \8820_9119 );
and \U$23617 ( \32393_32692 , RIfccaec8_7331, \8822_9121 );
and \U$23618 ( \32394_32693 , RIfc44cd8_5805, \8824_9123 );
and \U$23619 ( \32395_32694 , RIe224940_4706, \8826_9125 );
and \U$23620 ( \32396_32695 , RIfcb6180_7094, \8828_9127 );
and \U$23621 ( \32397_32696 , RIe221c40_4674, \8830_9129 );
and \U$23622 ( \32398_32697 , RIfc55ad8_5997, \8832_9131 );
and \U$23623 ( \32399_32698 , RIe21ef40_4642, \8834_9133 );
and \U$23624 ( \32400_32699 , RIe219540_4578, \8836_9135 );
and \U$23625 ( \32401_32700 , RIe216840_4546, \8838_9137 );
and \U$23626 ( \32402_32701 , RIfc4dc48_5907, \8840_9139 );
and \U$23627 ( \32403_32702 , RIe213b40_4514, \8842_9141 );
and \U$23628 ( \32404_32703 , RIfcdcf10_7536, \8844_9143 );
and \U$23629 ( \32405_32704 , RIe210e40_4482, \8846_9145 );
and \U$23630 ( \32406_32705 , RIfcab1b8_6969, \8848_9147 );
and \U$23631 ( \32407_32706 , RIe20e140_4450, \8850_9149 );
and \U$23632 ( \32408_32707 , RIe20b440_4418, \8852_9151 );
and \U$23633 ( \32409_32708 , RIe208740_4386, \8854_9153 );
and \U$23634 ( \32410_32709 , RIfce3720_7610, \8856_9155 );
and \U$23635 ( \32411_32710 , RIfc64178_6161, \8858_9157 );
and \U$23636 ( \32412_32711 , RIe203178_4325, \8860_9159 );
and \U$23637 ( \32413_32712 , RIe201558_4305, \8862_9161 );
and \U$23638 ( \32414_32713 , RIfcd2ec0_7422, \8864_9163 );
and \U$23639 ( \32415_32714 , RIf164828_5603, \8866_9165 );
and \U$23640 ( \32416_32715 , RIfc7f838_6473, \8868_9167 );
and \U$23641 ( \32417_32716 , RIf162398_5577, \8870_9169 );
and \U$23642 ( \32418_32717 , RIfcc9c80_7318, \8872_9171 );
and \U$23643 ( \32419_32718 , RIfca8bc0_6942, \8874_9173 );
and \U$23644 ( \32420_32719 , RIfea2ac8_8195, \8876_9175 );
and \U$23645 ( \32421_32720 , RIfea2c30_8196, \8878_9177 );
and \U$23646 ( \32422_32721 , RIfc59318_6037, \8880_9179 );
and \U$23647 ( \32423_32722 , RIfc4f160_5922, \8882_9181 );
and \U$23648 ( \32424_32723 , RIf15ac10_5492, \8884_9183 );
and \U$23649 ( \32425_32724 , RIfcebf88_7707, \8886_9185 );
or \U$23650 ( \32426_32725 , \32362_32661 , \32363_32662 , \32364_32663 , \32365_32664 , \32366_32665 , \32367_32666 , \32368_32667 , \32369_32668 , \32370_32669 , \32371_32670 , \32372_32671 , \32373_32672 , \32374_32673 , \32375_32674 , \32376_32675 , \32377_32676 , \32378_32677 , \32379_32678 , \32380_32679 , \32381_32680 , \32382_32681 , \32383_32682 , \32384_32683 , \32385_32684 , \32386_32685 , \32387_32686 , \32388_32687 , \32389_32688 , \32390_32689 , \32391_32690 , \32392_32691 , \32393_32692 , \32394_32693 , \32395_32694 , \32396_32695 , \32397_32696 , \32398_32697 , \32399_32698 , \32400_32699 , \32401_32700 , \32402_32701 , \32403_32702 , \32404_32703 , \32405_32704 , \32406_32705 , \32407_32706 , \32408_32707 , \32409_32708 , \32410_32709 , \32411_32710 , \32412_32711 , \32413_32712 , \32414_32713 , \32415_32714 , \32416_32715 , \32417_32716 , \32418_32717 , \32419_32718 , \32420_32719 , \32421_32720 , \32422_32721 , \32423_32722 , \32424_32723 , \32425_32724 );
and \U$23651 ( \32427_32726 , RIfcbb040_7150, \8889_9188 );
and \U$23652 ( \32428_32727 , RIfca1870_6860, \8891_9190 );
and \U$23653 ( \32429_32728 , RIfc93d10_6704, \8893_9192 );
and \U$23654 ( \32430_32729 , RIe1faeb0_4232, \8895_9194 );
and \U$23655 ( \32431_32730 , RIf1565c0_5442, \8897_9196 );
and \U$23656 ( \32432_32731 , RIf155a80_5434, \8899_9198 );
and \U$23657 ( \32433_32732 , RIfc45c50_5816, \8901_9200 );
and \U$23658 ( \32434_32733 , RIe1f6428_4179, \8903_9202 );
and \U$23659 ( \32435_32734 , RIfccdbc8_7363, \8905_9204 );
and \U$23660 ( \32436_32735 , RIfcccae8_7351, \8907_9206 );
and \U$23661 ( \32437_32736 , RIfca6cd0_6920, \8909_9208 );
and \U$23662 ( \32438_32737 , RIfec6018_8373, \8911_9210 );
and \U$23663 ( \32439_32738 , RIfc64010_6160, \8913_9212 );
and \U$23664 ( \32440_32739 , RIfc434f0_5788, \8915_9214 );
and \U$23665 ( \32441_32740 , RIfc4c028_5887, \8917_9216 );
and \U$23666 ( \32442_32741 , RIe1eee08_4095, \8919_9218 );
and \U$23667 ( \32443_32742 , RIe1ec6a8_4067, \8921_9220 );
and \U$23668 ( \32444_32743 , RIe1e99a8_4035, \8923_9222 );
and \U$23669 ( \32445_32744 , RIe1e6ca8_4003, \8925_9224 );
and \U$23670 ( \32446_32745 , RIe1e3fa8_3971, \8927_9226 );
and \U$23671 ( \32447_32746 , RIe1e12a8_3939, \8929_9228 );
and \U$23672 ( \32448_32747 , RIe1de5a8_3907, \8931_9230 );
and \U$23673 ( \32449_32748 , RIe1db8a8_3875, \8933_9232 );
and \U$23674 ( \32450_32749 , RIe1d8ba8_3843, \8935_9234 );
and \U$23675 ( \32451_32750 , RIe1d31a8_3779, \8937_9236 );
and \U$23676 ( \32452_32751 , RIe1d04a8_3747, \8939_9238 );
and \U$23677 ( \32453_32752 , RIe1cd7a8_3715, \8941_9240 );
and \U$23678 ( \32454_32753 , RIe1caaa8_3683, \8943_9242 );
and \U$23679 ( \32455_32754 , RIe1c7da8_3651, \8945_9244 );
and \U$23680 ( \32456_32755 , RIe1c50a8_3619, \8947_9246 );
and \U$23681 ( \32457_32756 , RIe1c23a8_3587, \8949_9248 );
and \U$23682 ( \32458_32757 , RIe1bf6a8_3555, \8951_9250 );
and \U$23683 ( \32459_32758 , RIfc63908_6155, \8953_9252 );
and \U$23684 ( \32460_32759 , RIfc6bd38_6249, \8955_9254 );
and \U$23685 ( \32461_32760 , RIe1ba0e0_3494, \8957_9256 );
and \U$23686 ( \32462_32761 , RIe1b7f20_3470, \8959_9258 );
and \U$23687 ( \32463_32762 , RIfc66fe0_6194, \8961_9260 );
and \U$23688 ( \32464_32763 , RIfc92ac8_6691, \8963_9262 );
and \U$23689 ( \32465_32764 , RIe1b5d60_3446, \8965_9264 );
and \U$23690 ( \32466_32765 , RIfea2f00_8198, \8967_9266 );
and \U$23691 ( \32467_32766 , RIfc9bfd8_6797, \8969_9268 );
and \U$23692 ( \32468_32767 , RIfc50d80_5942, \8971_9270 );
and \U$23693 ( \32469_32768 , RIe1b31c8_3415, \8973_9272 );
and \U$23694 ( \32470_32769 , RIe1b1878_3397, \8975_9274 );
and \U$23695 ( \32471_32770 , RIfc4df18_5909, \8977_9276 );
and \U$23696 ( \32472_32771 , RIfc9d658_6813, \8979_9278 );
and \U$23697 ( \32473_32772 , RIe1ad0c0_3346, \8981_9280 );
and \U$23698 ( \32474_32773 , RIe1ab8d8_3329, \8983_9282 );
and \U$23699 ( \32475_32774 , RIe1a99e8_3307, \8985_9284 );
and \U$23700 ( \32476_32775 , RIe1a6ce8_3275, \8987_9286 );
and \U$23701 ( \32477_32776 , RIe1a3fe8_3243, \8989_9288 );
and \U$23702 ( \32478_32777 , RIe1a12e8_3211, \8991_9290 );
and \U$23703 ( \32479_32778 , RIe18d7e8_2987, \8993_9292 );
and \U$23704 ( \32480_32779 , RIe179ce8_2763, \8995_9294 );
and \U$23705 ( \32481_32780 , RIe227640_4738, \8997_9296 );
and \U$23706 ( \32482_32781 , RIe21c240_4610, \8999_9298 );
and \U$23707 ( \32483_32782 , RIe205a40_4354, \9001_9300 );
and \U$23708 ( \32484_32783 , RIe1ffaa0_4286, \9003_9302 );
and \U$23709 ( \32485_32784 , RIe1f8e58_4209, \9005_9304 );
and \U$23710 ( \32486_32785 , RIe1f19a0_4126, \9007_9306 );
and \U$23711 ( \32487_32786 , RIe1d5ea8_3811, \9009_9308 );
and \U$23712 ( \32488_32787 , RIe1bc9a8_3523, \9011_9310 );
and \U$23713 ( \32489_32788 , RIe1af820_3374, \9013_9312 );
and \U$23714 ( \32490_32789 , RIe171e58_2673, \9015_9314 );
or \U$23715 ( \32491_32790 , \32427_32726 , \32428_32727 , \32429_32728 , \32430_32729 , \32431_32730 , \32432_32731 , \32433_32732 , \32434_32733 , \32435_32734 , \32436_32735 , \32437_32736 , \32438_32737 , \32439_32738 , \32440_32739 , \32441_32740 , \32442_32741 , \32443_32742 , \32444_32743 , \32445_32744 , \32446_32745 , \32447_32746 , \32448_32747 , \32449_32748 , \32450_32749 , \32451_32750 , \32452_32751 , \32453_32752 , \32454_32753 , \32455_32754 , \32456_32755 , \32457_32756 , \32458_32757 , \32459_32758 , \32460_32759 , \32461_32760 , \32462_32761 , \32463_32762 , \32464_32763 , \32465_32764 , \32466_32765 , \32467_32766 , \32468_32767 , \32469_32768 , \32470_32769 , \32471_32770 , \32472_32771 , \32473_32772 , \32474_32773 , \32475_32774 , \32476_32775 , \32477_32776 , \32478_32777 , \32479_32778 , \32480_32779 , \32481_32780 , \32482_32781 , \32483_32782 , \32484_32783 , \32485_32784 , \32486_32785 , \32487_32786 , \32488_32787 , \32489_32788 , \32490_32789 );
or \U$23716 ( \32492_32791 , \32426_32725 , \32491_32790 );
_DC \g65d5/U$1 ( \32493 , \32492_32791 , \9024_9323 );
and g65d6_GF_PartitionCandidate( \32494_32793_nG65d6 , \32361 , \32493 );
buf \U$23717 ( \32495_32794 , \32494_32793_nG65d6 );
and \U$23718 ( \32496_32795 , \32495_32794 , \10389_10691 );
nor \U$23719 ( \32497_32796 , \32229_32528 , \32496_32795 );
xnor \U$23720 ( \32498_32797 , \32497_32796 , \10678_10980 );
not \U$23721 ( \32499_32798 , \31766_32068 );
_DC \g64f1/U$1 ( \32500 , \32360_32659 , \9298_9597 );
_DC \g6575/U$1 ( \32501 , \32492_32791 , \9024_9323 );
xor g6576_GF_PartitionCandidate( \32502_32801_nG6576 , \32500 , \32501 );
buf \U$23722 ( \32503_32802 , \32502_32801_nG6576 );
and \U$23723 ( \32504_32803 , \31764_32066 , \30508_30810 );
not \U$23724 ( \32505_32804 , \32504_32803 );
and \U$23725 ( \32506_32805 , \32503_32802 , \32505_32804 );
and \U$23726 ( \32507_32806 , \32499_32798 , \32506_32805 );
xor \U$23727 ( \32508_32807 , \32498_32797 , \32507_32806 );
and \U$23728 ( \32509_32808 , \31755_32057 , \31759_32061 );
and \U$23729 ( \32510_32809 , \31759_32061 , \31766_32068 );
and \U$23730 ( \32511_32810 , \31755_32057 , \31766_32068 );
or \U$23731 ( \32512_32811 , \32509_32808 , \32510_32809 , \32511_32810 );
xor \U$23732 ( \32513_32812 , \32508_32807 , \32512_32811 );
and \U$23733 ( \32514_32813 , \31853_32155 , \31857_32159 );
and \U$23734 ( \32515_32814 , \31857_32159 , \31862_32164 );
and \U$23735 ( \32516_32815 , \31853_32155 , \31862_32164 );
or \U$23736 ( \32517_32816 , \32514_32813 , \32515_32814 , \32516_32815 );
xor \U$23737 ( \32518_32817 , \32513_32812 , \32517_32816 );
xor \U$23738 ( \32519_32818 , \32228_32527 , \32518_32817 );
xor \U$23739 ( \32520_32819 , \32209_32508 , \32519_32818 );
and \U$23740 ( \32521_32820 , \31485_31787 , \31767_32069 );
and \U$23741 ( \32522_32821 , \31767_32069 , \31782_32084 );
and \U$23742 ( \32523_32822 , \31485_31787 , \31782_32084 );
or \U$23743 ( \32524_32823 , \32521_32820 , \32522_32821 , \32523_32822 );
and \U$23744 ( \32525_32824 , \31834_32136 , \31848_32150 );
and \U$23745 ( \32526_32825 , \31848_32150 , \31863_32165 );
and \U$23746 ( \32527_32826 , \31834_32136 , \31863_32165 );
or \U$23747 ( \32528_32827 , \32525_32824 , \32526_32825 , \32527_32826 );
xor \U$23748 ( \32529_32828 , \32524_32823 , \32528_32827 );
and \U$23749 ( \32530_32829 , \21788_22090 , \17791_18090 );
and \U$23750 ( \32531_32830 , \22257_22556 , \17353_17655 );
nor \U$23751 ( \32532_32831 , \32530_32829 , \32531_32830 );
xnor \U$23752 ( \32533_32832 , \32532_32831 , \17747_18046 );
and \U$23753 ( \32534_32833 , \12146_12448 , \28768_29070 );
and \U$23754 ( \32535_32834 , \12470_12769 , \28224_28526 );
nor \U$23755 ( \32536_32835 , \32534_32833 , \32535_32834 );
xnor \U$23756 ( \32537_32836 , \32536_32835 , \28774_29076 );
xor \U$23757 ( \32538_32837 , \32533_32832 , \32537_32836 );
and \U$23758 ( \32539_32838 , \10968_11270 , \30521_30823 );
and \U$23759 ( \32540_32839 , \11287_11586 , \29944_30246 );
nor \U$23760 ( \32541_32840 , \32539_32838 , \32540_32839 );
xnor \U$23761 ( \32542_32841 , \32541_32840 , \30511_30813 );
xor \U$23762 ( \32543_32842 , \32538_32837 , \32542_32841 );
and \U$23763 ( \32544_32843 , \29966_30268 , \11275_11574 );
and \U$23764 ( \32545_32844 , \30500_30802 , \10976_11278 );
nor \U$23765 ( \32546_32845 , \32544_32843 , \32545_32844 );
xnor \U$23766 ( \32547_32846 , \32546_32845 , \11281_11580 );
and \U$23767 ( \32548_32847 , \26527_26829 , \13755_14054 );
and \U$23768 ( \32549_32848 , \27011_27313 , \13390_13692 );
nor \U$23769 ( \32550_32849 , \32548_32847 , \32549_32848 );
xnor \U$23770 ( \32551_32850 , \32550_32849 , \13736_14035 );
xor \U$23771 ( \32552_32851 , \32547_32846 , \32551_32850 );
xor \U$23772 ( \32553_32852 , \32503_32802 , \31764_32066 );
not \U$23773 ( \32554_32853 , \31765_32067 );
and \U$23774 ( \32555_32854 , \32553_32852 , \32554_32853 );
and \U$23775 ( \32556_32855 , \10385_10687 , \32555_32854 );
and \U$23776 ( \32557_32856 , \10686_10988 , \31765_32067 );
nor \U$23777 ( \32558_32857 , \32556_32855 , \32557_32856 );
xnor \U$23778 ( \32559_32858 , \32558_32857 , \32506_32805 );
xor \U$23779 ( \32560_32859 , \32552_32851 , \32559_32858 );
xor \U$23780 ( \32561_32860 , \32543_32842 , \32560_32859 );
and \U$23781 ( \32562_32861 , \24970_25272 , \15037_15336 );
and \U$23782 ( \32563_32862 , \25516_25815 , \14661_14963 );
nor \U$23783 ( \32564_32863 , \32562_32861 , \32563_32862 );
xnor \U$23784 ( \32565_32864 , \32564_32863 , \15043_15342 );
and \U$23785 ( \32566_32865 , \20242_20544 , \19235_19534 );
and \U$23786 ( \32567_32866 , \20734_21033 , \18743_19045 );
nor \U$23787 ( \32568_32867 , \32566_32865 , \32567_32866 );
xnor \U$23788 ( \32569_32868 , \32568_32867 , \19241_19540 );
xor \U$23789 ( \32570_32869 , \32565_32864 , \32569_32868 );
and \U$23790 ( \32571_32870 , \18730_19032 , \20706_21005 );
and \U$23791 ( \32572_32871 , \19259_19558 , \20255_20557 );
nor \U$23792 ( \32573_32872 , \32571_32870 , \32572_32871 );
xnor \U$23793 ( \32574_32873 , \32573_32872 , \20712_21011 );
xor \U$23794 ( \32575_32874 , \32570_32869 , \32574_32873 );
xor \U$23795 ( \32576_32875 , \32561_32860 , \32575_32874 );
xor \U$23796 ( \32577_32876 , \32529_32828 , \32576_32875 );
xor \U$23797 ( \32578_32877 , \32520_32819 , \32577_32876 );
xor \U$23798 ( \32579_32878 , \32205_32504 , \32578_32877 );
and \U$23799 ( \32580_32879 , \31462_31764 , \31784_32086 );
and \U$23800 ( \32581_32880 , \31784_32086 , \31866_32168 );
and \U$23801 ( \32582_32881 , \31462_31764 , \31866_32168 );
or \U$23802 ( \32583_32882 , \32580_32879 , \32581_32880 , \32582_32881 );
xor \U$23803 ( \32584_32883 , \32579_32878 , \32583_32882 );
and \U$23804 ( \32585_32884 , \31867_32169 , \31871_32173 );
and \U$23805 ( \32586_32885 , \31872_32174 , \31875_32177 );
or \U$23806 ( \32587_32886 , \32585_32884 , \32586_32885 );
xor \U$23807 ( \32588_32887 , \32584_32883 , \32587_32886 );
buf g9bb1_GF_PartitionCandidate( \32589_32888_nG9bb1 , \32588_32887 );
and \U$23808 ( \32590_32889 , \10402_10704 , \32589_32888_nG9bb1 );
or \U$23809 ( \32591_32890 , \32156_32455 , \32590_32889 );
xor \U$23810 ( \32592_32891 , \10399_10703 , \32591_32890 );
buf \U$23811 ( \32593_32892 , \32592_32891 );
buf \U$23813 ( \32594_32893 , \32593_32892 );
xor \U$23814 ( \32595_32894 , \32155_32454 , \32594_32893 );
buf \U$23815 ( \32596_32895 , \32595_32894 );
xor \U$23816 ( \32597_32896 , \32143_32442 , \32596_32895 );
and \U$23817 ( \32598_32897 , \31410_31712 , \31456_31758 );
and \U$23818 ( \32599_32898 , \31410_31712 , \31882_32184 );
and \U$23819 ( \32600_32899 , \31456_31758 , \31882_32184 );
or \U$23820 ( \32601_32900 , \32598_32897 , \32599_32898 , \32600_32899 );
buf \U$23821 ( \32602_32901 , \32601_32900 );
xor \U$23822 ( \32603_32902 , \32597_32896 , \32602_32901 );
buf \U$23823 ( \32604_32903 , \32603_32902 );
xor \U$23824 ( \32605_32904 , \32085_32384 , \32604_32903 );
xor \U$23825 ( \32606_32905 , \31965_32267 , \32605_32904 );
and \U$23826 ( \32607_32906 , \31351_31653 , \31886_32188 );
and \U$23827 ( \32608_32907 , \31351_31653 , \31956_32258 );
and \U$23828 ( \32609_32908 , \31886_32188 , \31956_32258 );
or \U$23829 ( \32610_32909 , \32607_32906 , \32608_32907 , \32609_32908 );
and \U$23830 ( \32611_32910 , \32606_32905 , \32610_32909 );
and \U$23831 ( \32612_32911 , \31960_32262 , \31964_32266 );
and \U$23832 ( \32613_32912 , \31960_32262 , \32605_32904 );
and \U$23833 ( \32614_32913 , \31964_32266 , \32605_32904 );
or \U$23834 ( \32615_32914 , \32612_32911 , \32613_32912 , \32614_32913 );
xor \U$23835 ( \32616_32915 , \32611_32910 , \32615_32914 );
xor \U$23840 ( \32617_32916 , 1'b0 , \31328_31627_nG43fa );
and \U$23845 ( \32618_32918 , \32617_32916 , \10392_10694_nG9c0e );
or \U$23846 ( \32619_32919 , 1'b0 , \32618_32918 );
xor \U$23847 ( \32620_32920 , 1'b0 , \32619_32919 );
xor \U$23848 ( \32621_32921 , 1'b0 , \32620_32920 );
buf \U$23849 ( \32622_32922 , \32621_32921 );
buf \U$23850 ( \32623_32923 , \32622_32922 );
xor \U$23851 ( \32624_32924 , \32616_32915 , \32623_32923 );
and \U$23852 ( \32625_32925 , \32079_32378 , \32084_32383 );
and \U$23853 ( \32626_32926 , \32079_32378 , \32604_32903 );
and \U$23854 ( \32627_32927 , \32084_32383 , \32604_32903 );
or \U$23855 ( \32628_32928 , \32625_32925 , \32626_32926 , \32627_32927 );
and \U$23856 ( \32629_32929 , \32624_32924 , \32628_32928 );
and \U$23857 ( \32630_32930 , \32043_32342 , \32063_32362 );
and \U$23858 ( \32631_32931 , \32043_32342 , \32069_32368 );
and \U$23859 ( \32632_32932 , \32063_32362 , \32069_32368 );
or \U$23860 ( \32633_32933 , \32630_32930 , \32631_32931 , \32632_32932 );
buf \U$23861 ( \32634_32934 , \32633_32933 );
and \U$23862 ( \32635_32935 , \32090_32389 , \32107_32406 );
and \U$23863 ( \32636_32936 , \32090_32389 , \32114_32413 );
and \U$23864 ( \32637_32937 , \32107_32406 , \32114_32413 );
or \U$23865 ( \32638_32938 , \32635_32935 , \32636_32936 , \32637_32937 );
buf \U$23866 ( \32639_32939 , \32638_32938 );
and \U$23867 ( \32640_32940 , \31978_32280 , \31984_32286 );
buf \U$23868 ( \32641_32941 , \32640_32940 );
and \U$23869 ( \32642_32942 , \28946_28118 , \12502_12801_nG9bff );
and \U$23870 ( \32643_32943 , \27816_28115 , \13403_13705_nG9bfc );
or \U$23871 ( \32644_32944 , \32642_32942 , \32643_32943 );
xor \U$23872 ( \32645_32945 , \27815_28114 , \32644_32944 );
buf \U$23873 ( \32646_32946 , \32645_32945 );
buf \U$23875 ( \32647_32947 , \32646_32946 );
xor \U$23876 ( \32648_32948 , \32641_32941 , \32647_32947 );
and \U$23877 ( \32649_32949 , \27141_26431 , \13771_14070_nG9bf9 );
and \U$23878 ( \32650_32950 , \26129_26428 , \14682_14984_nG9bf6 );
or \U$23879 ( \32651_32951 , \32649_32949 , \32650_32950 );
xor \U$23880 ( \32652_32952 , \26128_26427 , \32651_32951 );
buf \U$23881 ( \32653_32953 , \32652_32952 );
buf \U$23883 ( \32654_32954 , \32653_32953 );
xor \U$23884 ( \32655_32955 , \32648_32948 , \32654_32954 );
buf \U$23885 ( \32656_32956 , \32655_32955 );
and \U$23886 ( \32657_32957 , \23495_23201 , \16378_16680_nG9bed );
and \U$23887 ( \32658_32958 , \22899_23198 , \17363_17665_nG9bea );
or \U$23888 ( \32659_32959 , \32657_32957 , \32658_32958 );
xor \U$23889 ( \32660_32960 , \22898_23197 , \32659_32959 );
buf \U$23890 ( \32661_32961 , \32660_32960 );
buf \U$23892 ( \32662_32962 , \32661_32961 );
xor \U$23893 ( \32663_32963 , \32656_32956 , \32662_32962 );
and \U$23894 ( \32664_32964 , \21908_21658 , \17808_18107_nG9be7 );
and \U$23895 ( \32665_32965 , \21356_21655 , \18789_19091_nG9be4 );
or \U$23896 ( \32666_32966 , \32664_32964 , \32665_32965 );
xor \U$23897 ( \32667_32967 , \21355_21654 , \32666_32966 );
buf \U$23898 ( \32668_32968 , \32667_32967 );
buf \U$23900 ( \32669_32969 , \32668_32968 );
xor \U$23901 ( \32670_32970 , \32663_32963 , \32669_32969 );
buf \U$23902 ( \32671_32971 , \32670_32970 );
xor \U$23903 ( \32672_32972 , \32639_32939 , \32671_32971 );
and \U$23904 ( \32673_32973 , \16405_15940 , \23927_24226_nG9bcf );
and \U$23905 ( \32674_32974 , \15638_15937 , \24996_25298_nG9bcc );
or \U$23906 ( \32675_32975 , \32673_32973 , \32674_32974 );
xor \U$23907 ( \32676_32976 , \15637_15936 , \32675_32975 );
buf \U$23908 ( \32677_32977 , \32676_32976 );
buf \U$23910 ( \32678_32978 , \32677_32977 );
xor \U$23911 ( \32679_32979 , \32672_32972 , \32678_32978 );
buf \U$23912 ( \32680_32980 , \32679_32979 );
and \U$23913 ( \32681_32981 , \31975_32277 , \32004_32303 );
and \U$23914 ( \32682_32982 , \31975_32277 , \32011_32310 );
and \U$23915 ( \32683_32983 , \32004_32303 , \32011_32310 );
or \U$23916 ( \32684_32984 , \32681_32981 , \32682_32982 , \32683_32983 );
buf \U$23917 ( \32685_32985 , \32684_32984 );
and \U$23918 ( \32686_32986 , \31986_32288 , \31995_32294 );
and \U$23919 ( \32687_32987 , \31986_32288 , \32002_32301 );
and \U$23920 ( \32688_32988 , \31995_32294 , \32002_32301 );
or \U$23921 ( \32689_32989 , \32686_32986 , \32687_32987 , \32688_32988 );
buf \U$23922 ( \32690_32990 , \32689_32989 );
and \U$23923 ( \32691_32991 , \31989_31636 , \10693_10995_nG9c0b );
and \U$23924 ( \32692_32992 , \31334_31633 , \10981_11283_nG9c08 );
or \U$23925 ( \32693_32993 , \32691_32991 , \32692_32992 );
xor \U$23926 ( \32694_32994 , \31333_31632 , \32693_32993 );
buf \U$23927 ( \32695_32995 , \32694_32994 );
buf \U$23929 ( \32696_32996 , \32695_32995 );
and \U$23930 ( \32697_32997 , \30670_29853 , \11299_11598_nG9c05 );
and \U$23931 ( \32698_32998 , \29551_29850 , \12168_12470_nG9c02 );
or \U$23932 ( \32699_32999 , \32697_32997 , \32698_32998 );
xor \U$23933 ( \32700_33000 , \29550_29849 , \32699_32999 );
buf \U$23934 ( \32701_33001 , \32700_33000 );
buf \U$23936 ( \32702_33002 , \32701_33001 );
xor \U$23937 ( \32703_33003 , \32696_32996 , \32702_33002 );
buf \U$23938 ( \32704_33004 , \32703_33003 );
xor \U$23939 ( \32705_33005 , \32690_32990 , \32704_33004 );
and \U$23940 ( \32706_33006 , \25044_24792 , \15074_15373_nG9bf3 );
and \U$23941 ( \32707_33007 , \24490_24789 , \16013_16315_nG9bf0 );
or \U$23942 ( \32708_33008 , \32706_33006 , \32707_33007 );
xor \U$23943 ( \32709_33009 , \24489_24788 , \32708_33008 );
buf \U$23944 ( \32710_33010 , \32709_33009 );
buf \U$23946 ( \32711_33011 , \32710_33010 );
xor \U$23947 ( \32712_33012 , \32705_33005 , \32711_33011 );
buf \U$23948 ( \32713_33013 , \32712_33012 );
xor \U$23949 ( \32714_33014 , \32685_32985 , \32713_33013 );
and \U$23950 ( \32715_33015 , \17437_17297 , \22330_22629_nG9bd5 );
and \U$23951 ( \32716_33016 , \16995_17294 , \23394_23696_nG9bd2 );
or \U$23952 ( \32717_33017 , \32715_33015 , \32716_33016 );
xor \U$23953 ( \32718_33018 , \16994_17293 , \32717_33017 );
buf \U$23954 ( \32719_33019 , \32718_33018 );
buf \U$23956 ( \32720_33020 , \32719_33019 );
xor \U$23957 ( \32721_33021 , \32714_33014 , \32720_33020 );
buf \U$23958 ( \32722_33022 , \32721_33021 );
xor \U$23959 ( \32723_33023 , \32680_32980 , \32722_33022 );
and \U$23960 ( \32724_33024 , \10411_10707 , \32589_32888_nG9bb1 );
and \U$23961 ( \32725_33025 , \32160_32459 , \32204_32503 );
and \U$23962 ( \32726_33026 , \32204_32503 , \32578_32877 );
and \U$23963 ( \32727_33027 , \32160_32459 , \32578_32877 );
or \U$23964 ( \32728_33028 , \32725_33025 , \32726_33026 , \32727_33027 );
and \U$23965 ( \32729_33029 , \32164_32463 , \32168_32467 );
and \U$23966 ( \32730_33030 , \32168_32467 , \32203_32502 );
and \U$23967 ( \32731_33031 , \32164_32463 , \32203_32502 );
or \U$23968 ( \32732_33032 , \32729_33029 , \32730_33030 , \32731_33031 );
and \U$23969 ( \32733_33033 , \32209_32508 , \32519_32818 );
and \U$23970 ( \32734_33034 , \32519_32818 , \32577_32876 );
and \U$23971 ( \32735_33035 , \32209_32508 , \32577_32876 );
or \U$23972 ( \32736_33036 , \32733_33033 , \32734_33034 , \32735_33035 );
xor \U$23973 ( \32737_33037 , \32732_33032 , \32736_33036 );
and \U$23974 ( \32738_33038 , \32508_32807 , \32512_32811 );
and \U$23975 ( \32739_33039 , \32512_32811 , \32517_32816 );
and \U$23976 ( \32740_33040 , \32508_32807 , \32517_32816 );
or \U$23977 ( \32741_33041 , \32738_33038 , \32739_33039 , \32740_33040 );
and \U$23978 ( \32742_33042 , \32543_32842 , \32560_32859 );
and \U$23979 ( \32743_33043 , \32560_32859 , \32575_32874 );
and \U$23980 ( \32744_33044 , \32543_32842 , \32575_32874 );
or \U$23981 ( \32745_33045 , \32742_33042 , \32743_33043 , \32744_33044 );
xor \U$23982 ( \32746_33046 , \32741_33041 , \32745_33045 );
and \U$23983 ( \32747_33047 , \32533_32832 , \32537_32836 );
and \U$23984 ( \32748_33048 , \32537_32836 , \32542_32841 );
and \U$23985 ( \32749_33049 , \32533_32832 , \32542_32841 );
or \U$23986 ( \32750_33050 , \32747_33047 , \32748_33048 , \32749_33049 );
and \U$23987 ( \32751_33051 , \32177_32476 , \32181_32480 );
and \U$23988 ( \32752_33052 , \32181_32480 , \32186_32485 );
and \U$23989 ( \32753_33053 , \32177_32476 , \32186_32485 );
or \U$23990 ( \32754_33054 , \32751_33051 , \32752_33052 , \32753_33053 );
xor \U$23991 ( \32755_33055 , \32750_33050 , \32754_33054 );
and \U$23992 ( \32756_33056 , \32495_32794 , \10681_10983 );
not \U$23993 ( \32757_33057 , \32756_33056 );
xnor \U$23994 ( \32758_33058 , \32757_33057 , \10678_10980 );
and \U$23995 ( \32759_33059 , \30500_30802 , \11275_11574 );
and \U$23996 ( \32760_33060 , \31752_32054 , \10976_11278 );
nor \U$23997 ( \32761_33061 , \32759_33059 , \32760_33060 );
xnor \U$23998 ( \32762_33062 , \32761_33061 , \11281_11580 );
xor \U$23999 ( \32763_33063 , \32758_33058 , \32762_33062 );
and \U$24000 ( \32764_33064 , \10385_10687 , \32503_32802 );
xor \U$24001 ( \32765_33065 , \32763_33063 , \32764_33064 );
xor \U$24002 ( \32766_33066 , \32755_33055 , \32765_33065 );
xor \U$24003 ( \32767_33067 , \32746_33046 , \32766_33066 );
and \U$24004 ( \32768_33068 , \32173_32472 , \32187_32486 );
and \U$24005 ( \32769_33069 , \32187_32486 , \32202_32501 );
and \U$24006 ( \32770_33070 , \32173_32472 , \32202_32501 );
or \U$24007 ( \32771_33071 , \32768_33068 , \32769_33069 , \32770_33070 );
and \U$24008 ( \32772_33072 , \32547_32846 , \32551_32850 );
and \U$24009 ( \32773_33073 , \32551_32850 , \32559_32858 );
and \U$24010 ( \32774_33074 , \32547_32846 , \32559_32858 );
or \U$24011 ( \32775_33075 , \32772_33072 , \32773_33073 , \32774_33074 );
and \U$24012 ( \32776_33076 , \32565_32864 , \32569_32868 );
and \U$24013 ( \32777_33077 , \32569_32868 , \32574_32873 );
and \U$24014 ( \32778_33078 , \32565_32864 , \32574_32873 );
or \U$24015 ( \32779_33079 , \32776_33076 , \32777_33077 , \32778_33078 );
xor \U$24016 ( \32780_33080 , \32775_33075 , \32779_33079 );
and \U$24017 ( \32781_33081 , \32192_32491 , \32196_32495 );
and \U$24018 ( \32782_33082 , \32196_32495 , \32201_32500 );
and \U$24019 ( \32783_33083 , \32192_32491 , \32201_32500 );
or \U$24020 ( \32784_33084 , \32781_33081 , \32782_33082 , \32783_33083 );
xor \U$24021 ( \32785_33085 , \32780_33080 , \32784_33084 );
xor \U$24022 ( \32786_33086 , \32771_33071 , \32785_33085 );
and \U$24023 ( \32787_33087 , \25516_25815 , \15037_15336 );
and \U$24024 ( \32788_33088 , \26527_26829 , \14661_14963 );
nor \U$24025 ( \32789_33089 , \32787_33087 , \32788_33088 );
xnor \U$24026 ( \32790_33090 , \32789_33089 , \15043_15342 );
and \U$24027 ( \32791_33091 , \19259_19558 , \20706_21005 );
and \U$24028 ( \32792_33092 , \20242_20544 , \20255_20557 );
nor \U$24029 ( \32793_33093 , \32791_33091 , \32792_33092 );
xnor \U$24030 ( \32794_33094 , \32793_33093 , \20712_21011 );
xor \U$24031 ( \32795_33095 , \32790_33090 , \32794_33094 );
and \U$24032 ( \32796_33096 , \17736_18035 , \22243_22542 );
and \U$24033 ( \32797_33097 , \18730_19032 , \21801_22103 );
nor \U$24034 ( \32798_33098 , \32796_33096 , \32797_33097 );
xnor \U$24035 ( \32799_33099 , \32798_33098 , \22249_22548 );
xor \U$24036 ( \32800_33100 , \32795_33095 , \32799_33099 );
and \U$24037 ( \32801_33101 , \28782_29084 , \12491_12790 );
and \U$24038 ( \32802_33102 , \29966_30268 , \12159_12461 );
nor \U$24039 ( \32803_33103 , \32801_33101 , \32802_33102 );
xnor \U$24040 ( \32804_33104 , \32803_33103 , \12481_12780 );
and \U$24041 ( \32805_33105 , \23900_24199 , \16333_16635 );
and \U$24042 ( \32806_33106 , \24970_25272 , \15999_16301 );
nor \U$24043 ( \32807_33107 , \32805_33105 , \32806_33106 );
xnor \U$24044 ( \32808_33108 , \32807_33107 , \16323_16625 );
xor \U$24045 ( \32809_33109 , \32804_33104 , \32808_33108 );
and \U$24046 ( \32810_33110 , \16353_16655 , \23839_24138 );
and \U$24047 ( \32811_33111 , \17325_17627 , \23328_23630 );
nor \U$24048 ( \32812_33112 , \32810_33110 , \32811_33111 );
xnor \U$24049 ( \32813_33113 , \32812_33112 , \23845_24144 );
xor \U$24050 ( \32814_33114 , \32809_33109 , \32813_33113 );
xor \U$24051 ( \32815_33115 , \32800_33100 , \32814_33114 );
and \U$24052 ( \32816_33116 , \22257_22556 , \17791_18090 );
and \U$24053 ( \32817_33117 , \23315_23617 , \17353_17655 );
nor \U$24054 ( \32818_33118 , \32816_33116 , \32817_33117 );
xnor \U$24055 ( \32819_33119 , \32818_33118 , \17747_18046 );
and \U$24056 ( \32820_33120 , \15022_15321 , \25527_25826 );
and \U$24057 ( \32821_33121 , \15965_16267 , \24962_25264 );
nor \U$24058 ( \32822_33122 , \32820_33120 , \32821_33121 );
xnor \U$24059 ( \32823_33123 , \32822_33122 , \25474_25773 );
xor \U$24060 ( \32824_33124 , \32819_33119 , \32823_33123 );
and \U$24061 ( \32825_33125 , \13725_14024 , \27095_27397 );
and \U$24062 ( \32826_33126 , \14648_14950 , \26505_26807 );
nor \U$24063 ( \32827_33127 , \32825_33125 , \32826_33126 );
xnor \U$24064 ( \32828_33128 , \32827_33127 , \26993_27295 );
xor \U$24065 ( \32829_33129 , \32824_33124 , \32828_33128 );
xor \U$24066 ( \32830_33130 , \32815_33115 , \32829_33129 );
xor \U$24067 ( \32831_33131 , \32786_33086 , \32830_33130 );
xor \U$24068 ( \32832_33132 , \32767_33067 , \32831_33131 );
and \U$24069 ( \32833_33133 , \32213_32512 , \32227_32526 );
and \U$24070 ( \32834_33134 , \32227_32526 , \32518_32817 );
and \U$24071 ( \32835_33135 , \32213_32512 , \32518_32817 );
or \U$24072 ( \32836_33136 , \32833_33133 , \32834_33134 , \32835_33135 );
and \U$24073 ( \32837_33137 , \32524_32823 , \32528_32827 );
and \U$24074 ( \32838_33138 , \32528_32827 , \32576_32875 );
and \U$24075 ( \32839_33139 , \32524_32823 , \32576_32875 );
or \U$24076 ( \32840_33140 , \32837_33137 , \32838_33138 , \32839_33139 );
xor \U$24077 ( \32841_33141 , \32836_33136 , \32840_33140 );
and \U$24078 ( \32842_33142 , \32217_32516 , \32221_32520 );
and \U$24079 ( \32843_33143 , \32221_32520 , \32226_32525 );
and \U$24080 ( \32844_33144 , \32217_32516 , \32226_32525 );
or \U$24081 ( \32845_33145 , \32842_33142 , \32843_33143 , \32844_33144 );
and \U$24082 ( \32846_33146 , \27011_27313 , \13755_14054 );
and \U$24083 ( \32847_33147 , \28232_28534 , \13390_13692 );
nor \U$24084 ( \32848_33148 , \32846_33146 , \32847_33147 );
xnor \U$24085 ( \32849_33149 , \32848_33148 , \13736_14035 );
and \U$24086 ( \32850_33150 , \20734_21033 , \19235_19534 );
and \U$24087 ( \32851_33151 , \21788_22090 , \18743_19045 );
nor \U$24088 ( \32852_33152 , \32850_33150 , \32851_33151 );
xnor \U$24089 ( \32853_33153 , \32852_33152 , \19241_19540 );
xor \U$24090 ( \32854_33154 , \32849_33149 , \32853_33153 );
and \U$24091 ( \32855_33155 , \10686_10988 , \32555_32854 );
and \U$24092 ( \32856_33156 , \10968_11270 , \31765_32067 );
nor \U$24093 ( \32857_33157 , \32855_33155 , \32856_33156 );
xnor \U$24094 ( \32858_33158 , \32857_33157 , \32506_32805 );
xor \U$24095 ( \32859_33159 , \32854_33154 , \32858_33158 );
xor \U$24096 ( \32860_33160 , \32845_33145 , \32859_33159 );
and \U$24097 ( \32861_33161 , \32498_32797 , \32507_32806 );
and \U$24098 ( \32862_33162 , \12470_12769 , \28768_29070 );
and \U$24099 ( \32863_33163 , \13377_13679 , \28224_28526 );
nor \U$24100 ( \32864_33164 , \32862_33162 , \32863_33163 );
xnor \U$24101 ( \32865_33165 , \32864_33164 , \28774_29076 );
xor \U$24102 ( \32866_33166 , \32861_33161 , \32865_33165 );
and \U$24103 ( \32867_33167 , \11287_11586 , \30521_30823 );
and \U$24104 ( \32868_33168 , \12146_12448 , \29944_30246 );
nor \U$24105 ( \32869_33169 , \32867_33167 , \32868_33168 );
xnor \U$24106 ( \32870_33170 , \32869_33169 , \30511_30813 );
xor \U$24107 ( \32871_33171 , \32866_33166 , \32870_33170 );
xor \U$24108 ( \32872_33172 , \32860_33160 , \32871_33171 );
xor \U$24109 ( \32873_33173 , \32841_33141 , \32872_33172 );
xor \U$24110 ( \32874_33174 , \32832_33132 , \32873_33173 );
xor \U$24111 ( \32875_33175 , \32737_33037 , \32874_33174 );
xor \U$24112 ( \32876_33176 , \32728_33028 , \32875_33175 );
and \U$24113 ( \32877_33177 , \32579_32878 , \32583_32882 );
and \U$24114 ( \32878_33178 , \32584_32883 , \32587_32886 );
or \U$24115 ( \32879_33179 , \32877_33177 , \32878_33178 );
xor \U$24116 ( \32880_33180 , \32876_33176 , \32879_33179 );
buf g9bae_GF_PartitionCandidate( \32881_33181_nG9bae , \32880_33180 );
and \U$24117 ( \32882_33182 , \10402_10704 , \32881_33181_nG9bae );
or \U$24118 ( \32883_33183 , \32724_33024 , \32882_33182 );
xor \U$24119 ( \32884_33184 , \10399_10703 , \32883_33183 );
buf \U$24120 ( \32885_33185 , \32884_33184 );
buf \U$24122 ( \32886_33186 , \32885_33185 );
xor \U$24123 ( \32887_33187 , \32723_33023 , \32886_33186 );
buf \U$24124 ( \32888_33188 , \32887_33187 );
xor \U$24125 ( \32889_33189 , \32634_32934 , \32888_33188 );
and \U$24126 ( \32890_33190 , \32130_32429 , \32135_32434 );
and \U$24127 ( \32891_33191 , \32130_32429 , \32141_32440 );
and \U$24128 ( \32892_33192 , \32135_32434 , \32141_32440 );
or \U$24129 ( \32893_33193 , \32890_33190 , \32891_33191 , \32892_33192 );
buf \U$24130 ( \32894_33194 , \32893_33193 );
xor \U$24131 ( \32895_33195 , \32889_33189 , \32894_33194 );
buf \U$24132 ( \32896_33196 , \32895_33195 );
and \U$24133 ( \32897_33197 , \31970_32272 , \32071_32370 );
and \U$24134 ( \32898_33198 , \31970_32272 , \32077_32376 );
and \U$24135 ( \32899_33199 , \32071_32370 , \32077_32376 );
or \U$24136 ( \32900_33200 , \32897_33197 , \32898_33198 , \32899_33199 );
buf \U$24137 ( \32901_33201 , \32900_33200 );
xor \U$24138 ( \32902_33202 , \32896_33196 , \32901_33201 );
and \U$24139 ( \32903_33203 , \32143_32442 , \32596_32895 );
and \U$24140 ( \32904_33204 , \32143_32442 , \32602_32901 );
and \U$24141 ( \32905_33205 , \32596_32895 , \32602_32901 );
or \U$24142 ( \32906_33206 , \32903_33203 , \32904_33204 , \32905_33205 );
buf \U$24143 ( \32907_33207 , \32906_33206 );
and \U$24144 ( \32908_33208 , \32028_32327 , \32034_32333 );
and \U$24145 ( \32909_33209 , \32028_32327 , \32041_32340 );
and \U$24146 ( \32910_33210 , \32034_32333 , \32041_32340 );
or \U$24147 ( \32911_33211 , \32908_33208 , \32909_33209 , \32910_33210 );
buf \U$24148 ( \32912_33212 , \32911_33211 );
and \U$24149 ( \32913_33213 , \32148_32447 , \32154_32453 );
and \U$24150 ( \32914_33214 , \32148_32447 , \32594_32893 );
and \U$24151 ( \32915_33215 , \32154_32453 , \32594_32893 );
or \U$24152 ( \32916_33216 , \32913_33213 , \32914_33214 , \32915_33215 );
buf \U$24153 ( \32917_33217 , \32916_33216 );
xor \U$24154 ( \32918_33218 , \32912_33212 , \32917_33217 );
and \U$24155 ( \32919_33219 , \13431_13370 , \27114_27416_nG9bc3 );
and \U$24156 ( \32920_33220 , \13068_13367 , \28300_28602_nG9bc0 );
or \U$24157 ( \32921_33221 , \32919_33219 , \32920_33220 );
xor \U$24158 ( \32922_33222 , \13067_13366 , \32921_33221 );
buf \U$24159 ( \32923_33223 , \32922_33222 );
buf \U$24161 ( \32924_33224 , \32923_33223 );
and \U$24162 ( \32925_33225 , \12183_12157 , \28877_29179_nG9bbd );
and \U$24163 ( \32926_33226 , \11855_12154 , \30064_30366_nG9bba );
or \U$24164 ( \32927_33227 , \32925_33225 , \32926_33226 );
xor \U$24165 ( \32928_33228 , \11854_12153 , \32927_33227 );
buf \U$24166 ( \32929_33229 , \32928_33228 );
buf \U$24168 ( \32930_33230 , \32929_33229 );
xor \U$24169 ( \32931_33231 , \32924_33224 , \32930_33230 );
and \U$24170 ( \32932_33232 , \10996_10421 , \30638_30940_nG9bb7 );
and \U$24171 ( \32933_33233 , \10119_10418 , \31877_32179_nG9bb4 );
or \U$24172 ( \32934_33234 , \32932_33232 , \32933_33233 );
xor \U$24173 ( \32935_33235 , \10118_10417 , \32934_33234 );
buf \U$24174 ( \32936_33236 , \32935_33235 );
buf \U$24176 ( \32937_33237 , \32936_33236 );
xor \U$24177 ( \32938_33238 , \32931_33231 , \32937_33237 );
buf \U$24178 ( \32939_33239 , \32938_33238 );
xor \U$24179 ( \32940_33240 , \32918_33218 , \32939_33239 );
buf \U$24180 ( \32941_33241 , \32940_33240 );
xor \U$24181 ( \32942_33242 , \32907_33207 , \32941_33241 );
and \U$24182 ( \32943_33243 , \32116_32415 , \32121_32420 );
and \U$24183 ( \32944_33244 , \32116_32415 , \32128_32427 );
and \U$24184 ( \32945_33245 , \32121_32420 , \32128_32427 );
or \U$24185 ( \32946_33246 , \32943_33243 , \32944_33244 , \32945_33245 );
buf \U$24186 ( \32947_33247 , \32946_33246 );
and \U$24187 ( \32948_33248 , \32013_32312 , \32019_32318 );
and \U$24188 ( \32949_33249 , \32013_32312 , \32026_32325 );
and \U$24189 ( \32950_33250 , \32019_32318 , \32026_32325 );
or \U$24190 ( \32951_33251 , \32948_33248 , \32949_33249 , \32950_33250 );
buf \U$24191 ( \32952_33252 , \32951_33251 );
and \U$24192 ( \32953_33253 , \32092_32391 , \32098_32397 );
and \U$24193 ( \32954_33254 , \32092_32391 , \32105_32404 );
and \U$24194 ( \32955_33255 , \32098_32397 , \32105_32404 );
or \U$24195 ( \32956_33256 , \32953_33253 , \32954_33254 , \32955_33255 );
buf \U$24196 ( \32957_33257 , \32956_33256 );
and \U$24197 ( \32958_33258 , \20353_20155 , \19287_19586_nG9be1 );
and \U$24198 ( \32959_33259 , \19853_20152 , \20306_20608_nG9bde );
or \U$24199 ( \32960_33260 , \32958_33258 , \32959_33259 );
xor \U$24200 ( \32961_33261 , \19852_20151 , \32960_33260 );
buf \U$24201 ( \32962_33262 , \32961_33261 );
buf \U$24203 ( \32963_33263 , \32962_33262 );
xor \U$24204 ( \32964_33264 , \32957_33257 , \32963_33263 );
and \U$24205 ( \32965_33265 , \18908_18702 , \20787_21086_nG9bdb );
and \U$24206 ( \32966_33266 , \18400_18699 , \21827_22129_nG9bd8 );
or \U$24207 ( \32967_33267 , \32965_33265 , \32966_33266 );
xor \U$24208 ( \32968_33268 , \18399_18698 , \32967_33267 );
buf \U$24209 ( \32969_33269 , \32968_33268 );
buf \U$24211 ( \32970_33270 , \32969_33269 );
xor \U$24212 ( \32971_33271 , \32964_33264 , \32970_33270 );
buf \U$24213 ( \32972_33272 , \32971_33271 );
xor \U$24214 ( \32973_33273 , \32952_33252 , \32972_33272 );
and \U$24215 ( \32974_33274 , \14710_14631 , \25561_25860_nG9bc9 );
and \U$24216 ( \32975_33275 , \14329_14628 , \26585_26887_nG9bc6 );
or \U$24217 ( \32976_33276 , \32974_33274 , \32975_33275 );
xor \U$24218 ( \32977_33277 , \14328_14627 , \32976_33276 );
buf \U$24219 ( \32978_33278 , \32977_33277 );
buf \U$24221 ( \32979_33279 , \32978_33278 );
xor \U$24222 ( \32980_33280 , \32973_33273 , \32979_33279 );
buf \U$24223 ( \32981_33281 , \32980_33280 );
xor \U$24224 ( \32982_33282 , \32947_33247 , \32981_33281 );
and \U$24225 ( \32983_33283 , \32048_32347 , \32054_32353 );
and \U$24226 ( \32984_33284 , \32048_32347 , \32061_32360 );
and \U$24227 ( \32985_33285 , \32054_32353 , \32061_32360 );
or \U$24228 ( \32986_33286 , \32983_33283 , \32984_33284 , \32985_33285 );
buf \U$24229 ( \32987_33287 , \32986_33286 );
xor \U$24230 ( \32988_33288 , \32982_33282 , \32987_33287 );
buf \U$24231 ( \32989_33289 , \32988_33288 );
xor \U$24232 ( \32990_33290 , \32942_33242 , \32989_33289 );
buf \U$24233 ( \32991_33291 , \32990_33290 );
xor \U$24234 ( \32992_33292 , \32902_33202 , \32991_33291 );
and \U$24235 ( \32993_33293 , \32624_32924 , \32992_33292 );
and \U$24236 ( \32994_33294 , \32628_32928 , \32992_33292 );
or \U$24237 ( \32995_33295 , \32629_32929 , \32993_33293 , \32994_33294 );
and \U$24238 ( \32996_33296 , \32611_32910 , \32615_32914 );
and \U$24239 ( \32997_33297 , \32611_32910 , \32623_32923 );
and \U$24240 ( \32998_33298 , \32615_32914 , \32623_32923 );
or \U$24241 ( \32999_33299 , \32996_33296 , \32997_33297 , \32998_33298 );
xor \U$24242 ( \33000_33300 , \32995_33295 , \32999_33299 );
xor \U$24246 ( \33001_33301 , \33000_33300 , 1'b0 );
and \U$24247 ( \33002_33302 , \32907_33207 , \32941_33241 );
and \U$24248 ( \33003_33303 , \32907_33207 , \32989_33289 );
and \U$24249 ( \33004_33304 , \32941_33241 , \32989_33289 );
or \U$24250 ( \33005_33305 , \33002_33302 , \33003_33303 , \33004_33304 );
buf \U$24251 ( \33006_33306 , \33005_33305 );
and \U$24252 ( \33007_33307 , \32690_32990 , \32704_33004 );
and \U$24253 ( \33008_33308 , \32690_32990 , \32711_33011 );
and \U$24254 ( \33009_33309 , \32704_33004 , \32711_33011 );
or \U$24255 ( \33010_33310 , \33007_33307 , \33008_33308 , \33009_33309 );
buf \U$24256 ( \33011_33311 , \33010_33310 );
and \U$24257 ( \33012_33312 , \32696_32996 , \32702_33002 );
buf \U$24258 ( \33013_33313 , \33012_33312 );
and \U$24259 ( \33014_33314 , \28946_28118 , \13403_13705_nG9bfc );
and \U$24260 ( \33015_33315 , \27816_28115 , \13771_14070_nG9bf9 );
or \U$24261 ( \33016_33316 , \33014_33314 , \33015_33315 );
xor \U$24262 ( \33017_33317 , \27815_28114 , \33016_33316 );
buf \U$24263 ( \33018_33318 , \33017_33317 );
buf \U$24265 ( \33019_33319 , \33018_33318 );
xor \U$24266 ( \33020_33320 , \33013_33313 , \33019_33319 );
and \U$24267 ( \33021_33321 , \27141_26431 , \14682_14984_nG9bf6 );
and \U$24268 ( \33022_33322 , \26129_26428 , \15074_15373_nG9bf3 );
or \U$24269 ( \33023_33323 , \33021_33321 , \33022_33322 );
xor \U$24270 ( \33024_33324 , \26128_26427 , \33023_33323 );
buf \U$24271 ( \33025_33325 , \33024_33324 );
buf \U$24273 ( \33026_33326 , \33025_33325 );
xor \U$24274 ( \33027_33327 , \33020_33320 , \33026_33326 );
buf \U$24275 ( \33028_33328 , \33027_33327 );
xor \U$24276 ( \33029_33329 , \33011_33311 , \33028_33328 );
and \U$24277 ( \33030_33330 , \23495_23201 , \17363_17665_nG9bea );
and \U$24278 ( \33031_33331 , \22899_23198 , \17808_18107_nG9be7 );
or \U$24279 ( \33032_33332 , \33030_33330 , \33031_33331 );
xor \U$24280 ( \33033_33333 , \22898_23197 , \33032_33332 );
buf \U$24281 ( \33034_33334 , \33033_33333 );
buf \U$24283 ( \33035_33335 , \33034_33334 );
xor \U$24284 ( \33036_33336 , \33029_33329 , \33035_33335 );
buf \U$24285 ( \33037_33337 , \33036_33336 );
and \U$24286 ( \33038_33338 , \32641_32941 , \32647_32947 );
and \U$24287 ( \33039_33339 , \32641_32941 , \32654_32954 );
and \U$24288 ( \33040_33340 , \32647_32947 , \32654_32954 );
or \U$24289 ( \33041_33341 , \33038_33338 , \33039_33339 , \33040_33340 );
buf \U$24290 ( \33042_33342 , \33041_33341 );
and \U$24292 ( \33043_33343 , \32617_32916 , \10693_10995_nG9c0b );
or \U$24293 ( \33044_33344 , 1'b0 , \33043_33343 );
xor \U$24294 ( \33045_33345 , 1'b0 , \33044_33344 );
buf \U$24295 ( \33046_33346 , \33045_33345 );
buf \U$24297 ( \33047_33347 , \33046_33346 );
and \U$24298 ( \33048_33348 , \31989_31636 , \10981_11283_nG9c08 );
and \U$24299 ( \33049_33349 , \31334_31633 , \11299_11598_nG9c05 );
or \U$24300 ( \33050_33350 , \33048_33348 , \33049_33349 );
xor \U$24301 ( \33051_33351 , \31333_31632 , \33050_33350 );
buf \U$24302 ( \33052_33352 , \33051_33351 );
buf \U$24304 ( \33053_33353 , \33052_33352 );
xor \U$24305 ( \33054_33354 , \33047_33347 , \33053_33353 );
and \U$24306 ( \33055_33355 , \30670_29853 , \12168_12470_nG9c02 );
and \U$24307 ( \33056_33356 , \29551_29850 , \12502_12801_nG9bff );
or \U$24308 ( \33057_33357 , \33055_33355 , \33056_33356 );
xor \U$24309 ( \33058_33358 , \29550_29849 , \33057_33357 );
buf \U$24310 ( \33059_33359 , \33058_33358 );
buf \U$24312 ( \33060_33360 , \33059_33359 );
xor \U$24313 ( \33061_33361 , \33054_33354 , \33060_33360 );
buf \U$24314 ( \33062_33362 , \33061_33361 );
xor \U$24315 ( \33063_33363 , \33042_33342 , \33062_33362 );
and \U$24316 ( \33064_33364 , \25044_24792 , \16013_16315_nG9bf0 );
and \U$24317 ( \33065_33365 , \24490_24789 , \16378_16680_nG9bed );
or \U$24318 ( \33066_33366 , \33064_33364 , \33065_33365 );
xor \U$24319 ( \33067_33367 , \24489_24788 , \33066_33366 );
buf \U$24320 ( \33068_33368 , \33067_33367 );
buf \U$24322 ( \33069_33369 , \33068_33368 );
xor \U$24323 ( \33070_33370 , \33063_33363 , \33069_33369 );
buf \U$24324 ( \33071_33371 , \33070_33370 );
and \U$24325 ( \33072_33372 , \21908_21658 , \18789_19091_nG9be4 );
and \U$24326 ( \33073_33373 , \21356_21655 , \19287_19586_nG9be1 );
or \U$24327 ( \33074_33374 , \33072_33372 , \33073_33373 );
xor \U$24328 ( \33075_33375 , \21355_21654 , \33074_33374 );
buf \U$24329 ( \33076_33376 , \33075_33375 );
buf \U$24331 ( \33077_33377 , \33076_33376 );
xor \U$24332 ( \33078_33378 , \33071_33371 , \33077_33377 );
and \U$24333 ( \33079_33379 , \20353_20155 , \20306_20608_nG9bde );
and \U$24334 ( \33080_33380 , \19853_20152 , \20787_21086_nG9bdb );
or \U$24335 ( \33081_33381 , \33079_33379 , \33080_33380 );
xor \U$24336 ( \33082_33382 , \19852_20151 , \33081_33381 );
buf \U$24337 ( \33083_33383 , \33082_33382 );
buf \U$24339 ( \33084_33384 , \33083_33383 );
xor \U$24340 ( \33085_33385 , \33078_33378 , \33084_33384 );
buf \U$24341 ( \33086_33386 , \33085_33385 );
xor \U$24342 ( \33087_33387 , \33037_33337 , \33086_33386 );
and \U$24343 ( \33088_33388 , \32957_33257 , \32963_33263 );
and \U$24344 ( \33089_33389 , \32957_33257 , \32970_33270 );
and \U$24345 ( \33090_33390 , \32963_33263 , \32970_33270 );
or \U$24346 ( \33091_33391 , \33088_33388 , \33089_33389 , \33090_33390 );
buf \U$24347 ( \33092_33392 , \33091_33391 );
xor \U$24348 ( \33093_33393 , \33087_33387 , \33092_33392 );
buf \U$24349 ( \33094_33394 , \33093_33393 );
and \U$24350 ( \33095_33395 , \32952_33252 , \32972_33272 );
and \U$24351 ( \33096_33396 , \32952_33252 , \32979_33279 );
and \U$24352 ( \33097_33397 , \32972_33272 , \32979_33279 );
or \U$24353 ( \33098_33398 , \33095_33395 , \33096_33396 , \33097_33397 );
buf \U$24354 ( \33099_33399 , \33098_33398 );
xor \U$24355 ( \33100_33400 , \33094_33394 , \33099_33399 );
and \U$24356 ( \33101_33401 , \16405_15940 , \24996_25298_nG9bcc );
and \U$24357 ( \33102_33402 , \15638_15937 , \25561_25860_nG9bc9 );
or \U$24358 ( \33103_33403 , \33101_33401 , \33102_33402 );
xor \U$24359 ( \33104_33404 , \15637_15936 , \33103_33403 );
buf \U$24360 ( \33105_33405 , \33104_33404 );
buf \U$24362 ( \33106_33406 , \33105_33405 );
and \U$24363 ( \33107_33407 , \14710_14631 , \26585_26887_nG9bc6 );
and \U$24364 ( \33108_33408 , \14329_14628 , \27114_27416_nG9bc3 );
or \U$24365 ( \33109_33409 , \33107_33407 , \33108_33408 );
xor \U$24366 ( \33110_33410 , \14328_14627 , \33109_33409 );
buf \U$24367 ( \33111_33411 , \33110_33410 );
buf \U$24369 ( \33112_33412 , \33111_33411 );
xor \U$24370 ( \33113_33413 , \33106_33406 , \33112_33412 );
and \U$24371 ( \33114_33414 , \12183_12157 , \30064_30366_nG9bba );
and \U$24372 ( \33115_33415 , \11855_12154 , \30638_30940_nG9bb7 );
or \U$24373 ( \33116_33416 , \33114_33414 , \33115_33415 );
xor \U$24374 ( \33117_33417 , \11854_12153 , \33116_33416 );
buf \U$24375 ( \33118_33418 , \33117_33417 );
buf \U$24377 ( \33119_33419 , \33118_33418 );
xor \U$24378 ( \33120_33420 , \33113_33413 , \33119_33419 );
buf \U$24379 ( \33121_33421 , \33120_33420 );
xor \U$24380 ( \33122_33422 , \33100_33400 , \33121_33421 );
buf \U$24381 ( \33123_33423 , \33122_33422 );
and \U$24382 ( \33124_33424 , \32947_33247 , \32981_33281 );
and \U$24383 ( \33125_33425 , \32947_33247 , \32987_33287 );
and \U$24384 ( \33126_33426 , \32981_33281 , \32987_33287 );
or \U$24385 ( \33127_33427 , \33124_33424 , \33125_33425 , \33126_33426 );
buf \U$24386 ( \33128_33428 , \33127_33427 );
xor \U$24387 ( \33129_33429 , \33123_33423 , \33128_33428 );
and \U$24388 ( \33130_33430 , \32656_32956 , \32662_32962 );
and \U$24389 ( \33131_33431 , \32656_32956 , \32669_32969 );
and \U$24390 ( \33132_33432 , \32662_32962 , \32669_32969 );
or \U$24391 ( \33133_33433 , \33130_33430 , \33131_33431 , \33132_33432 );
buf \U$24392 ( \33134_33434 , \33133_33433 );
and \U$24393 ( \33135_33435 , \18908_18702 , \21827_22129_nG9bd8 );
and \U$24394 ( \33136_33436 , \18400_18699 , \22330_22629_nG9bd5 );
or \U$24395 ( \33137_33437 , \33135_33435 , \33136_33436 );
xor \U$24396 ( \33138_33438 , \18399_18698 , \33137_33437 );
buf \U$24397 ( \33139_33439 , \33138_33438 );
buf \U$24399 ( \33140_33440 , \33139_33439 );
xor \U$24400 ( \33141_33441 , \33134_33434 , \33140_33440 );
and \U$24401 ( \33142_33442 , \17437_17297 , \23394_23696_nG9bd2 );
and \U$24402 ( \33143_33443 , \16995_17294 , \23927_24226_nG9bcf );
or \U$24403 ( \33144_33444 , \33142_33442 , \33143_33443 );
xor \U$24404 ( \33145_33445 , \16994_17293 , \33144_33444 );
buf \U$24405 ( \33146_33446 , \33145_33445 );
buf \U$24407 ( \33147_33447 , \33146_33446 );
xor \U$24408 ( \33148_33448 , \33141_33441 , \33147_33447 );
buf \U$24409 ( \33149_33449 , \33148_33448 );
and \U$24410 ( \33150_33450 , \32639_32939 , \32671_32971 );
and \U$24411 ( \33151_33451 , \32639_32939 , \32678_32978 );
and \U$24412 ( \33152_33452 , \32671_32971 , \32678_32978 );
or \U$24413 ( \33153_33453 , \33150_33450 , \33151_33451 , \33152_33452 );
buf \U$24414 ( \33154_33454 , \33153_33453 );
xor \U$24415 ( \33155_33455 , \33149_33449 , \33154_33454 );
and \U$24416 ( \33156_33456 , \10411_10707 , \32881_33181_nG9bae );
and \U$24417 ( \33157_33457 , \32767_33067 , \32831_33131 );
and \U$24418 ( \33158_33458 , \32831_33131 , \32873_33173 );
and \U$24419 ( \33159_33459 , \32767_33067 , \32873_33173 );
or \U$24420 ( \33160_33460 , \33157_33457 , \33158_33458 , \33159_33459 );
and \U$24421 ( \33161_33461 , \32741_33041 , \32745_33045 );
and \U$24422 ( \33162_33462 , \32745_33045 , \32766_33066 );
and \U$24423 ( \33163_33463 , \32741_33041 , \32766_33066 );
or \U$24424 ( \33164_33464 , \33161_33461 , \33162_33462 , \33163_33463 );
and \U$24425 ( \33165_33465 , \32861_33161 , \32865_33165 );
and \U$24426 ( \33166_33466 , \32865_33165 , \32870_33170 );
and \U$24427 ( \33167_33467 , \32861_33161 , \32870_33170 );
or \U$24428 ( \33168_33468 , \33165_33465 , \33166_33466 , \33167_33467 );
and \U$24429 ( \33169_33469 , \32775_33075 , \32779_33079 );
and \U$24430 ( \33170_33470 , \32779_33079 , \32784_33084 );
and \U$24431 ( \33171_33471 , \32775_33075 , \32784_33084 );
or \U$24432 ( \33172_33472 , \33169_33469 , \33170_33470 , \33171_33471 );
xor \U$24433 ( \33173_33473 , \33168_33468 , \33172_33472 );
and \U$24434 ( \33174_33474 , \32750_33050 , \32754_33054 );
and \U$24435 ( \33175_33475 , \32754_33054 , \32765_33065 );
and \U$24436 ( \33176_33476 , \32750_33050 , \32765_33065 );
or \U$24437 ( \33177_33477 , \33174_33474 , \33175_33475 , \33176_33476 );
xor \U$24438 ( \33178_33478 , \33173_33473 , \33177_33477 );
xor \U$24439 ( \33179_33479 , \33164_33464 , \33178_33478 );
and \U$24440 ( \33180_33480 , \32800_33100 , \32814_33114 );
and \U$24441 ( \33181_33481 , \32814_33114 , \32829_33129 );
and \U$24442 ( \33182_33482 , \32800_33100 , \32829_33129 );
or \U$24443 ( \33183_33483 , \33180_33480 , \33181_33481 , \33182_33482 );
and \U$24444 ( \33184_33484 , \32790_33090 , \32794_33094 );
and \U$24445 ( \33185_33485 , \32794_33094 , \32799_33099 );
and \U$24446 ( \33186_33486 , \32790_33090 , \32799_33099 );
or \U$24447 ( \33187_33487 , \33184_33484 , \33185_33485 , \33186_33486 );
and \U$24448 ( \33188_33488 , \32819_33119 , \32823_33123 );
and \U$24449 ( \33189_33489 , \32823_33123 , \32828_33128 );
and \U$24450 ( \33190_33490 , \32819_33119 , \32828_33128 );
or \U$24451 ( \33191_33491 , \33188_33488 , \33189_33489 , \33190_33490 );
xor \U$24452 ( \33192_33492 , \33187_33487 , \33191_33491 );
and \U$24453 ( \33193_33493 , \32849_33149 , \32853_33153 );
and \U$24454 ( \33194_33494 , \32853_33153 , \32858_33158 );
and \U$24455 ( \33195_33495 , \32849_33149 , \32858_33158 );
or \U$24456 ( \33196_33496 , \33193_33493 , \33194_33494 , \33195_33495 );
xor \U$24457 ( \33197_33497 , \33192_33492 , \33196_33496 );
xor \U$24458 ( \33198_33498 , \33183_33483 , \33197_33497 );
and \U$24459 ( \33199_33499 , \32758_33058 , \32762_33062 );
and \U$24460 ( \33200_33500 , \32762_33062 , \32764_33064 );
and \U$24461 ( \33201_33501 , \32758_33058 , \32764_33064 );
or \U$24462 ( \33202_33502 , \33199_33499 , \33200_33500 , \33201_33501 );
xor \U$24463 ( \33203_33503 , \33202_33502 , \10678_10980 );
and \U$24464 ( \33204_33504 , \12146_12448 , \30521_30823 );
and \U$24465 ( \33205_33505 , \12470_12769 , \29944_30246 );
nor \U$24466 ( \33206_33506 , \33204_33504 , \33205_33505 );
xnor \U$24467 ( \33207_33507 , \33206_33506 , \30511_30813 );
xor \U$24468 ( \33208_33508 , \33203_33503 , \33207_33507 );
xor \U$24469 ( \33209_33509 , \33198_33498 , \33208_33508 );
xor \U$24470 ( \33210_33510 , \33179_33479 , \33209_33509 );
xor \U$24471 ( \33211_33511 , \33160_33460 , \33210_33510 );
and \U$24472 ( \33212_33512 , \32771_33071 , \32785_33085 );
and \U$24473 ( \33213_33513 , \32785_33085 , \32830_33130 );
and \U$24474 ( \33214_33514 , \32771_33071 , \32830_33130 );
or \U$24475 ( \33215_33515 , \33212_33512 , \33213_33513 , \33214_33514 );
and \U$24476 ( \33216_33516 , \32836_33136 , \32840_33140 );
and \U$24477 ( \33217_33517 , \32840_33140 , \32872_33172 );
and \U$24478 ( \33218_33518 , \32836_33136 , \32872_33172 );
or \U$24479 ( \33219_33519 , \33216_33516 , \33217_33517 , \33218_33518 );
xor \U$24480 ( \33220_33520 , \33215_33515 , \33219_33519 );
and \U$24481 ( \33221_33521 , \32845_33145 , \32859_33159 );
and \U$24482 ( \33222_33522 , \32859_33159 , \32871_33171 );
and \U$24483 ( \33223_33523 , \32845_33145 , \32871_33171 );
or \U$24484 ( \33224_33524 , \33221_33521 , \33222_33522 , \33223_33523 );
and \U$24485 ( \33225_33525 , \32804_33104 , \32808_33108 );
and \U$24486 ( \33226_33526 , \32808_33108 , \32813_33113 );
and \U$24487 ( \33227_33527 , \32804_33104 , \32813_33113 );
or \U$24488 ( \33228_33528 , \33225_33525 , \33226_33526 , \33227_33527 );
and \U$24489 ( \33229_33529 , \21788_22090 , \19235_19534 );
and \U$24490 ( \33230_33530 , \22257_22556 , \18743_19045 );
nor \U$24491 ( \33231_33531 , \33229_33529 , \33230_33530 );
xnor \U$24492 ( \33232_33532 , \33231_33531 , \19241_19540 );
and \U$24493 ( \33233_33533 , \10968_11270 , \32555_32854 );
and \U$24494 ( \33234_33534 , \11287_11586 , \31765_32067 );
nor \U$24495 ( \33235_33535 , \33233_33533 , \33234_33534 );
xnor \U$24496 ( \33236_33536 , \33235_33535 , \32506_32805 );
xor \U$24497 ( \33237_33537 , \33232_33532 , \33236_33536 );
and \U$24498 ( \33238_33538 , \10686_10988 , \32503_32802 );
xor \U$24499 ( \33239_33539 , \33237_33537 , \33238_33538 );
xor \U$24500 ( \33240_33540 , \33228_33528 , \33239_33539 );
and \U$24501 ( \33241_33541 , \23315_23617 , \17791_18090 );
and \U$24502 ( \33242_33542 , \23900_24199 , \17353_17655 );
nor \U$24503 ( \33243_33543 , \33241_33541 , \33242_33542 );
xnor \U$24504 ( \33244_33544 , \33243_33543 , \17747_18046 );
and \U$24505 ( \33245_33545 , \14648_14950 , \27095_27397 );
and \U$24506 ( \33246_33546 , \15022_15321 , \26505_26807 );
nor \U$24507 ( \33247_33547 , \33245_33545 , \33246_33546 );
xnor \U$24508 ( \33248_33548 , \33247_33547 , \26993_27295 );
xor \U$24509 ( \33249_33549 , \33244_33544 , \33248_33548 );
and \U$24510 ( \33250_33550 , \13377_13679 , \28768_29070 );
and \U$24511 ( \33251_33551 , \13725_14024 , \28224_28526 );
nor \U$24512 ( \33252_33552 , \33250_33550 , \33251_33551 );
xnor \U$24513 ( \33253_33553 , \33252_33552 , \28774_29076 );
xor \U$24514 ( \33254_33554 , \33249_33549 , \33253_33553 );
xor \U$24515 ( \33255_33555 , \33240_33540 , \33254_33554 );
xor \U$24516 ( \33256_33556 , \33224_33524 , \33255_33555 );
and \U$24517 ( \33257_33557 , \31752_32054 , \11275_11574 );
and \U$24518 ( \33258_33558 , \32495_32794 , \10976_11278 );
nor \U$24519 ( \33259_33559 , \33257_33557 , \33258_33558 );
xnor \U$24520 ( \33260_33560 , \33259_33559 , \11281_11580 );
and \U$24521 ( \33261_33561 , \28232_28534 , \13755_14054 );
and \U$24522 ( \33262_33562 , \28782_29084 , \13390_13692 );
nor \U$24523 ( \33263_33563 , \33261_33561 , \33262_33562 );
xnor \U$24524 ( \33264_33564 , \33263_33563 , \13736_14035 );
xor \U$24525 ( \33265_33565 , \33260_33560 , \33264_33564 );
and \U$24526 ( \33266_33566 , \20242_20544 , \20706_21005 );
and \U$24527 ( \33267_33567 , \20734_21033 , \20255_20557 );
nor \U$24528 ( \33268_33568 , \33266_33566 , \33267_33567 );
xnor \U$24529 ( \33269_33569 , \33268_33568 , \20712_21011 );
xor \U$24530 ( \33270_33570 , \33265_33565 , \33269_33569 );
and \U$24531 ( \33271_33571 , \26527_26829 , \15037_15336 );
and \U$24532 ( \33272_33572 , \27011_27313 , \14661_14963 );
nor \U$24533 ( \33273_33573 , \33271_33571 , \33272_33572 );
xnor \U$24534 ( \33274_33574 , \33273_33573 , \15043_15342 );
and \U$24535 ( \33275_33575 , \18730_19032 , \22243_22542 );
and \U$24536 ( \33276_33576 , \19259_19558 , \21801_22103 );
nor \U$24537 ( \33277_33577 , \33275_33575 , \33276_33576 );
xnor \U$24538 ( \33278_33578 , \33277_33577 , \22249_22548 );
xor \U$24539 ( \33279_33579 , \33274_33574 , \33278_33578 );
and \U$24540 ( \33280_33580 , \17325_17627 , \23839_24138 );
and \U$24541 ( \33281_33581 , \17736_18035 , \23328_23630 );
nor \U$24542 ( \33282_33582 , \33280_33580 , \33281_33581 );
xnor \U$24543 ( \33283_33583 , \33282_33582 , \23845_24144 );
xor \U$24544 ( \33284_33584 , \33279_33579 , \33283_33583 );
xor \U$24545 ( \33285_33585 , \33270_33570 , \33284_33584 );
and \U$24546 ( \33286_33586 , \29966_30268 , \12491_12790 );
and \U$24547 ( \33287_33587 , \30500_30802 , \12159_12461 );
nor \U$24548 ( \33288_33588 , \33286_33586 , \33287_33587 );
xnor \U$24549 ( \33289_33589 , \33288_33588 , \12481_12780 );
and \U$24550 ( \33290_33590 , \24970_25272 , \16333_16635 );
and \U$24551 ( \33291_33591 , \25516_25815 , \15999_16301 );
nor \U$24552 ( \33292_33592 , \33290_33590 , \33291_33591 );
xnor \U$24553 ( \33293_33593 , \33292_33592 , \16323_16625 );
xor \U$24554 ( \33294_33594 , \33289_33589 , \33293_33593 );
and \U$24555 ( \33295_33595 , \15965_16267 , \25527_25826 );
and \U$24556 ( \33296_33596 , \16353_16655 , \24962_25264 );
nor \U$24557 ( \33297_33597 , \33295_33595 , \33296_33596 );
xnor \U$24558 ( \33298_33598 , \33297_33597 , \25474_25773 );
xor \U$24559 ( \33299_33599 , \33294_33594 , \33298_33598 );
xor \U$24560 ( \33300_33600 , \33285_33585 , \33299_33599 );
xor \U$24561 ( \33301_33601 , \33256_33556 , \33300_33600 );
xor \U$24562 ( \33302_33602 , \33220_33520 , \33301_33601 );
xor \U$24563 ( \33303_33603 , \33211_33511 , \33302_33602 );
and \U$24564 ( \33304_33604 , \32732_33032 , \32736_33036 );
and \U$24565 ( \33305_33605 , \32736_33036 , \32874_33174 );
and \U$24566 ( \33306_33606 , \32732_33032 , \32874_33174 );
or \U$24567 ( \33307_33607 , \33304_33604 , \33305_33605 , \33306_33606 );
xor \U$24568 ( \33308_33608 , \33303_33603 , \33307_33607 );
and \U$24569 ( \33309_33609 , \32728_33028 , \32875_33175 );
and \U$24570 ( \33310_33610 , \32876_33176 , \32879_33179 );
or \U$24571 ( \33311_33611 , \33309_33609 , \33310_33610 );
xor \U$24572 ( \33312_33612 , \33308_33608 , \33311_33611 );
buf g9bab_GF_PartitionCandidate( \33313_33613_nG9bab , \33312_33612 );
and \U$24573 ( \33314_33614 , \10402_10704 , \33313_33613_nG9bab );
or \U$24574 ( \33315_33615 , \33156_33456 , \33314_33614 );
xor \U$24575 ( \33316_33616 , \10399_10703 , \33315_33615 );
buf \U$24576 ( \33317_33617 , \33316_33616 );
buf \U$24578 ( \33318_33618 , \33317_33617 );
xor \U$24579 ( \33319_33619 , \33155_33455 , \33318_33618 );
buf \U$24580 ( \33320_33620 , \33319_33619 );
xor \U$24581 ( \33321_33621 , \33129_33429 , \33320_33620 );
buf \U$24582 ( \33322_33622 , \33321_33621 );
xor \U$24583 ( \33323_33623 , \33006_33306 , \33322_33622 );
and \U$24584 ( \33324_33624 , \32634_32934 , \32888_33188 );
and \U$24585 ( \33325_33625 , \32634_32934 , \32894_33194 );
and \U$24586 ( \33326_33626 , \32888_33188 , \32894_33194 );
or \U$24587 ( \33327_33627 , \33324_33624 , \33325_33625 , \33326_33626 );
buf \U$24588 ( \33328_33628 , \33327_33627 );
and \U$24589 ( \33329_33629 , \32680_32980 , \32722_33022 );
and \U$24590 ( \33330_33630 , \32680_32980 , \32886_33186 );
and \U$24591 ( \33331_33631 , \32722_33022 , \32886_33186 );
or \U$24592 ( \33332_33632 , \33329_33629 , \33330_33630 , \33331_33631 );
buf \U$24593 ( \33333_33633 , \33332_33632 );
and \U$24594 ( \33334_33634 , \32924_33224 , \32930_33230 );
and \U$24595 ( \33335_33635 , \32924_33224 , \32937_33237 );
and \U$24596 ( \33336_33636 , \32930_33230 , \32937_33237 );
or \U$24597 ( \33337_33637 , \33334_33634 , \33335_33635 , \33336_33636 );
buf \U$24598 ( \33338_33638 , \33337_33637 );
xor \U$24599 ( \33339_33639 , \33333_33633 , \33338_33638 );
and \U$24600 ( \33340_33640 , \32685_32985 , \32713_33013 );
and \U$24601 ( \33341_33641 , \32685_32985 , \32720_33020 );
and \U$24602 ( \33342_33642 , \32713_33013 , \32720_33020 );
or \U$24603 ( \33343_33643 , \33340_33640 , \33341_33641 , \33342_33642 );
buf \U$24604 ( \33344_33644 , \33343_33643 );
and \U$24605 ( \33345_33645 , \13431_13370 , \28300_28602_nG9bc0 );
and \U$24606 ( \33346_33646 , \13068_13367 , \28877_29179_nG9bbd );
or \U$24607 ( \33347_33647 , \33345_33645 , \33346_33646 );
xor \U$24608 ( \33348_33648 , \13067_13366 , \33347_33647 );
buf \U$24609 ( \33349_33649 , \33348_33648 );
buf \U$24611 ( \33350_33650 , \33349_33649 );
xor \U$24612 ( \33351_33651 , \33344_33644 , \33350_33650 );
and \U$24613 ( \33352_33652 , \10996_10421 , \31877_32179_nG9bb4 );
and \U$24614 ( \33353_33653 , \10119_10418 , \32589_32888_nG9bb1 );
or \U$24615 ( \33354_33654 , \33352_33652 , \33353_33653 );
xor \U$24616 ( \33355_33655 , \10118_10417 , \33354_33654 );
buf \U$24617 ( \33356_33656 , \33355_33655 );
buf \U$24619 ( \33357_33657 , \33356_33656 );
xor \U$24620 ( \33358_33658 , \33351_33651 , \33357_33657 );
buf \U$24621 ( \33359_33659 , \33358_33658 );
xor \U$24622 ( \33360_33660 , \33339_33639 , \33359_33659 );
buf \U$24623 ( \33361_33661 , \33360_33660 );
xor \U$24624 ( \33362_33662 , \33328_33628 , \33361_33661 );
and \U$24625 ( \33363_33663 , \32912_33212 , \32917_33217 );
and \U$24626 ( \33364_33664 , \32912_33212 , \32939_33239 );
and \U$24627 ( \33365_33665 , \32917_33217 , \32939_33239 );
or \U$24628 ( \33366_33666 , \33363_33663 , \33364_33664 , \33365_33665 );
buf \U$24629 ( \33367_33667 , \33366_33666 );
xor \U$24630 ( \33368_33668 , \33362_33662 , \33367_33667 );
buf \U$24631 ( \33369_33669 , \33368_33668 );
xor \U$24632 ( \33370_33670 , \33323_33623 , \33369_33669 );
and \U$24633 ( \33371_33671 , \33001_33301 , \33370_33670 );
and \U$24634 ( \33372_33672 , \32896_33196 , \32901_33201 );
and \U$24635 ( \33373_33673 , \32896_33196 , \32991_33291 );
and \U$24636 ( \33374_33674 , \32901_33201 , \32991_33291 );
or \U$24637 ( \33375_33675 , \33372_33672 , \33373_33673 , \33374_33674 );
and \U$24638 ( \33376_33676 , \33001_33301 , \33375_33675 );
and \U$24639 ( \33377_33677 , \33370_33670 , \33375_33675 );
or \U$24640 ( \33378_33678 , \33371_33671 , \33376_33676 , \33377_33677 );
and \U$24641 ( \33379_33679 , \32995_33295 , \32999_33299 );
or \U$24644 ( \33380_33680 , \33379_33679 , 1'b0 , 1'b0 );
xor \U$24645 ( \33381_33681 , \33378_33678 , \33380_33680 );
xor \U$24659 ( \33382_33682 , \33381_33681 , 1'b0 );
and \U$24660 ( \33383_33683 , \33006_33306 , \33322_33622 );
and \U$24661 ( \33384_33684 , \33006_33306 , \33369_33669 );
and \U$24662 ( \33385_33685 , \33322_33622 , \33369_33669 );
or \U$24663 ( \33386_33686 , \33383_33683 , \33384_33684 , \33385_33685 );
and \U$24664 ( \33387_33687 , \33382_33682 , \33386_33686 );
and \U$24665 ( \33388_33688 , \33123_33423 , \33128_33428 );
and \U$24666 ( \33389_33689 , \33123_33423 , \33320_33620 );
and \U$24667 ( \33390_33690 , \33128_33428 , \33320_33620 );
or \U$24668 ( \33391_33691 , \33388_33688 , \33389_33689 , \33390_33690 );
buf \U$24669 ( \33392_33692 , \33391_33691 );
and \U$24670 ( \33393_33693 , \33149_33449 , \33154_33454 );
and \U$24671 ( \33394_33694 , \33149_33449 , \33318_33618 );
and \U$24672 ( \33395_33695 , \33154_33454 , \33318_33618 );
or \U$24673 ( \33396_33696 , \33393_33693 , \33394_33694 , \33395_33695 );
buf \U$24674 ( \33397_33697 , \33396_33696 );
and \U$24675 ( \33398_33698 , \16405_15940 , \25561_25860_nG9bc9 );
and \U$24676 ( \33399_33699 , \15638_15937 , \26585_26887_nG9bc6 );
or \U$24677 ( \33400_33700 , \33398_33698 , \33399_33699 );
xor \U$24678 ( \33401_33701 , \15637_15936 , \33400_33700 );
buf \U$24679 ( \33402_33702 , \33401_33701 );
buf \U$24681 ( \33403_33703 , \33402_33702 );
and \U$24682 ( \33404_33704 , \13431_13370 , \28877_29179_nG9bbd );
and \U$24683 ( \33405_33705 , \13068_13367 , \30064_30366_nG9bba );
or \U$24684 ( \33406_33706 , \33404_33704 , \33405_33705 );
xor \U$24685 ( \33407_33707 , \13067_13366 , \33406_33706 );
buf \U$24686 ( \33408_33708 , \33407_33707 );
buf \U$24688 ( \33409_33709 , \33408_33708 );
xor \U$24689 ( \33410_33710 , \33403_33703 , \33409_33709 );
and \U$24690 ( \33411_33711 , \12183_12157 , \30638_30940_nG9bb7 );
and \U$24691 ( \33412_33712 , \11855_12154 , \31877_32179_nG9bb4 );
or \U$24692 ( \33413_33713 , \33411_33711 , \33412_33712 );
xor \U$24693 ( \33414_33714 , \11854_12153 , \33413_33713 );
buf \U$24694 ( \33415_33715 , \33414_33714 );
buf \U$24696 ( \33416_33716 , \33415_33715 );
xor \U$24697 ( \33417_33717 , \33410_33710 , \33416_33716 );
buf \U$24698 ( \33418_33718 , \33417_33717 );
xor \U$24699 ( \33419_33719 , \33397_33697 , \33418_33718 );
and \U$24700 ( \33420_33720 , \33011_33311 , \33028_33328 );
and \U$24701 ( \33421_33721 , \33011_33311 , \33035_33335 );
and \U$24702 ( \33422_33722 , \33028_33328 , \33035_33335 );
or \U$24703 ( \33423_33723 , \33420_33720 , \33421_33721 , \33422_33722 );
buf \U$24704 ( \33424_33724 , \33423_33723 );
and \U$24705 ( \33425_33725 , \33013_33313 , \33019_33319 );
and \U$24706 ( \33426_33726 , \33013_33313 , \33026_33326 );
and \U$24707 ( \33427_33727 , \33019_33319 , \33026_33326 );
or \U$24708 ( \33428_33728 , \33425_33725 , \33426_33726 , \33427_33727 );
buf \U$24709 ( \33429_33729 , \33428_33728 );
and \U$24711 ( \33430_33730 , \32617_32916 , \10981_11283_nG9c08 );
or \U$24712 ( \33431_33731 , 1'b0 , \33430_33730 );
xor \U$24713 ( \33432_33732 , 1'b0 , \33431_33731 );
buf \U$24714 ( \33433_33733 , \33432_33732 );
buf \U$24716 ( \33434_33734 , \33433_33733 );
and \U$24717 ( \33435_33735 , \31989_31636 , \11299_11598_nG9c05 );
and \U$24718 ( \33436_33736 , \31334_31633 , \12168_12470_nG9c02 );
or \U$24719 ( \33437_33737 , \33435_33735 , \33436_33736 );
xor \U$24720 ( \33438_33738 , \31333_31632 , \33437_33737 );
buf \U$24721 ( \33439_33739 , \33438_33738 );
buf \U$24723 ( \33440_33740 , \33439_33739 );
xor \U$24724 ( \33441_33741 , \33434_33734 , \33440_33740 );
buf \U$24725 ( \33442_33742 , \33441_33741 );
and \U$24726 ( \33443_33743 , \30670_29853 , \12502_12801_nG9bff );
and \U$24727 ( \33444_33744 , \29551_29850 , \13403_13705_nG9bfc );
or \U$24728 ( \33445_33745 , \33443_33743 , \33444_33744 );
xor \U$24729 ( \33446_33746 , \29550_29849 , \33445_33745 );
buf \U$24730 ( \33447_33747 , \33446_33746 );
buf \U$24732 ( \33448_33748 , \33447_33747 );
xor \U$24733 ( \33449_33749 , \33442_33742 , \33448_33748 );
buf \U$24734 ( \33450_33750 , \33449_33749 );
xor \U$24735 ( \33451_33751 , \33429_33729 , \33450_33750 );
and \U$24736 ( \33452_33752 , \25044_24792 , \16378_16680_nG9bed );
and \U$24737 ( \33453_33753 , \24490_24789 , \17363_17665_nG9bea );
or \U$24738 ( \33454_33754 , \33452_33752 , \33453_33753 );
xor \U$24739 ( \33455_33755 , \24489_24788 , \33454_33754 );
buf \U$24740 ( \33456_33756 , \33455_33755 );
buf \U$24742 ( \33457_33757 , \33456_33756 );
xor \U$24743 ( \33458_33758 , \33451_33751 , \33457_33757 );
buf \U$24744 ( \33459_33759 , \33458_33758 );
xor \U$24745 ( \33460_33760 , \33424_33724 , \33459_33759 );
and \U$24746 ( \33461_33761 , \17437_17297 , \23927_24226_nG9bcf );
and \U$24747 ( \33462_33762 , \16995_17294 , \24996_25298_nG9bcc );
or \U$24748 ( \33463_33763 , \33461_33761 , \33462_33762 );
xor \U$24749 ( \33464_33764 , \16994_17293 , \33463_33763 );
buf \U$24750 ( \33465_33765 , \33464_33764 );
buf \U$24752 ( \33466_33766 , \33465_33765 );
xor \U$24753 ( \33467_33767 , \33460_33760 , \33466_33766 );
buf \U$24754 ( \33468_33768 , \33467_33767 );
and \U$24755 ( \33469_33769 , \33042_33342 , \33062_33362 );
and \U$24756 ( \33470_33770 , \33042_33342 , \33069_33369 );
and \U$24757 ( \33471_33771 , \33062_33362 , \33069_33369 );
or \U$24758 ( \33472_33772 , \33469_33769 , \33470_33770 , \33471_33771 );
buf \U$24759 ( \33473_33773 , \33472_33772 );
and \U$24760 ( \33474_33774 , \33047_33347 , \33053_33353 );
and \U$24761 ( \33475_33775 , \33047_33347 , \33060_33360 );
and \U$24762 ( \33476_33776 , \33053_33353 , \33060_33360 );
or \U$24763 ( \33477_33777 , \33474_33774 , \33475_33775 , \33476_33776 );
buf \U$24764 ( \33478_33778 , \33477_33777 );
and \U$24765 ( \33479_33779 , \28946_28118 , \13771_14070_nG9bf9 );
and \U$24766 ( \33480_33780 , \27816_28115 , \14682_14984_nG9bf6 );
or \U$24767 ( \33481_33781 , \33479_33779 , \33480_33780 );
xor \U$24768 ( \33482_33782 , \27815_28114 , \33481_33781 );
buf \U$24769 ( \33483_33783 , \33482_33782 );
buf \U$24771 ( \33484_33784 , \33483_33783 );
xor \U$24772 ( \33485_33785 , \33478_33778 , \33484_33784 );
and \U$24773 ( \33486_33786 , \27141_26431 , \15074_15373_nG9bf3 );
and \U$24774 ( \33487_33787 , \26129_26428 , \16013_16315_nG9bf0 );
or \U$24775 ( \33488_33788 , \33486_33786 , \33487_33787 );
xor \U$24776 ( \33489_33789 , \26128_26427 , \33488_33788 );
buf \U$24777 ( \33490_33790 , \33489_33789 );
buf \U$24779 ( \33491_33791 , \33490_33790 );
xor \U$24780 ( \33492_33792 , \33485_33785 , \33491_33791 );
buf \U$24781 ( \33493_33793 , \33492_33792 );
xor \U$24782 ( \33494_33794 , \33473_33773 , \33493_33793 );
and \U$24783 ( \33495_33795 , \18908_18702 , \22330_22629_nG9bd5 );
and \U$24784 ( \33496_33796 , \18400_18699 , \23394_23696_nG9bd2 );
or \U$24785 ( \33497_33797 , \33495_33795 , \33496_33796 );
xor \U$24786 ( \33498_33798 , \18399_18698 , \33497_33797 );
buf \U$24787 ( \33499_33799 , \33498_33798 );
buf \U$24789 ( \33500_33800 , \33499_33799 );
xor \U$24790 ( \33501_33801 , \33494_33794 , \33500_33800 );
buf \U$24791 ( \33502_33802 , \33501_33801 );
xor \U$24792 ( \33503_33803 , \33468_33768 , \33502_33802 );
and \U$24793 ( \33504_33804 , \10996_10421 , \32589_32888_nG9bb1 );
and \U$24794 ( \33505_33805 , \10119_10418 , \32881_33181_nG9bae );
or \U$24795 ( \33506_33806 , \33504_33804 , \33505_33805 );
xor \U$24796 ( \33507_33807 , \10118_10417 , \33506_33806 );
buf \U$24797 ( \33508_33808 , \33507_33807 );
buf \U$24799 ( \33509_33809 , \33508_33808 );
xor \U$24800 ( \33510_33810 , \33503_33803 , \33509_33809 );
buf \U$24801 ( \33511_33811 , \33510_33810 );
xor \U$24802 ( \33512_33812 , \33419_33719 , \33511_33811 );
buf \U$24803 ( \33513_33813 , \33512_33812 );
xor \U$24804 ( \33514_33814 , \33392_33692 , \33513_33813 );
and \U$24805 ( \33515_33815 , \33106_33406 , \33112_33412 );
and \U$24806 ( \33516_33816 , \33106_33406 , \33119_33419 );
and \U$24807 ( \33517_33817 , \33112_33412 , \33119_33419 );
or \U$24808 ( \33518_33818 , \33515_33815 , \33516_33816 , \33517_33817 );
buf \U$24809 ( \33519_33819 , \33518_33818 );
and \U$24810 ( \33520_33820 , \33071_33371 , \33077_33377 );
and \U$24811 ( \33521_33821 , \33071_33371 , \33084_33384 );
and \U$24812 ( \33522_33822 , \33077_33377 , \33084_33384 );
or \U$24813 ( \33523_33823 , \33520_33820 , \33521_33821 , \33522_33822 );
buf \U$24814 ( \33524_33824 , \33523_33823 );
and \U$24815 ( \33525_33825 , \23495_23201 , \17808_18107_nG9be7 );
and \U$24816 ( \33526_33826 , \22899_23198 , \18789_19091_nG9be4 );
or \U$24817 ( \33527_33827 , \33525_33825 , \33526_33826 );
xor \U$24818 ( \33528_33828 , \22898_23197 , \33527_33827 );
buf \U$24819 ( \33529_33829 , \33528_33828 );
buf \U$24821 ( \33530_33830 , \33529_33829 );
and \U$24822 ( \33531_33831 , \21908_21658 , \19287_19586_nG9be1 );
and \U$24823 ( \33532_33832 , \21356_21655 , \20306_20608_nG9bde );
or \U$24824 ( \33533_33833 , \33531_33831 , \33532_33832 );
xor \U$24825 ( \33534_33834 , \21355_21654 , \33533_33833 );
buf \U$24826 ( \33535_33835 , \33534_33834 );
buf \U$24828 ( \33536_33836 , \33535_33835 );
xor \U$24829 ( \33537_33837 , \33530_33830 , \33536_33836 );
and \U$24830 ( \33538_33838 , \20353_20155 , \20787_21086_nG9bdb );
and \U$24831 ( \33539_33839 , \19853_20152 , \21827_22129_nG9bd8 );
or \U$24832 ( \33540_33840 , \33538_33838 , \33539_33839 );
xor \U$24833 ( \33541_33841 , \19852_20151 , \33540_33840 );
buf \U$24834 ( \33542_33842 , \33541_33841 );
buf \U$24836 ( \33543_33843 , \33542_33842 );
xor \U$24837 ( \33544_33844 , \33537_33837 , \33543_33843 );
buf \U$24838 ( \33545_33845 , \33544_33844 );
xor \U$24839 ( \33546_33846 , \33524_33824 , \33545_33845 );
and \U$24840 ( \33547_33847 , \14710_14631 , \27114_27416_nG9bc3 );
and \U$24841 ( \33548_33848 , \14329_14628 , \28300_28602_nG9bc0 );
or \U$24842 ( \33549_33849 , \33547_33847 , \33548_33848 );
xor \U$24843 ( \33550_33850 , \14328_14627 , \33549_33849 );
buf \U$24844 ( \33551_33851 , \33550_33850 );
buf \U$24846 ( \33552_33852 , \33551_33851 );
xor \U$24847 ( \33553_33853 , \33546_33846 , \33552_33852 );
buf \U$24848 ( \33554_33854 , \33553_33853 );
xor \U$24849 ( \33555_33855 , \33519_33819 , \33554_33854 );
and \U$24850 ( \33556_33856 , \33344_33644 , \33350_33650 );
and \U$24851 ( \33557_33857 , \33344_33644 , \33357_33657 );
and \U$24852 ( \33558_33858 , \33350_33650 , \33357_33657 );
or \U$24853 ( \33559_33859 , \33556_33856 , \33557_33857 , \33558_33858 );
buf \U$24854 ( \33560_33860 , \33559_33859 );
xor \U$24855 ( \33561_33861 , \33555_33855 , \33560_33860 );
buf \U$24856 ( \33562_33862 , \33561_33861 );
xor \U$24857 ( \33563_33863 , \33514_33814 , \33562_33862 );
buf \U$24858 ( \33564_33864 , \33563_33863 );
and \U$24859 ( \33565_33865 , \33328_33628 , \33361_33661 );
and \U$24860 ( \33566_33866 , \33328_33628 , \33367_33667 );
and \U$24861 ( \33567_33867 , \33361_33661 , \33367_33667 );
or \U$24862 ( \33568_33868 , \33565_33865 , \33566_33866 , \33567_33867 );
buf \U$24863 ( \33569_33869 , \33568_33868 );
xor \U$24864 ( \33570_33870 , \33564_33864 , \33569_33869 );
and \U$24865 ( \33571_33871 , \33037_33337 , \33086_33386 );
and \U$24866 ( \33572_33872 , \33037_33337 , \33092_33392 );
and \U$24867 ( \33573_33873 , \33086_33386 , \33092_33392 );
or \U$24868 ( \33574_33874 , \33571_33871 , \33572_33872 , \33573_33873 );
buf \U$24869 ( \33575_33875 , \33574_33874 );
and \U$24870 ( \33576_33876 , \33134_33434 , \33140_33440 );
and \U$24871 ( \33577_33877 , \33134_33434 , \33147_33447 );
and \U$24872 ( \33578_33878 , \33140_33440 , \33147_33447 );
or \U$24873 ( \33579_33879 , \33576_33876 , \33577_33877 , \33578_33878 );
buf \U$24874 ( \33580_33880 , \33579_33879 );
xor \U$24875 ( \33581_33881 , \33575_33875 , \33580_33880 );
and \U$24876 ( \33582_33882 , \10411_10707 , \33313_33613_nG9bab );
and \U$24877 ( \33583_33883 , \33215_33515 , \33219_33519 );
and \U$24878 ( \33584_33884 , \33219_33519 , \33301_33601 );
and \U$24879 ( \33585_33885 , \33215_33515 , \33301_33601 );
or \U$24880 ( \33586_33886 , \33583_33883 , \33584_33884 , \33585_33885 );
and \U$24881 ( \33587_33887 , \33168_33468 , \33172_33472 );
and \U$24882 ( \33588_33888 , \33172_33472 , \33177_33477 );
and \U$24883 ( \33589_33889 , \33168_33468 , \33177_33477 );
or \U$24884 ( \33590_33890 , \33587_33887 , \33588_33888 , \33589_33889 );
and \U$24885 ( \33591_33891 , \33187_33487 , \33191_33491 );
and \U$24886 ( \33592_33892 , \33191_33491 , \33196_33496 );
and \U$24887 ( \33593_33893 , \33187_33487 , \33196_33496 );
or \U$24888 ( \33594_33894 , \33591_33891 , \33592_33892 , \33593_33893 );
and \U$24889 ( \33595_33895 , \33202_33502 , \10678_10980 );
and \U$24890 ( \33596_33896 , \10678_10980 , \33207_33507 );
and \U$24891 ( \33597_33897 , \33202_33502 , \33207_33507 );
or \U$24892 ( \33598_33898 , \33595_33895 , \33596_33896 , \33597_33897 );
xor \U$24893 ( \33599_33899 , \33594_33894 , \33598_33898 );
and \U$24894 ( \33600_33900 , \33260_33560 , \33264_33564 );
and \U$24895 ( \33601_33901 , \33264_33564 , \33269_33569 );
and \U$24896 ( \33602_33902 , \33260_33560 , \33269_33569 );
or \U$24897 ( \33603_33903 , \33600_33900 , \33601_33901 , \33602_33902 );
and \U$24898 ( \33604_33904 , \33274_33574 , \33278_33578 );
and \U$24899 ( \33605_33905 , \33278_33578 , \33283_33583 );
and \U$24900 ( \33606_33906 , \33274_33574 , \33283_33583 );
or \U$24901 ( \33607_33907 , \33604_33904 , \33605_33905 , \33606_33906 );
xor \U$24902 ( \33608_33908 , \33603_33903 , \33607_33907 );
and \U$24903 ( \33609_33909 , \33289_33589 , \33293_33593 );
and \U$24904 ( \33610_33910 , \33293_33593 , \33298_33598 );
and \U$24905 ( \33611_33911 , \33289_33589 , \33298_33598 );
or \U$24906 ( \33612_33912 , \33609_33909 , \33610_33910 , \33611_33911 );
xor \U$24907 ( \33613_33913 , \33608_33908 , \33612_33912 );
xor \U$24908 ( \33614_33914 , \33599_33899 , \33613_33913 );
xor \U$24909 ( \33615_33915 , \33590_33890 , \33614_33914 );
and \U$24910 ( \33616_33916 , \33228_33528 , \33239_33539 );
and \U$24911 ( \33617_33917 , \33239_33539 , \33254_33554 );
and \U$24912 ( \33618_33918 , \33228_33528 , \33254_33554 );
or \U$24913 ( \33619_33919 , \33616_33916 , \33617_33917 , \33618_33918 );
and \U$24914 ( \33620_33920 , \33270_33570 , \33284_33584 );
and \U$24915 ( \33621_33921 , \33284_33584 , \33299_33599 );
and \U$24916 ( \33622_33922 , \33270_33570 , \33299_33599 );
or \U$24917 ( \33623_33923 , \33620_33920 , \33621_33921 , \33622_33922 );
xor \U$24918 ( \33624_33924 , \33619_33919 , \33623_33923 );
and \U$24919 ( \33625_33925 , \33232_33532 , \33236_33536 );
and \U$24920 ( \33626_33926 , \33236_33536 , \33238_33538 );
and \U$24921 ( \33627_33927 , \33232_33532 , \33238_33538 );
or \U$24922 ( \33628_33928 , \33625_33925 , \33626_33926 , \33627_33927 );
not \U$24923 ( \33629_33929 , \10678_10980 );
buf \U$24924 ( \33630_33930 , \33629_33929 );
xor \U$24925 ( \33631_33931 , \33628_33928 , \33630_33930 );
and \U$24926 ( \33632_33932 , \32495_32794 , \11275_11574 );
not \U$24927 ( \33633_33933 , \33632_33932 );
xnor \U$24928 ( \33634_33934 , \33633_33933 , \11281_11580 );
not \U$24929 ( \33635_33935 , \33634_33934 );
xor \U$24930 ( \33636_33936 , \33631_33931 , \33635_33935 );
xor \U$24931 ( \33637_33937 , \33624_33924 , \33636_33936 );
xor \U$24932 ( \33638_33938 , \33615_33915 , \33637_33937 );
xor \U$24933 ( \33639_33939 , \33586_33886 , \33638_33938 );
and \U$24934 ( \33640_33940 , \33224_33524 , \33255_33555 );
and \U$24935 ( \33641_33941 , \33255_33555 , \33300_33600 );
and \U$24936 ( \33642_33942 , \33224_33524 , \33300_33600 );
or \U$24937 ( \33643_33943 , \33640_33940 , \33641_33941 , \33642_33942 );
and \U$24938 ( \33644_33944 , \33164_33464 , \33178_33478 );
and \U$24939 ( \33645_33945 , \33178_33478 , \33209_33509 );
and \U$24940 ( \33646_33946 , \33164_33464 , \33209_33509 );
or \U$24941 ( \33647_33947 , \33644_33944 , \33645_33945 , \33646_33946 );
xor \U$24942 ( \33648_33948 , \33643_33943 , \33647_33947 );
and \U$24943 ( \33649_33949 , \33183_33483 , \33197_33497 );
and \U$24944 ( \33650_33950 , \33197_33497 , \33208_33508 );
and \U$24945 ( \33651_33951 , \33183_33483 , \33208_33508 );
or \U$24946 ( \33652_33952 , \33649_33949 , \33650_33950 , \33651_33951 );
and \U$24947 ( \33653_33953 , \30500_30802 , \12491_12790 );
and \U$24948 ( \33654_33954 , \31752_32054 , \12159_12461 );
nor \U$24949 ( \33655_33955 , \33653_33953 , \33654_33954 );
xnor \U$24950 ( \33656_33956 , \33655_33955 , \12481_12780 );
and \U$24951 ( \33657_33957 , \27011_27313 , \15037_15336 );
and \U$24952 ( \33658_33958 , \28232_28534 , \14661_14963 );
nor \U$24953 ( \33659_33959 , \33657_33957 , \33658_33958 );
xnor \U$24954 ( \33660_33960 , \33659_33959 , \15043_15342 );
xor \U$24955 ( \33661_33961 , \33656_33956 , \33660_33960 );
and \U$24956 ( \33662_33962 , \10968_11270 , \32503_32802 );
xor \U$24957 ( \33663_33963 , \33661_33961 , \33662_33962 );
and \U$24958 ( \33664_33964 , \23900_24199 , \17791_18090 );
and \U$24959 ( \33665_33965 , \24970_25272 , \17353_17655 );
nor \U$24960 ( \33666_33966 , \33664_33964 , \33665_33965 );
xnor \U$24961 ( \33667_33967 , \33666_33966 , \17747_18046 );
and \U$24962 ( \33668_33968 , \15022_15321 , \27095_27397 );
and \U$24963 ( \33669_33969 , \15965_16267 , \26505_26807 );
nor \U$24964 ( \33670_33970 , \33668_33968 , \33669_33969 );
xnor \U$24965 ( \33671_33971 , \33670_33970 , \26993_27295 );
xor \U$24966 ( \33672_33972 , \33667_33967 , \33671_33971 );
and \U$24967 ( \33673_33973 , \13725_14024 , \28768_29070 );
and \U$24968 ( \33674_33974 , \14648_14950 , \28224_28526 );
nor \U$24969 ( \33675_33975 , \33673_33973 , \33674_33974 );
xnor \U$24970 ( \33676_33976 , \33675_33975 , \28774_29076 );
xor \U$24971 ( \33677_33977 , \33672_33972 , \33676_33976 );
xor \U$24972 ( \33678_33978 , \33663_33963 , \33677_33977 );
and \U$24973 ( \33679_33979 , \28782_29084 , \13755_14054 );
and \U$24974 ( \33680_33980 , \29966_30268 , \13390_13692 );
nor \U$24975 ( \33681_33981 , \33679_33979 , \33680_33980 );
xnor \U$24976 ( \33682_33982 , \33681_33981 , \13736_14035 );
and \U$24977 ( \33683_33983 , \17736_18035 , \23839_24138 );
and \U$24978 ( \33684_33984 , \18730_19032 , \23328_23630 );
nor \U$24979 ( \33685_33985 , \33683_33983 , \33684_33984 );
xnor \U$24980 ( \33686_33986 , \33685_33985 , \23845_24144 );
xor \U$24981 ( \33687_33987 , \33682_33982 , \33686_33986 );
and \U$24982 ( \33688_33988 , \16353_16655 , \25527_25826 );
and \U$24983 ( \33689_33989 , \17325_17627 , \24962_25264 );
nor \U$24984 ( \33690_33990 , \33688_33988 , \33689_33989 );
xnor \U$24985 ( \33691_33991 , \33690_33990 , \25474_25773 );
xor \U$24986 ( \33692_33992 , \33687_33987 , \33691_33991 );
xor \U$24987 ( \33693_33993 , \33678_33978 , \33692_33992 );
xor \U$24988 ( \33694_33994 , \33652_33952 , \33693_33993 );
and \U$24989 ( \33695_33995 , \33244_33544 , \33248_33548 );
and \U$24990 ( \33696_33996 , \33248_33548 , \33253_33553 );
and \U$24991 ( \33697_33997 , \33244_33544 , \33253_33553 );
or \U$24992 ( \33698_33998 , \33695_33995 , \33696_33996 , \33697_33997 );
and \U$24993 ( \33699_33999 , \22257_22556 , \19235_19534 );
and \U$24994 ( \33700_34000 , \23315_23617 , \18743_19045 );
nor \U$24995 ( \33701_34001 , \33699_33999 , \33700_34000 );
xnor \U$24996 ( \33702_34002 , \33701_34001 , \19241_19540 );
and \U$24997 ( \33703_34003 , \12470_12769 , \30521_30823 );
and \U$24998 ( \33704_34004 , \13377_13679 , \29944_30246 );
nor \U$24999 ( \33705_34005 , \33703_34003 , \33704_34004 );
xnor \U$25000 ( \33706_34006 , \33705_34005 , \30511_30813 );
xor \U$25001 ( \33707_34007 , \33702_34002 , \33706_34006 );
and \U$25002 ( \33708_34008 , \11287_11586 , \32555_32854 );
and \U$25003 ( \33709_34009 , \12146_12448 , \31765_32067 );
nor \U$25004 ( \33710_34010 , \33708_34008 , \33709_34009 );
xnor \U$25005 ( \33711_34011 , \33710_34010 , \32506_32805 );
xor \U$25006 ( \33712_34012 , \33707_34007 , \33711_34011 );
xor \U$25007 ( \33713_34013 , \33698_33998 , \33712_34012 );
and \U$25008 ( \33714_34014 , \25516_25815 , \16333_16635 );
and \U$25009 ( \33715_34015 , \26527_26829 , \15999_16301 );
nor \U$25010 ( \33716_34016 , \33714_34014 , \33715_34015 );
xnor \U$25011 ( \33717_34017 , \33716_34016 , \16323_16625 );
and \U$25012 ( \33718_34018 , \20734_21033 , \20706_21005 );
and \U$25013 ( \33719_34019 , \21788_22090 , \20255_20557 );
nor \U$25014 ( \33720_34020 , \33718_34018 , \33719_34019 );
xnor \U$25015 ( \33721_34021 , \33720_34020 , \20712_21011 );
xor \U$25016 ( \33722_34022 , \33717_34017 , \33721_34021 );
and \U$25017 ( \33723_34023 , \19259_19558 , \22243_22542 );
and \U$25018 ( \33724_34024 , \20242_20544 , \21801_22103 );
nor \U$25019 ( \33725_34025 , \33723_34023 , \33724_34024 );
xnor \U$25020 ( \33726_34026 , \33725_34025 , \22249_22548 );
xor \U$25021 ( \33727_34027 , \33722_34022 , \33726_34026 );
xor \U$25022 ( \33728_34028 , \33713_34013 , \33727_34027 );
xor \U$25023 ( \33729_34029 , \33694_33994 , \33728_34028 );
xor \U$25024 ( \33730_34030 , \33648_33948 , \33729_34029 );
xor \U$25025 ( \33731_34031 , \33639_33939 , \33730_34030 );
and \U$25026 ( \33732_34032 , \33160_33460 , \33210_33510 );
and \U$25027 ( \33733_34033 , \33210_33510 , \33302_33602 );
and \U$25028 ( \33734_34034 , \33160_33460 , \33302_33602 );
or \U$25029 ( \33735_34035 , \33732_34032 , \33733_34033 , \33734_34034 );
xor \U$25030 ( \33736_34036 , \33731_34031 , \33735_34035 );
and \U$25031 ( \33737_34037 , \33303_33603 , \33307_33607 );
and \U$25032 ( \33738_34038 , \33308_33608 , \33311_33611 );
or \U$25033 ( \33739_34039 , \33737_34037 , \33738_34038 );
xor \U$25034 ( \33740_34040 , \33736_34036 , \33739_34039 );
buf g9ba8_GF_PartitionCandidate( \33741_34041_nG9ba8 , \33740_34040 );
and \U$25035 ( \33742_34042 , \10402_10704 , \33741_34041_nG9ba8 );
or \U$25036 ( \33743_34043 , \33582_33882 , \33742_34042 );
xor \U$25037 ( \33744_34044 , \10399_10703 , \33743_34043 );
buf \U$25038 ( \33745_34045 , \33744_34044 );
buf \U$25040 ( \33746_34046 , \33745_34045 );
xor \U$25041 ( \33747_34047 , \33581_33881 , \33746_34046 );
buf \U$25042 ( \33748_34048 , \33747_34047 );
and \U$25043 ( \33749_34049 , \33094_33394 , \33099_33399 );
and \U$25044 ( \33750_34050 , \33094_33394 , \33121_33421 );
and \U$25045 ( \33751_34051 , \33099_33399 , \33121_33421 );
or \U$25046 ( \33752_34052 , \33749_34049 , \33750_34050 , \33751_34051 );
buf \U$25047 ( \33753_34053 , \33752_34052 );
xor \U$25048 ( \33754_34054 , \33748_34048 , \33753_34053 );
and \U$25049 ( \33755_34055 , \33333_33633 , \33338_33638 );
and \U$25050 ( \33756_34056 , \33333_33633 , \33359_33659 );
and \U$25051 ( \33757_34057 , \33338_33638 , \33359_33659 );
or \U$25052 ( \33758_34058 , \33755_34055 , \33756_34056 , \33757_34057 );
buf \U$25053 ( \33759_34059 , \33758_34058 );
xor \U$25054 ( \33760_34060 , \33754_34054 , \33759_34059 );
buf \U$25055 ( \33761_34061 , \33760_34060 );
xor \U$25056 ( \33762_34062 , \33570_33870 , \33761_34061 );
and \U$25057 ( \33763_34063 , \33382_33682 , \33762_34062 );
and \U$25058 ( \33764_34064 , \33386_33686 , \33762_34062 );
or \U$25059 ( \33765_34065 , \33387_33687 , \33763_34063 , \33764_34064 );
and \U$25060 ( \33766_34066 , \33378_33678 , \33380_33680 );
or \U$25063 ( \33767_34067 , \33766_34066 , 1'b0 , 1'b0 );
xor \U$25064 ( \33768_34068 , \33765_34065 , \33767_34067 );
xor \U$25068 ( \33769_34069 , \33768_34068 , 1'b0 );
xor \U$25075 ( \33770_34070 , \33769_34069 , 1'b0 );
and \U$25076 ( \33771_34071 , \33564_33864 , \33569_33869 );
and \U$25077 ( \33772_34072 , \33564_33864 , \33761_34061 );
and \U$25078 ( \33773_34073 , \33569_33869 , \33761_34061 );
or \U$25079 ( \33774_34074 , \33771_34071 , \33772_34072 , \33773_34073 );
xor \U$25080 ( \33775_34075 , \33770_34070 , \33774_34074 );
and \U$25081 ( \33776_34076 , \33392_33692 , \33513_33813 );
and \U$25082 ( \33777_34077 , \33392_33692 , \33562_33862 );
and \U$25083 ( \33778_34078 , \33513_33813 , \33562_33862 );
or \U$25084 ( \33779_34079 , \33776_34076 , \33777_34077 , \33778_34078 );
buf \U$25085 ( \33780_34080 , \33779_34079 );
and \U$25086 ( \33781_34081 , \33478_33778 , \33484_33784 );
and \U$25087 ( \33782_34082 , \33478_33778 , \33491_33791 );
and \U$25088 ( \33783_34083 , \33484_33784 , \33491_33791 );
or \U$25089 ( \33784_34084 , \33781_34081 , \33782_34082 , \33783_34083 );
buf \U$25090 ( \33785_34085 , \33784_34084 );
and \U$25092 ( \33786_34086 , \32617_32916 , \11299_11598_nG9c05 );
or \U$25093 ( \33787_34087 , 1'b0 , \33786_34086 );
xor \U$25094 ( \33788_34088 , 1'b0 , \33787_34087 );
buf \U$25095 ( \33789_34089 , \33788_34088 );
buf \U$25097 ( \33790_34090 , \33789_34089 );
and \U$25098 ( \33791_34091 , \31989_31636 , \12168_12470_nG9c02 );
and \U$25099 ( \33792_34092 , \31334_31633 , \12502_12801_nG9bff );
or \U$25100 ( \33793_34093 , \33791_34091 , \33792_34092 );
xor \U$25101 ( \33794_34094 , \31333_31632 , \33793_34093 );
buf \U$25102 ( \33795_34095 , \33794_34094 );
buf \U$25104 ( \33796_34096 , \33795_34095 );
xor \U$25105 ( \33797_34097 , \33790_34090 , \33796_34096 );
buf \U$25106 ( \33798_34098 , \33797_34097 );
and \U$25107 ( \33799_34099 , \33434_33734 , \33440_33740 );
buf \U$25108 ( \33800_34100 , \33799_34099 );
xor \U$25109 ( \33801_34101 , \33798_34098 , \33800_34100 );
and \U$25110 ( \33802_34102 , \30670_29853 , \13403_13705_nG9bfc );
and \U$25111 ( \33803_34103 , \29551_29850 , \13771_14070_nG9bf9 );
or \U$25112 ( \33804_34104 , \33802_34102 , \33803_34103 );
xor \U$25113 ( \33805_34105 , \29550_29849 , \33804_34104 );
buf \U$25114 ( \33806_34106 , \33805_34105 );
buf \U$25116 ( \33807_34107 , \33806_34106 );
xor \U$25117 ( \33808_34108 , \33801_34101 , \33807_34107 );
buf \U$25118 ( \33809_34109 , \33808_34108 );
xor \U$25119 ( \33810_34110 , \33785_34085 , \33809_34109 );
and \U$25120 ( \33811_34111 , \25044_24792 , \17363_17665_nG9bea );
and \U$25121 ( \33812_34112 , \24490_24789 , \17808_18107_nG9be7 );
or \U$25122 ( \33813_34113 , \33811_34111 , \33812_34112 );
xor \U$25123 ( \33814_34114 , \24489_24788 , \33813_34113 );
buf \U$25124 ( \33815_34115 , \33814_34114 );
buf \U$25126 ( \33816_34116 , \33815_34115 );
xor \U$25127 ( \33817_34117 , \33810_34110 , \33816_34116 );
buf \U$25128 ( \33818_34118 , \33817_34117 );
and \U$25129 ( \33819_34119 , \33530_33830 , \33536_33836 );
and \U$25130 ( \33820_34120 , \33530_33830 , \33543_33843 );
and \U$25131 ( \33821_34121 , \33536_33836 , \33543_33843 );
or \U$25132 ( \33822_34122 , \33819_34119 , \33820_34120 , \33821_34121 );
buf \U$25133 ( \33823_34123 , \33822_34122 );
xor \U$25134 ( \33824_34124 , \33818_34118 , \33823_34123 );
and \U$25135 ( \33825_34125 , \16405_15940 , \26585_26887_nG9bc6 );
and \U$25136 ( \33826_34126 , \15638_15937 , \27114_27416_nG9bc3 );
or \U$25137 ( \33827_34127 , \33825_34125 , \33826_34126 );
xor \U$25138 ( \33828_34128 , \15637_15936 , \33827_34127 );
buf \U$25139 ( \33829_34129 , \33828_34128 );
buf \U$25141 ( \33830_34130 , \33829_34129 );
xor \U$25142 ( \33831_34131 , \33824_34124 , \33830_34130 );
buf \U$25143 ( \33832_34132 , \33831_34131 );
and \U$25144 ( \33833_34133 , \33524_33824 , \33545_33845 );
and \U$25145 ( \33834_34134 , \33524_33824 , \33552_33852 );
and \U$25146 ( \33835_34135 , \33545_33845 , \33552_33852 );
or \U$25147 ( \33836_34136 , \33833_34133 , \33834_34134 , \33835_34135 );
buf \U$25148 ( \33837_34137 , \33836_34136 );
xor \U$25149 ( \33838_34138 , \33832_34132 , \33837_34137 );
and \U$25150 ( \33839_34139 , \10411_10707 , \33741_34041_nG9ba8 );
and \U$25151 ( \33840_34140 , \33586_33886 , \33638_33938 );
and \U$25152 ( \33841_34141 , \33638_33938 , \33730_34030 );
and \U$25153 ( \33842_34142 , \33586_33886 , \33730_34030 );
or \U$25154 ( \33843_34143 , \33840_34140 , \33841_34141 , \33842_34142 );
and \U$25155 ( \33844_34144 , \33643_33943 , \33647_33947 );
and \U$25156 ( \33845_34145 , \33647_33947 , \33729_34029 );
and \U$25157 ( \33846_34146 , \33643_33943 , \33729_34029 );
or \U$25158 ( \33847_34147 , \33844_34144 , \33845_34145 , \33846_34146 );
and \U$25159 ( \33848_34148 , \33594_33894 , \33598_33898 );
and \U$25160 ( \33849_34149 , \33598_33898 , \33613_33913 );
and \U$25161 ( \33850_34150 , \33594_33894 , \33613_33913 );
or \U$25162 ( \33851_34151 , \33848_34148 , \33849_34149 , \33850_34150 );
and \U$25163 ( \33852_34152 , \33619_33919 , \33623_33923 );
and \U$25164 ( \33853_34153 , \33623_33923 , \33636_33936 );
and \U$25165 ( \33854_34154 , \33619_33919 , \33636_33936 );
or \U$25166 ( \33855_34155 , \33852_34152 , \33853_34153 , \33854_34154 );
xor \U$25167 ( \33856_34156 , \33851_34151 , \33855_34155 );
and \U$25168 ( \33857_34157 , \33663_33963 , \33677_33977 );
and \U$25169 ( \33858_34158 , \33677_33977 , \33692_33992 );
and \U$25170 ( \33859_34159 , \33663_33963 , \33692_33992 );
or \U$25171 ( \33860_34160 , \33857_34157 , \33858_34158 , \33859_34159 );
and \U$25172 ( \33861_34161 , \33698_33998 , \33712_34012 );
and \U$25173 ( \33862_34162 , \33712_34012 , \33727_34027 );
and \U$25174 ( \33863_34163 , \33698_33998 , \33727_34027 );
or \U$25175 ( \33864_34164 , \33861_34161 , \33862_34162 , \33863_34163 );
xor \U$25176 ( \33865_34165 , \33860_34160 , \33864_34164 );
and \U$25177 ( \33866_34166 , \33717_34017 , \33721_34021 );
and \U$25178 ( \33867_34167 , \33721_34021 , \33726_34026 );
and \U$25179 ( \33868_34168 , \33717_34017 , \33726_34026 );
or \U$25180 ( \33869_34169 , \33866_34166 , \33867_34167 , \33868_34168 );
and \U$25181 ( \33870_34170 , \33667_33967 , \33671_33971 );
and \U$25182 ( \33871_34171 , \33671_33971 , \33676_33976 );
and \U$25183 ( \33872_34172 , \33667_33967 , \33676_33976 );
or \U$25184 ( \33873_34173 , \33870_34170 , \33871_34171 , \33872_34172 );
xor \U$25185 ( \33874_34174 , \33869_34169 , \33873_34173 );
and \U$25186 ( \33875_34175 , \33682_33982 , \33686_33986 );
and \U$25187 ( \33876_34176 , \33686_33986 , \33691_33991 );
and \U$25188 ( \33877_34177 , \33682_33982 , \33691_33991 );
or \U$25189 ( \33878_34178 , \33875_34175 , \33876_34176 , \33877_34177 );
xor \U$25190 ( \33879_34179 , \33874_34174 , \33878_34178 );
xor \U$25191 ( \33880_34180 , \33865_34165 , \33879_34179 );
xor \U$25192 ( \33881_34181 , \33856_34156 , \33880_34180 );
xor \U$25193 ( \33882_34182 , \33847_34147 , \33881_34181 );
and \U$25194 ( \33883_34183 , \33652_33952 , \33693_33993 );
and \U$25195 ( \33884_34184 , \33693_33993 , \33728_34028 );
and \U$25196 ( \33885_34185 , \33652_33952 , \33728_34028 );
or \U$25197 ( \33886_34186 , \33883_34183 , \33884_34184 , \33885_34185 );
and \U$25198 ( \33887_34187 , \33590_33890 , \33614_33914 );
and \U$25199 ( \33888_34188 , \33614_33914 , \33637_33937 );
and \U$25200 ( \33889_34189 , \33590_33890 , \33637_33937 );
or \U$25201 ( \33890_34190 , \33887_34187 , \33888_34188 , \33889_34189 );
xor \U$25202 ( \33891_34191 , \33886_34186 , \33890_34190 );
and \U$25203 ( \33892_34192 , \23315_23617 , \19235_19534 );
and \U$25204 ( \33893_34193 , \23900_24199 , \18743_19045 );
nor \U$25205 ( \33894_34194 , \33892_34192 , \33893_34193 );
xnor \U$25206 ( \33895_34195 , \33894_34194 , \19241_19540 );
and \U$25207 ( \33896_34196 , \14648_14950 , \28768_29070 );
and \U$25208 ( \33897_34197 , \15022_15321 , \28224_28526 );
nor \U$25209 ( \33898_34198 , \33896_34196 , \33897_34197 );
xnor \U$25210 ( \33899_34199 , \33898_34198 , \28774_29076 );
xor \U$25211 ( \33900_34200 , \33895_34195 , \33899_34199 );
and \U$25212 ( \33901_34201 , \13377_13679 , \30521_30823 );
and \U$25213 ( \33902_34202 , \13725_14024 , \29944_30246 );
nor \U$25214 ( \33903_34203 , \33901_34201 , \33902_34202 );
xnor \U$25215 ( \33904_34204 , \33903_34203 , \30511_30813 );
xor \U$25216 ( \33905_34205 , \33900_34200 , \33904_34204 );
and \U$25217 ( \33906_34206 , \26527_26829 , \16333_16635 );
and \U$25218 ( \33907_34207 , \27011_27313 , \15999_16301 );
nor \U$25219 ( \33908_34208 , \33906_34206 , \33907_34207 );
xnor \U$25220 ( \33909_34209 , \33908_34208 , \16323_16625 );
and \U$25221 ( \33910_34210 , \18730_19032 , \23839_24138 );
and \U$25222 ( \33911_34211 , \19259_19558 , \23328_23630 );
nor \U$25223 ( \33912_34212 , \33910_34210 , \33911_34211 );
xnor \U$25224 ( \33913_34213 , \33912_34212 , \23845_24144 );
xor \U$25225 ( \33914_34214 , \33909_34209 , \33913_34213 );
and \U$25226 ( \33915_34215 , \17325_17627 , \25527_25826 );
and \U$25227 ( \33916_34216 , \17736_18035 , \24962_25264 );
nor \U$25228 ( \33917_34217 , \33915_34215 , \33916_34216 );
xnor \U$25229 ( \33918_34218 , \33917_34217 , \25474_25773 );
xor \U$25230 ( \33919_34219 , \33914_34214 , \33918_34218 );
xor \U$25231 ( \33920_34220 , \33905_34205 , \33919_34219 );
and \U$25232 ( \33921_34221 , \29966_30268 , \13755_14054 );
and \U$25233 ( \33922_34222 , \30500_30802 , \13390_13692 );
nor \U$25234 ( \33923_34223 , \33921_34221 , \33922_34222 );
xnor \U$25235 ( \33924_34224 , \33923_34223 , \13736_14035 );
and \U$25236 ( \33925_34225 , \24970_25272 , \17791_18090 );
and \U$25237 ( \33926_34226 , \25516_25815 , \17353_17655 );
nor \U$25238 ( \33927_34227 , \33925_34225 , \33926_34226 );
xnor \U$25239 ( \33928_34228 , \33927_34227 , \17747_18046 );
xor \U$25240 ( \33929_34229 , \33924_34224 , \33928_34228 );
and \U$25241 ( \33930_34230 , \15965_16267 , \27095_27397 );
and \U$25242 ( \33931_34231 , \16353_16655 , \26505_26807 );
nor \U$25243 ( \33932_34232 , \33930_34230 , \33931_34231 );
xnor \U$25244 ( \33933_34233 , \33932_34232 , \26993_27295 );
xor \U$25245 ( \33934_34234 , \33929_34229 , \33933_34233 );
xor \U$25246 ( \33935_34235 , \33920_34220 , \33934_34234 );
and \U$25247 ( \33936_34236 , \33702_34002 , \33706_34006 );
and \U$25248 ( \33937_34237 , \33706_34006 , \33711_34011 );
and \U$25249 ( \33938_34238 , \33702_34002 , \33711_34011 );
or \U$25250 ( \33939_34239 , \33936_34236 , \33937_34237 , \33938_34238 );
not \U$25251 ( \33940_34240 , \11281_11580 );
and \U$25252 ( \33941_34241 , \31752_32054 , \12491_12790 );
and \U$25253 ( \33942_34242 , \32495_32794 , \12159_12461 );
nor \U$25254 ( \33943_34243 , \33941_34241 , \33942_34242 );
xnor \U$25255 ( \33944_34244 , \33943_34243 , \12481_12780 );
xor \U$25256 ( \33945_34245 , \33940_34240 , \33944_34244 );
and \U$25257 ( \33946_34246 , \28232_28534 , \15037_15336 );
and \U$25258 ( \33947_34247 , \28782_29084 , \14661_14963 );
nor \U$25259 ( \33948_34248 , \33946_34246 , \33947_34247 );
xnor \U$25260 ( \33949_34249 , \33948_34248 , \15043_15342 );
xor \U$25261 ( \33950_34250 , \33945_34245 , \33949_34249 );
xor \U$25262 ( \33951_34251 , \33939_34239 , \33950_34250 );
and \U$25263 ( \33952_34252 , \21788_22090 , \20706_21005 );
and \U$25264 ( \33953_34253 , \22257_22556 , \20255_20557 );
nor \U$25265 ( \33954_34254 , \33952_34252 , \33953_34253 );
xnor \U$25266 ( \33955_34255 , \33954_34254 , \20712_21011 );
and \U$25267 ( \33956_34256 , \20242_20544 , \22243_22542 );
and \U$25268 ( \33957_34257 , \20734_21033 , \21801_22103 );
nor \U$25269 ( \33958_34258 , \33956_34256 , \33957_34257 );
xnor \U$25270 ( \33959_34259 , \33958_34258 , \22249_22548 );
xor \U$25271 ( \33960_34260 , \33955_34255 , \33959_34259 );
and \U$25272 ( \33961_34261 , \11287_11586 , \32503_32802 );
xor \U$25273 ( \33962_34262 , \33960_34260 , \33961_34261 );
xor \U$25274 ( \33963_34263 , \33951_34251 , \33962_34262 );
xor \U$25275 ( \33964_34264 , \33935_34235 , \33963_34263 );
and \U$25276 ( \33965_34265 , \33603_33903 , \33607_33907 );
and \U$25277 ( \33966_34266 , \33607_33907 , \33612_33912 );
and \U$25278 ( \33967_34267 , \33603_33903 , \33612_33912 );
or \U$25279 ( \33968_34268 , \33965_34265 , \33966_34266 , \33967_34267 );
and \U$25280 ( \33969_34269 , \33628_33928 , \33630_33930 );
and \U$25281 ( \33970_34270 , \33630_33930 , \33635_33935 );
and \U$25282 ( \33971_34271 , \33628_33928 , \33635_33935 );
or \U$25283 ( \33972_34272 , \33969_34269 , \33970_34270 , \33971_34271 );
xor \U$25284 ( \33973_34273 , \33968_34268 , \33972_34272 );
and \U$25285 ( \33974_34274 , \33656_33956 , \33660_33960 );
and \U$25286 ( \33975_34275 , \33660_33960 , \33662_33962 );
and \U$25287 ( \33976_34276 , \33656_33956 , \33662_33962 );
or \U$25288 ( \33977_34277 , \33974_34274 , \33975_34275 , \33976_34276 );
buf \U$25289 ( \33978_34278 , \33634_33934 );
xor \U$25290 ( \33979_34279 , \33977_34277 , \33978_34278 );
and \U$25291 ( \33980_34280 , \12146_12448 , \32555_32854 );
and \U$25292 ( \33981_34281 , \12470_12769 , \31765_32067 );
nor \U$25293 ( \33982_34282 , \33980_34280 , \33981_34281 );
xnor \U$25294 ( \33983_34283 , \33982_34282 , \32506_32805 );
xor \U$25295 ( \33984_34284 , \33979_34279 , \33983_34283 );
xor \U$25296 ( \33985_34285 , \33973_34273 , \33984_34284 );
xor \U$25297 ( \33986_34286 , \33964_34264 , \33985_34285 );
xor \U$25298 ( \33987_34287 , \33891_34191 , \33986_34286 );
xor \U$25299 ( \33988_34288 , \33882_34182 , \33987_34287 );
xor \U$25300 ( \33989_34289 , \33843_34143 , \33988_34288 );
and \U$25301 ( \33990_34290 , \33731_34031 , \33735_34035 );
and \U$25302 ( \33991_34291 , \33736_34036 , \33739_34039 );
or \U$25303 ( \33992_34292 , \33990_34290 , \33991_34291 );
xor \U$25304 ( \33993_34293 , \33989_34289 , \33992_34292 );
buf g9ba5_GF_PartitionCandidate( \33994_34294_nG9ba5 , \33993_34293 );
and \U$25305 ( \33995_34295 , \10402_10704 , \33994_34294_nG9ba5 );
or \U$25306 ( \33996_34296 , \33839_34139 , \33995_34295 );
xor \U$25307 ( \33997_34297 , \10399_10703 , \33996_34296 );
buf \U$25308 ( \33998_34298 , \33997_34297 );
buf \U$25310 ( \33999_34299 , \33998_34298 );
xor \U$25311 ( \34000_34300 , \33838_34138 , \33999_34299 );
buf \U$25312 ( \34001_34301 , \34000_34300 );
and \U$25313 ( \34002_34302 , \33519_33819 , \33554_33854 );
and \U$25314 ( \34003_34303 , \33519_33819 , \33560_33860 );
and \U$25315 ( \34004_34304 , \33554_33854 , \33560_33860 );
or \U$25316 ( \34005_34305 , \34002_34302 , \34003_34303 , \34004_34304 );
buf \U$25317 ( \34006_34306 , \34005_34305 );
xor \U$25318 ( \34007_34307 , \34001_34301 , \34006_34306 );
and \U$25319 ( \34008_34308 , \33424_33724 , \33459_33759 );
and \U$25320 ( \34009_34309 , \33424_33724 , \33466_33766 );
and \U$25321 ( \34010_34310 , \33459_33759 , \33466_33766 );
or \U$25322 ( \34011_34311 , \34008_34308 , \34009_34309 , \34010_34310 );
buf \U$25323 ( \34012_34312 , \34011_34311 );
and \U$25324 ( \34013_34313 , \33473_33773 , \33493_33793 );
and \U$25325 ( \34014_34314 , \33473_33773 , \33500_33800 );
and \U$25326 ( \34015_34315 , \33493_33793 , \33500_33800 );
or \U$25327 ( \34016_34316 , \34013_34313 , \34014_34314 , \34015_34315 );
buf \U$25328 ( \34017_34317 , \34016_34316 );
xor \U$25329 ( \34018_34318 , \34012_34312 , \34017_34317 );
and \U$25330 ( \34019_34319 , \13431_13370 , \30064_30366_nG9bba );
and \U$25331 ( \34020_34320 , \13068_13367 , \30638_30940_nG9bb7 );
or \U$25332 ( \34021_34321 , \34019_34319 , \34020_34320 );
xor \U$25333 ( \34022_34322 , \13067_13366 , \34021_34321 );
buf \U$25334 ( \34023_34323 , \34022_34322 );
buf \U$25336 ( \34024_34324 , \34023_34323 );
xor \U$25337 ( \34025_34325 , \34018_34318 , \34024_34324 );
buf \U$25338 ( \34026_34326 , \34025_34325 );
and \U$25339 ( \34027_34327 , \33442_33742 , \33448_33748 );
buf \U$25340 ( \34028_34328 , \34027_34327 );
and \U$25341 ( \34029_34329 , \28946_28118 , \14682_14984_nG9bf6 );
and \U$25342 ( \34030_34330 , \27816_28115 , \15074_15373_nG9bf3 );
or \U$25343 ( \34031_34331 , \34029_34329 , \34030_34330 );
xor \U$25344 ( \34032_34332 , \27815_28114 , \34031_34331 );
buf \U$25345 ( \34033_34333 , \34032_34332 );
buf \U$25347 ( \34034_34334 , \34033_34333 );
xor \U$25348 ( \34035_34335 , \34028_34328 , \34034_34334 );
and \U$25349 ( \34036_34336 , \27141_26431 , \16013_16315_nG9bf0 );
and \U$25350 ( \34037_34337 , \26129_26428 , \16378_16680_nG9bed );
or \U$25351 ( \34038_34338 , \34036_34336 , \34037_34337 );
xor \U$25352 ( \34039_34339 , \26128_26427 , \34038_34338 );
buf \U$25353 ( \34040_34340 , \34039_34339 );
buf \U$25355 ( \34041_34341 , \34040_34340 );
xor \U$25356 ( \34042_34342 , \34035_34335 , \34041_34341 );
buf \U$25357 ( \34043_34343 , \34042_34342 );
and \U$25358 ( \34044_34344 , \23495_23201 , \18789_19091_nG9be4 );
and \U$25359 ( \34045_34345 , \22899_23198 , \19287_19586_nG9be1 );
or \U$25360 ( \34046_34346 , \34044_34344 , \34045_34345 );
xor \U$25361 ( \34047_34347 , \22898_23197 , \34046_34346 );
buf \U$25362 ( \34048_34348 , \34047_34347 );
buf \U$25364 ( \34049_34349 , \34048_34348 );
xor \U$25365 ( \34050_34350 , \34043_34343 , \34049_34349 );
and \U$25366 ( \34051_34351 , \21908_21658 , \20306_20608_nG9bde );
and \U$25367 ( \34052_34352 , \21356_21655 , \20787_21086_nG9bdb );
or \U$25368 ( \34053_34353 , \34051_34351 , \34052_34352 );
xor \U$25369 ( \34054_34354 , \21355_21654 , \34053_34353 );
buf \U$25370 ( \34055_34355 , \34054_34354 );
buf \U$25372 ( \34056_34356 , \34055_34355 );
xor \U$25373 ( \34057_34357 , \34050_34350 , \34056_34356 );
buf \U$25374 ( \34058_34358 , \34057_34357 );
and \U$25375 ( \34059_34359 , \17437_17297 , \24996_25298_nG9bcc );
and \U$25376 ( \34060_34360 , \16995_17294 , \25561_25860_nG9bc9 );
or \U$25377 ( \34061_34361 , \34059_34359 , \34060_34360 );
xor \U$25378 ( \34062_34362 , \16994_17293 , \34061_34361 );
buf \U$25379 ( \34063_34363 , \34062_34362 );
buf \U$25381 ( \34064_34364 , \34063_34363 );
xor \U$25382 ( \34065_34365 , \34058_34358 , \34064_34364 );
and \U$25383 ( \34066_34366 , \14710_14631 , \28300_28602_nG9bc0 );
and \U$25384 ( \34067_34367 , \14329_14628 , \28877_29179_nG9bbd );
or \U$25385 ( \34068_34368 , \34066_34366 , \34067_34367 );
xor \U$25386 ( \34069_34369 , \14328_14627 , \34068_34368 );
buf \U$25387 ( \34070_34370 , \34069_34369 );
buf \U$25389 ( \34071_34371 , \34070_34370 );
xor \U$25390 ( \34072_34372 , \34065_34365 , \34071_34371 );
buf \U$25391 ( \34073_34373 , \34072_34372 );
xor \U$25392 ( \34074_34374 , \34026_34326 , \34073_34373 );
and \U$25393 ( \34075_34375 , \33403_33703 , \33409_33709 );
and \U$25394 ( \34076_34376 , \33403_33703 , \33416_33716 );
and \U$25395 ( \34077_34377 , \33409_33709 , \33416_33716 );
or \U$25396 ( \34078_34378 , \34075_34375 , \34076_34376 , \34077_34377 );
buf \U$25397 ( \34079_34379 , \34078_34378 );
xor \U$25398 ( \34080_34380 , \34074_34374 , \34079_34379 );
buf \U$25399 ( \34081_34381 , \34080_34380 );
xor \U$25400 ( \34082_34382 , \34007_34307 , \34081_34381 );
buf \U$25401 ( \34083_34383 , \34082_34382 );
xor \U$25402 ( \34084_34384 , \33780_34080 , \34083_34383 );
and \U$25403 ( \34085_34385 , \33397_33697 , \33418_33718 );
and \U$25404 ( \34086_34386 , \33397_33697 , \33511_33811 );
and \U$25405 ( \34087_34387 , \33418_33718 , \33511_33811 );
or \U$25406 ( \34088_34388 , \34085_34385 , \34086_34386 , \34087_34387 );
buf \U$25407 ( \34089_34389 , \34088_34388 );
and \U$25408 ( \34090_34390 , \33748_34048 , \33753_34053 );
and \U$25409 ( \34091_34391 , \33748_34048 , \33759_34059 );
and \U$25410 ( \34092_34392 , \33753_34053 , \33759_34059 );
or \U$25411 ( \34093_34393 , \34090_34390 , \34091_34391 , \34092_34392 );
buf \U$25412 ( \34094_34394 , \34093_34393 );
xor \U$25413 ( \34095_34395 , \34089_34389 , \34094_34394 );
and \U$25414 ( \34096_34396 , \33575_33875 , \33580_33880 );
and \U$25415 ( \34097_34397 , \33575_33875 , \33746_34046 );
and \U$25416 ( \34098_34398 , \33580_33880 , \33746_34046 );
or \U$25417 ( \34099_34399 , \34096_34396 , \34097_34397 , \34098_34398 );
buf \U$25418 ( \34100_34400 , \34099_34399 );
and \U$25419 ( \34101_34401 , \33429_33729 , \33450_33750 );
and \U$25420 ( \34102_34402 , \33429_33729 , \33457_33757 );
and \U$25421 ( \34103_34403 , \33450_33750 , \33457_33757 );
or \U$25422 ( \34104_34404 , \34101_34401 , \34102_34402 , \34103_34403 );
buf \U$25423 ( \34105_34405 , \34104_34404 );
and \U$25424 ( \34106_34406 , \20353_20155 , \21827_22129_nG9bd8 );
and \U$25425 ( \34107_34407 , \19853_20152 , \22330_22629_nG9bd5 );
or \U$25426 ( \34108_34408 , \34106_34406 , \34107_34407 );
xor \U$25427 ( \34109_34409 , \19852_20151 , \34108_34408 );
buf \U$25428 ( \34110_34410 , \34109_34409 );
buf \U$25430 ( \34111_34411 , \34110_34410 );
xor \U$25431 ( \34112_34412 , \34105_34405 , \34111_34411 );
and \U$25432 ( \34113_34413 , \18908_18702 , \23394_23696_nG9bd2 );
and \U$25433 ( \34114_34414 , \18400_18699 , \23927_24226_nG9bcf );
or \U$25434 ( \34115_34415 , \34113_34413 , \34114_34414 );
xor \U$25435 ( \34116_34416 , \18399_18698 , \34115_34415 );
buf \U$25436 ( \34117_34417 , \34116_34416 );
buf \U$25438 ( \34118_34418 , \34117_34417 );
xor \U$25439 ( \34119_34419 , \34112_34412 , \34118_34418 );
buf \U$25440 ( \34120_34420 , \34119_34419 );
and \U$25441 ( \34121_34421 , \12183_12157 , \31877_32179_nG9bb4 );
and \U$25442 ( \34122_34422 , \11855_12154 , \32589_32888_nG9bb1 );
or \U$25443 ( \34123_34423 , \34121_34421 , \34122_34422 );
xor \U$25444 ( \34124_34424 , \11854_12153 , \34123_34423 );
buf \U$25445 ( \34125_34425 , \34124_34424 );
buf \U$25447 ( \34126_34426 , \34125_34425 );
xor \U$25448 ( \34127_34427 , \34120_34420 , \34126_34426 );
and \U$25449 ( \34128_34428 , \10996_10421 , \32881_33181_nG9bae );
and \U$25450 ( \34129_34429 , \10119_10418 , \33313_33613_nG9bab );
or \U$25451 ( \34130_34430 , \34128_34428 , \34129_34429 );
xor \U$25452 ( \34131_34431 , \10118_10417 , \34130_34430 );
buf \U$25453 ( \34132_34432 , \34131_34431 );
buf \U$25455 ( \34133_34433 , \34132_34432 );
xor \U$25456 ( \34134_34434 , \34127_34427 , \34133_34433 );
buf \U$25457 ( \34135_34435 , \34134_34434 );
xor \U$25458 ( \34136_34436 , \34100_34400 , \34135_34435 );
and \U$25459 ( \34137_34437 , \33468_33768 , \33502_33802 );
and \U$25460 ( \34138_34438 , \33468_33768 , \33509_33809 );
and \U$25461 ( \34139_34439 , \33502_33802 , \33509_33809 );
or \U$25462 ( \34140_34440 , \34137_34437 , \34138_34438 , \34139_34439 );
buf \U$25463 ( \34141_34441 , \34140_34440 );
xor \U$25464 ( \34142_34442 , \34136_34436 , \34141_34441 );
buf \U$25465 ( \34143_34443 , \34142_34442 );
xor \U$25466 ( \34144_34444 , \34095_34395 , \34143_34443 );
buf \U$25467 ( \34145_34445 , \34144_34444 );
xor \U$25468 ( \34146_34446 , \34084_34384 , \34145_34445 );
and \U$25469 ( \34147_34447 , \33775_34075 , \34146_34446 );
and \U$25471 ( \34148_34448 , \33769_34069 , \33774_34074 );
or \U$25473 ( \34149_34449 , 1'b0 , \34148_34448 , 1'b0 );
xor \U$25474 ( \34150_34450 , \34147_34447 , \34149_34449 );
and \U$25475 ( \34151_34451 , \33765_34065 , \33767_34067 );
or \U$25478 ( \34152_34452 , \34151_34451 , 1'b0 , 1'b0 );
xor \U$25479 ( \34153_34453 , \34150_34450 , \34152_34452 );
xor \U$25486 ( \34154_34454 , \34153_34453 , 1'b0 );
and \U$25487 ( \34155_34455 , \33780_34080 , \34083_34383 );
and \U$25488 ( \34156_34456 , \33780_34080 , \34145_34445 );
and \U$25489 ( \34157_34457 , \34083_34383 , \34145_34445 );
or \U$25490 ( \34158_34458 , \34155_34455 , \34156_34456 , \34157_34457 );
xor \U$25491 ( \34159_34459 , \34154_34454 , \34158_34458 );
and \U$25492 ( \34160_34460 , \34001_34301 , \34006_34306 );
and \U$25493 ( \34161_34461 , \34001_34301 , \34081_34381 );
and \U$25494 ( \34162_34462 , \34006_34306 , \34081_34381 );
or \U$25495 ( \34163_34463 , \34160_34460 , \34161_34461 , \34162_34462 );
buf \U$25496 ( \34164_34464 , \34163_34463 );
and \U$25497 ( \34165_34465 , \33785_34085 , \33809_34109 );
and \U$25498 ( \34166_34466 , \33785_34085 , \33816_34116 );
and \U$25499 ( \34167_34467 , \33809_34109 , \33816_34116 );
or \U$25500 ( \34168_34468 , \34165_34465 , \34166_34466 , \34167_34467 );
buf \U$25501 ( \34169_34469 , \34168_34468 );
and \U$25502 ( \34170_34470 , \20353_20155 , \22330_22629_nG9bd5 );
and \U$25503 ( \34171_34471 , \19853_20152 , \23394_23696_nG9bd2 );
or \U$25504 ( \34172_34472 , \34170_34470 , \34171_34471 );
xor \U$25505 ( \34173_34473 , \19852_20151 , \34172_34472 );
buf \U$25506 ( \34174_34474 , \34173_34473 );
buf \U$25508 ( \34175_34475 , \34174_34474 );
xor \U$25509 ( \34176_34476 , \34169_34469 , \34175_34475 );
and \U$25510 ( \34177_34477 , \18908_18702 , \23927_24226_nG9bcf );
and \U$25511 ( \34178_34478 , \18400_18699 , \24996_25298_nG9bcc );
or \U$25512 ( \34179_34479 , \34177_34477 , \34178_34478 );
xor \U$25513 ( \34180_34480 , \18399_18698 , \34179_34479 );
buf \U$25514 ( \34181_34481 , \34180_34480 );
buf \U$25516 ( \34182_34482 , \34181_34481 );
xor \U$25517 ( \34183_34483 , \34176_34476 , \34182_34482 );
buf \U$25518 ( \34184_34484 , \34183_34483 );
and \U$25519 ( \34185_34485 , \12183_12157 , \32589_32888_nG9bb1 );
and \U$25520 ( \34186_34486 , \11855_12154 , \32881_33181_nG9bae );
or \U$25521 ( \34187_34487 , \34185_34485 , \34186_34486 );
xor \U$25522 ( \34188_34488 , \11854_12153 , \34187_34487 );
buf \U$25523 ( \34189_34489 , \34188_34488 );
buf \U$25525 ( \34190_34490 , \34189_34489 );
xor \U$25526 ( \34191_34491 , \34184_34484 , \34190_34490 );
and \U$25527 ( \34192_34492 , \10411_10707 , \33994_34294_nG9ba5 );
and \U$25528 ( \34193_34493 , \33886_34186 , \33890_34190 );
and \U$25529 ( \34194_34494 , \33890_34190 , \33986_34286 );
and \U$25530 ( \34195_34495 , \33886_34186 , \33986_34286 );
or \U$25531 ( \34196_34496 , \34193_34493 , \34194_34494 , \34195_34495 );
and \U$25532 ( \34197_34497 , \33860_34160 , \33864_34164 );
and \U$25533 ( \34198_34498 , \33864_34164 , \33879_34179 );
and \U$25534 ( \34199_34499 , \33860_34160 , \33879_34179 );
or \U$25535 ( \34200_34500 , \34197_34497 , \34198_34498 , \34199_34499 );
and \U$25536 ( \34201_34501 , \33869_34169 , \33873_34173 );
and \U$25537 ( \34202_34502 , \33873_34173 , \33878_34178 );
and \U$25538 ( \34203_34503 , \33869_34169 , \33878_34178 );
or \U$25539 ( \34204_34504 , \34201_34501 , \34202_34502 , \34203_34503 );
and \U$25540 ( \34205_34505 , \33977_34277 , \33978_34278 );
and \U$25541 ( \34206_34506 , \33978_34278 , \33983_34283 );
and \U$25542 ( \34207_34507 , \33977_34277 , \33983_34283 );
or \U$25543 ( \34208_34508 , \34205_34505 , \34206_34506 , \34207_34507 );
xor \U$25544 ( \34209_34509 , \34204_34504 , \34208_34508 );
and \U$25545 ( \34210_34510 , \32495_32794 , \12491_12790 );
not \U$25546 ( \34211_34511 , \34210_34510 );
xnor \U$25547 ( \34212_34512 , \34211_34511 , \12481_12780 );
not \U$25548 ( \34213_34513 , \34212_34512 );
and \U$25549 ( \34214_34514 , \12470_12769 , \32555_32854 );
and \U$25550 ( \34215_34515 , \13377_13679 , \31765_32067 );
nor \U$25551 ( \34216_34516 , \34214_34514 , \34215_34515 );
xnor \U$25552 ( \34217_34517 , \34216_34516 , \32506_32805 );
xor \U$25553 ( \34218_34518 , \34213_34513 , \34217_34517 );
and \U$25554 ( \34219_34519 , \12146_12448 , \32503_32802 );
xor \U$25555 ( \34220_34520 , \34218_34518 , \34219_34519 );
xor \U$25556 ( \34221_34521 , \34209_34509 , \34220_34520 );
xor \U$25557 ( \34222_34522 , \34200_34500 , \34221_34521 );
and \U$25558 ( \34223_34523 , \33939_34239 , \33950_34250 );
and \U$25559 ( \34224_34524 , \33950_34250 , \33962_34262 );
and \U$25560 ( \34225_34525 , \33939_34239 , \33962_34262 );
or \U$25561 ( \34226_34526 , \34223_34523 , \34224_34524 , \34225_34525 );
and \U$25562 ( \34227_34527 , \33940_34240 , \33944_34244 );
and \U$25563 ( \34228_34528 , \33944_34244 , \33949_34249 );
and \U$25564 ( \34229_34529 , \33940_34240 , \33949_34249 );
or \U$25565 ( \34230_34530 , \34227_34527 , \34228_34528 , \34229_34529 );
and \U$25566 ( \34231_34531 , \33955_34255 , \33959_34259 );
and \U$25567 ( \34232_34532 , \33959_34259 , \33961_34261 );
and \U$25568 ( \34233_34533 , \33955_34255 , \33961_34261 );
or \U$25569 ( \34234_34534 , \34231_34531 , \34232_34532 , \34233_34533 );
xor \U$25570 ( \34235_34535 , \34230_34530 , \34234_34534 );
and \U$25571 ( \34236_34536 , \33909_34209 , \33913_34213 );
and \U$25572 ( \34237_34537 , \33913_34213 , \33918_34218 );
and \U$25573 ( \34238_34538 , \33909_34209 , \33918_34218 );
or \U$25574 ( \34239_34539 , \34236_34536 , \34237_34537 , \34238_34538 );
xor \U$25575 ( \34240_34540 , \34235_34535 , \34239_34539 );
xor \U$25576 ( \34241_34541 , \34226_34526 , \34240_34540 );
and \U$25577 ( \34242_34542 , \33895_34195 , \33899_34199 );
and \U$25578 ( \34243_34543 , \33899_34199 , \33904_34204 );
and \U$25579 ( \34244_34544 , \33895_34195 , \33904_34204 );
or \U$25580 ( \34245_34545 , \34242_34542 , \34243_34543 , \34244_34544 );
and \U$25581 ( \34246_34546 , \33924_34224 , \33928_34228 );
and \U$25582 ( \34247_34547 , \33928_34228 , \33933_34233 );
and \U$25583 ( \34248_34548 , \33924_34224 , \33933_34233 );
or \U$25584 ( \34249_34549 , \34246_34546 , \34247_34547 , \34248_34548 );
xor \U$25585 ( \34250_34550 , \34245_34545 , \34249_34549 );
and \U$25586 ( \34251_34551 , \30500_30802 , \13755_14054 );
and \U$25587 ( \34252_34552 , \31752_32054 , \13390_13692 );
nor \U$25588 ( \34253_34553 , \34251_34551 , \34252_34552 );
xnor \U$25589 ( \34254_34554 , \34253_34553 , \13736_14035 );
and \U$25590 ( \34255_34555 , \27011_27313 , \16333_16635 );
and \U$25591 ( \34256_34556 , \28232_28534 , \15999_16301 );
nor \U$25592 ( \34257_34557 , \34255_34555 , \34256_34556 );
xnor \U$25593 ( \34258_34558 , \34257_34557 , \16323_16625 );
xor \U$25594 ( \34259_34559 , \34254_34554 , \34258_34558 );
and \U$25595 ( \34260_34560 , \20734_21033 , \22243_22542 );
and \U$25596 ( \34261_34561 , \21788_22090 , \21801_22103 );
nor \U$25597 ( \34262_34562 , \34260_34560 , \34261_34561 );
xnor \U$25598 ( \34263_34563 , \34262_34562 , \22249_22548 );
xor \U$25599 ( \34264_34564 , \34259_34559 , \34263_34563 );
xor \U$25600 ( \34265_34565 , \34250_34550 , \34264_34564 );
xor \U$25601 ( \34266_34566 , \34241_34541 , \34265_34565 );
xor \U$25602 ( \34267_34567 , \34222_34522 , \34266_34566 );
xor \U$25603 ( \34268_34568 , \34196_34496 , \34267_34567 );
and \U$25604 ( \34269_34569 , \33851_34151 , \33855_34155 );
and \U$25605 ( \34270_34570 , \33855_34155 , \33880_34180 );
and \U$25606 ( \34271_34571 , \33851_34151 , \33880_34180 );
or \U$25607 ( \34272_34572 , \34269_34569 , \34270_34570 , \34271_34571 );
and \U$25608 ( \34273_34573 , \33935_34235 , \33963_34263 );
and \U$25609 ( \34274_34574 , \33963_34263 , \33985_34285 );
and \U$25610 ( \34275_34575 , \33935_34235 , \33985_34285 );
or \U$25611 ( \34276_34576 , \34273_34573 , \34274_34574 , \34275_34575 );
xor \U$25612 ( \34277_34577 , \34272_34572 , \34276_34576 );
and \U$25613 ( \34278_34578 , \33905_34205 , \33919_34219 );
and \U$25614 ( \34279_34579 , \33919_34219 , \33934_34234 );
and \U$25615 ( \34280_34580 , \33905_34205 , \33934_34234 );
or \U$25616 ( \34281_34581 , \34278_34578 , \34279_34579 , \34280_34580 );
and \U$25617 ( \34282_34582 , \33968_34268 , \33972_34272 );
and \U$25618 ( \34283_34583 , \33972_34272 , \33984_34284 );
and \U$25619 ( \34284_34584 , \33968_34268 , \33984_34284 );
or \U$25620 ( \34285_34585 , \34282_34582 , \34283_34583 , \34284_34584 );
xor \U$25621 ( \34286_34586 , \34281_34581 , \34285_34585 );
and \U$25622 ( \34287_34587 , \22257_22556 , \20706_21005 );
and \U$25623 ( \34288_34588 , \23315_23617 , \20255_20557 );
nor \U$25624 ( \34289_34589 , \34287_34587 , \34288_34588 );
xnor \U$25625 ( \34290_34590 , \34289_34589 , \20712_21011 );
and \U$25626 ( \34291_34591 , \15022_15321 , \28768_29070 );
and \U$25627 ( \34292_34592 , \15965_16267 , \28224_28526 );
nor \U$25628 ( \34293_34593 , \34291_34591 , \34292_34592 );
xnor \U$25629 ( \34294_34594 , \34293_34593 , \28774_29076 );
xor \U$25630 ( \34295_34595 , \34290_34590 , \34294_34594 );
and \U$25631 ( \34296_34596 , \13725_14024 , \30521_30823 );
and \U$25632 ( \34297_34597 , \14648_14950 , \29944_30246 );
nor \U$25633 ( \34298_34598 , \34296_34596 , \34297_34597 );
xnor \U$25634 ( \34299_34599 , \34298_34598 , \30511_30813 );
xor \U$25635 ( \34300_34600 , \34295_34595 , \34299_34599 );
and \U$25636 ( \34301_34601 , \25516_25815 , \17791_18090 );
and \U$25637 ( \34302_34602 , \26527_26829 , \17353_17655 );
nor \U$25638 ( \34303_34603 , \34301_34601 , \34302_34602 );
xnor \U$25639 ( \34304_34604 , \34303_34603 , \17747_18046 );
and \U$25640 ( \34305_34605 , \19259_19558 , \23839_24138 );
and \U$25641 ( \34306_34606 , \20242_20544 , \23328_23630 );
nor \U$25642 ( \34307_34607 , \34305_34605 , \34306_34606 );
xnor \U$25643 ( \34308_34608 , \34307_34607 , \23845_24144 );
xor \U$25644 ( \34309_34609 , \34304_34604 , \34308_34608 );
and \U$25645 ( \34310_34610 , \17736_18035 , \25527_25826 );
and \U$25646 ( \34311_34611 , \18730_19032 , \24962_25264 );
nor \U$25647 ( \34312_34612 , \34310_34610 , \34311_34611 );
xnor \U$25648 ( \34313_34613 , \34312_34612 , \25474_25773 );
xor \U$25649 ( \34314_34614 , \34309_34609 , \34313_34613 );
xor \U$25650 ( \34315_34615 , \34300_34600 , \34314_34614 );
and \U$25651 ( \34316_34616 , \28782_29084 , \15037_15336 );
and \U$25652 ( \34317_34617 , \29966_30268 , \14661_14963 );
nor \U$25653 ( \34318_34618 , \34316_34616 , \34317_34617 );
xnor \U$25654 ( \34319_34619 , \34318_34618 , \15043_15342 );
and \U$25655 ( \34320_34620 , \23900_24199 , \19235_19534 );
and \U$25656 ( \34321_34621 , \24970_25272 , \18743_19045 );
nor \U$25657 ( \34322_34622 , \34320_34620 , \34321_34621 );
xnor \U$25658 ( \34323_34623 , \34322_34622 , \19241_19540 );
xor \U$25659 ( \34324_34624 , \34319_34619 , \34323_34623 );
and \U$25660 ( \34325_34625 , \16353_16655 , \27095_27397 );
and \U$25661 ( \34326_34626 , \17325_17627 , \26505_26807 );
nor \U$25662 ( \34327_34627 , \34325_34625 , \34326_34626 );
xnor \U$25663 ( \34328_34628 , \34327_34627 , \26993_27295 );
xor \U$25664 ( \34329_34629 , \34324_34624 , \34328_34628 );
xor \U$25665 ( \34330_34630 , \34315_34615 , \34329_34629 );
xor \U$25666 ( \34331_34631 , \34286_34586 , \34330_34630 );
xor \U$25667 ( \34332_34632 , \34277_34577 , \34331_34631 );
xor \U$25668 ( \34333_34633 , \34268_34568 , \34332_34632 );
and \U$25669 ( \34334_34634 , \33847_34147 , \33881_34181 );
and \U$25670 ( \34335_34635 , \33881_34181 , \33987_34287 );
and \U$25671 ( \34336_34636 , \33847_34147 , \33987_34287 );
or \U$25672 ( \34337_34637 , \34334_34634 , \34335_34635 , \34336_34636 );
xor \U$25673 ( \34338_34638 , \34333_34633 , \34337_34637 );
and \U$25674 ( \34339_34639 , \33843_34143 , \33988_34288 );
and \U$25675 ( \34340_34640 , \33989_34289 , \33992_34292 );
or \U$25676 ( \34341_34641 , \34339_34639 , \34340_34640 );
xor \U$25677 ( \34342_34642 , \34338_34638 , \34341_34641 );
buf g9ba2_GF_PartitionCandidate( \34343_34643_nG9ba2 , \34342_34642 );
and \U$25678 ( \34344_34644 , \10402_10704 , \34343_34643_nG9ba2 );
or \U$25679 ( \34345_34645 , \34192_34492 , \34344_34644 );
xor \U$25680 ( \34346_34646 , \10399_10703 , \34345_34645 );
buf \U$25681 ( \34347_34647 , \34346_34646 );
buf \U$25683 ( \34348_34648 , \34347_34647 );
xor \U$25684 ( \34349_34649 , \34191_34491 , \34348_34648 );
buf \U$25685 ( \34350_34650 , \34349_34649 );
and \U$25686 ( \34351_34651 , \33832_34132 , \33837_34137 );
and \U$25687 ( \34352_34652 , \33832_34132 , \33999_34299 );
and \U$25688 ( \34353_34653 , \33837_34137 , \33999_34299 );
or \U$25689 ( \34354_34654 , \34351_34651 , \34352_34652 , \34353_34653 );
buf \U$25690 ( \34355_34655 , \34354_34654 );
xor \U$25691 ( \34356_34656 , \34350_34650 , \34355_34655 );
and \U$25692 ( \34357_34657 , \34105_34405 , \34111_34411 );
and \U$25693 ( \34358_34658 , \34105_34405 , \34118_34418 );
and \U$25694 ( \34359_34659 , \34111_34411 , \34118_34418 );
or \U$25695 ( \34360_34660 , \34357_34657 , \34358_34658 , \34359_34659 );
buf \U$25696 ( \34361_34661 , \34360_34660 );
and \U$25697 ( \34362_34662 , \13431_13370 , \30638_30940_nG9bb7 );
and \U$25698 ( \34363_34663 , \13068_13367 , \31877_32179_nG9bb4 );
or \U$25699 ( \34364_34664 , \34362_34662 , \34363_34663 );
xor \U$25700 ( \34365_34665 , \13067_13366 , \34364_34664 );
buf \U$25701 ( \34366_34666 , \34365_34665 );
buf \U$25703 ( \34367_34667 , \34366_34666 );
xor \U$25704 ( \34368_34668 , \34361_34661 , \34367_34667 );
and \U$25705 ( \34369_34669 , \10996_10421 , \33313_33613_nG9bab );
and \U$25706 ( \34370_34670 , \10119_10418 , \33741_34041_nG9ba8 );
or \U$25707 ( \34371_34671 , \34369_34669 , \34370_34670 );
xor \U$25708 ( \34372_34672 , \10118_10417 , \34371_34671 );
buf \U$25709 ( \34373_34673 , \34372_34672 );
buf \U$25711 ( \34374_34674 , \34373_34673 );
xor \U$25712 ( \34375_34675 , \34368_34668 , \34374_34674 );
buf \U$25713 ( \34376_34676 , \34375_34675 );
xor \U$25714 ( \34377_34677 , \34356_34656 , \34376_34676 );
buf \U$25715 ( \34378_34678 , \34377_34677 );
xor \U$25716 ( \34379_34679 , \34164_34464 , \34378_34678 );
and \U$25717 ( \34380_34680 , \34100_34400 , \34135_34435 );
and \U$25718 ( \34381_34681 , \34100_34400 , \34141_34441 );
and \U$25719 ( \34382_34682 , \34135_34435 , \34141_34441 );
or \U$25720 ( \34383_34683 , \34380_34680 , \34381_34681 , \34382_34682 );
buf \U$25721 ( \34384_34684 , \34383_34683 );
xor \U$25722 ( \34385_34685 , \34379_34679 , \34384_34684 );
buf \U$25723 ( \34386_34686 , \34385_34685 );
and \U$25724 ( \34387_34687 , \34089_34389 , \34094_34394 );
and \U$25725 ( \34388_34688 , \34089_34389 , \34143_34443 );
and \U$25726 ( \34389_34689 , \34094_34394 , \34143_34443 );
or \U$25727 ( \34390_34690 , \34387_34687 , \34388_34688 , \34389_34689 );
buf \U$25728 ( \34391_34691 , \34390_34690 );
xor \U$25729 ( \34392_34692 , \34386_34686 , \34391_34691 );
and \U$25730 ( \34393_34693 , \34120_34420 , \34126_34426 );
and \U$25731 ( \34394_34694 , \34120_34420 , \34133_34433 );
and \U$25732 ( \34395_34695 , \34126_34426 , \34133_34433 );
or \U$25733 ( \34396_34696 , \34393_34693 , \34394_34694 , \34395_34695 );
buf \U$25734 ( \34397_34697 , \34396_34696 );
and \U$25735 ( \34398_34698 , \34012_34312 , \34017_34317 );
and \U$25736 ( \34399_34699 , \34012_34312 , \34024_34324 );
and \U$25737 ( \34400_34700 , \34017_34317 , \34024_34324 );
or \U$25738 ( \34401_34701 , \34398_34698 , \34399_34699 , \34400_34700 );
buf \U$25739 ( \34402_34702 , \34401_34701 );
xor \U$25740 ( \34403_34703 , \34397_34697 , \34402_34702 );
and \U$25741 ( \34404_34704 , \34058_34358 , \34064_34364 );
and \U$25742 ( \34405_34705 , \34058_34358 , \34071_34371 );
and \U$25743 ( \34406_34706 , \34064_34364 , \34071_34371 );
or \U$25744 ( \34407_34707 , \34404_34704 , \34405_34705 , \34406_34706 );
buf \U$25745 ( \34408_34708 , \34407_34707 );
xor \U$25746 ( \34409_34709 , \34403_34703 , \34408_34708 );
buf \U$25747 ( \34410_34710 , \34409_34709 );
and \U$25748 ( \34411_34711 , \34026_34326 , \34073_34373 );
and \U$25749 ( \34412_34712 , \34026_34326 , \34079_34379 );
and \U$25750 ( \34413_34713 , \34073_34373 , \34079_34379 );
or \U$25751 ( \34414_34714 , \34411_34711 , \34412_34712 , \34413_34713 );
buf \U$25752 ( \34415_34715 , \34414_34714 );
xor \U$25753 ( \34416_34716 , \34410_34710 , \34415_34715 );
and \U$25754 ( \34417_34717 , \33798_34098 , \33800_34100 );
and \U$25755 ( \34418_34718 , \33798_34098 , \33807_34107 );
and \U$25756 ( \34419_34719 , \33800_34100 , \33807_34107 );
or \U$25757 ( \34420_34720 , \34417_34717 , \34418_34718 , \34419_34719 );
buf \U$25758 ( \34421_34721 , \34420_34720 );
and \U$25759 ( \34422_34722 , \28946_28118 , \15074_15373_nG9bf3 );
and \U$25760 ( \34423_34723 , \27816_28115 , \16013_16315_nG9bf0 );
or \U$25761 ( \34424_34724 , \34422_34722 , \34423_34723 );
xor \U$25762 ( \34425_34725 , \27815_28114 , \34424_34724 );
buf \U$25763 ( \34426_34726 , \34425_34725 );
buf \U$25765 ( \34427_34727 , \34426_34726 );
xor \U$25766 ( \34428_34728 , \34421_34721 , \34427_34727 );
and \U$25767 ( \34429_34729 , \27141_26431 , \16378_16680_nG9bed );
and \U$25768 ( \34430_34730 , \26129_26428 , \17363_17665_nG9bea );
or \U$25769 ( \34431_34731 , \34429_34729 , \34430_34730 );
xor \U$25770 ( \34432_34732 , \26128_26427 , \34431_34731 );
buf \U$25771 ( \34433_34733 , \34432_34732 );
buf \U$25773 ( \34434_34734 , \34433_34733 );
xor \U$25774 ( \34435_34735 , \34428_34728 , \34434_34734 );
buf \U$25775 ( \34436_34736 , \34435_34735 );
and \U$25776 ( \34437_34737 , \34028_34328 , \34034_34334 );
and \U$25777 ( \34438_34738 , \34028_34328 , \34041_34341 );
and \U$25778 ( \34439_34739 , \34034_34334 , \34041_34341 );
or \U$25779 ( \34440_34740 , \34437_34737 , \34438_34738 , \34439_34739 );
buf \U$25780 ( \34441_34741 , \34440_34740 );
xor \U$25781 ( \34442_34742 , \34436_34736 , \34441_34741 );
and \U$25782 ( \34443_34743 , \21908_21658 , \20787_21086_nG9bdb );
and \U$25783 ( \34444_34744 , \21356_21655 , \21827_22129_nG9bd8 );
or \U$25784 ( \34445_34745 , \34443_34743 , \34444_34744 );
xor \U$25785 ( \34446_34746 , \21355_21654 , \34445_34745 );
buf \U$25786 ( \34447_34747 , \34446_34746 );
buf \U$25788 ( \34448_34748 , \34447_34747 );
xor \U$25789 ( \34449_34749 , \34442_34742 , \34448_34748 );
buf \U$25790 ( \34450_34750 , \34449_34749 );
and \U$25791 ( \34451_34751 , \17437_17297 , \25561_25860_nG9bc9 );
and \U$25792 ( \34452_34752 , \16995_17294 , \26585_26887_nG9bc6 );
or \U$25793 ( \34453_34753 , \34451_34751 , \34452_34752 );
xor \U$25794 ( \34454_34754 , \16994_17293 , \34453_34753 );
buf \U$25795 ( \34455_34755 , \34454_34754 );
buf \U$25797 ( \34456_34756 , \34455_34755 );
xor \U$25798 ( \34457_34757 , \34450_34750 , \34456_34756 );
and \U$25799 ( \34458_34758 , \14710_14631 , \28877_29179_nG9bbd );
and \U$25800 ( \34459_34759 , \14329_14628 , \30064_30366_nG9bba );
or \U$25801 ( \34460_34760 , \34458_34758 , \34459_34759 );
xor \U$25802 ( \34461_34761 , \14328_14627 , \34460_34760 );
buf \U$25803 ( \34462_34762 , \34461_34761 );
buf \U$25805 ( \34463_34763 , \34462_34762 );
xor \U$25806 ( \34464_34764 , \34457_34757 , \34463_34763 );
buf \U$25807 ( \34465_34765 , \34464_34764 );
and \U$25809 ( \34466_34766 , \32617_32916 , \12168_12470_nG9c02 );
or \U$25810 ( \34467_34767 , 1'b0 , \34466_34766 );
xor \U$25811 ( \34468_34768 , 1'b0 , \34467_34767 );
buf \U$25812 ( \34469_34769 , \34468_34768 );
buf \U$25814 ( \34470_34770 , \34469_34769 );
and \U$25815 ( \34471_34771 , \31989_31636 , \12502_12801_nG9bff );
and \U$25816 ( \34472_34772 , \31334_31633 , \13403_13705_nG9bfc );
or \U$25817 ( \34473_34773 , \34471_34771 , \34472_34772 );
xor \U$25818 ( \34474_34774 , \31333_31632 , \34473_34773 );
buf \U$25819 ( \34475_34775 , \34474_34774 );
buf \U$25821 ( \34476_34776 , \34475_34775 );
xor \U$25822 ( \34477_34777 , \34470_34770 , \34476_34776 );
buf \U$25823 ( \34478_34778 , \34477_34777 );
and \U$25824 ( \34479_34779 , \33790_34090 , \33796_34096 );
buf \U$25825 ( \34480_34780 , \34479_34779 );
xor \U$25826 ( \34481_34781 , \34478_34778 , \34480_34780 );
and \U$25827 ( \34482_34782 , \30670_29853 , \13771_14070_nG9bf9 );
and \U$25828 ( \34483_34783 , \29551_29850 , \14682_14984_nG9bf6 );
or \U$25829 ( \34484_34784 , \34482_34782 , \34483_34783 );
xor \U$25830 ( \34485_34785 , \29550_29849 , \34484_34784 );
buf \U$25831 ( \34486_34786 , \34485_34785 );
buf \U$25833 ( \34487_34787 , \34486_34786 );
xor \U$25834 ( \34488_34788 , \34481_34781 , \34487_34787 );
buf \U$25835 ( \34489_34789 , \34488_34788 );
and \U$25836 ( \34490_34790 , \25044_24792 , \17808_18107_nG9be7 );
and \U$25837 ( \34491_34791 , \24490_24789 , \18789_19091_nG9be4 );
or \U$25838 ( \34492_34792 , \34490_34790 , \34491_34791 );
xor \U$25839 ( \34493_34793 , \24489_24788 , \34492_34792 );
buf \U$25840 ( \34494_34794 , \34493_34793 );
buf \U$25842 ( \34495_34795 , \34494_34794 );
xor \U$25843 ( \34496_34796 , \34489_34789 , \34495_34795 );
and \U$25844 ( \34497_34797 , \23495_23201 , \19287_19586_nG9be1 );
and \U$25845 ( \34498_34798 , \22899_23198 , \20306_20608_nG9bde );
or \U$25846 ( \34499_34799 , \34497_34797 , \34498_34798 );
xor \U$25847 ( \34500_34800 , \22898_23197 , \34499_34799 );
buf \U$25848 ( \34501_34801 , \34500_34800 );
buf \U$25850 ( \34502_34802 , \34501_34801 );
xor \U$25851 ( \34503_34803 , \34496_34796 , \34502_34802 );
buf \U$25852 ( \34504_34804 , \34503_34803 );
and \U$25853 ( \34505_34805 , \34043_34343 , \34049_34349 );
and \U$25854 ( \34506_34806 , \34043_34343 , \34056_34356 );
and \U$25855 ( \34507_34807 , \34049_34349 , \34056_34356 );
or \U$25856 ( \34508_34808 , \34505_34805 , \34506_34806 , \34507_34807 );
buf \U$25857 ( \34509_34809 , \34508_34808 );
xor \U$25858 ( \34510_34810 , \34504_34804 , \34509_34809 );
and \U$25859 ( \34511_34811 , \16405_15940 , \27114_27416_nG9bc3 );
and \U$25860 ( \34512_34812 , \15638_15937 , \28300_28602_nG9bc0 );
or \U$25861 ( \34513_34813 , \34511_34811 , \34512_34812 );
xor \U$25862 ( \34514_34814 , \15637_15936 , \34513_34813 );
buf \U$25863 ( \34515_34815 , \34514_34814 );
buf \U$25865 ( \34516_34816 , \34515_34815 );
xor \U$25866 ( \34517_34817 , \34510_34810 , \34516_34816 );
buf \U$25867 ( \34518_34818 , \34517_34817 );
xor \U$25868 ( \34519_34819 , \34465_34765 , \34518_34818 );
and \U$25869 ( \34520_34820 , \33818_34118 , \33823_34123 );
and \U$25870 ( \34521_34821 , \33818_34118 , \33830_34130 );
and \U$25871 ( \34522_34822 , \33823_34123 , \33830_34130 );
or \U$25872 ( \34523_34823 , \34520_34820 , \34521_34821 , \34522_34822 );
buf \U$25873 ( \34524_34824 , \34523_34823 );
xor \U$25874 ( \34525_34825 , \34519_34819 , \34524_34824 );
buf \U$25875 ( \34526_34826 , \34525_34825 );
xor \U$25876 ( \34527_34827 , \34416_34716 , \34526_34826 );
buf \U$25877 ( \34528_34828 , \34527_34827 );
xor \U$25878 ( \34529_34829 , \34392_34692 , \34528_34828 );
and \U$25879 ( \34530_34830 , \34159_34459 , \34529_34829 );
and \U$25881 ( \34531_34831 , \34153_34453 , \34158_34458 );
or \U$25883 ( \34532_34832 , 1'b0 , \34531_34831 , 1'b0 );
xor \U$25884 ( \34533_34833 , \34530_34830 , \34532_34832 );
and \U$25886 ( \34534_34834 , \34147_34447 , \34152_34452 );
or \U$25888 ( \34535_34835 , 1'b0 , \34534_34834 , 1'b0 );
xor \U$25889 ( \34536_34836 , \34533_34833 , \34535_34835 );
xor \U$25896 ( \34537_34837 , \34536_34836 , 1'b0 );
and \U$25897 ( \34538_34838 , \34386_34686 , \34391_34691 );
and \U$25898 ( \34539_34839 , \34386_34686 , \34528_34828 );
and \U$25899 ( \34540_34840 , \34391_34691 , \34528_34828 );
or \U$25900 ( \34541_34841 , \34538_34838 , \34539_34839 , \34540_34840 );
xor \U$25901 ( \34542_34842 , \34537_34837 , \34541_34841 );
and \U$25902 ( \34543_34843 , \34350_34650 , \34355_34655 );
and \U$25903 ( \34544_34844 , \34350_34650 , \34376_34676 );
and \U$25904 ( \34545_34845 , \34355_34655 , \34376_34676 );
or \U$25905 ( \34546_34846 , \34543_34843 , \34544_34844 , \34545_34845 );
buf \U$25906 ( \34547_34847 , \34546_34846 );
and \U$25907 ( \34548_34848 , \34397_34697 , \34402_34702 );
and \U$25908 ( \34549_34849 , \34397_34697 , \34408_34708 );
and \U$25909 ( \34550_34850 , \34402_34702 , \34408_34708 );
or \U$25910 ( \34551_34851 , \34548_34848 , \34549_34849 , \34550_34850 );
buf \U$25911 ( \34552_34852 , \34551_34851 );
xor \U$25912 ( \34553_34853 , \34547_34847 , \34552_34852 );
and \U$25913 ( \34554_34854 , \34450_34750 , \34456_34756 );
and \U$25914 ( \34555_34855 , \34450_34750 , \34463_34763 );
and \U$25915 ( \34556_34856 , \34456_34756 , \34463_34763 );
or \U$25916 ( \34557_34857 , \34554_34854 , \34555_34855 , \34556_34856 );
buf \U$25917 ( \34558_34858 , \34557_34857 );
and \U$25918 ( \34559_34859 , \34504_34804 , \34509_34809 );
and \U$25919 ( \34560_34860 , \34504_34804 , \34516_34816 );
and \U$25920 ( \34561_34861 , \34509_34809 , \34516_34816 );
or \U$25921 ( \34562_34862 , \34559_34859 , \34560_34860 , \34561_34861 );
buf \U$25922 ( \34563_34863 , \34562_34862 );
xor \U$25923 ( \34564_34864 , \34558_34858 , \34563_34863 );
and \U$25924 ( \34565_34865 , \34436_34736 , \34441_34741 );
and \U$25925 ( \34566_34866 , \34436_34736 , \34448_34748 );
and \U$25926 ( \34567_34867 , \34441_34741 , \34448_34748 );
or \U$25927 ( \34568_34868 , \34565_34865 , \34566_34866 , \34567_34867 );
buf \U$25928 ( \34569_34869 , \34568_34868 );
and \U$25930 ( \34570_34870 , \32617_32916 , \12502_12801_nG9bff );
or \U$25931 ( \34571_34871 , 1'b0 , \34570_34870 );
xor \U$25932 ( \34572_34872 , 1'b0 , \34571_34871 );
buf \U$25933 ( \34573_34873 , \34572_34872 );
buf \U$25935 ( \34574_34874 , \34573_34873 );
and \U$25936 ( \34575_34875 , \31989_31636 , \13403_13705_nG9bfc );
and \U$25937 ( \34576_34876 , \31334_31633 , \13771_14070_nG9bf9 );
or \U$25938 ( \34577_34877 , \34575_34875 , \34576_34876 );
xor \U$25939 ( \34578_34878 , \31333_31632 , \34577_34877 );
buf \U$25940 ( \34579_34879 , \34578_34878 );
buf \U$25942 ( \34580_34880 , \34579_34879 );
xor \U$25943 ( \34581_34881 , \34574_34874 , \34580_34880 );
buf \U$25944 ( \34582_34882 , \34581_34881 );
and \U$25945 ( \34583_34883 , \34470_34770 , \34476_34776 );
buf \U$25946 ( \34584_34884 , \34583_34883 );
xor \U$25947 ( \34585_34885 , \34582_34882 , \34584_34884 );
and \U$25948 ( \34586_34886 , \30670_29853 , \14682_14984_nG9bf6 );
and \U$25949 ( \34587_34887 , \29551_29850 , \15074_15373_nG9bf3 );
or \U$25950 ( \34588_34888 , \34586_34886 , \34587_34887 );
xor \U$25951 ( \34589_34889 , \29550_29849 , \34588_34888 );
buf \U$25952 ( \34590_34890 , \34589_34889 );
buf \U$25954 ( \34591_34891 , \34590_34890 );
xor \U$25955 ( \34592_34892 , \34585_34885 , \34591_34891 );
buf \U$25956 ( \34593_34893 , \34592_34892 );
and \U$25957 ( \34594_34894 , \25044_24792 , \18789_19091_nG9be4 );
and \U$25958 ( \34595_34895 , \24490_24789 , \19287_19586_nG9be1 );
or \U$25959 ( \34596_34896 , \34594_34894 , \34595_34895 );
xor \U$25960 ( \34597_34897 , \24489_24788 , \34596_34896 );
buf \U$25961 ( \34598_34898 , \34597_34897 );
buf \U$25963 ( \34599_34899 , \34598_34898 );
xor \U$25964 ( \34600_34900 , \34593_34893 , \34599_34899 );
and \U$25965 ( \34601_34901 , \23495_23201 , \20306_20608_nG9bde );
and \U$25966 ( \34602_34902 , \22899_23198 , \20787_21086_nG9bdb );
or \U$25967 ( \34603_34903 , \34601_34901 , \34602_34902 );
xor \U$25968 ( \34604_34904 , \22898_23197 , \34603_34903 );
buf \U$25969 ( \34605_34905 , \34604_34904 );
buf \U$25971 ( \34606_34906 , \34605_34905 );
xor \U$25972 ( \34607_34907 , \34600_34900 , \34606_34906 );
buf \U$25973 ( \34608_34908 , \34607_34907 );
xor \U$25974 ( \34609_34909 , \34569_34869 , \34608_34908 );
and \U$25975 ( \34610_34910 , \17437_17297 , \26585_26887_nG9bc6 );
and \U$25976 ( \34611_34911 , \16995_17294 , \27114_27416_nG9bc3 );
or \U$25977 ( \34612_34912 , \34610_34910 , \34611_34911 );
xor \U$25978 ( \34613_34913 , \16994_17293 , \34612_34912 );
buf \U$25979 ( \34614_34914 , \34613_34913 );
buf \U$25981 ( \34615_34915 , \34614_34914 );
xor \U$25982 ( \34616_34916 , \34609_34909 , \34615_34915 );
buf \U$25983 ( \34617_34917 , \34616_34916 );
xor \U$25984 ( \34618_34918 , \34564_34864 , \34617_34917 );
buf \U$25985 ( \34619_34919 , \34618_34918 );
xor \U$25986 ( \34620_34920 , \34553_34853 , \34619_34919 );
buf \U$25987 ( \34621_34921 , \34620_34920 );
and \U$25988 ( \34622_34922 , \34489_34789 , \34495_34795 );
and \U$25989 ( \34623_34923 , \34489_34789 , \34502_34802 );
and \U$25990 ( \34624_34924 , \34495_34795 , \34502_34802 );
or \U$25991 ( \34625_34925 , \34622_34922 , \34623_34923 , \34624_34924 );
buf \U$25992 ( \34626_34926 , \34625_34925 );
and \U$25993 ( \34627_34927 , \20353_20155 , \23394_23696_nG9bd2 );
and \U$25994 ( \34628_34928 , \19853_20152 , \23927_24226_nG9bcf );
or \U$25995 ( \34629_34929 , \34627_34927 , \34628_34928 );
xor \U$25996 ( \34630_34930 , \19852_20151 , \34629_34929 );
buf \U$25997 ( \34631_34931 , \34630_34930 );
buf \U$25999 ( \34632_34932 , \34631_34931 );
xor \U$26000 ( \34633_34933 , \34626_34926 , \34632_34932 );
and \U$26001 ( \34634_34934 , \18908_18702 , \24996_25298_nG9bcc );
and \U$26002 ( \34635_34935 , \18400_18699 , \25561_25860_nG9bc9 );
or \U$26003 ( \34636_34936 , \34634_34934 , \34635_34935 );
xor \U$26004 ( \34637_34937 , \18399_18698 , \34636_34936 );
buf \U$26005 ( \34638_34938 , \34637_34937 );
buf \U$26007 ( \34639_34939 , \34638_34938 );
xor \U$26008 ( \34640_34940 , \34633_34933 , \34639_34939 );
buf \U$26009 ( \34641_34941 , \34640_34940 );
and \U$26010 ( \34642_34942 , \10996_10421 , \33741_34041_nG9ba8 );
and \U$26011 ( \34643_34943 , \10119_10418 , \33994_34294_nG9ba5 );
or \U$26012 ( \34644_34944 , \34642_34942 , \34643_34943 );
xor \U$26013 ( \34645_34945 , \10118_10417 , \34644_34944 );
buf \U$26014 ( \34646_34946 , \34645_34945 );
buf \U$26016 ( \34647_34947 , \34646_34946 );
xor \U$26017 ( \34648_34948 , \34641_34941 , \34647_34947 );
and \U$26018 ( \34649_34949 , \10411_10707 , \34343_34643_nG9ba2 );
and \U$26019 ( \34650_34950 , \34272_34572 , \34276_34576 );
and \U$26020 ( \34651_34951 , \34276_34576 , \34331_34631 );
and \U$26021 ( \34652_34952 , \34272_34572 , \34331_34631 );
or \U$26022 ( \34653_34953 , \34650_34950 , \34651_34951 , \34652_34952 );
and \U$26023 ( \34654_34954 , \34204_34504 , \34208_34508 );
and \U$26024 ( \34655_34955 , \34208_34508 , \34220_34520 );
and \U$26025 ( \34656_34956 , \34204_34504 , \34220_34520 );
or \U$26026 ( \34657_34957 , \34654_34954 , \34655_34955 , \34656_34956 );
and \U$26027 ( \34658_34958 , \34226_34526 , \34240_34540 );
and \U$26028 ( \34659_34959 , \34240_34540 , \34265_34565 );
and \U$26029 ( \34660_34960 , \34226_34526 , \34265_34565 );
or \U$26030 ( \34661_34961 , \34658_34958 , \34659_34959 , \34660_34960 );
xor \U$26031 ( \34662_34962 , \34657_34957 , \34661_34961 );
and \U$26032 ( \34663_34963 , \34245_34545 , \34249_34549 );
and \U$26033 ( \34664_34964 , \34249_34549 , \34264_34564 );
and \U$26034 ( \34665_34965 , \34245_34545 , \34264_34564 );
or \U$26035 ( \34666_34966 , \34663_34963 , \34664_34964 , \34665_34965 );
and \U$26036 ( \34667_34967 , \34254_34554 , \34258_34558 );
and \U$26037 ( \34668_34968 , \34258_34558 , \34263_34563 );
and \U$26038 ( \34669_34969 , \34254_34554 , \34263_34563 );
or \U$26039 ( \34670_34970 , \34667_34967 , \34668_34968 , \34669_34969 );
and \U$26040 ( \34671_34971 , \34304_34604 , \34308_34608 );
and \U$26041 ( \34672_34972 , \34308_34608 , \34313_34613 );
and \U$26042 ( \34673_34973 , \34304_34604 , \34313_34613 );
or \U$26043 ( \34674_34974 , \34671_34971 , \34672_34972 , \34673_34973 );
xor \U$26044 ( \34675_34975 , \34670_34970 , \34674_34974 );
buf \U$26045 ( \34676_34976 , \34212_34512 );
xor \U$26046 ( \34677_34977 , \34675_34975 , \34676_34976 );
xor \U$26047 ( \34678_34978 , \34666_34966 , \34677_34977 );
and \U$26048 ( \34679_34979 , \34290_34590 , \34294_34594 );
and \U$26049 ( \34680_34980 , \34294_34594 , \34299_34599 );
and \U$26050 ( \34681_34981 , \34290_34590 , \34299_34599 );
or \U$26051 ( \34682_34982 , \34679_34979 , \34680_34980 , \34681_34981 );
and \U$26052 ( \34683_34983 , \34319_34619 , \34323_34623 );
and \U$26053 ( \34684_34984 , \34323_34623 , \34328_34628 );
and \U$26054 ( \34685_34985 , \34319_34619 , \34328_34628 );
or \U$26055 ( \34686_34986 , \34683_34983 , \34684_34984 , \34685_34985 );
xor \U$26056 ( \34687_34987 , \34682_34982 , \34686_34986 );
and \U$26057 ( \34688_34988 , \26527_26829 , \17791_18090 );
and \U$26058 ( \34689_34989 , \27011_27313 , \17353_17655 );
nor \U$26059 ( \34690_34990 , \34688_34988 , \34689_34989 );
xnor \U$26060 ( \34691_34991 , \34690_34990 , \17747_18046 );
and \U$26061 ( \34692_34992 , \21788_22090 , \22243_22542 );
and \U$26062 ( \34693_34993 , \22257_22556 , \21801_22103 );
nor \U$26063 ( \34694_34994 , \34692_34992 , \34693_34993 );
xnor \U$26064 ( \34695_34995 , \34694_34994 , \22249_22548 );
xor \U$26065 ( \34696_34996 , \34691_34991 , \34695_34995 );
and \U$26066 ( \34697_34997 , \20242_20544 , \23839_24138 );
and \U$26067 ( \34698_34998 , \20734_21033 , \23328_23630 );
nor \U$26068 ( \34699_34999 , \34697_34997 , \34698_34998 );
xnor \U$26069 ( \34700_35000 , \34699_34999 , \23845_24144 );
xor \U$26070 ( \34701_35001 , \34696_34996 , \34700_35000 );
xor \U$26071 ( \34702_35002 , \34687_34987 , \34701_35001 );
xor \U$26072 ( \34703_35003 , \34678_34978 , \34702_35002 );
xor \U$26073 ( \34704_35004 , \34662_34962 , \34703_35003 );
xor \U$26074 ( \34705_35005 , \34653_34953 , \34704_35004 );
and \U$26075 ( \34706_35006 , \34281_34581 , \34285_34585 );
and \U$26076 ( \34707_35007 , \34285_34585 , \34330_34630 );
and \U$26077 ( \34708_35008 , \34281_34581 , \34330_34630 );
or \U$26078 ( \34709_35009 , \34706_35006 , \34707_35007 , \34708_35008 );
and \U$26079 ( \34710_35010 , \34200_34500 , \34221_34521 );
and \U$26080 ( \34711_35011 , \34221_34521 , \34266_34566 );
and \U$26081 ( \34712_35012 , \34200_34500 , \34266_34566 );
or \U$26082 ( \34713_35013 , \34710_35010 , \34711_35011 , \34712_35012 );
xor \U$26083 ( \34714_35014 , \34709_35009 , \34713_35013 );
and \U$26084 ( \34715_35015 , \34300_34600 , \34314_34614 );
and \U$26085 ( \34716_35016 , \34314_34614 , \34329_34629 );
and \U$26086 ( \34717_35017 , \34300_34600 , \34329_34629 );
or \U$26087 ( \34718_35018 , \34715_35015 , \34716_35016 , \34717_35017 );
not \U$26088 ( \34719_35019 , \12481_12780 );
and \U$26089 ( \34720_35020 , \31752_32054 , \13755_14054 );
and \U$26090 ( \34721_35021 , \32495_32794 , \13390_13692 );
nor \U$26091 ( \34722_35022 , \34720_35020 , \34721_35021 );
xnor \U$26092 ( \34723_35023 , \34722_35022 , \13736_14035 );
xor \U$26093 ( \34724_35024 , \34719_35019 , \34723_35023 );
and \U$26094 ( \34725_35025 , \28232_28534 , \16333_16635 );
and \U$26095 ( \34726_35026 , \28782_29084 , \15999_16301 );
nor \U$26096 ( \34727_35027 , \34725_35025 , \34726_35026 );
xnor \U$26097 ( \34728_35028 , \34727_35027 , \16323_16625 );
xor \U$26098 ( \34729_35029 , \34724_35024 , \34728_35028 );
and \U$26099 ( \34730_35030 , \24970_25272 , \19235_19534 );
and \U$26100 ( \34731_35031 , \25516_25815 , \18743_19045 );
nor \U$26101 ( \34732_35032 , \34730_35030 , \34731_35031 );
xnor \U$26102 ( \34733_35033 , \34732_35032 , \19241_19540 );
and \U$26103 ( \34734_35034 , \15965_16267 , \28768_29070 );
and \U$26104 ( \34735_35035 , \16353_16655 , \28224_28526 );
nor \U$26105 ( \34736_35036 , \34734_35034 , \34735_35035 );
xnor \U$26106 ( \34737_35037 , \34736_35036 , \28774_29076 );
xor \U$26107 ( \34738_35038 , \34733_35033 , \34737_35037 );
and \U$26108 ( \34739_35039 , \14648_14950 , \30521_30823 );
and \U$26109 ( \34740_35040 , \15022_15321 , \29944_30246 );
nor \U$26110 ( \34741_35041 , \34739_35039 , \34740_35040 );
xnor \U$26111 ( \34742_35042 , \34741_35041 , \30511_30813 );
xor \U$26112 ( \34743_35043 , \34738_35038 , \34742_35042 );
xor \U$26113 ( \34744_35044 , \34729_35029 , \34743_35043 );
and \U$26114 ( \34745_35045 , \23315_23617 , \20706_21005 );
and \U$26115 ( \34746_35046 , \23900_24199 , \20255_20557 );
nor \U$26116 ( \34747_35047 , \34745_35045 , \34746_35046 );
xnor \U$26117 ( \34748_35048 , \34747_35047 , \20712_21011 );
and \U$26118 ( \34749_35049 , \13377_13679 , \32555_32854 );
and \U$26119 ( \34750_35050 , \13725_14024 , \31765_32067 );
nor \U$26120 ( \34751_35051 , \34749_35049 , \34750_35050 );
xnor \U$26121 ( \34752_35052 , \34751_35051 , \32506_32805 );
xor \U$26122 ( \34753_35053 , \34748_35048 , \34752_35052 );
and \U$26123 ( \34754_35054 , \12470_12769 , \32503_32802 );
xor \U$26124 ( \34755_35055 , \34753_35053 , \34754_35054 );
xor \U$26125 ( \34756_35056 , \34744_35044 , \34755_35055 );
xor \U$26126 ( \34757_35057 , \34718_35018 , \34756_35056 );
and \U$26127 ( \34758_35058 , \34230_34530 , \34234_34534 );
and \U$26128 ( \34759_35059 , \34234_34534 , \34239_34539 );
and \U$26129 ( \34760_35060 , \34230_34530 , \34239_34539 );
or \U$26130 ( \34761_35061 , \34758_35058 , \34759_35059 , \34760_35060 );
and \U$26131 ( \34762_35062 , \34213_34513 , \34217_34517 );
and \U$26132 ( \34763_35063 , \34217_34517 , \34219_34519 );
and \U$26133 ( \34764_35064 , \34213_34513 , \34219_34519 );
or \U$26134 ( \34765_35065 , \34762_35062 , \34763_35063 , \34764_35064 );
xor \U$26135 ( \34766_35066 , \34761_35061 , \34765_35065 );
and \U$26136 ( \34767_35067 , \29966_30268 , \15037_15336 );
and \U$26137 ( \34768_35068 , \30500_30802 , \14661_14963 );
nor \U$26138 ( \34769_35069 , \34767_35067 , \34768_35068 );
xnor \U$26139 ( \34770_35070 , \34769_35069 , \15043_15342 );
and \U$26140 ( \34771_35071 , \18730_19032 , \25527_25826 );
and \U$26141 ( \34772_35072 , \19259_19558 , \24962_25264 );
nor \U$26142 ( \34773_35073 , \34771_35071 , \34772_35072 );
xnor \U$26143 ( \34774_35074 , \34773_35073 , \25474_25773 );
xor \U$26144 ( \34775_35075 , \34770_35070 , \34774_35074 );
and \U$26145 ( \34776_35076 , \17325_17627 , \27095_27397 );
and \U$26146 ( \34777_35077 , \17736_18035 , \26505_26807 );
nor \U$26147 ( \34778_35078 , \34776_35076 , \34777_35077 );
xnor \U$26148 ( \34779_35079 , \34778_35078 , \26993_27295 );
xor \U$26149 ( \34780_35080 , \34775_35075 , \34779_35079 );
xor \U$26150 ( \34781_35081 , \34766_35066 , \34780_35080 );
xor \U$26151 ( \34782_35082 , \34757_35057 , \34781_35081 );
xor \U$26152 ( \34783_35083 , \34714_35014 , \34782_35082 );
xor \U$26153 ( \34784_35084 , \34705_35005 , \34783_35083 );
and \U$26154 ( \34785_35085 , \34196_34496 , \34267_34567 );
and \U$26155 ( \34786_35086 , \34267_34567 , \34332_34632 );
and \U$26156 ( \34787_35087 , \34196_34496 , \34332_34632 );
or \U$26157 ( \34788_35088 , \34785_35085 , \34786_35086 , \34787_35087 );
xor \U$26158 ( \34789_35089 , \34784_35084 , \34788_35088 );
and \U$26159 ( \34790_35090 , \34333_34633 , \34337_34637 );
and \U$26160 ( \34791_35091 , \34338_34638 , \34341_34641 );
or \U$26161 ( \34792_35092 , \34790_35090 , \34791_35091 );
xor \U$26162 ( \34793_35093 , \34789_35089 , \34792_35092 );
buf g9b9f_GF_PartitionCandidate( \34794_35094_nG9b9f , \34793_35093 );
and \U$26163 ( \34795_35095 , \10402_10704 , \34794_35094_nG9b9f );
or \U$26164 ( \34796_35096 , \34649_34949 , \34795_35095 );
xor \U$26165 ( \34797_35097 , \10399_10703 , \34796_35096 );
buf \U$26166 ( \34798_35098 , \34797_35097 );
buf \U$26168 ( \34799_35099 , \34798_35098 );
xor \U$26169 ( \34800_35100 , \34648_34948 , \34799_35099 );
buf \U$26170 ( \34801_35101 , \34800_35100 );
and \U$26171 ( \34802_35102 , \34465_34765 , \34518_34818 );
and \U$26172 ( \34803_35103 , \34465_34765 , \34524_34824 );
and \U$26173 ( \34804_35104 , \34518_34818 , \34524_34824 );
or \U$26174 ( \34805_35105 , \34802_35102 , \34803_35103 , \34804_35104 );
buf \U$26175 ( \34806_35106 , \34805_35105 );
xor \U$26176 ( \34807_35107 , \34801_35101 , \34806_35106 );
and \U$26177 ( \34808_35108 , \34169_34469 , \34175_34475 );
and \U$26178 ( \34809_35109 , \34169_34469 , \34182_34482 );
and \U$26179 ( \34810_35110 , \34175_34475 , \34182_34482 );
or \U$26180 ( \34811_35111 , \34808_35108 , \34809_35109 , \34810_35110 );
buf \U$26181 ( \34812_35112 , \34811_35111 );
and \U$26182 ( \34813_35113 , \34421_34721 , \34427_34727 );
and \U$26183 ( \34814_35114 , \34421_34721 , \34434_34734 );
and \U$26184 ( \34815_35115 , \34427_34727 , \34434_34734 );
or \U$26185 ( \34816_35116 , \34813_35113 , \34814_35114 , \34815_35115 );
buf \U$26186 ( \34817_35117 , \34816_35116 );
and \U$26187 ( \34818_35118 , \34478_34778 , \34480_34780 );
and \U$26188 ( \34819_35119 , \34478_34778 , \34487_34787 );
and \U$26189 ( \34820_35120 , \34480_34780 , \34487_34787 );
or \U$26190 ( \34821_35121 , \34818_35118 , \34819_35119 , \34820_35120 );
buf \U$26191 ( \34822_35122 , \34821_35121 );
and \U$26192 ( \34823_35123 , \28946_28118 , \16013_16315_nG9bf0 );
and \U$26193 ( \34824_35124 , \27816_28115 , \16378_16680_nG9bed );
or \U$26194 ( \34825_35125 , \34823_35123 , \34824_35124 );
xor \U$26195 ( \34826_35126 , \27815_28114 , \34825_35125 );
buf \U$26196 ( \34827_35127 , \34826_35126 );
buf \U$26198 ( \34828_35128 , \34827_35127 );
xor \U$26199 ( \34829_35129 , \34822_35122 , \34828_35128 );
and \U$26200 ( \34830_35130 , \27141_26431 , \17363_17665_nG9bea );
and \U$26201 ( \34831_35131 , \26129_26428 , \17808_18107_nG9be7 );
or \U$26202 ( \34832_35132 , \34830_35130 , \34831_35131 );
xor \U$26203 ( \34833_35133 , \26128_26427 , \34832_35132 );
buf \U$26204 ( \34834_35134 , \34833_35133 );
buf \U$26206 ( \34835_35135 , \34834_35134 );
xor \U$26207 ( \34836_35136 , \34829_35129 , \34835_35135 );
buf \U$26208 ( \34837_35137 , \34836_35136 );
xor \U$26209 ( \34838_35138 , \34817_35117 , \34837_35137 );
and \U$26210 ( \34839_35139 , \21908_21658 , \21827_22129_nG9bd8 );
and \U$26211 ( \34840_35140 , \21356_21655 , \22330_22629_nG9bd5 );
or \U$26212 ( \34841_35141 , \34839_35139 , \34840_35140 );
xor \U$26213 ( \34842_35142 , \21355_21654 , \34841_35141 );
buf \U$26214 ( \34843_35143 , \34842_35142 );
buf \U$26216 ( \34844_35144 , \34843_35143 );
xor \U$26217 ( \34845_35145 , \34838_35138 , \34844_35144 );
buf \U$26218 ( \34846_35146 , \34845_35145 );
xor \U$26219 ( \34847_35147 , \34812_35112 , \34846_35146 );
and \U$26220 ( \34848_35148 , \13431_13370 , \31877_32179_nG9bb4 );
and \U$26221 ( \34849_35149 , \13068_13367 , \32589_32888_nG9bb1 );
or \U$26222 ( \34850_35150 , \34848_35148 , \34849_35149 );
xor \U$26223 ( \34851_35151 , \13067_13366 , \34850_35150 );
buf \U$26224 ( \34852_35152 , \34851_35151 );
buf \U$26226 ( \34853_35153 , \34852_35152 );
xor \U$26227 ( \34854_35154 , \34847_35147 , \34853_35153 );
buf \U$26228 ( \34855_35155 , \34854_35154 );
xor \U$26229 ( \34856_35156 , \34807_35107 , \34855_35155 );
buf \U$26230 ( \34857_35157 , \34856_35156 );
xor \U$26231 ( \34858_35158 , \34621_34921 , \34857_35157 );
and \U$26232 ( \34859_35159 , \34184_34484 , \34190_34490 );
and \U$26233 ( \34860_35160 , \34184_34484 , \34348_34648 );
and \U$26234 ( \34861_35161 , \34190_34490 , \34348_34648 );
or \U$26235 ( \34862_35162 , \34859_35159 , \34860_35160 , \34861_35161 );
buf \U$26236 ( \34863_35163 , \34862_35162 );
and \U$26237 ( \34864_35164 , \34361_34661 , \34367_34667 );
and \U$26238 ( \34865_35165 , \34361_34661 , \34374_34674 );
and \U$26239 ( \34866_35166 , \34367_34667 , \34374_34674 );
or \U$26240 ( \34867_35167 , \34864_35164 , \34865_35165 , \34866_35166 );
buf \U$26241 ( \34868_35168 , \34867_35167 );
xor \U$26242 ( \34869_35169 , \34863_35163 , \34868_35168 );
and \U$26243 ( \34870_35170 , \16405_15940 , \28300_28602_nG9bc0 );
and \U$26244 ( \34871_35171 , \15638_15937 , \28877_29179_nG9bbd );
or \U$26245 ( \34872_35172 , \34870_35170 , \34871_35171 );
xor \U$26246 ( \34873_35173 , \15637_15936 , \34872_35172 );
buf \U$26247 ( \34874_35174 , \34873_35173 );
buf \U$26249 ( \34875_35175 , \34874_35174 );
and \U$26250 ( \34876_35176 , \14710_14631 , \30064_30366_nG9bba );
and \U$26251 ( \34877_35177 , \14329_14628 , \30638_30940_nG9bb7 );
or \U$26252 ( \34878_35178 , \34876_35176 , \34877_35177 );
xor \U$26253 ( \34879_35179 , \14328_14627 , \34878_35178 );
buf \U$26254 ( \34880_35180 , \34879_35179 );
buf \U$26256 ( \34881_35181 , \34880_35180 );
xor \U$26257 ( \34882_35182 , \34875_35175 , \34881_35181 );
and \U$26258 ( \34883_35183 , \12183_12157 , \32881_33181_nG9bae );
and \U$26259 ( \34884_35184 , \11855_12154 , \33313_33613_nG9bab );
or \U$26260 ( \34885_35185 , \34883_35183 , \34884_35184 );
xor \U$26261 ( \34886_35186 , \11854_12153 , \34885_35185 );
buf \U$26262 ( \34887_35187 , \34886_35186 );
buf \U$26264 ( \34888_35188 , \34887_35187 );
xor \U$26265 ( \34889_35189 , \34882_35182 , \34888_35188 );
buf \U$26266 ( \34890_35190 , \34889_35189 );
xor \U$26267 ( \34891_35191 , \34869_35169 , \34890_35190 );
buf \U$26268 ( \34892_35192 , \34891_35191 );
xor \U$26269 ( \34893_35193 , \34858_35158 , \34892_35192 );
buf \U$26270 ( \34894_35194 , \34893_35193 );
and \U$26271 ( \34895_35195 , \34164_34464 , \34378_34678 );
and \U$26272 ( \34896_35196 , \34164_34464 , \34384_34684 );
and \U$26273 ( \34897_35197 , \34378_34678 , \34384_34684 );
or \U$26274 ( \34898_35198 , \34895_35195 , \34896_35196 , \34897_35197 );
buf \U$26275 ( \34899_35199 , \34898_35198 );
xor \U$26276 ( \34900_35200 , \34894_35194 , \34899_35199 );
and \U$26277 ( \34901_35201 , \34410_34710 , \34415_34715 );
and \U$26278 ( \34902_35202 , \34410_34710 , \34526_34826 );
and \U$26279 ( \34903_35203 , \34415_34715 , \34526_34826 );
or \U$26280 ( \34904_35204 , \34901_35201 , \34902_35202 , \34903_35203 );
buf \U$26281 ( \34905_35205 , \34904_35204 );
xor \U$26282 ( \34906_35206 , \34900_35200 , \34905_35205 );
and \U$26283 ( \34907_35207 , \34542_34842 , \34906_35206 );
and \U$26285 ( \34908_35208 , \34536_34836 , \34541_34841 );
or \U$26287 ( \34909_35209 , 1'b0 , \34908_35208 , 1'b0 );
xor \U$26288 ( \34910_35210 , \34907_35207 , \34909_35209 );
and \U$26290 ( \34911_35211 , \34530_34830 , \34535_34835 );
and \U$26291 ( \34912_35212 , \34532_34832 , \34535_34835 );
or \U$26292 ( \34913_35213 , 1'b0 , \34911_35211 , \34912_35212 );
xor \U$26293 ( \34914_35214 , \34910_35210 , \34913_35213 );
xor \U$26300 ( \34915_35215 , \34914_35214 , 1'b0 );
and \U$26301 ( \34916_35216 , \34894_35194 , \34899_35199 );
and \U$26302 ( \34917_35217 , \34894_35194 , \34905_35205 );
and \U$26303 ( \34918_35218 , \34899_35199 , \34905_35205 );
or \U$26304 ( \34919_35219 , \34916_35216 , \34917_35217 , \34918_35218 );
xor \U$26305 ( \34920_35220 , \34915_35215 , \34919_35219 );
and \U$26306 ( \34921_35221 , \34621_34921 , \34857_35157 );
and \U$26307 ( \34922_35222 , \34621_34921 , \34892_35192 );
and \U$26308 ( \34923_35223 , \34857_35157 , \34892_35192 );
or \U$26309 ( \34924_35224 , \34921_35221 , \34922_35222 , \34923_35223 );
buf \U$26310 ( \34925_35225 , \34924_35224 );
and \U$26311 ( \34926_35226 , \34641_34941 , \34647_34947 );
and \U$26312 ( \34927_35227 , \34641_34941 , \34799_35099 );
and \U$26313 ( \34928_35228 , \34647_34947 , \34799_35099 );
or \U$26314 ( \34929_35229 , \34926_35226 , \34927_35227 , \34928_35228 );
buf \U$26315 ( \34930_35230 , \34929_35229 );
and \U$26316 ( \34931_35231 , \34558_34858 , \34563_34863 );
and \U$26317 ( \34932_35232 , \34558_34858 , \34617_34917 );
and \U$26318 ( \34933_35233 , \34563_34863 , \34617_34917 );
or \U$26319 ( \34934_35234 , \34931_35231 , \34932_35232 , \34933_35233 );
buf \U$26320 ( \34935_35235 , \34934_35234 );
xor \U$26321 ( \34936_35236 , \34930_35230 , \34935_35235 );
and \U$26322 ( \34937_35237 , \34569_34869 , \34608_34908 );
and \U$26323 ( \34938_35238 , \34569_34869 , \34615_34915 );
and \U$26324 ( \34939_35239 , \34608_34908 , \34615_34915 );
or \U$26325 ( \34940_35240 , \34937_35237 , \34938_35238 , \34939_35239 );
buf \U$26326 ( \34941_35241 , \34940_35240 );
and \U$26327 ( \34942_35242 , \34626_34926 , \34632_34932 );
and \U$26328 ( \34943_35243 , \34626_34926 , \34639_34939 );
and \U$26329 ( \34944_35244 , \34632_34932 , \34639_34939 );
or \U$26330 ( \34945_35245 , \34942_35242 , \34943_35243 , \34944_35244 );
buf \U$26331 ( \34946_35246 , \34945_35245 );
xor \U$26332 ( \34947_35247 , \34941_35241 , \34946_35246 );
and \U$26333 ( \34948_35248 , \34593_34893 , \34599_34899 );
and \U$26334 ( \34949_35249 , \34593_34893 , \34606_34906 );
and \U$26335 ( \34950_35250 , \34599_34899 , \34606_34906 );
or \U$26336 ( \34951_35251 , \34948_35248 , \34949_35249 , \34950_35250 );
buf \U$26337 ( \34952_35252 , \34951_35251 );
and \U$26338 ( \34953_35253 , \34582_34882 , \34584_34884 );
and \U$26339 ( \34954_35254 , \34582_34882 , \34591_34891 );
and \U$26340 ( \34955_35255 , \34584_34884 , \34591_34891 );
or \U$26341 ( \34956_35256 , \34953_35253 , \34954_35254 , \34955_35255 );
buf \U$26342 ( \34957_35257 , \34956_35256 );
and \U$26343 ( \34958_35258 , \28946_28118 , \16378_16680_nG9bed );
and \U$26344 ( \34959_35259 , \27816_28115 , \17363_17665_nG9bea );
or \U$26345 ( \34960_35260 , \34958_35258 , \34959_35259 );
xor \U$26346 ( \34961_35261 , \27815_28114 , \34960_35260 );
buf \U$26347 ( \34962_35262 , \34961_35261 );
buf \U$26349 ( \34963_35263 , \34962_35262 );
xor \U$26350 ( \34964_35264 , \34957_35257 , \34963_35263 );
and \U$26351 ( \34965_35265 , \27141_26431 , \17808_18107_nG9be7 );
and \U$26352 ( \34966_35266 , \26129_26428 , \18789_19091_nG9be4 );
or \U$26353 ( \34967_35267 , \34965_35265 , \34966_35266 );
xor \U$26354 ( \34968_35268 , \26128_26427 , \34967_35267 );
buf \U$26355 ( \34969_35269 , \34968_35268 );
buf \U$26357 ( \34970_35270 , \34969_35269 );
xor \U$26358 ( \34971_35271 , \34964_35264 , \34970_35270 );
buf \U$26359 ( \34972_35272 , \34971_35271 );
xor \U$26360 ( \34973_35273 , \34952_35252 , \34972_35272 );
and \U$26361 ( \34974_35274 , \18908_18702 , \25561_25860_nG9bc9 );
and \U$26362 ( \34975_35275 , \18400_18699 , \26585_26887_nG9bc6 );
or \U$26363 ( \34976_35276 , \34974_35274 , \34975_35275 );
xor \U$26364 ( \34977_35277 , \18399_18698 , \34976_35276 );
buf \U$26365 ( \34978_35278 , \34977_35277 );
buf \U$26367 ( \34979_35279 , \34978_35278 );
xor \U$26368 ( \34980_35280 , \34973_35273 , \34979_35279 );
buf \U$26369 ( \34981_35281 , \34980_35280 );
xor \U$26370 ( \34982_35282 , \34947_35247 , \34981_35281 );
buf \U$26371 ( \34983_35283 , \34982_35282 );
xor \U$26372 ( \34984_35284 , \34936_35236 , \34983_35283 );
buf \U$26373 ( \34985_35285 , \34984_35284 );
and \U$26374 ( \34986_35286 , \34801_35101 , \34806_35106 );
and \U$26375 ( \34987_35287 , \34801_35101 , \34855_35155 );
and \U$26376 ( \34988_35288 , \34806_35106 , \34855_35155 );
or \U$26377 ( \34989_35289 , \34986_35286 , \34987_35287 , \34988_35288 );
buf \U$26378 ( \34990_35290 , \34989_35289 );
xor \U$26379 ( \34991_35291 , \34985_35285 , \34990_35290 );
and \U$26380 ( \34992_35292 , \34547_34847 , \34552_34852 );
and \U$26381 ( \34993_35293 , \34547_34847 , \34619_34919 );
and \U$26382 ( \34994_35294 , \34552_34852 , \34619_34919 );
or \U$26383 ( \34995_35295 , \34992_35292 , \34993_35293 , \34994_35294 );
buf \U$26384 ( \34996_35296 , \34995_35295 );
xor \U$26385 ( \34997_35297 , \34991_35291 , \34996_35296 );
buf \U$26386 ( \34998_35298 , \34997_35297 );
xor \U$26387 ( \34999_35299 , \34925_35225 , \34998_35298 );
and \U$26388 ( \35000_35300 , \34822_35122 , \34828_35128 );
and \U$26389 ( \35001_35301 , \34822_35122 , \34835_35135 );
and \U$26390 ( \35002_35302 , \34828_35128 , \34835_35135 );
or \U$26391 ( \35003_35303 , \35000_35300 , \35001_35301 , \35002_35302 );
buf \U$26392 ( \35004_35304 , \35003_35303 );
and \U$26393 ( \35005_35305 , \21908_21658 , \22330_22629_nG9bd5 );
and \U$26394 ( \35006_35306 , \21356_21655 , \23394_23696_nG9bd2 );
or \U$26395 ( \35007_35307 , \35005_35305 , \35006_35306 );
xor \U$26396 ( \35008_35308 , \21355_21654 , \35007_35307 );
buf \U$26397 ( \35009_35309 , \35008_35308 );
buf \U$26399 ( \35010_35310 , \35009_35309 );
xor \U$26400 ( \35011_35311 , \35004_35304 , \35010_35310 );
and \U$26401 ( \35012_35312 , \20353_20155 , \23927_24226_nG9bcf );
and \U$26402 ( \35013_35313 , \19853_20152 , \24996_25298_nG9bcc );
or \U$26403 ( \35014_35314 , \35012_35312 , \35013_35313 );
xor \U$26404 ( \35015_35315 , \19852_20151 , \35014_35314 );
buf \U$26405 ( \35016_35316 , \35015_35315 );
buf \U$26407 ( \35017_35317 , \35016_35316 );
xor \U$26408 ( \35018_35318 , \35011_35311 , \35017_35317 );
buf \U$26409 ( \35019_35319 , \35018_35318 );
and \U$26410 ( \35020_35320 , \13431_13370 , \32589_32888_nG9bb1 );
and \U$26411 ( \35021_35321 , \13068_13367 , \32881_33181_nG9bae );
or \U$26412 ( \35022_35322 , \35020_35320 , \35021_35321 );
xor \U$26413 ( \35023_35323 , \13067_13366 , \35022_35322 );
buf \U$26414 ( \35024_35324 , \35023_35323 );
buf \U$26416 ( \35025_35325 , \35024_35324 );
xor \U$26417 ( \35026_35326 , \35019_35319 , \35025_35325 );
and \U$26418 ( \35027_35327 , \10996_10421 , \33994_34294_nG9ba5 );
and \U$26419 ( \35028_35328 , \10119_10418 , \34343_34643_nG9ba2 );
or \U$26420 ( \35029_35329 , \35027_35327 , \35028_35328 );
xor \U$26421 ( \35030_35330 , \10118_10417 , \35029_35329 );
buf \U$26422 ( \35031_35331 , \35030_35330 );
buf \U$26424 ( \35032_35332 , \35031_35331 );
xor \U$26425 ( \35033_35333 , \35026_35326 , \35032_35332 );
buf \U$26426 ( \35034_35334 , \35033_35333 );
and \U$26427 ( \35035_35335 , \34812_35112 , \34846_35146 );
and \U$26428 ( \35036_35336 , \34812_35112 , \34853_35153 );
and \U$26429 ( \35037_35337 , \34846_35146 , \34853_35153 );
or \U$26430 ( \35038_35338 , \35035_35335 , \35036_35336 , \35037_35337 );
buf \U$26431 ( \35039_35339 , \35038_35338 );
xor \U$26432 ( \35040_35340 , \35034_35334 , \35039_35339 );
and \U$26433 ( \35041_35341 , \34875_35175 , \34881_35181 );
and \U$26434 ( \35042_35342 , \34875_35175 , \34888_35188 );
and \U$26435 ( \35043_35343 , \34881_35181 , \34888_35188 );
or \U$26436 ( \35044_35344 , \35041_35341 , \35042_35342 , \35043_35343 );
buf \U$26437 ( \35045_35345 , \35044_35344 );
xor \U$26438 ( \35046_35346 , \35040_35340 , \35045_35345 );
buf \U$26439 ( \35047_35347 , \35046_35346 );
and \U$26440 ( \35048_35348 , \34863_35163 , \34868_35168 );
and \U$26441 ( \35049_35349 , \34863_35163 , \34890_35190 );
and \U$26442 ( \35050_35350 , \34868_35168 , \34890_35190 );
or \U$26443 ( \35051_35351 , \35048_35348 , \35049_35349 , \35050_35350 );
buf \U$26444 ( \35052_35352 , \35051_35351 );
xor \U$26445 ( \35053_35353 , \35047_35347 , \35052_35352 );
and \U$26446 ( \35054_35354 , \16405_15940 , \28877_29179_nG9bbd );
and \U$26447 ( \35055_35355 , \15638_15937 , \30064_30366_nG9bba );
or \U$26448 ( \35056_35356 , \35054_35354 , \35055_35355 );
xor \U$26449 ( \35057_35357 , \15637_15936 , \35056_35356 );
buf \U$26450 ( \35058_35358 , \35057_35357 );
buf \U$26452 ( \35059_35359 , \35058_35358 );
and \U$26453 ( \35060_35360 , \14710_14631 , \30638_30940_nG9bb7 );
and \U$26454 ( \35061_35361 , \14329_14628 , \31877_32179_nG9bb4 );
or \U$26455 ( \35062_35362 , \35060_35360 , \35061_35361 );
xor \U$26456 ( \35063_35363 , \14328_14627 , \35062_35362 );
buf \U$26457 ( \35064_35364 , \35063_35363 );
buf \U$26459 ( \35065_35365 , \35064_35364 );
xor \U$26460 ( \35066_35366 , \35059_35359 , \35065_35365 );
and \U$26461 ( \35067_35367 , \12183_12157 , \33313_33613_nG9bab );
and \U$26462 ( \35068_35368 , \11855_12154 , \33741_34041_nG9ba8 );
or \U$26463 ( \35069_35369 , \35067_35367 , \35068_35368 );
xor \U$26464 ( \35070_35370 , \11854_12153 , \35069_35369 );
buf \U$26465 ( \35071_35371 , \35070_35370 );
buf \U$26467 ( \35072_35372 , \35071_35371 );
xor \U$26468 ( \35073_35373 , \35066_35366 , \35072_35372 );
buf \U$26469 ( \35074_35374 , \35073_35373 );
and \U$26470 ( \35075_35375 , \34817_35117 , \34837_35137 );
and \U$26471 ( \35076_35376 , \34817_35117 , \34844_35144 );
and \U$26472 ( \35077_35377 , \34837_35137 , \34844_35144 );
or \U$26473 ( \35078_35378 , \35075_35375 , \35076_35376 , \35077_35377 );
buf \U$26474 ( \35079_35379 , \35078_35378 );
and \U$26476 ( \35080_35380 , \32617_32916 , \13403_13705_nG9bfc );
or \U$26477 ( \35081_35381 , 1'b0 , \35080_35380 );
xor \U$26478 ( \35082_35382 , 1'b0 , \35081_35381 );
buf \U$26479 ( \35083_35383 , \35082_35382 );
buf \U$26481 ( \35084_35384 , \35083_35383 );
and \U$26482 ( \35085_35385 , \31989_31636 , \13771_14070_nG9bf9 );
and \U$26483 ( \35086_35386 , \31334_31633 , \14682_14984_nG9bf6 );
or \U$26484 ( \35087_35387 , \35085_35385 , \35086_35386 );
xor \U$26485 ( \35088_35388 , \31333_31632 , \35087_35387 );
buf \U$26486 ( \35089_35389 , \35088_35388 );
buf \U$26488 ( \35090_35390 , \35089_35389 );
xor \U$26489 ( \35091_35391 , \35084_35384 , \35090_35390 );
buf \U$26490 ( \35092_35392 , \35091_35391 );
and \U$26491 ( \35093_35393 , \34574_34874 , \34580_34880 );
buf \U$26492 ( \35094_35394 , \35093_35393 );
xor \U$26493 ( \35095_35395 , \35092_35392 , \35094_35394 );
and \U$26494 ( \35096_35396 , \30670_29853 , \15074_15373_nG9bf3 );
and \U$26495 ( \35097_35397 , \29551_29850 , \16013_16315_nG9bf0 );
or \U$26496 ( \35098_35398 , \35096_35396 , \35097_35397 );
xor \U$26497 ( \35099_35399 , \29550_29849 , \35098_35398 );
buf \U$26498 ( \35100_35400 , \35099_35399 );
buf \U$26500 ( \35101_35401 , \35100_35400 );
xor \U$26501 ( \35102_35402 , \35095_35395 , \35101_35401 );
buf \U$26502 ( \35103_35403 , \35102_35402 );
and \U$26503 ( \35104_35404 , \25044_24792 , \19287_19586_nG9be1 );
and \U$26504 ( \35105_35405 , \24490_24789 , \20306_20608_nG9bde );
or \U$26505 ( \35106_35406 , \35104_35404 , \35105_35405 );
xor \U$26506 ( \35107_35407 , \24489_24788 , \35106_35406 );
buf \U$26507 ( \35108_35408 , \35107_35407 );
buf \U$26509 ( \35109_35409 , \35108_35408 );
xor \U$26510 ( \35110_35410 , \35103_35403 , \35109_35409 );
and \U$26511 ( \35111_35411 , \23495_23201 , \20787_21086_nG9bdb );
and \U$26512 ( \35112_35412 , \22899_23198 , \21827_22129_nG9bd8 );
or \U$26513 ( \35113_35413 , \35111_35411 , \35112_35412 );
xor \U$26514 ( \35114_35414 , \22898_23197 , \35113_35413 );
buf \U$26515 ( \35115_35415 , \35114_35414 );
buf \U$26517 ( \35116_35416 , \35115_35415 );
xor \U$26518 ( \35117_35417 , \35110_35410 , \35116_35416 );
buf \U$26519 ( \35118_35418 , \35117_35417 );
xor \U$26520 ( \35119_35419 , \35079_35379 , \35118_35418 );
and \U$26521 ( \35120_35420 , \17437_17297 , \27114_27416_nG9bc3 );
and \U$26522 ( \35121_35421 , \16995_17294 , \28300_28602_nG9bc0 );
or \U$26523 ( \35122_35422 , \35120_35420 , \35121_35421 );
xor \U$26524 ( \35123_35423 , \16994_17293 , \35122_35422 );
buf \U$26525 ( \35124_35424 , \35123_35423 );
buf \U$26527 ( \35125_35425 , \35124_35424 );
xor \U$26528 ( \35126_35426 , \35119_35419 , \35125_35425 );
buf \U$26529 ( \35127_35427 , \35126_35426 );
xor \U$26530 ( \35128_35428 , \35074_35374 , \35127_35427 );
and \U$26531 ( \35129_35429 , \10411_10707 , \34794_35094_nG9b9f );
and \U$26532 ( \35130_35430 , \34657_34957 , \34661_34961 );
and \U$26533 ( \35131_35431 , \34661_34961 , \34703_35003 );
and \U$26534 ( \35132_35432 , \34657_34957 , \34703_35003 );
or \U$26535 ( \35133_35433 , \35130_35430 , \35131_35431 , \35132_35432 );
and \U$26536 ( \35134_35434 , \34709_35009 , \34713_35013 );
and \U$26537 ( \35135_35435 , \34713_35013 , \34782_35082 );
and \U$26538 ( \35136_35436 , \34709_35009 , \34782_35082 );
or \U$26539 ( \35137_35437 , \35134_35434 , \35135_35435 , \35136_35436 );
xor \U$26540 ( \35138_35438 , \35133_35433 , \35137_35437 );
and \U$26541 ( \35139_35439 , \34718_35018 , \34756_35056 );
and \U$26542 ( \35140_35440 , \34756_35056 , \34781_35081 );
and \U$26543 ( \35141_35441 , \34718_35018 , \34781_35081 );
or \U$26544 ( \35142_35442 , \35139_35439 , \35140_35440 , \35141_35441 );
and \U$26545 ( \35143_35443 , \34729_35029 , \34743_35043 );
and \U$26546 ( \35144_35444 , \34743_35043 , \34755_35055 );
and \U$26547 ( \35145_35445 , \34729_35029 , \34755_35055 );
or \U$26548 ( \35146_35446 , \35143_35443 , \35144_35444 , \35145_35445 );
and \U$26549 ( \35147_35447 , \34761_35061 , \34765_35065 );
and \U$26550 ( \35148_35448 , \34765_35065 , \34780_35080 );
and \U$26551 ( \35149_35449 , \34761_35061 , \34780_35080 );
or \U$26552 ( \35150_35450 , \35147_35447 , \35148_35448 , \35149_35449 );
xor \U$26553 ( \35151_35451 , \35146_35446 , \35150_35450 );
and \U$26554 ( \35152_35452 , \34748_35048 , \34752_35052 );
and \U$26555 ( \35153_35453 , \34752_35052 , \34754_35054 );
and \U$26556 ( \35154_35454 , \34748_35048 , \34754_35054 );
or \U$26557 ( \35155_35455 , \35152_35452 , \35153_35453 , \35154_35454 );
and \U$26558 ( \35156_35456 , \28782_29084 , \16333_16635 );
and \U$26559 ( \35157_35457 , \29966_30268 , \15999_16301 );
nor \U$26560 ( \35158_35458 , \35156_35456 , \35157_35457 );
xnor \U$26561 ( \35159_35459 , \35158_35458 , \16323_16625 );
and \U$26562 ( \35160_35460 , \13725_14024 , \32555_32854 );
and \U$26563 ( \35161_35461 , \14648_14950 , \31765_32067 );
nor \U$26564 ( \35162_35462 , \35160_35460 , \35161_35461 );
xnor \U$26565 ( \35163_35463 , \35162_35462 , \32506_32805 );
xor \U$26566 ( \35164_35464 , \35159_35459 , \35163_35463 );
and \U$26567 ( \35165_35465 , \13377_13679 , \32503_32802 );
xor \U$26568 ( \35166_35466 , \35164_35464 , \35165_35465 );
xor \U$26569 ( \35167_35467 , \35155_35455 , \35166_35466 );
and \U$26570 ( \35168_35468 , \27011_27313 , \17791_18090 );
and \U$26571 ( \35169_35469 , \28232_28534 , \17353_17655 );
nor \U$26572 ( \35170_35470 , \35168_35468 , \35169_35469 );
xnor \U$26573 ( \35171_35471 , \35170_35470 , \17747_18046 );
and \U$26574 ( \35172_35472 , \20734_21033 , \23839_24138 );
and \U$26575 ( \35173_35473 , \21788_22090 , \23328_23630 );
nor \U$26576 ( \35174_35474 , \35172_35472 , \35173_35473 );
xnor \U$26577 ( \35175_35475 , \35174_35474 , \23845_24144 );
xor \U$26578 ( \35176_35476 , \35171_35471 , \35175_35475 );
and \U$26579 ( \35177_35477 , \19259_19558 , \25527_25826 );
and \U$26580 ( \35178_35478 , \20242_20544 , \24962_25264 );
nor \U$26581 ( \35179_35479 , \35177_35477 , \35178_35478 );
xnor \U$26582 ( \35180_35480 , \35179_35479 , \25474_25773 );
xor \U$26583 ( \35181_35481 , \35176_35476 , \35180_35480 );
xor \U$26584 ( \35182_35482 , \35167_35467 , \35181_35481 );
xor \U$26585 ( \35183_35483 , \35151_35451 , \35182_35482 );
xor \U$26586 ( \35184_35484 , \35142_35442 , \35183_35483 );
and \U$26587 ( \35185_35485 , \34666_34966 , \34677_34977 );
and \U$26588 ( \35186_35486 , \34677_34977 , \34702_35002 );
and \U$26589 ( \35187_35487 , \34666_34966 , \34702_35002 );
or \U$26590 ( \35188_35488 , \35185_35485 , \35186_35486 , \35187_35487 );
and \U$26591 ( \35189_35489 , \32495_32794 , \13755_14054 );
not \U$26592 ( \35190_35490 , \35189_35489 );
xnor \U$26593 ( \35191_35491 , \35190_35490 , \13736_14035 );
and \U$26594 ( \35192_35492 , \23900_24199 , \20706_21005 );
and \U$26595 ( \35193_35493 , \24970_25272 , \20255_20557 );
nor \U$26596 ( \35194_35494 , \35192_35492 , \35193_35493 );
xnor \U$26597 ( \35195_35495 , \35194_35494 , \20712_21011 );
xor \U$26598 ( \35196_35496 , \35191_35491 , \35195_35495 );
and \U$26599 ( \35197_35497 , \15022_15321 , \30521_30823 );
and \U$26600 ( \35198_35498 , \15965_16267 , \29944_30246 );
nor \U$26601 ( \35199_35499 , \35197_35497 , \35198_35498 );
xnor \U$26602 ( \35200_35500 , \35199_35499 , \30511_30813 );
xor \U$26603 ( \35201_35501 , \35196_35496 , \35200_35500 );
and \U$26604 ( \35202_35502 , \25516_25815 , \19235_19534 );
and \U$26605 ( \35203_35503 , \26527_26829 , \18743_19045 );
nor \U$26606 ( \35204_35504 , \35202_35502 , \35203_35503 );
xnor \U$26607 ( \35205_35505 , \35204_35504 , \19241_19540 );
and \U$26608 ( \35206_35506 , \17736_18035 , \27095_27397 );
and \U$26609 ( \35207_35507 , \18730_19032 , \26505_26807 );
nor \U$26610 ( \35208_35508 , \35206_35506 , \35207_35507 );
xnor \U$26611 ( \35209_35509 , \35208_35508 , \26993_27295 );
xor \U$26612 ( \35210_35510 , \35205_35505 , \35209_35509 );
and \U$26613 ( \35211_35511 , \16353_16655 , \28768_29070 );
and \U$26614 ( \35212_35512 , \17325_17627 , \28224_28526 );
nor \U$26615 ( \35213_35513 , \35211_35511 , \35212_35512 );
xnor \U$26616 ( \35214_35514 , \35213_35513 , \28774_29076 );
xor \U$26617 ( \35215_35515 , \35210_35510 , \35214_35514 );
xor \U$26618 ( \35216_35516 , \35201_35501 , \35215_35515 );
and \U$26619 ( \35217_35517 , \34733_35033 , \34737_35037 );
and \U$26620 ( \35218_35518 , \34737_35037 , \34742_35042 );
and \U$26621 ( \35219_35519 , \34733_35033 , \34742_35042 );
or \U$26622 ( \35220_35520 , \35217_35517 , \35218_35518 , \35219_35519 );
and \U$26623 ( \35221_35521 , \30500_30802 , \15037_15336 );
and \U$26624 ( \35222_35522 , \31752_32054 , \14661_14963 );
nor \U$26625 ( \35223_35523 , \35221_35521 , \35222_35522 );
xnor \U$26626 ( \35224_35524 , \35223_35523 , \15043_15342 );
not \U$26627 ( \35225_35525 , \35224_35524 );
xor \U$26628 ( \35226_35526 , \35220_35520 , \35225_35525 );
and \U$26629 ( \35227_35527 , \22257_22556 , \22243_22542 );
and \U$26630 ( \35228_35528 , \23315_23617 , \21801_22103 );
nor \U$26631 ( \35229_35529 , \35227_35527 , \35228_35528 );
xnor \U$26632 ( \35230_35530 , \35229_35529 , \22249_22548 );
xor \U$26633 ( \35231_35531 , \35226_35526 , \35230_35530 );
xor \U$26634 ( \35232_35532 , \35216_35516 , \35231_35531 );
xor \U$26635 ( \35233_35533 , \35188_35488 , \35232_35532 );
and \U$26636 ( \35234_35534 , \34670_34970 , \34674_34974 );
and \U$26637 ( \35235_35535 , \34674_34974 , \34676_34976 );
and \U$26638 ( \35236_35536 , \34670_34970 , \34676_34976 );
or \U$26639 ( \35237_35537 , \35234_35534 , \35235_35535 , \35236_35536 );
and \U$26640 ( \35238_35538 , \34682_34982 , \34686_34986 );
and \U$26641 ( \35239_35539 , \34686_34986 , \34701_35001 );
and \U$26642 ( \35240_35540 , \34682_34982 , \34701_35001 );
or \U$26643 ( \35241_35541 , \35238_35538 , \35239_35539 , \35240_35540 );
xor \U$26644 ( \35242_35542 , \35237_35537 , \35241_35541 );
and \U$26645 ( \35243_35543 , \34691_34991 , \34695_34995 );
and \U$26646 ( \35244_35544 , \34695_34995 , \34700_35000 );
and \U$26647 ( \35245_35545 , \34691_34991 , \34700_35000 );
or \U$26648 ( \35246_35546 , \35243_35543 , \35244_35544 , \35245_35545 );
and \U$26649 ( \35247_35547 , \34770_35070 , \34774_35074 );
and \U$26650 ( \35248_35548 , \34774_35074 , \34779_35079 );
and \U$26651 ( \35249_35549 , \34770_35070 , \34779_35079 );
or \U$26652 ( \35250_35550 , \35247_35547 , \35248_35548 , \35249_35549 );
xor \U$26653 ( \35251_35551 , \35246_35546 , \35250_35550 );
and \U$26654 ( \35252_35552 , \34719_35019 , \34723_35023 );
and \U$26655 ( \35253_35553 , \34723_35023 , \34728_35028 );
and \U$26656 ( \35254_35554 , \34719_35019 , \34728_35028 );
or \U$26657 ( \35255_35555 , \35252_35552 , \35253_35553 , \35254_35554 );
xor \U$26658 ( \35256_35556 , \35251_35551 , \35255_35555 );
xor \U$26659 ( \35257_35557 , \35242_35542 , \35256_35556 );
xor \U$26660 ( \35258_35558 , \35233_35533 , \35257_35557 );
xor \U$26661 ( \35259_35559 , \35184_35484 , \35258_35558 );
xor \U$26662 ( \35260_35560 , \35138_35438 , \35259_35559 );
and \U$26663 ( \35261_35561 , \34653_34953 , \34704_35004 );
and \U$26664 ( \35262_35562 , \34704_35004 , \34783_35083 );
and \U$26665 ( \35263_35563 , \34653_34953 , \34783_35083 );
or \U$26666 ( \35264_35564 , \35261_35561 , \35262_35562 , \35263_35563 );
xor \U$26667 ( \35265_35565 , \35260_35560 , \35264_35564 );
and \U$26668 ( \35266_35566 , \34784_35084 , \34788_35088 );
and \U$26669 ( \35267_35567 , \34789_35089 , \34792_35092 );
or \U$26670 ( \35268_35568 , \35266_35566 , \35267_35567 );
xor \U$26671 ( \35269_35569 , \35265_35565 , \35268_35568 );
buf g9b9c_GF_PartitionCandidate( \35270_35570_nG9b9c , \35269_35569 );
and \U$26672 ( \35271_35571 , \10402_10704 , \35270_35570_nG9b9c );
or \U$26673 ( \35272_35572 , \35129_35429 , \35271_35571 );
xor \U$26674 ( \35273_35573 , \10399_10703 , \35272_35572 );
buf \U$26675 ( \35274_35574 , \35273_35573 );
buf \U$26677 ( \35275_35575 , \35274_35574 );
xor \U$26678 ( \35276_35576 , \35128_35428 , \35275_35575 );
buf \U$26679 ( \35277_35577 , \35276_35576 );
xor \U$26680 ( \35278_35578 , \35053_35353 , \35277_35577 );
buf \U$26681 ( \35279_35579 , \35278_35578 );
xor \U$26682 ( \35280_35580 , \34999_35299 , \35279_35579 );
and \U$26683 ( \35281_35581 , \34920_35220 , \35280_35580 );
and \U$26685 ( \35282_35582 , \34914_35214 , \34919_35219 );
or \U$26687 ( \35283_35583 , 1'b0 , \35282_35582 , 1'b0 );
xor \U$26688 ( \35284_35584 , \35281_35581 , \35283_35583 );
and \U$26690 ( \35285_35585 , \34907_35207 , \34913_35213 );
and \U$26691 ( \35286_35586 , \34909_35209 , \34913_35213 );
or \U$26692 ( \35287_35587 , 1'b0 , \35285_35585 , \35286_35586 );
xor \U$26693 ( \35288_35588 , \35284_35584 , \35287_35587 );
xor \U$26700 ( \35289_35589 , \35288_35588 , 1'b0 );
and \U$26701 ( \35290_35590 , \34925_35225 , \34998_35298 );
and \U$26702 ( \35291_35591 , \34925_35225 , \35279_35579 );
and \U$26703 ( \35292_35592 , \34998_35298 , \35279_35579 );
or \U$26704 ( \35293_35593 , \35290_35590 , \35291_35591 , \35292_35592 );
xor \U$26705 ( \35294_35594 , \35289_35589 , \35293_35593 );
and \U$26706 ( \35295_35595 , \35047_35347 , \35052_35352 );
and \U$26707 ( \35296_35596 , \35047_35347 , \35277_35577 );
and \U$26708 ( \35297_35597 , \35052_35352 , \35277_35577 );
or \U$26709 ( \35298_35598 , \35295_35595 , \35296_35596 , \35297_35597 );
buf \U$26710 ( \35299_35599 , \35298_35598 );
and \U$26711 ( \35300_35600 , \35019_35319 , \35025_35325 );
and \U$26712 ( \35301_35601 , \35019_35319 , \35032_35332 );
and \U$26713 ( \35302_35602 , \35025_35325 , \35032_35332 );
or \U$26714 ( \35303_35603 , \35300_35600 , \35301_35601 , \35302_35602 );
buf \U$26715 ( \35304_35604 , \35303_35603 );
and \U$26716 ( \35305_35605 , \35004_35304 , \35010_35310 );
and \U$26717 ( \35306_35606 , \35004_35304 , \35017_35317 );
and \U$26718 ( \35307_35607 , \35010_35310 , \35017_35317 );
or \U$26719 ( \35308_35608 , \35305_35605 , \35306_35606 , \35307_35607 );
buf \U$26720 ( \35309_35609 , \35308_35608 );
and \U$26721 ( \35310_35610 , \14710_14631 , \31877_32179_nG9bb4 );
and \U$26722 ( \35311_35611 , \14329_14628 , \32589_32888_nG9bb1 );
or \U$26723 ( \35312_35612 , \35310_35610 , \35311_35611 );
xor \U$26724 ( \35313_35613 , \14328_14627 , \35312_35612 );
buf \U$26725 ( \35314_35614 , \35313_35613 );
buf \U$26727 ( \35315_35615 , \35314_35614 );
xor \U$26728 ( \35316_35616 , \35309_35609 , \35315_35615 );
and \U$26729 ( \35317_35617 , \13431_13370 , \32881_33181_nG9bae );
and \U$26730 ( \35318_35618 , \13068_13367 , \33313_33613_nG9bab );
or \U$26731 ( \35319_35619 , \35317_35617 , \35318_35618 );
xor \U$26732 ( \35320_35620 , \13067_13366 , \35319_35619 );
buf \U$26733 ( \35321_35621 , \35320_35620 );
buf \U$26735 ( \35322_35622 , \35321_35621 );
xor \U$26736 ( \35323_35623 , \35316_35616 , \35322_35622 );
buf \U$26737 ( \35324_35624 , \35323_35623 );
xor \U$26738 ( \35325_35625 , \35304_35604 , \35324_35624 );
and \U$26739 ( \35326_35626 , \34941_35241 , \34946_35246 );
and \U$26740 ( \35327_35627 , \34941_35241 , \34981_35281 );
and \U$26741 ( \35328_35628 , \34946_35246 , \34981_35281 );
or \U$26742 ( \35329_35629 , \35326_35626 , \35327_35627 , \35328_35628 );
buf \U$26743 ( \35330_35630 , \35329_35629 );
xor \U$26744 ( \35331_35631 , \35325_35625 , \35330_35630 );
buf \U$26745 ( \35332_35632 , \35331_35631 );
xor \U$26746 ( \35333_35633 , \35299_35599 , \35332_35632 );
and \U$26747 ( \35334_35634 , \35074_35374 , \35127_35427 );
and \U$26748 ( \35335_35635 , \35074_35374 , \35275_35575 );
and \U$26749 ( \35336_35636 , \35127_35427 , \35275_35575 );
or \U$26750 ( \35337_35637 , \35334_35634 , \35335_35635 , \35336_35636 );
buf \U$26751 ( \35338_35638 , \35337_35637 );
and \U$26752 ( \35339_35639 , \35103_35403 , \35109_35409 );
and \U$26753 ( \35340_35640 , \35103_35403 , \35116_35416 );
and \U$26754 ( \35341_35641 , \35109_35409 , \35116_35416 );
or \U$26755 ( \35342_35642 , \35339_35639 , \35340_35640 , \35341_35641 );
buf \U$26756 ( \35343_35643 , \35342_35642 );
and \U$26757 ( \35344_35644 , \23495_23201 , \21827_22129_nG9bd8 );
and \U$26758 ( \35345_35645 , \22899_23198 , \22330_22629_nG9bd5 );
or \U$26759 ( \35346_35646 , \35344_35644 , \35345_35645 );
xor \U$26760 ( \35347_35647 , \22898_23197 , \35346_35646 );
buf \U$26761 ( \35348_35648 , \35347_35647 );
buf \U$26763 ( \35349_35649 , \35348_35648 );
xor \U$26764 ( \35350_35650 , \35343_35643 , \35349_35649 );
and \U$26765 ( \35351_35651 , \21908_21658 , \23394_23696_nG9bd2 );
and \U$26766 ( \35352_35652 , \21356_21655 , \23927_24226_nG9bcf );
or \U$26767 ( \35353_35653 , \35351_35651 , \35352_35652 );
xor \U$26768 ( \35354_35654 , \21355_21654 , \35353_35653 );
buf \U$26769 ( \35355_35655 , \35354_35654 );
buf \U$26771 ( \35356_35656 , \35355_35655 );
xor \U$26772 ( \35357_35657 , \35350_35650 , \35356_35656 );
buf \U$26773 ( \35358_35658 , \35357_35657 );
and \U$26774 ( \35359_35659 , \10996_10421 , \34343_34643_nG9ba2 );
and \U$26775 ( \35360_35660 , \10119_10418 , \34794_35094_nG9b9f );
or \U$26776 ( \35361_35661 , \35359_35659 , \35360_35660 );
xor \U$26777 ( \35362_35662 , \10118_10417 , \35361_35661 );
buf \U$26778 ( \35363_35663 , \35362_35662 );
buf \U$26780 ( \35364_35664 , \35363_35663 );
xor \U$26781 ( \35365_35665 , \35358_35658 , \35364_35664 );
and \U$26782 ( \35366_35666 , \10411_10707 , \35270_35570_nG9b9c );
and \U$26783 ( \35367_35667 , \35188_35488 , \35232_35532 );
and \U$26784 ( \35368_35668 , \35232_35532 , \35257_35557 );
and \U$26785 ( \35369_35669 , \35188_35488 , \35257_35557 );
or \U$26786 ( \35370_35670 , \35367_35667 , \35368_35668 , \35369_35669 );
and \U$26787 ( \35371_35671 , \35142_35442 , \35183_35483 );
and \U$26788 ( \35372_35672 , \35183_35483 , \35258_35558 );
and \U$26789 ( \35373_35673 , \35142_35442 , \35258_35558 );
or \U$26790 ( \35374_35674 , \35371_35671 , \35372_35672 , \35373_35673 );
xor \U$26791 ( \35375_35675 , \35370_35670 , \35374_35674 );
and \U$26792 ( \35376_35676 , \35146_35446 , \35150_35450 );
and \U$26793 ( \35377_35677 , \35150_35450 , \35182_35482 );
and \U$26794 ( \35378_35678 , \35146_35446 , \35182_35482 );
or \U$26795 ( \35379_35679 , \35376_35676 , \35377_35677 , \35378_35678 );
and \U$26796 ( \35380_35680 , \35201_35501 , \35215_35515 );
and \U$26797 ( \35381_35681 , \35215_35515 , \35231_35531 );
and \U$26798 ( \35382_35682 , \35201_35501 , \35231_35531 );
or \U$26799 ( \35383_35683 , \35380_35680 , \35381_35681 , \35382_35682 );
and \U$26800 ( \35384_35684 , \35237_35537 , \35241_35541 );
and \U$26801 ( \35385_35685 , \35241_35541 , \35256_35556 );
and \U$26802 ( \35386_35686 , \35237_35537 , \35256_35556 );
or \U$26803 ( \35387_35687 , \35384_35684 , \35385_35685 , \35386_35686 );
xor \U$26804 ( \35388_35688 , \35383_35683 , \35387_35687 );
and \U$26805 ( \35389_35689 , \35246_35546 , \35250_35550 );
and \U$26806 ( \35390_35690 , \35250_35550 , \35255_35555 );
and \U$26807 ( \35391_35691 , \35246_35546 , \35255_35555 );
or \U$26808 ( \35392_35692 , \35389_35689 , \35390_35690 , \35391_35691 );
and \U$26809 ( \35393_35693 , \35220_35520 , \35225_35525 );
and \U$26810 ( \35394_35694 , \35225_35525 , \35230_35530 );
and \U$26811 ( \35395_35695 , \35220_35520 , \35230_35530 );
or \U$26812 ( \35396_35696 , \35393_35693 , \35394_35694 , \35395_35695 );
xor \U$26813 ( \35397_35697 , \35392_35692 , \35396_35696 );
and \U$26814 ( \35398_35698 , \35191_35491 , \35195_35495 );
and \U$26815 ( \35399_35699 , \35195_35495 , \35200_35500 );
and \U$26816 ( \35400_35700 , \35191_35491 , \35200_35500 );
or \U$26817 ( \35401_35701 , \35398_35698 , \35399_35699 , \35400_35700 );
and \U$26818 ( \35402_35702 , \35205_35505 , \35209_35509 );
and \U$26819 ( \35403_35703 , \35209_35509 , \35214_35514 );
and \U$26820 ( \35404_35704 , \35205_35505 , \35214_35514 );
or \U$26821 ( \35405_35705 , \35402_35702 , \35403_35703 , \35404_35704 );
xor \U$26822 ( \35406_35706 , \35401_35701 , \35405_35705 );
and \U$26823 ( \35407_35707 , \35171_35471 , \35175_35475 );
and \U$26824 ( \35408_35708 , \35175_35475 , \35180_35480 );
and \U$26825 ( \35409_35709 , \35171_35471 , \35180_35480 );
or \U$26826 ( \35410_35710 , \35407_35707 , \35408_35708 , \35409_35709 );
xor \U$26827 ( \35411_35711 , \35406_35706 , \35410_35710 );
xor \U$26828 ( \35412_35712 , \35397_35697 , \35411_35711 );
xor \U$26829 ( \35413_35713 , \35388_35688 , \35412_35712 );
xor \U$26830 ( \35414_35714 , \35379_35679 , \35413_35713 );
and \U$26831 ( \35415_35715 , \35155_35455 , \35166_35466 );
and \U$26832 ( \35416_35716 , \35166_35466 , \35181_35481 );
and \U$26833 ( \35417_35717 , \35155_35455 , \35181_35481 );
or \U$26834 ( \35418_35718 , \35415_35715 , \35416_35716 , \35417_35717 );
and \U$26835 ( \35419_35719 , \35159_35459 , \35163_35463 );
and \U$26836 ( \35420_35720 , \35163_35463 , \35165_35465 );
and \U$26837 ( \35421_35721 , \35159_35459 , \35165_35465 );
or \U$26838 ( \35422_35722 , \35419_35719 , \35420_35720 , \35421_35721 );
and \U$26839 ( \35423_35723 , \26527_26829 , \19235_19534 );
and \U$26840 ( \35424_35724 , \27011_27313 , \18743_19045 );
nor \U$26841 ( \35425_35725 , \35423_35723 , \35424_35724 );
xnor \U$26842 ( \35426_35726 , \35425_35725 , \19241_19540 );
and \U$26843 ( \35427_35727 , \21788_22090 , \23839_24138 );
and \U$26844 ( \35428_35728 , \22257_22556 , \23328_23630 );
nor \U$26845 ( \35429_35729 , \35427_35727 , \35428_35728 );
xnor \U$26846 ( \35430_35730 , \35429_35729 , \23845_24144 );
xor \U$26847 ( \35431_35731 , \35426_35726 , \35430_35730 );
and \U$26848 ( \35432_35732 , \20242_20544 , \25527_25826 );
and \U$26849 ( \35433_35733 , \20734_21033 , \24962_25264 );
nor \U$26850 ( \35434_35734 , \35432_35732 , \35433_35733 );
xnor \U$26851 ( \35435_35735 , \35434_35734 , \25474_25773 );
xor \U$26852 ( \35436_35736 , \35431_35731 , \35435_35735 );
xor \U$26853 ( \35437_35737 , \35422_35722 , \35436_35736 );
not \U$26854 ( \35438_35738 , \13736_14035 );
and \U$26855 ( \35439_35739 , \31752_32054 , \15037_15336 );
and \U$26856 ( \35440_35740 , \32495_32794 , \14661_14963 );
nor \U$26857 ( \35441_35741 , \35439_35739 , \35440_35740 );
xnor \U$26858 ( \35442_35742 , \35441_35741 , \15043_15342 );
xor \U$26859 ( \35443_35743 , \35438_35738 , \35442_35742 );
and \U$26860 ( \35444_35744 , \28232_28534 , \17791_18090 );
and \U$26861 ( \35445_35745 , \28782_29084 , \17353_17655 );
nor \U$26862 ( \35446_35746 , \35444_35744 , \35445_35745 );
xnor \U$26863 ( \35447_35747 , \35446_35746 , \17747_18046 );
xor \U$26864 ( \35448_35748 , \35443_35743 , \35447_35747 );
xor \U$26865 ( \35449_35749 , \35437_35737 , \35448_35748 );
xor \U$26866 ( \35450_35750 , \35418_35718 , \35449_35749 );
and \U$26867 ( \35451_35751 , \24970_25272 , \20706_21005 );
and \U$26868 ( \35452_35752 , \25516_25815 , \20255_20557 );
nor \U$26869 ( \35453_35753 , \35451_35751 , \35452_35752 );
xnor \U$26870 ( \35454_35754 , \35453_35753 , \20712_21011 );
and \U$26871 ( \35455_35755 , \15965_16267 , \30521_30823 );
and \U$26872 ( \35456_35756 , \16353_16655 , \29944_30246 );
nor \U$26873 ( \35457_35757 , \35455_35755 , \35456_35756 );
xnor \U$26874 ( \35458_35758 , \35457_35757 , \30511_30813 );
xor \U$26875 ( \35459_35759 , \35454_35754 , \35458_35758 );
and \U$26876 ( \35460_35760 , \14648_14950 , \32555_32854 );
and \U$26877 ( \35461_35761 , \15022_15321 , \31765_32067 );
nor \U$26878 ( \35462_35762 , \35460_35760 , \35461_35761 );
xnor \U$26879 ( \35463_35763 , \35462_35762 , \32506_32805 );
xor \U$26880 ( \35464_35764 , \35459_35759 , \35463_35763 );
and \U$26881 ( \35465_35765 , \29966_30268 , \16333_16635 );
and \U$26882 ( \35466_35766 , \30500_30802 , \15999_16301 );
nor \U$26883 ( \35467_35767 , \35465_35765 , \35466_35766 );
xnor \U$26884 ( \35468_35768 , \35467_35767 , \16323_16625 );
and \U$26885 ( \35469_35769 , \18730_19032 , \27095_27397 );
and \U$26886 ( \35470_35770 , \19259_19558 , \26505_26807 );
nor \U$26887 ( \35471_35771 , \35469_35769 , \35470_35770 );
xnor \U$26888 ( \35472_35772 , \35471_35771 , \26993_27295 );
xor \U$26889 ( \35473_35773 , \35468_35768 , \35472_35772 );
and \U$26890 ( \35474_35774 , \17325_17627 , \28768_29070 );
and \U$26891 ( \35475_35775 , \17736_18035 , \28224_28526 );
nor \U$26892 ( \35476_35776 , \35474_35774 , \35475_35775 );
xnor \U$26893 ( \35477_35777 , \35476_35776 , \28774_29076 );
xor \U$26894 ( \35478_35778 , \35473_35773 , \35477_35777 );
xor \U$26895 ( \35479_35779 , \35464_35764 , \35478_35778 );
buf \U$26896 ( \35480_35780 , \35224_35524 );
and \U$26897 ( \35481_35781 , \23315_23617 , \22243_22542 );
and \U$26898 ( \35482_35782 , \23900_24199 , \21801_22103 );
nor \U$26899 ( \35483_35783 , \35481_35781 , \35482_35782 );
xnor \U$26900 ( \35484_35784 , \35483_35783 , \22249_22548 );
xor \U$26901 ( \35485_35785 , \35480_35780 , \35484_35784 );
and \U$26902 ( \35486_35786 , \13725_14024 , \32503_32802 );
xor \U$26903 ( \35487_35787 , \35485_35785 , \35486_35786 );
xor \U$26904 ( \35488_35788 , \35479_35779 , \35487_35787 );
xor \U$26905 ( \35489_35789 , \35450_35750 , \35488_35788 );
xor \U$26906 ( \35490_35790 , \35414_35714 , \35489_35789 );
xor \U$26907 ( \35491_35791 , \35375_35675 , \35490_35790 );
and \U$26908 ( \35492_35792 , \35133_35433 , \35137_35437 );
and \U$26909 ( \35493_35793 , \35137_35437 , \35259_35559 );
and \U$26910 ( \35494_35794 , \35133_35433 , \35259_35559 );
or \U$26911 ( \35495_35795 , \35492_35792 , \35493_35793 , \35494_35794 );
xor \U$26912 ( \35496_35796 , \35491_35791 , \35495_35795 );
and \U$26913 ( \35497_35797 , \35260_35560 , \35264_35564 );
and \U$26914 ( \35498_35798 , \35265_35565 , \35268_35568 );
or \U$26915 ( \35499_35799 , \35497_35797 , \35498_35798 );
xor \U$26916 ( \35500_35800 , \35496_35796 , \35499_35799 );
buf g9b99_GF_PartitionCandidate( \35501_35801_nG9b99 , \35500_35800 );
and \U$26917 ( \35502_35802 , \10402_10704 , \35501_35801_nG9b99 );
or \U$26918 ( \35503_35803 , \35366_35666 , \35502_35802 );
xor \U$26919 ( \35504_35804 , \10399_10703 , \35503_35803 );
buf \U$26920 ( \35505_35805 , \35504_35804 );
buf \U$26922 ( \35506_35806 , \35505_35805 );
xor \U$26923 ( \35507_35807 , \35365_35665 , \35506_35806 );
buf \U$26924 ( \35508_35808 , \35507_35807 );
xor \U$26925 ( \35509_35809 , \35338_35638 , \35508_35808 );
and \U$26926 ( \35510_35810 , \35092_35392 , \35094_35394 );
and \U$26927 ( \35511_35811 , \35092_35392 , \35101_35401 );
and \U$26928 ( \35512_35812 , \35094_35394 , \35101_35401 );
or \U$26929 ( \35513_35813 , \35510_35810 , \35511_35811 , \35512_35812 );
buf \U$26930 ( \35514_35814 , \35513_35813 );
and \U$26931 ( \35515_35815 , \28946_28118 , \17363_17665_nG9bea );
and \U$26932 ( \35516_35816 , \27816_28115 , \17808_18107_nG9be7 );
or \U$26933 ( \35517_35817 , \35515_35815 , \35516_35816 );
xor \U$26934 ( \35518_35818 , \27815_28114 , \35517_35817 );
buf \U$26935 ( \35519_35819 , \35518_35818 );
buf \U$26937 ( \35520_35820 , \35519_35819 );
xor \U$26938 ( \35521_35821 , \35514_35814 , \35520_35820 );
and \U$26939 ( \35522_35822 , \25044_24792 , \20306_20608_nG9bde );
and \U$26940 ( \35523_35823 , \24490_24789 , \20787_21086_nG9bdb );
or \U$26941 ( \35524_35824 , \35522_35822 , \35523_35823 );
xor \U$26942 ( \35525_35825 , \24489_24788 , \35524_35824 );
buf \U$26943 ( \35526_35826 , \35525_35825 );
buf \U$26945 ( \35527_35827 , \35526_35826 );
xor \U$26946 ( \35528_35828 , \35521_35821 , \35527_35827 );
buf \U$26947 ( \35529_35829 , \35528_35828 );
and \U$26948 ( \35530_35830 , \20353_20155 , \24996_25298_nG9bcc );
and \U$26949 ( \35531_35831 , \19853_20152 , \25561_25860_nG9bc9 );
or \U$26950 ( \35532_35832 , \35530_35830 , \35531_35831 );
xor \U$26951 ( \35533_35833 , \19852_20151 , \35532_35832 );
buf \U$26952 ( \35534_35834 , \35533_35833 );
buf \U$26954 ( \35535_35835 , \35534_35834 );
xor \U$26955 ( \35536_35836 , \35529_35829 , \35535_35835 );
and \U$26956 ( \35537_35837 , \18908_18702 , \26585_26887_nG9bc6 );
and \U$26957 ( \35538_35838 , \18400_18699 , \27114_27416_nG9bc3 );
or \U$26958 ( \35539_35839 , \35537_35837 , \35538_35838 );
xor \U$26959 ( \35540_35840 , \18399_18698 , \35539_35839 );
buf \U$26960 ( \35541_35841 , \35540_35840 );
buf \U$26962 ( \35542_35842 , \35541_35841 );
xor \U$26963 ( \35543_35843 , \35536_35836 , \35542_35842 );
buf \U$26964 ( \35544_35844 , \35543_35843 );
and \U$26965 ( \35545_35845 , \34952_35252 , \34972_35272 );
and \U$26966 ( \35546_35846 , \34952_35252 , \34979_35279 );
and \U$26967 ( \35547_35847 , \34972_35272 , \34979_35279 );
or \U$26968 ( \35548_35848 , \35545_35845 , \35546_35846 , \35547_35847 );
buf \U$26969 ( \35549_35849 , \35548_35848 );
xor \U$26970 ( \35550_35850 , \35544_35844 , \35549_35849 );
and \U$26971 ( \35551_35851 , \12183_12157 , \33741_34041_nG9ba8 );
and \U$26972 ( \35552_35852 , \11855_12154 , \33994_34294_nG9ba5 );
or \U$26973 ( \35553_35853 , \35551_35851 , \35552_35852 );
xor \U$26974 ( \35554_35854 , \11854_12153 , \35553_35853 );
buf \U$26975 ( \35555_35855 , \35554_35854 );
buf \U$26977 ( \35556_35856 , \35555_35855 );
xor \U$26978 ( \35557_35857 , \35550_35850 , \35556_35856 );
buf \U$26979 ( \35558_35858 , \35557_35857 );
xor \U$26980 ( \35559_35859 , \35509_35809 , \35558_35858 );
buf \U$26981 ( \35560_35860 , \35559_35859 );
xor \U$26982 ( \35561_35861 , \35333_35633 , \35560_35860 );
buf \U$26983 ( \35562_35862 , \35561_35861 );
and \U$26984 ( \35563_35863 , \34985_35285 , \34990_35290 );
and \U$26985 ( \35564_35864 , \34985_35285 , \34996_35296 );
and \U$26986 ( \35565_35865 , \34990_35290 , \34996_35296 );
or \U$26987 ( \35566_35866 , \35563_35863 , \35564_35864 , \35565_35865 );
buf \U$26988 ( \35567_35867 , \35566_35866 );
xor \U$26989 ( \35568_35868 , \35562_35862 , \35567_35867 );
and \U$26990 ( \35569_35869 , \35034_35334 , \35039_35339 );
and \U$26991 ( \35570_35870 , \35034_35334 , \35045_35345 );
and \U$26992 ( \35571_35871 , \35039_35339 , \35045_35345 );
or \U$26993 ( \35572_35872 , \35569_35869 , \35570_35870 , \35571_35871 );
buf \U$26994 ( \35573_35873 , \35572_35872 );
and \U$26995 ( \35574_35874 , \34930_35230 , \34935_35235 );
and \U$26996 ( \35575_35875 , \34930_35230 , \34983_35283 );
and \U$26997 ( \35576_35876 , \34935_35235 , \34983_35283 );
or \U$26998 ( \35577_35877 , \35574_35874 , \35575_35875 , \35576_35876 );
buf \U$26999 ( \35578_35878 , \35577_35877 );
xor \U$27000 ( \35579_35879 , \35573_35873 , \35578_35878 );
and \U$27001 ( \35580_35880 , \35059_35359 , \35065_35365 );
and \U$27002 ( \35581_35881 , \35059_35359 , \35072_35372 );
and \U$27003 ( \35582_35882 , \35065_35365 , \35072_35372 );
or \U$27004 ( \35583_35883 , \35580_35880 , \35581_35881 , \35582_35882 );
buf \U$27005 ( \35584_35884 , \35583_35883 );
and \U$27006 ( \35585_35885 , \34957_35257 , \34963_35263 );
and \U$27007 ( \35586_35886 , \34957_35257 , \34970_35270 );
and \U$27008 ( \35587_35887 , \34963_35263 , \34970_35270 );
or \U$27009 ( \35588_35888 , \35585_35885 , \35586_35886 , \35587_35887 );
buf \U$27010 ( \35589_35889 , \35588_35888 );
and \U$27012 ( \35590_35890 , \32617_32916 , \13771_14070_nG9bf9 );
or \U$27013 ( \35591_35891 , 1'b0 , \35590_35890 );
xor \U$27014 ( \35592_35892 , 1'b0 , \35591_35891 );
buf \U$27015 ( \35593_35893 , \35592_35892 );
buf \U$27017 ( \35594_35894 , \35593_35893 );
and \U$27018 ( \35595_35895 , \31989_31636 , \14682_14984_nG9bf6 );
and \U$27019 ( \35596_35896 , \31334_31633 , \15074_15373_nG9bf3 );
or \U$27020 ( \35597_35897 , \35595_35895 , \35596_35896 );
xor \U$27021 ( \35598_35898 , \31333_31632 , \35597_35897 );
buf \U$27022 ( \35599_35899 , \35598_35898 );
buf \U$27024 ( \35600_35900 , \35599_35899 );
xor \U$27025 ( \35601_35901 , \35594_35894 , \35600_35900 );
buf \U$27026 ( \35602_35902 , \35601_35901 );
and \U$27027 ( \35603_35903 , \35084_35384 , \35090_35390 );
buf \U$27028 ( \35604_35904 , \35603_35903 );
xor \U$27029 ( \35605_35905 , \35602_35902 , \35604_35904 );
and \U$27030 ( \35606_35906 , \30670_29853 , \16013_16315_nG9bf0 );
and \U$27031 ( \35607_35907 , \29551_29850 , \16378_16680_nG9bed );
or \U$27032 ( \35608_35908 , \35606_35906 , \35607_35907 );
xor \U$27033 ( \35609_35909 , \29550_29849 , \35608_35908 );
buf \U$27034 ( \35610_35910 , \35609_35909 );
buf \U$27036 ( \35611_35911 , \35610_35910 );
xor \U$27037 ( \35612_35912 , \35605_35905 , \35611_35911 );
buf \U$27038 ( \35613_35913 , \35612_35912 );
xor \U$27039 ( \35614_35914 , \35589_35889 , \35613_35913 );
and \U$27040 ( \35615_35915 , \27141_26431 , \18789_19091_nG9be4 );
and \U$27041 ( \35616_35916 , \26129_26428 , \19287_19586_nG9be1 );
or \U$27042 ( \35617_35917 , \35615_35915 , \35616_35916 );
xor \U$27043 ( \35618_35918 , \26128_26427 , \35617_35917 );
buf \U$27044 ( \35619_35919 , \35618_35918 );
buf \U$27046 ( \35620_35920 , \35619_35919 );
xor \U$27047 ( \35621_35921 , \35614_35914 , \35620_35920 );
buf \U$27048 ( \35622_35922 , \35621_35921 );
and \U$27049 ( \35623_35923 , \17437_17297 , \28300_28602_nG9bc0 );
and \U$27050 ( \35624_35924 , \16995_17294 , \28877_29179_nG9bbd );
or \U$27051 ( \35625_35925 , \35623_35923 , \35624_35924 );
xor \U$27052 ( \35626_35926 , \16994_17293 , \35625_35925 );
buf \U$27053 ( \35627_35927 , \35626_35926 );
buf \U$27055 ( \35628_35928 , \35627_35927 );
xor \U$27056 ( \35629_35929 , \35622_35922 , \35628_35928 );
and \U$27057 ( \35630_35930 , \16405_15940 , \30064_30366_nG9bba );
and \U$27058 ( \35631_35931 , \15638_15937 , \30638_30940_nG9bb7 );
or \U$27059 ( \35632_35932 , \35630_35930 , \35631_35931 );
xor \U$27060 ( \35633_35933 , \15637_15936 , \35632_35932 );
buf \U$27061 ( \35634_35934 , \35633_35933 );
buf \U$27063 ( \35635_35935 , \35634_35934 );
xor \U$27064 ( \35636_35936 , \35629_35929 , \35635_35935 );
buf \U$27065 ( \35637_35937 , \35636_35936 );
xor \U$27066 ( \35638_35938 , \35584_35884 , \35637_35937 );
and \U$27067 ( \35639_35939 , \35079_35379 , \35118_35418 );
and \U$27068 ( \35640_35940 , \35079_35379 , \35125_35425 );
and \U$27069 ( \35641_35941 , \35118_35418 , \35125_35425 );
or \U$27070 ( \35642_35942 , \35639_35939 , \35640_35940 , \35641_35941 );
buf \U$27071 ( \35643_35943 , \35642_35942 );
xor \U$27072 ( \35644_35944 , \35638_35938 , \35643_35943 );
buf \U$27073 ( \35645_35945 , \35644_35944 );
xor \U$27074 ( \35646_35946 , \35579_35879 , \35645_35945 );
buf \U$27075 ( \35647_35947 , \35646_35946 );
xor \U$27076 ( \35648_35948 , \35568_35868 , \35647_35947 );
and \U$27077 ( \35649_35949 , \35294_35594 , \35648_35948 );
and \U$27079 ( \35650_35950 , \35288_35588 , \35293_35593 );
or \U$27081 ( \35651_35951 , 1'b0 , \35650_35950 , 1'b0 );
xor \U$27082 ( \35652_35952 , \35649_35949 , \35651_35951 );
and \U$27084 ( \35653_35953 , \35281_35581 , \35287_35587 );
and \U$27085 ( \35654_35954 , \35283_35583 , \35287_35587 );
or \U$27086 ( \35655_35955 , 1'b0 , \35653_35953 , \35654_35954 );
xor \U$27087 ( \35656_35956 , \35652_35952 , \35655_35955 );
xor \U$27094 ( \35657_35957 , \35656_35956 , 1'b0 );
and \U$27095 ( \35658_35958 , \35562_35862 , \35567_35867 );
and \U$27096 ( \35659_35959 , \35562_35862 , \35647_35947 );
and \U$27097 ( \35660_35960 , \35567_35867 , \35647_35947 );
or \U$27098 ( \35661_35961 , \35658_35958 , \35659_35959 , \35660_35960 );
xor \U$27099 ( \35662_35962 , \35657_35957 , \35661_35961 );
and \U$27100 ( \35663_35963 , \35573_35873 , \35578_35878 );
and \U$27101 ( \35664_35964 , \35573_35873 , \35645_35945 );
and \U$27102 ( \35665_35965 , \35578_35878 , \35645_35945 );
or \U$27103 ( \35666_35966 , \35663_35963 , \35664_35964 , \35665_35965 );
buf \U$27104 ( \35667_35967 , \35666_35966 );
and \U$27105 ( \35668_35968 , \35338_35638 , \35508_35808 );
and \U$27106 ( \35669_35969 , \35338_35638 , \35558_35858 );
and \U$27107 ( \35670_35970 , \35508_35808 , \35558_35858 );
or \U$27108 ( \35671_35971 , \35668_35968 , \35669_35969 , \35670_35970 );
buf \U$27109 ( \35672_35972 , \35671_35971 );
xor \U$27110 ( \35673_35973 , \35667_35967 , \35672_35972 );
and \U$27111 ( \35674_35974 , \35584_35884 , \35637_35937 );
and \U$27112 ( \35675_35975 , \35584_35884 , \35643_35943 );
and \U$27113 ( \35676_35976 , \35637_35937 , \35643_35943 );
or \U$27114 ( \35677_35977 , \35674_35974 , \35675_35975 , \35676_35976 );
buf \U$27115 ( \35678_35978 , \35677_35977 );
and \U$27116 ( \35679_35979 , \35622_35922 , \35628_35928 );
and \U$27117 ( \35680_35980 , \35622_35922 , \35635_35935 );
and \U$27118 ( \35681_35981 , \35628_35928 , \35635_35935 );
or \U$27119 ( \35682_35982 , \35679_35979 , \35680_35980 , \35681_35981 );
buf \U$27120 ( \35683_35983 , \35682_35982 );
and \U$27121 ( \35684_35984 , \35514_35814 , \35520_35820 );
and \U$27122 ( \35685_35985 , \35514_35814 , \35527_35827 );
and \U$27123 ( \35686_35986 , \35520_35820 , \35527_35827 );
or \U$27124 ( \35687_35987 , \35684_35984 , \35685_35985 , \35686_35986 );
buf \U$27125 ( \35688_35988 , \35687_35987 );
and \U$27126 ( \35689_35989 , \21908_21658 , \23927_24226_nG9bcf );
and \U$27127 ( \35690_35990 , \21356_21655 , \24996_25298_nG9bcc );
or \U$27128 ( \35691_35991 , \35689_35989 , \35690_35990 );
xor \U$27129 ( \35692_35992 , \21355_21654 , \35691_35991 );
buf \U$27130 ( \35693_35993 , \35692_35992 );
buf \U$27132 ( \35694_35994 , \35693_35993 );
xor \U$27133 ( \35695_35995 , \35688_35988 , \35694_35994 );
and \U$27134 ( \35696_35996 , \18908_18702 , \27114_27416_nG9bc3 );
and \U$27135 ( \35697_35997 , \18400_18699 , \28300_28602_nG9bc0 );
or \U$27136 ( \35698_35998 , \35696_35996 , \35697_35997 );
xor \U$27137 ( \35699_35999 , \18399_18698 , \35698_35998 );
buf \U$27138 ( \35700_36000 , \35699_35999 );
buf \U$27140 ( \35701_36001 , \35700_36000 );
xor \U$27141 ( \35702_36002 , \35695_35995 , \35701_36001 );
buf \U$27142 ( \35703_36003 , \35702_36002 );
xor \U$27143 ( \35704_36004 , \35683_35983 , \35703_36003 );
and \U$27144 ( \35705_36005 , \12183_12157 , \33994_34294_nG9ba5 );
and \U$27145 ( \35706_36006 , \11855_12154 , \34343_34643_nG9ba2 );
or \U$27146 ( \35707_36007 , \35705_36005 , \35706_36006 );
xor \U$27147 ( \35708_36008 , \11854_12153 , \35707_36007 );
buf \U$27148 ( \35709_36009 , \35708_36008 );
buf \U$27150 ( \35710_36010 , \35709_36009 );
xor \U$27151 ( \35711_36011 , \35704_36004 , \35710_36010 );
buf \U$27152 ( \35712_36012 , \35711_36011 );
xor \U$27153 ( \35713_36013 , \35678_35978 , \35712_36012 );
and \U$27154 ( \35714_36014 , \35544_35844 , \35549_35849 );
and \U$27155 ( \35715_36015 , \35544_35844 , \35556_35856 );
and \U$27156 ( \35716_36016 , \35549_35849 , \35556_35856 );
or \U$27157 ( \35717_36017 , \35714_36014 , \35715_36015 , \35716_36016 );
buf \U$27158 ( \35718_36018 , \35717_36017 );
xor \U$27159 ( \35719_36019 , \35713_36013 , \35718_36018 );
buf \U$27160 ( \35720_36020 , \35719_36019 );
xor \U$27161 ( \35721_36021 , \35673_35973 , \35720_36020 );
buf \U$27162 ( \35722_36022 , \35721_36021 );
and \U$27163 ( \35723_36023 , \35299_35599 , \35332_35632 );
and \U$27164 ( \35724_36024 , \35299_35599 , \35560_35860 );
and \U$27165 ( \35725_36025 , \35332_35632 , \35560_35860 );
or \U$27166 ( \35726_36026 , \35723_36023 , \35724_36024 , \35725_36025 );
buf \U$27167 ( \35727_36027 , \35726_36026 );
xor \U$27168 ( \35728_36028 , \35722_36022 , \35727_36027 );
and \U$27169 ( \35729_36029 , \35529_35829 , \35535_35835 );
and \U$27170 ( \35730_36030 , \35529_35829 , \35542_35842 );
and \U$27171 ( \35731_36031 , \35535_35835 , \35542_35842 );
or \U$27172 ( \35732_36032 , \35729_36029 , \35730_36030 , \35731_36031 );
buf \U$27173 ( \35733_36033 , \35732_36032 );
and \U$27174 ( \35734_36034 , \10996_10421 , \34794_35094_nG9b9f );
and \U$27175 ( \35735_36035 , \10119_10418 , \35270_35570_nG9b9c );
or \U$27176 ( \35736_36036 , \35734_36034 , \35735_36035 );
xor \U$27177 ( \35737_36037 , \10118_10417 , \35736_36036 );
buf \U$27178 ( \35738_36038 , \35737_36037 );
buf \U$27180 ( \35739_36039 , \35738_36038 );
xor \U$27181 ( \35740_36040 , \35733_36033 , \35739_36039 );
and \U$27182 ( \35741_36041 , \10411_10707 , \35501_35801_nG9b99 );
and \U$27183 ( \35742_36042 , \35379_35679 , \35413_35713 );
and \U$27184 ( \35743_36043 , \35413_35713 , \35489_35789 );
and \U$27185 ( \35744_36044 , \35379_35679 , \35489_35789 );
or \U$27186 ( \35745_36045 , \35742_36042 , \35743_36043 , \35744_36044 );
and \U$27187 ( \35746_36046 , \35392_35692 , \35396_35696 );
and \U$27188 ( \35747_36047 , \35396_35696 , \35411_35711 );
and \U$27189 ( \35748_36048 , \35392_35692 , \35411_35711 );
or \U$27190 ( \35749_36049 , \35746_36046 , \35747_36047 , \35748_36048 );
and \U$27191 ( \35750_36050 , \27011_27313 , \19235_19534 );
and \U$27192 ( \35751_36051 , \28232_28534 , \18743_19045 );
nor \U$27193 ( \35752_36052 , \35750_36050 , \35751_36051 );
xnor \U$27194 ( \35753_36053 , \35752_36052 , \19241_19540 );
and \U$27195 ( \35754_36054 , \20734_21033 , \25527_25826 );
and \U$27196 ( \35755_36055 , \21788_22090 , \24962_25264 );
nor \U$27197 ( \35756_36056 , \35754_36054 , \35755_36055 );
xnor \U$27198 ( \35757_36057 , \35756_36056 , \25474_25773 );
xor \U$27199 ( \35758_36058 , \35753_36053 , \35757_36057 );
and \U$27200 ( \35759_36059 , \19259_19558 , \27095_27397 );
and \U$27201 ( \35760_36060 , \20242_20544 , \26505_26807 );
nor \U$27202 ( \35761_36061 , \35759_36059 , \35760_36060 );
xnor \U$27203 ( \35762_36062 , \35761_36061 , \26993_27295 );
xor \U$27204 ( \35763_36063 , \35758_36058 , \35762_36062 );
and \U$27205 ( \35764_36064 , \32495_32794 , \15037_15336 );
not \U$27206 ( \35765_36065 , \35764_36064 );
xnor \U$27207 ( \35766_36066 , \35765_36065 , \15043_15342 );
and \U$27208 ( \35767_36067 , \23900_24199 , \22243_22542 );
and \U$27209 ( \35768_36068 , \24970_25272 , \21801_22103 );
nor \U$27210 ( \35769_36069 , \35767_36067 , \35768_36068 );
xnor \U$27211 ( \35770_36070 , \35769_36069 , \22249_22548 );
xor \U$27212 ( \35771_36071 , \35766_36066 , \35770_36070 );
and \U$27213 ( \35772_36072 , \15022_15321 , \32555_32854 );
and \U$27214 ( \35773_36073 , \15965_16267 , \31765_32067 );
nor \U$27215 ( \35774_36074 , \35772_36072 , \35773_36073 );
xnor \U$27216 ( \35775_36075 , \35774_36074 , \32506_32805 );
xor \U$27217 ( \35776_36076 , \35771_36071 , \35775_36075 );
xor \U$27218 ( \35777_36077 , \35763_36063 , \35776_36076 );
and \U$27219 ( \35778_36078 , \25516_25815 , \20706_21005 );
and \U$27220 ( \35779_36079 , \26527_26829 , \20255_20557 );
nor \U$27221 ( \35780_36080 , \35778_36078 , \35779_36079 );
xnor \U$27222 ( \35781_36081 , \35780_36080 , \20712_21011 );
and \U$27223 ( \35782_36082 , \17736_18035 , \28768_29070 );
and \U$27224 ( \35783_36083 , \18730_19032 , \28224_28526 );
nor \U$27225 ( \35784_36084 , \35782_36082 , \35783_36083 );
xnor \U$27226 ( \35785_36085 , \35784_36084 , \28774_29076 );
xor \U$27227 ( \35786_36086 , \35781_36081 , \35785_36085 );
and \U$27228 ( \35787_36087 , \16353_16655 , \30521_30823 );
and \U$27229 ( \35788_36088 , \17325_17627 , \29944_30246 );
nor \U$27230 ( \35789_36089 , \35787_36087 , \35788_36088 );
xnor \U$27231 ( \35790_36090 , \35789_36089 , \30511_30813 );
xor \U$27232 ( \35791_36091 , \35786_36086 , \35790_36090 );
xor \U$27233 ( \35792_36092 , \35777_36077 , \35791_36091 );
xor \U$27234 ( \35793_36093 , \35749_36049 , \35792_36092 );
and \U$27235 ( \35794_36094 , \35401_35701 , \35405_35705 );
and \U$27236 ( \35795_36095 , \35405_35705 , \35410_35710 );
and \U$27237 ( \35796_36096 , \35401_35701 , \35410_35710 );
or \U$27238 ( \35797_36097 , \35794_36094 , \35795_36095 , \35796_36096 );
and \U$27239 ( \35798_36098 , \35480_35780 , \35484_35784 );
and \U$27240 ( \35799_36099 , \35484_35784 , \35486_35786 );
and \U$27241 ( \35800_36100 , \35480_35780 , \35486_35786 );
or \U$27242 ( \35801_36101 , \35798_36098 , \35799_36099 , \35800_36100 );
xor \U$27243 ( \35802_36102 , \35797_36097 , \35801_36101 );
and \U$27244 ( \35803_36103 , \35426_35726 , \35430_35730 );
and \U$27245 ( \35804_36104 , \35430_35730 , \35435_35735 );
and \U$27246 ( \35805_36105 , \35426_35726 , \35435_35735 );
or \U$27247 ( \35806_36106 , \35803_36103 , \35804_36104 , \35805_36105 );
and \U$27248 ( \35807_36107 , \35468_35768 , \35472_35772 );
and \U$27249 ( \35808_36108 , \35472_35772 , \35477_35777 );
and \U$27250 ( \35809_36109 , \35468_35768 , \35477_35777 );
or \U$27251 ( \35810_36110 , \35807_36107 , \35808_36108 , \35809_36109 );
xor \U$27252 ( \35811_36111 , \35806_36106 , \35810_36110 );
and \U$27253 ( \35812_36112 , \30500_30802 , \16333_16635 );
and \U$27254 ( \35813_36113 , \31752_32054 , \15999_16301 );
nor \U$27255 ( \35814_36114 , \35812_36112 , \35813_36113 );
xnor \U$27256 ( \35815_36115 , \35814_36114 , \16323_16625 );
not \U$27257 ( \35816_36116 , \35815_36115 );
xor \U$27258 ( \35817_36117 , \35811_36111 , \35816_36116 );
xor \U$27259 ( \35818_36118 , \35802_36102 , \35817_36117 );
xor \U$27260 ( \35819_36119 , \35793_36093 , \35818_36118 );
xor \U$27261 ( \35820_36120 , \35745_36045 , \35819_36119 );
and \U$27262 ( \35821_36121 , \35383_35683 , \35387_35687 );
and \U$27263 ( \35822_36122 , \35387_35687 , \35412_35712 );
and \U$27264 ( \35823_36123 , \35383_35683 , \35412_35712 );
or \U$27265 ( \35824_36124 , \35821_36121 , \35822_36122 , \35823_36123 );
and \U$27266 ( \35825_36125 , \35418_35718 , \35449_35749 );
and \U$27267 ( \35826_36126 , \35449_35749 , \35488_35788 );
and \U$27268 ( \35827_36127 , \35418_35718 , \35488_35788 );
or \U$27269 ( \35828_36128 , \35825_36125 , \35826_36126 , \35827_36127 );
xor \U$27270 ( \35829_36129 , \35824_36124 , \35828_36128 );
and \U$27271 ( \35830_36130 , \35422_35722 , \35436_35736 );
and \U$27272 ( \35831_36131 , \35436_35736 , \35448_35748 );
and \U$27273 ( \35832_36132 , \35422_35722 , \35448_35748 );
or \U$27274 ( \35833_36133 , \35830_36130 , \35831_36131 , \35832_36132 );
and \U$27275 ( \35834_36134 , \35464_35764 , \35478_35778 );
and \U$27276 ( \35835_36135 , \35478_35778 , \35487_35787 );
and \U$27277 ( \35836_36136 , \35464_35764 , \35487_35787 );
or \U$27278 ( \35837_36137 , \35834_36134 , \35835_36135 , \35836_36136 );
xor \U$27279 ( \35838_36138 , \35833_36133 , \35837_36137 );
and \U$27280 ( \35839_36139 , \35438_35738 , \35442_35742 );
and \U$27281 ( \35840_36140 , \35442_35742 , \35447_35747 );
and \U$27282 ( \35841_36141 , \35438_35738 , \35447_35747 );
or \U$27283 ( \35842_36142 , \35839_36139 , \35840_36140 , \35841_36141 );
and \U$27284 ( \35843_36143 , \35454_35754 , \35458_35758 );
and \U$27285 ( \35844_36144 , \35458_35758 , \35463_35763 );
and \U$27286 ( \35845_36145 , \35454_35754 , \35463_35763 );
or \U$27287 ( \35846_36146 , \35843_36143 , \35844_36144 , \35845_36145 );
xor \U$27288 ( \35847_36147 , \35842_36142 , \35846_36146 );
and \U$27289 ( \35848_36148 , \28782_29084 , \17791_18090 );
and \U$27290 ( \35849_36149 , \29966_30268 , \17353_17655 );
nor \U$27291 ( \35850_36150 , \35848_36148 , \35849_36149 );
xnor \U$27292 ( \35851_36151 , \35850_36150 , \17747_18046 );
and \U$27293 ( \35852_36152 , \22257_22556 , \23839_24138 );
and \U$27294 ( \35853_36153 , \23315_23617 , \23328_23630 );
nor \U$27295 ( \35854_36154 , \35852_36152 , \35853_36153 );
xnor \U$27296 ( \35855_36155 , \35854_36154 , \23845_24144 );
xor \U$27297 ( \35856_36156 , \35851_36151 , \35855_36155 );
and \U$27298 ( \35857_36157 , \14648_14950 , \32503_32802 );
xor \U$27299 ( \35858_36158 , \35856_36156 , \35857_36157 );
xor \U$27300 ( \35859_36159 , \35847_36147 , \35858_36158 );
xor \U$27301 ( \35860_36160 , \35838_36138 , \35859_36159 );
xor \U$27302 ( \35861_36161 , \35829_36129 , \35860_36160 );
xor \U$27303 ( \35862_36162 , \35820_36120 , \35861_36161 );
and \U$27304 ( \35863_36163 , \35370_35670 , \35374_35674 );
and \U$27305 ( \35864_36164 , \35374_35674 , \35490_35790 );
and \U$27306 ( \35865_36165 , \35370_35670 , \35490_35790 );
or \U$27307 ( \35866_36166 , \35863_36163 , \35864_36164 , \35865_36165 );
xor \U$27308 ( \35867_36167 , \35862_36162 , \35866_36166 );
and \U$27309 ( \35868_36168 , \35491_35791 , \35495_35795 );
and \U$27310 ( \35869_36169 , \35496_35796 , \35499_35799 );
or \U$27311 ( \35870_36170 , \35868_36168 , \35869_36169 );
xor \U$27312 ( \35871_36171 , \35867_36167 , \35870_36170 );
buf g9b96_GF_PartitionCandidate( \35872_36172_nG9b96 , \35871_36171 );
and \U$27313 ( \35873_36173 , \10402_10704 , \35872_36172_nG9b96 );
or \U$27314 ( \35874_36174 , \35741_36041 , \35873_36173 );
xor \U$27315 ( \35875_36175 , \10399_10703 , \35874_36174 );
buf \U$27316 ( \35876_36176 , \35875_36175 );
buf \U$27318 ( \35877_36177 , \35876_36176 );
xor \U$27319 ( \35878_36178 , \35740_36040 , \35877_36177 );
buf \U$27320 ( \35879_36179 , \35878_36178 );
and \U$27321 ( \35880_36180 , \35358_35658 , \35364_35664 );
and \U$27322 ( \35881_36181 , \35358_35658 , \35506_35806 );
and \U$27323 ( \35882_36182 , \35364_35664 , \35506_35806 );
or \U$27324 ( \35883_36183 , \35880_36180 , \35881_36181 , \35882_36182 );
buf \U$27325 ( \35884_36184 , \35883_36183 );
xor \U$27326 ( \35885_36185 , \35879_36179 , \35884_36184 );
and \U$27327 ( \35886_36186 , \35343_35643 , \35349_35649 );
and \U$27328 ( \35887_36187 , \35343_35643 , \35356_35656 );
and \U$27329 ( \35888_36188 , \35349_35649 , \35356_35656 );
or \U$27330 ( \35889_36189 , \35886_36186 , \35887_36187 , \35888_36188 );
buf \U$27331 ( \35890_36190 , \35889_36189 );
and \U$27333 ( \35891_36191 , \32617_32916 , \14682_14984_nG9bf6 );
or \U$27334 ( \35892_36192 , 1'b0 , \35891_36191 );
xor \U$27335 ( \35893_36193 , 1'b0 , \35892_36192 );
buf \U$27336 ( \35894_36194 , \35893_36193 );
buf \U$27338 ( \35895_36195 , \35894_36194 );
and \U$27339 ( \35896_36196 , \31989_31636 , \15074_15373_nG9bf3 );
and \U$27340 ( \35897_36197 , \31334_31633 , \16013_16315_nG9bf0 );
or \U$27341 ( \35898_36198 , \35896_36196 , \35897_36197 );
xor \U$27342 ( \35899_36199 , \31333_31632 , \35898_36198 );
buf \U$27343 ( \35900_36200 , \35899_36199 );
buf \U$27345 ( \35901_36201 , \35900_36200 );
xor \U$27346 ( \35902_36202 , \35895_36195 , \35901_36201 );
buf \U$27347 ( \35903_36203 , \35902_36202 );
and \U$27348 ( \35904_36204 , \35594_35894 , \35600_35900 );
buf \U$27349 ( \35905_36205 , \35904_36204 );
xor \U$27350 ( \35906_36206 , \35903_36203 , \35905_36205 );
and \U$27351 ( \35907_36207 , \30670_29853 , \16378_16680_nG9bed );
and \U$27352 ( \35908_36208 , \29551_29850 , \17363_17665_nG9bea );
or \U$27353 ( \35909_36209 , \35907_36207 , \35908_36208 );
xor \U$27354 ( \35910_36210 , \29550_29849 , \35909_36209 );
buf \U$27355 ( \35911_36211 , \35910_36210 );
buf \U$27357 ( \35912_36212 , \35911_36211 );
xor \U$27358 ( \35913_36213 , \35906_36206 , \35912_36212 );
buf \U$27359 ( \35914_36214 , \35913_36213 );
and \U$27360 ( \35915_36215 , \35602_35902 , \35604_35904 );
and \U$27361 ( \35916_36216 , \35602_35902 , \35611_35911 );
and \U$27362 ( \35917_36217 , \35604_35904 , \35611_35911 );
or \U$27363 ( \35918_36218 , \35915_36215 , \35916_36216 , \35917_36217 );
buf \U$27364 ( \35919_36219 , \35918_36218 );
xor \U$27365 ( \35920_36220 , \35914_36214 , \35919_36219 );
and \U$27366 ( \35921_36221 , \23495_23201 , \22330_22629_nG9bd5 );
and \U$27367 ( \35922_36222 , \22899_23198 , \23394_23696_nG9bd2 );
or \U$27368 ( \35923_36223 , \35921_36221 , \35922_36222 );
xor \U$27369 ( \35924_36224 , \22898_23197 , \35923_36223 );
buf \U$27370 ( \35925_36225 , \35924_36224 );
buf \U$27372 ( \35926_36226 , \35925_36225 );
xor \U$27373 ( \35927_36227 , \35920_36220 , \35926_36226 );
buf \U$27374 ( \35928_36228 , \35927_36227 );
xor \U$27375 ( \35929_36229 , \35890_36190 , \35928_36228 );
and \U$27376 ( \35930_36230 , \13431_13370 , \33313_33613_nG9bab );
and \U$27377 ( \35931_36231 , \13068_13367 , \33741_34041_nG9ba8 );
or \U$27378 ( \35932_36232 , \35930_36230 , \35931_36231 );
xor \U$27379 ( \35933_36233 , \13067_13366 , \35932_36232 );
buf \U$27380 ( \35934_36234 , \35933_36233 );
buf \U$27382 ( \35935_36235 , \35934_36234 );
xor \U$27383 ( \35936_36236 , \35929_36229 , \35935_36235 );
buf \U$27384 ( \35937_36237 , \35936_36236 );
xor \U$27385 ( \35938_36238 , \35885_36185 , \35937_36237 );
buf \U$27386 ( \35939_36239 , \35938_36238 );
and \U$27387 ( \35940_36240 , \35304_35604 , \35324_35624 );
and \U$27388 ( \35941_36241 , \35304_35604 , \35330_35630 );
and \U$27389 ( \35942_36242 , \35324_35624 , \35330_35630 );
or \U$27390 ( \35943_36243 , \35940_36240 , \35941_36241 , \35942_36242 );
buf \U$27391 ( \35944_36244 , \35943_36243 );
xor \U$27392 ( \35945_36245 , \35939_36239 , \35944_36244 );
and \U$27393 ( \35946_36246 , \35589_35889 , \35613_35913 );
and \U$27394 ( \35947_36247 , \35589_35889 , \35620_35920 );
and \U$27395 ( \35948_36248 , \35613_35913 , \35620_35920 );
or \U$27396 ( \35949_36249 , \35946_36246 , \35947_36247 , \35948_36248 );
buf \U$27397 ( \35950_36250 , \35949_36249 );
and \U$27398 ( \35951_36251 , \17437_17297 , \28877_29179_nG9bbd );
and \U$27399 ( \35952_36252 , \16995_17294 , \30064_30366_nG9bba );
or \U$27400 ( \35953_36253 , \35951_36251 , \35952_36252 );
xor \U$27401 ( \35954_36254 , \16994_17293 , \35953_36253 );
buf \U$27402 ( \35955_36255 , \35954_36254 );
buf \U$27404 ( \35956_36256 , \35955_36255 );
xor \U$27405 ( \35957_36257 , \35950_36250 , \35956_36256 );
and \U$27406 ( \35958_36258 , \14710_14631 , \32589_32888_nG9bb1 );
and \U$27407 ( \35959_36259 , \14329_14628 , \32881_33181_nG9bae );
or \U$27408 ( \35960_36260 , \35958_36258 , \35959_36259 );
xor \U$27409 ( \35961_36261 , \14328_14627 , \35960_36260 );
buf \U$27410 ( \35962_36262 , \35961_36261 );
buf \U$27412 ( \35963_36263 , \35962_36262 );
xor \U$27413 ( \35964_36264 , \35957_36257 , \35963_36263 );
buf \U$27414 ( \35965_36265 , \35964_36264 );
and \U$27415 ( \35966_36266 , \35309_35609 , \35315_35615 );
and \U$27416 ( \35967_36267 , \35309_35609 , \35322_35622 );
and \U$27417 ( \35968_36268 , \35315_35615 , \35322_35622 );
or \U$27418 ( \35969_36269 , \35966_36266 , \35967_36267 , \35968_36268 );
buf \U$27419 ( \35970_36270 , \35969_36269 );
xor \U$27420 ( \35971_36271 , \35965_36265 , \35970_36270 );
and \U$27421 ( \35972_36272 , \28946_28118 , \17808_18107_nG9be7 );
and \U$27422 ( \35973_36273 , \27816_28115 , \18789_19091_nG9be4 );
or \U$27423 ( \35974_36274 , \35972_36272 , \35973_36273 );
xor \U$27424 ( \35975_36275 , \27815_28114 , \35974_36274 );
buf \U$27425 ( \35976_36276 , \35975_36275 );
buf \U$27427 ( \35977_36277 , \35976_36276 );
and \U$27428 ( \35978_36278 , \27141_26431 , \19287_19586_nG9be1 );
and \U$27429 ( \35979_36279 , \26129_26428 , \20306_20608_nG9bde );
or \U$27430 ( \35980_36280 , \35978_36278 , \35979_36279 );
xor \U$27431 ( \35981_36281 , \26128_26427 , \35980_36280 );
buf \U$27432 ( \35982_36282 , \35981_36281 );
buf \U$27434 ( \35983_36283 , \35982_36282 );
xor \U$27435 ( \35984_36284 , \35977_36277 , \35983_36283 );
and \U$27436 ( \35985_36285 , \25044_24792 , \20787_21086_nG9bdb );
and \U$27437 ( \35986_36286 , \24490_24789 , \21827_22129_nG9bd8 );
or \U$27438 ( \35987_36287 , \35985_36285 , \35986_36286 );
xor \U$27439 ( \35988_36288 , \24489_24788 , \35987_36287 );
buf \U$27440 ( \35989_36289 , \35988_36288 );
buf \U$27442 ( \35990_36290 , \35989_36289 );
xor \U$27443 ( \35991_36291 , \35984_36284 , \35990_36290 );
buf \U$27444 ( \35992_36292 , \35991_36291 );
and \U$27445 ( \35993_36293 , \20353_20155 , \25561_25860_nG9bc9 );
and \U$27446 ( \35994_36294 , \19853_20152 , \26585_26887_nG9bc6 );
or \U$27447 ( \35995_36295 , \35993_36293 , \35994_36294 );
xor \U$27448 ( \35996_36296 , \19852_20151 , \35995_36295 );
buf \U$27449 ( \35997_36297 , \35996_36296 );
buf \U$27451 ( \35998_36298 , \35997_36297 );
xor \U$27452 ( \35999_36299 , \35992_36292 , \35998_36298 );
and \U$27453 ( \36000_36300 , \16405_15940 , \30638_30940_nG9bb7 );
and \U$27454 ( \36001_36301 , \15638_15937 , \31877_32179_nG9bb4 );
or \U$27455 ( \36002_36302 , \36000_36300 , \36001_36301 );
xor \U$27456 ( \36003_36303 , \15637_15936 , \36002_36302 );
buf \U$27457 ( \36004_36304 , \36003_36303 );
buf \U$27459 ( \36005_36305 , \36004_36304 );
xor \U$27460 ( \36006_36306 , \35999_36299 , \36005_36305 );
buf \U$27461 ( \36007_36307 , \36006_36306 );
xor \U$27462 ( \36008_36308 , \35971_36271 , \36007_36307 );
buf \U$27463 ( \36009_36309 , \36008_36308 );
xor \U$27464 ( \36010_36310 , \35945_36245 , \36009_36309 );
buf \U$27465 ( \36011_36311 , \36010_36310 );
xor \U$27466 ( \36012_36312 , \35728_36028 , \36011_36311 );
and \U$27467 ( \36013_36313 , \35662_35962 , \36012_36312 );
and \U$27469 ( \36014_36314 , \35656_35956 , \35661_35961 );
or \U$27471 ( \36015_36315 , 1'b0 , \36014_36314 , 1'b0 );
xor \U$27472 ( \36016_36316 , \36013_36313 , \36015_36315 );
and \U$27474 ( \36017_36317 , \35649_35949 , \35655_35955 );
and \U$27475 ( \36018_36318 , \35651_35951 , \35655_35955 );
or \U$27476 ( \36019_36319 , 1'b0 , \36017_36317 , \36018_36318 );
xor \U$27477 ( \36020_36320 , \36016_36316 , \36019_36319 );
xor \U$27484 ( \36021_36321 , \36020_36320 , 1'b0 );
and \U$27485 ( \36022_36322 , \35722_36022 , \35727_36027 );
and \U$27486 ( \36023_36323 , \35722_36022 , \36011_36311 );
and \U$27487 ( \36024_36324 , \35727_36027 , \36011_36311 );
or \U$27488 ( \36025_36325 , \36022_36322 , \36023_36323 , \36024_36324 );
xor \U$27489 ( \36026_36326 , \36021_36321 , \36025_36325 );
and \U$27490 ( \36027_36327 , \35667_35967 , \35672_35972 );
and \U$27491 ( \36028_36328 , \35667_35967 , \35720_36020 );
and \U$27492 ( \36029_36329 , \35672_35972 , \35720_36020 );
or \U$27493 ( \36030_36330 , \36027_36327 , \36028_36328 , \36029_36329 );
buf \U$27494 ( \36031_36331 , \36030_36330 );
and \U$27495 ( \36032_36332 , \35939_36239 , \35944_36244 );
and \U$27496 ( \36033_36333 , \35939_36239 , \36009_36309 );
and \U$27497 ( \36034_36334 , \35944_36244 , \36009_36309 );
or \U$27498 ( \36035_36335 , \36032_36332 , \36033_36333 , \36034_36334 );
buf \U$27499 ( \36036_36336 , \36035_36335 );
and \U$27500 ( \36037_36337 , \35914_36214 , \35919_36219 );
and \U$27501 ( \36038_36338 , \35914_36214 , \35926_36226 );
and \U$27502 ( \36039_36339 , \35919_36219 , \35926_36226 );
or \U$27503 ( \36040_36340 , \36037_36337 , \36038_36338 , \36039_36339 );
buf \U$27504 ( \36041_36341 , \36040_36340 );
and \U$27505 ( \36042_36342 , \35903_36203 , \35905_36205 );
and \U$27506 ( \36043_36343 , \35903_36203 , \35912_36212 );
and \U$27507 ( \36044_36344 , \35905_36205 , \35912_36212 );
or \U$27508 ( \36045_36345 , \36042_36342 , \36043_36343 , \36044_36344 );
buf \U$27509 ( \36046_36346 , \36045_36345 );
and \U$27510 ( \36047_36347 , \28946_28118 , \18789_19091_nG9be4 );
and \U$27511 ( \36048_36348 , \27816_28115 , \19287_19586_nG9be1 );
or \U$27512 ( \36049_36349 , \36047_36347 , \36048_36348 );
xor \U$27513 ( \36050_36350 , \27815_28114 , \36049_36349 );
buf \U$27514 ( \36051_36351 , \36050_36350 );
buf \U$27516 ( \36052_36352 , \36051_36351 );
xor \U$27517 ( \36053_36353 , \36046_36346 , \36052_36352 );
and \U$27518 ( \36054_36354 , \27141_26431 , \20306_20608_nG9bde );
and \U$27519 ( \36055_36355 , \26129_26428 , \20787_21086_nG9bdb );
or \U$27520 ( \36056_36356 , \36054_36354 , \36055_36355 );
xor \U$27521 ( \36057_36357 , \26128_26427 , \36056_36356 );
buf \U$27522 ( \36058_36358 , \36057_36357 );
buf \U$27524 ( \36059_36359 , \36058_36358 );
xor \U$27525 ( \36060_36360 , \36053_36353 , \36059_36359 );
buf \U$27526 ( \36061_36361 , \36060_36360 );
xor \U$27527 ( \36062_36362 , \36041_36341 , \36061_36361 );
and \U$27528 ( \36063_36363 , \18908_18702 , \28300_28602_nG9bc0 );
and \U$27529 ( \36064_36364 , \18400_18699 , \28877_29179_nG9bbd );
or \U$27530 ( \36065_36365 , \36063_36363 , \36064_36364 );
xor \U$27531 ( \36066_36366 , \18399_18698 , \36065_36365 );
buf \U$27532 ( \36067_36367 , \36066_36366 );
buf \U$27534 ( \36068_36368 , \36067_36367 );
xor \U$27535 ( \36069_36369 , \36062_36362 , \36068_36368 );
buf \U$27536 ( \36070_36370 , \36069_36369 );
and \U$27537 ( \36071_36371 , \35992_36292 , \35998_36298 );
and \U$27538 ( \36072_36372 , \35992_36292 , \36005_36305 );
and \U$27539 ( \36073_36373 , \35998_36298 , \36005_36305 );
or \U$27540 ( \36074_36374 , \36071_36371 , \36072_36372 , \36073_36373 );
buf \U$27541 ( \36075_36375 , \36074_36374 );
xor \U$27542 ( \36076_36376 , \36070_36370 , \36075_36375 );
and \U$27544 ( \36077_36377 , \32617_32916 , \15074_15373_nG9bf3 );
or \U$27545 ( \36078_36378 , 1'b0 , \36077_36377 );
xor \U$27546 ( \36079_36379 , 1'b0 , \36078_36378 );
buf \U$27547 ( \36080_36380 , \36079_36379 );
buf \U$27549 ( \36081_36381 , \36080_36380 );
and \U$27550 ( \36082_36382 , \31989_31636 , \16013_16315_nG9bf0 );
and \U$27551 ( \36083_36383 , \31334_31633 , \16378_16680_nG9bed );
or \U$27552 ( \36084_36384 , \36082_36382 , \36083_36383 );
xor \U$27553 ( \36085_36385 , \31333_31632 , \36084_36384 );
buf \U$27554 ( \36086_36386 , \36085_36385 );
buf \U$27556 ( \36087_36387 , \36086_36386 );
xor \U$27557 ( \36088_36388 , \36081_36381 , \36087_36387 );
buf \U$27558 ( \36089_36389 , \36088_36388 );
and \U$27559 ( \36090_36390 , \35895_36195 , \35901_36201 );
buf \U$27560 ( \36091_36391 , \36090_36390 );
xor \U$27561 ( \36092_36392 , \36089_36389 , \36091_36391 );
and \U$27562 ( \36093_36393 , \30670_29853 , \17363_17665_nG9bea );
and \U$27563 ( \36094_36394 , \29551_29850 , \17808_18107_nG9be7 );
or \U$27564 ( \36095_36395 , \36093_36393 , \36094_36394 );
xor \U$27565 ( \36096_36396 , \29550_29849 , \36095_36395 );
buf \U$27566 ( \36097_36397 , \36096_36396 );
buf \U$27568 ( \36098_36398 , \36097_36397 );
xor \U$27569 ( \36099_36399 , \36092_36392 , \36098_36398 );
buf \U$27570 ( \36100_36400 , \36099_36399 );
and \U$27571 ( \36101_36401 , \21908_21658 , \24996_25298_nG9bcc );
and \U$27572 ( \36102_36402 , \21356_21655 , \25561_25860_nG9bc9 );
or \U$27573 ( \36103_36403 , \36101_36401 , \36102_36402 );
xor \U$27574 ( \36104_36404 , \21355_21654 , \36103_36403 );
buf \U$27575 ( \36105_36405 , \36104_36404 );
buf \U$27577 ( \36106_36406 , \36105_36405 );
xor \U$27578 ( \36107_36407 , \36100_36400 , \36106_36406 );
and \U$27579 ( \36108_36408 , \20353_20155 , \26585_26887_nG9bc6 );
and \U$27580 ( \36109_36409 , \19853_20152 , \27114_27416_nG9bc3 );
or \U$27581 ( \36110_36410 , \36108_36408 , \36109_36409 );
xor \U$27582 ( \36111_36411 , \19852_20151 , \36110_36410 );
buf \U$27583 ( \36112_36412 , \36111_36411 );
buf \U$27585 ( \36113_36413 , \36112_36412 );
xor \U$27586 ( \36114_36414 , \36107_36407 , \36113_36413 );
buf \U$27587 ( \36115_36415 , \36114_36414 );
xor \U$27588 ( \36116_36416 , \36076_36376 , \36115_36415 );
buf \U$27589 ( \36117_36417 , \36116_36416 );
and \U$27590 ( \36118_36418 , \35683_35983 , \35703_36003 );
and \U$27591 ( \36119_36419 , \35683_35983 , \35710_36010 );
and \U$27592 ( \36120_36420 , \35703_36003 , \35710_36010 );
or \U$27593 ( \36121_36421 , \36118_36418 , \36119_36419 , \36120_36420 );
buf \U$27594 ( \36122_36422 , \36121_36421 );
xor \U$27595 ( \36123_36423 , \36117_36417 , \36122_36422 );
and \U$27596 ( \36124_36424 , \35965_36265 , \35970_36270 );
and \U$27597 ( \36125_36425 , \35965_36265 , \36007_36307 );
and \U$27598 ( \36126_36426 , \35970_36270 , \36007_36307 );
or \U$27599 ( \36127_36427 , \36124_36424 , \36125_36425 , \36126_36426 );
buf \U$27600 ( \36128_36428 , \36127_36427 );
xor \U$27601 ( \36129_36429 , \36123_36423 , \36128_36428 );
buf \U$27602 ( \36130_36430 , \36129_36429 );
xor \U$27603 ( \36131_36431 , \36036_36336 , \36130_36430 );
and \U$27604 ( \36132_36432 , \35733_36033 , \35739_36039 );
and \U$27605 ( \36133_36433 , \35733_36033 , \35877_36177 );
and \U$27606 ( \36134_36434 , \35739_36039 , \35877_36177 );
or \U$27607 ( \36135_36435 , \36132_36432 , \36133_36433 , \36134_36434 );
buf \U$27608 ( \36136_36436 , \36135_36435 );
and \U$27609 ( \36137_36437 , \35977_36277 , \35983_36283 );
and \U$27610 ( \36138_36438 , \35977_36277 , \35990_36290 );
and \U$27611 ( \36139_36439 , \35983_36283 , \35990_36290 );
or \U$27612 ( \36140_36440 , \36137_36437 , \36138_36438 , \36139_36439 );
buf \U$27613 ( \36141_36441 , \36140_36440 );
and \U$27614 ( \36142_36442 , \25044_24792 , \21827_22129_nG9bd8 );
and \U$27615 ( \36143_36443 , \24490_24789 , \22330_22629_nG9bd5 );
or \U$27616 ( \36144_36444 , \36142_36442 , \36143_36443 );
xor \U$27617 ( \36145_36445 , \24489_24788 , \36144_36444 );
buf \U$27618 ( \36146_36446 , \36145_36445 );
buf \U$27620 ( \36147_36447 , \36146_36446 );
xor \U$27621 ( \36148_36448 , \36141_36441 , \36147_36447 );
and \U$27622 ( \36149_36449 , \23495_23201 , \23394_23696_nG9bd2 );
and \U$27623 ( \36150_36450 , \22899_23198 , \23927_24226_nG9bcf );
or \U$27624 ( \36151_36451 , \36149_36449 , \36150_36450 );
xor \U$27625 ( \36152_36452 , \22898_23197 , \36151_36451 );
buf \U$27626 ( \36153_36453 , \36152_36452 );
buf \U$27628 ( \36154_36454 , \36153_36453 );
xor \U$27629 ( \36155_36455 , \36148_36448 , \36154_36454 );
buf \U$27630 ( \36156_36456 , \36155_36455 );
and \U$27631 ( \36157_36457 , \12183_12157 , \34343_34643_nG9ba2 );
and \U$27632 ( \36158_36458 , \11855_12154 , \34794_35094_nG9b9f );
or \U$27633 ( \36159_36459 , \36157_36457 , \36158_36458 );
xor \U$27634 ( \36160_36460 , \11854_12153 , \36159_36459 );
buf \U$27635 ( \36161_36461 , \36160_36460 );
buf \U$27637 ( \36162_36462 , \36161_36461 );
xor \U$27638 ( \36163_36463 , \36156_36456 , \36162_36462 );
and \U$27639 ( \36164_36464 , \10411_10707 , \35872_36172_nG9b96 );
and \U$27640 ( \36165_36465 , \35824_36124 , \35828_36128 );
and \U$27641 ( \36166_36466 , \35828_36128 , \35860_36160 );
and \U$27642 ( \36167_36467 , \35824_36124 , \35860_36160 );
or \U$27643 ( \36168_36468 , \36165_36465 , \36166_36466 , \36167_36467 );
and \U$27644 ( \36169_36469 , \35797_36097 , \35801_36101 );
and \U$27645 ( \36170_36470 , \35801_36101 , \35817_36117 );
and \U$27646 ( \36171_36471 , \35797_36097 , \35817_36117 );
or \U$27647 ( \36172_36472 , \36169_36469 , \36170_36470 , \36171_36471 );
and \U$27648 ( \36173_36473 , \26527_26829 , \20706_21005 );
and \U$27649 ( \36174_36474 , \27011_27313 , \20255_20557 );
nor \U$27650 ( \36175_36475 , \36173_36473 , \36174_36474 );
xnor \U$27651 ( \36176_36476 , \36175_36475 , \20712_21011 );
and \U$27652 ( \36177_36477 , \21788_22090 , \25527_25826 );
and \U$27653 ( \36178_36478 , \22257_22556 , \24962_25264 );
nor \U$27654 ( \36179_36479 , \36177_36477 , \36178_36478 );
xnor \U$27655 ( \36180_36480 , \36179_36479 , \25474_25773 );
xor \U$27656 ( \36181_36481 , \36176_36476 , \36180_36480 );
and \U$27657 ( \36182_36482 , \20242_20544 , \27095_27397 );
and \U$27658 ( \36183_36483 , \20734_21033 , \26505_26807 );
nor \U$27659 ( \36184_36484 , \36182_36482 , \36183_36483 );
xnor \U$27660 ( \36185_36485 , \36184_36484 , \26993_27295 );
xor \U$27661 ( \36186_36486 , \36181_36481 , \36185_36485 );
not \U$27662 ( \36187_36487 , \15043_15342 );
and \U$27663 ( \36188_36488 , \31752_32054 , \16333_16635 );
and \U$27664 ( \36189_36489 , \32495_32794 , \15999_16301 );
nor \U$27665 ( \36190_36490 , \36188_36488 , \36189_36489 );
xnor \U$27666 ( \36191_36491 , \36190_36490 , \16323_16625 );
xor \U$27667 ( \36192_36492 , \36187_36487 , \36191_36491 );
and \U$27668 ( \36193_36493 , \28232_28534 , \19235_19534 );
and \U$27669 ( \36194_36494 , \28782_29084 , \18743_19045 );
nor \U$27670 ( \36195_36495 , \36193_36493 , \36194_36494 );
xnor \U$27671 ( \36196_36496 , \36195_36495 , \19241_19540 );
xor \U$27672 ( \36197_36497 , \36192_36492 , \36196_36496 );
xor \U$27673 ( \36198_36498 , \36186_36486 , \36197_36497 );
and \U$27674 ( \36199_36499 , \29966_30268 , \17791_18090 );
and \U$27675 ( \36200_36500 , \30500_30802 , \17353_17655 );
nor \U$27676 ( \36201_36501 , \36199_36499 , \36200_36500 );
xnor \U$27677 ( \36202_36502 , \36201_36501 , \17747_18046 );
and \U$27678 ( \36203_36503 , \18730_19032 , \28768_29070 );
and \U$27679 ( \36204_36504 , \19259_19558 , \28224_28526 );
nor \U$27680 ( \36205_36505 , \36203_36503 , \36204_36504 );
xnor \U$27681 ( \36206_36506 , \36205_36505 , \28774_29076 );
xor \U$27682 ( \36207_36507 , \36202_36502 , \36206_36506 );
and \U$27683 ( \36208_36508 , \17325_17627 , \30521_30823 );
and \U$27684 ( \36209_36509 , \17736_18035 , \29944_30246 );
nor \U$27685 ( \36210_36510 , \36208_36508 , \36209_36509 );
xnor \U$27686 ( \36211_36511 , \36210_36510 , \30511_30813 );
xor \U$27687 ( \36212_36512 , \36207_36507 , \36211_36511 );
xor \U$27688 ( \36213_36513 , \36198_36498 , \36212_36512 );
xor \U$27689 ( \36214_36514 , \36172_36472 , \36213_36513 );
and \U$27690 ( \36215_36515 , \35806_36106 , \35810_36110 );
and \U$27691 ( \36216_36516 , \35810_36110 , \35816_36116 );
and \U$27692 ( \36217_36517 , \35806_36106 , \35816_36116 );
or \U$27693 ( \36218_36518 , \36215_36515 , \36216_36516 , \36217_36517 );
and \U$27694 ( \36219_36519 , \24970_25272 , \22243_22542 );
and \U$27695 ( \36220_36520 , \25516_25815 , \21801_22103 );
nor \U$27696 ( \36221_36521 , \36219_36519 , \36220_36520 );
xnor \U$27697 ( \36222_36522 , \36221_36521 , \22249_22548 );
and \U$27698 ( \36223_36523 , \15965_16267 , \32555_32854 );
and \U$27699 ( \36224_36524 , \16353_16655 , \31765_32067 );
nor \U$27700 ( \36225_36525 , \36223_36523 , \36224_36524 );
xnor \U$27701 ( \36226_36526 , \36225_36525 , \32506_32805 );
xor \U$27702 ( \36227_36527 , \36222_36522 , \36226_36526 );
and \U$27703 ( \36228_36528 , \15022_15321 , \32503_32802 );
xor \U$27704 ( \36229_36529 , \36227_36527 , \36228_36528 );
xor \U$27705 ( \36230_36530 , \36218_36518 , \36229_36529 );
and \U$27706 ( \36231_36531 , \35781_36081 , \35785_36085 );
and \U$27707 ( \36232_36532 , \35785_36085 , \35790_36090 );
and \U$27708 ( \36233_36533 , \35781_36081 , \35790_36090 );
or \U$27709 ( \36234_36534 , \36231_36531 , \36232_36532 , \36233_36533 );
buf \U$27710 ( \36235_36535 , \35815_36115 );
xor \U$27711 ( \36236_36536 , \36234_36534 , \36235_36535 );
and \U$27712 ( \36237_36537 , \23315_23617 , \23839_24138 );
and \U$27713 ( \36238_36538 , \23900_24199 , \23328_23630 );
nor \U$27714 ( \36239_36539 , \36237_36537 , \36238_36538 );
xnor \U$27715 ( \36240_36540 , \36239_36539 , \23845_24144 );
xor \U$27716 ( \36241_36541 , \36236_36536 , \36240_36540 );
xor \U$27717 ( \36242_36542 , \36230_36530 , \36241_36541 );
xor \U$27718 ( \36243_36543 , \36214_36514 , \36242_36542 );
xor \U$27719 ( \36244_36544 , \36168_36468 , \36243_36543 );
and \U$27720 ( \36245_36545 , \35833_36133 , \35837_36137 );
and \U$27721 ( \36246_36546 , \35837_36137 , \35859_36159 );
and \U$27722 ( \36247_36547 , \35833_36133 , \35859_36159 );
or \U$27723 ( \36248_36548 , \36245_36545 , \36246_36546 , \36247_36547 );
and \U$27724 ( \36249_36549 , \35749_36049 , \35792_36092 );
and \U$27725 ( \36250_36550 , \35792_36092 , \35818_36118 );
and \U$27726 ( \36251_36551 , \35749_36049 , \35818_36118 );
or \U$27727 ( \36252_36552 , \36249_36549 , \36250_36550 , \36251_36551 );
xor \U$27728 ( \36253_36553 , \36248_36548 , \36252_36552 );
and \U$27729 ( \36254_36554 , \35842_36142 , \35846_36146 );
and \U$27730 ( \36255_36555 , \35846_36146 , \35858_36158 );
and \U$27731 ( \36256_36556 , \35842_36142 , \35858_36158 );
or \U$27732 ( \36257_36557 , \36254_36554 , \36255_36555 , \36256_36556 );
and \U$27733 ( \36258_36558 , \35763_36063 , \35776_36076 );
and \U$27734 ( \36259_36559 , \35776_36076 , \35791_36091 );
and \U$27735 ( \36260_36560 , \35763_36063 , \35791_36091 );
or \U$27736 ( \36261_36561 , \36258_36558 , \36259_36559 , \36260_36560 );
xor \U$27737 ( \36262_36562 , \36257_36557 , \36261_36561 );
and \U$27738 ( \36263_36563 , \35851_36151 , \35855_36155 );
and \U$27739 ( \36264_36564 , \35855_36155 , \35857_36157 );
and \U$27740 ( \36265_36565 , \35851_36151 , \35857_36157 );
or \U$27741 ( \36266_36566 , \36263_36563 , \36264_36564 , \36265_36565 );
and \U$27742 ( \36267_36567 , \35753_36053 , \35757_36057 );
and \U$27743 ( \36268_36568 , \35757_36057 , \35762_36062 );
and \U$27744 ( \36269_36569 , \35753_36053 , \35762_36062 );
or \U$27745 ( \36270_36570 , \36267_36567 , \36268_36568 , \36269_36569 );
xor \U$27746 ( \36271_36571 , \36266_36566 , \36270_36570 );
and \U$27747 ( \36272_36572 , \35766_36066 , \35770_36070 );
and \U$27748 ( \36273_36573 , \35770_36070 , \35775_36075 );
and \U$27749 ( \36274_36574 , \35766_36066 , \35775_36075 );
or \U$27750 ( \36275_36575 , \36272_36572 , \36273_36573 , \36274_36574 );
xor \U$27751 ( \36276_36576 , \36271_36571 , \36275_36575 );
xor \U$27752 ( \36277_36577 , \36262_36562 , \36276_36576 );
xor \U$27753 ( \36278_36578 , \36253_36553 , \36277_36577 );
xor \U$27754 ( \36279_36579 , \36244_36544 , \36278_36578 );
and \U$27755 ( \36280_36580 , \35745_36045 , \35819_36119 );
and \U$27756 ( \36281_36581 , \35819_36119 , \35861_36161 );
and \U$27757 ( \36282_36582 , \35745_36045 , \35861_36161 );
or \U$27758 ( \36283_36583 , \36280_36580 , \36281_36581 , \36282_36582 );
xor \U$27759 ( \36284_36584 , \36279_36579 , \36283_36583 );
and \U$27760 ( \36285_36585 , \35862_36162 , \35866_36166 );
and \U$27761 ( \36286_36586 , \35867_36167 , \35870_36170 );
or \U$27762 ( \36287_36587 , \36285_36585 , \36286_36586 );
xor \U$27763 ( \36288_36588 , \36284_36584 , \36287_36587 );
buf g9b93_GF_PartitionCandidate( \36289_36589_nG9b93 , \36288_36588 );
and \U$27764 ( \36290_36590 , \10402_10704 , \36289_36589_nG9b93 );
or \U$27765 ( \36291_36591 , \36164_36464 , \36290_36590 );
xor \U$27766 ( \36292_36592 , \10399_10703 , \36291_36591 );
buf \U$27767 ( \36293_36593 , \36292_36592 );
buf \U$27769 ( \36294_36594 , \36293_36593 );
xor \U$27770 ( \36295_36595 , \36163_36463 , \36294_36594 );
buf \U$27771 ( \36296_36596 , \36295_36595 );
xor \U$27772 ( \36297_36597 , \36136_36436 , \36296_36596 );
and \U$27773 ( \36298_36598 , \35688_35988 , \35694_35994 );
and \U$27774 ( \36299_36599 , \35688_35988 , \35701_36001 );
and \U$27775 ( \36300_36600 , \35694_35994 , \35701_36001 );
or \U$27776 ( \36301_36601 , \36298_36598 , \36299_36599 , \36300_36600 );
buf \U$27777 ( \36302_36602 , \36301_36601 );
and \U$27778 ( \36303_36603 , \13431_13370 , \33741_34041_nG9ba8 );
and \U$27779 ( \36304_36604 , \13068_13367 , \33994_34294_nG9ba5 );
or \U$27780 ( \36305_36605 , \36303_36603 , \36304_36604 );
xor \U$27781 ( \36306_36606 , \13067_13366 , \36305_36605 );
buf \U$27782 ( \36307_36607 , \36306_36606 );
buf \U$27784 ( \36308_36608 , \36307_36607 );
xor \U$27785 ( \36309_36609 , \36302_36602 , \36308_36608 );
and \U$27786 ( \36310_36610 , \10996_10421 , \35270_35570_nG9b9c );
and \U$27787 ( \36311_36611 , \10119_10418 , \35501_35801_nG9b99 );
or \U$27788 ( \36312_36612 , \36310_36610 , \36311_36611 );
xor \U$27789 ( \36313_36613 , \10118_10417 , \36312_36612 );
buf \U$27790 ( \36314_36614 , \36313_36613 );
buf \U$27792 ( \36315_36615 , \36314_36614 );
xor \U$27793 ( \36316_36616 , \36309_36609 , \36315_36615 );
buf \U$27794 ( \36317_36617 , \36316_36616 );
xor \U$27795 ( \36318_36618 , \36297_36597 , \36317_36617 );
buf \U$27796 ( \36319_36619 , \36318_36618 );
xor \U$27797 ( \36320_36620 , \36131_36431 , \36319_36619 );
buf \U$27798 ( \36321_36621 , \36320_36620 );
xor \U$27799 ( \36322_36622 , \36031_36331 , \36321_36621 );
and \U$27800 ( \36323_36623 , \35678_35978 , \35712_36012 );
and \U$27801 ( \36324_36624 , \35678_35978 , \35718_36018 );
and \U$27802 ( \36325_36625 , \35712_36012 , \35718_36018 );
or \U$27803 ( \36326_36626 , \36323_36623 , \36324_36624 , \36325_36625 );
buf \U$27804 ( \36327_36627 , \36326_36626 );
and \U$27805 ( \36328_36628 , \35879_36179 , \35884_36184 );
and \U$27806 ( \36329_36629 , \35879_36179 , \35937_36237 );
and \U$27807 ( \36330_36630 , \35884_36184 , \35937_36237 );
or \U$27808 ( \36331_36631 , \36328_36628 , \36329_36629 , \36330_36630 );
buf \U$27809 ( \36332_36632 , \36331_36631 );
xor \U$27810 ( \36333_36633 , \36327_36627 , \36332_36632 );
and \U$27811 ( \36334_36634 , \17437_17297 , \30064_30366_nG9bba );
and \U$27812 ( \36335_36635 , \16995_17294 , \30638_30940_nG9bb7 );
or \U$27813 ( \36336_36636 , \36334_36634 , \36335_36635 );
xor \U$27814 ( \36337_36637 , \16994_17293 , \36336_36636 );
buf \U$27815 ( \36338_36638 , \36337_36637 );
buf \U$27817 ( \36339_36639 , \36338_36638 );
and \U$27818 ( \36340_36640 , \16405_15940 , \31877_32179_nG9bb4 );
and \U$27819 ( \36341_36641 , \15638_15937 , \32589_32888_nG9bb1 );
or \U$27820 ( \36342_36642 , \36340_36640 , \36341_36641 );
xor \U$27821 ( \36343_36643 , \15637_15936 , \36342_36642 );
buf \U$27822 ( \36344_36644 , \36343_36643 );
buf \U$27824 ( \36345_36645 , \36344_36644 );
xor \U$27825 ( \36346_36646 , \36339_36639 , \36345_36645 );
and \U$27826 ( \36347_36647 , \14710_14631 , \32881_33181_nG9bae );
and \U$27827 ( \36348_36648 , \14329_14628 , \33313_33613_nG9bab );
or \U$27828 ( \36349_36649 , \36347_36647 , \36348_36648 );
xor \U$27829 ( \36350_36650 , \14328_14627 , \36349_36649 );
buf \U$27830 ( \36351_36651 , \36350_36650 );
buf \U$27832 ( \36352_36652 , \36351_36651 );
xor \U$27833 ( \36353_36653 , \36346_36646 , \36352_36652 );
buf \U$27834 ( \36354_36654 , \36353_36653 );
and \U$27835 ( \36355_36655 , \35890_36190 , \35928_36228 );
and \U$27836 ( \36356_36656 , \35890_36190 , \35935_36235 );
and \U$27837 ( \36357_36657 , \35928_36228 , \35935_36235 );
or \U$27838 ( \36358_36658 , \36355_36655 , \36356_36656 , \36357_36657 );
buf \U$27839 ( \36359_36659 , \36358_36658 );
xor \U$27840 ( \36360_36660 , \36354_36654 , \36359_36659 );
and \U$27841 ( \36361_36661 , \35950_36250 , \35956_36256 );
and \U$27842 ( \36362_36662 , \35950_36250 , \35963_36263 );
and \U$27843 ( \36363_36663 , \35956_36256 , \35963_36263 );
or \U$27844 ( \36364_36664 , \36361_36661 , \36362_36662 , \36363_36663 );
buf \U$27845 ( \36365_36665 , \36364_36664 );
xor \U$27846 ( \36366_36666 , \36360_36660 , \36365_36665 );
buf \U$27847 ( \36367_36667 , \36366_36666 );
xor \U$27848 ( \36368_36668 , \36333_36633 , \36367_36667 );
buf \U$27849 ( \36369_36669 , \36368_36668 );
xor \U$27850 ( \36370_36670 , \36322_36622 , \36369_36669 );
and \U$27851 ( \36371_36671 , \36026_36326 , \36370_36670 );
and \U$27853 ( \36372_36672 , \36020_36320 , \36025_36325 );
or \U$27855 ( \36373_36673 , 1'b0 , \36372_36672 , 1'b0 );
xor \U$27856 ( \36374_36674 , \36371_36671 , \36373_36673 );
and \U$27858 ( \36375_36675 , \36013_36313 , \36019_36319 );
and \U$27859 ( \36376_36676 , \36015_36315 , \36019_36319 );
or \U$27860 ( \36377_36677 , 1'b0 , \36375_36675 , \36376_36676 );
xor \U$27861 ( \36378_36678 , \36374_36674 , \36377_36677 );
xor \U$27868 ( \36379_36679 , \36378_36678 , 1'b0 );
and \U$27869 ( \36380_36680 , \36031_36331 , \36321_36621 );
and \U$27870 ( \36381_36681 , \36031_36331 , \36369_36669 );
and \U$27871 ( \36382_36682 , \36321_36621 , \36369_36669 );
or \U$27872 ( \36383_36683 , \36380_36680 , \36381_36681 , \36382_36682 );
xor \U$27873 ( \36384_36684 , \36379_36679 , \36383_36683 );
and \U$27874 ( \36385_36685 , \36036_36336 , \36130_36430 );
and \U$27875 ( \36386_36686 , \36036_36336 , \36319_36619 );
and \U$27876 ( \36387_36687 , \36130_36430 , \36319_36619 );
or \U$27877 ( \36388_36688 , \36385_36685 , \36386_36686 , \36387_36687 );
buf \U$27878 ( \36389_36689 , \36388_36688 );
and \U$27879 ( \36390_36690 , \36117_36417 , \36122_36422 );
and \U$27880 ( \36391_36691 , \36117_36417 , \36128_36428 );
and \U$27881 ( \36392_36692 , \36122_36422 , \36128_36428 );
or \U$27882 ( \36393_36693 , \36390_36690 , \36391_36691 , \36392_36692 );
buf \U$27883 ( \36394_36694 , \36393_36693 );
and \U$27884 ( \36395_36695 , \36136_36436 , \36296_36596 );
and \U$27885 ( \36396_36696 , \36136_36436 , \36317_36617 );
and \U$27886 ( \36397_36697 , \36296_36596 , \36317_36617 );
or \U$27887 ( \36398_36698 , \36395_36695 , \36396_36696 , \36397_36697 );
buf \U$27888 ( \36399_36699 , \36398_36698 );
xor \U$27889 ( \36400_36700 , \36394_36694 , \36399_36699 );
and \U$27890 ( \36401_36701 , \36141_36441 , \36147_36447 );
and \U$27891 ( \36402_36702 , \36141_36441 , \36154_36454 );
and \U$27892 ( \36403_36703 , \36147_36447 , \36154_36454 );
or \U$27893 ( \36404_36704 , \36401_36701 , \36402_36702 , \36403_36703 );
buf \U$27894 ( \36405_36705 , \36404_36704 );
and \U$27895 ( \36406_36706 , \16405_15940 , \32589_32888_nG9bb1 );
and \U$27896 ( \36407_36707 , \15638_15937 , \32881_33181_nG9bae );
or \U$27897 ( \36408_36708 , \36406_36706 , \36407_36707 );
xor \U$27898 ( \36409_36709 , \15637_15936 , \36408_36708 );
buf \U$27899 ( \36410_36710 , \36409_36709 );
buf \U$27901 ( \36411_36711 , \36410_36710 );
xor \U$27902 ( \36412_36712 , \36405_36705 , \36411_36711 );
and \U$27903 ( \36413_36713 , \14710_14631 , \33313_33613_nG9bab );
and \U$27904 ( \36414_36714 , \14329_14628 , \33741_34041_nG9ba8 );
or \U$27905 ( \36415_36715 , \36413_36713 , \36414_36714 );
xor \U$27906 ( \36416_36716 , \14328_14627 , \36415_36715 );
buf \U$27907 ( \36417_36717 , \36416_36716 );
buf \U$27909 ( \36418_36718 , \36417_36717 );
xor \U$27910 ( \36419_36719 , \36412_36712 , \36418_36718 );
buf \U$27911 ( \36420_36720 , \36419_36719 );
and \U$27912 ( \36421_36721 , \36089_36389 , \36091_36391 );
and \U$27913 ( \36422_36722 , \36089_36389 , \36098_36398 );
and \U$27914 ( \36423_36723 , \36091_36391 , \36098_36398 );
or \U$27915 ( \36424_36724 , \36421_36721 , \36422_36722 , \36423_36723 );
buf \U$27916 ( \36425_36725 , \36424_36724 );
and \U$27917 ( \36426_36726 , \28946_28118 , \19287_19586_nG9be1 );
and \U$27918 ( \36427_36727 , \27816_28115 , \20306_20608_nG9bde );
or \U$27919 ( \36428_36728 , \36426_36726 , \36427_36727 );
xor \U$27920 ( \36429_36729 , \27815_28114 , \36428_36728 );
buf \U$27921 ( \36430_36730 , \36429_36729 );
buf \U$27923 ( \36431_36731 , \36430_36730 );
xor \U$27924 ( \36432_36732 , \36425_36725 , \36431_36731 );
and \U$27925 ( \36433_36733 , \27141_26431 , \20787_21086_nG9bdb );
and \U$27926 ( \36434_36734 , \26129_26428 , \21827_22129_nG9bd8 );
or \U$27927 ( \36435_36735 , \36433_36733 , \36434_36734 );
xor \U$27928 ( \36436_36736 , \26128_26427 , \36435_36735 );
buf \U$27929 ( \36437_36737 , \36436_36736 );
buf \U$27931 ( \36438_36738 , \36437_36737 );
xor \U$27932 ( \36439_36739 , \36432_36732 , \36438_36738 );
buf \U$27933 ( \36440_36740 , \36439_36739 );
and \U$27934 ( \36441_36741 , \18908_18702 , \28877_29179_nG9bbd );
and \U$27935 ( \36442_36742 , \18400_18699 , \30064_30366_nG9bba );
or \U$27936 ( \36443_36743 , \36441_36741 , \36442_36742 );
xor \U$27937 ( \36444_36744 , \18399_18698 , \36443_36743 );
buf \U$27938 ( \36445_36745 , \36444_36744 );
buf \U$27940 ( \36446_36746 , \36445_36745 );
xor \U$27941 ( \36447_36747 , \36440_36740 , \36446_36746 );
and \U$27942 ( \36448_36748 , \17437_17297 , \30638_30940_nG9bb7 );
and \U$27943 ( \36449_36749 , \16995_17294 , \31877_32179_nG9bb4 );
or \U$27944 ( \36450_36750 , \36448_36748 , \36449_36749 );
xor \U$27945 ( \36451_36751 , \16994_17293 , \36450_36750 );
buf \U$27946 ( \36452_36752 , \36451_36751 );
buf \U$27948 ( \36453_36753 , \36452_36752 );
xor \U$27949 ( \36454_36754 , \36447_36747 , \36453_36753 );
buf \U$27950 ( \36455_36755 , \36454_36754 );
xor \U$27951 ( \36456_36756 , \36420_36720 , \36455_36755 );
and \U$27952 ( \36457_36757 , \36302_36602 , \36308_36608 );
and \U$27953 ( \36458_36758 , \36302_36602 , \36315_36615 );
and \U$27954 ( \36459_36759 , \36308_36608 , \36315_36615 );
or \U$27955 ( \36460_36760 , \36457_36757 , \36458_36758 , \36459_36759 );
buf \U$27956 ( \36461_36761 , \36460_36760 );
xor \U$27957 ( \36462_36762 , \36456_36756 , \36461_36761 );
buf \U$27958 ( \36463_36763 , \36462_36762 );
xor \U$27959 ( \36464_36764 , \36400_36700 , \36463_36763 );
buf \U$27960 ( \36465_36765 , \36464_36764 );
xor \U$27961 ( \36466_36766 , \36389_36689 , \36465_36765 );
and \U$27962 ( \36467_36767 , \36327_36627 , \36332_36632 );
and \U$27963 ( \36468_36768 , \36327_36627 , \36367_36667 );
and \U$27964 ( \36469_36769 , \36332_36632 , \36367_36667 );
or \U$27965 ( \36470_36770 , \36467_36767 , \36468_36768 , \36469_36769 );
buf \U$27966 ( \36471_36771 , \36470_36770 );
and \U$27967 ( \36472_36772 , \36354_36654 , \36359_36659 );
and \U$27968 ( \36473_36773 , \36354_36654 , \36365_36665 );
and \U$27969 ( \36474_36774 , \36359_36659 , \36365_36665 );
or \U$27970 ( \36475_36775 , \36472_36772 , \36473_36773 , \36474_36774 );
buf \U$27971 ( \36476_36776 , \36475_36775 );
and \U$27972 ( \36477_36777 , \36339_36639 , \36345_36645 );
and \U$27973 ( \36478_36778 , \36339_36639 , \36352_36652 );
and \U$27974 ( \36479_36779 , \36345_36645 , \36352_36652 );
or \U$27975 ( \36480_36780 , \36477_36777 , \36478_36778 , \36479_36779 );
buf \U$27976 ( \36481_36781 , \36480_36780 );
and \U$27977 ( \36482_36782 , \36041_36341 , \36061_36361 );
and \U$27978 ( \36483_36783 , \36041_36341 , \36068_36368 );
and \U$27979 ( \36484_36784 , \36061_36361 , \36068_36368 );
or \U$27980 ( \36485_36785 , \36482_36782 , \36483_36783 , \36484_36784 );
buf \U$27981 ( \36486_36786 , \36485_36785 );
xor \U$27982 ( \36487_36787 , \36481_36781 , \36486_36786 );
and \U$27983 ( \36488_36788 , \36046_36346 , \36052_36352 );
and \U$27984 ( \36489_36789 , \36046_36346 , \36059_36359 );
and \U$27985 ( \36490_36790 , \36052_36352 , \36059_36359 );
or \U$27986 ( \36491_36791 , \36488_36788 , \36489_36789 , \36490_36790 );
buf \U$27987 ( \36492_36792 , \36491_36791 );
and \U$27988 ( \36493_36793 , \21908_21658 , \25561_25860_nG9bc9 );
and \U$27989 ( \36494_36794 , \21356_21655 , \26585_26887_nG9bc6 );
or \U$27990 ( \36495_36795 , \36493_36793 , \36494_36794 );
xor \U$27991 ( \36496_36796 , \21355_21654 , \36495_36795 );
buf \U$27992 ( \36497_36797 , \36496_36796 );
buf \U$27994 ( \36498_36798 , \36497_36797 );
xor \U$27995 ( \36499_36799 , \36492_36792 , \36498_36798 );
and \U$27996 ( \36500_36800 , \20353_20155 , \27114_27416_nG9bc3 );
and \U$27997 ( \36501_36801 , \19853_20152 , \28300_28602_nG9bc0 );
or \U$27998 ( \36502_36802 , \36500_36800 , \36501_36801 );
xor \U$27999 ( \36503_36803 , \19852_20151 , \36502_36802 );
buf \U$28000 ( \36504_36804 , \36503_36803 );
buf \U$28002 ( \36505_36805 , \36504_36804 );
xor \U$28003 ( \36506_36806 , \36499_36799 , \36505_36805 );
buf \U$28004 ( \36507_36807 , \36506_36806 );
xor \U$28005 ( \36508_36808 , \36487_36787 , \36507_36807 );
buf \U$28006 ( \36509_36809 , \36508_36808 );
xor \U$28007 ( \36510_36810 , \36476_36776 , \36509_36809 );
and \U$28008 ( \36511_36811 , \36070_36370 , \36075_36375 );
and \U$28009 ( \36512_36812 , \36070_36370 , \36115_36415 );
and \U$28010 ( \36513_36813 , \36075_36375 , \36115_36415 );
or \U$28011 ( \36514_36814 , \36511_36811 , \36512_36812 , \36513_36813 );
buf \U$28012 ( \36515_36815 , \36514_36814 );
xor \U$28013 ( \36516_36816 , \36510_36810 , \36515_36815 );
buf \U$28014 ( \36517_36817 , \36516_36816 );
xor \U$28015 ( \36518_36818 , \36471_36771 , \36517_36817 );
and \U$28017 ( \36519_36819 , \32617_32916 , \16013_16315_nG9bf0 );
or \U$28018 ( \36520_36820 , 1'b0 , \36519_36819 );
xor \U$28019 ( \36521_36821 , 1'b0 , \36520_36820 );
buf \U$28020 ( \36522_36822 , \36521_36821 );
buf \U$28022 ( \36523_36823 , \36522_36822 );
and \U$28023 ( \36524_36824 , \31989_31636 , \16378_16680_nG9bed );
and \U$28024 ( \36525_36825 , \31334_31633 , \17363_17665_nG9bea );
or \U$28025 ( \36526_36826 , \36524_36824 , \36525_36825 );
xor \U$28026 ( \36527_36827 , \31333_31632 , \36526_36826 );
buf \U$28027 ( \36528_36828 , \36527_36827 );
buf \U$28029 ( \36529_36829 , \36528_36828 );
xor \U$28030 ( \36530_36830 , \36523_36823 , \36529_36829 );
buf \U$28031 ( \36531_36831 , \36530_36830 );
and \U$28032 ( \36532_36832 , \36081_36381 , \36087_36387 );
buf \U$28033 ( \36533_36833 , \36532_36832 );
xor \U$28034 ( \36534_36834 , \36531_36831 , \36533_36833 );
and \U$28035 ( \36535_36835 , \30670_29853 , \17808_18107_nG9be7 );
and \U$28036 ( \36536_36836 , \29551_29850 , \18789_19091_nG9be4 );
or \U$28037 ( \36537_36837 , \36535_36835 , \36536_36836 );
xor \U$28038 ( \36538_36838 , \29550_29849 , \36537_36837 );
buf \U$28039 ( \36539_36839 , \36538_36838 );
buf \U$28041 ( \36540_36840 , \36539_36839 );
xor \U$28042 ( \36541_36841 , \36534_36834 , \36540_36840 );
buf \U$28043 ( \36542_36842 , \36541_36841 );
and \U$28044 ( \36543_36843 , \25044_24792 , \22330_22629_nG9bd5 );
and \U$28045 ( \36544_36844 , \24490_24789 , \23394_23696_nG9bd2 );
or \U$28046 ( \36545_36845 , \36543_36843 , \36544_36844 );
xor \U$28047 ( \36546_36846 , \24489_24788 , \36545_36845 );
buf \U$28048 ( \36547_36847 , \36546_36846 );
buf \U$28050 ( \36548_36848 , \36547_36847 );
xor \U$28051 ( \36549_36849 , \36542_36842 , \36548_36848 );
and \U$28052 ( \36550_36850 , \23495_23201 , \23927_24226_nG9bcf );
and \U$28053 ( \36551_36851 , \22899_23198 , \24996_25298_nG9bcc );
or \U$28054 ( \36552_36852 , \36550_36850 , \36551_36851 );
xor \U$28055 ( \36553_36853 , \22898_23197 , \36552_36852 );
buf \U$28056 ( \36554_36854 , \36553_36853 );
buf \U$28058 ( \36555_36855 , \36554_36854 );
xor \U$28059 ( \36556_36856 , \36549_36849 , \36555_36855 );
buf \U$28060 ( \36557_36857 , \36556_36856 );
and \U$28061 ( \36558_36858 , \12183_12157 , \34794_35094_nG9b9f );
and \U$28062 ( \36559_36859 , \11855_12154 , \35270_35570_nG9b9c );
or \U$28063 ( \36560_36860 , \36558_36858 , \36559_36859 );
xor \U$28064 ( \36561_36861 , \11854_12153 , \36560_36860 );
buf \U$28065 ( \36562_36862 , \36561_36861 );
buf \U$28067 ( \36563_36863 , \36562_36862 );
xor \U$28068 ( \36564_36864 , \36557_36857 , \36563_36863 );
and \U$28069 ( \36565_36865 , \10411_10707 , \36289_36589_nG9b93 );
and \U$28070 ( \36566_36866 , \36248_36548 , \36252_36552 );
and \U$28071 ( \36567_36867 , \36252_36552 , \36277_36577 );
and \U$28072 ( \36568_36868 , \36248_36548 , \36277_36577 );
or \U$28073 ( \36569_36869 , \36566_36866 , \36567_36867 , \36568_36868 );
and \U$28074 ( \36570_36870 , \36218_36518 , \36229_36529 );
and \U$28075 ( \36571_36871 , \36229_36529 , \36241_36541 );
and \U$28076 ( \36572_36872 , \36218_36518 , \36241_36541 );
or \U$28077 ( \36573_36873 , \36570_36870 , \36571_36871 , \36572_36872 );
and \U$28078 ( \36574_36874 , \36176_36476 , \36180_36480 );
and \U$28079 ( \36575_36875 , \36180_36480 , \36185_36485 );
and \U$28080 ( \36576_36876 , \36176_36476 , \36185_36485 );
or \U$28081 ( \36577_36877 , \36574_36874 , \36575_36875 , \36576_36876 );
and \U$28082 ( \36578_36878 , \32495_32794 , \16333_16635 );
not \U$28083 ( \36579_36879 , \36578_36878 );
xnor \U$28084 ( \36580_36880 , \36579_36879 , \16323_16625 );
and \U$28085 ( \36581_36881 , \28782_29084 , \19235_19534 );
and \U$28086 ( \36582_36882 , \29966_30268 , \18743_19045 );
nor \U$28087 ( \36583_36883 , \36581_36881 , \36582_36882 );
xnor \U$28088 ( \36584_36884 , \36583_36883 , \19241_19540 );
xor \U$28089 ( \36585_36885 , \36580_36880 , \36584_36884 );
and \U$28090 ( \36586_36886 , \15965_16267 , \32503_32802 );
xor \U$28091 ( \36587_36887 , \36585_36885 , \36586_36886 );
xor \U$28092 ( \36588_36888 , \36577_36877 , \36587_36887 );
and \U$28093 ( \36589_36889 , \27011_27313 , \20706_21005 );
and \U$28094 ( \36590_36890 , \28232_28534 , \20255_20557 );
nor \U$28095 ( \36591_36891 , \36589_36889 , \36590_36890 );
xnor \U$28096 ( \36592_36892 , \36591_36891 , \20712_21011 );
and \U$28097 ( \36593_36893 , \20734_21033 , \27095_27397 );
and \U$28098 ( \36594_36894 , \21788_22090 , \26505_26807 );
nor \U$28099 ( \36595_36895 , \36593_36893 , \36594_36894 );
xnor \U$28100 ( \36596_36896 , \36595_36895 , \26993_27295 );
xor \U$28101 ( \36597_36897 , \36592_36892 , \36596_36896 );
and \U$28102 ( \36598_36898 , \19259_19558 , \28768_29070 );
and \U$28103 ( \36599_36899 , \20242_20544 , \28224_28526 );
nor \U$28104 ( \36600_36900 , \36598_36898 , \36599_36899 );
xnor \U$28105 ( \36601_36901 , \36600_36900 , \28774_29076 );
xor \U$28106 ( \36602_36902 , \36597_36897 , \36601_36901 );
xor \U$28107 ( \36603_36903 , \36588_36888 , \36602_36902 );
xor \U$28108 ( \36604_36904 , \36573_36873 , \36603_36903 );
and \U$28109 ( \36605_36905 , \36266_36566 , \36270_36570 );
and \U$28110 ( \36606_36906 , \36270_36570 , \36275_36575 );
and \U$28111 ( \36607_36907 , \36266_36566 , \36275_36575 );
or \U$28112 ( \36608_36908 , \36605_36905 , \36606_36906 , \36607_36907 );
and \U$28113 ( \36609_36909 , \25516_25815 , \22243_22542 );
and \U$28114 ( \36610_36910 , \26527_26829 , \21801_22103 );
nor \U$28115 ( \36611_36911 , \36609_36909 , \36610_36910 );
xnor \U$28116 ( \36612_36912 , \36611_36911 , \22249_22548 );
and \U$28117 ( \36613_36913 , \17736_18035 , \30521_30823 );
and \U$28118 ( \36614_36914 , \18730_19032 , \29944_30246 );
nor \U$28119 ( \36615_36915 , \36613_36913 , \36614_36914 );
xnor \U$28120 ( \36616_36916 , \36615_36915 , \30511_30813 );
xor \U$28121 ( \36617_36917 , \36612_36912 , \36616_36916 );
and \U$28122 ( \36618_36918 , \16353_16655 , \32555_32854 );
and \U$28123 ( \36619_36919 , \17325_17627 , \31765_32067 );
nor \U$28124 ( \36620_36920 , \36618_36918 , \36619_36919 );
xnor \U$28125 ( \36621_36921 , \36620_36920 , \32506_32805 );
xor \U$28126 ( \36622_36922 , \36617_36917 , \36621_36921 );
xor \U$28127 ( \36623_36923 , \36608_36908 , \36622_36922 );
and \U$28128 ( \36624_36924 , \30500_30802 , \17791_18090 );
and \U$28129 ( \36625_36925 , \31752_32054 , \17353_17655 );
nor \U$28130 ( \36626_36926 , \36624_36924 , \36625_36925 );
xnor \U$28131 ( \36627_36927 , \36626_36926 , \17747_18046 );
not \U$28132 ( \36628_36928 , \36627_36927 );
and \U$28133 ( \36629_36929 , \23900_24199 , \23839_24138 );
and \U$28134 ( \36630_36930 , \24970_25272 , \23328_23630 );
nor \U$28135 ( \36631_36931 , \36629_36929 , \36630_36930 );
xnor \U$28136 ( \36632_36932 , \36631_36931 , \23845_24144 );
xor \U$28137 ( \36633_36933 , \36628_36928 , \36632_36932 );
and \U$28138 ( \36634_36934 , \22257_22556 , \25527_25826 );
and \U$28139 ( \36635_36935 , \23315_23617 , \24962_25264 );
nor \U$28140 ( \36636_36936 , \36634_36934 , \36635_36935 );
xnor \U$28141 ( \36637_36937 , \36636_36936 , \25474_25773 );
xor \U$28142 ( \36638_36938 , \36633_36933 , \36637_36937 );
xor \U$28143 ( \36639_36939 , \36623_36923 , \36638_36938 );
xor \U$28144 ( \36640_36940 , \36604_36904 , \36639_36939 );
xor \U$28145 ( \36641_36941 , \36569_36869 , \36640_36940 );
and \U$28146 ( \36642_36942 , \36257_36557 , \36261_36561 );
and \U$28147 ( \36643_36943 , \36261_36561 , \36276_36576 );
and \U$28148 ( \36644_36944 , \36257_36557 , \36276_36576 );
or \U$28149 ( \36645_36945 , \36642_36942 , \36643_36943 , \36644_36944 );
and \U$28150 ( \36646_36946 , \36172_36472 , \36213_36513 );
and \U$28151 ( \36647_36947 , \36213_36513 , \36242_36542 );
and \U$28152 ( \36648_36948 , \36172_36472 , \36242_36542 );
or \U$28153 ( \36649_36949 , \36646_36946 , \36647_36947 , \36648_36948 );
xor \U$28154 ( \36650_36950 , \36645_36945 , \36649_36949 );
and \U$28155 ( \36651_36951 , \36234_36534 , \36235_36535 );
and \U$28156 ( \36652_36952 , \36235_36535 , \36240_36540 );
and \U$28157 ( \36653_36953 , \36234_36534 , \36240_36540 );
or \U$28158 ( \36654_36954 , \36651_36951 , \36652_36952 , \36653_36953 );
and \U$28159 ( \36655_36955 , \36186_36486 , \36197_36497 );
and \U$28160 ( \36656_36956 , \36197_36497 , \36212_36512 );
and \U$28161 ( \36657_36957 , \36186_36486 , \36212_36512 );
or \U$28162 ( \36658_36958 , \36655_36955 , \36656_36956 , \36657_36957 );
xor \U$28163 ( \36659_36959 , \36654_36954 , \36658_36958 );
and \U$28164 ( \36660_36960 , \36222_36522 , \36226_36526 );
and \U$28165 ( \36661_36961 , \36226_36526 , \36228_36528 );
and \U$28166 ( \36662_36962 , \36222_36522 , \36228_36528 );
or \U$28167 ( \36663_36963 , \36660_36960 , \36661_36961 , \36662_36962 );
and \U$28168 ( \36664_36964 , \36187_36487 , \36191_36491 );
and \U$28169 ( \36665_36965 , \36191_36491 , \36196_36496 );
and \U$28170 ( \36666_36966 , \36187_36487 , \36196_36496 );
or \U$28171 ( \36667_36967 , \36664_36964 , \36665_36965 , \36666_36966 );
xor \U$28172 ( \36668_36968 , \36663_36963 , \36667_36967 );
and \U$28173 ( \36669_36969 , \36202_36502 , \36206_36506 );
and \U$28174 ( \36670_36970 , \36206_36506 , \36211_36511 );
and \U$28175 ( \36671_36971 , \36202_36502 , \36211_36511 );
or \U$28176 ( \36672_36972 , \36669_36969 , \36670_36970 , \36671_36971 );
xor \U$28177 ( \36673_36973 , \36668_36968 , \36672_36972 );
xor \U$28178 ( \36674_36974 , \36659_36959 , \36673_36973 );
xor \U$28179 ( \36675_36975 , \36650_36950 , \36674_36974 );
xor \U$28180 ( \36676_36976 , \36641_36941 , \36675_36975 );
and \U$28181 ( \36677_36977 , \36168_36468 , \36243_36543 );
and \U$28182 ( \36678_36978 , \36243_36543 , \36278_36578 );
and \U$28183 ( \36679_36979 , \36168_36468 , \36278_36578 );
or \U$28184 ( \36680_36980 , \36677_36977 , \36678_36978 , \36679_36979 );
xor \U$28185 ( \36681_36981 , \36676_36976 , \36680_36980 );
and \U$28186 ( \36682_36982 , \36279_36579 , \36283_36583 );
and \U$28187 ( \36683_36983 , \36284_36584 , \36287_36587 );
or \U$28188 ( \36684_36984 , \36682_36982 , \36683_36983 );
xor \U$28189 ( \36685_36985 , \36681_36981 , \36684_36984 );
buf g9b90_GF_PartitionCandidate( \36686_36986_nG9b90 , \36685_36985 );
and \U$28190 ( \36687_36987 , \10402_10704 , \36686_36986_nG9b90 );
or \U$28191 ( \36688_36988 , \36565_36865 , \36687_36987 );
xor \U$28192 ( \36689_36989 , \10399_10703 , \36688_36988 );
buf \U$28193 ( \36690_36990 , \36689_36989 );
buf \U$28195 ( \36691_36991 , \36690_36990 );
xor \U$28196 ( \36692_36992 , \36564_36864 , \36691_36991 );
buf \U$28197 ( \36693_36993 , \36692_36992 );
and \U$28198 ( \36694_36994 , \36100_36400 , \36106_36406 );
and \U$28199 ( \36695_36995 , \36100_36400 , \36113_36413 );
and \U$28200 ( \36696_36996 , \36106_36406 , \36113_36413 );
or \U$28201 ( \36697_36997 , \36694_36994 , \36695_36995 , \36696_36996 );
buf \U$28202 ( \36698_36998 , \36697_36997 );
and \U$28203 ( \36699_36999 , \13431_13370 , \33994_34294_nG9ba5 );
and \U$28204 ( \36700_37000 , \13068_13367 , \34343_34643_nG9ba2 );
or \U$28205 ( \36701_37001 , \36699_36999 , \36700_37000 );
xor \U$28206 ( \36702_37002 , \13067_13366 , \36701_37001 );
buf \U$28207 ( \36703_37003 , \36702_37002 );
buf \U$28209 ( \36704_37004 , \36703_37003 );
xor \U$28210 ( \36705_37005 , \36698_36998 , \36704_37004 );
and \U$28211 ( \36706_37006 , \10996_10421 , \35501_35801_nG9b99 );
and \U$28212 ( \36707_37007 , \10119_10418 , \35872_36172_nG9b96 );
or \U$28213 ( \36708_37008 , \36706_37006 , \36707_37007 );
xor \U$28214 ( \36709_37009 , \10118_10417 , \36708_37008 );
buf \U$28215 ( \36710_37010 , \36709_37009 );
buf \U$28217 ( \36711_37011 , \36710_37010 );
xor \U$28218 ( \36712_37012 , \36705_37005 , \36711_37011 );
buf \U$28219 ( \36713_37013 , \36712_37012 );
xor \U$28220 ( \36714_37014 , \36693_36993 , \36713_37013 );
and \U$28221 ( \36715_37015 , \36156_36456 , \36162_36462 );
and \U$28222 ( \36716_37016 , \36156_36456 , \36294_36594 );
and \U$28223 ( \36717_37017 , \36162_36462 , \36294_36594 );
or \U$28224 ( \36718_37018 , \36715_37015 , \36716_37016 , \36717_37017 );
buf \U$28225 ( \36719_37019 , \36718_37018 );
xor \U$28226 ( \36720_37020 , \36714_37014 , \36719_37019 );
buf \U$28227 ( \36721_37021 , \36720_37020 );
xor \U$28228 ( \36722_37022 , \36518_36818 , \36721_37021 );
buf \U$28229 ( \36723_37023 , \36722_37022 );
xor \U$28230 ( \36724_37024 , \36466_36766 , \36723_37023 );
and \U$28231 ( \36725_37025 , \36384_36684 , \36724_37024 );
and \U$28233 ( \36726_37026 , \36378_36678 , \36383_36683 );
or \U$28235 ( \36727_37027 , 1'b0 , \36726_37026 , 1'b0 );
xor \U$28236 ( \36728_37028 , \36725_37025 , \36727_37027 );
and \U$28238 ( \36729_37029 , \36371_36671 , \36377_36677 );
and \U$28239 ( \36730_37030 , \36373_36673 , \36377_36677 );
or \U$28240 ( \36731_37031 , 1'b0 , \36729_37029 , \36730_37030 );
xor \U$28241 ( \36732_37032 , \36728_37028 , \36731_37031 );
xor \U$28248 ( \36733_37033 , \36732_37032 , 1'b0 );
and \U$28249 ( \36734_37034 , \36389_36689 , \36465_36765 );
and \U$28250 ( \36735_37035 , \36389_36689 , \36723_37023 );
and \U$28251 ( \36736_37036 , \36465_36765 , \36723_37023 );
or \U$28252 ( \36737_37037 , \36734_37034 , \36735_37035 , \36736_37036 );
xor \U$28253 ( \36738_37038 , \36733_37033 , \36737_37037 );
and \U$28254 ( \36739_37039 , \36471_36771 , \36517_36817 );
and \U$28255 ( \36740_37040 , \36471_36771 , \36721_37021 );
and \U$28256 ( \36741_37041 , \36517_36817 , \36721_37021 );
or \U$28257 ( \36742_37042 , \36739_37039 , \36740_37040 , \36741_37041 );
buf \U$28258 ( \36743_37043 , \36742_37042 );
and \U$28259 ( \36744_37044 , \36481_36781 , \36486_36786 );
and \U$28260 ( \36745_37045 , \36481_36781 , \36507_36807 );
and \U$28261 ( \36746_37046 , \36486_36786 , \36507_36807 );
or \U$28262 ( \36747_37047 , \36744_37044 , \36745_37045 , \36746_37046 );
buf \U$28263 ( \36748_37048 , \36747_37047 );
and \U$28264 ( \36749_37049 , \36425_36725 , \36431_36731 );
and \U$28265 ( \36750_37050 , \36425_36725 , \36438_36738 );
and \U$28266 ( \36751_37051 , \36431_36731 , \36438_36738 );
or \U$28267 ( \36752_37052 , \36749_37049 , \36750_37050 , \36751_37051 );
buf \U$28268 ( \36753_37053 , \36752_37052 );
and \U$28269 ( \36754_37054 , \36523_36823 , \36529_36829 );
buf \U$28270 ( \36755_37055 , \36754_37054 );
and \U$28271 ( \36756_37056 , \30670_29853 , \18789_19091_nG9be4 );
and \U$28272 ( \36757_37057 , \29551_29850 , \19287_19586_nG9be1 );
or \U$28273 ( \36758_37058 , \36756_37056 , \36757_37057 );
xor \U$28274 ( \36759_37059 , \29550_29849 , \36758_37058 );
buf \U$28275 ( \36760_37060 , \36759_37059 );
buf \U$28277 ( \36761_37061 , \36760_37060 );
xor \U$28278 ( \36762_37062 , \36755_37055 , \36761_37061 );
and \U$28279 ( \36763_37063 , \28946_28118 , \20306_20608_nG9bde );
and \U$28280 ( \36764_37064 , \27816_28115 , \20787_21086_nG9bdb );
or \U$28281 ( \36765_37065 , \36763_37063 , \36764_37064 );
xor \U$28282 ( \36766_37066 , \27815_28114 , \36765_37065 );
buf \U$28283 ( \36767_37067 , \36766_37066 );
buf \U$28285 ( \36768_37068 , \36767_37067 );
xor \U$28286 ( \36769_37069 , \36762_37062 , \36768_37068 );
buf \U$28287 ( \36770_37070 , \36769_37069 );
xor \U$28288 ( \36771_37071 , \36753_37053 , \36770_37070 );
and \U$28289 ( \36772_37072 , \18908_18702 , \30064_30366_nG9bba );
and \U$28290 ( \36773_37073 , \18400_18699 , \30638_30940_nG9bb7 );
or \U$28291 ( \36774_37074 , \36772_37072 , \36773_37073 );
xor \U$28292 ( \36775_37075 , \18399_18698 , \36774_37074 );
buf \U$28293 ( \36776_37076 , \36775_37075 );
buf \U$28295 ( \36777_37077 , \36776_37076 );
xor \U$28296 ( \36778_37078 , \36771_37071 , \36777_37077 );
buf \U$28297 ( \36779_37079 , \36778_37078 );
and \U$28298 ( \36780_37080 , \25044_24792 , \23394_23696_nG9bd2 );
and \U$28299 ( \36781_37081 , \24490_24789 , \23927_24226_nG9bcf );
or \U$28300 ( \36782_37082 , \36780_37080 , \36781_37081 );
xor \U$28301 ( \36783_37083 , \24489_24788 , \36782_37082 );
buf \U$28302 ( \36784_37084 , \36783_37083 );
buf \U$28304 ( \36785_37085 , \36784_37084 );
and \U$28305 ( \36786_37086 , \23495_23201 , \24996_25298_nG9bcc );
and \U$28306 ( \36787_37087 , \22899_23198 , \25561_25860_nG9bc9 );
or \U$28307 ( \36788_37088 , \36786_37086 , \36787_37087 );
xor \U$28308 ( \36789_37089 , \22898_23197 , \36788_37088 );
buf \U$28309 ( \36790_37090 , \36789_37089 );
buf \U$28311 ( \36791_37091 , \36790_37090 );
xor \U$28312 ( \36792_37092 , \36785_37085 , \36791_37091 );
and \U$28313 ( \36793_37093 , \21908_21658 , \26585_26887_nG9bc6 );
and \U$28314 ( \36794_37094 , \21356_21655 , \27114_27416_nG9bc3 );
or \U$28315 ( \36795_37095 , \36793_37093 , \36794_37094 );
xor \U$28316 ( \36796_37096 , \21355_21654 , \36795_37095 );
buf \U$28317 ( \36797_37097 , \36796_37096 );
buf \U$28319 ( \36798_37098 , \36797_37097 );
xor \U$28320 ( \36799_37099 , \36792_37092 , \36798_37098 );
buf \U$28321 ( \36800_37100 , \36799_37099 );
xor \U$28322 ( \36801_37101 , \36779_37079 , \36800_37100 );
and \U$28323 ( \36802_37102 , \36405_36705 , \36411_36711 );
and \U$28324 ( \36803_37103 , \36405_36705 , \36418_36718 );
and \U$28325 ( \36804_37104 , \36411_36711 , \36418_36718 );
or \U$28326 ( \36805_37105 , \36802_37102 , \36803_37103 , \36804_37104 );
buf \U$28327 ( \36806_37106 , \36805_37105 );
xor \U$28328 ( \36807_37107 , \36801_37101 , \36806_37106 );
buf \U$28329 ( \36808_37108 , \36807_37107 );
xor \U$28330 ( \36809_37109 , \36748_37048 , \36808_37108 );
and \U$28331 ( \36810_37110 , \36420_36720 , \36455_36755 );
and \U$28332 ( \36811_37111 , \36420_36720 , \36461_36761 );
and \U$28333 ( \36812_37112 , \36455_36755 , \36461_36761 );
or \U$28334 ( \36813_37113 , \36810_37110 , \36811_37111 , \36812_37112 );
buf \U$28335 ( \36814_37114 , \36813_37113 );
xor \U$28336 ( \36815_37115 , \36809_37109 , \36814_37114 );
buf \U$28337 ( \36816_37116 , \36815_37115 );
and \U$28338 ( \36817_37117 , \36476_36776 , \36509_36809 );
and \U$28339 ( \36818_37118 , \36476_36776 , \36515_36815 );
and \U$28340 ( \36819_37119 , \36509_36809 , \36515_36815 );
or \U$28341 ( \36820_37120 , \36817_37117 , \36818_37118 , \36819_37119 );
buf \U$28342 ( \36821_37121 , \36820_37120 );
xor \U$28343 ( \36822_37122 , \36816_37116 , \36821_37121 );
and \U$28344 ( \36823_37123 , \36440_36740 , \36446_36746 );
and \U$28345 ( \36824_37124 , \36440_36740 , \36453_36753 );
and \U$28346 ( \36825_37125 , \36446_36746 , \36453_36753 );
or \U$28347 ( \36826_37126 , \36823_37123 , \36824_37124 , \36825_37125 );
buf \U$28348 ( \36827_37127 , \36826_37126 );
and \U$28349 ( \36828_37128 , \10996_10421 , \35872_36172_nG9b96 );
and \U$28350 ( \36829_37129 , \10119_10418 , \36289_36589_nG9b93 );
or \U$28351 ( \36830_37130 , \36828_37128 , \36829_37129 );
xor \U$28352 ( \36831_37131 , \10118_10417 , \36830_37130 );
buf \U$28353 ( \36832_37132 , \36831_37131 );
buf \U$28355 ( \36833_37133 , \36832_37132 );
xor \U$28356 ( \36834_37134 , \36827_37127 , \36833_37133 );
and \U$28357 ( \36835_37135 , \10411_10707 , \36686_36986_nG9b90 );
and \U$28358 ( \36836_37136 , \36645_36945 , \36649_36949 );
and \U$28359 ( \36837_37137 , \36649_36949 , \36674_36974 );
and \U$28360 ( \36838_37138 , \36645_36945 , \36674_36974 );
or \U$28361 ( \36839_37139 , \36836_37136 , \36837_37137 , \36838_37138 );
and \U$28362 ( \36840_37140 , \36608_36908 , \36622_36922 );
and \U$28363 ( \36841_37141 , \36622_36922 , \36638_36938 );
and \U$28364 ( \36842_37142 , \36608_36908 , \36638_36938 );
or \U$28365 ( \36843_37143 , \36840_37140 , \36841_37141 , \36842_37142 );
and \U$28366 ( \36844_37144 , \36628_36928 , \36632_36932 );
and \U$28367 ( \36845_37145 , \36632_36932 , \36637_36937 );
and \U$28368 ( \36846_37146 , \36628_36928 , \36637_36937 );
or \U$28369 ( \36847_37147 , \36844_37144 , \36845_37145 , \36846_37146 );
not \U$28370 ( \36848_37148 , \16323_16625 );
and \U$28371 ( \36849_37149 , \31752_32054 , \17791_18090 );
and \U$28372 ( \36850_37150 , \32495_32794 , \17353_17655 );
nor \U$28373 ( \36851_37151 , \36849_37149 , \36850_37150 );
xnor \U$28374 ( \36852_37152 , \36851_37151 , \17747_18046 );
xor \U$28375 ( \36853_37153 , \36848_37148 , \36852_37152 );
and \U$28376 ( \36854_37154 , \28232_28534 , \20706_21005 );
and \U$28377 ( \36855_37155 , \28782_29084 , \20255_20557 );
nor \U$28378 ( \36856_37156 , \36854_37154 , \36855_37155 );
xnor \U$28379 ( \36857_37157 , \36856_37156 , \20712_21011 );
xor \U$28380 ( \36858_37158 , \36853_37153 , \36857_37157 );
xor \U$28381 ( \36859_37159 , \36847_37147 , \36858_37158 );
and \U$28382 ( \36860_37160 , \26527_26829 , \22243_22542 );
and \U$28383 ( \36861_37161 , \27011_27313 , \21801_22103 );
nor \U$28384 ( \36862_37162 , \36860_37160 , \36861_37161 );
xnor \U$28385 ( \36863_37163 , \36862_37162 , \22249_22548 );
and \U$28386 ( \36864_37164 , \21788_22090 , \27095_27397 );
and \U$28387 ( \36865_37165 , \22257_22556 , \26505_26807 );
nor \U$28388 ( \36866_37166 , \36864_37164 , \36865_37165 );
xnor \U$28389 ( \36867_37167 , \36866_37166 , \26993_27295 );
xor \U$28390 ( \36868_37168 , \36863_37163 , \36867_37167 );
and \U$28391 ( \36869_37169 , \20242_20544 , \28768_29070 );
and \U$28392 ( \36870_37170 , \20734_21033 , \28224_28526 );
nor \U$28393 ( \36871_37171 , \36869_37169 , \36870_37170 );
xnor \U$28394 ( \36872_37172 , \36871_37171 , \28774_29076 );
xor \U$28395 ( \36873_37173 , \36868_37168 , \36872_37172 );
xor \U$28396 ( \36874_37174 , \36859_37159 , \36873_37173 );
xor \U$28397 ( \36875_37175 , \36843_37143 , \36874_37174 );
and \U$28398 ( \36876_37176 , \36612_36912 , \36616_36916 );
and \U$28399 ( \36877_37177 , \36616_36916 , \36621_36921 );
and \U$28400 ( \36878_37178 , \36612_36912 , \36621_36921 );
or \U$28401 ( \36879_37179 , \36876_37176 , \36877_37177 , \36878_37178 );
and \U$28402 ( \36880_37180 , \29966_30268 , \19235_19534 );
and \U$28403 ( \36881_37181 , \30500_30802 , \18743_19045 );
nor \U$28404 ( \36882_37182 , \36880_37180 , \36881_37181 );
xnor \U$28405 ( \36883_37183 , \36882_37182 , \19241_19540 );
and \U$28406 ( \36884_37184 , \18730_19032 , \30521_30823 );
and \U$28407 ( \36885_37185 , \19259_19558 , \29944_30246 );
nor \U$28408 ( \36886_37186 , \36884_37184 , \36885_37185 );
xnor \U$28409 ( \36887_37187 , \36886_37186 , \30511_30813 );
xor \U$28410 ( \36888_37188 , \36883_37183 , \36887_37187 );
and \U$28411 ( \36889_37189 , \17325_17627 , \32555_32854 );
and \U$28412 ( \36890_37190 , \17736_18035 , \31765_32067 );
nor \U$28413 ( \36891_37191 , \36889_37189 , \36890_37190 );
xnor \U$28414 ( \36892_37192 , \36891_37191 , \32506_32805 );
xor \U$28415 ( \36893_37193 , \36888_37188 , \36892_37192 );
xor \U$28416 ( \36894_37194 , \36879_37179 , \36893_37193 );
and \U$28417 ( \36895_37195 , \24970_25272 , \23839_24138 );
and \U$28418 ( \36896_37196 , \25516_25815 , \23328_23630 );
nor \U$28419 ( \36897_37197 , \36895_37195 , \36896_37196 );
xnor \U$28420 ( \36898_37198 , \36897_37197 , \23845_24144 );
and \U$28421 ( \36899_37199 , \23315_23617 , \25527_25826 );
and \U$28422 ( \36900_37200 , \23900_24199 , \24962_25264 );
nor \U$28423 ( \36901_37201 , \36899_37199 , \36900_37200 );
xnor \U$28424 ( \36902_37202 , \36901_37201 , \25474_25773 );
xor \U$28425 ( \36903_37203 , \36898_37198 , \36902_37202 );
and \U$28426 ( \36904_37204 , \16353_16655 , \32503_32802 );
xor \U$28427 ( \36905_37205 , \36903_37203 , \36904_37204 );
xor \U$28428 ( \36906_37206 , \36894_37194 , \36905_37205 );
xor \U$28429 ( \36907_37207 , \36875_37175 , \36906_37206 );
xor \U$28430 ( \36908_37208 , \36839_37139 , \36907_37207 );
and \U$28431 ( \36909_37209 , \36654_36954 , \36658_36958 );
and \U$28432 ( \36910_37210 , \36658_36958 , \36673_36973 );
and \U$28433 ( \36911_37211 , \36654_36954 , \36673_36973 );
or \U$28434 ( \36912_37212 , \36909_37209 , \36910_37210 , \36911_37211 );
and \U$28435 ( \36913_37213 , \36573_36873 , \36603_36903 );
and \U$28436 ( \36914_37214 , \36603_36903 , \36639_36939 );
and \U$28437 ( \36915_37215 , \36573_36873 , \36639_36939 );
or \U$28438 ( \36916_37216 , \36913_37213 , \36914_37214 , \36915_37215 );
xor \U$28439 ( \36917_37217 , \36912_37212 , \36916_37216 );
and \U$28440 ( \36918_37218 , \36663_36963 , \36667_36967 );
and \U$28441 ( \36919_37219 , \36667_36967 , \36672_36972 );
and \U$28442 ( \36920_37220 , \36663_36963 , \36672_36972 );
or \U$28443 ( \36921_37221 , \36918_37218 , \36919_37219 , \36920_37220 );
and \U$28444 ( \36922_37222 , \36577_36877 , \36587_36887 );
and \U$28445 ( \36923_37223 , \36587_36887 , \36602_36902 );
and \U$28446 ( \36924_37224 , \36577_36877 , \36602_36902 );
or \U$28447 ( \36925_37225 , \36922_37222 , \36923_37223 , \36924_37224 );
xor \U$28448 ( \36926_37226 , \36921_37221 , \36925_37225 );
and \U$28449 ( \36927_37227 , \36580_36880 , \36584_36884 );
and \U$28450 ( \36928_37228 , \36584_36884 , \36586_36886 );
and \U$28451 ( \36929_37229 , \36580_36880 , \36586_36886 );
or \U$28452 ( \36930_37230 , \36927_37227 , \36928_37228 , \36929_37229 );
and \U$28453 ( \36931_37231 , \36592_36892 , \36596_36896 );
and \U$28454 ( \36932_37232 , \36596_36896 , \36601_36901 );
and \U$28455 ( \36933_37233 , \36592_36892 , \36601_36901 );
or \U$28456 ( \36934_37234 , \36931_37231 , \36932_37232 , \36933_37233 );
xor \U$28457 ( \36935_37235 , \36930_37230 , \36934_37234 );
buf \U$28458 ( \36936_37236 , \36627_36927 );
xor \U$28459 ( \36937_37237 , \36935_37235 , \36936_37236 );
xor \U$28460 ( \36938_37238 , \36926_37226 , \36937_37237 );
xor \U$28461 ( \36939_37239 , \36917_37217 , \36938_37238 );
xor \U$28462 ( \36940_37240 , \36908_37208 , \36939_37239 );
and \U$28463 ( \36941_37241 , \36569_36869 , \36640_36940 );
and \U$28464 ( \36942_37242 , \36640_36940 , \36675_36975 );
and \U$28465 ( \36943_37243 , \36569_36869 , \36675_36975 );
or \U$28466 ( \36944_37244 , \36941_37241 , \36942_37242 , \36943_37243 );
xor \U$28467 ( \36945_37245 , \36940_37240 , \36944_37244 );
and \U$28468 ( \36946_37246 , \36676_36976 , \36680_36980 );
and \U$28469 ( \36947_37247 , \36681_36981 , \36684_36984 );
or \U$28470 ( \36948_37248 , \36946_37246 , \36947_37247 );
xor \U$28471 ( \36949_37249 , \36945_37245 , \36948_37248 );
buf g9b8d_GF_PartitionCandidate( \36950_37250_nG9b8d , \36949_37249 );
and \U$28472 ( \36951_37251 , \10402_10704 , \36950_37250_nG9b8d );
or \U$28473 ( \36952_37252 , \36835_37135 , \36951_37251 );
xor \U$28474 ( \36953_37253 , \10399_10703 , \36952_37252 );
buf \U$28475 ( \36954_37254 , \36953_37253 );
buf \U$28477 ( \36955_37255 , \36954_37254 );
xor \U$28478 ( \36956_37256 , \36834_37134 , \36955_37255 );
buf \U$28479 ( \36957_37257 , \36956_37256 );
and \U$28480 ( \36958_37258 , \36557_36857 , \36563_36863 );
and \U$28481 ( \36959_37259 , \36557_36857 , \36691_36991 );
and \U$28482 ( \36960_37260 , \36563_36863 , \36691_36991 );
or \U$28483 ( \36961_37261 , \36958_37258 , \36959_37259 , \36960_37260 );
buf \U$28484 ( \36962_37262 , \36961_37261 );
xor \U$28485 ( \36963_37263 , \36957_37257 , \36962_37262 );
and \U$28486 ( \36964_37264 , \36492_36792 , \36498_36798 );
and \U$28487 ( \36965_37265 , \36492_36792 , \36505_36805 );
and \U$28488 ( \36966_37266 , \36498_36798 , \36505_36805 );
or \U$28489 ( \36967_37267 , \36964_37264 , \36965_37265 , \36966_37266 );
buf \U$28490 ( \36968_37268 , \36967_37267 );
and \U$28491 ( \36969_37269 , \14710_14631 , \33741_34041_nG9ba8 );
and \U$28492 ( \36970_37270 , \14329_14628 , \33994_34294_nG9ba5 );
or \U$28493 ( \36971_37271 , \36969_37269 , \36970_37270 );
xor \U$28494 ( \36972_37272 , \14328_14627 , \36971_37271 );
buf \U$28495 ( \36973_37273 , \36972_37272 );
buf \U$28497 ( \36974_37274 , \36973_37273 );
xor \U$28498 ( \36975_37275 , \36968_37268 , \36974_37274 );
and \U$28499 ( \36976_37276 , \12183_12157 , \35270_35570_nG9b9c );
and \U$28500 ( \36977_37277 , \11855_12154 , \35501_35801_nG9b99 );
or \U$28501 ( \36978_37278 , \36976_37276 , \36977_37277 );
xor \U$28502 ( \36979_37279 , \11854_12153 , \36978_37278 );
buf \U$28503 ( \36980_37280 , \36979_37279 );
buf \U$28505 ( \36981_37281 , \36980_37280 );
xor \U$28506 ( \36982_37282 , \36975_37275 , \36981_37281 );
buf \U$28507 ( \36983_37283 , \36982_37282 );
xor \U$28508 ( \36984_37284 , \36963_37263 , \36983_37283 );
buf \U$28509 ( \36985_37285 , \36984_37284 );
and \U$28510 ( \36986_37286 , \36698_36998 , \36704_37004 );
and \U$28511 ( \36987_37287 , \36698_36998 , \36711_37011 );
and \U$28512 ( \36988_37288 , \36704_37004 , \36711_37011 );
or \U$28513 ( \36989_37289 , \36986_37286 , \36987_37287 , \36988_37288 );
buf \U$28514 ( \36990_37290 , \36989_37289 );
and \U$28515 ( \36991_37291 , \36531_36831 , \36533_36833 );
and \U$28516 ( \36992_37292 , \36531_36831 , \36540_36840 );
and \U$28517 ( \36993_37293 , \36533_36833 , \36540_36840 );
or \U$28518 ( \36994_37294 , \36991_37291 , \36992_37292 , \36993_37293 );
buf \U$28519 ( \36995_37295 , \36994_37294 );
and \U$28521 ( \36996_37296 , \32617_32916 , \16378_16680_nG9bed );
or \U$28522 ( \36997_37297 , 1'b0 , \36996_37296 );
xor \U$28523 ( \36998_37298 , 1'b0 , \36997_37297 );
buf \U$28524 ( \36999_37299 , \36998_37298 );
buf \U$28526 ( \37000_37300 , \36999_37299 );
and \U$28527 ( \37001_37301 , \31989_31636 , \17363_17665_nG9bea );
and \U$28528 ( \37002_37302 , \31334_31633 , \17808_18107_nG9be7 );
or \U$28529 ( \37003_37303 , \37001_37301 , \37002_37302 );
xor \U$28530 ( \37004_37304 , \31333_31632 , \37003_37303 );
buf \U$28531 ( \37005_37305 , \37004_37304 );
buf \U$28533 ( \37006_37306 , \37005_37305 );
xor \U$28534 ( \37007_37307 , \37000_37300 , \37006_37306 );
buf \U$28535 ( \37008_37308 , \37007_37307 );
xor \U$28536 ( \37009_37309 , \36995_37295 , \37008_37308 );
and \U$28537 ( \37010_37310 , \27141_26431 , \21827_22129_nG9bd8 );
and \U$28538 ( \37011_37311 , \26129_26428 , \22330_22629_nG9bd5 );
or \U$28539 ( \37012_37312 , \37010_37310 , \37011_37311 );
xor \U$28540 ( \37013_37313 , \26128_26427 , \37012_37312 );
buf \U$28541 ( \37014_37314 , \37013_37313 );
buf \U$28543 ( \37015_37315 , \37014_37314 );
xor \U$28544 ( \37016_37316 , \37009_37309 , \37015_37315 );
buf \U$28545 ( \37017_37317 , \37016_37316 );
and \U$28546 ( \37018_37318 , \17437_17297 , \31877_32179_nG9bb4 );
and \U$28547 ( \37019_37319 , \16995_17294 , \32589_32888_nG9bb1 );
or \U$28548 ( \37020_37320 , \37018_37318 , \37019_37319 );
xor \U$28549 ( \37021_37321 , \16994_17293 , \37020_37320 );
buf \U$28550 ( \37022_37322 , \37021_37321 );
buf \U$28552 ( \37023_37323 , \37022_37322 );
xor \U$28553 ( \37024_37324 , \37017_37317 , \37023_37323 );
and \U$28554 ( \37025_37325 , \13431_13370 , \34343_34643_nG9ba2 );
and \U$28555 ( \37026_37326 , \13068_13367 , \34794_35094_nG9b9f );
or \U$28556 ( \37027_37327 , \37025_37325 , \37026_37326 );
xor \U$28557 ( \37028_37328 , \13067_13366 , \37027_37327 );
buf \U$28558 ( \37029_37329 , \37028_37328 );
buf \U$28560 ( \37030_37330 , \37029_37329 );
xor \U$28561 ( \37031_37331 , \37024_37324 , \37030_37330 );
buf \U$28562 ( \37032_37332 , \37031_37331 );
xor \U$28563 ( \37033_37333 , \36990_37290 , \37032_37332 );
and \U$28564 ( \37034_37334 , \36542_36842 , \36548_36848 );
and \U$28565 ( \37035_37335 , \36542_36842 , \36555_36855 );
and \U$28566 ( \37036_37336 , \36548_36848 , \36555_36855 );
or \U$28567 ( \37037_37337 , \37034_37334 , \37035_37335 , \37036_37336 );
buf \U$28568 ( \37038_37338 , \37037_37337 );
and \U$28569 ( \37039_37339 , \20353_20155 , \28300_28602_nG9bc0 );
and \U$28570 ( \37040_37340 , \19853_20152 , \28877_29179_nG9bbd );
or \U$28571 ( \37041_37341 , \37039_37339 , \37040_37340 );
xor \U$28572 ( \37042_37342 , \19852_20151 , \37041_37341 );
buf \U$28573 ( \37043_37343 , \37042_37342 );
buf \U$28575 ( \37044_37344 , \37043_37343 );
xor \U$28576 ( \37045_37345 , \37038_37338 , \37044_37344 );
and \U$28577 ( \37046_37346 , \16405_15940 , \32881_33181_nG9bae );
and \U$28578 ( \37047_37347 , \15638_15937 , \33313_33613_nG9bab );
or \U$28579 ( \37048_37348 , \37046_37346 , \37047_37347 );
xor \U$28580 ( \37049_37349 , \15637_15936 , \37048_37348 );
buf \U$28581 ( \37050_37350 , \37049_37349 );
buf \U$28583 ( \37051_37351 , \37050_37350 );
xor \U$28584 ( \37052_37352 , \37045_37345 , \37051_37351 );
buf \U$28585 ( \37053_37353 , \37052_37352 );
xor \U$28586 ( \37054_37354 , \37033_37333 , \37053_37353 );
buf \U$28587 ( \37055_37355 , \37054_37354 );
xor \U$28588 ( \37056_37356 , \36985_37285 , \37055_37355 );
and \U$28589 ( \37057_37357 , \36693_36993 , \36713_37013 );
and \U$28590 ( \37058_37358 , \36693_36993 , \36719_37019 );
and \U$28591 ( \37059_37359 , \36713_37013 , \36719_37019 );
or \U$28592 ( \37060_37360 , \37057_37357 , \37058_37358 , \37059_37359 );
buf \U$28593 ( \37061_37361 , \37060_37360 );
xor \U$28594 ( \37062_37362 , \37056_37356 , \37061_37361 );
buf \U$28595 ( \37063_37363 , \37062_37362 );
xor \U$28596 ( \37064_37364 , \36822_37122 , \37063_37363 );
buf \U$28597 ( \37065_37365 , \37064_37364 );
xor \U$28598 ( \37066_37366 , \36743_37043 , \37065_37365 );
and \U$28599 ( \37067_37367 , \36394_36694 , \36399_36699 );
and \U$28600 ( \37068_37368 , \36394_36694 , \36463_36763 );
and \U$28601 ( \37069_37369 , \36399_36699 , \36463_36763 );
or \U$28602 ( \37070_37370 , \37067_37367 , \37068_37368 , \37069_37369 );
buf \U$28603 ( \37071_37371 , \37070_37370 );
xor \U$28604 ( \37072_37372 , \37066_37366 , \37071_37371 );
and \U$28605 ( \37073_37373 , \36738_37038 , \37072_37372 );
and \U$28607 ( \37074_37374 , \36732_37032 , \36737_37037 );
or \U$28609 ( \37075_37375 , 1'b0 , \37074_37374 , 1'b0 );
xor \U$28610 ( \37076_37376 , \37073_37373 , \37075_37375 );
and \U$28612 ( \37077_37377 , \36725_37025 , \36731_37031 );
and \U$28613 ( \37078_37378 , \36727_37027 , \36731_37031 );
or \U$28614 ( \37079_37379 , 1'b0 , \37077_37377 , \37078_37378 );
xor \U$28615 ( \37080_37380 , \37076_37376 , \37079_37379 );
xor \U$28622 ( \37081_37381 , \37080_37380 , 1'b0 );
and \U$28623 ( \37082_37382 , \36743_37043 , \37065_37365 );
and \U$28624 ( \37083_37383 , \36743_37043 , \37071_37371 );
and \U$28625 ( \37084_37384 , \37065_37365 , \37071_37371 );
or \U$28626 ( \37085_37385 , \37082_37382 , \37083_37383 , \37084_37384 );
xor \U$28627 ( \37086_37386 , \37081_37381 , \37085_37385 );
and \U$28628 ( \37087_37387 , \36985_37285 , \37055_37355 );
and \U$28629 ( \37088_37388 , \36985_37285 , \37061_37361 );
and \U$28630 ( \37089_37389 , \37055_37355 , \37061_37361 );
or \U$28631 ( \37090_37390 , \37087_37387 , \37088_37388 , \37089_37389 );
buf \U$28632 ( \37091_37391 , \37090_37390 );
and \U$28633 ( \37092_37392 , \36990_37290 , \37032_37332 );
and \U$28634 ( \37093_37393 , \36990_37290 , \37053_37353 );
and \U$28635 ( \37094_37394 , \37032_37332 , \37053_37353 );
or \U$28636 ( \37095_37395 , \37092_37392 , \37093_37393 , \37094_37394 );
buf \U$28637 ( \37096_37396 , \37095_37395 );
and \U$28638 ( \37097_37397 , \37038_37338 , \37044_37344 );
and \U$28639 ( \37098_37398 , \37038_37338 , \37051_37351 );
and \U$28640 ( \37099_37399 , \37044_37344 , \37051_37351 );
or \U$28641 ( \37100_37400 , \37097_37397 , \37098_37398 , \37099_37399 );
buf \U$28642 ( \37101_37401 , \37100_37400 );
and \U$28643 ( \37102_37402 , \37000_37300 , \37006_37306 );
buf \U$28644 ( \37103_37403 , \37102_37402 );
and \U$28645 ( \37104_37404 , \30670_29853 , \19287_19586_nG9be1 );
and \U$28646 ( \37105_37405 , \29551_29850 , \20306_20608_nG9bde );
or \U$28647 ( \37106_37406 , \37104_37404 , \37105_37405 );
xor \U$28648 ( \37107_37407 , \29550_29849 , \37106_37406 );
buf \U$28649 ( \37108_37408 , \37107_37407 );
buf \U$28651 ( \37109_37409 , \37108_37408 );
xor \U$28652 ( \37110_37410 , \37103_37403 , \37109_37409 );
and \U$28653 ( \37111_37411 , \28946_28118 , \20787_21086_nG9bdb );
and \U$28654 ( \37112_37412 , \27816_28115 , \21827_22129_nG9bd8 );
or \U$28655 ( \37113_37413 , \37111_37411 , \37112_37412 );
xor \U$28656 ( \37114_37414 , \27815_28114 , \37113_37413 );
buf \U$28657 ( \37115_37415 , \37114_37414 );
buf \U$28659 ( \37116_37416 , \37115_37415 );
xor \U$28660 ( \37117_37417 , \37110_37410 , \37116_37416 );
buf \U$28661 ( \37118_37418 , \37117_37417 );
and \U$28662 ( \37119_37419 , \20353_20155 , \28877_29179_nG9bbd );
and \U$28663 ( \37120_37420 , \19853_20152 , \30064_30366_nG9bba );
or \U$28664 ( \37121_37421 , \37119_37419 , \37120_37420 );
xor \U$28665 ( \37122_37422 , \19852_20151 , \37121_37421 );
buf \U$28666 ( \37123_37423 , \37122_37422 );
buf \U$28668 ( \37124_37424 , \37123_37423 );
xor \U$28669 ( \37125_37425 , \37118_37418 , \37124_37424 );
and \U$28670 ( \37126_37426 , \18908_18702 , \30638_30940_nG9bb7 );
and \U$28671 ( \37127_37427 , \18400_18699 , \31877_32179_nG9bb4 );
or \U$28672 ( \37128_37428 , \37126_37426 , \37127_37427 );
xor \U$28673 ( \37129_37429 , \18399_18698 , \37128_37428 );
buf \U$28674 ( \37130_37430 , \37129_37429 );
buf \U$28676 ( \37131_37431 , \37130_37430 );
xor \U$28677 ( \37132_37432 , \37125_37425 , \37131_37431 );
buf \U$28678 ( \37133_37433 , \37132_37432 );
xor \U$28679 ( \37134_37434 , \37101_37401 , \37133_37433 );
and \U$28680 ( \37135_37435 , \37017_37317 , \37023_37323 );
and \U$28681 ( \37136_37436 , \37017_37317 , \37030_37330 );
and \U$28682 ( \37137_37437 , \37023_37323 , \37030_37330 );
or \U$28683 ( \37138_37438 , \37135_37435 , \37136_37436 , \37137_37437 );
buf \U$28684 ( \37139_37439 , \37138_37438 );
xor \U$28685 ( \37140_37440 , \37134_37434 , \37139_37439 );
buf \U$28686 ( \37141_37441 , \37140_37440 );
xor \U$28687 ( \37142_37442 , \37096_37396 , \37141_37441 );
and \U$28688 ( \37143_37443 , \36779_37079 , \36800_37100 );
and \U$28689 ( \37144_37444 , \36779_37079 , \36806_37106 );
and \U$28690 ( \37145_37445 , \36800_37100 , \36806_37106 );
or \U$28691 ( \37146_37446 , \37143_37443 , \37144_37444 , \37145_37445 );
buf \U$28692 ( \37147_37447 , \37146_37446 );
xor \U$28693 ( \37148_37448 , \37142_37442 , \37147_37447 );
buf \U$28694 ( \37149_37449 , \37148_37448 );
xor \U$28695 ( \37150_37450 , \37091_37391 , \37149_37449 );
and \U$28696 ( \37151_37451 , \36748_37048 , \36808_37108 );
and \U$28697 ( \37152_37452 , \36748_37048 , \36814_37114 );
and \U$28698 ( \37153_37453 , \36808_37108 , \36814_37114 );
or \U$28699 ( \37154_37454 , \37151_37451 , \37152_37452 , \37153_37453 );
buf \U$28700 ( \37155_37455 , \37154_37454 );
xor \U$28701 ( \37156_37456 , \37150_37450 , \37155_37455 );
buf \U$28702 ( \37157_37457 , \37156_37456 );
and \U$28703 ( \37158_37458 , \36957_37257 , \36962_37262 );
and \U$28704 ( \37159_37459 , \36957_37257 , \36983_37283 );
and \U$28705 ( \37160_37460 , \36962_37262 , \36983_37283 );
or \U$28706 ( \37161_37461 , \37158_37458 , \37159_37459 , \37160_37460 );
buf \U$28707 ( \37162_37462 , \37161_37461 );
and \U$28708 ( \37163_37463 , \36827_37127 , \36833_37133 );
and \U$28709 ( \37164_37464 , \36827_37127 , \36955_37255 );
and \U$28710 ( \37165_37465 , \36833_37133 , \36955_37255 );
or \U$28711 ( \37166_37466 , \37163_37463 , \37164_37464 , \37165_37465 );
buf \U$28712 ( \37167_37467 , \37166_37466 );
and \U$28713 ( \37168_37468 , \25044_24792 , \23927_24226_nG9bcf );
and \U$28714 ( \37169_37469 , \24490_24789 , \24996_25298_nG9bcc );
or \U$28715 ( \37170_37470 , \37168_37468 , \37169_37469 );
xor \U$28716 ( \37171_37471 , \24489_24788 , \37170_37470 );
buf \U$28717 ( \37172_37472 , \37171_37471 );
buf \U$28719 ( \37173_37473 , \37172_37472 );
and \U$28720 ( \37174_37474 , \23495_23201 , \25561_25860_nG9bc9 );
and \U$28721 ( \37175_37475 , \22899_23198 , \26585_26887_nG9bc6 );
or \U$28722 ( \37176_37476 , \37174_37474 , \37175_37475 );
xor \U$28723 ( \37177_37477 , \22898_23197 , \37176_37476 );
buf \U$28724 ( \37178_37478 , \37177_37477 );
buf \U$28726 ( \37179_37479 , \37178_37478 );
xor \U$28727 ( \37180_37480 , \37173_37473 , \37179_37479 );
and \U$28728 ( \37181_37481 , \21908_21658 , \27114_27416_nG9bc3 );
and \U$28729 ( \37182_37482 , \21356_21655 , \28300_28602_nG9bc0 );
or \U$28730 ( \37183_37483 , \37181_37481 , \37182_37482 );
xor \U$28731 ( \37184_37484 , \21355_21654 , \37183_37483 );
buf \U$28732 ( \37185_37485 , \37184_37484 );
buf \U$28734 ( \37186_37486 , \37185_37485 );
xor \U$28735 ( \37187_37487 , \37180_37480 , \37186_37486 );
buf \U$28736 ( \37188_37488 , \37187_37487 );
and \U$28737 ( \37189_37489 , \10996_10421 , \36289_36589_nG9b93 );
and \U$28738 ( \37190_37490 , \10119_10418 , \36686_36986_nG9b90 );
or \U$28739 ( \37191_37491 , \37189_37489 , \37190_37490 );
xor \U$28740 ( \37192_37492 , \10118_10417 , \37191_37491 );
buf \U$28741 ( \37193_37493 , \37192_37492 );
buf \U$28743 ( \37194_37494 , \37193_37493 );
xor \U$28744 ( \37195_37495 , \37188_37488 , \37194_37494 );
and \U$28745 ( \37196_37496 , \10411_10707 , \36950_37250_nG9b8d );
and \U$28746 ( \37197_37497 , \36912_37212 , \36916_37216 );
and \U$28747 ( \37198_37498 , \36916_37216 , \36938_37238 );
and \U$28748 ( \37199_37499 , \36912_37212 , \36938_37238 );
or \U$28749 ( \37200_37500 , \37197_37497 , \37198_37498 , \37199_37499 );
and \U$28750 ( \37201_37501 , \36847_37147 , \36858_37158 );
and \U$28751 ( \37202_37502 , \36858_37158 , \36873_37173 );
and \U$28752 ( \37203_37503 , \36847_37147 , \36873_37173 );
or \U$28753 ( \37204_37504 , \37201_37501 , \37202_37502 , \37203_37503 );
and \U$28754 ( \37205_37505 , \36879_37179 , \36893_37193 );
and \U$28755 ( \37206_37506 , \36893_37193 , \36905_37205 );
and \U$28756 ( \37207_37507 , \36879_37179 , \36905_37205 );
or \U$28757 ( \37208_37508 , \37205_37505 , \37206_37506 , \37207_37507 );
xor \U$28758 ( \37209_37509 , \37204_37504 , \37208_37508 );
and \U$28759 ( \37210_37510 , \27011_27313 , \22243_22542 );
and \U$28760 ( \37211_37511 , \28232_28534 , \21801_22103 );
nor \U$28761 ( \37212_37512 , \37210_37510 , \37211_37511 );
xnor \U$28762 ( \37213_37513 , \37212_37512 , \22249_22548 );
and \U$28763 ( \37214_37514 , \20734_21033 , \28768_29070 );
and \U$28764 ( \37215_37515 , \21788_22090 , \28224_28526 );
nor \U$28765 ( \37216_37516 , \37214_37514 , \37215_37515 );
xnor \U$28766 ( \37217_37517 , \37216_37516 , \28774_29076 );
xor \U$28767 ( \37218_37518 , \37213_37513 , \37217_37517 );
and \U$28768 ( \37219_37519 , \19259_19558 , \30521_30823 );
and \U$28769 ( \37220_37520 , \20242_20544 , \29944_30246 );
nor \U$28770 ( \37221_37521 , \37219_37519 , \37220_37520 );
xnor \U$28771 ( \37222_37522 , \37221_37521 , \30511_30813 );
xor \U$28772 ( \37223_37523 , \37218_37518 , \37222_37522 );
and \U$28773 ( \37224_37524 , \25516_25815 , \23839_24138 );
and \U$28774 ( \37225_37525 , \26527_26829 , \23328_23630 );
nor \U$28775 ( \37226_37526 , \37224_37524 , \37225_37525 );
xnor \U$28776 ( \37227_37527 , \37226_37526 , \23845_24144 );
and \U$28777 ( \37228_37528 , \17736_18035 , \32555_32854 );
and \U$28778 ( \37229_37529 , \18730_19032 , \31765_32067 );
nor \U$28779 ( \37230_37530 , \37228_37528 , \37229_37529 );
xnor \U$28780 ( \37231_37531 , \37230_37530 , \32506_32805 );
xor \U$28781 ( \37232_37532 , \37227_37527 , \37231_37531 );
and \U$28782 ( \37233_37533 , \17325_17627 , \32503_32802 );
xor \U$28783 ( \37234_37534 , \37232_37532 , \37233_37533 );
xor \U$28784 ( \37235_37535 , \37223_37523 , \37234_37534 );
and \U$28785 ( \37236_37536 , \32495_32794 , \17791_18090 );
not \U$28786 ( \37237_37537 , \37236_37536 );
xnor \U$28787 ( \37238_37538 , \37237_37537 , \17747_18046 );
and \U$28788 ( \37239_37539 , \28782_29084 , \20706_21005 );
and \U$28789 ( \37240_37540 , \29966_30268 , \20255_20557 );
nor \U$28790 ( \37241_37541 , \37239_37539 , \37240_37540 );
xnor \U$28791 ( \37242_37542 , \37241_37541 , \20712_21011 );
xor \U$28792 ( \37243_37543 , \37238_37538 , \37242_37542 );
and \U$28793 ( \37244_37544 , \23900_24199 , \25527_25826 );
and \U$28794 ( \37245_37545 , \24970_25272 , \24962_25264 );
nor \U$28795 ( \37246_37546 , \37244_37544 , \37245_37545 );
xnor \U$28796 ( \37247_37547 , \37246_37546 , \25474_25773 );
xor \U$28797 ( \37248_37548 , \37243_37543 , \37247_37547 );
xor \U$28798 ( \37249_37549 , \37235_37535 , \37248_37548 );
xor \U$28799 ( \37250_37550 , \37209_37509 , \37249_37549 );
xor \U$28800 ( \37251_37551 , \37200_37500 , \37250_37550 );
and \U$28801 ( \37252_37552 , \36921_37221 , \36925_37225 );
and \U$28802 ( \37253_37553 , \36925_37225 , \36937_37237 );
and \U$28803 ( \37254_37554 , \36921_37221 , \36937_37237 );
or \U$28804 ( \37255_37555 , \37252_37552 , \37253_37553 , \37254_37554 );
and \U$28805 ( \37256_37556 , \36843_37143 , \36874_37174 );
and \U$28806 ( \37257_37557 , \36874_37174 , \36906_37206 );
and \U$28807 ( \37258_37558 , \36843_37143 , \36906_37206 );
or \U$28808 ( \37259_37559 , \37256_37556 , \37257_37557 , \37258_37558 );
xor \U$28809 ( \37260_37560 , \37255_37555 , \37259_37559 );
and \U$28810 ( \37261_37561 , \36930_37230 , \36934_37234 );
and \U$28811 ( \37262_37562 , \36934_37234 , \36936_37236 );
and \U$28812 ( \37263_37563 , \36930_37230 , \36936_37236 );
or \U$28813 ( \37264_37564 , \37261_37561 , \37262_37562 , \37263_37563 );
and \U$28814 ( \37265_37565 , \36898_37198 , \36902_37202 );
and \U$28815 ( \37266_37566 , \36902_37202 , \36904_37204 );
and \U$28816 ( \37267_37567 , \36898_37198 , \36904_37204 );
or \U$28817 ( \37268_37568 , \37265_37565 , \37266_37566 , \37267_37567 );
and \U$28818 ( \37269_37569 , \36848_37148 , \36852_37152 );
and \U$28819 ( \37270_37570 , \36852_37152 , \36857_37157 );
and \U$28820 ( \37271_37571 , \36848_37148 , \36857_37157 );
or \U$28821 ( \37272_37572 , \37269_37569 , \37270_37570 , \37271_37571 );
xor \U$28822 ( \37273_37573 , \37268_37568 , \37272_37572 );
and \U$28823 ( \37274_37574 , \36863_37163 , \36867_37167 );
and \U$28824 ( \37275_37575 , \36867_37167 , \36872_37172 );
and \U$28825 ( \37276_37576 , \36863_37163 , \36872_37172 );
or \U$28826 ( \37277_37577 , \37274_37574 , \37275_37575 , \37276_37576 );
xor \U$28827 ( \37278_37578 , \37273_37573 , \37277_37577 );
xor \U$28828 ( \37279_37579 , \37264_37564 , \37278_37578 );
and \U$28829 ( \37280_37580 , \36883_37183 , \36887_37187 );
and \U$28830 ( \37281_37581 , \36887_37187 , \36892_37192 );
and \U$28831 ( \37282_37582 , \36883_37183 , \36892_37192 );
or \U$28832 ( \37283_37583 , \37280_37580 , \37281_37581 , \37282_37582 );
and \U$28833 ( \37284_37584 , \30500_30802 , \19235_19534 );
and \U$28834 ( \37285_37585 , \31752_32054 , \18743_19045 );
nor \U$28835 ( \37286_37586 , \37284_37584 , \37285_37585 );
xnor \U$28836 ( \37287_37587 , \37286_37586 , \19241_19540 );
not \U$28837 ( \37288_37588 , \37287_37587 );
xor \U$28838 ( \37289_37589 , \37283_37583 , \37288_37588 );
and \U$28839 ( \37290_37590 , \22257_22556 , \27095_27397 );
and \U$28840 ( \37291_37591 , \23315_23617 , \26505_26807 );
nor \U$28841 ( \37292_37592 , \37290_37590 , \37291_37591 );
xnor \U$28842 ( \37293_37593 , \37292_37592 , \26993_27295 );
xor \U$28843 ( \37294_37594 , \37289_37589 , \37293_37593 );
xor \U$28844 ( \37295_37595 , \37279_37579 , \37294_37594 );
xor \U$28845 ( \37296_37596 , \37260_37560 , \37295_37595 );
xor \U$28846 ( \37297_37597 , \37251_37551 , \37296_37596 );
and \U$28847 ( \37298_37598 , \36839_37139 , \36907_37207 );
and \U$28848 ( \37299_37599 , \36907_37207 , \36939_37239 );
and \U$28849 ( \37300_37600 , \36839_37139 , \36939_37239 );
or \U$28850 ( \37301_37601 , \37298_37598 , \37299_37599 , \37300_37600 );
xor \U$28851 ( \37302_37602 , \37297_37597 , \37301_37601 );
and \U$28852 ( \37303_37603 , \36940_37240 , \36944_37244 );
and \U$28853 ( \37304_37604 , \36945_37245 , \36948_37248 );
or \U$28854 ( \37305_37605 , \37303_37603 , \37304_37604 );
xor \U$28855 ( \37306_37606 , \37302_37602 , \37305_37605 );
buf g9b8a_GF_PartitionCandidate( \37307_37607_nG9b8a , \37306_37606 );
and \U$28856 ( \37308_37608 , \10402_10704 , \37307_37607_nG9b8a );
or \U$28857 ( \37309_37609 , \37196_37496 , \37308_37608 );
xor \U$28858 ( \37310_37610 , \10399_10703 , \37309_37609 );
buf \U$28859 ( \37311_37611 , \37310_37610 );
buf \U$28861 ( \37312_37612 , \37311_37611 );
xor \U$28862 ( \37313_37613 , \37195_37495 , \37312_37612 );
buf \U$28863 ( \37314_37614 , \37313_37613 );
xor \U$28864 ( \37315_37615 , \37167_37467 , \37314_37614 );
and \U$28865 ( \37316_37616 , \36753_37053 , \36770_37070 );
and \U$28866 ( \37317_37617 , \36753_37053 , \36777_37077 );
and \U$28867 ( \37318_37618 , \36770_37070 , \36777_37077 );
or \U$28868 ( \37319_37619 , \37316_37616 , \37317_37617 , \37318_37618 );
buf \U$28869 ( \37320_37620 , \37319_37619 );
and \U$28870 ( \37321_37621 , \36785_37085 , \36791_37091 );
and \U$28871 ( \37322_37622 , \36785_37085 , \36798_37098 );
and \U$28872 ( \37323_37623 , \36791_37091 , \36798_37098 );
or \U$28873 ( \37324_37624 , \37321_37621 , \37322_37622 , \37323_37623 );
buf \U$28874 ( \37325_37625 , \37324_37624 );
xor \U$28875 ( \37326_37626 , \37320_37620 , \37325_37625 );
and \U$28876 ( \37327_37627 , \12183_12157 , \35501_35801_nG9b99 );
and \U$28877 ( \37328_37628 , \11855_12154 , \35872_36172_nG9b96 );
or \U$28878 ( \37329_37629 , \37327_37627 , \37328_37628 );
xor \U$28879 ( \37330_37630 , \11854_12153 , \37329_37629 );
buf \U$28880 ( \37331_37631 , \37330_37630 );
buf \U$28882 ( \37332_37632 , \37331_37631 );
xor \U$28883 ( \37333_37633 , \37326_37626 , \37332_37632 );
buf \U$28884 ( \37334_37634 , \37333_37633 );
xor \U$28885 ( \37335_37635 , \37315_37615 , \37334_37634 );
buf \U$28886 ( \37336_37636 , \37335_37635 );
xor \U$28887 ( \37337_37637 , \37162_37462 , \37336_37636 );
and \U$28888 ( \37338_37638 , \36968_37268 , \36974_37274 );
and \U$28889 ( \37339_37639 , \36968_37268 , \36981_37281 );
and \U$28890 ( \37340_37640 , \36974_37274 , \36981_37281 );
or \U$28891 ( \37341_37641 , \37338_37638 , \37339_37639 , \37340_37640 );
buf \U$28892 ( \37342_37642 , \37341_37641 );
and \U$28893 ( \37343_37643 , \36995_37295 , \37008_37308 );
and \U$28894 ( \37344_37644 , \36995_37295 , \37015_37315 );
and \U$28895 ( \37345_37645 , \37008_37308 , \37015_37315 );
or \U$28896 ( \37346_37646 , \37343_37643 , \37344_37644 , \37345_37645 );
buf \U$28897 ( \37347_37647 , \37346_37646 );
and \U$28898 ( \37348_37648 , \17437_17297 , \32589_32888_nG9bb1 );
and \U$28899 ( \37349_37649 , \16995_17294 , \32881_33181_nG9bae );
or \U$28900 ( \37350_37650 , \37348_37648 , \37349_37649 );
xor \U$28901 ( \37351_37651 , \16994_17293 , \37350_37650 );
buf \U$28902 ( \37352_37652 , \37351_37651 );
buf \U$28904 ( \37353_37653 , \37352_37652 );
xor \U$28905 ( \37354_37654 , \37347_37647 , \37353_37653 );
and \U$28906 ( \37355_37655 , \16405_15940 , \33313_33613_nG9bab );
and \U$28907 ( \37356_37656 , \15638_15937 , \33741_34041_nG9ba8 );
or \U$28908 ( \37357_37657 , \37355_37655 , \37356_37656 );
xor \U$28909 ( \37358_37658 , \15637_15936 , \37357_37657 );
buf \U$28910 ( \37359_37659 , \37358_37658 );
buf \U$28912 ( \37360_37660 , \37359_37659 );
xor \U$28913 ( \37361_37661 , \37354_37654 , \37360_37660 );
buf \U$28914 ( \37362_37662 , \37361_37661 );
xor \U$28915 ( \37363_37663 , \37342_37642 , \37362_37662 );
and \U$28916 ( \37364_37664 , \36755_37055 , \36761_37061 );
and \U$28917 ( \37365_37665 , \36755_37055 , \36768_37068 );
and \U$28918 ( \37366_37666 , \36761_37061 , \36768_37068 );
or \U$28919 ( \37367_37667 , \37364_37664 , \37365_37665 , \37366_37666 );
buf \U$28920 ( \37368_37668 , \37367_37667 );
and \U$28922 ( \37369_37669 , \32617_32916 , \17363_17665_nG9bea );
or \U$28923 ( \37370_37670 , 1'b0 , \37369_37669 );
xor \U$28924 ( \37371_37671 , 1'b0 , \37370_37670 );
buf \U$28925 ( \37372_37672 , \37371_37671 );
buf \U$28927 ( \37373_37673 , \37372_37672 );
and \U$28928 ( \37374_37674 , \31989_31636 , \17808_18107_nG9be7 );
and \U$28929 ( \37375_37675 , \31334_31633 , \18789_19091_nG9be4 );
or \U$28930 ( \37376_37676 , \37374_37674 , \37375_37675 );
xor \U$28931 ( \37377_37677 , \31333_31632 , \37376_37676 );
buf \U$28932 ( \37378_37678 , \37377_37677 );
buf \U$28934 ( \37379_37679 , \37378_37678 );
xor \U$28935 ( \37380_37680 , \37373_37673 , \37379_37679 );
buf \U$28936 ( \37381_37681 , \37380_37680 );
xor \U$28937 ( \37382_37682 , \37368_37668 , \37381_37681 );
and \U$28938 ( \37383_37683 , \27141_26431 , \22330_22629_nG9bd5 );
and \U$28939 ( \37384_37684 , \26129_26428 , \23394_23696_nG9bd2 );
or \U$28940 ( \37385_37685 , \37383_37683 , \37384_37684 );
xor \U$28941 ( \37386_37686 , \26128_26427 , \37385_37685 );
buf \U$28942 ( \37387_37687 , \37386_37686 );
buf \U$28944 ( \37388_37688 , \37387_37687 );
xor \U$28945 ( \37389_37689 , \37382_37682 , \37388_37688 );
buf \U$28946 ( \37390_37690 , \37389_37689 );
and \U$28947 ( \37391_37691 , \14710_14631 , \33994_34294_nG9ba5 );
and \U$28948 ( \37392_37692 , \14329_14628 , \34343_34643_nG9ba2 );
or \U$28949 ( \37393_37693 , \37391_37691 , \37392_37692 );
xor \U$28950 ( \37394_37694 , \14328_14627 , \37393_37693 );
buf \U$28951 ( \37395_37695 , \37394_37694 );
buf \U$28953 ( \37396_37696 , \37395_37695 );
xor \U$28954 ( \37397_37697 , \37390_37690 , \37396_37696 );
and \U$28955 ( \37398_37698 , \13431_13370 , \34794_35094_nG9b9f );
and \U$28956 ( \37399_37699 , \13068_13367 , \35270_35570_nG9b9c );
or \U$28957 ( \37400_37700 , \37398_37698 , \37399_37699 );
xor \U$28958 ( \37401_37701 , \13067_13366 , \37400_37700 );
buf \U$28959 ( \37402_37702 , \37401_37701 );
buf \U$28961 ( \37403_37703 , \37402_37702 );
xor \U$28962 ( \37404_37704 , \37397_37697 , \37403_37703 );
buf \U$28963 ( \37405_37705 , \37404_37704 );
xor \U$28964 ( \37406_37706 , \37363_37663 , \37405_37705 );
buf \U$28965 ( \37407_37707 , \37406_37706 );
xor \U$28966 ( \37408_37708 , \37337_37637 , \37407_37707 );
buf \U$28967 ( \37409_37709 , \37408_37708 );
xor \U$28968 ( \37410_37710 , \37157_37457 , \37409_37709 );
and \U$28969 ( \37411_37711 , \36816_37116 , \36821_37121 );
and \U$28970 ( \37412_37712 , \36816_37116 , \37063_37363 );
and \U$28971 ( \37413_37713 , \36821_37121 , \37063_37363 );
or \U$28972 ( \37414_37714 , \37411_37711 , \37412_37712 , \37413_37713 );
buf \U$28973 ( \37415_37715 , \37414_37714 );
xor \U$28974 ( \37416_37716 , \37410_37710 , \37415_37715 );
and \U$28975 ( \37417_37717 , \37086_37386 , \37416_37716 );
and \U$28977 ( \37418_37718 , \37080_37380 , \37085_37385 );
or \U$28979 ( \37419_37719 , 1'b0 , \37418_37718 , 1'b0 );
xor \U$28980 ( \37420_37720 , \37417_37717 , \37419_37719 );
and \U$28982 ( \37421_37721 , \37073_37373 , \37079_37379 );
and \U$28983 ( \37422_37722 , \37075_37375 , \37079_37379 );
or \U$28984 ( \37423_37723 , 1'b0 , \37421_37721 , \37422_37722 );
xor \U$28985 ( \37424_37724 , \37420_37720 , \37423_37723 );
xor \U$28992 ( \37425_37725 , \37424_37724 , 1'b0 );
and \U$28993 ( \37426_37726 , \37157_37457 , \37409_37709 );
and \U$28994 ( \37427_37727 , \37157_37457 , \37415_37715 );
and \U$28995 ( \37428_37728 , \37409_37709 , \37415_37715 );
or \U$28996 ( \37429_37729 , \37426_37726 , \37427_37727 , \37428_37728 );
xor \U$28997 ( \37430_37730 , \37425_37725 , \37429_37729 );
and \U$28998 ( \37431_37731 , \37091_37391 , \37149_37449 );
and \U$28999 ( \37432_37732 , \37091_37391 , \37155_37455 );
and \U$29000 ( \37433_37733 , \37149_37449 , \37155_37455 );
or \U$29001 ( \37434_37734 , \37431_37731 , \37432_37732 , \37433_37733 );
buf \U$29002 ( \37435_37735 , \37434_37734 );
and \U$29003 ( \37436_37736 , \37096_37396 , \37141_37441 );
and \U$29004 ( \37437_37737 , \37096_37396 , \37147_37447 );
and \U$29005 ( \37438_37738 , \37141_37441 , \37147_37447 );
or \U$29006 ( \37439_37739 , \37436_37736 , \37437_37737 , \37438_37738 );
buf \U$29007 ( \37440_37740 , \37439_37739 );
and \U$29008 ( \37441_37741 , \37162_37462 , \37336_37636 );
and \U$29009 ( \37442_37742 , \37162_37462 , \37407_37707 );
and \U$29010 ( \37443_37743 , \37336_37636 , \37407_37707 );
or \U$29011 ( \37444_37744 , \37441_37741 , \37442_37742 , \37443_37743 );
buf \U$29012 ( \37445_37745 , \37444_37744 );
xor \U$29013 ( \37446_37746 , \37440_37740 , \37445_37745 );
and \U$29014 ( \37447_37747 , \37101_37401 , \37133_37433 );
and \U$29015 ( \37448_37748 , \37101_37401 , \37139_37439 );
and \U$29016 ( \37449_37749 , \37133_37433 , \37139_37439 );
or \U$29017 ( \37450_37750 , \37447_37747 , \37448_37748 , \37449_37749 );
buf \U$29018 ( \37451_37751 , \37450_37750 );
and \U$29019 ( \37452_37752 , \37342_37642 , \37362_37662 );
and \U$29020 ( \37453_37753 , \37342_37642 , \37405_37705 );
and \U$29021 ( \37454_37754 , \37362_37662 , \37405_37705 );
or \U$29022 ( \37455_37755 , \37452_37752 , \37453_37753 , \37454_37754 );
buf \U$29023 ( \37456_37756 , \37455_37755 );
xor \U$29024 ( \37457_37757 , \37451_37751 , \37456_37756 );
and \U$29026 ( \37458_37758 , \32617_32916 , \17808_18107_nG9be7 );
or \U$29027 ( \37459_37759 , 1'b0 , \37458_37758 );
xor \U$29028 ( \37460_37760 , 1'b0 , \37459_37759 );
buf \U$29029 ( \37461_37761 , \37460_37760 );
buf \U$29031 ( \37462_37762 , \37461_37761 );
and \U$29032 ( \37463_37763 , \30670_29853 , \20306_20608_nG9bde );
and \U$29033 ( \37464_37764 , \29551_29850 , \20787_21086_nG9bdb );
or \U$29034 ( \37465_37765 , \37463_37763 , \37464_37764 );
xor \U$29035 ( \37466_37766 , \29550_29849 , \37465_37765 );
buf \U$29036 ( \37467_37767 , \37466_37766 );
buf \U$29038 ( \37468_37768 , \37467_37767 );
xor \U$29039 ( \37469_37769 , \37462_37762 , \37468_37768 );
buf \U$29040 ( \37470_37770 , \37469_37769 );
and \U$29041 ( \37471_37771 , \37373_37673 , \37379_37679 );
buf \U$29042 ( \37472_37772 , \37471_37771 );
xor \U$29043 ( \37473_37773 , \37470_37770 , \37472_37772 );
and \U$29044 ( \37474_37774 , \31989_31636 , \18789_19091_nG9be4 );
and \U$29045 ( \37475_37775 , \31334_31633 , \19287_19586_nG9be1 );
or \U$29046 ( \37476_37776 , \37474_37774 , \37475_37775 );
xor \U$29047 ( \37477_37777 , \31333_31632 , \37476_37776 );
buf \U$29048 ( \37478_37778 , \37477_37777 );
buf \U$29050 ( \37479_37779 , \37478_37778 );
xor \U$29051 ( \37480_37780 , \37473_37773 , \37479_37779 );
buf \U$29052 ( \37481_37781 , \37480_37780 );
and \U$29053 ( \37482_37782 , \21908_21658 , \28300_28602_nG9bc0 );
and \U$29054 ( \37483_37783 , \21356_21655 , \28877_29179_nG9bbd );
or \U$29055 ( \37484_37784 , \37482_37782 , \37483_37783 );
xor \U$29056 ( \37485_37785 , \21355_21654 , \37484_37784 );
buf \U$29057 ( \37486_37786 , \37485_37785 );
buf \U$29059 ( \37487_37787 , \37486_37786 );
xor \U$29060 ( \37488_37788 , \37481_37781 , \37487_37787 );
and \U$29061 ( \37489_37789 , \18908_18702 , \31877_32179_nG9bb4 );
and \U$29062 ( \37490_37790 , \18400_18699 , \32589_32888_nG9bb1 );
or \U$29063 ( \37491_37791 , \37489_37789 , \37490_37790 );
xor \U$29064 ( \37492_37792 , \18399_18698 , \37491_37791 );
buf \U$29065 ( \37493_37793 , \37492_37792 );
buf \U$29067 ( \37494_37794 , \37493_37793 );
xor \U$29068 ( \37495_37795 , \37488_37788 , \37494_37794 );
buf \U$29069 ( \37496_37796 , \37495_37795 );
and \U$29070 ( \37497_37797 , \37390_37690 , \37396_37696 );
and \U$29071 ( \37498_37798 , \37390_37690 , \37403_37703 );
and \U$29072 ( \37499_37799 , \37396_37696 , \37403_37703 );
or \U$29073 ( \37500_37800 , \37497_37797 , \37498_37798 , \37499_37799 );
buf \U$29074 ( \37501_37801 , \37500_37800 );
xor \U$29075 ( \37502_37802 , \37496_37796 , \37501_37801 );
and \U$29076 ( \37503_37803 , \37347_37647 , \37353_37653 );
and \U$29077 ( \37504_37804 , \37347_37647 , \37360_37660 );
and \U$29078 ( \37505_37805 , \37353_37653 , \37360_37660 );
or \U$29079 ( \37506_37806 , \37503_37803 , \37504_37804 , \37505_37805 );
buf \U$29080 ( \37507_37807 , \37506_37806 );
xor \U$29081 ( \37508_37808 , \37502_37802 , \37507_37807 );
buf \U$29082 ( \37509_37809 , \37508_37808 );
xor \U$29083 ( \37510_37810 , \37457_37757 , \37509_37809 );
buf \U$29084 ( \37511_37811 , \37510_37810 );
xor \U$29085 ( \37512_37812 , \37446_37746 , \37511_37811 );
buf \U$29086 ( \37513_37813 , \37512_37812 );
xor \U$29087 ( \37514_37814 , \37435_37735 , \37513_37813 );
and \U$29088 ( \37515_37815 , \37118_37418 , \37124_37424 );
and \U$29089 ( \37516_37816 , \37118_37418 , \37131_37431 );
and \U$29090 ( \37517_37817 , \37124_37424 , \37131_37431 );
or \U$29091 ( \37518_37818 , \37515_37815 , \37516_37816 , \37517_37817 );
buf \U$29092 ( \37519_37819 , \37518_37818 );
and \U$29093 ( \37520_37820 , \25044_24792 , \24996_25298_nG9bcc );
and \U$29094 ( \37521_37821 , \24490_24789 , \25561_25860_nG9bc9 );
or \U$29095 ( \37522_37822 , \37520_37820 , \37521_37821 );
xor \U$29096 ( \37523_37823 , \24489_24788 , \37522_37822 );
buf \U$29097 ( \37524_37824 , \37523_37823 );
buf \U$29099 ( \37525_37825 , \37524_37824 );
and \U$29100 ( \37526_37826 , \23495_23201 , \26585_26887_nG9bc6 );
and \U$29101 ( \37527_37827 , \22899_23198 , \27114_27416_nG9bc3 );
or \U$29102 ( \37528_37828 , \37526_37826 , \37527_37827 );
xor \U$29103 ( \37529_37829 , \22898_23197 , \37528_37828 );
buf \U$29104 ( \37530_37830 , \37529_37829 );
buf \U$29106 ( \37531_37831 , \37530_37830 );
xor \U$29107 ( \37532_37832 , \37525_37825 , \37531_37831 );
and \U$29108 ( \37533_37833 , \20353_20155 , \30064_30366_nG9bba );
and \U$29109 ( \37534_37834 , \19853_20152 , \30638_30940_nG9bb7 );
or \U$29110 ( \37535_37835 , \37533_37833 , \37534_37834 );
xor \U$29111 ( \37536_37836 , \19852_20151 , \37535_37835 );
buf \U$29112 ( \37537_37837 , \37536_37836 );
buf \U$29114 ( \37538_37838 , \37537_37837 );
xor \U$29115 ( \37539_37839 , \37532_37832 , \37538_37838 );
buf \U$29116 ( \37540_37840 , \37539_37839 );
xor \U$29117 ( \37541_37841 , \37519_37819 , \37540_37840 );
and \U$29118 ( \37542_37842 , \12183_12157 , \35872_36172_nG9b96 );
and \U$29119 ( \37543_37843 , \11855_12154 , \36289_36589_nG9b93 );
or \U$29120 ( \37544_37844 , \37542_37842 , \37543_37843 );
xor \U$29121 ( \37545_37845 , \11854_12153 , \37544_37844 );
buf \U$29122 ( \37546_37846 , \37545_37845 );
buf \U$29124 ( \37547_37847 , \37546_37846 );
xor \U$29125 ( \37548_37848 , \37541_37841 , \37547_37847 );
buf \U$29126 ( \37549_37849 , \37548_37848 );
and \U$29127 ( \37550_37850 , \37188_37488 , \37194_37494 );
and \U$29128 ( \37551_37851 , \37188_37488 , \37312_37612 );
and \U$29129 ( \37552_37852 , \37194_37494 , \37312_37612 );
or \U$29130 ( \37553_37853 , \37550_37850 , \37551_37851 , \37552_37852 );
buf \U$29131 ( \37554_37854 , \37553_37853 );
xor \U$29132 ( \37555_37855 , \37549_37849 , \37554_37854 );
and \U$29133 ( \37556_37856 , \16405_15940 , \33741_34041_nG9ba8 );
and \U$29134 ( \37557_37857 , \15638_15937 , \33994_34294_nG9ba5 );
or \U$29135 ( \37558_37858 , \37556_37856 , \37557_37857 );
xor \U$29136 ( \37559_37859 , \15637_15936 , \37558_37858 );
buf \U$29137 ( \37560_37860 , \37559_37859 );
buf \U$29139 ( \37561_37861 , \37560_37860 );
and \U$29140 ( \37562_37862 , \10996_10421 , \36686_36986_nG9b90 );
and \U$29141 ( \37563_37863 , \10119_10418 , \36950_37250_nG9b8d );
or \U$29142 ( \37564_37864 , \37562_37862 , \37563_37863 );
xor \U$29143 ( \37565_37865 , \10118_10417 , \37564_37864 );
buf \U$29144 ( \37566_37866 , \37565_37865 );
buf \U$29146 ( \37567_37867 , \37566_37866 );
xor \U$29147 ( \37568_37868 , \37561_37861 , \37567_37867 );
and \U$29148 ( \37569_37869 , \10411_10707 , \37307_37607_nG9b8a );
and \U$29149 ( \37570_37870 , \37204_37504 , \37208_37508 );
and \U$29150 ( \37571_37871 , \37208_37508 , \37249_37549 );
and \U$29151 ( \37572_37872 , \37204_37504 , \37249_37549 );
or \U$29152 ( \37573_37873 , \37570_37870 , \37571_37871 , \37572_37872 );
and \U$29153 ( \37574_37874 , \37255_37555 , \37259_37559 );
and \U$29154 ( \37575_37875 , \37259_37559 , \37295_37595 );
and \U$29155 ( \37576_37876 , \37255_37555 , \37295_37595 );
or \U$29156 ( \37577_37877 , \37574_37874 , \37575_37875 , \37576_37876 );
xor \U$29157 ( \37578_37878 , \37573_37873 , \37577_37877 );
and \U$29158 ( \37579_37879 , \37264_37564 , \37278_37578 );
and \U$29159 ( \37580_37880 , \37278_37578 , \37294_37594 );
and \U$29160 ( \37581_37881 , \37264_37564 , \37294_37594 );
or \U$29161 ( \37582_37882 , \37579_37879 , \37580_37880 , \37581_37881 );
and \U$29162 ( \37583_37883 , \37268_37568 , \37272_37572 );
and \U$29163 ( \37584_37884 , \37272_37572 , \37277_37577 );
and \U$29164 ( \37585_37885 , \37268_37568 , \37277_37577 );
or \U$29165 ( \37586_37886 , \37583_37883 , \37584_37884 , \37585_37885 );
and \U$29166 ( \37587_37887 , \37283_37583 , \37288_37588 );
and \U$29167 ( \37588_37888 , \37288_37588 , \37293_37593 );
and \U$29168 ( \37589_37889 , \37283_37583 , \37293_37593 );
or \U$29169 ( \37590_37890 , \37587_37887 , \37588_37888 , \37589_37889 );
xor \U$29170 ( \37591_37891 , \37586_37886 , \37590_37890 );
buf \U$29171 ( \37592_37892 , \37287_37587 );
and \U$29172 ( \37593_37893 , \24970_25272 , \25527_25826 );
and \U$29173 ( \37594_37894 , \25516_25815 , \24962_25264 );
nor \U$29174 ( \37595_37895 , \37593_37893 , \37594_37894 );
xnor \U$29175 ( \37596_37896 , \37595_37895 , \25474_25773 );
xor \U$29176 ( \37597_37897 , \37592_37892 , \37596_37896 );
and \U$29177 ( \37598_37898 , \23315_23617 , \27095_27397 );
and \U$29178 ( \37599_37899 , \23900_24199 , \26505_26807 );
nor \U$29179 ( \37600_37900 , \37598_37898 , \37599_37899 );
xnor \U$29180 ( \37601_37901 , \37600_37900 , \26993_27295 );
xor \U$29181 ( \37602_37902 , \37597_37897 , \37601_37901 );
xor \U$29182 ( \37603_37903 , \37591_37891 , \37602_37902 );
xor \U$29183 ( \37604_37904 , \37582_37882 , \37603_37903 );
and \U$29184 ( \37605_37905 , \37223_37523 , \37234_37534 );
and \U$29185 ( \37606_37906 , \37234_37534 , \37248_37548 );
and \U$29186 ( \37607_37907 , \37223_37523 , \37248_37548 );
or \U$29187 ( \37608_37908 , \37605_37905 , \37606_37906 , \37607_37907 );
and \U$29188 ( \37609_37909 , \37213_37513 , \37217_37517 );
and \U$29189 ( \37610_37910 , \37217_37517 , \37222_37522 );
and \U$29190 ( \37611_37911 , \37213_37513 , \37222_37522 );
or \U$29191 ( \37612_37912 , \37609_37909 , \37610_37910 , \37611_37911 );
and \U$29192 ( \37613_37913 , \37227_37527 , \37231_37531 );
and \U$29193 ( \37614_37914 , \37231_37531 , \37233_37533 );
and \U$29194 ( \37615_37915 , \37227_37527 , \37233_37533 );
or \U$29195 ( \37616_37916 , \37613_37913 , \37614_37914 , \37615_37915 );
xor \U$29196 ( \37617_37917 , \37612_37912 , \37616_37916 );
and \U$29197 ( \37618_37918 , \37238_37538 , \37242_37542 );
and \U$29198 ( \37619_37919 , \37242_37542 , \37247_37547 );
and \U$29199 ( \37620_37920 , \37238_37538 , \37247_37547 );
or \U$29200 ( \37621_37921 , \37618_37918 , \37619_37919 , \37620_37920 );
xor \U$29201 ( \37622_37922 , \37617_37917 , \37621_37921 );
xor \U$29202 ( \37623_37923 , \37608_37908 , \37622_37922 );
and \U$29203 ( \37624_37924 , \29966_30268 , \20706_21005 );
and \U$29204 ( \37625_37925 , \30500_30802 , \20255_20557 );
nor \U$29205 ( \37626_37926 , \37624_37924 , \37625_37925 );
xnor \U$29206 ( \37627_37927 , \37626_37926 , \20712_21011 );
and \U$29207 ( \37628_37928 , \18730_19032 , \32555_32854 );
and \U$29208 ( \37629_37929 , \19259_19558 , \31765_32067 );
nor \U$29209 ( \37630_37930 , \37628_37928 , \37629_37929 );
xnor \U$29210 ( \37631_37931 , \37630_37930 , \32506_32805 );
xor \U$29211 ( \37632_37932 , \37627_37927 , \37631_37931 );
and \U$29212 ( \37633_37933 , \17736_18035 , \32503_32802 );
xor \U$29213 ( \37634_37934 , \37632_37932 , \37633_37933 );
and \U$29214 ( \37635_37935 , \26527_26829 , \23839_24138 );
and \U$29215 ( \37636_37936 , \27011_27313 , \23328_23630 );
nor \U$29216 ( \37637_37937 , \37635_37935 , \37636_37936 );
xnor \U$29217 ( \37638_37938 , \37637_37937 , \23845_24144 );
and \U$29218 ( \37639_37939 , \21788_22090 , \28768_29070 );
and \U$29219 ( \37640_37940 , \22257_22556 , \28224_28526 );
nor \U$29220 ( \37641_37941 , \37639_37939 , \37640_37940 );
xnor \U$29221 ( \37642_37942 , \37641_37941 , \28774_29076 );
xor \U$29222 ( \37643_37943 , \37638_37938 , \37642_37942 );
and \U$29223 ( \37644_37944 , \20242_20544 , \30521_30823 );
and \U$29224 ( \37645_37945 , \20734_21033 , \29944_30246 );
nor \U$29225 ( \37646_37946 , \37644_37944 , \37645_37945 );
xnor \U$29226 ( \37647_37947 , \37646_37946 , \30511_30813 );
xor \U$29227 ( \37648_37948 , \37643_37943 , \37647_37947 );
xor \U$29228 ( \37649_37949 , \37634_37934 , \37648_37948 );
not \U$29229 ( \37650_37950 , \17747_18046 );
and \U$29230 ( \37651_37951 , \31752_32054 , \19235_19534 );
and \U$29231 ( \37652_37952 , \32495_32794 , \18743_19045 );
nor \U$29232 ( \37653_37953 , \37651_37951 , \37652_37952 );
xnor \U$29233 ( \37654_37954 , \37653_37953 , \19241_19540 );
xor \U$29234 ( \37655_37955 , \37650_37950 , \37654_37954 );
and \U$29235 ( \37656_37956 , \28232_28534 , \22243_22542 );
and \U$29236 ( \37657_37957 , \28782_29084 , \21801_22103 );
nor \U$29237 ( \37658_37958 , \37656_37956 , \37657_37957 );
xnor \U$29238 ( \37659_37959 , \37658_37958 , \22249_22548 );
xor \U$29239 ( \37660_37960 , \37655_37955 , \37659_37959 );
xor \U$29240 ( \37661_37961 , \37649_37949 , \37660_37960 );
xor \U$29241 ( \37662_37962 , \37623_37923 , \37661_37961 );
xor \U$29242 ( \37663_37963 , \37604_37904 , \37662_37962 );
xor \U$29243 ( \37664_37964 , \37578_37878 , \37663_37963 );
and \U$29244 ( \37665_37965 , \37200_37500 , \37250_37550 );
and \U$29245 ( \37666_37966 , \37250_37550 , \37296_37596 );
and \U$29246 ( \37667_37967 , \37200_37500 , \37296_37596 );
or \U$29247 ( \37668_37968 , \37665_37965 , \37666_37966 , \37667_37967 );
xor \U$29248 ( \37669_37969 , \37664_37964 , \37668_37968 );
and \U$29249 ( \37670_37970 , \37297_37597 , \37301_37601 );
and \U$29250 ( \37671_37971 , \37302_37602 , \37305_37605 );
or \U$29251 ( \37672_37972 , \37670_37970 , \37671_37971 );
xor \U$29252 ( \37673_37973 , \37669_37969 , \37672_37972 );
buf g9b87_GF_PartitionCandidate( \37674_37974_nG9b87 , \37673_37973 );
and \U$29253 ( \37675_37975 , \10402_10704 , \37674_37974_nG9b87 );
or \U$29254 ( \37676_37976 , \37569_37869 , \37675_37975 );
xor \U$29255 ( \37677_37977 , \10399_10703 , \37676_37976 );
buf \U$29256 ( \37678_37978 , \37677_37977 );
buf \U$29258 ( \37679_37979 , \37678_37978 );
xor \U$29259 ( \37680_37980 , \37568_37868 , \37679_37979 );
buf \U$29260 ( \37681_37981 , \37680_37980 );
xor \U$29261 ( \37682_37982 , \37555_37855 , \37681_37981 );
buf \U$29262 ( \37683_37983 , \37682_37982 );
and \U$29263 ( \37684_37984 , \37320_37620 , \37325_37625 );
and \U$29264 ( \37685_37985 , \37320_37620 , \37332_37632 );
and \U$29265 ( \37686_37986 , \37325_37625 , \37332_37632 );
or \U$29266 ( \37687_37987 , \37684_37984 , \37685_37985 , \37686_37986 );
buf \U$29267 ( \37688_37988 , \37687_37987 );
and \U$29268 ( \37689_37989 , \37368_37668 , \37381_37681 );
and \U$29269 ( \37690_37990 , \37368_37668 , \37388_37688 );
and \U$29270 ( \37691_37991 , \37381_37681 , \37388_37688 );
or \U$29271 ( \37692_37992 , \37689_37989 , \37690_37990 , \37691_37991 );
buf \U$29272 ( \37693_37993 , \37692_37992 );
and \U$29273 ( \37694_37994 , \17437_17297 , \32881_33181_nG9bae );
and \U$29274 ( \37695_37995 , \16995_17294 , \33313_33613_nG9bab );
or \U$29275 ( \37696_37996 , \37694_37994 , \37695_37995 );
xor \U$29276 ( \37697_37997 , \16994_17293 , \37696_37996 );
buf \U$29277 ( \37698_37998 , \37697_37997 );
buf \U$29279 ( \37699_37999 , \37698_37998 );
xor \U$29280 ( \37700_38000 , \37693_37993 , \37699_37999 );
and \U$29281 ( \37701_38001 , \14710_14631 , \34343_34643_nG9ba2 );
and \U$29282 ( \37702_38002 , \14329_14628 , \34794_35094_nG9b9f );
or \U$29283 ( \37703_38003 , \37701_38001 , \37702_38002 );
xor \U$29284 ( \37704_38004 , \14328_14627 , \37703_38003 );
buf \U$29285 ( \37705_38005 , \37704_38004 );
buf \U$29287 ( \37706_38006 , \37705_38005 );
xor \U$29288 ( \37707_38007 , \37700_38000 , \37706_38006 );
buf \U$29289 ( \37708_38008 , \37707_38007 );
xor \U$29290 ( \37709_38009 , \37688_37988 , \37708_38008 );
and \U$29291 ( \37710_38010 , \37173_37473 , \37179_37479 );
and \U$29292 ( \37711_38011 , \37173_37473 , \37186_37486 );
and \U$29293 ( \37712_38012 , \37179_37479 , \37186_37486 );
or \U$29294 ( \37713_38013 , \37710_38010 , \37711_38011 , \37712_38012 );
buf \U$29295 ( \37714_38014 , \37713_38013 );
and \U$29296 ( \37715_38015 , \37103_37403 , \37109_37409 );
and \U$29297 ( \37716_38016 , \37103_37403 , \37116_37416 );
and \U$29298 ( \37717_38017 , \37109_37409 , \37116_37416 );
or \U$29299 ( \37718_38018 , \37715_38015 , \37716_38016 , \37717_38017 );
buf \U$29300 ( \37719_38019 , \37718_38018 );
and \U$29301 ( \37720_38020 , \28946_28118 , \21827_22129_nG9bd8 );
and \U$29302 ( \37721_38021 , \27816_28115 , \22330_22629_nG9bd5 );
or \U$29303 ( \37722_38022 , \37720_38020 , \37721_38021 );
xor \U$29304 ( \37723_38023 , \27815_28114 , \37722_38022 );
buf \U$29305 ( \37724_38024 , \37723_38023 );
buf \U$29307 ( \37725_38025 , \37724_38024 );
xor \U$29308 ( \37726_38026 , \37719_38019 , \37725_38025 );
and \U$29309 ( \37727_38027 , \27141_26431 , \23394_23696_nG9bd2 );
and \U$29310 ( \37728_38028 , \26129_26428 , \23927_24226_nG9bcf );
or \U$29311 ( \37729_38029 , \37727_38027 , \37728_38028 );
xor \U$29312 ( \37730_38030 , \26128_26427 , \37729_38029 );
buf \U$29313 ( \37731_38031 , \37730_38030 );
buf \U$29315 ( \37732_38032 , \37731_38031 );
xor \U$29316 ( \37733_38033 , \37726_38026 , \37732_38032 );
buf \U$29317 ( \37734_38034 , \37733_38033 );
xor \U$29318 ( \37735_38035 , \37714_38014 , \37734_38034 );
and \U$29319 ( \37736_38036 , \13431_13370 , \35270_35570_nG9b9c );
and \U$29320 ( \37737_38037 , \13068_13367 , \35501_35801_nG9b99 );
or \U$29321 ( \37738_38038 , \37736_38036 , \37737_38037 );
xor \U$29322 ( \37739_38039 , \13067_13366 , \37738_38038 );
buf \U$29323 ( \37740_38040 , \37739_38039 );
buf \U$29325 ( \37741_38041 , \37740_38040 );
xor \U$29326 ( \37742_38042 , \37735_38035 , \37741_38041 );
buf \U$29327 ( \37743_38043 , \37742_38042 );
xor \U$29328 ( \37744_38044 , \37709_38009 , \37743_38043 );
buf \U$29329 ( \37745_38045 , \37744_38044 );
xor \U$29330 ( \37746_38046 , \37683_37983 , \37745_38045 );
and \U$29331 ( \37747_38047 , \37167_37467 , \37314_37614 );
and \U$29332 ( \37748_38048 , \37167_37467 , \37334_37634 );
and \U$29333 ( \37749_38049 , \37314_37614 , \37334_37634 );
or \U$29334 ( \37750_38050 , \37747_38047 , \37748_38048 , \37749_38049 );
buf \U$29335 ( \37751_38051 , \37750_38050 );
xor \U$29336 ( \37752_38052 , \37746_38046 , \37751_38051 );
buf \U$29337 ( \37753_38053 , \37752_38052 );
xor \U$29338 ( \37754_38054 , \37514_37814 , \37753_38053 );
and \U$29339 ( \37755_38055 , \37430_37730 , \37754_38054 );
and \U$29341 ( \37756_38056 , \37424_37724 , \37429_37729 );
or \U$29343 ( \37757_38057 , 1'b0 , \37756_38056 , 1'b0 );
xor \U$29344 ( \37758_38058 , \37755_38055 , \37757_38057 );
and \U$29346 ( \37759_38059 , \37417_37717 , \37423_37723 );
and \U$29347 ( \37760_38060 , \37419_37719 , \37423_37723 );
or \U$29348 ( \37761_38061 , 1'b0 , \37759_38059 , \37760_38060 );
xor \U$29349 ( \37762_38062 , \37758_38058 , \37761_38061 );
xor \U$29356 ( \37763_38063 , \37762_38062 , 1'b0 );
and \U$29357 ( \37764_38064 , \37435_37735 , \37513_37813 );
and \U$29358 ( \37765_38065 , \37435_37735 , \37753_38053 );
and \U$29359 ( \37766_38066 , \37513_37813 , \37753_38053 );
or \U$29360 ( \37767_38067 , \37764_38064 , \37765_38065 , \37766_38066 );
xor \U$29361 ( \37768_38068 , \37763_38063 , \37767_38067 );
and \U$29362 ( \37769_38069 , \37683_37983 , \37745_38045 );
and \U$29363 ( \37770_38070 , \37683_37983 , \37751_38051 );
and \U$29364 ( \37771_38071 , \37745_38045 , \37751_38051 );
or \U$29365 ( \37772_38072 , \37769_38069 , \37770_38070 , \37771_38071 );
buf \U$29366 ( \37773_38073 , \37772_38072 );
and \U$29367 ( \37774_38074 , \37496_37796 , \37501_37801 );
and \U$29368 ( \37775_38075 , \37496_37796 , \37507_37807 );
and \U$29369 ( \37776_38076 , \37501_37801 , \37507_37807 );
or \U$29370 ( \37777_38077 , \37774_38074 , \37775_38075 , \37776_38076 );
buf \U$29371 ( \37778_38078 , \37777_38077 );
and \U$29372 ( \37779_38079 , \21908_21658 , \28877_29179_nG9bbd );
and \U$29373 ( \37780_38080 , \21356_21655 , \30064_30366_nG9bba );
or \U$29374 ( \37781_38081 , \37779_38079 , \37780_38080 );
xor \U$29375 ( \37782_38082 , \21355_21654 , \37781_38081 );
buf \U$29376 ( \37783_38083 , \37782_38082 );
buf \U$29378 ( \37784_38084 , \37783_38083 );
and \U$29379 ( \37785_38085 , \18908_18702 , \32589_32888_nG9bb1 );
and \U$29380 ( \37786_38086 , \18400_18699 , \32881_33181_nG9bae );
or \U$29381 ( \37787_38087 , \37785_38085 , \37786_38086 );
xor \U$29382 ( \37788_38088 , \18399_18698 , \37787_38087 );
buf \U$29383 ( \37789_38089 , \37788_38088 );
buf \U$29385 ( \37790_38090 , \37789_38089 );
xor \U$29386 ( \37791_38091 , \37784_38084 , \37790_38090 );
and \U$29387 ( \37792_38092 , \17437_17297 , \33313_33613_nG9bab );
and \U$29388 ( \37793_38093 , \16995_17294 , \33741_34041_nG9ba8 );
or \U$29389 ( \37794_38094 , \37792_38092 , \37793_38093 );
xor \U$29390 ( \37795_38095 , \16994_17293 , \37794_38094 );
buf \U$29391 ( \37796_38096 , \37795_38095 );
buf \U$29393 ( \37797_38097 , \37796_38096 );
xor \U$29394 ( \37798_38098 , \37791_38091 , \37797_38097 );
buf \U$29395 ( \37799_38099 , \37798_38098 );
and \U$29396 ( \37800_38100 , \37714_38014 , \37734_38034 );
and \U$29397 ( \37801_38101 , \37714_38014 , \37741_38041 );
and \U$29398 ( \37802_38102 , \37734_38034 , \37741_38041 );
or \U$29399 ( \37803_38103 , \37800_38100 , \37801_38101 , \37802_38102 );
buf \U$29400 ( \37804_38104 , \37803_38103 );
xor \U$29401 ( \37805_38105 , \37799_38099 , \37804_38104 );
and \U$29402 ( \37806_38106 , \37693_37993 , \37699_37999 );
and \U$29403 ( \37807_38107 , \37693_37993 , \37706_38006 );
and \U$29404 ( \37808_38108 , \37699_37999 , \37706_38006 );
or \U$29405 ( \37809_38109 , \37806_38106 , \37807_38107 , \37808_38108 );
buf \U$29406 ( \37810_38110 , \37809_38109 );
xor \U$29407 ( \37811_38111 , \37805_38105 , \37810_38110 );
buf \U$29408 ( \37812_38112 , \37811_38111 );
xor \U$29409 ( \37813_38113 , \37778_38078 , \37812_38112 );
and \U$29410 ( \37814_38114 , \37688_37988 , \37708_38008 );
and \U$29411 ( \37815_38115 , \37688_37988 , \37743_38043 );
and \U$29412 ( \37816_38116 , \37708_38008 , \37743_38043 );
or \U$29413 ( \37817_38117 , \37814_38114 , \37815_38115 , \37816_38116 );
buf \U$29414 ( \37818_38118 , \37817_38117 );
xor \U$29415 ( \37819_38119 , \37813_38113 , \37818_38118 );
buf \U$29416 ( \37820_38120 , \37819_38119 );
xor \U$29417 ( \37821_38121 , \37773_38073 , \37820_38120 );
and \U$29418 ( \37822_38122 , \37451_37751 , \37456_37756 );
and \U$29419 ( \37823_38123 , \37451_37751 , \37509_37809 );
and \U$29420 ( \37824_38124 , \37456_37756 , \37509_37809 );
or \U$29421 ( \37825_38125 , \37822_38122 , \37823_38123 , \37824_38124 );
buf \U$29422 ( \37826_38126 , \37825_38125 );
xor \U$29423 ( \37827_38127 , \37821_38121 , \37826_38126 );
buf \U$29424 ( \37828_38128 , \37827_38127 );
and \U$29425 ( \37829_38129 , \37440_37740 , \37445_37745 );
and \U$29426 ( \37830_38130 , \37440_37740 , \37511_37811 );
and \U$29427 ( \37831_38131 , \37445_37745 , \37511_37811 );
or \U$29428 ( \37832_38132 , \37829_38129 , \37830_38130 , \37831_38131 );
buf \U$29429 ( \37833_38133 , \37832_38132 );
xor \U$29430 ( \37834_38134 , \37828_38128 , \37833_38133 );
and \U$29431 ( \37835_38135 , \37549_37849 , \37554_37854 );
and \U$29432 ( \37836_38136 , \37549_37849 , \37681_37981 );
and \U$29433 ( \37837_38137 , \37554_37854 , \37681_37981 );
or \U$29434 ( \37838_38138 , \37835_38135 , \37836_38136 , \37837_38137 );
buf \U$29435 ( \37839_38139 , \37838_38138 );
and \U$29436 ( \37840_38140 , \37561_37861 , \37567_37867 );
and \U$29437 ( \37841_38141 , \37561_37861 , \37679_37979 );
and \U$29438 ( \37842_38142 , \37567_37867 , \37679_37979 );
or \U$29439 ( \37843_38143 , \37840_38140 , \37841_38141 , \37842_38142 );
buf \U$29440 ( \37844_38144 , \37843_38143 );
and \U$29441 ( \37845_38145 , \28946_28118 , \22330_22629_nG9bd5 );
and \U$29442 ( \37846_38146 , \27816_28115 , \23394_23696_nG9bd2 );
or \U$29443 ( \37847_38147 , \37845_38145 , \37846_38146 );
xor \U$29444 ( \37848_38148 , \27815_28114 , \37847_38147 );
buf \U$29445 ( \37849_38149 , \37848_38148 );
buf \U$29447 ( \37850_38150 , \37849_38149 );
and \U$29448 ( \37851_38151 , \27141_26431 , \23927_24226_nG9bcf );
and \U$29449 ( \37852_38152 , \26129_26428 , \24996_25298_nG9bcc );
or \U$29450 ( \37853_38153 , \37851_38151 , \37852_38152 );
xor \U$29451 ( \37854_38154 , \26128_26427 , \37853_38153 );
buf \U$29452 ( \37855_38155 , \37854_38154 );
buf \U$29454 ( \37856_38156 , \37855_38155 );
xor \U$29455 ( \37857_38157 , \37850_38150 , \37856_38156 );
and \U$29456 ( \37858_38158 , \25044_24792 , \25561_25860_nG9bc9 );
and \U$29457 ( \37859_38159 , \24490_24789 , \26585_26887_nG9bc6 );
or \U$29458 ( \37860_38160 , \37858_38158 , \37859_38159 );
xor \U$29459 ( \37861_38161 , \24489_24788 , \37860_38160 );
buf \U$29460 ( \37862_38162 , \37861_38161 );
buf \U$29462 ( \37863_38163 , \37862_38162 );
xor \U$29463 ( \37864_38164 , \37857_38157 , \37863_38163 );
buf \U$29464 ( \37865_38165 , \37864_38164 );
and \U$29465 ( \37866_38166 , \16405_15940 , \33994_34294_nG9ba5 );
and \U$29466 ( \37867_38167 , \15638_15937 , \34343_34643_nG9ba2 );
or \U$29467 ( \37868_38168 , \37866_38166 , \37867_38167 );
xor \U$29468 ( \37869_38169 , \15637_15936 , \37868_38168 );
buf \U$29469 ( \37870_38170 , \37869_38169 );
buf \U$29471 ( \37871_38171 , \37870_38170 );
xor \U$29472 ( \37872_38172 , \37865_38165 , \37871_38171 );
and \U$29473 ( \37873_38173 , \13431_13370 , \35501_35801_nG9b99 );
and \U$29474 ( \37874_38174 , \13068_13367 , \35872_36172_nG9b96 );
or \U$29475 ( \37875_38175 , \37873_38173 , \37874_38174 );
xor \U$29476 ( \37876_38176 , \13067_13366 , \37875_38175 );
buf \U$29477 ( \37877_38177 , \37876_38176 );
buf \U$29479 ( \37878_38178 , \37877_38177 );
xor \U$29480 ( \37879_38179 , \37872_38172 , \37878_38178 );
buf \U$29481 ( \37880_38180 , \37879_38179 );
xor \U$29482 ( \37881_38181 , \37844_38144 , \37880_38180 );
and \U$29483 ( \37882_38182 , \37519_37819 , \37540_37840 );
and \U$29484 ( \37883_38183 , \37519_37819 , \37547_37847 );
and \U$29485 ( \37884_38184 , \37540_37840 , \37547_37847 );
or \U$29486 ( \37885_38185 , \37882_38182 , \37883_38183 , \37884_38184 );
buf \U$29487 ( \37886_38186 , \37885_38185 );
xor \U$29488 ( \37887_38187 , \37881_38181 , \37886_38186 );
buf \U$29489 ( \37888_38188 , \37887_38187 );
xor \U$29490 ( \37889_38189 , \37839_38139 , \37888_38188 );
and \U$29491 ( \37890_38190 , \37481_37781 , \37487_37787 );
and \U$29492 ( \37891_38191 , \37481_37781 , \37494_37794 );
and \U$29493 ( \37892_38192 , \37487_37787 , \37494_37794 );
or \U$29494 ( \37893_38193 , \37890_38190 , \37891_38191 , \37892_38192 );
buf \U$29495 ( \37894_38194 , \37893_38193 );
and \U$29496 ( \37895_38195 , \37470_37770 , \37472_37772 );
and \U$29497 ( \37896_38196 , \37470_37770 , \37479_37779 );
and \U$29498 ( \37897_38197 , \37472_37772 , \37479_37779 );
or \U$29499 ( \37898_38198 , \37895_38195 , \37896_38196 , \37897_38197 );
buf \U$29500 ( \37899_38199 , \37898_38198 );
and \U$29501 ( \37900_38200 , \23495_23201 , \27114_27416_nG9bc3 );
and \U$29502 ( \37901_38201 , \22899_23198 , \28300_28602_nG9bc0 );
or \U$29503 ( \37902_38202 , \37900_38200 , \37901_38201 );
xor \U$29504 ( \37903_38203 , \22898_23197 , \37902_38202 );
buf \U$29505 ( \37904_38204 , \37903_38203 );
buf \U$29507 ( \37905_38205 , \37904_38204 );
xor \U$29508 ( \37906_38206 , \37899_38199 , \37905_38205 );
and \U$29509 ( \37907_38207 , \20353_20155 , \30638_30940_nG9bb7 );
and \U$29510 ( \37908_38208 , \19853_20152 , \31877_32179_nG9bb4 );
or \U$29511 ( \37909_38209 , \37907_38207 , \37908_38208 );
xor \U$29512 ( \37910_38210 , \19852_20151 , \37909_38209 );
buf \U$29513 ( \37911_38211 , \37910_38210 );
buf \U$29515 ( \37912_38212 , \37911_38211 );
xor \U$29516 ( \37913_38213 , \37906_38206 , \37912_38212 );
buf \U$29517 ( \37914_38214 , \37913_38213 );
xor \U$29518 ( \37915_38215 , \37894_38194 , \37914_38214 );
and \U$29519 ( \37916_38216 , \12183_12157 , \36289_36589_nG9b93 );
and \U$29520 ( \37917_38217 , \11855_12154 , \36686_36986_nG9b90 );
or \U$29521 ( \37918_38218 , \37916_38216 , \37917_38217 );
xor \U$29522 ( \37919_38219 , \11854_12153 , \37918_38218 );
buf \U$29523 ( \37920_38220 , \37919_38219 );
buf \U$29525 ( \37921_38221 , \37920_38220 );
xor \U$29526 ( \37922_38222 , \37915_38215 , \37921_38221 );
buf \U$29527 ( \37923_38223 , \37922_38222 );
and \U$29528 ( \37924_38224 , \37525_37825 , \37531_37831 );
and \U$29529 ( \37925_38225 , \37525_37825 , \37538_37838 );
and \U$29530 ( \37926_38226 , \37531_37831 , \37538_37838 );
or \U$29531 ( \37927_38227 , \37924_38224 , \37925_38225 , \37926_38226 );
buf \U$29532 ( \37928_38228 , \37927_38227 );
and \U$29533 ( \37929_38229 , \10996_10421 , \36950_37250_nG9b8d );
and \U$29534 ( \37930_38230 , \10119_10418 , \37307_37607_nG9b8a );
or \U$29535 ( \37931_38231 , \37929_38229 , \37930_38230 );
xor \U$29536 ( \37932_38232 , \10118_10417 , \37931_38231 );
buf \U$29537 ( \37933_38233 , \37932_38232 );
buf \U$29539 ( \37934_38234 , \37933_38233 );
xor \U$29540 ( \37935_38235 , \37928_38228 , \37934_38234 );
and \U$29541 ( \37936_38236 , \10411_10707 , \37674_37974_nG9b87 );
and \U$29542 ( \37937_38237 , \37582_37882 , \37603_37903 );
and \U$29543 ( \37938_38238 , \37603_37903 , \37662_37962 );
and \U$29544 ( \37939_38239 , \37582_37882 , \37662_37962 );
or \U$29545 ( \37940_38240 , \37937_38237 , \37938_38238 , \37939_38239 );
and \U$29546 ( \37941_38241 , \37634_37934 , \37648_37948 );
and \U$29547 ( \37942_38242 , \37648_37948 , \37660_37960 );
and \U$29548 ( \37943_38243 , \37634_37934 , \37660_37960 );
or \U$29549 ( \37944_38244 , \37941_38241 , \37942_38242 , \37943_38243 );
and \U$29550 ( \37945_38245 , \37638_37938 , \37642_37942 );
and \U$29551 ( \37946_38246 , \37642_37942 , \37647_37947 );
and \U$29552 ( \37947_38247 , \37638_37938 , \37647_37947 );
or \U$29553 ( \37948_38248 , \37945_38245 , \37946_38246 , \37947_38247 );
and \U$29554 ( \37949_38249 , \37650_37950 , \37654_37954 );
and \U$29555 ( \37950_38250 , \37654_37954 , \37659_37959 );
and \U$29556 ( \37951_38251 , \37650_37950 , \37659_37959 );
or \U$29557 ( \37952_38252 , \37949_38249 , \37950_38250 , \37951_38251 );
xor \U$29558 ( \37953_38253 , \37948_38248 , \37952_38252 );
and \U$29559 ( \37954_38254 , \32495_32794 , \19235_19534 );
not \U$29560 ( \37955_38255 , \37954_38254 );
xnor \U$29561 ( \37956_38256 , \37955_38255 , \19241_19540 );
not \U$29562 ( \37957_38257 , \37956_38256 );
xor \U$29563 ( \37958_38258 , \37953_38253 , \37957_38257 );
xor \U$29564 ( \37959_38259 , \37944_38244 , \37958_38258 );
and \U$29565 ( \37960_38260 , \37627_37927 , \37631_37931 );
and \U$29566 ( \37961_38261 , \37631_37931 , \37633_37933 );
and \U$29567 ( \37962_38262 , \37627_37927 , \37633_37933 );
or \U$29568 ( \37963_38263 , \37960_38260 , \37961_38261 , \37962_38262 );
and \U$29569 ( \37964_38264 , \30500_30802 , \20706_21005 );
and \U$29570 ( \37965_38265 , \31752_32054 , \20255_20557 );
nor \U$29571 ( \37966_38266 , \37964_38264 , \37965_38265 );
xnor \U$29572 ( \37967_38267 , \37966_38266 , \20712_21011 );
and \U$29573 ( \37968_38268 , \25516_25815 , \25527_25826 );
and \U$29574 ( \37969_38269 , \26527_26829 , \24962_25264 );
nor \U$29575 ( \37970_38270 , \37968_38268 , \37969_38269 );
xnor \U$29576 ( \37971_38271 , \37970_38270 , \25474_25773 );
xor \U$29577 ( \37972_38272 , \37967_38267 , \37971_38271 );
and \U$29578 ( \37973_38273 , \18730_19032 , \32503_32802 );
xor \U$29579 ( \37974_38274 , \37972_38272 , \37973_38273 );
xor \U$29580 ( \37975_38275 , \37963_38263 , \37974_38274 );
and \U$29581 ( \37976_38276 , \27011_27313 , \23839_24138 );
and \U$29582 ( \37977_38277 , \28232_28534 , \23328_23630 );
nor \U$29583 ( \37978_38278 , \37976_38276 , \37977_38277 );
xnor \U$29584 ( \37979_38279 , \37978_38278 , \23845_24144 );
and \U$29585 ( \37980_38280 , \20734_21033 , \30521_30823 );
and \U$29586 ( \37981_38281 , \21788_22090 , \29944_30246 );
nor \U$29587 ( \37982_38282 , \37980_38280 , \37981_38281 );
xnor \U$29588 ( \37983_38283 , \37982_38282 , \30511_30813 );
xor \U$29589 ( \37984_38284 , \37979_38279 , \37983_38283 );
and \U$29590 ( \37985_38285 , \19259_19558 , \32555_32854 );
and \U$29591 ( \37986_38286 , \20242_20544 , \31765_32067 );
nor \U$29592 ( \37987_38287 , \37985_38285 , \37986_38286 );
xnor \U$29593 ( \37988_38288 , \37987_38287 , \32506_32805 );
xor \U$29594 ( \37989_38289 , \37984_38284 , \37988_38288 );
xor \U$29595 ( \37990_38290 , \37975_38275 , \37989_38289 );
xor \U$29596 ( \37991_38291 , \37959_38259 , \37990_38290 );
xor \U$29597 ( \37992_38292 , \37940_38240 , \37991_38291 );
and \U$29598 ( \37993_38293 , \37586_37886 , \37590_37890 );
and \U$29599 ( \37994_38294 , \37590_37890 , \37602_37902 );
and \U$29600 ( \37995_38295 , \37586_37886 , \37602_37902 );
or \U$29601 ( \37996_38296 , \37993_38293 , \37994_38294 , \37995_38295 );
and \U$29602 ( \37997_38297 , \37608_37908 , \37622_37922 );
and \U$29603 ( \37998_38298 , \37622_37922 , \37661_37961 );
and \U$29604 ( \37999_38299 , \37608_37908 , \37661_37961 );
or \U$29605 ( \38000_38300 , \37997_38297 , \37998_38298 , \37999_38299 );
xor \U$29606 ( \38001_38301 , \37996_38296 , \38000_38300 );
and \U$29607 ( \38002_38302 , \37612_37912 , \37616_37916 );
and \U$29608 ( \38003_38303 , \37616_37916 , \37621_37921 );
and \U$29609 ( \38004_38304 , \37612_37912 , \37621_37921 );
or \U$29610 ( \38005_38305 , \38002_38302 , \38003_38303 , \38004_38304 );
and \U$29611 ( \38006_38306 , \37592_37892 , \37596_37896 );
and \U$29612 ( \38007_38307 , \37596_37896 , \37601_37901 );
and \U$29613 ( \38008_38308 , \37592_37892 , \37601_37901 );
or \U$29614 ( \38009_38309 , \38006_38306 , \38007_38307 , \38008_38308 );
xor \U$29615 ( \38010_38310 , \38005_38305 , \38009_38309 );
and \U$29616 ( \38011_38311 , \28782_29084 , \22243_22542 );
and \U$29617 ( \38012_38312 , \29966_30268 , \21801_22103 );
nor \U$29618 ( \38013_38313 , \38011_38311 , \38012_38312 );
xnor \U$29619 ( \38014_38314 , \38013_38313 , \22249_22548 );
and \U$29620 ( \38015_38315 , \23900_24199 , \27095_27397 );
and \U$29621 ( \38016_38316 , \24970_25272 , \26505_26807 );
nor \U$29622 ( \38017_38317 , \38015_38315 , \38016_38316 );
xnor \U$29623 ( \38018_38318 , \38017_38317 , \26993_27295 );
xor \U$29624 ( \38019_38319 , \38014_38314 , \38018_38318 );
and \U$29625 ( \38020_38320 , \22257_22556 , \28768_29070 );
and \U$29626 ( \38021_38321 , \23315_23617 , \28224_28526 );
nor \U$29627 ( \38022_38322 , \38020_38320 , \38021_38321 );
xnor \U$29628 ( \38023_38323 , \38022_38322 , \28774_29076 );
xor \U$29629 ( \38024_38324 , \38019_38319 , \38023_38323 );
xor \U$29630 ( \38025_38325 , \38010_38310 , \38024_38324 );
xor \U$29631 ( \38026_38326 , \38001_38301 , \38025_38325 );
xor \U$29632 ( \38027_38327 , \37992_38292 , \38026_38326 );
and \U$29633 ( \38028_38328 , \37573_37873 , \37577_37877 );
and \U$29634 ( \38029_38329 , \37577_37877 , \37663_37963 );
and \U$29635 ( \38030_38330 , \37573_37873 , \37663_37963 );
or \U$29636 ( \38031_38331 , \38028_38328 , \38029_38329 , \38030_38330 );
xor \U$29637 ( \38032_38332 , \38027_38327 , \38031_38331 );
and \U$29638 ( \38033_38333 , \37664_37964 , \37668_37968 );
and \U$29639 ( \38034_38334 , \37669_37969 , \37672_37972 );
or \U$29640 ( \38035_38335 , \38033_38333 , \38034_38334 );
xor \U$29641 ( \38036_38336 , \38032_38332 , \38035_38335 );
buf g9b84_GF_PartitionCandidate( \38037_38337_nG9b84 , \38036_38336 );
and \U$29642 ( \38038_38338 , \10402_10704 , \38037_38337_nG9b84 );
or \U$29643 ( \38039_38339 , \37936_38236 , \38038_38338 );
xor \U$29644 ( \38040_38340 , \10399_10703 , \38039_38339 );
buf \U$29645 ( \38041_38341 , \38040_38340 );
buf \U$29647 ( \38042_38342 , \38041_38341 );
xor \U$29648 ( \38043_38343 , \37935_38235 , \38042_38342 );
buf \U$29649 ( \38044_38344 , \38043_38343 );
xor \U$29650 ( \38045_38345 , \37923_38223 , \38044_38344 );
and \U$29651 ( \38046_38346 , \37719_38019 , \37725_38025 );
and \U$29652 ( \38047_38347 , \37719_38019 , \37732_38032 );
and \U$29653 ( \38048_38348 , \37725_38025 , \37732_38032 );
or \U$29654 ( \38049_38349 , \38046_38346 , \38047_38347 , \38048_38348 );
buf \U$29655 ( \38050_38350 , \38049_38349 );
and \U$29657 ( \38051_38351 , \32617_32916 , \18789_19091_nG9be4 );
or \U$29658 ( \38052_38352 , 1'b0 , \38051_38351 );
xor \U$29659 ( \38053_38353 , 1'b0 , \38052_38352 );
buf \U$29660 ( \38054_38354 , \38053_38353 );
buf \U$29662 ( \38055_38355 , \38054_38354 );
and \U$29663 ( \38056_38356 , \30670_29853 , \20787_21086_nG9bdb );
and \U$29664 ( \38057_38357 , \29551_29850 , \21827_22129_nG9bd8 );
or \U$29665 ( \38058_38358 , \38056_38356 , \38057_38357 );
xor \U$29666 ( \38059_38359 , \29550_29849 , \38058_38358 );
buf \U$29667 ( \38060_38360 , \38059_38359 );
buf \U$29669 ( \38061_38361 , \38060_38360 );
xor \U$29670 ( \38062_38362 , \38055_38355 , \38061_38361 );
buf \U$29671 ( \38063_38363 , \38062_38362 );
and \U$29672 ( \38064_38364 , \37462_37762 , \37468_37768 );
buf \U$29673 ( \38065_38365 , \38064_38364 );
xor \U$29674 ( \38066_38366 , \38063_38363 , \38065_38365 );
and \U$29675 ( \38067_38367 , \31989_31636 , \19287_19586_nG9be1 );
and \U$29676 ( \38068_38368 , \31334_31633 , \20306_20608_nG9bde );
or \U$29677 ( \38069_38369 , \38067_38367 , \38068_38368 );
xor \U$29678 ( \38070_38370 , \31333_31632 , \38069_38369 );
buf \U$29679 ( \38071_38371 , \38070_38370 );
buf \U$29681 ( \38072_38372 , \38071_38371 );
xor \U$29682 ( \38073_38373 , \38066_38366 , \38072_38372 );
buf \U$29683 ( \38074_38374 , \38073_38373 );
xor \U$29684 ( \38075_38375 , \38050_38350 , \38074_38374 );
and \U$29685 ( \38076_38376 , \14710_14631 , \34794_35094_nG9b9f );
and \U$29686 ( \38077_38377 , \14329_14628 , \35270_35570_nG9b9c );
or \U$29687 ( \38078_38378 , \38076_38376 , \38077_38377 );
xor \U$29688 ( \38079_38379 , \14328_14627 , \38078_38378 );
buf \U$29689 ( \38080_38380 , \38079_38379 );
buf \U$29691 ( \38081_38381 , \38080_38380 );
xor \U$29692 ( \38082_38382 , \38075_38375 , \38081_38381 );
buf \U$29693 ( \38083_38383 , \38082_38382 );
xor \U$29694 ( \38084_38384 , \38045_38345 , \38083_38383 );
buf \U$29695 ( \38085_38385 , \38084_38384 );
xor \U$29696 ( \38086_38386 , \37889_38189 , \38085_38385 );
buf \U$29697 ( \38087_38387 , \38086_38386 );
xor \U$29698 ( \38088_38388 , \37834_38134 , \38087_38387 );
and \U$29699 ( \38089_38389 , \37768_38068 , \38088_38388 );
and \U$29701 ( \38090_38390 , \37762_38062 , \37767_38067 );
or \U$29703 ( \38091_38391 , 1'b0 , \38090_38390 , 1'b0 );
xor \U$29704 ( \38092_38392 , \38089_38389 , \38091_38391 );
and \U$29706 ( \38093_38393 , \37755_38055 , \37761_38061 );
and \U$29707 ( \38094_38394 , \37757_38057 , \37761_38061 );
or \U$29708 ( \38095_38395 , 1'b0 , \38093_38393 , \38094_38394 );
xor \U$29709 ( \38096_38396 , \38092_38392 , \38095_38395 );
xor \U$29716 ( \38097_38397 , \38096_38396 , 1'b0 );
and \U$29717 ( \38098_38398 , \37865_38165 , \37871_38171 );
and \U$29718 ( \38099_38399 , \37865_38165 , \37878_38178 );
and \U$29719 ( \38100_38400 , \37871_38171 , \37878_38178 );
or \U$29720 ( \38101_38401 , \38098_38398 , \38099_38399 , \38100_38400 );
buf \U$29721 ( \38102_38402 , \38101_38401 );
and \U$29722 ( \38103_38403 , \38050_38350 , \38074_38374 );
and \U$29723 ( \38104_38404 , \38050_38350 , \38081_38381 );
and \U$29724 ( \38105_38405 , \38074_38374 , \38081_38381 );
or \U$29725 ( \38106_38406 , \38103_38403 , \38104_38404 , \38105_38405 );
buf \U$29726 ( \38107_38407 , \38106_38406 );
xor \U$29727 ( \38108_38408 , \38102_38402 , \38107_38407 );
and \U$29729 ( \38109_38409 , \32617_32916 , \19287_19586_nG9be1 );
or \U$29730 ( \38110_38410 , 1'b0 , \38109_38409 );
xor \U$29731 ( \38111_38411 , 1'b0 , \38110_38410 );
buf \U$29732 ( \38112_38412 , \38111_38411 );
buf \U$29734 ( \38113_38413 , \38112_38412 );
and \U$29735 ( \38114_38414 , \31989_31636 , \20306_20608_nG9bde );
and \U$29736 ( \38115_38415 , \31334_31633 , \20787_21086_nG9bdb );
or \U$29737 ( \38116_38416 , \38114_38414 , \38115_38415 );
xor \U$29738 ( \38117_38417 , \31333_31632 , \38116_38416 );
buf \U$29739 ( \38118_38418 , \38117_38417 );
buf \U$29741 ( \38119_38419 , \38118_38418 );
xor \U$29742 ( \38120_38420 , \38113_38413 , \38119_38419 );
buf \U$29743 ( \38121_38421 , \38120_38420 );
and \U$29744 ( \38122_38422 , \38055_38355 , \38061_38361 );
buf \U$29745 ( \38123_38423 , \38122_38422 );
xor \U$29746 ( \38124_38424 , \38121_38421 , \38123_38423 );
and \U$29747 ( \38125_38425 , \30670_29853 , \21827_22129_nG9bd8 );
and \U$29748 ( \38126_38426 , \29551_29850 , \22330_22629_nG9bd5 );
or \U$29749 ( \38127_38427 , \38125_38425 , \38126_38426 );
xor \U$29750 ( \38128_38428 , \29550_29849 , \38127_38427 );
buf \U$29751 ( \38129_38429 , \38128_38428 );
buf \U$29753 ( \38130_38430 , \38129_38429 );
xor \U$29754 ( \38131_38431 , \38124_38424 , \38130_38430 );
buf \U$29755 ( \38132_38432 , \38131_38431 );
and \U$29756 ( \38133_38433 , \20353_20155 , \31877_32179_nG9bb4 );
and \U$29757 ( \38134_38434 , \19853_20152 , \32589_32888_nG9bb1 );
or \U$29758 ( \38135_38435 , \38133_38433 , \38134_38434 );
xor \U$29759 ( \38136_38436 , \19852_20151 , \38135_38435 );
buf \U$29760 ( \38137_38437 , \38136_38436 );
buf \U$29762 ( \38138_38438 , \38137_38437 );
xor \U$29763 ( \38139_38439 , \38132_38432 , \38138_38438 );
and \U$29764 ( \38140_38440 , \18908_18702 , \32881_33181_nG9bae );
and \U$29765 ( \38141_38441 , \18400_18699 , \33313_33613_nG9bab );
or \U$29766 ( \38142_38442 , \38140_38440 , \38141_38441 );
xor \U$29767 ( \38143_38443 , \18399_18698 , \38142_38442 );
buf \U$29768 ( \38144_38444 , \38143_38443 );
buf \U$29770 ( \38145_38445 , \38144_38444 );
xor \U$29771 ( \38146_38446 , \38139_38439 , \38145_38445 );
buf \U$29772 ( \38147_38447 , \38146_38446 );
xor \U$29773 ( \38148_38448 , \38108_38408 , \38147_38447 );
buf \U$29774 ( \38149_38449 , \38148_38448 );
and \U$29775 ( \38150_38450 , \37844_38144 , \37880_38180 );
and \U$29776 ( \38151_38451 , \37844_38144 , \37886_38186 );
and \U$29777 ( \38152_38452 , \37880_38180 , \37886_38186 );
or \U$29778 ( \38153_38453 , \38150_38450 , \38151_38451 , \38152_38452 );
buf \U$29779 ( \38154_38454 , \38153_38453 );
xor \U$29780 ( \38155_38455 , \38149_38449 , \38154_38454 );
and \U$29781 ( \38156_38456 , \37799_38099 , \37804_38104 );
and \U$29782 ( \38157_38457 , \37799_38099 , \37810_38110 );
and \U$29783 ( \38158_38458 , \37804_38104 , \37810_38110 );
or \U$29784 ( \38159_38459 , \38156_38456 , \38157_38457 , \38158_38458 );
buf \U$29785 ( \38160_38460 , \38159_38459 );
xor \U$29786 ( \38161_38461 , \38155_38455 , \38160_38460 );
buf \U$29787 ( \38162_38462 , \38161_38461 );
and \U$29788 ( \38163_38463 , \37778_38078 , \37812_38112 );
and \U$29789 ( \38164_38464 , \37778_38078 , \37818_38118 );
and \U$29790 ( \38165_38465 , \37812_38112 , \37818_38118 );
or \U$29791 ( \38166_38466 , \38163_38463 , \38164_38464 , \38165_38465 );
buf \U$29792 ( \38167_38467 , \38166_38466 );
xor \U$29793 ( \38168_38468 , \38162_38462 , \38167_38467 );
and \U$29794 ( \38169_38469 , \37839_38139 , \37888_38188 );
and \U$29795 ( \38170_38470 , \37839_38139 , \38085_38385 );
and \U$29796 ( \38171_38471 , \37888_38188 , \38085_38385 );
or \U$29797 ( \38172_38472 , \38169_38469 , \38170_38470 , \38171_38471 );
buf \U$29798 ( \38173_38473 , \38172_38472 );
xor \U$29799 ( \38174_38474 , \38168_38468 , \38173_38473 );
buf \U$29800 ( \38175_38475 , \38174_38474 );
and \U$29801 ( \38176_38476 , \37773_38073 , \37820_38120 );
and \U$29802 ( \38177_38477 , \37773_38073 , \37826_38126 );
and \U$29803 ( \38178_38478 , \37820_38120 , \37826_38126 );
or \U$29804 ( \38179_38479 , \38176_38476 , \38177_38477 , \38178_38478 );
buf \U$29805 ( \38180_38480 , \38179_38479 );
xor \U$29806 ( \38181_38481 , \38175_38475 , \38180_38480 );
and \U$29807 ( \38182_38482 , \37923_38223 , \38044_38344 );
and \U$29808 ( \38183_38483 , \37923_38223 , \38083_38383 );
and \U$29809 ( \38184_38484 , \38044_38344 , \38083_38383 );
or \U$29810 ( \38185_38485 , \38182_38482 , \38183_38483 , \38184_38484 );
buf \U$29811 ( \38186_38486 , \38185_38485 );
and \U$29812 ( \38187_38487 , \37894_38194 , \37914_38214 );
and \U$29813 ( \38188_38488 , \37894_38194 , \37921_38221 );
and \U$29814 ( \38189_38489 , \37914_38214 , \37921_38221 );
or \U$29815 ( \38190_38490 , \38187_38487 , \38188_38488 , \38189_38489 );
buf \U$29816 ( \38191_38491 , \38190_38490 );
and \U$29817 ( \38192_38492 , \37928_38228 , \37934_38234 );
and \U$29818 ( \38193_38493 , \37928_38228 , \38042_38342 );
and \U$29819 ( \38194_38494 , \37934_38234 , \38042_38342 );
or \U$29820 ( \38195_38495 , \38192_38492 , \38193_38493 , \38194_38494 );
buf \U$29821 ( \38196_38496 , \38195_38495 );
xor \U$29822 ( \38197_38497 , \38191_38491 , \38196_38496 );
and \U$29823 ( \38198_38498 , \37850_38150 , \37856_38156 );
and \U$29824 ( \38199_38499 , \37850_38150 , \37863_38163 );
and \U$29825 ( \38200_38500 , \37856_38156 , \37863_38163 );
or \U$29826 ( \38201_38501 , \38198_38498 , \38199_38499 , \38200_38500 );
buf \U$29827 ( \38202_38502 , \38201_38501 );
and \U$29828 ( \38203_38503 , \16405_15940 , \34343_34643_nG9ba2 );
and \U$29829 ( \38204_38504 , \15638_15937 , \34794_35094_nG9b9f );
or \U$29830 ( \38205_38505 , \38203_38503 , \38204_38504 );
xor \U$29831 ( \38206_38506 , \15637_15936 , \38205_38505 );
buf \U$29832 ( \38207_38507 , \38206_38506 );
buf \U$29834 ( \38208_38508 , \38207_38507 );
xor \U$29835 ( \38209_38509 , \38202_38502 , \38208_38508 );
and \U$29836 ( \38210_38510 , \14710_14631 , \35270_35570_nG9b9c );
and \U$29837 ( \38211_38511 , \14329_14628 , \35501_35801_nG9b99 );
or \U$29838 ( \38212_38512 , \38210_38510 , \38211_38511 );
xor \U$29839 ( \38213_38513 , \14328_14627 , \38212_38512 );
buf \U$29840 ( \38214_38514 , \38213_38513 );
buf \U$29842 ( \38215_38515 , \38214_38514 );
xor \U$29843 ( \38216_38516 , \38209_38509 , \38215_38515 );
buf \U$29844 ( \38217_38517 , \38216_38516 );
xor \U$29845 ( \38218_38518 , \38197_38497 , \38217_38517 );
buf \U$29846 ( \38219_38519 , \38218_38518 );
xor \U$29847 ( \38220_38520 , \38186_38486 , \38219_38519 );
and \U$29848 ( \38221_38521 , \37784_38084 , \37790_38090 );
and \U$29849 ( \38222_38522 , \37784_38084 , \37797_38097 );
and \U$29850 ( \38223_38523 , \37790_38090 , \37797_38097 );
or \U$29851 ( \38224_38524 , \38221_38521 , \38222_38522 , \38223_38523 );
buf \U$29852 ( \38225_38525 , \38224_38524 );
and \U$29853 ( \38226_38526 , \38063_38363 , \38065_38365 );
and \U$29854 ( \38227_38527 , \38063_38363 , \38072_38372 );
and \U$29855 ( \38228_38528 , \38065_38365 , \38072_38372 );
or \U$29856 ( \38229_38529 , \38226_38526 , \38227_38527 , \38228_38528 );
buf \U$29857 ( \38230_38530 , \38229_38529 );
and \U$29858 ( \38231_38531 , \23495_23201 , \28300_28602_nG9bc0 );
and \U$29859 ( \38232_38532 , \22899_23198 , \28877_29179_nG9bbd );
or \U$29860 ( \38233_38533 , \38231_38531 , \38232_38532 );
xor \U$29861 ( \38234_38534 , \22898_23197 , \38233_38533 );
buf \U$29862 ( \38235_38535 , \38234_38534 );
buf \U$29864 ( \38236_38536 , \38235_38535 );
xor \U$29865 ( \38237_38537 , \38230_38530 , \38236_38536 );
and \U$29866 ( \38238_38538 , \21908_21658 , \30064_30366_nG9bba );
and \U$29867 ( \38239_38539 , \21356_21655 , \30638_30940_nG9bb7 );
or \U$29868 ( \38240_38540 , \38238_38538 , \38239_38539 );
xor \U$29869 ( \38241_38541 , \21355_21654 , \38240_38540 );
buf \U$29870 ( \38242_38542 , \38241_38541 );
buf \U$29872 ( \38243_38543 , \38242_38542 );
xor \U$29873 ( \38244_38544 , \38237_38537 , \38243_38543 );
buf \U$29874 ( \38245_38545 , \38244_38544 );
xor \U$29875 ( \38246_38546 , \38225_38525 , \38245_38545 );
and \U$29876 ( \38247_38547 , \12183_12157 , \36686_36986_nG9b90 );
and \U$29877 ( \38248_38548 , \11855_12154 , \36950_37250_nG9b8d );
or \U$29878 ( \38249_38549 , \38247_38547 , \38248_38548 );
xor \U$29879 ( \38250_38550 , \11854_12153 , \38249_38549 );
buf \U$29880 ( \38251_38551 , \38250_38550 );
buf \U$29882 ( \38252_38552 , \38251_38551 );
xor \U$29883 ( \38253_38553 , \38246_38546 , \38252_38552 );
buf \U$29884 ( \38254_38554 , \38253_38553 );
and \U$29885 ( \38255_38555 , \17437_17297 , \33741_34041_nG9ba8 );
and \U$29886 ( \38256_38556 , \16995_17294 , \33994_34294_nG9ba5 );
or \U$29887 ( \38257_38557 , \38255_38555 , \38256_38556 );
xor \U$29888 ( \38258_38558 , \16994_17293 , \38257_38557 );
buf \U$29889 ( \38259_38559 , \38258_38558 );
buf \U$29891 ( \38260_38560 , \38259_38559 );
and \U$29892 ( \38261_38561 , \13431_13370 , \35872_36172_nG9b96 );
and \U$29893 ( \38262_38562 , \13068_13367 , \36289_36589_nG9b93 );
or \U$29894 ( \38263_38563 , \38261_38561 , \38262_38562 );
xor \U$29895 ( \38264_38564 , \13067_13366 , \38263_38563 );
buf \U$29896 ( \38265_38565 , \38264_38564 );
buf \U$29898 ( \38266_38566 , \38265_38565 );
xor \U$29899 ( \38267_38567 , \38260_38560 , \38266_38566 );
and \U$29900 ( \38268_38568 , \10411_10707 , \38037_38337_nG9b84 );
and \U$29901 ( \38269_38569 , \37996_38296 , \38000_38300 );
and \U$29902 ( \38270_38570 , \38000_38300 , \38025_38325 );
and \U$29903 ( \38271_38571 , \37996_38296 , \38025_38325 );
or \U$29904 ( \38272_38572 , \38269_38569 , \38270_38570 , \38271_38571 );
and \U$29905 ( \38273_38573 , \37948_38248 , \37952_38252 );
and \U$29906 ( \38274_38574 , \37952_38252 , \37957_38257 );
and \U$29907 ( \38275_38575 , \37948_38248 , \37957_38257 );
or \U$29908 ( \38276_38576 , \38273_38573 , \38274_38574 , \38275_38575 );
and \U$29909 ( \38277_38577 , \37963_38263 , \37974_38274 );
and \U$29910 ( \38278_38578 , \37974_38274 , \37989_38289 );
and \U$29911 ( \38279_38579 , \37963_38263 , \37989_38289 );
or \U$29912 ( \38280_38580 , \38277_38577 , \38278_38578 , \38279_38579 );
xor \U$29913 ( \38281_38581 , \38276_38576 , \38280_38580 );
and \U$29914 ( \38282_38582 , \37967_38267 , \37971_38271 );
and \U$29915 ( \38283_38583 , \37971_38271 , \37973_38273 );
and \U$29916 ( \38284_38584 , \37967_38267 , \37973_38273 );
or \U$29917 ( \38285_38585 , \38282_38582 , \38283_38583 , \38284_38584 );
and \U$29918 ( \38286_38586 , \38014_38314 , \38018_38318 );
and \U$29919 ( \38287_38587 , \38018_38318 , \38023_38323 );
and \U$29920 ( \38288_38588 , \38014_38314 , \38023_38323 );
or \U$29921 ( \38289_38589 , \38286_38586 , \38287_38587 , \38288_38588 );
xor \U$29922 ( \38290_38590 , \38285_38585 , \38289_38589 );
and \U$29923 ( \38291_38591 , \29966_30268 , \22243_22542 );
and \U$29924 ( \38292_38592 , \30500_30802 , \21801_22103 );
nor \U$29925 ( \38293_38593 , \38291_38591 , \38292_38592 );
xnor \U$29926 ( \38294_38594 , \38293_38593 , \22249_22548 );
and \U$29927 ( \38295_38595 , \24970_25272 , \27095_27397 );
and \U$29928 ( \38296_38596 , \25516_25815 , \26505_26807 );
nor \U$29929 ( \38297_38597 , \38295_38595 , \38296_38596 );
xnor \U$29930 ( \38298_38598 , \38297_38597 , \26993_27295 );
xor \U$29931 ( \38299_38599 , \38294_38594 , \38298_38598 );
and \U$29932 ( \38300_38600 , \19259_19558 , \32503_32802 );
xor \U$29933 ( \38301_38601 , \38299_38599 , \38300_38600 );
xor \U$29934 ( \38302_38602 , \38290_38590 , \38301_38601 );
xor \U$29935 ( \38303_38603 , \38281_38581 , \38302_38602 );
xor \U$29936 ( \38304_38604 , \38272_38572 , \38303_38603 );
and \U$29937 ( \38305_38605 , \38005_38305 , \38009_38309 );
and \U$29938 ( \38306_38606 , \38009_38309 , \38024_38324 );
and \U$29939 ( \38307_38607 , \38005_38305 , \38024_38324 );
or \U$29940 ( \38308_38608 , \38305_38605 , \38306_38606 , \38307_38607 );
and \U$29941 ( \38309_38609 , \37944_38244 , \37958_38258 );
and \U$29942 ( \38310_38610 , \37958_38258 , \37990_38290 );
and \U$29943 ( \38311_38611 , \37944_38244 , \37990_38290 );
or \U$29944 ( \38312_38612 , \38309_38609 , \38310_38610 , \38311_38611 );
xor \U$29945 ( \38313_38613 , \38308_38608 , \38312_38612 );
not \U$29946 ( \38314_38614 , \19241_19540 );
and \U$29947 ( \38315_38615 , \31752_32054 , \20706_21005 );
and \U$29948 ( \38316_38616 , \32495_32794 , \20255_20557 );
nor \U$29949 ( \38317_38617 , \38315_38615 , \38316_38616 );
xnor \U$29950 ( \38318_38618 , \38317_38617 , \20712_21011 );
xor \U$29951 ( \38319_38619 , \38314_38614 , \38318_38618 );
and \U$29952 ( \38320_38620 , \28232_28534 , \23839_24138 );
and \U$29953 ( \38321_38621 , \28782_29084 , \23328_23630 );
nor \U$29954 ( \38322_38622 , \38320_38620 , \38321_38621 );
xnor \U$29955 ( \38323_38623 , \38322_38622 , \23845_24144 );
xor \U$29956 ( \38324_38624 , \38319_38619 , \38323_38623 );
and \U$29957 ( \38325_38625 , \26527_26829 , \25527_25826 );
and \U$29958 ( \38326_38626 , \27011_27313 , \24962_25264 );
nor \U$29959 ( \38327_38627 , \38325_38625 , \38326_38626 );
xnor \U$29960 ( \38328_38628 , \38327_38627 , \25474_25773 );
and \U$29961 ( \38329_38629 , \21788_22090 , \30521_30823 );
and \U$29962 ( \38330_38630 , \22257_22556 , \29944_30246 );
nor \U$29963 ( \38331_38631 , \38329_38629 , \38330_38630 );
xnor \U$29964 ( \38332_38632 , \38331_38631 , \30511_30813 );
xor \U$29965 ( \38333_38633 , \38328_38628 , \38332_38632 );
and \U$29966 ( \38334_38634 , \20242_20544 , \32555_32854 );
and \U$29967 ( \38335_38635 , \20734_21033 , \31765_32067 );
nor \U$29968 ( \38336_38636 , \38334_38634 , \38335_38635 );
xnor \U$29969 ( \38337_38637 , \38336_38636 , \32506_32805 );
xor \U$29970 ( \38338_38638 , \38333_38633 , \38337_38637 );
xor \U$29971 ( \38339_38639 , \38324_38624 , \38338_38638 );
and \U$29972 ( \38340_38640 , \37979_38279 , \37983_38283 );
and \U$29973 ( \38341_38641 , \37983_38283 , \37988_38288 );
and \U$29974 ( \38342_38642 , \37979_38279 , \37988_38288 );
or \U$29975 ( \38343_38643 , \38340_38640 , \38341_38641 , \38342_38642 );
buf \U$29976 ( \38344_38644 , \37956_38256 );
xor \U$29977 ( \38345_38645 , \38343_38643 , \38344_38644 );
and \U$29978 ( \38346_38646 , \23315_23617 , \28768_29070 );
and \U$29979 ( \38347_38647 , \23900_24199 , \28224_28526 );
nor \U$29980 ( \38348_38648 , \38346_38646 , \38347_38647 );
xnor \U$29981 ( \38349_38649 , \38348_38648 , \28774_29076 );
xor \U$29982 ( \38350_38650 , \38345_38645 , \38349_38649 );
xor \U$29983 ( \38351_38651 , \38339_38639 , \38350_38650 );
xor \U$29984 ( \38352_38652 , \38313_38613 , \38351_38651 );
xor \U$29985 ( \38353_38653 , \38304_38604 , \38352_38652 );
and \U$29986 ( \38354_38654 , \37940_38240 , \37991_38291 );
and \U$29987 ( \38355_38655 , \37991_38291 , \38026_38326 );
and \U$29988 ( \38356_38656 , \37940_38240 , \38026_38326 );
or \U$29989 ( \38357_38657 , \38354_38654 , \38355_38655 , \38356_38656 );
xor \U$29990 ( \38358_38658 , \38353_38653 , \38357_38657 );
and \U$29991 ( \38359_38659 , \38027_38327 , \38031_38331 );
and \U$29992 ( \38360_38660 , \38032_38332 , \38035_38335 );
or \U$29993 ( \38361_38661 , \38359_38659 , \38360_38660 );
xor \U$29994 ( \38362_38662 , \38358_38658 , \38361_38661 );
buf g9b81_GF_PartitionCandidate( \38363_38663_nG9b81 , \38362_38662 );
and \U$29995 ( \38364_38664 , \10402_10704 , \38363_38663_nG9b81 );
or \U$29996 ( \38365_38665 , \38268_38568 , \38364_38664 );
xor \U$29997 ( \38366_38666 , \10399_10703 , \38365_38665 );
buf \U$29998 ( \38367_38667 , \38366_38666 );
buf \U$30000 ( \38368_38668 , \38367_38667 );
xor \U$30001 ( \38369_38669 , \38267_38567 , \38368_38668 );
buf \U$30002 ( \38370_38670 , \38369_38669 );
xor \U$30003 ( \38371_38671 , \38254_38554 , \38370_38670 );
and \U$30004 ( \38372_38672 , \37899_38199 , \37905_38205 );
and \U$30005 ( \38373_38673 , \37899_38199 , \37912_38212 );
and \U$30006 ( \38374_38674 , \37905_38205 , \37912_38212 );
or \U$30007 ( \38375_38675 , \38372_38672 , \38373_38673 , \38374_38674 );
buf \U$30008 ( \38376_38676 , \38375_38675 );
and \U$30009 ( \38377_38677 , \28946_28118 , \23394_23696_nG9bd2 );
and \U$30010 ( \38378_38678 , \27816_28115 , \23927_24226_nG9bcf );
or \U$30011 ( \38379_38679 , \38377_38677 , \38378_38678 );
xor \U$30012 ( \38380_38680 , \27815_28114 , \38379_38679 );
buf \U$30013 ( \38381_38681 , \38380_38680 );
buf \U$30015 ( \38382_38682 , \38381_38681 );
and \U$30016 ( \38383_38683 , \27141_26431 , \24996_25298_nG9bcc );
and \U$30017 ( \38384_38684 , \26129_26428 , \25561_25860_nG9bc9 );
or \U$30018 ( \38385_38685 , \38383_38683 , \38384_38684 );
xor \U$30019 ( \38386_38686 , \26128_26427 , \38385_38685 );
buf \U$30020 ( \38387_38687 , \38386_38686 );
buf \U$30022 ( \38388_38688 , \38387_38687 );
xor \U$30023 ( \38389_38689 , \38382_38682 , \38388_38688 );
and \U$30024 ( \38390_38690 , \25044_24792 , \26585_26887_nG9bc6 );
and \U$30025 ( \38391_38691 , \24490_24789 , \27114_27416_nG9bc3 );
or \U$30026 ( \38392_38692 , \38390_38690 , \38391_38691 );
xor \U$30027 ( \38393_38693 , \24489_24788 , \38392_38692 );
buf \U$30028 ( \38394_38694 , \38393_38693 );
buf \U$30030 ( \38395_38695 , \38394_38694 );
xor \U$30031 ( \38396_38696 , \38389_38689 , \38395_38695 );
buf \U$30032 ( \38397_38697 , \38396_38696 );
xor \U$30033 ( \38398_38698 , \38376_38676 , \38397_38697 );
and \U$30034 ( \38399_38699 , \10996_10421 , \37307_37607_nG9b8a );
and \U$30035 ( \38400_38700 , \10119_10418 , \37674_37974_nG9b87 );
or \U$30036 ( \38401_38701 , \38399_38699 , \38400_38700 );
xor \U$30037 ( \38402_38702 , \10118_10417 , \38401_38701 );
buf \U$30038 ( \38403_38703 , \38402_38702 );
buf \U$30040 ( \38404_38704 , \38403_38703 );
xor \U$30041 ( \38405_38705 , \38398_38698 , \38404_38704 );
buf \U$30042 ( \38406_38706 , \38405_38705 );
xor \U$30043 ( \38407_38707 , \38371_38671 , \38406_38706 );
buf \U$30044 ( \38408_38708 , \38407_38707 );
xor \U$30045 ( \38409_38709 , \38220_38520 , \38408_38708 );
buf \U$30046 ( \38410_38710 , \38409_38709 );
xor \U$30047 ( \38411_38711 , \38181_38481 , \38410_38710 );
xor \U$30048 ( \38412_38712 , \38097_38397 , \38411_38711 );
and \U$30049 ( \38413_38713 , \37828_38128 , \37833_38133 );
and \U$30050 ( \38414_38714 , \37828_38128 , \38087_38387 );
and \U$30051 ( \38415_38715 , \37833_38133 , \38087_38387 );
or \U$30052 ( \38416_38716 , \38413_38713 , \38414_38714 , \38415_38715 );
and \U$30053 ( \38417_38717 , \38412_38712 , \38416_38716 );
and \U$30055 ( \38418_38718 , \38096_38396 , \38411_38711 );
or \U$30057 ( \38419_38719 , 1'b0 , \38418_38718 , 1'b0 );
xor \U$30058 ( \38420_38720 , \38417_38717 , \38419_38719 );
and \U$30060 ( \38421_38721 , \38089_38389 , \38095_38395 );
and \U$30061 ( \38422_38722 , \38091_38391 , \38095_38395 );
or \U$30062 ( \38423_38723 , 1'b0 , \38421_38721 , \38422_38722 );
xor \U$30063 ( \38424_38724 , \38420_38720 , \38423_38723 );
xor \U$30070 ( \38425_38725 , \38424_38724 , 1'b0 );
and \U$30071 ( \38426_38726 , \38175_38475 , \38180_38480 );
and \U$30072 ( \38427_38727 , \38175_38475 , \38410_38710 );
and \U$30073 ( \38428_38728 , \38180_38480 , \38410_38710 );
or \U$30074 ( \38429_38729 , \38426_38726 , \38427_38727 , \38428_38728 );
xor \U$30075 ( \38430_38730 , \38425_38725 , \38429_38729 );
and \U$30076 ( \38431_38731 , \38186_38486 , \38219_38519 );
and \U$30077 ( \38432_38732 , \38186_38486 , \38408_38708 );
and \U$30078 ( \38433_38733 , \38219_38519 , \38408_38708 );
or \U$30079 ( \38434_38734 , \38431_38731 , \38432_38732 , \38433_38733 );
buf \U$30080 ( \38435_38735 , \38434_38734 );
and \U$30081 ( \38436_38736 , \38191_38491 , \38196_38496 );
and \U$30082 ( \38437_38737 , \38191_38491 , \38217_38517 );
and \U$30083 ( \38438_38738 , \38196_38496 , \38217_38517 );
or \U$30084 ( \38439_38739 , \38436_38736 , \38437_38737 , \38438_38738 );
buf \U$30085 ( \38440_38740 , \38439_38739 );
and \U$30086 ( \38441_38741 , \38382_38682 , \38388_38688 );
and \U$30087 ( \38442_38742 , \38382_38682 , \38395_38695 );
and \U$30088 ( \38443_38743 , \38388_38688 , \38395_38695 );
or \U$30089 ( \38444_38744 , \38441_38741 , \38442_38742 , \38443_38743 );
buf \U$30090 ( \38445_38745 , \38444_38744 );
and \U$30091 ( \38446_38746 , \16405_15940 , \34794_35094_nG9b9f );
and \U$30092 ( \38447_38747 , \15638_15937 , \35270_35570_nG9b9c );
or \U$30093 ( \38448_38748 , \38446_38746 , \38447_38747 );
xor \U$30094 ( \38449_38749 , \15637_15936 , \38448_38748 );
buf \U$30095 ( \38450_38750 , \38449_38749 );
buf \U$30097 ( \38451_38751 , \38450_38750 );
xor \U$30098 ( \38452_38752 , \38445_38745 , \38451_38751 );
and \U$30099 ( \38453_38753 , \14710_14631 , \35501_35801_nG9b99 );
and \U$30100 ( \38454_38754 , \14329_14628 , \35872_36172_nG9b96 );
or \U$30101 ( \38455_38755 , \38453_38753 , \38454_38754 );
xor \U$30102 ( \38456_38756 , \14328_14627 , \38455_38755 );
buf \U$30103 ( \38457_38757 , \38456_38756 );
buf \U$30105 ( \38458_38758 , \38457_38757 );
xor \U$30106 ( \38459_38759 , \38452_38752 , \38458_38758 );
buf \U$30107 ( \38460_38760 , \38459_38759 );
and \U$30109 ( \38461_38761 , \32617_32916 , \20306_20608_nG9bde );
or \U$30110 ( \38462_38762 , 1'b0 , \38461_38761 );
xor \U$30111 ( \38463_38763 , 1'b0 , \38462_38762 );
buf \U$30112 ( \38464_38764 , \38463_38763 );
buf \U$30114 ( \38465_38765 , \38464_38764 );
and \U$30115 ( \38466_38766 , \31989_31636 , \20787_21086_nG9bdb );
and \U$30116 ( \38467_38767 , \31334_31633 , \21827_22129_nG9bd8 );
or \U$30117 ( \38468_38768 , \38466_38766 , \38467_38767 );
xor \U$30118 ( \38469_38769 , \31333_31632 , \38468_38768 );
buf \U$30119 ( \38470_38770 , \38469_38769 );
buf \U$30121 ( \38471_38771 , \38470_38770 );
xor \U$30122 ( \38472_38772 , \38465_38765 , \38471_38771 );
buf \U$30123 ( \38473_38773 , \38472_38772 );
and \U$30124 ( \38474_38774 , \38113_38413 , \38119_38419 );
buf \U$30125 ( \38475_38775 , \38474_38774 );
xor \U$30126 ( \38476_38776 , \38473_38773 , \38475_38775 );
and \U$30127 ( \38477_38777 , \30670_29853 , \22330_22629_nG9bd5 );
and \U$30128 ( \38478_38778 , \29551_29850 , \23394_23696_nG9bd2 );
or \U$30129 ( \38479_38779 , \38477_38777 , \38478_38778 );
xor \U$30130 ( \38480_38780 , \29550_29849 , \38479_38779 );
buf \U$30131 ( \38481_38781 , \38480_38780 );
buf \U$30133 ( \38482_38782 , \38481_38781 );
xor \U$30134 ( \38483_38783 , \38476_38776 , \38482_38782 );
buf \U$30135 ( \38484_38784 , \38483_38783 );
and \U$30136 ( \38485_38785 , \20353_20155 , \32589_32888_nG9bb1 );
and \U$30137 ( \38486_38786 , \19853_20152 , \32881_33181_nG9bae );
or \U$30138 ( \38487_38787 , \38485_38785 , \38486_38786 );
xor \U$30139 ( \38488_38788 , \19852_20151 , \38487_38787 );
buf \U$30140 ( \38489_38789 , \38488_38788 );
buf \U$30142 ( \38490_38790 , \38489_38789 );
xor \U$30143 ( \38491_38791 , \38484_38784 , \38490_38790 );
and \U$30144 ( \38492_38792 , \18908_18702 , \33313_33613_nG9bab );
and \U$30145 ( \38493_38793 , \18400_18699 , \33741_34041_nG9ba8 );
or \U$30146 ( \38494_38794 , \38492_38792 , \38493_38793 );
xor \U$30147 ( \38495_38795 , \18399_18698 , \38494_38794 );
buf \U$30148 ( \38496_38796 , \38495_38795 );
buf \U$30150 ( \38497_38797 , \38496_38796 );
xor \U$30151 ( \38498_38798 , \38491_38791 , \38497_38797 );
buf \U$30152 ( \38499_38799 , \38498_38798 );
xor \U$30153 ( \38500_38800 , \38460_38760 , \38499_38799 );
and \U$30154 ( \38501_38801 , \38202_38502 , \38208_38508 );
and \U$30155 ( \38502_38802 , \38202_38502 , \38215_38515 );
and \U$30156 ( \38503_38803 , \38208_38508 , \38215_38515 );
or \U$30157 ( \38504_38804 , \38501_38801 , \38502_38802 , \38503_38803 );
buf \U$30158 ( \38505_38805 , \38504_38804 );
xor \U$30159 ( \38506_38806 , \38500_38800 , \38505_38805 );
buf \U$30160 ( \38507_38807 , \38506_38806 );
xor \U$30161 ( \38508_38808 , \38440_38740 , \38507_38807 );
and \U$30162 ( \38509_38809 , \38102_38402 , \38107_38407 );
and \U$30163 ( \38510_38810 , \38102_38402 , \38147_38447 );
and \U$30164 ( \38511_38811 , \38107_38407 , \38147_38447 );
or \U$30165 ( \38512_38812 , \38509_38809 , \38510_38810 , \38511_38811 );
buf \U$30166 ( \38513_38813 , \38512_38812 );
xor \U$30167 ( \38514_38814 , \38508_38808 , \38513_38813 );
buf \U$30168 ( \38515_38815 , \38514_38814 );
xor \U$30169 ( \38516_38816 , \38435_38735 , \38515_38815 );
and \U$30170 ( \38517_38817 , \38149_38449 , \38154_38454 );
and \U$30171 ( \38518_38818 , \38149_38449 , \38160_38460 );
and \U$30172 ( \38519_38819 , \38154_38454 , \38160_38460 );
or \U$30173 ( \38520_38820 , \38517_38817 , \38518_38818 , \38519_38819 );
buf \U$30174 ( \38521_38821 , \38520_38820 );
xor \U$30175 ( \38522_38822 , \38516_38816 , \38521_38821 );
buf \U$30176 ( \38523_38823 , \38522_38822 );
and \U$30177 ( \38524_38824 , \38162_38462 , \38167_38467 );
and \U$30178 ( \38525_38825 , \38162_38462 , \38173_38473 );
and \U$30179 ( \38526_38826 , \38167_38467 , \38173_38473 );
or \U$30180 ( \38527_38827 , \38524_38824 , \38525_38825 , \38526_38826 );
buf \U$30181 ( \38528_38828 , \38527_38827 );
xor \U$30182 ( \38529_38829 , \38523_38823 , \38528_38828 );
and \U$30183 ( \38530_38830 , \38132_38432 , \38138_38438 );
and \U$30184 ( \38531_38831 , \38132_38432 , \38145_38445 );
and \U$30185 ( \38532_38832 , \38138_38438 , \38145_38445 );
or \U$30186 ( \38533_38833 , \38530_38830 , \38531_38831 , \38532_38832 );
buf \U$30187 ( \38534_38834 , \38533_38833 );
and \U$30188 ( \38535_38835 , \38121_38421 , \38123_38423 );
and \U$30189 ( \38536_38836 , \38121_38421 , \38130_38430 );
and \U$30190 ( \38537_38837 , \38123_38423 , \38130_38430 );
or \U$30191 ( \38538_38838 , \38535_38835 , \38536_38836 , \38537_38837 );
buf \U$30192 ( \38539_38839 , \38538_38838 );
and \U$30193 ( \38540_38840 , \23495_23201 , \28877_29179_nG9bbd );
and \U$30194 ( \38541_38841 , \22899_23198 , \30064_30366_nG9bba );
or \U$30195 ( \38542_38842 , \38540_38840 , \38541_38841 );
xor \U$30196 ( \38543_38843 , \22898_23197 , \38542_38842 );
buf \U$30197 ( \38544_38844 , \38543_38843 );
buf \U$30199 ( \38545_38845 , \38544_38844 );
xor \U$30200 ( \38546_38846 , \38539_38839 , \38545_38845 );
and \U$30201 ( \38547_38847 , \21908_21658 , \30638_30940_nG9bb7 );
and \U$30202 ( \38548_38848 , \21356_21655 , \31877_32179_nG9bb4 );
or \U$30203 ( \38549_38849 , \38547_38847 , \38548_38848 );
xor \U$30204 ( \38550_38850 , \21355_21654 , \38549_38849 );
buf \U$30205 ( \38551_38851 , \38550_38850 );
buf \U$30207 ( \38552_38852 , \38551_38851 );
xor \U$30208 ( \38553_38853 , \38546_38846 , \38552_38852 );
buf \U$30209 ( \38554_38854 , \38553_38853 );
xor \U$30210 ( \38555_38855 , \38534_38834 , \38554_38854 );
and \U$30211 ( \38556_38856 , \12183_12157 , \36950_37250_nG9b8d );
and \U$30212 ( \38557_38857 , \11855_12154 , \37307_37607_nG9b8a );
or \U$30213 ( \38558_38858 , \38556_38856 , \38557_38857 );
xor \U$30214 ( \38559_38859 , \11854_12153 , \38558_38858 );
buf \U$30215 ( \38560_38860 , \38559_38859 );
buf \U$30217 ( \38561_38861 , \38560_38860 );
xor \U$30218 ( \38562_38862 , \38555_38855 , \38561_38861 );
buf \U$30219 ( \38563_38863 , \38562_38862 );
and \U$30220 ( \38564_38864 , \17437_17297 , \33994_34294_nG9ba5 );
and \U$30221 ( \38565_38865 , \16995_17294 , \34343_34643_nG9ba2 );
or \U$30222 ( \38566_38866 , \38564_38864 , \38565_38865 );
xor \U$30223 ( \38567_38867 , \16994_17293 , \38566_38866 );
buf \U$30224 ( \38568_38868 , \38567_38867 );
buf \U$30226 ( \38569_38869 , \38568_38868 );
and \U$30227 ( \38570_38870 , \13431_13370 , \36289_36589_nG9b93 );
and \U$30228 ( \38571_38871 , \13068_13367 , \36686_36986_nG9b90 );
or \U$30229 ( \38572_38872 , \38570_38870 , \38571_38871 );
xor \U$30230 ( \38573_38873 , \13067_13366 , \38572_38872 );
buf \U$30231 ( \38574_38874 , \38573_38873 );
buf \U$30233 ( \38575_38875 , \38574_38874 );
xor \U$30234 ( \38576_38876 , \38569_38869 , \38575_38875 );
and \U$30235 ( \38577_38877 , \10411_10707 , \38363_38663_nG9b81 );
and \U$30236 ( \38578_38878 , \38308_38608 , \38312_38612 );
and \U$30237 ( \38579_38879 , \38312_38612 , \38351_38651 );
and \U$30238 ( \38580_38880 , \38308_38608 , \38351_38651 );
or \U$30239 ( \38581_38881 , \38578_38878 , \38579_38879 , \38580_38880 );
and \U$30240 ( \38582_38882 , \38343_38643 , \38344_38644 );
and \U$30241 ( \38583_38883 , \38344_38644 , \38349_38649 );
and \U$30242 ( \38584_38884 , \38343_38643 , \38349_38649 );
or \U$30243 ( \38585_38885 , \38582_38882 , \38583_38883 , \38584_38884 );
and \U$30244 ( \38586_38886 , \38285_38585 , \38289_38589 );
and \U$30245 ( \38587_38887 , \38289_38589 , \38301_38601 );
and \U$30246 ( \38588_38888 , \38285_38585 , \38301_38601 );
or \U$30247 ( \38589_38889 , \38586_38886 , \38587_38887 , \38588_38888 );
xor \U$30248 ( \38590_38890 , \38585_38885 , \38589_38889 );
and \U$30249 ( \38591_38891 , \38294_38594 , \38298_38598 );
and \U$30250 ( \38592_38892 , \38298_38598 , \38300_38600 );
and \U$30251 ( \38593_38893 , \38294_38594 , \38300_38600 );
or \U$30252 ( \38594_38894 , \38591_38891 , \38592_38892 , \38593_38893 );
and \U$30253 ( \38595_38895 , \38314_38614 , \38318_38618 );
and \U$30254 ( \38596_38896 , \38318_38618 , \38323_38623 );
and \U$30255 ( \38597_38897 , \38314_38614 , \38323_38623 );
or \U$30256 ( \38598_38898 , \38595_38895 , \38596_38896 , \38597_38897 );
xor \U$30257 ( \38599_38899 , \38594_38894 , \38598_38898 );
and \U$30258 ( \38600_38900 , \38328_38628 , \38332_38632 );
and \U$30259 ( \38601_38901 , \38332_38632 , \38337_38637 );
and \U$30260 ( \38602_38902 , \38328_38628 , \38337_38637 );
or \U$30261 ( \38603_38903 , \38600_38900 , \38601_38901 , \38602_38902 );
xor \U$30262 ( \38604_38904 , \38599_38899 , \38603_38903 );
xor \U$30263 ( \38605_38905 , \38590_38890 , \38604_38904 );
xor \U$30264 ( \38606_38906 , \38581_38881 , \38605_38905 );
and \U$30265 ( \38607_38907 , \38324_38624 , \38338_38638 );
and \U$30266 ( \38608_38908 , \38338_38638 , \38350_38650 );
and \U$30267 ( \38609_38909 , \38324_38624 , \38350_38650 );
or \U$30268 ( \38610_38910 , \38607_38907 , \38608_38908 , \38609_38909 );
and \U$30269 ( \38611_38911 , \38276_38576 , \38280_38580 );
and \U$30270 ( \38612_38912 , \38280_38580 , \38302_38602 );
and \U$30271 ( \38613_38913 , \38276_38576 , \38302_38602 );
or \U$30272 ( \38614_38914 , \38611_38911 , \38612_38912 , \38613_38913 );
xor \U$30273 ( \38615_38915 , \38610_38910 , \38614_38914 );
and \U$30274 ( \38616_38916 , \30500_30802 , \22243_22542 );
and \U$30275 ( \38617_38917 , \31752_32054 , \21801_22103 );
nor \U$30276 ( \38618_38918 , \38616_38916 , \38617_38917 );
xnor \U$30277 ( \38619_38919 , \38618_38918 , \22249_22548 );
and \U$30278 ( \38620_38920 , \28782_29084 , \23839_24138 );
and \U$30279 ( \38621_38921 , \29966_30268 , \23328_23630 );
nor \U$30280 ( \38622_38922 , \38620_38920 , \38621_38921 );
xnor \U$30281 ( \38623_38923 , \38622_38922 , \23845_24144 );
xor \U$30282 ( \38624_38924 , \38619_38919 , \38623_38923 );
and \U$30283 ( \38625_38925 , \25516_25815 , \27095_27397 );
and \U$30284 ( \38626_38926 , \26527_26829 , \26505_26807 );
nor \U$30285 ( \38627_38927 , \38625_38925 , \38626_38926 );
xnor \U$30286 ( \38628_38928 , \38627_38927 , \26993_27295 );
xor \U$30287 ( \38629_38929 , \38624_38924 , \38628_38928 );
and \U$30288 ( \38630_38930 , \27011_27313 , \25527_25826 );
and \U$30289 ( \38631_38931 , \28232_28534 , \24962_25264 );
nor \U$30290 ( \38632_38932 , \38630_38930 , \38631_38931 );
xnor \U$30291 ( \38633_38933 , \38632_38932 , \25474_25773 );
and \U$30292 ( \38634_38934 , \20734_21033 , \32555_32854 );
and \U$30293 ( \38635_38935 , \21788_22090 , \31765_32067 );
nor \U$30294 ( \38636_38936 , \38634_38934 , \38635_38935 );
xnor \U$30295 ( \38637_38937 , \38636_38936 , \32506_32805 );
xor \U$30296 ( \38638_38938 , \38633_38933 , \38637_38937 );
and \U$30297 ( \38639_38939 , \20242_20544 , \32503_32802 );
xor \U$30298 ( \38640_38940 , \38638_38938 , \38639_38939 );
xor \U$30299 ( \38641_38941 , \38629_38929 , \38640_38940 );
and \U$30300 ( \38642_38942 , \32495_32794 , \20706_21005 );
not \U$30301 ( \38643_38943 , \38642_38942 );
xnor \U$30302 ( \38644_38944 , \38643_38943 , \20712_21011 );
not \U$30303 ( \38645_38945 , \38644_38944 );
and \U$30304 ( \38646_38946 , \23900_24199 , \28768_29070 );
and \U$30305 ( \38647_38947 , \24970_25272 , \28224_28526 );
nor \U$30306 ( \38648_38948 , \38646_38946 , \38647_38947 );
xnor \U$30307 ( \38649_38949 , \38648_38948 , \28774_29076 );
xor \U$30308 ( \38650_38950 , \38645_38945 , \38649_38949 );
and \U$30309 ( \38651_38951 , \22257_22556 , \30521_30823 );
and \U$30310 ( \38652_38952 , \23315_23617 , \29944_30246 );
nor \U$30311 ( \38653_38953 , \38651_38951 , \38652_38952 );
xnor \U$30312 ( \38654_38954 , \38653_38953 , \30511_30813 );
xor \U$30313 ( \38655_38955 , \38650_38950 , \38654_38954 );
xor \U$30314 ( \38656_38956 , \38641_38941 , \38655_38955 );
xor \U$30315 ( \38657_38957 , \38615_38915 , \38656_38956 );
xor \U$30316 ( \38658_38958 , \38606_38906 , \38657_38957 );
and \U$30317 ( \38659_38959 , \38272_38572 , \38303_38603 );
and \U$30318 ( \38660_38960 , \38303_38603 , \38352_38652 );
and \U$30319 ( \38661_38961 , \38272_38572 , \38352_38652 );
or \U$30320 ( \38662_38962 , \38659_38959 , \38660_38960 , \38661_38961 );
xor \U$30321 ( \38663_38963 , \38658_38958 , \38662_38962 );
and \U$30322 ( \38664_38964 , \38353_38653 , \38357_38657 );
and \U$30323 ( \38665_38965 , \38358_38658 , \38361_38661 );
or \U$30324 ( \38666_38966 , \38664_38964 , \38665_38965 );
xor \U$30325 ( \38667_38967 , \38663_38963 , \38666_38966 );
buf g9b7e_GF_PartitionCandidate( \38668_38968_nG9b7e , \38667_38967 );
and \U$30326 ( \38669_38969 , \10402_10704 , \38668_38968_nG9b7e );
or \U$30327 ( \38670_38970 , \38577_38877 , \38669_38969 );
xor \U$30328 ( \38671_38971 , \10399_10703 , \38670_38970 );
buf \U$30329 ( \38672_38972 , \38671_38971 );
buf \U$30331 ( \38673_38973 , \38672_38972 );
xor \U$30332 ( \38674_38974 , \38576_38876 , \38673_38973 );
buf \U$30333 ( \38675_38975 , \38674_38974 );
xor \U$30334 ( \38676_38976 , \38563_38863 , \38675_38975 );
and \U$30335 ( \38677_38977 , \38230_38530 , \38236_38536 );
and \U$30336 ( \38678_38978 , \38230_38530 , \38243_38543 );
and \U$30337 ( \38679_38979 , \38236_38536 , \38243_38543 );
or \U$30338 ( \38680_38980 , \38677_38977 , \38678_38978 , \38679_38979 );
buf \U$30339 ( \38681_38981 , \38680_38980 );
and \U$30340 ( \38682_38982 , \28946_28118 , \23927_24226_nG9bcf );
and \U$30341 ( \38683_38983 , \27816_28115 , \24996_25298_nG9bcc );
or \U$30342 ( \38684_38984 , \38682_38982 , \38683_38983 );
xor \U$30343 ( \38685_38985 , \27815_28114 , \38684_38984 );
buf \U$30344 ( \38686_38986 , \38685_38985 );
buf \U$30346 ( \38687_38987 , \38686_38986 );
and \U$30347 ( \38688_38988 , \27141_26431 , \25561_25860_nG9bc9 );
and \U$30348 ( \38689_38989 , \26129_26428 , \26585_26887_nG9bc6 );
or \U$30349 ( \38690_38990 , \38688_38988 , \38689_38989 );
xor \U$30350 ( \38691_38991 , \26128_26427 , \38690_38990 );
buf \U$30351 ( \38692_38992 , \38691_38991 );
buf \U$30353 ( \38693_38993 , \38692_38992 );
xor \U$30354 ( \38694_38994 , \38687_38987 , \38693_38993 );
and \U$30355 ( \38695_38995 , \25044_24792 , \27114_27416_nG9bc3 );
and \U$30356 ( \38696_38996 , \24490_24789 , \28300_28602_nG9bc0 );
or \U$30357 ( \38697_38997 , \38695_38995 , \38696_38996 );
xor \U$30358 ( \38698_38998 , \24489_24788 , \38697_38997 );
buf \U$30359 ( \38699_38999 , \38698_38998 );
buf \U$30361 ( \38700_39000 , \38699_38999 );
xor \U$30362 ( \38701_39001 , \38694_38994 , \38700_39000 );
buf \U$30363 ( \38702_39002 , \38701_39001 );
xor \U$30364 ( \38703_39003 , \38681_38981 , \38702_39002 );
and \U$30365 ( \38704_39004 , \10996_10421 , \37674_37974_nG9b87 );
and \U$30366 ( \38705_39005 , \10119_10418 , \38037_38337_nG9b84 );
or \U$30367 ( \38706_39006 , \38704_39004 , \38705_39005 );
xor \U$30368 ( \38707_39007 , \10118_10417 , \38706_39006 );
buf \U$30369 ( \38708_39008 , \38707_39007 );
buf \U$30371 ( \38709_39009 , \38708_39008 );
xor \U$30372 ( \38710_39010 , \38703_39003 , \38709_39009 );
buf \U$30373 ( \38711_39011 , \38710_39010 );
xor \U$30374 ( \38712_39012 , \38676_38976 , \38711_39011 );
buf \U$30375 ( \38713_39013 , \38712_39012 );
and \U$30376 ( \38714_39014 , \38225_38525 , \38245_38545 );
and \U$30377 ( \38715_39015 , \38225_38525 , \38252_38552 );
and \U$30378 ( \38716_39016 , \38245_38545 , \38252_38552 );
or \U$30379 ( \38717_39017 , \38714_39014 , \38715_39015 , \38716_39016 );
buf \U$30380 ( \38718_39018 , \38717_39017 );
and \U$30381 ( \38719_39019 , \38260_38560 , \38266_38566 );
and \U$30382 ( \38720_39020 , \38260_38560 , \38368_38668 );
and \U$30383 ( \38721_39021 , \38266_38566 , \38368_38668 );
or \U$30384 ( \38722_39022 , \38719_39019 , \38720_39020 , \38721_39021 );
buf \U$30385 ( \38723_39023 , \38722_39022 );
xor \U$30386 ( \38724_39024 , \38718_39018 , \38723_39023 );
and \U$30387 ( \38725_39025 , \38376_38676 , \38397_38697 );
and \U$30388 ( \38726_39026 , \38376_38676 , \38404_38704 );
and \U$30389 ( \38727_39027 , \38397_38697 , \38404_38704 );
or \U$30390 ( \38728_39028 , \38725_39025 , \38726_39026 , \38727_39027 );
buf \U$30391 ( \38729_39029 , \38728_39028 );
xor \U$30392 ( \38730_39030 , \38724_39024 , \38729_39029 );
buf \U$30393 ( \38731_39031 , \38730_39030 );
xor \U$30394 ( \38732_39032 , \38713_39013 , \38731_39031 );
and \U$30395 ( \38733_39033 , \38254_38554 , \38370_38670 );
and \U$30396 ( \38734_39034 , \38254_38554 , \38406_38706 );
and \U$30397 ( \38735_39035 , \38370_38670 , \38406_38706 );
or \U$30398 ( \38736_39036 , \38733_39033 , \38734_39034 , \38735_39035 );
buf \U$30399 ( \38737_39037 , \38736_39036 );
xor \U$30400 ( \38738_39038 , \38732_39032 , \38737_39037 );
buf \U$30401 ( \38739_39039 , \38738_39038 );
xor \U$30402 ( \38740_39040 , \38529_38829 , \38739_39039 );
and \U$30403 ( \38741_39041 , \38430_38730 , \38740_39040 );
and \U$30405 ( \38742_39042 , \38424_38724 , \38429_38729 );
or \U$30407 ( \38743_39043 , 1'b0 , \38742_39042 , 1'b0 );
xor \U$30408 ( \38744_39044 , \38741_39041 , \38743_39043 );
and \U$30410 ( \38745_39045 , \38417_38717 , \38423_38723 );
and \U$30411 ( \38746_39046 , \38419_38719 , \38423_38723 );
or \U$30412 ( \38747_39047 , 1'b0 , \38745_39045 , \38746_39046 );
xor \U$30413 ( \38748_39048 , \38744_39044 , \38747_39047 );
xor \U$30420 ( \38749_39049 , \38748_39048 , 1'b0 );
and \U$30421 ( \38750_39050 , \38523_38823 , \38528_38828 );
and \U$30422 ( \38751_39051 , \38523_38823 , \38739_39039 );
and \U$30423 ( \38752_39052 , \38528_38828 , \38739_39039 );
or \U$30424 ( \38753_39053 , \38750_39050 , \38751_39051 , \38752_39052 );
xor \U$30425 ( \38754_39054 , \38749_39049 , \38753_39053 );
and \U$30426 ( \38755_39055 , \38460_38760 , \38499_38799 );
and \U$30427 ( \38756_39056 , \38460_38760 , \38505_38805 );
and \U$30428 ( \38757_39057 , \38499_38799 , \38505_38805 );
or \U$30429 ( \38758_39058 , \38755_39055 , \38756_39056 , \38757_39057 );
buf \U$30430 ( \38759_39059 , \38758_39058 );
and \U$30431 ( \38760_39060 , \38539_38839 , \38545_38845 );
and \U$30432 ( \38761_39061 , \38539_38839 , \38552_38852 );
and \U$30433 ( \38762_39062 , \38545_38845 , \38552_38852 );
or \U$30434 ( \38763_39063 , \38760_39060 , \38761_39061 , \38762_39062 );
buf \U$30435 ( \38764_39064 , \38763_39063 );
and \U$30436 ( \38765_39065 , \38473_38773 , \38475_38775 );
and \U$30437 ( \38766_39066 , \38473_38773 , \38482_38782 );
and \U$30438 ( \38767_39067 , \38475_38775 , \38482_38782 );
or \U$30439 ( \38768_39068 , \38765_39065 , \38766_39066 , \38767_39067 );
buf \U$30440 ( \38769_39069 , \38768_39068 );
and \U$30441 ( \38770_39070 , \28946_28118 , \24996_25298_nG9bcc );
and \U$30442 ( \38771_39071 , \27816_28115 , \25561_25860_nG9bc9 );
or \U$30443 ( \38772_39072 , \38770_39070 , \38771_39071 );
xor \U$30444 ( \38773_39073 , \27815_28114 , \38772_39072 );
buf \U$30445 ( \38774_39074 , \38773_39073 );
buf \U$30447 ( \38775_39075 , \38774_39074 );
xor \U$30448 ( \38776_39076 , \38769_39069 , \38775_39075 );
and \U$30449 ( \38777_39077 , \27141_26431 , \26585_26887_nG9bc6 );
and \U$30450 ( \38778_39078 , \26129_26428 , \27114_27416_nG9bc3 );
or \U$30451 ( \38779_39079 , \38777_39077 , \38778_39078 );
xor \U$30452 ( \38780_39080 , \26128_26427 , \38779_39079 );
buf \U$30453 ( \38781_39081 , \38780_39080 );
buf \U$30455 ( \38782_39082 , \38781_39081 );
xor \U$30456 ( \38783_39083 , \38776_39076 , \38782_39082 );
buf \U$30457 ( \38784_39084 , \38783_39083 );
xor \U$30458 ( \38785_39085 , \38764_39064 , \38784_39084 );
and \U$30459 ( \38786_39086 , \12183_12157 , \37307_37607_nG9b8a );
and \U$30460 ( \38787_39087 , \11855_12154 , \37674_37974_nG9b87 );
or \U$30461 ( \38788_39088 , \38786_39086 , \38787_39087 );
xor \U$30462 ( \38789_39089 , \11854_12153 , \38788_39088 );
buf \U$30463 ( \38790_39090 , \38789_39089 );
buf \U$30465 ( \38791_39091 , \38790_39090 );
xor \U$30466 ( \38792_39092 , \38785_39085 , \38791_39091 );
buf \U$30467 ( \38793_39093 , \38792_39092 );
and \U$30468 ( \38794_39094 , \38681_38981 , \38702_39002 );
and \U$30469 ( \38795_39095 , \38681_38981 , \38709_39009 );
and \U$30470 ( \38796_39096 , \38702_39002 , \38709_39009 );
or \U$30471 ( \38797_39097 , \38794_39094 , \38795_39095 , \38796_39096 );
buf \U$30472 ( \38798_39098 , \38797_39097 );
xor \U$30473 ( \38799_39099 , \38793_39093 , \38798_39098 );
and \U$30474 ( \38800_39100 , \38687_38987 , \38693_38993 );
and \U$30475 ( \38801_39101 , \38687_38987 , \38700_39000 );
and \U$30476 ( \38802_39102 , \38693_38993 , \38700_39000 );
or \U$30477 ( \38803_39103 , \38800_39100 , \38801_39101 , \38802_39102 );
buf \U$30478 ( \38804_39104 , \38803_39103 );
and \U$30479 ( \38805_39105 , \21908_21658 , \31877_32179_nG9bb4 );
and \U$30480 ( \38806_39106 , \21356_21655 , \32589_32888_nG9bb1 );
or \U$30481 ( \38807_39107 , \38805_39105 , \38806_39106 );
xor \U$30482 ( \38808_39108 , \21355_21654 , \38807_39107 );
buf \U$30483 ( \38809_39109 , \38808_39108 );
buf \U$30485 ( \38810_39110 , \38809_39109 );
xor \U$30486 ( \38811_39111 , \38804_39104 , \38810_39110 );
and \U$30487 ( \38812_39112 , \18908_18702 , \33741_34041_nG9ba8 );
and \U$30488 ( \38813_39113 , \18400_18699 , \33994_34294_nG9ba5 );
or \U$30489 ( \38814_39114 , \38812_39112 , \38813_39113 );
xor \U$30490 ( \38815_39115 , \18399_18698 , \38814_39114 );
buf \U$30491 ( \38816_39116 , \38815_39115 );
buf \U$30493 ( \38817_39117 , \38816_39116 );
xor \U$30494 ( \38818_39118 , \38811_39111 , \38817_39117 );
buf \U$30495 ( \38819_39119 , \38818_39118 );
xor \U$30496 ( \38820_39120 , \38799_39099 , \38819_39119 );
buf \U$30497 ( \38821_39121 , \38820_39120 );
xor \U$30498 ( \38822_39122 , \38759_39059 , \38821_39121 );
and \U$30500 ( \38823_39123 , \32617_32916 , \20787_21086_nG9bdb );
or \U$30501 ( \38824_39124 , 1'b0 , \38823_39123 );
xor \U$30502 ( \38825_39125 , 1'b0 , \38824_39124 );
buf \U$30503 ( \38826_39126 , \38825_39125 );
buf \U$30505 ( \38827_39127 , \38826_39126 );
and \U$30506 ( \38828_39128 , \31989_31636 , \21827_22129_nG9bd8 );
and \U$30507 ( \38829_39129 , \31334_31633 , \22330_22629_nG9bd5 );
or \U$30508 ( \38830_39130 , \38828_39128 , \38829_39129 );
xor \U$30509 ( \38831_39131 , \31333_31632 , \38830_39130 );
buf \U$30510 ( \38832_39132 , \38831_39131 );
buf \U$30512 ( \38833_39133 , \38832_39132 );
xor \U$30513 ( \38834_39134 , \38827_39127 , \38833_39133 );
buf \U$30514 ( \38835_39135 , \38834_39134 );
and \U$30515 ( \38836_39136 , \38465_38765 , \38471_38771 );
buf \U$30516 ( \38837_39137 , \38836_39136 );
xor \U$30517 ( \38838_39138 , \38835_39135 , \38837_39137 );
and \U$30518 ( \38839_39139 , \30670_29853 , \23394_23696_nG9bd2 );
and \U$30519 ( \38840_39140 , \29551_29850 , \23927_24226_nG9bcf );
or \U$30520 ( \38841_39141 , \38839_39139 , \38840_39140 );
xor \U$30521 ( \38842_39142 , \29550_29849 , \38841_39141 );
buf \U$30522 ( \38843_39143 , \38842_39142 );
buf \U$30524 ( \38844_39144 , \38843_39143 );
xor \U$30525 ( \38845_39145 , \38838_39138 , \38844_39144 );
buf \U$30526 ( \38846_39146 , \38845_39145 );
and \U$30527 ( \38847_39147 , \17437_17297 , \34343_34643_nG9ba2 );
and \U$30528 ( \38848_39148 , \16995_17294 , \34794_35094_nG9b9f );
or \U$30529 ( \38849_39149 , \38847_39147 , \38848_39148 );
xor \U$30530 ( \38850_39150 , \16994_17293 , \38849_39149 );
buf \U$30531 ( \38851_39151 , \38850_39150 );
buf \U$30533 ( \38852_39152 , \38851_39151 );
xor \U$30534 ( \38853_39153 , \38846_39146 , \38852_39152 );
and \U$30535 ( \38854_39154 , \16405_15940 , \35270_35570_nG9b9c );
and \U$30536 ( \38855_39155 , \15638_15937 , \35501_35801_nG9b99 );
or \U$30537 ( \38856_39156 , \38854_39154 , \38855_39155 );
xor \U$30538 ( \38857_39157 , \15637_15936 , \38856_39156 );
buf \U$30539 ( \38858_39158 , \38857_39157 );
buf \U$30541 ( \38859_39159 , \38858_39158 );
xor \U$30542 ( \38860_39160 , \38853_39153 , \38859_39159 );
buf \U$30543 ( \38861_39161 , \38860_39160 );
and \U$30544 ( \38862_39162 , \38445_38745 , \38451_38751 );
and \U$30545 ( \38863_39163 , \38445_38745 , \38458_38758 );
and \U$30546 ( \38864_39164 , \38451_38751 , \38458_38758 );
or \U$30547 ( \38865_39165 , \38862_39162 , \38863_39163 , \38864_39164 );
buf \U$30548 ( \38866_39166 , \38865_39165 );
xor \U$30549 ( \38867_39167 , \38861_39161 , \38866_39166 );
and \U$30550 ( \38868_39168 , \38569_38869 , \38575_38875 );
and \U$30551 ( \38869_39169 , \38569_38869 , \38673_38973 );
and \U$30552 ( \38870_39170 , \38575_38875 , \38673_38973 );
or \U$30553 ( \38871_39171 , \38868_39168 , \38869_39169 , \38870_39170 );
buf \U$30554 ( \38872_39172 , \38871_39171 );
xor \U$30555 ( \38873_39173 , \38867_39167 , \38872_39172 );
buf \U$30556 ( \38874_39174 , \38873_39173 );
xor \U$30557 ( \38875_39175 , \38822_39122 , \38874_39174 );
buf \U$30558 ( \38876_39176 , \38875_39175 );
and \U$30559 ( \38877_39177 , \38713_39013 , \38731_39031 );
and \U$30560 ( \38878_39178 , \38713_39013 , \38737_39037 );
and \U$30561 ( \38879_39179 , \38731_39031 , \38737_39037 );
or \U$30562 ( \38880_39180 , \38877_39177 , \38878_39178 , \38879_39179 );
buf \U$30563 ( \38881_39181 , \38880_39180 );
xor \U$30564 ( \38882_39182 , \38876_39176 , \38881_39181 );
and \U$30565 ( \38883_39183 , \38440_38740 , \38507_38807 );
and \U$30566 ( \38884_39184 , \38440_38740 , \38513_38813 );
and \U$30567 ( \38885_39185 , \38507_38807 , \38513_38813 );
or \U$30568 ( \38886_39186 , \38883_39183 , \38884_39184 , \38885_39185 );
buf \U$30569 ( \38887_39187 , \38886_39186 );
xor \U$30570 ( \38888_39188 , \38882_39182 , \38887_39187 );
buf \U$30571 ( \38889_39189 , \38888_39188 );
and \U$30572 ( \38890_39190 , \38435_38735 , \38515_38815 );
and \U$30573 ( \38891_39191 , \38435_38735 , \38521_38821 );
and \U$30574 ( \38892_39192 , \38515_38815 , \38521_38821 );
or \U$30575 ( \38893_39193 , \38890_39190 , \38891_39191 , \38892_39192 );
buf \U$30576 ( \38894_39194 , \38893_39193 );
xor \U$30577 ( \38895_39195 , \38889_39189 , \38894_39194 );
and \U$30578 ( \38896_39196 , \38563_38863 , \38675_38975 );
and \U$30579 ( \38897_39197 , \38563_38863 , \38711_39011 );
and \U$30580 ( \38898_39198 , \38675_38975 , \38711_39011 );
or \U$30581 ( \38899_39199 , \38896_39196 , \38897_39197 , \38898_39198 );
buf \U$30582 ( \38900_39200 , \38899_39199 );
and \U$30583 ( \38901_39201 , \14710_14631 , \35872_36172_nG9b96 );
and \U$30584 ( \38902_39202 , \14329_14628 , \36289_36589_nG9b93 );
or \U$30585 ( \38903_39203 , \38901_39201 , \38902_39202 );
xor \U$30586 ( \38904_39204 , \14328_14627 , \38903_39203 );
buf \U$30587 ( \38905_39205 , \38904_39204 );
buf \U$30589 ( \38906_39206 , \38905_39205 );
and \U$30590 ( \38907_39207 , \13431_13370 , \36686_36986_nG9b90 );
and \U$30591 ( \38908_39208 , \13068_13367 , \36950_37250_nG9b8d );
or \U$30592 ( \38909_39209 , \38907_39207 , \38908_39208 );
xor \U$30593 ( \38910_39210 , \13067_13366 , \38909_39209 );
buf \U$30594 ( \38911_39211 , \38910_39210 );
buf \U$30596 ( \38912_39212 , \38911_39211 );
xor \U$30597 ( \38913_39213 , \38906_39206 , \38912_39212 );
and \U$30598 ( \38914_39214 , \10996_10421 , \38037_38337_nG9b84 );
and \U$30599 ( \38915_39215 , \10119_10418 , \38363_38663_nG9b81 );
or \U$30600 ( \38916_39216 , \38914_39214 , \38915_39215 );
xor \U$30601 ( \38917_39217 , \10118_10417 , \38916_39216 );
buf \U$30602 ( \38918_39218 , \38917_39217 );
buf \U$30604 ( \38919_39219 , \38918_39218 );
xor \U$30605 ( \38920_39220 , \38913_39213 , \38919_39219 );
buf \U$30606 ( \38921_39221 , \38920_39220 );
and \U$30607 ( \38922_39222 , \38484_38784 , \38490_38790 );
and \U$30608 ( \38923_39223 , \38484_38784 , \38497_38797 );
and \U$30609 ( \38924_39224 , \38490_38790 , \38497_38797 );
or \U$30610 ( \38925_39225 , \38922_39222 , \38923_39223 , \38924_39224 );
buf \U$30611 ( \38926_39226 , \38925_39225 );
and \U$30612 ( \38927_39227 , \25044_24792 , \28300_28602_nG9bc0 );
and \U$30613 ( \38928_39228 , \24490_24789 , \28877_29179_nG9bbd );
or \U$30614 ( \38929_39229 , \38927_39227 , \38928_39228 );
xor \U$30615 ( \38930_39230 , \24489_24788 , \38929_39229 );
buf \U$30616 ( \38931_39231 , \38930_39230 );
buf \U$30618 ( \38932_39232 , \38931_39231 );
and \U$30619 ( \38933_39233 , \23495_23201 , \30064_30366_nG9bba );
and \U$30620 ( \38934_39234 , \22899_23198 , \30638_30940_nG9bb7 );
or \U$30621 ( \38935_39235 , \38933_39233 , \38934_39234 );
xor \U$30622 ( \38936_39236 , \22898_23197 , \38935_39235 );
buf \U$30623 ( \38937_39237 , \38936_39236 );
buf \U$30625 ( \38938_39238 , \38937_39237 );
xor \U$30626 ( \38939_39239 , \38932_39232 , \38938_39238 );
and \U$30627 ( \38940_39240 , \20353_20155 , \32881_33181_nG9bae );
and \U$30628 ( \38941_39241 , \19853_20152 , \33313_33613_nG9bab );
or \U$30629 ( \38942_39242 , \38940_39240 , \38941_39241 );
xor \U$30630 ( \38943_39243 , \19852_20151 , \38942_39242 );
buf \U$30631 ( \38944_39244 , \38943_39243 );
buf \U$30633 ( \38945_39245 , \38944_39244 );
xor \U$30634 ( \38946_39246 , \38939_39239 , \38945_39245 );
buf \U$30635 ( \38947_39247 , \38946_39246 );
xor \U$30636 ( \38948_39248 , \38926_39226 , \38947_39247 );
and \U$30637 ( \38949_39249 , \10411_10707 , \38668_38968_nG9b7e );
and \U$30638 ( \38950_39250 , \38610_38910 , \38614_38914 );
and \U$30639 ( \38951_39251 , \38614_38914 , \38656_38956 );
and \U$30640 ( \38952_39252 , \38610_38910 , \38656_38956 );
or \U$30641 ( \38953_39253 , \38950_39250 , \38951_39251 , \38952_39252 );
and \U$30642 ( \38954_39254 , \38594_38894 , \38598_38898 );
and \U$30643 ( \38955_39255 , \38598_38898 , \38603_38903 );
and \U$30644 ( \38956_39256 , \38594_38894 , \38603_38903 );
or \U$30645 ( \38957_39257 , \38954_39254 , \38955_39255 , \38956_39256 );
and \U$30646 ( \38958_39258 , \38645_38945 , \38649_38949 );
and \U$30647 ( \38959_39259 , \38649_38949 , \38654_38954 );
and \U$30648 ( \38960_39260 , \38645_38945 , \38654_38954 );
or \U$30649 ( \38961_39261 , \38958_39258 , \38959_39259 , \38960_39260 );
xor \U$30650 ( \38962_39262 , \38957_39257 , \38961_39261 );
and \U$30651 ( \38963_39263 , \38619_38919 , \38623_38923 );
and \U$30652 ( \38964_39264 , \38623_38923 , \38628_38928 );
and \U$30653 ( \38965_39265 , \38619_38919 , \38628_38928 );
or \U$30654 ( \38966_39266 , \38963_39263 , \38964_39264 , \38965_39265 );
and \U$30655 ( \38967_39267 , \38633_38933 , \38637_38937 );
and \U$30656 ( \38968_39268 , \38637_38937 , \38639_38939 );
and \U$30657 ( \38969_39269 , \38633_38933 , \38639_38939 );
or \U$30658 ( \38970_39270 , \38967_39267 , \38968_39268 , \38969_39269 );
xor \U$30659 ( \38971_39271 , \38966_39266 , \38970_39270 );
buf \U$30660 ( \38972_39272 , \38644_38944 );
xor \U$30661 ( \38973_39273 , \38971_39271 , \38972_39272 );
xor \U$30662 ( \38974_39274 , \38962_39262 , \38973_39273 );
xor \U$30663 ( \38975_39275 , \38953_39253 , \38974_39274 );
and \U$30664 ( \38976_39276 , \38629_38929 , \38640_38940 );
and \U$30665 ( \38977_39277 , \38640_38940 , \38655_38955 );
and \U$30666 ( \38978_39278 , \38629_38929 , \38655_38955 );
or \U$30667 ( \38979_39279 , \38976_39276 , \38977_39277 , \38978_39278 );
and \U$30668 ( \38980_39280 , \38585_38885 , \38589_38889 );
and \U$30669 ( \38981_39281 , \38589_38889 , \38604_38904 );
and \U$30670 ( \38982_39282 , \38585_38885 , \38604_38904 );
or \U$30671 ( \38983_39283 , \38980_39280 , \38981_39281 , \38982_39282 );
xor \U$30672 ( \38984_39284 , \38979_39279 , \38983_39283 );
and \U$30673 ( \38985_39285 , \26527_26829 , \27095_27397 );
and \U$30674 ( \38986_39286 , \27011_27313 , \26505_26807 );
nor \U$30675 ( \38987_39287 , \38985_39285 , \38986_39286 );
xnor \U$30676 ( \38988_39288 , \38987_39287 , \26993_27295 );
and \U$30677 ( \38989_39289 , \21788_22090 , \32555_32854 );
and \U$30678 ( \38990_39290 , \22257_22556 , \31765_32067 );
nor \U$30679 ( \38991_39291 , \38989_39289 , \38990_39290 );
xnor \U$30680 ( \38992_39292 , \38991_39291 , \32506_32805 );
xor \U$30681 ( \38993_39293 , \38988_39288 , \38992_39292 );
and \U$30682 ( \38994_39294 , \20734_21033 , \32503_32802 );
xor \U$30683 ( \38995_39295 , \38993_39293 , \38994_39294 );
not \U$30684 ( \38996_39296 , \20712_21011 );
and \U$30685 ( \38997_39297 , \31752_32054 , \22243_22542 );
and \U$30686 ( \38998_39298 , \32495_32794 , \21801_22103 );
nor \U$30687 ( \38999_39299 , \38997_39297 , \38998_39298 );
xnor \U$30688 ( \39000_39300 , \38999_39299 , \22249_22548 );
xor \U$30689 ( \39001_39301 , \38996_39296 , \39000_39300 );
and \U$30690 ( \39002_39302 , \28232_28534 , \25527_25826 );
and \U$30691 ( \39003_39303 , \28782_29084 , \24962_25264 );
nor \U$30692 ( \39004_39304 , \39002_39302 , \39003_39303 );
xnor \U$30693 ( \39005_39305 , \39004_39304 , \25474_25773 );
xor \U$30694 ( \39006_39306 , \39001_39301 , \39005_39305 );
xor \U$30695 ( \39007_39307 , \38995_39295 , \39006_39306 );
and \U$30696 ( \39008_39308 , \29966_30268 , \23839_24138 );
and \U$30697 ( \39009_39309 , \30500_30802 , \23328_23630 );
nor \U$30698 ( \39010_39310 , \39008_39308 , \39009_39309 );
xnor \U$30699 ( \39011_39311 , \39010_39310 , \23845_24144 );
and \U$30700 ( \39012_39312 , \24970_25272 , \28768_29070 );
and \U$30701 ( \39013_39313 , \25516_25815 , \28224_28526 );
nor \U$30702 ( \39014_39314 , \39012_39312 , \39013_39313 );
xnor \U$30703 ( \39015_39315 , \39014_39314 , \28774_29076 );
xor \U$30704 ( \39016_39316 , \39011_39311 , \39015_39315 );
and \U$30705 ( \39017_39317 , \23315_23617 , \30521_30823 );
and \U$30706 ( \39018_39318 , \23900_24199 , \29944_30246 );
nor \U$30707 ( \39019_39319 , \39017_39317 , \39018_39318 );
xnor \U$30708 ( \39020_39320 , \39019_39319 , \30511_30813 );
xor \U$30709 ( \39021_39321 , \39016_39316 , \39020_39320 );
xor \U$30710 ( \39022_39322 , \39007_39307 , \39021_39321 );
xor \U$30711 ( \39023_39323 , \38984_39284 , \39022_39322 );
xor \U$30712 ( \39024_39324 , \38975_39275 , \39023_39323 );
and \U$30713 ( \39025_39325 , \38581_38881 , \38605_38905 );
and \U$30714 ( \39026_39326 , \38605_38905 , \38657_38957 );
and \U$30715 ( \39027_39327 , \38581_38881 , \38657_38957 );
or \U$30716 ( \39028_39328 , \39025_39325 , \39026_39326 , \39027_39327 );
xor \U$30717 ( \39029_39329 , \39024_39324 , \39028_39328 );
and \U$30718 ( \39030_39330 , \38658_38958 , \38662_38962 );
and \U$30719 ( \39031_39331 , \38663_38963 , \38666_38966 );
or \U$30720 ( \39032_39332 , \39030_39330 , \39031_39331 );
xor \U$30721 ( \39033_39333 , \39029_39329 , \39032_39332 );
buf g9b7b_GF_PartitionCandidate( \39034_39334_nG9b7b , \39033_39333 );
and \U$30722 ( \39035_39335 , \10402_10704 , \39034_39334_nG9b7b );
or \U$30723 ( \39036_39336 , \38949_39249 , \39035_39335 );
xor \U$30724 ( \39037_39337 , \10399_10703 , \39036_39336 );
buf \U$30725 ( \39038_39338 , \39037_39337 );
buf \U$30727 ( \39039_39339 , \39038_39338 );
xor \U$30728 ( \39040_39340 , \38948_39248 , \39039_39339 );
buf \U$30729 ( \39041_39341 , \39040_39340 );
xor \U$30730 ( \39042_39342 , \38921_39221 , \39041_39341 );
and \U$30731 ( \39043_39343 , \38534_38834 , \38554_38854 );
and \U$30732 ( \39044_39344 , \38534_38834 , \38561_38861 );
and \U$30733 ( \39045_39345 , \38554_38854 , \38561_38861 );
or \U$30734 ( \39046_39346 , \39043_39343 , \39044_39344 , \39045_39345 );
buf \U$30735 ( \39047_39347 , \39046_39346 );
xor \U$30736 ( \39048_39348 , \39042_39342 , \39047_39347 );
buf \U$30737 ( \39049_39349 , \39048_39348 );
xor \U$30738 ( \39050_39350 , \38900_39200 , \39049_39349 );
and \U$30739 ( \39051_39351 , \38718_39018 , \38723_39023 );
and \U$30740 ( \39052_39352 , \38718_39018 , \38729_39029 );
and \U$30741 ( \39053_39353 , \38723_39023 , \38729_39029 );
or \U$30742 ( \39054_39354 , \39051_39351 , \39052_39352 , \39053_39353 );
buf \U$30743 ( \39055_39355 , \39054_39354 );
xor \U$30744 ( \39056_39356 , \39050_39350 , \39055_39355 );
buf \U$30745 ( \39057_39357 , \39056_39356 );
xor \U$30746 ( \39058_39358 , \38895_39195 , \39057_39357 );
and \U$30747 ( \39059_39359 , \38754_39054 , \39058_39358 );
and \U$30749 ( \39060_39360 , \38748_39048 , \38753_39053 );
or \U$30751 ( \39061_39361 , 1'b0 , \39060_39360 , 1'b0 );
xor \U$30752 ( \39062_39362 , \39059_39359 , \39061_39361 );
and \U$30754 ( \39063_39363 , \38741_39041 , \38747_39047 );
and \U$30755 ( \39064_39364 , \38743_39043 , \38747_39047 );
or \U$30756 ( \39065_39365 , 1'b0 , \39063_39363 , \39064_39364 );
xor \U$30757 ( \39066_39366 , \39062_39362 , \39065_39365 );
xor \U$30764 ( \39067_39367 , \39066_39366 , 1'b0 );
and \U$30765 ( \39068_39368 , \38889_39189 , \38894_39194 );
and \U$30766 ( \39069_39369 , \38889_39189 , \39057_39357 );
and \U$30767 ( \39070_39370 , \38894_39194 , \39057_39357 );
or \U$30768 ( \39071_39371 , \39068_39368 , \39069_39369 , \39070_39370 );
xor \U$30769 ( \39072_39372 , \39067_39367 , \39071_39371 );
and \U$30770 ( \39073_39373 , \38900_39200 , \39049_39349 );
and \U$30771 ( \39074_39374 , \38900_39200 , \39055_39355 );
and \U$30772 ( \39075_39375 , \39049_39349 , \39055_39355 );
or \U$30773 ( \39076_39376 , \39073_39373 , \39074_39374 , \39075_39375 );
buf \U$30774 ( \39077_39377 , \39076_39376 );
and \U$30775 ( \39078_39378 , \38861_39161 , \38866_39166 );
and \U$30776 ( \39079_39379 , \38861_39161 , \38872_39172 );
and \U$30777 ( \39080_39380 , \38866_39166 , \38872_39172 );
or \U$30778 ( \39081_39381 , \39078_39378 , \39079_39379 , \39080_39380 );
buf \U$30779 ( \39082_39382 , \39081_39381 );
and \U$30780 ( \39083_39383 , \38793_39093 , \38798_39098 );
and \U$30781 ( \39084_39384 , \38793_39093 , \38819_39119 );
and \U$30782 ( \39085_39385 , \38798_39098 , \38819_39119 );
or \U$30783 ( \39086_39386 , \39083_39383 , \39084_39384 , \39085_39385 );
buf \U$30784 ( \39087_39387 , \39086_39386 );
xor \U$30785 ( \39088_39388 , \39082_39382 , \39087_39387 );
and \U$30786 ( \39089_39389 , \38764_39064 , \38784_39084 );
and \U$30787 ( \39090_39390 , \38764_39064 , \38791_39091 );
and \U$30788 ( \39091_39391 , \38784_39084 , \38791_39091 );
or \U$30789 ( \39092_39392 , \39089_39389 , \39090_39390 , \39091_39391 );
buf \U$30790 ( \39093_39393 , \39092_39392 );
and \U$30791 ( \39094_39394 , \38835_39135 , \38837_39137 );
and \U$30792 ( \39095_39395 , \38835_39135 , \38844_39144 );
and \U$30793 ( \39096_39396 , \38837_39137 , \38844_39144 );
or \U$30794 ( \39097_39397 , \39094_39394 , \39095_39395 , \39096_39396 );
buf \U$30795 ( \39098_39398 , \39097_39397 );
and \U$30796 ( \39099_39399 , \18908_18702 , \33994_34294_nG9ba5 );
and \U$30797 ( \39100_39400 , \18400_18699 , \34343_34643_nG9ba2 );
or \U$30798 ( \39101_39401 , \39099_39399 , \39100_39400 );
xor \U$30799 ( \39102_39402 , \18399_18698 , \39101_39401 );
buf \U$30800 ( \39103_39403 , \39102_39402 );
buf \U$30802 ( \39104_39404 , \39103_39403 );
xor \U$30803 ( \39105_39405 , \39098_39398 , \39104_39404 );
and \U$30804 ( \39106_39406 , \16405_15940 , \35501_35801_nG9b99 );
and \U$30805 ( \39107_39407 , \15638_15937 , \35872_36172_nG9b96 );
or \U$30806 ( \39108_39408 , \39106_39406 , \39107_39407 );
xor \U$30807 ( \39109_39409 , \15637_15936 , \39108_39408 );
buf \U$30808 ( \39110_39410 , \39109_39409 );
buf \U$30810 ( \39111_39411 , \39110_39410 );
xor \U$30811 ( \39112_39412 , \39105_39405 , \39111_39411 );
buf \U$30812 ( \39113_39413 , \39112_39412 );
xor \U$30813 ( \39114_39414 , \39093_39393 , \39113_39413 );
and \U$30814 ( \39115_39415 , \23495_23201 , \30638_30940_nG9bb7 );
and \U$30815 ( \39116_39416 , \22899_23198 , \31877_32179_nG9bb4 );
or \U$30816 ( \39117_39417 , \39115_39415 , \39116_39416 );
xor \U$30817 ( \39118_39418 , \22898_23197 , \39117_39417 );
buf \U$30818 ( \39119_39419 , \39118_39418 );
buf \U$30820 ( \39120_39420 , \39119_39419 );
and \U$30821 ( \39121_39421 , \21908_21658 , \32589_32888_nG9bb1 );
and \U$30822 ( \39122_39422 , \21356_21655 , \32881_33181_nG9bae );
or \U$30823 ( \39123_39423 , \39121_39421 , \39122_39422 );
xor \U$30824 ( \39124_39424 , \21355_21654 , \39123_39423 );
buf \U$30825 ( \39125_39425 , \39124_39424 );
buf \U$30827 ( \39126_39426 , \39125_39425 );
xor \U$30828 ( \39127_39427 , \39120_39420 , \39126_39426 );
and \U$30829 ( \39128_39428 , \20353_20155 , \33313_33613_nG9bab );
and \U$30830 ( \39129_39429 , \19853_20152 , \33741_34041_nG9ba8 );
or \U$30831 ( \39130_39430 , \39128_39428 , \39129_39429 );
xor \U$30832 ( \39131_39431 , \19852_20151 , \39130_39430 );
buf \U$30833 ( \39132_39432 , \39131_39431 );
buf \U$30835 ( \39133_39433 , \39132_39432 );
xor \U$30836 ( \39134_39434 , \39127_39427 , \39133_39433 );
buf \U$30837 ( \39135_39435 , \39134_39434 );
xor \U$30838 ( \39136_39436 , \39114_39414 , \39135_39435 );
buf \U$30839 ( \39137_39437 , \39136_39436 );
xor \U$30840 ( \39138_39438 , \39088_39388 , \39137_39437 );
buf \U$30841 ( \39139_39439 , \39138_39438 );
xor \U$30842 ( \39140_39440 , \39077_39377 , \39139_39439 );
and \U$30843 ( \39141_39441 , \38759_39059 , \38821_39121 );
and \U$30844 ( \39142_39442 , \38759_39059 , \38874_39174 );
and \U$30845 ( \39143_39443 , \38821_39121 , \38874_39174 );
or \U$30846 ( \39144_39444 , \39141_39441 , \39142_39442 , \39143_39443 );
buf \U$30847 ( \39145_39445 , \39144_39444 );
xor \U$30848 ( \39146_39446 , \39140_39440 , \39145_39445 );
buf \U$30849 ( \39147_39447 , \39146_39446 );
and \U$30850 ( \39148_39448 , \38876_39176 , \38881_39181 );
and \U$30851 ( \39149_39449 , \38876_39176 , \38887_39187 );
and \U$30852 ( \39150_39450 , \38881_39181 , \38887_39187 );
or \U$30853 ( \39151_39451 , \39148_39448 , \39149_39449 , \39150_39450 );
buf \U$30854 ( \39152_39452 , \39151_39451 );
xor \U$30855 ( \39153_39453 , \39147_39447 , \39152_39452 );
and \U$30856 ( \39154_39454 , \38921_39221 , \39041_39341 );
and \U$30857 ( \39155_39455 , \38921_39221 , \39047_39347 );
and \U$30858 ( \39156_39456 , \39041_39341 , \39047_39347 );
or \U$30859 ( \39157_39457 , \39154_39454 , \39155_39455 , \39156_39456 );
buf \U$30860 ( \39158_39458 , \39157_39457 );
and \U$30861 ( \39159_39459 , \38926_39226 , \38947_39247 );
and \U$30862 ( \39160_39460 , \38926_39226 , \39039_39339 );
and \U$30863 ( \39161_39461 , \38947_39247 , \39039_39339 );
or \U$30864 ( \39162_39462 , \39159_39459 , \39160_39460 , \39161_39461 );
buf \U$30865 ( \39163_39463 , \39162_39462 );
and \U$30866 ( \39164_39464 , \28946_28118 , \25561_25860_nG9bc9 );
and \U$30867 ( \39165_39465 , \27816_28115 , \26585_26887_nG9bc6 );
or \U$30868 ( \39166_39466 , \39164_39464 , \39165_39465 );
xor \U$30869 ( \39167_39467 , \27815_28114 , \39166_39466 );
buf \U$30870 ( \39168_39468 , \39167_39467 );
buf \U$30872 ( \39169_39469 , \39168_39468 );
and \U$30873 ( \39170_39470 , \27141_26431 , \27114_27416_nG9bc3 );
and \U$30874 ( \39171_39471 , \26129_26428 , \28300_28602_nG9bc0 );
or \U$30875 ( \39172_39472 , \39170_39470 , \39171_39471 );
xor \U$30876 ( \39173_39473 , \26128_26427 , \39172_39472 );
buf \U$30877 ( \39174_39474 , \39173_39473 );
buf \U$30879 ( \39175_39475 , \39174_39474 );
xor \U$30880 ( \39176_39476 , \39169_39469 , \39175_39475 );
and \U$30881 ( \39177_39477 , \25044_24792 , \28877_29179_nG9bbd );
and \U$30882 ( \39178_39478 , \24490_24789 , \30064_30366_nG9bba );
or \U$30883 ( \39179_39479 , \39177_39477 , \39178_39478 );
xor \U$30884 ( \39180_39480 , \24489_24788 , \39179_39479 );
buf \U$30885 ( \39181_39481 , \39180_39480 );
buf \U$30887 ( \39182_39482 , \39181_39481 );
xor \U$30888 ( \39183_39483 , \39176_39476 , \39182_39482 );
buf \U$30889 ( \39184_39484 , \39183_39483 );
and \U$30891 ( \39185_39485 , \32617_32916 , \21827_22129_nG9bd8 );
or \U$30892 ( \39186_39486 , 1'b0 , \39185_39485 );
xor \U$30893 ( \39187_39487 , 1'b0 , \39186_39486 );
buf \U$30894 ( \39188_39488 , \39187_39487 );
buf \U$30896 ( \39189_39489 , \39188_39488 );
and \U$30897 ( \39190_39490 , \31989_31636 , \22330_22629_nG9bd5 );
and \U$30898 ( \39191_39491 , \31334_31633 , \23394_23696_nG9bd2 );
or \U$30899 ( \39192_39492 , \39190_39490 , \39191_39491 );
xor \U$30900 ( \39193_39493 , \31333_31632 , \39192_39492 );
buf \U$30901 ( \39194_39494 , \39193_39493 );
buf \U$30903 ( \39195_39495 , \39194_39494 );
xor \U$30904 ( \39196_39496 , \39189_39489 , \39195_39495 );
buf \U$30905 ( \39197_39497 , \39196_39496 );
and \U$30906 ( \39198_39498 , \38827_39127 , \38833_39133 );
buf \U$30907 ( \39199_39499 , \39198_39498 );
xor \U$30908 ( \39200_39500 , \39197_39497 , \39199_39499 );
and \U$30909 ( \39201_39501 , \30670_29853 , \23927_24226_nG9bcf );
and \U$30910 ( \39202_39502 , \29551_29850 , \24996_25298_nG9bcc );
or \U$30911 ( \39203_39503 , \39201_39501 , \39202_39502 );
xor \U$30912 ( \39204_39504 , \29550_29849 , \39203_39503 );
buf \U$30913 ( \39205_39505 , \39204_39504 );
buf \U$30915 ( \39206_39506 , \39205_39505 );
xor \U$30916 ( \39207_39507 , \39200_39500 , \39206_39506 );
buf \U$30917 ( \39208_39508 , \39207_39507 );
xor \U$30918 ( \39209_39509 , \39184_39484 , \39208_39508 );
and \U$30919 ( \39210_39510 , \10411_10707 , \39034_39334_nG9b7b );
and \U$30920 ( \39211_39511 , \38957_39257 , \38961_39261 );
and \U$30921 ( \39212_39512 , \38961_39261 , \38973_39273 );
and \U$30922 ( \39213_39513 , \38957_39257 , \38973_39273 );
or \U$30923 ( \39214_39514 , \39211_39511 , \39212_39512 , \39213_39513 );
and \U$30924 ( \39215_39515 , \38979_39279 , \38983_39283 );
and \U$30925 ( \39216_39516 , \38983_39283 , \39022_39322 );
and \U$30926 ( \39217_39517 , \38979_39279 , \39022_39322 );
or \U$30927 ( \39218_39518 , \39215_39515 , \39216_39516 , \39217_39517 );
xor \U$30928 ( \39219_39519 , \39214_39514 , \39218_39518 );
and \U$30929 ( \39220_39520 , \38995_39295 , \39006_39306 );
and \U$30930 ( \39221_39521 , \39006_39306 , \39021_39321 );
and \U$30931 ( \39222_39522 , \38995_39295 , \39021_39321 );
or \U$30932 ( \39223_39523 , \39220_39520 , \39221_39521 , \39222_39522 );
and \U$30933 ( \39224_39524 , \38988_39288 , \38992_39292 );
and \U$30934 ( \39225_39525 , \38992_39292 , \38994_39294 );
and \U$30935 ( \39226_39526 , \38988_39288 , \38994_39294 );
or \U$30936 ( \39227_39527 , \39224_39524 , \39225_39525 , \39226_39526 );
and \U$30937 ( \39228_39528 , \39011_39311 , \39015_39315 );
and \U$30938 ( \39229_39529 , \39015_39315 , \39020_39320 );
and \U$30939 ( \39230_39530 , \39011_39311 , \39020_39320 );
or \U$30940 ( \39231_39531 , \39228_39528 , \39229_39529 , \39230_39530 );
xor \U$30941 ( \39232_39532 , \39227_39527 , \39231_39531 );
and \U$30942 ( \39233_39533 , \28782_29084 , \25527_25826 );
and \U$30943 ( \39234_39534 , \29966_30268 , \24962_25264 );
nor \U$30944 ( \39235_39535 , \39233_39533 , \39234_39534 );
xnor \U$30945 ( \39236_39536 , \39235_39535 , \25474_25773 );
and \U$30946 ( \39237_39537 , \25516_25815 , \28768_29070 );
and \U$30947 ( \39238_39538 , \26527_26829 , \28224_28526 );
nor \U$30948 ( \39239_39539 , \39237_39537 , \39238_39538 );
xnor \U$30949 ( \39240_39540 , \39239_39539 , \28774_29076 );
xor \U$30950 ( \39241_39541 , \39236_39536 , \39240_39540 );
and \U$30951 ( \39242_39542 , \23900_24199 , \30521_30823 );
and \U$30952 ( \39243_39543 , \24970_25272 , \29944_30246 );
nor \U$30953 ( \39244_39544 , \39242_39542 , \39243_39543 );
xnor \U$30954 ( \39245_39545 , \39244_39544 , \30511_30813 );
xor \U$30955 ( \39246_39546 , \39241_39541 , \39245_39545 );
xor \U$30956 ( \39247_39547 , \39232_39532 , \39246_39546 );
xor \U$30957 ( \39248_39548 , \39223_39523 , \39247_39547 );
and \U$30958 ( \39249_39549 , \38966_39266 , \38970_39270 );
and \U$30959 ( \39250_39550 , \38970_39270 , \38972_39272 );
and \U$30960 ( \39251_39551 , \38966_39266 , \38972_39272 );
or \U$30961 ( \39252_39552 , \39249_39549 , \39250_39550 , \39251_39551 );
and \U$30962 ( \39253_39553 , \30500_30802 , \23839_24138 );
and \U$30963 ( \39254_39554 , \31752_32054 , \23328_23630 );
nor \U$30964 ( \39255_39555 , \39253_39553 , \39254_39554 );
xnor \U$30965 ( \39256_39556 , \39255_39555 , \23845_24144 );
and \U$30966 ( \39257_39557 , \27011_27313 , \27095_27397 );
and \U$30967 ( \39258_39558 , \28232_28534 , \26505_26807 );
nor \U$30968 ( \39259_39559 , \39257_39557 , \39258_39558 );
xnor \U$30969 ( \39260_39560 , \39259_39559 , \26993_27295 );
xor \U$30970 ( \39261_39561 , \39256_39556 , \39260_39560 );
and \U$30971 ( \39262_39562 , \21788_22090 , \32503_32802 );
xor \U$30972 ( \39263_39563 , \39261_39561 , \39262_39562 );
xor \U$30973 ( \39264_39564 , \39252_39552 , \39263_39563 );
and \U$30974 ( \39265_39565 , \38996_39296 , \39000_39300 );
and \U$30975 ( \39266_39566 , \39000_39300 , \39005_39305 );
and \U$30976 ( \39267_39567 , \38996_39296 , \39005_39305 );
or \U$30977 ( \39268_39568 , \39265_39565 , \39266_39566 , \39267_39567 );
and \U$30978 ( \39269_39569 , \32495_32794 , \22243_22542 );
not \U$30979 ( \39270_39570 , \39269_39569 );
xnor \U$30980 ( \39271_39571 , \39270_39570 , \22249_22548 );
not \U$30981 ( \39272_39572 , \39271_39571 );
xor \U$30982 ( \39273_39573 , \39268_39568 , \39272_39572 );
and \U$30983 ( \39274_39574 , \22257_22556 , \32555_32854 );
and \U$30984 ( \39275_39575 , \23315_23617 , \31765_32067 );
nor \U$30985 ( \39276_39576 , \39274_39574 , \39275_39575 );
xnor \U$30986 ( \39277_39577 , \39276_39576 , \32506_32805 );
xor \U$30987 ( \39278_39578 , \39273_39573 , \39277_39577 );
xor \U$30988 ( \39279_39579 , \39264_39564 , \39278_39578 );
xor \U$30989 ( \39280_39580 , \39248_39548 , \39279_39579 );
xor \U$30990 ( \39281_39581 , \39219_39519 , \39280_39580 );
and \U$30991 ( \39282_39582 , \38953_39253 , \38974_39274 );
and \U$30992 ( \39283_39583 , \38974_39274 , \39023_39323 );
and \U$30993 ( \39284_39584 , \38953_39253 , \39023_39323 );
or \U$30994 ( \39285_39585 , \39282_39582 , \39283_39583 , \39284_39584 );
xor \U$30995 ( \39286_39586 , \39281_39581 , \39285_39585 );
and \U$30996 ( \39287_39587 , \39024_39324 , \39028_39328 );
and \U$30997 ( \39288_39588 , \39029_39329 , \39032_39332 );
or \U$30998 ( \39289_39589 , \39287_39587 , \39288_39588 );
xor \U$30999 ( \39290_39590 , \39286_39586 , \39289_39589 );
buf g9b78_GF_PartitionCandidate( \39291_39591_nG9b78 , \39290_39590 );
and \U$31000 ( \39292_39592 , \10402_10704 , \39291_39591_nG9b78 );
or \U$31001 ( \39293_39593 , \39210_39510 , \39292_39592 );
xor \U$31002 ( \39294_39594 , \10399_10703 , \39293_39593 );
buf \U$31003 ( \39295_39595 , \39294_39594 );
buf \U$31005 ( \39296_39596 , \39295_39595 );
xor \U$31006 ( \39297_39597 , \39209_39509 , \39296_39596 );
buf \U$31007 ( \39298_39598 , \39297_39597 );
xor \U$31008 ( \39299_39599 , \39163_39463 , \39298_39598 );
and \U$31009 ( \39300_39600 , \38906_39206 , \38912_39212 );
and \U$31010 ( \39301_39601 , \38906_39206 , \38919_39219 );
and \U$31011 ( \39302_39602 , \38912_39212 , \38919_39219 );
or \U$31012 ( \39303_39603 , \39300_39600 , \39301_39601 , \39302_39602 );
buf \U$31013 ( \39304_39604 , \39303_39603 );
xor \U$31014 ( \39305_39605 , \39299_39599 , \39304_39604 );
buf \U$31015 ( \39306_39606 , \39305_39605 );
xor \U$31016 ( \39307_39607 , \39158_39458 , \39306_39606 );
and \U$31017 ( \39308_39608 , \38846_39146 , \38852_39152 );
and \U$31018 ( \39309_39609 , \38846_39146 , \38859_39159 );
and \U$31019 ( \39310_39610 , \38852_39152 , \38859_39159 );
or \U$31020 ( \39311_39611 , \39308_39608 , \39309_39609 , \39310_39610 );
buf \U$31021 ( \39312_39612 , \39311_39611 );
and \U$31022 ( \39313_39613 , \38804_39104 , \38810_39110 );
and \U$31023 ( \39314_39614 , \38804_39104 , \38817_39117 );
and \U$31024 ( \39315_39615 , \38810_39110 , \38817_39117 );
or \U$31025 ( \39316_39616 , \39313_39613 , \39314_39614 , \39315_39615 );
buf \U$31026 ( \39317_39617 , \39316_39616 );
xor \U$31027 ( \39318_39618 , \39312_39612 , \39317_39617 );
and \U$31028 ( \39319_39619 , \38932_39232 , \38938_39238 );
and \U$31029 ( \39320_39620 , \38932_39232 , \38945_39245 );
and \U$31030 ( \39321_39621 , \38938_39238 , \38945_39245 );
or \U$31031 ( \39322_39622 , \39319_39619 , \39320_39620 , \39321_39621 );
buf \U$31032 ( \39323_39623 , \39322_39622 );
xor \U$31033 ( \39324_39624 , \39318_39618 , \39323_39623 );
buf \U$31034 ( \39325_39625 , \39324_39624 );
and \U$31035 ( \39326_39626 , \17437_17297 , \34794_35094_nG9b9f );
and \U$31036 ( \39327_39627 , \16995_17294 , \35270_35570_nG9b9c );
or \U$31037 ( \39328_39628 , \39326_39626 , \39327_39627 );
xor \U$31038 ( \39329_39629 , \16994_17293 , \39328_39628 );
buf \U$31039 ( \39330_39630 , \39329_39629 );
buf \U$31041 ( \39331_39631 , \39330_39630 );
and \U$31042 ( \39332_39632 , \13431_13370 , \36950_37250_nG9b8d );
and \U$31043 ( \39333_39633 , \13068_13367 , \37307_37607_nG9b8a );
or \U$31044 ( \39334_39634 , \39332_39632 , \39333_39633 );
xor \U$31045 ( \39335_39635 , \13067_13366 , \39334_39634 );
buf \U$31046 ( \39336_39636 , \39335_39635 );
buf \U$31048 ( \39337_39637 , \39336_39636 );
xor \U$31049 ( \39338_39638 , \39331_39631 , \39337_39637 );
and \U$31050 ( \39339_39639 , \10996_10421 , \38363_38663_nG9b81 );
and \U$31051 ( \39340_39640 , \10119_10418 , \38668_38968_nG9b7e );
or \U$31052 ( \39341_39641 , \39339_39639 , \39340_39640 );
xor \U$31053 ( \39342_39642 , \10118_10417 , \39341_39641 );
buf \U$31054 ( \39343_39643 , \39342_39642 );
buf \U$31056 ( \39344_39644 , \39343_39643 );
xor \U$31057 ( \39345_39645 , \39338_39638 , \39344_39644 );
buf \U$31058 ( \39346_39646 , \39345_39645 );
xor \U$31059 ( \39347_39647 , \39325_39625 , \39346_39646 );
and \U$31060 ( \39348_39648 , \38769_39069 , \38775_39075 );
and \U$31061 ( \39349_39649 , \38769_39069 , \38782_39082 );
and \U$31062 ( \39350_39650 , \38775_39075 , \38782_39082 );
or \U$31063 ( \39351_39651 , \39348_39648 , \39349_39649 , \39350_39650 );
buf \U$31064 ( \39352_39652 , \39351_39651 );
and \U$31065 ( \39353_39653 , \14710_14631 , \36289_36589_nG9b93 );
and \U$31066 ( \39354_39654 , \14329_14628 , \36686_36986_nG9b90 );
or \U$31067 ( \39355_39655 , \39353_39653 , \39354_39654 );
xor \U$31068 ( \39356_39656 , \14328_14627 , \39355_39655 );
buf \U$31069 ( \39357_39657 , \39356_39656 );
buf \U$31071 ( \39358_39658 , \39357_39657 );
xor \U$31072 ( \39359_39659 , \39352_39652 , \39358_39658 );
and \U$31073 ( \39360_39660 , \12183_12157 , \37674_37974_nG9b87 );
and \U$31074 ( \39361_39661 , \11855_12154 , \38037_38337_nG9b84 );
or \U$31075 ( \39362_39662 , \39360_39660 , \39361_39661 );
xor \U$31076 ( \39363_39663 , \11854_12153 , \39362_39662 );
buf \U$31077 ( \39364_39664 , \39363_39663 );
buf \U$31079 ( \39365_39665 , \39364_39664 );
xor \U$31080 ( \39366_39666 , \39359_39659 , \39365_39665 );
buf \U$31081 ( \39367_39667 , \39366_39666 );
xor \U$31082 ( \39368_39668 , \39347_39647 , \39367_39667 );
buf \U$31083 ( \39369_39669 , \39368_39668 );
xor \U$31084 ( \39370_39670 , \39307_39607 , \39369_39669 );
buf \U$31085 ( \39371_39671 , \39370_39670 );
xor \U$31086 ( \39372_39672 , \39153_39453 , \39371_39671 );
and \U$31087 ( \39373_39673 , \39072_39372 , \39372_39672 );
and \U$31089 ( \39374_39674 , \39066_39366 , \39071_39371 );
or \U$31091 ( \39375_39675 , 1'b0 , \39374_39674 , 1'b0 );
xor \U$31092 ( \39376_39676 , \39373_39673 , \39375_39675 );
and \U$31094 ( \39377_39677 , \39059_39359 , \39065_39365 );
and \U$31095 ( \39378_39678 , \39061_39361 , \39065_39365 );
or \U$31096 ( \39379_39679 , 1'b0 , \39377_39677 , \39378_39678 );
xor \U$31097 ( \39380_39680 , \39376_39676 , \39379_39679 );
xor \U$31104 ( \39381_39681 , \39380_39680 , 1'b0 );
and \U$31105 ( \39382_39682 , \39158_39458 , \39306_39606 );
and \U$31106 ( \39383_39683 , \39158_39458 , \39369_39669 );
and \U$31107 ( \39384_39684 , \39306_39606 , \39369_39669 );
or \U$31108 ( \39385_39685 , \39382_39682 , \39383_39683 , \39384_39684 );
buf \U$31109 ( \39386_39686 , \39385_39685 );
and \U$31110 ( \39387_39687 , \39163_39463 , \39298_39598 );
and \U$31111 ( \39388_39688 , \39163_39463 , \39304_39604 );
and \U$31112 ( \39389_39689 , \39298_39598 , \39304_39604 );
or \U$31113 ( \39390_39690 , \39387_39687 , \39388_39688 , \39389_39689 );
buf \U$31114 ( \39391_39691 , \39390_39690 );
and \U$31115 ( \39392_39692 , \39184_39484 , \39208_39508 );
and \U$31116 ( \39393_39693 , \39184_39484 , \39296_39596 );
and \U$31117 ( \39394_39694 , \39208_39508 , \39296_39596 );
or \U$31118 ( \39395_39695 , \39392_39692 , \39393_39693 , \39394_39694 );
buf \U$31119 ( \39396_39696 , \39395_39695 );
and \U$31120 ( \39397_39697 , \39331_39631 , \39337_39637 );
and \U$31121 ( \39398_39698 , \39331_39631 , \39344_39644 );
and \U$31122 ( \39399_39699 , \39337_39637 , \39344_39644 );
or \U$31123 ( \39400_39700 , \39397_39697 , \39398_39698 , \39399_39699 );
buf \U$31124 ( \39401_39701 , \39400_39700 );
xor \U$31125 ( \39402_39702 , \39396_39696 , \39401_39701 );
and \U$31126 ( \39403_39703 , \39352_39652 , \39358_39658 );
and \U$31127 ( \39404_39704 , \39352_39652 , \39365_39665 );
and \U$31128 ( \39405_39705 , \39358_39658 , \39365_39665 );
or \U$31129 ( \39406_39706 , \39403_39703 , \39404_39704 , \39405_39705 );
buf \U$31130 ( \39407_39707 , \39406_39706 );
xor \U$31131 ( \39408_39708 , \39402_39702 , \39407_39707 );
buf \U$31132 ( \39409_39709 , \39408_39708 );
xor \U$31133 ( \39410_39710 , \39391_39691 , \39409_39709 );
and \U$31134 ( \39411_39711 , \39093_39393 , \39113_39413 );
and \U$31135 ( \39412_39712 , \39093_39393 , \39135_39435 );
and \U$31136 ( \39413_39713 , \39113_39413 , \39135_39435 );
or \U$31137 ( \39414_39714 , \39411_39711 , \39412_39712 , \39413_39713 );
buf \U$31138 ( \39415_39715 , \39414_39714 );
xor \U$31139 ( \39416_39716 , \39410_39710 , \39415_39715 );
buf \U$31140 ( \39417_39717 , \39416_39716 );
xor \U$31141 ( \39418_39718 , \39386_39686 , \39417_39717 );
and \U$31142 ( \39419_39719 , \39082_39382 , \39087_39387 );
and \U$31143 ( \39420_39720 , \39082_39382 , \39137_39437 );
and \U$31144 ( \39421_39721 , \39087_39387 , \39137_39437 );
or \U$31145 ( \39422_39722 , \39419_39719 , \39420_39720 , \39421_39721 );
buf \U$31146 ( \39423_39723 , \39422_39722 );
xor \U$31147 ( \39424_39724 , \39418_39718 , \39423_39723 );
buf \U$31148 ( \39425_39725 , \39424_39724 );
and \U$31149 ( \39426_39726 , \39077_39377 , \39139_39439 );
and \U$31150 ( \39427_39727 , \39077_39377 , \39145_39445 );
and \U$31151 ( \39428_39728 , \39139_39439 , \39145_39445 );
or \U$31152 ( \39429_39729 , \39426_39726 , \39427_39727 , \39428_39728 );
buf \U$31153 ( \39430_39730 , \39429_39729 );
xor \U$31154 ( \39431_39731 , \39425_39725 , \39430_39730 );
and \U$31155 ( \39432_39732 , \39325_39625 , \39346_39646 );
and \U$31156 ( \39433_39733 , \39325_39625 , \39367_39667 );
and \U$31157 ( \39434_39734 , \39346_39646 , \39367_39667 );
or \U$31158 ( \39435_39735 , \39432_39732 , \39433_39733 , \39434_39734 );
buf \U$31159 ( \39436_39736 , \39435_39735 );
and \U$31160 ( \39437_39737 , \39189_39489 , \39195_39495 );
buf \U$31161 ( \39438_39738 , \39437_39737 );
and \U$31162 ( \39439_39739 , \30670_29853 , \24996_25298_nG9bcc );
and \U$31163 ( \39440_39740 , \29551_29850 , \25561_25860_nG9bc9 );
or \U$31164 ( \39441_39741 , \39439_39739 , \39440_39740 );
xor \U$31165 ( \39442_39742 , \29550_29849 , \39441_39741 );
buf \U$31166 ( \39443_39743 , \39442_39742 );
buf \U$31168 ( \39444_39744 , \39443_39743 );
xor \U$31169 ( \39445_39745 , \39438_39738 , \39444_39744 );
and \U$31170 ( \39446_39746 , \28946_28118 , \26585_26887_nG9bc6 );
and \U$31171 ( \39447_39747 , \27816_28115 , \27114_27416_nG9bc3 );
or \U$31172 ( \39448_39748 , \39446_39746 , \39447_39747 );
xor \U$31173 ( \39449_39749 , \27815_28114 , \39448_39748 );
buf \U$31174 ( \39450_39750 , \39449_39749 );
buf \U$31176 ( \39451_39751 , \39450_39750 );
xor \U$31177 ( \39452_39752 , \39445_39745 , \39451_39751 );
buf \U$31178 ( \39453_39753 , \39452_39752 );
and \U$31179 ( \39454_39754 , \39120_39420 , \39126_39426 );
and \U$31180 ( \39455_39755 , \39120_39420 , \39133_39433 );
and \U$31181 ( \39456_39756 , \39126_39426 , \39133_39433 );
or \U$31182 ( \39457_39757 , \39454_39754 , \39455_39755 , \39456_39756 );
buf \U$31183 ( \39458_39758 , \39457_39757 );
xor \U$31184 ( \39459_39759 , \39453_39753 , \39458_39758 );
and \U$31185 ( \39460_39760 , \12183_12157 , \38037_38337_nG9b84 );
and \U$31186 ( \39461_39761 , \11855_12154 , \38363_38663_nG9b81 );
or \U$31187 ( \39462_39762 , \39460_39760 , \39461_39761 );
xor \U$31188 ( \39463_39763 , \11854_12153 , \39462_39762 );
buf \U$31189 ( \39464_39764 , \39463_39763 );
buf \U$31191 ( \39465_39765 , \39464_39764 );
xor \U$31192 ( \39466_39766 , \39459_39759 , \39465_39765 );
buf \U$31193 ( \39467_39767 , \39466_39766 );
and \U$31194 ( \39468_39768 , \14710_14631 , \36686_36986_nG9b90 );
and \U$31195 ( \39469_39769 , \14329_14628 , \36950_37250_nG9b8d );
or \U$31196 ( \39470_39770 , \39468_39768 , \39469_39769 );
xor \U$31197 ( \39471_39771 , \14328_14627 , \39470_39770 );
buf \U$31198 ( \39472_39772 , \39471_39771 );
buf \U$31200 ( \39473_39773 , \39472_39772 );
and \U$31201 ( \39474_39774 , \13431_13370 , \37307_37607_nG9b8a );
and \U$31202 ( \39475_39775 , \13068_13367 , \37674_37974_nG9b87 );
or \U$31203 ( \39476_39776 , \39474_39774 , \39475_39775 );
xor \U$31204 ( \39477_39777 , \13067_13366 , \39476_39776 );
buf \U$31205 ( \39478_39778 , \39477_39777 );
buf \U$31207 ( \39479_39779 , \39478_39778 );
xor \U$31208 ( \39480_39780 , \39473_39773 , \39479_39779 );
and \U$31209 ( \39481_39781 , \10996_10421 , \38668_38968_nG9b7e );
and \U$31210 ( \39482_39782 , \10119_10418 , \39034_39334_nG9b7b );
or \U$31211 ( \39483_39783 , \39481_39781 , \39482_39782 );
xor \U$31212 ( \39484_39784 , \10118_10417 , \39483_39783 );
buf \U$31213 ( \39485_39785 , \39484_39784 );
buf \U$31215 ( \39486_39786 , \39485_39785 );
xor \U$31216 ( \39487_39787 , \39480_39780 , \39486_39786 );
buf \U$31217 ( \39488_39788 , \39487_39787 );
xor \U$31218 ( \39489_39789 , \39467_39767 , \39488_39788 );
and \U$31219 ( \39490_39790 , \39197_39497 , \39199_39499 );
and \U$31220 ( \39491_39791 , \39197_39497 , \39206_39506 );
and \U$31221 ( \39492_39792 , \39199_39499 , \39206_39506 );
or \U$31222 ( \39493_39793 , \39490_39790 , \39491_39791 , \39492_39792 );
buf \U$31223 ( \39494_39794 , \39493_39793 );
and \U$31224 ( \39495_39795 , \18908_18702 , \34343_34643_nG9ba2 );
and \U$31225 ( \39496_39796 , \18400_18699 , \34794_35094_nG9b9f );
or \U$31226 ( \39497_39797 , \39495_39795 , \39496_39796 );
xor \U$31227 ( \39498_39798 , \18399_18698 , \39497_39797 );
buf \U$31228 ( \39499_39799 , \39498_39798 );
buf \U$31230 ( \39500_39800 , \39499_39799 );
xor \U$31231 ( \39501_39801 , \39494_39794 , \39500_39800 );
and \U$31232 ( \39502_39802 , \17437_17297 , \35270_35570_nG9b9c );
and \U$31233 ( \39503_39803 , \16995_17294 , \35501_35801_nG9b99 );
or \U$31234 ( \39504_39804 , \39502_39802 , \39503_39803 );
xor \U$31235 ( \39505_39805 , \16994_17293 , \39504_39804 );
buf \U$31236 ( \39506_39806 , \39505_39805 );
buf \U$31238 ( \39507_39807 , \39506_39806 );
xor \U$31239 ( \39508_39808 , \39501_39801 , \39507_39807 );
buf \U$31240 ( \39509_39809 , \39508_39808 );
xor \U$31241 ( \39510_39810 , \39489_39789 , \39509_39809 );
buf \U$31242 ( \39511_39811 , \39510_39810 );
xor \U$31243 ( \39512_39812 , \39436_39736 , \39511_39811 );
and \U$31244 ( \39513_39813 , \39098_39398 , \39104_39404 );
and \U$31245 ( \39514_39814 , \39098_39398 , \39111_39411 );
and \U$31246 ( \39515_39815 , \39104_39404 , \39111_39411 );
or \U$31247 ( \39516_39816 , \39513_39813 , \39514_39814 , \39515_39815 );
buf \U$31248 ( \39517_39817 , \39516_39816 );
and \U$31249 ( \39518_39818 , \23495_23201 , \31877_32179_nG9bb4 );
and \U$31250 ( \39519_39819 , \22899_23198 , \32589_32888_nG9bb1 );
or \U$31251 ( \39520_39820 , \39518_39818 , \39519_39819 );
xor \U$31252 ( \39521_39821 , \22898_23197 , \39520_39820 );
buf \U$31253 ( \39522_39822 , \39521_39821 );
buf \U$31255 ( \39523_39823 , \39522_39822 );
and \U$31256 ( \39524_39824 , \21908_21658 , \32881_33181_nG9bae );
and \U$31257 ( \39525_39825 , \21356_21655 , \33313_33613_nG9bab );
or \U$31258 ( \39526_39826 , \39524_39824 , \39525_39825 );
xor \U$31259 ( \39527_39827 , \21355_21654 , \39526_39826 );
buf \U$31260 ( \39528_39828 , \39527_39827 );
buf \U$31262 ( \39529_39829 , \39528_39828 );
xor \U$31263 ( \39530_39830 , \39523_39823 , \39529_39829 );
and \U$31264 ( \39531_39831 , \20353_20155 , \33741_34041_nG9ba8 );
and \U$31265 ( \39532_39832 , \19853_20152 , \33994_34294_nG9ba5 );
or \U$31266 ( \39533_39833 , \39531_39831 , \39532_39832 );
xor \U$31267 ( \39534_39834 , \19852_20151 , \39533_39833 );
buf \U$31268 ( \39535_39835 , \39534_39834 );
buf \U$31270 ( \39536_39836 , \39535_39835 );
xor \U$31271 ( \39537_39837 , \39530_39830 , \39536_39836 );
buf \U$31272 ( \39538_39838 , \39537_39837 );
xor \U$31273 ( \39539_39839 , \39517_39817 , \39538_39838 );
and \U$31275 ( \39540_39840 , \32617_32916 , \22330_22629_nG9bd5 );
or \U$31276 ( \39541_39841 , 1'b0 , \39540_39840 );
xor \U$31277 ( \39542_39842 , 1'b0 , \39541_39841 );
buf \U$31278 ( \39543_39843 , \39542_39842 );
buf \U$31280 ( \39544_39844 , \39543_39843 );
and \U$31281 ( \39545_39845 , \31989_31636 , \23394_23696_nG9bd2 );
and \U$31282 ( \39546_39846 , \31334_31633 , \23927_24226_nG9bcf );
or \U$31283 ( \39547_39847 , \39545_39845 , \39546_39846 );
xor \U$31284 ( \39548_39848 , \31333_31632 , \39547_39847 );
buf \U$31285 ( \39549_39849 , \39548_39848 );
buf \U$31287 ( \39550_39850 , \39549_39849 );
xor \U$31288 ( \39551_39851 , \39544_39844 , \39550_39850 );
buf \U$31289 ( \39552_39852 , \39551_39851 );
and \U$31290 ( \39553_39853 , \27141_26431 , \28300_28602_nG9bc0 );
and \U$31291 ( \39554_39854 , \26129_26428 , \28877_29179_nG9bbd );
or \U$31292 ( \39555_39855 , \39553_39853 , \39554_39854 );
xor \U$31293 ( \39556_39856 , \26128_26427 , \39555_39855 );
buf \U$31294 ( \39557_39857 , \39556_39856 );
buf \U$31296 ( \39558_39858 , \39557_39857 );
xor \U$31297 ( \39559_39859 , \39552_39852 , \39558_39858 );
and \U$31298 ( \39560_39860 , \25044_24792 , \30064_30366_nG9bba );
and \U$31299 ( \39561_39861 , \24490_24789 , \30638_30940_nG9bb7 );
or \U$31300 ( \39562_39862 , \39560_39860 , \39561_39861 );
xor \U$31301 ( \39563_39863 , \24489_24788 , \39562_39862 );
buf \U$31302 ( \39564_39864 , \39563_39863 );
buf \U$31304 ( \39565_39865 , \39564_39864 );
xor \U$31305 ( \39566_39866 , \39559_39859 , \39565_39865 );
buf \U$31306 ( \39567_39867 , \39566_39866 );
xor \U$31307 ( \39568_39868 , \39539_39839 , \39567_39867 );
buf \U$31308 ( \39569_39869 , \39568_39868 );
and \U$31309 ( \39570_39870 , \39312_39612 , \39317_39617 );
and \U$31310 ( \39571_39871 , \39312_39612 , \39323_39623 );
and \U$31311 ( \39572_39872 , \39317_39617 , \39323_39623 );
or \U$31312 ( \39573_39873 , \39570_39870 , \39571_39871 , \39572_39872 );
buf \U$31313 ( \39574_39874 , \39573_39873 );
xor \U$31314 ( \39575_39875 , \39569_39869 , \39574_39874 );
and \U$31315 ( \39576_39876 , \39169_39469 , \39175_39475 );
and \U$31316 ( \39577_39877 , \39169_39469 , \39182_39482 );
and \U$31317 ( \39578_39878 , \39175_39475 , \39182_39482 );
or \U$31318 ( \39579_39879 , \39576_39876 , \39577_39877 , \39578_39878 );
buf \U$31319 ( \39580_39880 , \39579_39879 );
and \U$31320 ( \39581_39881 , \16405_15940 , \35872_36172_nG9b96 );
and \U$31321 ( \39582_39882 , \15638_15937 , \36289_36589_nG9b93 );
or \U$31322 ( \39583_39883 , \39581_39881 , \39582_39882 );
xor \U$31323 ( \39584_39884 , \15637_15936 , \39583_39883 );
buf \U$31324 ( \39585_39885 , \39584_39884 );
buf \U$31326 ( \39586_39886 , \39585_39885 );
xor \U$31327 ( \39587_39887 , \39580_39880 , \39586_39886 );
and \U$31328 ( \39588_39888 , \10411_10707 , \39291_39591_nG9b78 );
and \U$31329 ( \39589_39889 , \39223_39523 , \39247_39547 );
and \U$31330 ( \39590_39890 , \39247_39547 , \39279_39579 );
and \U$31331 ( \39591_39891 , \39223_39523 , \39279_39579 );
or \U$31332 ( \39592_39892 , \39589_39889 , \39590_39890 , \39591_39891 );
and \U$31333 ( \39593_39893 , \39268_39568 , \39272_39572 );
and \U$31334 ( \39594_39894 , \39272_39572 , \39277_39577 );
and \U$31335 ( \39595_39895 , \39268_39568 , \39277_39577 );
or \U$31336 ( \39596_39896 , \39593_39893 , \39594_39894 , \39595_39895 );
and \U$31337 ( \39597_39897 , \29966_30268 , \25527_25826 );
and \U$31338 ( \39598_39898 , \30500_30802 , \24962_25264 );
nor \U$31339 ( \39599_39899 , \39597_39897 , \39598_39898 );
xnor \U$31340 ( \39600_39900 , \39599_39899 , \25474_25773 );
and \U$31341 ( \39601_39901 , \26527_26829 , \28768_29070 );
and \U$31342 ( \39602_39902 , \27011_27313 , \28224_28526 );
nor \U$31343 ( \39603_39903 , \39601_39901 , \39602_39902 );
xnor \U$31344 ( \39604_39904 , \39603_39903 , \28774_29076 );
xor \U$31345 ( \39605_39905 , \39600_39900 , \39604_39904 );
and \U$31346 ( \39606_39906 , \22257_22556 , \32503_32802 );
xor \U$31347 ( \39607_39907 , \39605_39905 , \39606_39906 );
xor \U$31348 ( \39608_39908 , \39596_39896 , \39607_39907 );
buf \U$31349 ( \39609_39909 , \39271_39571 );
and \U$31350 ( \39610_39910 , \24970_25272 , \30521_30823 );
and \U$31351 ( \39611_39911 , \25516_25815 , \29944_30246 );
nor \U$31352 ( \39612_39912 , \39610_39910 , \39611_39911 );
xnor \U$31353 ( \39613_39913 , \39612_39912 , \30511_30813 );
xor \U$31354 ( \39614_39914 , \39609_39909 , \39613_39913 );
and \U$31355 ( \39615_39915 , \23315_23617 , \32555_32854 );
and \U$31356 ( \39616_39916 , \23900_24199 , \31765_32067 );
nor \U$31357 ( \39617_39917 , \39615_39915 , \39616_39916 );
xnor \U$31358 ( \39618_39918 , \39617_39917 , \32506_32805 );
xor \U$31359 ( \39619_39919 , \39614_39914 , \39618_39918 );
xor \U$31360 ( \39620_39920 , \39608_39908 , \39619_39919 );
xor \U$31361 ( \39621_39921 , \39592_39892 , \39620_39920 );
and \U$31362 ( \39622_39922 , \39227_39527 , \39231_39531 );
and \U$31363 ( \39623_39923 , \39231_39531 , \39246_39546 );
and \U$31364 ( \39624_39924 , \39227_39527 , \39246_39546 );
or \U$31365 ( \39625_39925 , \39622_39922 , \39623_39923 , \39624_39924 );
and \U$31366 ( \39626_39926 , \39252_39552 , \39263_39563 );
and \U$31367 ( \39627_39927 , \39263_39563 , \39278_39578 );
and \U$31368 ( \39628_39928 , \39252_39552 , \39278_39578 );
or \U$31369 ( \39629_39929 , \39626_39926 , \39627_39927 , \39628_39928 );
xor \U$31370 ( \39630_39930 , \39625_39925 , \39629_39929 );
and \U$31371 ( \39631_39931 , \39236_39536 , \39240_39540 );
and \U$31372 ( \39632_39932 , \39240_39540 , \39245_39545 );
and \U$31373 ( \39633_39933 , \39236_39536 , \39245_39545 );
or \U$31374 ( \39634_39934 , \39631_39931 , \39632_39932 , \39633_39933 );
and \U$31375 ( \39635_39935 , \39256_39556 , \39260_39560 );
and \U$31376 ( \39636_39936 , \39260_39560 , \39262_39562 );
and \U$31377 ( \39637_39937 , \39256_39556 , \39262_39562 );
or \U$31378 ( \39638_39938 , \39635_39935 , \39636_39936 , \39637_39937 );
xor \U$31379 ( \39639_39939 , \39634_39934 , \39638_39938 );
not \U$31380 ( \39640_39940 , \22249_22548 );
and \U$31381 ( \39641_39941 , \31752_32054 , \23839_24138 );
and \U$31382 ( \39642_39942 , \32495_32794 , \23328_23630 );
nor \U$31383 ( \39643_39943 , \39641_39941 , \39642_39942 );
xnor \U$31384 ( \39644_39944 , \39643_39943 , \23845_24144 );
xor \U$31385 ( \39645_39945 , \39640_39940 , \39644_39944 );
and \U$31386 ( \39646_39946 , \28232_28534 , \27095_27397 );
and \U$31387 ( \39647_39947 , \28782_29084 , \26505_26807 );
nor \U$31388 ( \39648_39948 , \39646_39946 , \39647_39947 );
xnor \U$31389 ( \39649_39949 , \39648_39948 , \26993_27295 );
xor \U$31390 ( \39650_39950 , \39645_39945 , \39649_39949 );
xor \U$31391 ( \39651_39951 , \39639_39939 , \39650_39950 );
xor \U$31392 ( \39652_39952 , \39630_39930 , \39651_39951 );
xor \U$31393 ( \39653_39953 , \39621_39921 , \39652_39952 );
and \U$31394 ( \39654_39954 , \39214_39514 , \39218_39518 );
and \U$31395 ( \39655_39955 , \39218_39518 , \39280_39580 );
and \U$31396 ( \39656_39956 , \39214_39514 , \39280_39580 );
or \U$31397 ( \39657_39957 , \39654_39954 , \39655_39955 , \39656_39956 );
xor \U$31398 ( \39658_39958 , \39653_39953 , \39657_39957 );
and \U$31399 ( \39659_39959 , \39281_39581 , \39285_39585 );
and \U$31400 ( \39660_39960 , \39286_39586 , \39289_39589 );
or \U$31401 ( \39661_39961 , \39659_39959 , \39660_39960 );
xor \U$31402 ( \39662_39962 , \39658_39958 , \39661_39961 );
buf g9b75_GF_PartitionCandidate( \39663_39963_nG9b75 , \39662_39962 );
and \U$31403 ( \39664_39964 , \10402_10704 , \39663_39963_nG9b75 );
or \U$31404 ( \39665_39965 , \39588_39888 , \39664_39964 );
xor \U$31405 ( \39666_39966 , \10399_10703 , \39665_39965 );
buf \U$31406 ( \39667_39967 , \39666_39966 );
buf \U$31408 ( \39668_39968 , \39667_39967 );
xor \U$31409 ( \39669_39969 , \39587_39887 , \39668_39968 );
buf \U$31410 ( \39670_39970 , \39669_39969 );
xor \U$31411 ( \39671_39971 , \39575_39875 , \39670_39970 );
buf \U$31412 ( \39672_39972 , \39671_39971 );
xor \U$31413 ( \39673_39973 , \39512_39812 , \39672_39972 );
buf \U$31414 ( \39674_39974 , \39673_39973 );
xor \U$31415 ( \39675_39975 , \39431_39731 , \39674_39974 );
xor \U$31416 ( \39676_39976 , \39381_39681 , \39675_39975 );
and \U$31417 ( \39677_39977 , \39147_39447 , \39152_39452 );
and \U$31418 ( \39678_39978 , \39147_39447 , \39371_39671 );
and \U$31419 ( \39679_39979 , \39152_39452 , \39371_39671 );
or \U$31420 ( \39680_39980 , \39677_39977 , \39678_39978 , \39679_39979 );
and \U$31421 ( \39681_39981 , \39676_39976 , \39680_39980 );
and \U$31423 ( \39682_39982 , \39380_39680 , \39675_39975 );
or \U$31425 ( \39683_39983 , 1'b0 , \39682_39982 , 1'b0 );
xor \U$31426 ( \39684_39984 , \39681_39981 , \39683_39983 );
and \U$31428 ( \39685_39985 , \39373_39673 , \39379_39679 );
and \U$31429 ( \39686_39986 , \39375_39675 , \39379_39679 );
or \U$31430 ( \39687_39987 , 1'b0 , \39685_39985 , \39686_39986 );
xor \U$31431 ( \39688_39988 , \39684_39984 , \39687_39987 );
xor \U$31438 ( \39689_39989 , \39688_39988 , 1'b0 );
and \U$31439 ( \39690_39990 , \39425_39725 , \39430_39730 );
and \U$31440 ( \39691_39991 , \39425_39725 , \39674_39974 );
and \U$31441 ( \39692_39992 , \39430_39730 , \39674_39974 );
or \U$31442 ( \39693_39993 , \39690_39990 , \39691_39991 , \39692_39992 );
xor \U$31443 ( \39694_39994 , \39689_39989 , \39693_39993 );
and \U$31444 ( \39695_39995 , \39436_39736 , \39511_39811 );
and \U$31445 ( \39696_39996 , \39436_39736 , \39672_39972 );
and \U$31446 ( \39697_39997 , \39511_39811 , \39672_39972 );
or \U$31447 ( \39698_39998 , \39695_39995 , \39696_39996 , \39697_39997 );
buf \U$31448 ( \39699_39999 , \39698_39998 );
and \U$31449 ( \39700_40000 , \39391_39691 , \39409_39709 );
and \U$31450 ( \39701_40001 , \39391_39691 , \39415_39715 );
and \U$31451 ( \39702_40002 , \39409_39709 , \39415_39715 );
or \U$31452 ( \39703_40003 , \39700_40000 , \39701_40001 , \39702_40002 );
buf \U$31453 ( \39704_40004 , \39703_40003 );
xor \U$31454 ( \39705_40005 , \39699_39999 , \39704_40004 );
and \U$31455 ( \39706_40006 , \39396_39696 , \39401_39701 );
and \U$31456 ( \39707_40007 , \39396_39696 , \39407_39707 );
and \U$31457 ( \39708_40008 , \39401_39701 , \39407_39707 );
or \U$31458 ( \39709_40009 , \39706_40006 , \39707_40007 , \39708_40008 );
buf \U$31459 ( \39710_40010 , \39709_40009 );
and \U$31460 ( \39711_40011 , \39467_39767 , \39488_39788 );
and \U$31461 ( \39712_40012 , \39467_39767 , \39509_39809 );
and \U$31462 ( \39713_40013 , \39488_39788 , \39509_39809 );
or \U$31463 ( \39714_40014 , \39711_40011 , \39712_40012 , \39713_40013 );
buf \U$31464 ( \39715_40015 , \39714_40014 );
xor \U$31465 ( \39716_40016 , \39710_40010 , \39715_40015 );
and \U$31466 ( \39717_40017 , \39580_39880 , \39586_39886 );
and \U$31467 ( \39718_40018 , \39580_39880 , \39668_39968 );
and \U$31468 ( \39719_40019 , \39586_39886 , \39668_39968 );
or \U$31469 ( \39720_40020 , \39717_40017 , \39718_40018 , \39719_40019 );
buf \U$31470 ( \39721_40021 , \39720_40020 );
and \U$31471 ( \39722_40022 , \39473_39773 , \39479_39779 );
and \U$31472 ( \39723_40023 , \39473_39773 , \39486_39786 );
and \U$31473 ( \39724_40024 , \39479_39779 , \39486_39786 );
or \U$31474 ( \39725_40025 , \39722_40022 , \39723_40023 , \39724_40024 );
buf \U$31475 ( \39726_40026 , \39725_40025 );
xor \U$31476 ( \39727_40027 , \39721_40021 , \39726_40026 );
and \U$31477 ( \39728_40028 , \39438_39738 , \39444_39744 );
and \U$31478 ( \39729_40029 , \39438_39738 , \39451_39751 );
and \U$31479 ( \39730_40030 , \39444_39744 , \39451_39751 );
or \U$31480 ( \39731_40031 , \39728_40028 , \39729_40029 , \39730_40030 );
buf \U$31481 ( \39732_40032 , \39731_40031 );
and \U$31482 ( \39733_40033 , \18908_18702 , \34794_35094_nG9b9f );
and \U$31483 ( \39734_40034 , \18400_18699 , \35270_35570_nG9b9c );
or \U$31484 ( \39735_40035 , \39733_40033 , \39734_40034 );
xor \U$31485 ( \39736_40036 , \18399_18698 , \39735_40035 );
buf \U$31486 ( \39737_40037 , \39736_40036 );
buf \U$31488 ( \39738_40038 , \39737_40037 );
xor \U$31489 ( \39739_40039 , \39732_40032 , \39738_40038 );
and \U$31490 ( \39740_40040 , \17437_17297 , \35501_35801_nG9b99 );
and \U$31491 ( \39741_40041 , \16995_17294 , \35872_36172_nG9b96 );
or \U$31492 ( \39742_40042 , \39740_40040 , \39741_40041 );
xor \U$31493 ( \39743_40043 , \16994_17293 , \39742_40042 );
buf \U$31494 ( \39744_40044 , \39743_40043 );
buf \U$31496 ( \39745_40045 , \39744_40044 );
xor \U$31497 ( \39746_40046 , \39739_40039 , \39745_40045 );
buf \U$31498 ( \39747_40047 , \39746_40046 );
xor \U$31499 ( \39748_40048 , \39727_40027 , \39747_40047 );
buf \U$31500 ( \39749_40049 , \39748_40048 );
xor \U$31501 ( \39750_40050 , \39716_40016 , \39749_40049 );
buf \U$31502 ( \39751_40051 , \39750_40050 );
xor \U$31503 ( \39752_40052 , \39705_40005 , \39751_40051 );
buf \U$31504 ( \39753_40053 , \39752_40052 );
and \U$31505 ( \39754_40054 , \39386_39686 , \39417_39717 );
and \U$31506 ( \39755_40055 , \39386_39686 , \39423_39723 );
and \U$31507 ( \39756_40056 , \39417_39717 , \39423_39723 );
or \U$31508 ( \39757_40057 , \39754_40054 , \39755_40055 , \39756_40056 );
buf \U$31509 ( \39758_40058 , \39757_40057 );
xor \U$31510 ( \39759_40059 , \39753_40053 , \39758_40058 );
and \U$31512 ( \39760_40060 , \32617_32916 , \23394_23696_nG9bd2 );
or \U$31513 ( \39761_40061 , 1'b0 , \39760_40060 );
xor \U$31514 ( \39762_40062 , 1'b0 , \39761_40061 );
buf \U$31515 ( \39763_40063 , \39762_40062 );
buf \U$31517 ( \39764_40064 , \39763_40063 );
and \U$31518 ( \39765_40065 , \31989_31636 , \23927_24226_nG9bcf );
and \U$31519 ( \39766_40066 , \31334_31633 , \24996_25298_nG9bcc );
or \U$31520 ( \39767_40067 , \39765_40065 , \39766_40066 );
xor \U$31521 ( \39768_40068 , \31333_31632 , \39767_40067 );
buf \U$31522 ( \39769_40069 , \39768_40068 );
buf \U$31524 ( \39770_40070 , \39769_40069 );
xor \U$31525 ( \39771_40071 , \39764_40064 , \39770_40070 );
buf \U$31526 ( \39772_40072 , \39771_40071 );
and \U$31527 ( \39773_40073 , \27141_26431 , \28877_29179_nG9bbd );
and \U$31528 ( \39774_40074 , \26129_26428 , \30064_30366_nG9bba );
or \U$31529 ( \39775_40075 , \39773_40073 , \39774_40074 );
xor \U$31530 ( \39776_40076 , \26128_26427 , \39775_40075 );
buf \U$31531 ( \39777_40077 , \39776_40076 );
buf \U$31533 ( \39778_40078 , \39777_40077 );
xor \U$31534 ( \39779_40079 , \39772_40072 , \39778_40078 );
and \U$31535 ( \39780_40080 , \25044_24792 , \30638_30940_nG9bb7 );
and \U$31536 ( \39781_40081 , \24490_24789 , \31877_32179_nG9bb4 );
or \U$31537 ( \39782_40082 , \39780_40080 , \39781_40081 );
xor \U$31538 ( \39783_40083 , \24489_24788 , \39782_40082 );
buf \U$31539 ( \39784_40084 , \39783_40083 );
buf \U$31541 ( \39785_40085 , \39784_40084 );
xor \U$31542 ( \39786_40086 , \39779_40079 , \39785_40085 );
buf \U$31543 ( \39787_40087 , \39786_40086 );
and \U$31544 ( \39788_40088 , \13431_13370 , \37674_37974_nG9b87 );
and \U$31545 ( \39789_40089 , \13068_13367 , \38037_38337_nG9b84 );
or \U$31546 ( \39790_40090 , \39788_40088 , \39789_40089 );
xor \U$31547 ( \39791_40091 , \13067_13366 , \39790_40090 );
buf \U$31548 ( \39792_40092 , \39791_40091 );
buf \U$31550 ( \39793_40093 , \39792_40092 );
xor \U$31551 ( \39794_40094 , \39787_40087 , \39793_40093 );
and \U$31552 ( \39795_40095 , \12183_12157 , \38363_38663_nG9b81 );
and \U$31553 ( \39796_40096 , \11855_12154 , \38668_38968_nG9b7e );
or \U$31554 ( \39797_40097 , \39795_40095 , \39796_40096 );
xor \U$31555 ( \39798_40098 , \11854_12153 , \39797_40097 );
buf \U$31556 ( \39799_40099 , \39798_40098 );
buf \U$31558 ( \39800_40100 , \39799_40099 );
xor \U$31559 ( \39801_40101 , \39794_40094 , \39800_40100 );
buf \U$31560 ( \39802_40102 , \39801_40101 );
and \U$31561 ( \39803_40103 , \39453_39753 , \39458_39758 );
and \U$31562 ( \39804_40104 , \39453_39753 , \39465_39765 );
and \U$31563 ( \39805_40105 , \39458_39758 , \39465_39765 );
or \U$31564 ( \39806_40106 , \39803_40103 , \39804_40104 , \39805_40105 );
buf \U$31565 ( \39807_40107 , \39806_40106 );
xor \U$31566 ( \39808_40108 , \39802_40102 , \39807_40107 );
and \U$31567 ( \39809_40109 , \39544_39844 , \39550_39850 );
buf \U$31568 ( \39810_40110 , \39809_40109 );
and \U$31569 ( \39811_40111 , \30670_29853 , \25561_25860_nG9bc9 );
and \U$31570 ( \39812_40112 , \29551_29850 , \26585_26887_nG9bc6 );
or \U$31571 ( \39813_40113 , \39811_40111 , \39812_40112 );
xor \U$31572 ( \39814_40114 , \29550_29849 , \39813_40113 );
buf \U$31573 ( \39815_40115 , \39814_40114 );
buf \U$31575 ( \39816_40116 , \39815_40115 );
xor \U$31576 ( \39817_40117 , \39810_40110 , \39816_40116 );
and \U$31577 ( \39818_40118 , \28946_28118 , \27114_27416_nG9bc3 );
and \U$31578 ( \39819_40119 , \27816_28115 , \28300_28602_nG9bc0 );
or \U$31579 ( \39820_40120 , \39818_40118 , \39819_40119 );
xor \U$31580 ( \39821_40121 , \27815_28114 , \39820_40120 );
buf \U$31581 ( \39822_40122 , \39821_40121 );
buf \U$31583 ( \39823_40123 , \39822_40122 );
xor \U$31584 ( \39824_40124 , \39817_40117 , \39823_40123 );
buf \U$31585 ( \39825_40125 , \39824_40124 );
and \U$31586 ( \39826_40126 , \16405_15940 , \36289_36589_nG9b93 );
and \U$31587 ( \39827_40127 , \15638_15937 , \36686_36986_nG9b90 );
or \U$31588 ( \39828_40128 , \39826_40126 , \39827_40127 );
xor \U$31589 ( \39829_40129 , \15637_15936 , \39828_40128 );
buf \U$31590 ( \39830_40130 , \39829_40129 );
buf \U$31592 ( \39831_40131 , \39830_40130 );
xor \U$31593 ( \39832_40132 , \39825_40125 , \39831_40131 );
and \U$31594 ( \39833_40133 , \10411_10707 , \39663_39963_nG9b75 );
and \U$31595 ( \39834_40134 , \39592_39892 , \39620_39920 );
and \U$31596 ( \39835_40135 , \39620_39920 , \39652_39952 );
and \U$31597 ( \39836_40136 , \39592_39892 , \39652_39952 );
or \U$31598 ( \39837_40137 , \39834_40134 , \39835_40135 , \39836_40136 );
and \U$31599 ( \39838_40138 , \39596_39896 , \39607_39907 );
and \U$31600 ( \39839_40139 , \39607_39907 , \39619_39919 );
and \U$31601 ( \39840_40140 , \39596_39896 , \39619_39919 );
or \U$31602 ( \39841_40141 , \39838_40138 , \39839_40139 , \39840_40140 );
and \U$31603 ( \39842_40142 , \39625_39925 , \39629_39929 );
and \U$31604 ( \39843_40143 , \39629_39929 , \39651_39951 );
and \U$31605 ( \39844_40144 , \39625_39925 , \39651_39951 );
or \U$31606 ( \39845_40145 , \39842_40142 , \39843_40143 , \39844_40144 );
xor \U$31607 ( \39846_40146 , \39841_40141 , \39845_40145 );
and \U$31608 ( \39847_40147 , \39634_39934 , \39638_39938 );
and \U$31609 ( \39848_40148 , \39638_39938 , \39650_39950 );
and \U$31610 ( \39849_40149 , \39634_39934 , \39650_39950 );
or \U$31611 ( \39850_40150 , \39847_40147 , \39848_40148 , \39849_40149 );
and \U$31612 ( \39851_40151 , \39600_39900 , \39604_39904 );
and \U$31613 ( \39852_40152 , \39604_39904 , \39606_39906 );
and \U$31614 ( \39853_40153 , \39600_39900 , \39606_39906 );
or \U$31615 ( \39854_40154 , \39851_40151 , \39852_40152 , \39853_40153 );
and \U$31616 ( \39855_40155 , \39640_39940 , \39644_39944 );
and \U$31617 ( \39856_40156 , \39644_39944 , \39649_39949 );
and \U$31618 ( \39857_40157 , \39640_39940 , \39649_39949 );
or \U$31619 ( \39858_40158 , \39855_40155 , \39856_40156 , \39857_40157 );
xor \U$31620 ( \39859_40159 , \39854_40154 , \39858_40158 );
and \U$31621 ( \39860_40160 , \32495_32794 , \23839_24138 );
not \U$31622 ( \39861_40161 , \39860_40160 );
xnor \U$31623 ( \39862_40162 , \39861_40161 , \23845_24144 );
not \U$31624 ( \39863_40163 , \39862_40162 );
xor \U$31625 ( \39864_40164 , \39859_40159 , \39863_40163 );
xor \U$31626 ( \39865_40165 , \39850_40150 , \39864_40164 );
and \U$31627 ( \39866_40166 , \39609_39909 , \39613_39913 );
and \U$31628 ( \39867_40167 , \39613_39913 , \39618_39918 );
and \U$31629 ( \39868_40168 , \39609_39909 , \39618_39918 );
or \U$31630 ( \39869_40169 , \39866_40166 , \39867_40167 , \39868_40168 );
and \U$31631 ( \39870_40170 , \30500_30802 , \25527_25826 );
and \U$31632 ( \39871_40171 , \31752_32054 , \24962_25264 );
nor \U$31633 ( \39872_40172 , \39870_40170 , \39871_40171 );
xnor \U$31634 ( \39873_40173 , \39872_40172 , \25474_25773 );
and \U$31635 ( \39874_40174 , \27011_27313 , \28768_29070 );
and \U$31636 ( \39875_40175 , \28232_28534 , \28224_28526 );
nor \U$31637 ( \39876_40176 , \39874_40174 , \39875_40175 );
xnor \U$31638 ( \39877_40177 , \39876_40176 , \28774_29076 );
xor \U$31639 ( \39878_40178 , \39873_40173 , \39877_40177 );
and \U$31640 ( \39879_40179 , \25516_25815 , \30521_30823 );
and \U$31641 ( \39880_40180 , \26527_26829 , \29944_30246 );
nor \U$31642 ( \39881_40181 , \39879_40179 , \39880_40180 );
xnor \U$31643 ( \39882_40182 , \39881_40181 , \30511_30813 );
xor \U$31644 ( \39883_40183 , \39878_40178 , \39882_40182 );
xor \U$31645 ( \39884_40184 , \39869_40169 , \39883_40183 );
and \U$31646 ( \39885_40185 , \28782_29084 , \27095_27397 );
and \U$31647 ( \39886_40186 , \29966_30268 , \26505_26807 );
nor \U$31648 ( \39887_40187 , \39885_40185 , \39886_40186 );
xnor \U$31649 ( \39888_40188 , \39887_40187 , \26993_27295 );
and \U$31650 ( \39889_40189 , \23900_24199 , \32555_32854 );
and \U$31651 ( \39890_40190 , \24970_25272 , \31765_32067 );
nor \U$31652 ( \39891_40191 , \39889_40189 , \39890_40190 );
xnor \U$31653 ( \39892_40192 , \39891_40191 , \32506_32805 );
xor \U$31654 ( \39893_40193 , \39888_40188 , \39892_40192 );
and \U$31655 ( \39894_40194 , \23315_23617 , \32503_32802 );
xor \U$31656 ( \39895_40195 , \39893_40193 , \39894_40194 );
xor \U$31657 ( \39896_40196 , \39884_40184 , \39895_40195 );
xor \U$31658 ( \39897_40197 , \39865_40165 , \39896_40196 );
xor \U$31659 ( \39898_40198 , \39846_40146 , \39897_40197 );
xor \U$31660 ( \39899_40199 , \39837_40137 , \39898_40198 );
and \U$31661 ( \39900_40200 , \39653_39953 , \39657_39957 );
and \U$31662 ( \39901_40201 , \39658_39958 , \39661_39961 );
or \U$31663 ( \39902_40202 , \39900_40200 , \39901_40201 );
xor \U$31664 ( \39903_40203 , \39899_40199 , \39902_40202 );
buf g9b72_GF_PartitionCandidate( \39904_40204_nG9b72 , \39903_40203 );
and \U$31665 ( \39905_40205 , \10402_10704 , \39904_40204_nG9b72 );
or \U$31666 ( \39906_40206 , \39833_40133 , \39905_40205 );
xor \U$31667 ( \39907_40207 , \10399_10703 , \39906_40206 );
buf \U$31668 ( \39908_40208 , \39907_40207 );
buf \U$31670 ( \39909_40209 , \39908_40208 );
xor \U$31671 ( \39910_40210 , \39832_40132 , \39909_40209 );
buf \U$31672 ( \39911_40211 , \39910_40210 );
xor \U$31673 ( \39912_40212 , \39808_40108 , \39911_40211 );
buf \U$31674 ( \39913_40213 , \39912_40212 );
and \U$31675 ( \39914_40214 , \39569_39869 , \39574_39874 );
and \U$31676 ( \39915_40215 , \39569_39869 , \39670_39970 );
and \U$31677 ( \39916_40216 , \39574_39874 , \39670_39970 );
or \U$31678 ( \39917_40217 , \39914_40214 , \39915_40215 , \39916_40216 );
buf \U$31679 ( \39918_40218 , \39917_40217 );
xor \U$31680 ( \39919_40219 , \39913_40213 , \39918_40218 );
and \U$31681 ( \39920_40220 , \39494_39794 , \39500_39800 );
and \U$31682 ( \39921_40221 , \39494_39794 , \39507_39807 );
and \U$31683 ( \39922_40222 , \39500_39800 , \39507_39807 );
or \U$31684 ( \39923_40223 , \39920_40220 , \39921_40221 , \39922_40222 );
buf \U$31685 ( \39924_40224 , \39923_40223 );
and \U$31686 ( \39925_40225 , \39523_39823 , \39529_39829 );
and \U$31687 ( \39926_40226 , \39523_39823 , \39536_39836 );
and \U$31688 ( \39927_40227 , \39529_39829 , \39536_39836 );
or \U$31689 ( \39928_40228 , \39925_40225 , \39926_40226 , \39927_40227 );
buf \U$31690 ( \39929_40229 , \39928_40228 );
xor \U$31691 ( \39930_40230 , \39924_40224 , \39929_40229 );
and \U$31692 ( \39931_40231 , \23495_23201 , \32589_32888_nG9bb1 );
and \U$31693 ( \39932_40232 , \22899_23198 , \32881_33181_nG9bae );
or \U$31694 ( \39933_40233 , \39931_40231 , \39932_40232 );
xor \U$31695 ( \39934_40234 , \22898_23197 , \39933_40233 );
buf \U$31696 ( \39935_40235 , \39934_40234 );
buf \U$31698 ( \39936_40236 , \39935_40235 );
and \U$31699 ( \39937_40237 , \21908_21658 , \33313_33613_nG9bab );
and \U$31700 ( \39938_40238 , \21356_21655 , \33741_34041_nG9ba8 );
or \U$31701 ( \39939_40239 , \39937_40237 , \39938_40238 );
xor \U$31702 ( \39940_40240 , \21355_21654 , \39939_40239 );
buf \U$31703 ( \39941_40241 , \39940_40240 );
buf \U$31705 ( \39942_40242 , \39941_40241 );
xor \U$31706 ( \39943_40243 , \39936_40236 , \39942_40242 );
and \U$31707 ( \39944_40244 , \20353_20155 , \33994_34294_nG9ba5 );
and \U$31708 ( \39945_40245 , \19853_20152 , \34343_34643_nG9ba2 );
or \U$31709 ( \39946_40246 , \39944_40244 , \39945_40245 );
xor \U$31710 ( \39947_40247 , \19852_20151 , \39946_40246 );
buf \U$31711 ( \39948_40248 , \39947_40247 );
buf \U$31713 ( \39949_40249 , \39948_40248 );
xor \U$31714 ( \39950_40250 , \39943_40243 , \39949_40249 );
buf \U$31715 ( \39951_40251 , \39950_40250 );
xor \U$31716 ( \39952_40252 , \39930_40230 , \39951_40251 );
buf \U$31717 ( \39953_40253 , \39952_40252 );
and \U$31718 ( \39954_40254 , \39552_39852 , \39558_39858 );
and \U$31719 ( \39955_40255 , \39552_39852 , \39565_39865 );
and \U$31720 ( \39956_40256 , \39558_39858 , \39565_39865 );
or \U$31721 ( \39957_40257 , \39954_40254 , \39955_40255 , \39956_40256 );
buf \U$31722 ( \39958_40258 , \39957_40257 );
and \U$31723 ( \39959_40259 , \14710_14631 , \36950_37250_nG9b8d );
and \U$31724 ( \39960_40260 , \14329_14628 , \37307_37607_nG9b8a );
or \U$31725 ( \39961_40261 , \39959_40259 , \39960_40260 );
xor \U$31726 ( \39962_40262 , \14328_14627 , \39961_40261 );
buf \U$31727 ( \39963_40263 , \39962_40262 );
buf \U$31729 ( \39964_40264 , \39963_40263 );
xor \U$31730 ( \39965_40265 , \39958_40258 , \39964_40264 );
and \U$31731 ( \39966_40266 , \10996_10421 , \39034_39334_nG9b7b );
and \U$31732 ( \39967_40267 , \10119_10418 , \39291_39591_nG9b78 );
or \U$31733 ( \39968_40268 , \39966_40266 , \39967_40267 );
xor \U$31734 ( \39969_40269 , \10118_10417 , \39968_40268 );
buf \U$31735 ( \39970_40270 , \39969_40269 );
buf \U$31737 ( \39971_40271 , \39970_40270 );
xor \U$31738 ( \39972_40272 , \39965_40265 , \39971_40271 );
buf \U$31739 ( \39973_40273 , \39972_40272 );
xor \U$31740 ( \39974_40274 , \39953_40253 , \39973_40273 );
and \U$31741 ( \39975_40275 , \39517_39817 , \39538_39838 );
and \U$31742 ( \39976_40276 , \39517_39817 , \39567_39867 );
and \U$31743 ( \39977_40277 , \39538_39838 , \39567_39867 );
or \U$31744 ( \39978_40278 , \39975_40275 , \39976_40276 , \39977_40277 );
buf \U$31745 ( \39979_40279 , \39978_40278 );
xor \U$31746 ( \39980_40280 , \39974_40274 , \39979_40279 );
buf \U$31747 ( \39981_40281 , \39980_40280 );
xor \U$31748 ( \39982_40282 , \39919_40219 , \39981_40281 );
buf \U$31749 ( \39983_40283 , \39982_40282 );
xor \U$31750 ( \39984_40284 , \39759_40059 , \39983_40283 );
and \U$31751 ( \39985_40285 , \39694_39994 , \39984_40284 );
and \U$31753 ( \39986_40286 , \39688_39988 , \39693_39993 );
or \U$31755 ( \39987_40287 , 1'b0 , \39986_40286 , 1'b0 );
xor \U$31756 ( \39988_40288 , \39985_40285 , \39987_40287 );
and \U$31758 ( \39989_40289 , \39681_39981 , \39687_39987 );
and \U$31759 ( \39990_40290 , \39683_39983 , \39687_39987 );
or \U$31760 ( \39991_40291 , 1'b0 , \39989_40289 , \39990_40290 );
xor \U$31761 ( \39992_40292 , \39988_40288 , \39991_40291 );
xor \U$31768 ( \39993_40293 , \39992_40292 , 1'b0 );
and \U$31769 ( \39994_40294 , \39753_40053 , \39758_40058 );
and \U$31770 ( \39995_40295 , \39753_40053 , \39983_40283 );
and \U$31771 ( \39996_40296 , \39758_40058 , \39983_40283 );
or \U$31772 ( \39997_40297 , \39994_40294 , \39995_40295 , \39996_40296 );
xor \U$31773 ( \39998_40298 , \39993_40293 , \39997_40297 );
and \U$31774 ( \39999_40299 , \39699_39999 , \39704_40004 );
and \U$31775 ( \40000_40300 , \39699_39999 , \39751_40051 );
and \U$31776 ( \40001_40301 , \39704_40004 , \39751_40051 );
or \U$31777 ( \40002_40302 , \39999_40299 , \40000_40300 , \40001_40301 );
buf \U$31778 ( \40003_40303 , \40002_40302 );
and \U$31779 ( \40004_40304 , \39721_40021 , \39726_40026 );
and \U$31780 ( \40005_40305 , \39721_40021 , \39747_40047 );
and \U$31781 ( \40006_40306 , \39726_40026 , \39747_40047 );
or \U$31782 ( \40007_40307 , \40004_40304 , \40005_40305 , \40006_40306 );
buf \U$31783 ( \40008_40308 , \40007_40307 );
and \U$31784 ( \40009_40309 , \39764_40064 , \39770_40070 );
buf \U$31785 ( \40010_40310 , \40009_40309 );
and \U$31786 ( \40011_40311 , \31989_31636 , \24996_25298_nG9bcc );
and \U$31787 ( \40012_40312 , \31334_31633 , \25561_25860_nG9bc9 );
or \U$31788 ( \40013_40313 , \40011_40311 , \40012_40312 );
xor \U$31789 ( \40014_40314 , \31333_31632 , \40013_40313 );
buf \U$31790 ( \40015_40315 , \40014_40314 );
buf \U$31792 ( \40016_40316 , \40015_40315 );
xor \U$31793 ( \40017_40317 , \40010_40310 , \40016_40316 );
and \U$31794 ( \40018_40318 , \27141_26431 , \30064_30366_nG9bba );
and \U$31795 ( \40019_40319 , \26129_26428 , \30638_30940_nG9bb7 );
or \U$31796 ( \40020_40320 , \40018_40318 , \40019_40319 );
xor \U$31797 ( \40021_40321 , \26128_26427 , \40020_40320 );
buf \U$31798 ( \40022_40322 , \40021_40321 );
buf \U$31800 ( \40023_40323 , \40022_40322 );
xor \U$31801 ( \40024_40324 , \40017_40317 , \40023_40323 );
buf \U$31802 ( \40025_40325 , \40024_40324 );
and \U$31803 ( \40026_40326 , \39936_40236 , \39942_40242 );
and \U$31804 ( \40027_40327 , \39936_40236 , \39949_40249 );
and \U$31805 ( \40028_40328 , \39942_40242 , \39949_40249 );
or \U$31806 ( \40029_40329 , \40026_40326 , \40027_40327 , \40028_40328 );
buf \U$31807 ( \40030_40330 , \40029_40329 );
xor \U$31808 ( \40031_40331 , \40025_40325 , \40030_40330 );
and \U$31809 ( \40032_40332 , \17437_17297 , \35872_36172_nG9b96 );
and \U$31810 ( \40033_40333 , \16995_17294 , \36289_36589_nG9b93 );
or \U$31811 ( \40034_40334 , \40032_40332 , \40033_40333 );
xor \U$31812 ( \40035_40335 , \16994_17293 , \40034_40334 );
buf \U$31813 ( \40036_40336 , \40035_40335 );
buf \U$31815 ( \40037_40337 , \40036_40336 );
xor \U$31816 ( \40038_40338 , \40031_40331 , \40037_40337 );
buf \U$31817 ( \40039_40339 , \40038_40338 );
xor \U$31818 ( \40040_40340 , \40008_40308 , \40039_40339 );
and \U$31819 ( \40041_40341 , \39924_40224 , \39929_40229 );
and \U$31820 ( \40042_40342 , \39924_40224 , \39951_40251 );
and \U$31821 ( \40043_40343 , \39929_40229 , \39951_40251 );
or \U$31822 ( \40044_40344 , \40041_40341 , \40042_40342 , \40043_40343 );
buf \U$31823 ( \40045_40345 , \40044_40344 );
xor \U$31824 ( \40046_40346 , \40040_40340 , \40045_40345 );
buf \U$31825 ( \40047_40347 , \40046_40346 );
and \U$31826 ( \40048_40348 , \39953_40253 , \39973_40273 );
and \U$31827 ( \40049_40349 , \39953_40253 , \39979_40279 );
and \U$31828 ( \40050_40350 , \39973_40273 , \39979_40279 );
or \U$31829 ( \40051_40351 , \40048_40348 , \40049_40349 , \40050_40350 );
buf \U$31830 ( \40052_40352 , \40051_40351 );
xor \U$31831 ( \40053_40353 , \40047_40347 , \40052_40352 );
and \U$31832 ( \40054_40354 , \39772_40072 , \39778_40078 );
and \U$31833 ( \40055_40355 , \39772_40072 , \39785_40085 );
and \U$31834 ( \40056_40356 , \39778_40078 , \39785_40085 );
or \U$31835 ( \40057_40357 , \40054_40354 , \40055_40355 , \40056_40356 );
buf \U$31836 ( \40058_40358 , \40057_40357 );
and \U$31837 ( \40059_40359 , \16405_15940 , \36686_36986_nG9b90 );
and \U$31838 ( \40060_40360 , \15638_15937 , \36950_37250_nG9b8d );
or \U$31839 ( \40061_40361 , \40059_40359 , \40060_40360 );
xor \U$31840 ( \40062_40362 , \15637_15936 , \40061_40361 );
buf \U$31841 ( \40063_40363 , \40062_40362 );
buf \U$31843 ( \40064_40364 , \40063_40363 );
xor \U$31844 ( \40065_40365 , \40058_40358 , \40064_40364 );
and \U$31845 ( \40066_40366 , \12183_12157 , \38668_38968_nG9b7e );
and \U$31846 ( \40067_40367 , \11855_12154 , \39034_39334_nG9b7b );
or \U$31847 ( \40068_40368 , \40066_40366 , \40067_40367 );
xor \U$31848 ( \40069_40369 , \11854_12153 , \40068_40368 );
buf \U$31849 ( \40070_40370 , \40069_40369 );
buf \U$31851 ( \40071_40371 , \40070_40370 );
xor \U$31852 ( \40072_40372 , \40065_40365 , \40071_40371 );
buf \U$31853 ( \40073_40373 , \40072_40372 );
and \U$31854 ( \40074_40374 , \21908_21658 , \33741_34041_nG9ba8 );
and \U$31855 ( \40075_40375 , \21356_21655 , \33994_34294_nG9ba5 );
or \U$31856 ( \40076_40376 , \40074_40374 , \40075_40375 );
xor \U$31857 ( \40077_40377 , \21355_21654 , \40076_40376 );
buf \U$31858 ( \40078_40378 , \40077_40377 );
buf \U$31860 ( \40079_40379 , \40078_40378 );
and \U$31861 ( \40080_40380 , \13431_13370 , \38037_38337_nG9b84 );
and \U$31862 ( \40081_40381 , \13068_13367 , \38363_38663_nG9b81 );
or \U$31863 ( \40082_40382 , \40080_40380 , \40081_40381 );
xor \U$31864 ( \40083_40383 , \13067_13366 , \40082_40382 );
buf \U$31865 ( \40084_40384 , \40083_40383 );
buf \U$31867 ( \40085_40385 , \40084_40384 );
xor \U$31868 ( \40086_40386 , \40079_40379 , \40085_40385 );
and \U$31869 ( \40087_40387 , \10411_10707 , \39904_40204_nG9b72 );
and \U$31870 ( \40088_40388 , \39850_40150 , \39864_40164 );
and \U$31871 ( \40089_40389 , \39864_40164 , \39896_40196 );
and \U$31872 ( \40090_40390 , \39850_40150 , \39896_40196 );
or \U$31873 ( \40091_40391 , \40088_40388 , \40089_40389 , \40090_40390 );
and \U$31874 ( \40092_40392 , \39888_40188 , \39892_40192 );
and \U$31875 ( \40093_40393 , \39892_40192 , \39894_40194 );
and \U$31876 ( \40094_40394 , \39888_40188 , \39894_40194 );
or \U$31877 ( \40095_40395 , \40092_40392 , \40093_40393 , \40094_40394 );
not \U$31878 ( \40096_40396 , \23845_24144 );
and \U$31879 ( \40097_40397 , \31752_32054 , \25527_25826 );
and \U$31880 ( \40098_40398 , \32495_32794 , \24962_25264 );
nor \U$31881 ( \40099_40399 , \40097_40397 , \40098_40398 );
xnor \U$31882 ( \40100_40400 , \40099_40399 , \25474_25773 );
xor \U$31883 ( \40101_40401 , \40096_40396 , \40100_40400 );
and \U$31884 ( \40102_40402 , \28232_28534 , \28768_29070 );
and \U$31885 ( \40103_40403 , \28782_29084 , \28224_28526 );
nor \U$31886 ( \40104_40404 , \40102_40402 , \40103_40403 );
xnor \U$31887 ( \40105_40405 , \40104_40404 , \28774_29076 );
xor \U$31888 ( \40106_40406 , \40101_40401 , \40105_40405 );
xor \U$31889 ( \40107_40407 , \40095_40395 , \40106_40406 );
and \U$31890 ( \40108_40408 , \29966_30268 , \27095_27397 );
and \U$31891 ( \40109_40409 , \30500_30802 , \26505_26807 );
nor \U$31892 ( \40110_40410 , \40108_40408 , \40109_40409 );
xnor \U$31893 ( \40111_40411 , \40110_40410 , \26993_27295 );
and \U$31894 ( \40112_40412 , \26527_26829 , \30521_30823 );
and \U$31895 ( \40113_40413 , \27011_27313 , \29944_30246 );
nor \U$31896 ( \40114_40414 , \40112_40412 , \40113_40413 );
xnor \U$31897 ( \40115_40415 , \40114_40414 , \30511_30813 );
xor \U$31898 ( \40116_40416 , \40111_40411 , \40115_40415 );
and \U$31899 ( \40117_40417 , \24970_25272 , \32555_32854 );
and \U$31900 ( \40118_40418 , \25516_25815 , \31765_32067 );
nor \U$31901 ( \40119_40419 , \40117_40417 , \40118_40418 );
xnor \U$31902 ( \40120_40420 , \40119_40419 , \32506_32805 );
xor \U$31903 ( \40121_40421 , \40116_40416 , \40120_40420 );
xor \U$31904 ( \40122_40422 , \40107_40407 , \40121_40421 );
xor \U$31905 ( \40123_40423 , \40091_40391 , \40122_40422 );
and \U$31906 ( \40124_40424 , \39854_40154 , \39858_40158 );
and \U$31907 ( \40125_40425 , \39858_40158 , \39863_40163 );
and \U$31908 ( \40126_40426 , \39854_40154 , \39863_40163 );
or \U$31909 ( \40127_40427 , \40124_40424 , \40125_40425 , \40126_40426 );
and \U$31910 ( \40128_40428 , \39869_40169 , \39883_40183 );
and \U$31911 ( \40129_40429 , \39883_40183 , \39895_40195 );
and \U$31912 ( \40130_40430 , \39869_40169 , \39895_40195 );
or \U$31913 ( \40131_40431 , \40128_40428 , \40129_40429 , \40130_40430 );
xor \U$31914 ( \40132_40432 , \40127_40427 , \40131_40431 );
and \U$31915 ( \40133_40433 , \39873_40173 , \39877_40177 );
and \U$31916 ( \40134_40434 , \39877_40177 , \39882_40182 );
and \U$31917 ( \40135_40435 , \39873_40173 , \39882_40182 );
or \U$31918 ( \40136_40436 , \40133_40433 , \40134_40434 , \40135_40435 );
buf \U$31919 ( \40137_40437 , \39862_40162 );
xor \U$31920 ( \40138_40438 , \40136_40436 , \40137_40437 );
and \U$31921 ( \40139_40439 , \23900_24199 , \32503_32802 );
xor \U$31922 ( \40140_40440 , \40138_40438 , \40139_40439 );
xor \U$31923 ( \40141_40441 , \40132_40432 , \40140_40440 );
xor \U$31924 ( \40142_40442 , \40123_40423 , \40141_40441 );
and \U$31925 ( \40143_40443 , \39841_40141 , \39845_40145 );
and \U$31926 ( \40144_40444 , \39845_40145 , \39897_40197 );
and \U$31927 ( \40145_40445 , \39841_40141 , \39897_40197 );
or \U$31928 ( \40146_40446 , \40143_40443 , \40144_40444 , \40145_40445 );
xor \U$31929 ( \40147_40447 , \40142_40442 , \40146_40446 );
and \U$31930 ( \40148_40448 , \39837_40137 , \39898_40198 );
and \U$31931 ( \40149_40449 , \39899_40199 , \39902_40202 );
or \U$31932 ( \40150_40450 , \40148_40448 , \40149_40449 );
xor \U$31933 ( \40151_40451 , \40147_40447 , \40150_40450 );
buf g9b6f_GF_PartitionCandidate( \40152_40452_nG9b6f , \40151_40451 );
and \U$31934 ( \40153_40453 , \10402_10704 , \40152_40452_nG9b6f );
or \U$31935 ( \40154_40454 , \40087_40387 , \40153_40453 );
xor \U$31936 ( \40155_40455 , \10399_10703 , \40154_40454 );
buf \U$31937 ( \40156_40456 , \40155_40455 );
buf \U$31939 ( \40157_40457 , \40156_40456 );
xor \U$31940 ( \40158_40458 , \40086_40386 , \40157_40457 );
buf \U$31941 ( \40159_40459 , \40158_40458 );
xor \U$31942 ( \40160_40460 , \40073_40373 , \40159_40459 );
and \U$31943 ( \40161_40461 , \39810_40110 , \39816_40116 );
and \U$31944 ( \40162_40462 , \39810_40110 , \39823_40123 );
and \U$31945 ( \40163_40463 , \39816_40116 , \39823_40123 );
or \U$31946 ( \40164_40464 , \40161_40461 , \40162_40462 , \40163_40463 );
buf \U$31947 ( \40165_40465 , \40164_40464 );
and \U$31948 ( \40166_40466 , \14710_14631 , \37307_37607_nG9b8a );
and \U$31949 ( \40167_40467 , \14329_14628 , \37674_37974_nG9b87 );
or \U$31950 ( \40168_40468 , \40166_40466 , \40167_40467 );
xor \U$31951 ( \40169_40469 , \14328_14627 , \40168_40468 );
buf \U$31952 ( \40170_40470 , \40169_40469 );
buf \U$31954 ( \40171_40471 , \40170_40470 );
xor \U$31955 ( \40172_40472 , \40165_40465 , \40171_40471 );
and \U$31956 ( \40173_40473 , \10996_10421 , \39291_39591_nG9b78 );
and \U$31957 ( \40174_40474 , \10119_10418 , \39663_39963_nG9b75 );
or \U$31958 ( \40175_40475 , \40173_40473 , \40174_40474 );
xor \U$31959 ( \40176_40476 , \10118_10417 , \40175_40475 );
buf \U$31960 ( \40177_40477 , \40176_40476 );
buf \U$31962 ( \40178_40478 , \40177_40477 );
xor \U$31963 ( \40179_40479 , \40172_40472 , \40178_40478 );
buf \U$31964 ( \40180_40480 , \40179_40479 );
xor \U$31965 ( \40181_40481 , \40160_40460 , \40180_40480 );
buf \U$31966 ( \40182_40482 , \40181_40481 );
xor \U$31967 ( \40183_40483 , \40053_40353 , \40182_40482 );
buf \U$31968 ( \40184_40484 , \40183_40483 );
xor \U$31969 ( \40185_40485 , \40003_40303 , \40184_40484 );
and \U$31970 ( \40186_40486 , \39913_40213 , \39918_40218 );
and \U$31971 ( \40187_40487 , \39913_40213 , \39981_40281 );
and \U$31972 ( \40188_40488 , \39918_40218 , \39981_40281 );
or \U$31973 ( \40189_40489 , \40186_40486 , \40187_40487 , \40188_40488 );
buf \U$31974 ( \40190_40490 , \40189_40489 );
and \U$31975 ( \40191_40491 , \39802_40102 , \39807_40107 );
and \U$31976 ( \40192_40492 , \39802_40102 , \39911_40211 );
and \U$31977 ( \40193_40493 , \39807_40107 , \39911_40211 );
or \U$31978 ( \40194_40494 , \40191_40491 , \40192_40492 , \40193_40493 );
buf \U$31979 ( \40195_40495 , \40194_40494 );
and \U$31980 ( \40196_40496 , \39787_40087 , \39793_40093 );
and \U$31981 ( \40197_40497 , \39787_40087 , \39800_40100 );
and \U$31982 ( \40198_40498 , \39793_40093 , \39800_40100 );
or \U$31983 ( \40199_40499 , \40196_40496 , \40197_40497 , \40198_40498 );
buf \U$31984 ( \40200_40500 , \40199_40499 );
and \U$31985 ( \40201_40501 , \39825_40125 , \39831_40131 );
and \U$31986 ( \40202_40502 , \39825_40125 , \39909_40209 );
and \U$31987 ( \40203_40503 , \39831_40131 , \39909_40209 );
or \U$31988 ( \40204_40504 , \40201_40501 , \40202_40502 , \40203_40503 );
buf \U$31989 ( \40205_40505 , \40204_40504 );
xor \U$31990 ( \40206_40506 , \40200_40500 , \40205_40505 );
and \U$31991 ( \40207_40507 , \23495_23201 , \32881_33181_nG9bae );
and \U$31992 ( \40208_40508 , \22899_23198 , \33313_33613_nG9bab );
or \U$31993 ( \40209_40509 , \40207_40507 , \40208_40508 );
xor \U$31994 ( \40210_40510 , \22898_23197 , \40209_40509 );
buf \U$31995 ( \40211_40511 , \40210_40510 );
buf \U$31997 ( \40212_40512 , \40211_40511 );
and \U$31998 ( \40213_40513 , \20353_20155 , \34343_34643_nG9ba2 );
and \U$31999 ( \40214_40514 , \19853_20152 , \34794_35094_nG9b9f );
or \U$32000 ( \40215_40515 , \40213_40513 , \40214_40514 );
xor \U$32001 ( \40216_40516 , \19852_20151 , \40215_40515 );
buf \U$32002 ( \40217_40517 , \40216_40516 );
buf \U$32004 ( \40218_40518 , \40217_40517 );
xor \U$32005 ( \40219_40519 , \40212_40512 , \40218_40518 );
and \U$32006 ( \40220_40520 , \18908_18702 , \35270_35570_nG9b9c );
and \U$32007 ( \40221_40521 , \18400_18699 , \35501_35801_nG9b99 );
or \U$32008 ( \40222_40522 , \40220_40520 , \40221_40521 );
xor \U$32009 ( \40223_40523 , \18399_18698 , \40222_40522 );
buf \U$32010 ( \40224_40524 , \40223_40523 );
buf \U$32012 ( \40225_40525 , \40224_40524 );
xor \U$32013 ( \40226_40526 , \40219_40519 , \40225_40525 );
buf \U$32014 ( \40227_40527 , \40226_40526 );
xor \U$32015 ( \40228_40528 , \40206_40506 , \40227_40527 );
buf \U$32016 ( \40229_40529 , \40228_40528 );
xor \U$32017 ( \40230_40530 , \40195_40495 , \40229_40529 );
and \U$32018 ( \40231_40531 , \39958_40258 , \39964_40264 );
and \U$32019 ( \40232_40532 , \39958_40258 , \39971_40271 );
and \U$32020 ( \40233_40533 , \39964_40264 , \39971_40271 );
or \U$32021 ( \40234_40534 , \40231_40531 , \40232_40532 , \40233_40533 );
buf \U$32022 ( \40235_40535 , \40234_40534 );
and \U$32023 ( \40236_40536 , \39732_40032 , \39738_40038 );
and \U$32024 ( \40237_40537 , \39732_40032 , \39745_40045 );
and \U$32025 ( \40238_40538 , \39738_40038 , \39745_40045 );
or \U$32026 ( \40239_40539 , \40236_40536 , \40237_40537 , \40238_40538 );
buf \U$32027 ( \40240_40540 , \40239_40539 );
xor \U$32028 ( \40241_40541 , \40235_40535 , \40240_40540 );
and \U$32030 ( \40242_40542 , \32617_32916 , \23927_24226_nG9bcf );
or \U$32031 ( \40243_40543 , 1'b0 , \40242_40542 );
xor \U$32032 ( \40244_40544 , 1'b0 , \40243_40543 );
buf \U$32033 ( \40245_40545 , \40244_40544 );
buf \U$32035 ( \40246_40546 , \40245_40545 );
and \U$32036 ( \40247_40547 , \30670_29853 , \26585_26887_nG9bc6 );
and \U$32037 ( \40248_40548 , \29551_29850 , \27114_27416_nG9bc3 );
or \U$32038 ( \40249_40549 , \40247_40547 , \40248_40548 );
xor \U$32039 ( \40250_40550 , \29550_29849 , \40249_40549 );
buf \U$32040 ( \40251_40551 , \40250_40550 );
buf \U$32042 ( \40252_40552 , \40251_40551 );
xor \U$32043 ( \40253_40553 , \40246_40546 , \40252_40552 );
buf \U$32044 ( \40254_40554 , \40253_40553 );
and \U$32045 ( \40255_40555 , \28946_28118 , \28300_28602_nG9bc0 );
and \U$32046 ( \40256_40556 , \27816_28115 , \28877_29179_nG9bbd );
or \U$32047 ( \40257_40557 , \40255_40555 , \40256_40556 );
xor \U$32048 ( \40258_40558 , \27815_28114 , \40257_40557 );
buf \U$32049 ( \40259_40559 , \40258_40558 );
buf \U$32051 ( \40260_40560 , \40259_40559 );
xor \U$32052 ( \40261_40561 , \40254_40554 , \40260_40560 );
and \U$32053 ( \40262_40562 , \25044_24792 , \31877_32179_nG9bb4 );
and \U$32054 ( \40263_40563 , \24490_24789 , \32589_32888_nG9bb1 );
or \U$32055 ( \40264_40564 , \40262_40562 , \40263_40563 );
xor \U$32056 ( \40265_40565 , \24489_24788 , \40264_40564 );
buf \U$32057 ( \40266_40566 , \40265_40565 );
buf \U$32059 ( \40267_40567 , \40266_40566 );
xor \U$32060 ( \40268_40568 , \40261_40561 , \40267_40567 );
buf \U$32061 ( \40269_40569 , \40268_40568 );
xor \U$32062 ( \40270_40570 , \40241_40541 , \40269_40569 );
buf \U$32063 ( \40271_40571 , \40270_40570 );
xor \U$32064 ( \40272_40572 , \40230_40530 , \40271_40571 );
buf \U$32065 ( \40273_40573 , \40272_40572 );
xor \U$32066 ( \40274_40574 , \40190_40490 , \40273_40573 );
and \U$32067 ( \40275_40575 , \39710_40010 , \39715_40015 );
and \U$32068 ( \40276_40576 , \39710_40010 , \39749_40049 );
and \U$32069 ( \40277_40577 , \39715_40015 , \39749_40049 );
or \U$32070 ( \40278_40578 , \40275_40575 , \40276_40576 , \40277_40577 );
buf \U$32071 ( \40279_40579 , \40278_40578 );
xor \U$32072 ( \40280_40580 , \40274_40574 , \40279_40579 );
buf \U$32073 ( \40281_40581 , \40280_40580 );
xor \U$32074 ( \40282_40582 , \40185_40485 , \40281_40581 );
and \U$32075 ( \40283_40583 , \39998_40298 , \40282_40582 );
and \U$32077 ( \40284_40584 , \39992_40292 , \39997_40297 );
or \U$32079 ( \40285_40585 , 1'b0 , \40284_40584 , 1'b0 );
xor \U$32080 ( \40286_40586 , \40283_40583 , \40285_40585 );
and \U$32082 ( \40287_40587 , \39985_40285 , \39991_40291 );
and \U$32083 ( \40288_40588 , \39987_40287 , \39991_40291 );
or \U$32084 ( \40289_40589 , 1'b0 , \40287_40587 , \40288_40588 );
xor \U$32085 ( \40290_40590 , \40286_40586 , \40289_40589 );
xor \U$32092 ( \40291_40591 , \40290_40590 , 1'b0 );
and \U$32093 ( \40292_40592 , \40003_40303 , \40184_40484 );
and \U$32094 ( \40293_40593 , \40003_40303 , \40281_40581 );
and \U$32095 ( \40294_40594 , \40184_40484 , \40281_40581 );
or \U$32096 ( \40295_40595 , \40292_40592 , \40293_40593 , \40294_40594 );
xor \U$32097 ( \40296_40596 , \40291_40591 , \40295_40595 );
and \U$32098 ( \40297_40597 , \40047_40347 , \40052_40352 );
and \U$32099 ( \40298_40598 , \40047_40347 , \40182_40482 );
and \U$32100 ( \40299_40599 , \40052_40352 , \40182_40482 );
or \U$32101 ( \40300_40600 , \40297_40597 , \40298_40598 , \40299_40599 );
buf \U$32102 ( \40301_40601 , \40300_40600 );
and \U$32103 ( \40302_40602 , \40073_40373 , \40159_40459 );
and \U$32104 ( \40303_40603 , \40073_40373 , \40180_40480 );
and \U$32105 ( \40304_40604 , \40159_40459 , \40180_40480 );
or \U$32106 ( \40305_40605 , \40302_40602 , \40303_40603 , \40304_40604 );
buf \U$32107 ( \40306_40606 , \40305_40605 );
and \U$32108 ( \40307_40607 , \17437_17297 , \36289_36589_nG9b93 );
and \U$32109 ( \40308_40608 , \16995_17294 , \36686_36986_nG9b90 );
or \U$32110 ( \40309_40609 , \40307_40607 , \40308_40608 );
xor \U$32111 ( \40310_40610 , \16994_17293 , \40309_40609 );
buf \U$32112 ( \40311_40611 , \40310_40610 );
buf \U$32114 ( \40312_40612 , \40311_40611 );
and \U$32115 ( \40313_40613 , \16405_15940 , \36950_37250_nG9b8d );
and \U$32116 ( \40314_40614 , \15638_15937 , \37307_37607_nG9b8a );
or \U$32117 ( \40315_40615 , \40313_40613 , \40314_40614 );
xor \U$32118 ( \40316_40616 , \15637_15936 , \40315_40615 );
buf \U$32119 ( \40317_40617 , \40316_40616 );
buf \U$32121 ( \40318_40618 , \40317_40617 );
xor \U$32122 ( \40319_40619 , \40312_40612 , \40318_40618 );
and \U$32123 ( \40320_40620 , \12183_12157 , \39034_39334_nG9b7b );
and \U$32124 ( \40321_40621 , \11855_12154 , \39291_39591_nG9b78 );
or \U$32125 ( \40322_40622 , \40320_40620 , \40321_40621 );
xor \U$32126 ( \40323_40623 , \11854_12153 , \40322_40622 );
buf \U$32127 ( \40324_40624 , \40323_40623 );
buf \U$32129 ( \40325_40625 , \40324_40624 );
xor \U$32130 ( \40326_40626 , \40319_40619 , \40325_40625 );
buf \U$32131 ( \40327_40627 , \40326_40626 );
and \U$32132 ( \40328_40628 , \23495_23201 , \33313_33613_nG9bab );
and \U$32133 ( \40329_40629 , \22899_23198 , \33741_34041_nG9ba8 );
or \U$32134 ( \40330_40630 , \40328_40628 , \40329_40629 );
xor \U$32135 ( \40331_40631 , \22898_23197 , \40330_40630 );
buf \U$32136 ( \40332_40632 , \40331_40631 );
buf \U$32138 ( \40333_40633 , \40332_40632 );
and \U$32139 ( \40334_40634 , \20353_20155 , \34794_35094_nG9b9f );
and \U$32140 ( \40335_40635 , \19853_20152 , \35270_35570_nG9b9c );
or \U$32141 ( \40336_40636 , \40334_40634 , \40335_40635 );
xor \U$32142 ( \40337_40637 , \19852_20151 , \40336_40636 );
buf \U$32143 ( \40338_40638 , \40337_40637 );
buf \U$32145 ( \40339_40639 , \40338_40638 );
xor \U$32146 ( \40340_40640 , \40333_40633 , \40339_40639 );
and \U$32147 ( \40341_40641 , \18908_18702 , \35501_35801_nG9b99 );
and \U$32148 ( \40342_40642 , \18400_18699 , \35872_36172_nG9b96 );
or \U$32149 ( \40343_40643 , \40341_40641 , \40342_40642 );
xor \U$32150 ( \40344_40644 , \18399_18698 , \40343_40643 );
buf \U$32151 ( \40345_40645 , \40344_40644 );
buf \U$32153 ( \40346_40646 , \40345_40645 );
xor \U$32154 ( \40347_40647 , \40340_40640 , \40346_40646 );
buf \U$32155 ( \40348_40648 , \40347_40647 );
xor \U$32156 ( \40349_40649 , \40327_40627 , \40348_40648 );
and \U$32157 ( \40350_40650 , \40058_40358 , \40064_40364 );
and \U$32158 ( \40351_40651 , \40058_40358 , \40071_40371 );
and \U$32159 ( \40352_40652 , \40064_40364 , \40071_40371 );
or \U$32160 ( \40353_40653 , \40350_40650 , \40351_40651 , \40352_40652 );
buf \U$32161 ( \40354_40654 , \40353_40653 );
xor \U$32162 ( \40355_40655 , \40349_40649 , \40354_40654 );
buf \U$32163 ( \40356_40656 , \40355_40655 );
xor \U$32164 ( \40357_40657 , \40306_40606 , \40356_40656 );
and \U$32165 ( \40358_40658 , \40200_40500 , \40205_40505 );
and \U$32166 ( \40359_40659 , \40200_40500 , \40227_40527 );
and \U$32167 ( \40360_40660 , \40205_40505 , \40227_40527 );
or \U$32168 ( \40361_40661 , \40358_40658 , \40359_40659 , \40360_40660 );
buf \U$32169 ( \40362_40662 , \40361_40661 );
xor \U$32170 ( \40363_40663 , \40357_40657 , \40362_40662 );
buf \U$32171 ( \40364_40664 , \40363_40663 );
xor \U$32172 ( \40365_40665 , \40301_40601 , \40364_40664 );
and \U$32173 ( \40366_40666 , \40079_40379 , \40085_40385 );
and \U$32174 ( \40367_40667 , \40079_40379 , \40157_40457 );
and \U$32175 ( \40368_40668 , \40085_40385 , \40157_40457 );
or \U$32176 ( \40369_40669 , \40366_40666 , \40367_40667 , \40368_40668 );
buf \U$32177 ( \40370_40670 , \40369_40669 );
and \U$32178 ( \40371_40671 , \40165_40465 , \40171_40471 );
and \U$32179 ( \40372_40672 , \40165_40465 , \40178_40478 );
and \U$32180 ( \40373_40673 , \40171_40471 , \40178_40478 );
or \U$32181 ( \40374_40674 , \40371_40671 , \40372_40672 , \40373_40673 );
buf \U$32182 ( \40375_40675 , \40374_40674 );
xor \U$32183 ( \40376_40676 , \40370_40670 , \40375_40675 );
and \U$32185 ( \40377_40677 , \32617_32916 , \24996_25298_nG9bcc );
or \U$32186 ( \40378_40678 , 1'b0 , \40377_40677 );
xor \U$32187 ( \40379_40679 , 1'b0 , \40378_40678 );
buf \U$32188 ( \40380_40680 , \40379_40679 );
buf \U$32190 ( \40381_40681 , \40380_40680 );
and \U$32191 ( \40382_40682 , \30670_29853 , \27114_27416_nG9bc3 );
and \U$32192 ( \40383_40683 , \29551_29850 , \28300_28602_nG9bc0 );
or \U$32193 ( \40384_40684 , \40382_40682 , \40383_40683 );
xor \U$32194 ( \40385_40685 , \29550_29849 , \40384_40684 );
buf \U$32195 ( \40386_40686 , \40385_40685 );
buf \U$32197 ( \40387_40687 , \40386_40686 );
xor \U$32198 ( \40388_40688 , \40381_40681 , \40387_40687 );
buf \U$32199 ( \40389_40689 , \40388_40688 );
and \U$32200 ( \40390_40690 , \40246_40546 , \40252_40552 );
buf \U$32201 ( \40391_40691 , \40390_40690 );
xor \U$32202 ( \40392_40692 , \40389_40689 , \40391_40691 );
and \U$32203 ( \40393_40693 , \25044_24792 , \32589_32888_nG9bb1 );
and \U$32204 ( \40394_40694 , \24490_24789 , \32881_33181_nG9bae );
or \U$32205 ( \40395_40695 , \40393_40693 , \40394_40694 );
xor \U$32206 ( \40396_40696 , \24489_24788 , \40395_40695 );
buf \U$32207 ( \40397_40697 , \40396_40696 );
buf \U$32209 ( \40398_40698 , \40397_40697 );
xor \U$32210 ( \40399_40699 , \40392_40692 , \40398_40698 );
buf \U$32211 ( \40400_40700 , \40399_40699 );
xor \U$32212 ( \40401_40701 , \40376_40676 , \40400_40700 );
buf \U$32213 ( \40402_40702 , \40401_40701 );
and \U$32214 ( \40403_40703 , \40235_40535 , \40240_40540 );
and \U$32215 ( \40404_40704 , \40235_40535 , \40269_40569 );
and \U$32216 ( \40405_40705 , \40240_40540 , \40269_40569 );
or \U$32217 ( \40406_40706 , \40403_40703 , \40404_40704 , \40405_40705 );
buf \U$32218 ( \40407_40707 , \40406_40706 );
xor \U$32219 ( \40408_40708 , \40402_40702 , \40407_40707 );
and \U$32220 ( \40409_40709 , \40212_40512 , \40218_40518 );
and \U$32221 ( \40410_40710 , \40212_40512 , \40225_40525 );
and \U$32222 ( \40411_40711 , \40218_40518 , \40225_40525 );
or \U$32223 ( \40412_40712 , \40409_40709 , \40410_40710 , \40411_40711 );
buf \U$32224 ( \40413_40713 , \40412_40712 );
and \U$32225 ( \40414_40714 , \40254_40554 , \40260_40560 );
and \U$32226 ( \40415_40715 , \40254_40554 , \40267_40567 );
and \U$32227 ( \40416_40716 , \40260_40560 , \40267_40567 );
or \U$32228 ( \40417_40717 , \40414_40714 , \40415_40715 , \40416_40716 );
buf \U$32229 ( \40418_40718 , \40417_40717 );
xor \U$32230 ( \40419_40719 , \40413_40713 , \40418_40718 );
and \U$32231 ( \40420_40720 , \31989_31636 , \25561_25860_nG9bc9 );
and \U$32232 ( \40421_40721 , \31334_31633 , \26585_26887_nG9bc6 );
or \U$32233 ( \40422_40722 , \40420_40720 , \40421_40721 );
xor \U$32234 ( \40423_40723 , \31333_31632 , \40422_40722 );
buf \U$32235 ( \40424_40724 , \40423_40723 );
buf \U$32237 ( \40425_40725 , \40424_40724 );
and \U$32238 ( \40426_40726 , \28946_28118 , \28877_29179_nG9bbd );
and \U$32239 ( \40427_40727 , \27816_28115 , \30064_30366_nG9bba );
or \U$32240 ( \40428_40728 , \40426_40726 , \40427_40727 );
xor \U$32241 ( \40429_40729 , \27815_28114 , \40428_40728 );
buf \U$32242 ( \40430_40730 , \40429_40729 );
buf \U$32244 ( \40431_40731 , \40430_40730 );
xor \U$32245 ( \40432_40732 , \40425_40725 , \40431_40731 );
and \U$32246 ( \40433_40733 , \27141_26431 , \30638_30940_nG9bb7 );
and \U$32247 ( \40434_40734 , \26129_26428 , \31877_32179_nG9bb4 );
or \U$32248 ( \40435_40735 , \40433_40733 , \40434_40734 );
xor \U$32249 ( \40436_40736 , \26128_26427 , \40435_40735 );
buf \U$32250 ( \40437_40737 , \40436_40736 );
buf \U$32252 ( \40438_40738 , \40437_40737 );
xor \U$32253 ( \40439_40739 , \40432_40732 , \40438_40738 );
buf \U$32254 ( \40440_40740 , \40439_40739 );
xor \U$32255 ( \40441_40741 , \40419_40719 , \40440_40740 );
buf \U$32256 ( \40442_40742 , \40441_40741 );
xor \U$32257 ( \40443_40743 , \40408_40708 , \40442_40742 );
buf \U$32258 ( \40444_40744 , \40443_40743 );
xor \U$32259 ( \40445_40745 , \40365_40665 , \40444_40744 );
buf \U$32260 ( \40446_40746 , \40445_40745 );
and \U$32261 ( \40447_40747 , \40190_40490 , \40273_40573 );
and \U$32262 ( \40448_40748 , \40190_40490 , \40279_40579 );
and \U$32263 ( \40449_40749 , \40273_40573 , \40279_40579 );
or \U$32264 ( \40450_40750 , \40447_40747 , \40448_40748 , \40449_40749 );
buf \U$32265 ( \40451_40751 , \40450_40750 );
xor \U$32266 ( \40452_40752 , \40446_40746 , \40451_40751 );
and \U$32267 ( \40453_40753 , \40195_40495 , \40229_40529 );
and \U$32268 ( \40454_40754 , \40195_40495 , \40271_40571 );
and \U$32269 ( \40455_40755 , \40229_40529 , \40271_40571 );
or \U$32270 ( \40456_40756 , \40453_40753 , \40454_40754 , \40455_40755 );
buf \U$32271 ( \40457_40757 , \40456_40756 );
and \U$32272 ( \40458_40758 , \40008_40308 , \40039_40339 );
and \U$32273 ( \40459_40759 , \40008_40308 , \40045_40345 );
and \U$32274 ( \40460_40760 , \40039_40339 , \40045_40345 );
or \U$32275 ( \40461_40761 , \40458_40758 , \40459_40759 , \40460_40760 );
buf \U$32276 ( \40462_40762 , \40461_40761 );
xor \U$32277 ( \40463_40763 , \40457_40757 , \40462_40762 );
and \U$32278 ( \40464_40764 , \40025_40325 , \40030_40330 );
and \U$32279 ( \40465_40765 , \40025_40325 , \40037_40337 );
and \U$32280 ( \40466_40766 , \40030_40330 , \40037_40337 );
or \U$32281 ( \40467_40767 , \40464_40764 , \40465_40765 , \40466_40766 );
buf \U$32282 ( \40468_40768 , \40467_40767 );
and \U$32283 ( \40469_40769 , \21908_21658 , \33994_34294_nG9ba5 );
and \U$32284 ( \40470_40770 , \21356_21655 , \34343_34643_nG9ba2 );
or \U$32285 ( \40471_40771 , \40469_40769 , \40470_40770 );
xor \U$32286 ( \40472_40772 , \21355_21654 , \40471_40771 );
buf \U$32287 ( \40473_40773 , \40472_40772 );
buf \U$32289 ( \40474_40774 , \40473_40773 );
and \U$32290 ( \40475_40775 , \13431_13370 , \38363_38663_nG9b81 );
and \U$32291 ( \40476_40776 , \13068_13367 , \38668_38968_nG9b7e );
or \U$32292 ( \40477_40777 , \40475_40775 , \40476_40776 );
xor \U$32293 ( \40478_40778 , \13067_13366 , \40477_40777 );
buf \U$32294 ( \40479_40779 , \40478_40778 );
buf \U$32296 ( \40480_40780 , \40479_40779 );
xor \U$32297 ( \40481_40781 , \40474_40774 , \40480_40780 );
and \U$32298 ( \40482_40782 , \10411_10707 , \40152_40452_nG9b6f );
and \U$32299 ( \40483_40783 , \40127_40427 , \40131_40431 );
and \U$32300 ( \40484_40784 , \40131_40431 , \40140_40440 );
and \U$32301 ( \40485_40785 , \40127_40427 , \40140_40440 );
or \U$32302 ( \40486_40786 , \40483_40783 , \40484_40784 , \40485_40785 );
and \U$32303 ( \40487_40787 , \40096_40396 , \40100_40400 );
and \U$32304 ( \40488_40788 , \40100_40400 , \40105_40405 );
and \U$32305 ( \40489_40789 , \40096_40396 , \40105_40405 );
or \U$32306 ( \40490_40790 , \40487_40787 , \40488_40788 , \40489_40789 );
and \U$32307 ( \40491_40791 , \40111_40411 , \40115_40415 );
and \U$32308 ( \40492_40792 , \40115_40415 , \40120_40420 );
and \U$32309 ( \40493_40793 , \40111_40411 , \40120_40420 );
or \U$32310 ( \40494_40794 , \40491_40791 , \40492_40792 , \40493_40793 );
xor \U$32311 ( \40495_40795 , \40490_40790 , \40494_40794 );
and \U$32312 ( \40496_40796 , \32495_32794 , \25527_25826 );
not \U$32313 ( \40497_40797 , \40496_40796 );
xnor \U$32314 ( \40498_40798 , \40497_40797 , \25474_25773 );
and \U$32315 ( \40499_40799 , \27011_27313 , \30521_30823 );
and \U$32316 ( \40500_40800 , \28232_28534 , \29944_30246 );
nor \U$32317 ( \40501_40801 , \40499_40799 , \40500_40800 );
xnor \U$32318 ( \40502_40802 , \40501_40801 , \30511_30813 );
xor \U$32319 ( \40503_40803 , \40498_40798 , \40502_40802 );
and \U$32320 ( \40504_40804 , \25516_25815 , \32555_32854 );
and \U$32321 ( \40505_40805 , \26527_26829 , \31765_32067 );
nor \U$32322 ( \40506_40806 , \40504_40804 , \40505_40805 );
xnor \U$32323 ( \40507_40807 , \40506_40806 , \32506_32805 );
xor \U$32324 ( \40508_40808 , \40503_40803 , \40507_40807 );
xor \U$32325 ( \40509_40809 , \40495_40795 , \40508_40808 );
xor \U$32326 ( \40510_40810 , \40486_40786 , \40509_40809 );
and \U$32327 ( \40511_40811 , \40136_40436 , \40137_40437 );
and \U$32328 ( \40512_40812 , \40137_40437 , \40139_40439 );
and \U$32329 ( \40513_40813 , \40136_40436 , \40139_40439 );
or \U$32330 ( \40514_40814 , \40511_40811 , \40512_40812 , \40513_40813 );
and \U$32331 ( \40515_40815 , \40095_40395 , \40106_40406 );
and \U$32332 ( \40516_40816 , \40106_40406 , \40121_40421 );
and \U$32333 ( \40517_40817 , \40095_40395 , \40121_40421 );
or \U$32334 ( \40518_40818 , \40515_40815 , \40516_40816 , \40517_40817 );
xor \U$32335 ( \40519_40819 , \40514_40814 , \40518_40818 );
and \U$32336 ( \40520_40820 , \30500_30802 , \27095_27397 );
and \U$32337 ( \40521_40821 , \31752_32054 , \26505_26807 );
nor \U$32338 ( \40522_40822 , \40520_40820 , \40521_40821 );
xnor \U$32339 ( \40523_40823 , \40522_40822 , \26993_27295 );
not \U$32340 ( \40524_40824 , \40523_40823 );
and \U$32341 ( \40525_40825 , \28782_29084 , \28768_29070 );
and \U$32342 ( \40526_40826 , \29966_30268 , \28224_28526 );
nor \U$32343 ( \40527_40827 , \40525_40825 , \40526_40826 );
xnor \U$32344 ( \40528_40828 , \40527_40827 , \28774_29076 );
xor \U$32345 ( \40529_40829 , \40524_40824 , \40528_40828 );
and \U$32346 ( \40530_40830 , \24970_25272 , \32503_32802 );
xor \U$32347 ( \40531_40831 , \40529_40829 , \40530_40830 );
xor \U$32348 ( \40532_40832 , \40519_40819 , \40531_40831 );
xor \U$32349 ( \40533_40833 , \40510_40810 , \40532_40832 );
and \U$32350 ( \40534_40834 , \40091_40391 , \40122_40422 );
and \U$32351 ( \40535_40835 , \40122_40422 , \40141_40441 );
and \U$32352 ( \40536_40836 , \40091_40391 , \40141_40441 );
or \U$32353 ( \40537_40837 , \40534_40834 , \40535_40835 , \40536_40836 );
xor \U$32354 ( \40538_40838 , \40533_40833 , \40537_40837 );
and \U$32355 ( \40539_40839 , \40142_40442 , \40146_40446 );
and \U$32356 ( \40540_40840 , \40147_40447 , \40150_40450 );
or \U$32357 ( \40541_40841 , \40539_40839 , \40540_40840 );
xor \U$32358 ( \40542_40842 , \40538_40838 , \40541_40841 );
buf g9b6c_GF_PartitionCandidate( \40543_40843_nG9b6c , \40542_40842 );
and \U$32359 ( \40544_40844 , \10402_10704 , \40543_40843_nG9b6c );
or \U$32360 ( \40545_40845 , \40482_40782 , \40544_40844 );
xor \U$32361 ( \40546_40846 , \10399_10703 , \40545_40845 );
buf \U$32362 ( \40547_40847 , \40546_40846 );
buf \U$32364 ( \40548_40848 , \40547_40847 );
xor \U$32365 ( \40549_40849 , \40481_40781 , \40548_40848 );
buf \U$32366 ( \40550_40850 , \40549_40849 );
xor \U$32367 ( \40551_40851 , \40468_40768 , \40550_40850 );
and \U$32368 ( \40552_40852 , \40010_40310 , \40016_40316 );
and \U$32369 ( \40553_40853 , \40010_40310 , \40023_40323 );
and \U$32370 ( \40554_40854 , \40016_40316 , \40023_40323 );
or \U$32371 ( \40555_40855 , \40552_40852 , \40553_40853 , \40554_40854 );
buf \U$32372 ( \40556_40856 , \40555_40855 );
and \U$32373 ( \40557_40857 , \14710_14631 , \37674_37974_nG9b87 );
and \U$32374 ( \40558_40858 , \14329_14628 , \38037_38337_nG9b84 );
or \U$32375 ( \40559_40859 , \40557_40857 , \40558_40858 );
xor \U$32376 ( \40560_40860 , \14328_14627 , \40559_40859 );
buf \U$32377 ( \40561_40861 , \40560_40860 );
buf \U$32379 ( \40562_40862 , \40561_40861 );
xor \U$32380 ( \40563_40863 , \40556_40856 , \40562_40862 );
and \U$32381 ( \40564_40864 , \10996_10421 , \39663_39963_nG9b75 );
and \U$32382 ( \40565_40865 , \10119_10418 , \39904_40204_nG9b72 );
or \U$32383 ( \40566_40866 , \40564_40864 , \40565_40865 );
xor \U$32384 ( \40567_40867 , \10118_10417 , \40566_40866 );
buf \U$32385 ( \40568_40868 , \40567_40867 );
buf \U$32387 ( \40569_40869 , \40568_40868 );
xor \U$32388 ( \40570_40870 , \40563_40863 , \40569_40869 );
buf \U$32389 ( \40571_40871 , \40570_40870 );
xor \U$32390 ( \40572_40872 , \40551_40851 , \40571_40871 );
buf \U$32391 ( \40573_40873 , \40572_40872 );
xor \U$32392 ( \40574_40874 , \40463_40763 , \40573_40873 );
buf \U$32393 ( \40575_40875 , \40574_40874 );
xor \U$32394 ( \40576_40876 , \40452_40752 , \40575_40875 );
and \U$32395 ( \40577_40877 , \40296_40596 , \40576_40876 );
and \U$32397 ( \40578_40878 , \40290_40590 , \40295_40595 );
or \U$32399 ( \40579_40879 , 1'b0 , \40578_40878 , 1'b0 );
xor \U$32400 ( \40580_40880 , \40577_40877 , \40579_40879 );
and \U$32402 ( \40581_40881 , \40283_40583 , \40289_40589 );
and \U$32403 ( \40582_40882 , \40285_40585 , \40289_40589 );
or \U$32404 ( \40583_40883 , 1'b0 , \40581_40881 , \40582_40882 );
xor \U$32405 ( \40584_40884 , \40580_40880 , \40583_40883 );
xor \U$32412 ( \40585_40885 , \40584_40884 , 1'b0 );
and \U$32413 ( \40586_40886 , \40446_40746 , \40451_40751 );
and \U$32414 ( \40587_40887 , \40446_40746 , \40575_40875 );
and \U$32415 ( \40588_40888 , \40451_40751 , \40575_40875 );
or \U$32416 ( \40589_40889 , \40586_40886 , \40587_40887 , \40588_40888 );
xor \U$32417 ( \40590_40890 , \40585_40885 , \40589_40889 );
and \U$32418 ( \40591_40891 , \40457_40757 , \40462_40762 );
and \U$32419 ( \40592_40892 , \40457_40757 , \40573_40873 );
and \U$32420 ( \40593_40893 , \40462_40762 , \40573_40873 );
or \U$32421 ( \40594_40894 , \40591_40891 , \40592_40892 , \40593_40893 );
buf \U$32422 ( \40595_40895 , \40594_40894 );
and \U$32423 ( \40596_40896 , \40468_40768 , \40550_40850 );
and \U$32424 ( \40597_40897 , \40468_40768 , \40571_40871 );
and \U$32425 ( \40598_40898 , \40550_40850 , \40571_40871 );
or \U$32426 ( \40599_40899 , \40596_40896 , \40597_40897 , \40598_40898 );
buf \U$32427 ( \40600_40900 , \40599_40899 );
and \U$32428 ( \40601_40901 , \17437_17297 , \36686_36986_nG9b90 );
and \U$32429 ( \40602_40902 , \16995_17294 , \36950_37250_nG9b8d );
or \U$32430 ( \40603_40903 , \40601_40901 , \40602_40902 );
xor \U$32431 ( \40604_40904 , \16994_17293 , \40603_40903 );
buf \U$32432 ( \40605_40905 , \40604_40904 );
buf \U$32434 ( \40606_40906 , \40605_40905 );
and \U$32435 ( \40607_40907 , \16405_15940 , \37307_37607_nG9b8a );
and \U$32436 ( \40608_40908 , \15638_15937 , \37674_37974_nG9b87 );
or \U$32437 ( \40609_40909 , \40607_40907 , \40608_40908 );
xor \U$32438 ( \40610_40910 , \15637_15936 , \40609_40909 );
buf \U$32439 ( \40611_40911 , \40610_40910 );
buf \U$32441 ( \40612_40912 , \40611_40911 );
xor \U$32442 ( \40613_40913 , \40606_40906 , \40612_40912 );
and \U$32443 ( \40614_40914 , \12183_12157 , \39291_39591_nG9b78 );
and \U$32444 ( \40615_40915 , \11855_12154 , \39663_39963_nG9b75 );
or \U$32445 ( \40616_40916 , \40614_40914 , \40615_40915 );
xor \U$32446 ( \40617_40917 , \11854_12153 , \40616_40916 );
buf \U$32447 ( \40618_40918 , \40617_40917 );
buf \U$32449 ( \40619_40919 , \40618_40918 );
xor \U$32450 ( \40620_40920 , \40613_40913 , \40619_40919 );
buf \U$32451 ( \40621_40921 , \40620_40920 );
and \U$32452 ( \40622_40922 , \23495_23201 , \33741_34041_nG9ba8 );
and \U$32453 ( \40623_40923 , \22899_23198 , \33994_34294_nG9ba5 );
or \U$32454 ( \40624_40924 , \40622_40922 , \40623_40923 );
xor \U$32455 ( \40625_40925 , \22898_23197 , \40624_40924 );
buf \U$32456 ( \40626_40926 , \40625_40925 );
buf \U$32458 ( \40627_40927 , \40626_40926 );
and \U$32459 ( \40628_40928 , \21908_21658 , \34343_34643_nG9ba2 );
and \U$32460 ( \40629_40929 , \21356_21655 , \34794_35094_nG9b9f );
or \U$32461 ( \40630_40930 , \40628_40928 , \40629_40929 );
xor \U$32462 ( \40631_40931 , \21355_21654 , \40630_40930 );
buf \U$32463 ( \40632_40932 , \40631_40931 );
buf \U$32465 ( \40633_40933 , \40632_40932 );
xor \U$32466 ( \40634_40934 , \40627_40927 , \40633_40933 );
and \U$32467 ( \40635_40935 , \20353_20155 , \35270_35570_nG9b9c );
and \U$32468 ( \40636_40936 , \19853_20152 , \35501_35801_nG9b99 );
or \U$32469 ( \40637_40937 , \40635_40935 , \40636_40936 );
xor \U$32470 ( \40638_40938 , \19852_20151 , \40637_40937 );
buf \U$32471 ( \40639_40939 , \40638_40938 );
buf \U$32473 ( \40640_40940 , \40639_40939 );
xor \U$32474 ( \40641_40941 , \40634_40934 , \40640_40940 );
buf \U$32475 ( \40642_40942 , \40641_40941 );
xor \U$32476 ( \40643_40943 , \40621_40921 , \40642_40942 );
and \U$32477 ( \40644_40944 , \40312_40612 , \40318_40618 );
and \U$32478 ( \40645_40945 , \40312_40612 , \40325_40625 );
and \U$32479 ( \40646_40946 , \40318_40618 , \40325_40625 );
or \U$32480 ( \40647_40947 , \40644_40944 , \40645_40945 , \40646_40946 );
buf \U$32481 ( \40648_40948 , \40647_40947 );
xor \U$32482 ( \40649_40949 , \40643_40943 , \40648_40948 );
buf \U$32483 ( \40650_40950 , \40649_40949 );
xor \U$32484 ( \40651_40951 , \40600_40900 , \40650_40950 );
and \U$32485 ( \40652_40952 , \40327_40627 , \40348_40648 );
and \U$32486 ( \40653_40953 , \40327_40627 , \40354_40654 );
and \U$32487 ( \40654_40954 , \40348_40648 , \40354_40654 );
or \U$32488 ( \40655_40955 , \40652_40952 , \40653_40953 , \40654_40954 );
buf \U$32489 ( \40656_40956 , \40655_40955 );
xor \U$32490 ( \40657_40957 , \40651_40951 , \40656_40956 );
buf \U$32491 ( \40658_40958 , \40657_40957 );
xor \U$32492 ( \40659_40959 , \40595_40895 , \40658_40958 );
and \U$32493 ( \40660_40960 , \40306_40606 , \40356_40656 );
and \U$32494 ( \40661_40961 , \40306_40606 , \40362_40662 );
and \U$32495 ( \40662_40962 , \40356_40656 , \40362_40662 );
or \U$32496 ( \40663_40963 , \40660_40960 , \40661_40961 , \40662_40962 );
buf \U$32497 ( \40664_40964 , \40663_40963 );
xor \U$32498 ( \40665_40965 , \40659_40959 , \40664_40964 );
buf \U$32499 ( \40666_40966 , \40665_40965 );
and \U$32500 ( \40667_40967 , \40301_40601 , \40364_40664 );
and \U$32501 ( \40668_40968 , \40301_40601 , \40444_40744 );
and \U$32502 ( \40669_40969 , \40364_40664 , \40444_40744 );
or \U$32503 ( \40670_40970 , \40667_40967 , \40668_40968 , \40669_40969 );
buf \U$32504 ( \40671_40971 , \40670_40970 );
xor \U$32505 ( \40672_40972 , \40666_40966 , \40671_40971 );
and \U$32506 ( \40673_40973 , \40425_40725 , \40431_40731 );
and \U$32507 ( \40674_40974 , \40425_40725 , \40438_40738 );
and \U$32508 ( \40675_40975 , \40431_40731 , \40438_40738 );
or \U$32509 ( \40676_40976 , \40673_40973 , \40674_40974 , \40675_40975 );
buf \U$32510 ( \40677_40977 , \40676_40976 );
and \U$32511 ( \40678_40978 , \14710_14631 , \38037_38337_nG9b84 );
and \U$32512 ( \40679_40979 , \14329_14628 , \38363_38663_nG9b81 );
or \U$32513 ( \40680_40980 , \40678_40978 , \40679_40979 );
xor \U$32514 ( \40681_40981 , \14328_14627 , \40680_40980 );
buf \U$32515 ( \40682_40982 , \40681_40981 );
buf \U$32517 ( \40683_40983 , \40682_40982 );
xor \U$32518 ( \40684_40984 , \40677_40977 , \40683_40983 );
and \U$32519 ( \40685_40985 , \10411_10707 , \40543_40843_nG9b6c );
and \U$32520 ( \40686_40986 , \40490_40790 , \40494_40794 );
and \U$32521 ( \40687_40987 , \40494_40794 , \40508_40808 );
and \U$32522 ( \40688_40988 , \40490_40790 , \40508_40808 );
or \U$32523 ( \40689_40989 , \40686_40986 , \40687_40987 , \40688_40988 );
and \U$32524 ( \40690_40990 , \40514_40814 , \40518_40818 );
and \U$32525 ( \40691_40991 , \40518_40818 , \40531_40831 );
and \U$32526 ( \40692_40992 , \40514_40814 , \40531_40831 );
or \U$32527 ( \40693_40993 , \40690_40990 , \40691_40991 , \40692_40992 );
xor \U$32528 ( \40694_40994 , \40689_40989 , \40693_40993 );
and \U$32529 ( \40695_40995 , \40524_40824 , \40528_40828 );
and \U$32530 ( \40696_40996 , \40528_40828 , \40530_40830 );
and \U$32531 ( \40697_40997 , \40524_40824 , \40530_40830 );
or \U$32532 ( \40698_40998 , \40695_40995 , \40696_40996 , \40697_40997 );
not \U$32533 ( \40699_40999 , \25474_25773 );
and \U$32534 ( \40700_41000 , \31752_32054 , \27095_27397 );
and \U$32535 ( \40701_41001 , \32495_32794 , \26505_26807 );
nor \U$32536 ( \40702_41002 , \40700_41000 , \40701_41001 );
xnor \U$32537 ( \40703_41003 , \40702_41002 , \26993_27295 );
xor \U$32538 ( \40704_41004 , \40699_40999 , \40703_41003 );
and \U$32539 ( \40705_41005 , \28232_28534 , \30521_30823 );
and \U$32540 ( \40706_41006 , \28782_29084 , \29944_30246 );
nor \U$32541 ( \40707_41007 , \40705_41005 , \40706_41006 );
xnor \U$32542 ( \40708_41008 , \40707_41007 , \30511_30813 );
xor \U$32543 ( \40709_41009 , \40704_41004 , \40708_41008 );
xor \U$32544 ( \40710_41010 , \40698_40998 , \40709_41009 );
and \U$32545 ( \40711_41011 , \40498_40798 , \40502_40802 );
and \U$32546 ( \40712_41012 , \40502_40802 , \40507_40807 );
and \U$32547 ( \40713_41013 , \40498_40798 , \40507_40807 );
or \U$32548 ( \40714_41014 , \40711_41011 , \40712_41012 , \40713_41013 );
buf \U$32549 ( \40715_41015 , \40523_40823 );
xor \U$32550 ( \40716_41016 , \40714_41014 , \40715_41015 );
and \U$32551 ( \40717_41017 , \29966_30268 , \28768_29070 );
and \U$32552 ( \40718_41018 , \30500_30802 , \28224_28526 );
nor \U$32553 ( \40719_41019 , \40717_41017 , \40718_41018 );
xnor \U$32554 ( \40720_41020 , \40719_41019 , \28774_29076 );
and \U$32555 ( \40721_41021 , \26527_26829 , \32555_32854 );
and \U$32556 ( \40722_41022 , \27011_27313 , \31765_32067 );
nor \U$32557 ( \40723_41023 , \40721_41021 , \40722_41022 );
xnor \U$32558 ( \40724_41024 , \40723_41023 , \32506_32805 );
xor \U$32559 ( \40725_41025 , \40720_41020 , \40724_41024 );
and \U$32560 ( \40726_41026 , \25516_25815 , \32503_32802 );
xor \U$32561 ( \40727_41027 , \40725_41025 , \40726_41026 );
xor \U$32562 ( \40728_41028 , \40716_41016 , \40727_41027 );
xor \U$32563 ( \40729_41029 , \40710_41010 , \40728_41028 );
xor \U$32564 ( \40730_41030 , \40694_40994 , \40729_41029 );
and \U$32565 ( \40731_41031 , \40486_40786 , \40509_40809 );
and \U$32566 ( \40732_41032 , \40509_40809 , \40532_40832 );
and \U$32567 ( \40733_41033 , \40486_40786 , \40532_40832 );
or \U$32568 ( \40734_41034 , \40731_41031 , \40732_41032 , \40733_41033 );
xor \U$32569 ( \40735_41035 , \40730_41030 , \40734_41034 );
and \U$32570 ( \40736_41036 , \40533_40833 , \40537_40837 );
and \U$32571 ( \40737_41037 , \40538_40838 , \40541_40841 );
or \U$32572 ( \40738_41038 , \40736_41036 , \40737_41037 );
xor \U$32573 ( \40739_41039 , \40735_41035 , \40738_41038 );
buf g9b69_GF_PartitionCandidate( \40740_41040_nG9b69 , \40739_41039 );
and \U$32574 ( \40741_41041 , \10402_10704 , \40740_41040_nG9b69 );
or \U$32575 ( \40742_41042 , \40685_40985 , \40741_41041 );
xor \U$32576 ( \40743_41043 , \10399_10703 , \40742_41042 );
buf \U$32577 ( \40744_41044 , \40743_41043 );
buf \U$32579 ( \40745_41045 , \40744_41044 );
xor \U$32580 ( \40746_41046 , \40684_40984 , \40745_41045 );
buf \U$32581 ( \40747_41047 , \40746_41046 );
and \U$32582 ( \40748_41048 , \40413_40713 , \40418_40718 );
and \U$32583 ( \40749_41049 , \40413_40713 , \40440_40740 );
and \U$32584 ( \40750_41050 , \40418_40718 , \40440_40740 );
or \U$32585 ( \40751_41051 , \40748_41048 , \40749_41049 , \40750_41050 );
buf \U$32586 ( \40752_41052 , \40751_41051 );
xor \U$32587 ( \40753_41053 , \40747_41047 , \40752_41052 );
and \U$32588 ( \40754_41054 , \18908_18702 , \35872_36172_nG9b96 );
and \U$32589 ( \40755_41055 , \18400_18699 , \36289_36589_nG9b93 );
or \U$32590 ( \40756_41056 , \40754_41054 , \40755_41055 );
xor \U$32591 ( \40757_41057 , \18399_18698 , \40756_41056 );
buf \U$32592 ( \40758_41058 , \40757_41057 );
buf \U$32594 ( \40759_41059 , \40758_41058 );
and \U$32595 ( \40760_41060 , \13431_13370 , \38668_38968_nG9b7e );
and \U$32596 ( \40761_41061 , \13068_13367 , \39034_39334_nG9b7b );
or \U$32597 ( \40762_41062 , \40760_41060 , \40761_41061 );
xor \U$32598 ( \40763_41063 , \13067_13366 , \40762_41062 );
buf \U$32599 ( \40764_41064 , \40763_41063 );
buf \U$32601 ( \40765_41065 , \40764_41064 );
xor \U$32602 ( \40766_41066 , \40759_41059 , \40765_41065 );
and \U$32603 ( \40767_41067 , \10996_10421 , \39904_40204_nG9b72 );
and \U$32604 ( \40768_41068 , \10119_10418 , \40152_40452_nG9b6f );
or \U$32605 ( \40769_41069 , \40767_41067 , \40768_41068 );
xor \U$32606 ( \40770_41070 , \10118_10417 , \40769_41069 );
buf \U$32607 ( \40771_41071 , \40770_41070 );
buf \U$32609 ( \40772_41072 , \40771_41071 );
xor \U$32610 ( \40773_41073 , \40766_41066 , \40772_41072 );
buf \U$32611 ( \40774_41074 , \40773_41073 );
xor \U$32612 ( \40775_41075 , \40753_41053 , \40774_41074 );
buf \U$32613 ( \40776_41076 , \40775_41075 );
and \U$32614 ( \40777_41077 , \40402_40702 , \40407_40707 );
and \U$32615 ( \40778_41078 , \40402_40702 , \40442_40742 );
and \U$32616 ( \40779_41079 , \40407_40707 , \40442_40742 );
or \U$32617 ( \40780_41080 , \40777_41077 , \40778_41078 , \40779_41079 );
buf \U$32618 ( \40781_41081 , \40780_41080 );
xor \U$32619 ( \40782_41082 , \40776_41076 , \40781_41081 );
and \U$32620 ( \40783_41083 , \40474_40774 , \40480_40780 );
and \U$32621 ( \40784_41084 , \40474_40774 , \40548_40848 );
and \U$32622 ( \40785_41085 , \40480_40780 , \40548_40848 );
or \U$32623 ( \40786_41086 , \40783_41083 , \40784_41084 , \40785_41085 );
buf \U$32624 ( \40787_41087 , \40786_41086 );
and \U$32625 ( \40788_41088 , \40556_40856 , \40562_40862 );
and \U$32626 ( \40789_41089 , \40556_40856 , \40569_40869 );
and \U$32627 ( \40790_41090 , \40562_40862 , \40569_40869 );
or \U$32628 ( \40791_41091 , \40788_41088 , \40789_41089 , \40790_41090 );
buf \U$32629 ( \40792_41092 , \40791_41091 );
xor \U$32630 ( \40793_41093 , \40787_41087 , \40792_41092 );
and \U$32632 ( \40794_41094 , \32617_32916 , \25561_25860_nG9bc9 );
or \U$32633 ( \40795_41095 , 1'b0 , \40794_41094 );
xor \U$32634 ( \40796_41096 , 1'b0 , \40795_41095 );
buf \U$32635 ( \40797_41097 , \40796_41096 );
buf \U$32637 ( \40798_41098 , \40797_41097 );
and \U$32638 ( \40799_41099 , \31989_31636 , \26585_26887_nG9bc6 );
and \U$32639 ( \40800_41100 , \31334_31633 , \27114_27416_nG9bc3 );
or \U$32640 ( \40801_41101 , \40799_41099 , \40800_41100 );
xor \U$32641 ( \40802_41102 , \31333_31632 , \40801_41101 );
buf \U$32642 ( \40803_41103 , \40802_41102 );
buf \U$32644 ( \40804_41104 , \40803_41103 );
xor \U$32645 ( \40805_41105 , \40798_41098 , \40804_41104 );
buf \U$32646 ( \40806_41106 , \40805_41105 );
and \U$32647 ( \40807_41107 , \27141_26431 , \31877_32179_nG9bb4 );
and \U$32648 ( \40808_41108 , \26129_26428 , \32589_32888_nG9bb1 );
or \U$32649 ( \40809_41109 , \40807_41107 , \40808_41108 );
xor \U$32650 ( \40810_41110 , \26128_26427 , \40809_41109 );
buf \U$32651 ( \40811_41111 , \40810_41110 );
buf \U$32653 ( \40812_41112 , \40811_41111 );
xor \U$32654 ( \40813_41113 , \40806_41106 , \40812_41112 );
and \U$32655 ( \40814_41114 , \25044_24792 , \32881_33181_nG9bae );
and \U$32656 ( \40815_41115 , \24490_24789 , \33313_33613_nG9bab );
or \U$32657 ( \40816_41116 , \40814_41114 , \40815_41115 );
xor \U$32658 ( \40817_41117 , \24489_24788 , \40816_41116 );
buf \U$32659 ( \40818_41118 , \40817_41117 );
buf \U$32661 ( \40819_41119 , \40818_41118 );
xor \U$32662 ( \40820_41120 , \40813_41113 , \40819_41119 );
buf \U$32663 ( \40821_41121 , \40820_41120 );
xor \U$32664 ( \40822_41122 , \40793_41093 , \40821_41121 );
buf \U$32665 ( \40823_41123 , \40822_41122 );
and \U$32666 ( \40824_41124 , \40370_40670 , \40375_40675 );
and \U$32667 ( \40825_41125 , \40370_40670 , \40400_40700 );
and \U$32668 ( \40826_41126 , \40375_40675 , \40400_40700 );
or \U$32669 ( \40827_41127 , \40824_41124 , \40825_41125 , \40826_41126 );
buf \U$32670 ( \40828_41128 , \40827_41127 );
xor \U$32671 ( \40829_41129 , \40823_41123 , \40828_41128 );
and \U$32672 ( \40830_41130 , \40333_40633 , \40339_40639 );
and \U$32673 ( \40831_41131 , \40333_40633 , \40346_40646 );
and \U$32674 ( \40832_41132 , \40339_40639 , \40346_40646 );
or \U$32675 ( \40833_41133 , \40830_41130 , \40831_41131 , \40832_41132 );
buf \U$32676 ( \40834_41134 , \40833_41133 );
and \U$32677 ( \40835_41135 , \40389_40689 , \40391_40691 );
and \U$32678 ( \40836_41136 , \40389_40689 , \40398_40698 );
and \U$32679 ( \40837_41137 , \40391_40691 , \40398_40698 );
or \U$32680 ( \40838_41138 , \40835_41135 , \40836_41136 , \40837_41137 );
buf \U$32681 ( \40839_41139 , \40838_41138 );
xor \U$32682 ( \40840_41140 , \40834_41134 , \40839_41139 );
and \U$32683 ( \40841_41141 , \40381_40681 , \40387_40687 );
buf \U$32684 ( \40842_41142 , \40841_41141 );
and \U$32685 ( \40843_41143 , \30670_29853 , \28300_28602_nG9bc0 );
and \U$32686 ( \40844_41144 , \29551_29850 , \28877_29179_nG9bbd );
or \U$32687 ( \40845_41145 , \40843_41143 , \40844_41144 );
xor \U$32688 ( \40846_41146 , \29550_29849 , \40845_41145 );
buf \U$32689 ( \40847_41147 , \40846_41146 );
buf \U$32691 ( \40848_41148 , \40847_41147 );
xor \U$32692 ( \40849_41149 , \40842_41142 , \40848_41148 );
and \U$32693 ( \40850_41150 , \28946_28118 , \30064_30366_nG9bba );
and \U$32694 ( \40851_41151 , \27816_28115 , \30638_30940_nG9bb7 );
or \U$32695 ( \40852_41152 , \40850_41150 , \40851_41151 );
xor \U$32696 ( \40853_41153 , \27815_28114 , \40852_41152 );
buf \U$32697 ( \40854_41154 , \40853_41153 );
buf \U$32699 ( \40855_41155 , \40854_41154 );
xor \U$32700 ( \40856_41156 , \40849_41149 , \40855_41155 );
buf \U$32701 ( \40857_41157 , \40856_41156 );
xor \U$32702 ( \40858_41158 , \40840_41140 , \40857_41157 );
buf \U$32703 ( \40859_41159 , \40858_41158 );
xor \U$32704 ( \40860_41160 , \40829_41129 , \40859_41159 );
buf \U$32705 ( \40861_41161 , \40860_41160 );
xor \U$32706 ( \40862_41162 , \40782_41082 , \40861_41161 );
buf \U$32707 ( \40863_41163 , \40862_41162 );
xor \U$32708 ( \40864_41164 , \40672_40972 , \40863_41163 );
and \U$32709 ( \40865_41165 , \40590_40890 , \40864_41164 );
and \U$32711 ( \40866_41166 , \40584_40884 , \40589_40889 );
or \U$32713 ( \40867_41167 , 1'b0 , \40866_41166 , 1'b0 );
xor \U$32714 ( \40868_41168 , \40865_41165 , \40867_41167 );
and \U$32716 ( \40869_41169 , \40577_40877 , \40583_40883 );
and \U$32717 ( \40870_41170 , \40579_40879 , \40583_40883 );
or \U$32718 ( \40871_41171 , 1'b0 , \40869_41169 , \40870_41170 );
xor \U$32719 ( \40872_41172 , \40868_41168 , \40871_41171 );
xor \U$32726 ( \40873_41173 , \40872_41172 , 1'b0 );
and \U$32727 ( \40874_41174 , \40666_40966 , \40671_40971 );
and \U$32728 ( \40875_41175 , \40666_40966 , \40863_41163 );
and \U$32729 ( \40876_41176 , \40671_40971 , \40863_41163 );
or \U$32730 ( \40877_41177 , \40874_41174 , \40875_41175 , \40876_41176 );
xor \U$32731 ( \40878_41178 , \40873_41173 , \40877_41177 );
and \U$32732 ( \40879_41179 , \40776_41076 , \40781_41081 );
and \U$32733 ( \40880_41180 , \40776_41076 , \40861_41161 );
and \U$32734 ( \40881_41181 , \40781_41081 , \40861_41161 );
or \U$32735 ( \40882_41182 , \40879_41179 , \40880_41180 , \40881_41181 );
buf \U$32736 ( \40883_41183 , \40882_41182 );
and \U$32737 ( \40884_41184 , \40747_41047 , \40752_41052 );
and \U$32738 ( \40885_41185 , \40747_41047 , \40774_41074 );
and \U$32739 ( \40886_41186 , \40752_41052 , \40774_41074 );
or \U$32740 ( \40887_41187 , \40884_41184 , \40885_41185 , \40886_41186 );
buf \U$32741 ( \40888_41188 , \40887_41187 );
and \U$32742 ( \40889_41189 , \18908_18702 , \36289_36589_nG9b93 );
and \U$32743 ( \40890_41190 , \18400_18699 , \36686_36986_nG9b90 );
or \U$32744 ( \40891_41191 , \40889_41189 , \40890_41190 );
xor \U$32745 ( \40892_41192 , \18399_18698 , \40891_41191 );
buf \U$32746 ( \40893_41193 , \40892_41192 );
buf \U$32748 ( \40894_41194 , \40893_41193 );
and \U$32749 ( \40895_41195 , \13431_13370 , \39034_39334_nG9b7b );
and \U$32750 ( \40896_41196 , \13068_13367 , \39291_39591_nG9b78 );
or \U$32751 ( \40897_41197 , \40895_41195 , \40896_41196 );
xor \U$32752 ( \40898_41198 , \13067_13366 , \40897_41197 );
buf \U$32753 ( \40899_41199 , \40898_41198 );
buf \U$32755 ( \40900_41200 , \40899_41199 );
xor \U$32756 ( \40901_41201 , \40894_41194 , \40900_41200 );
and \U$32757 ( \40902_41202 , \10996_10421 , \40152_40452_nG9b6f );
and \U$32758 ( \40903_41203 , \10119_10418 , \40543_40843_nG9b6c );
or \U$32759 ( \40904_41204 , \40902_41202 , \40903_41203 );
xor \U$32760 ( \40905_41205 , \10118_10417 , \40904_41204 );
buf \U$32761 ( \40906_41206 , \40905_41205 );
buf \U$32763 ( \40907_41207 , \40906_41206 );
xor \U$32764 ( \40908_41208 , \40901_41201 , \40907_41207 );
buf \U$32765 ( \40909_41209 , \40908_41208 );
and \U$32766 ( \40910_41210 , \40606_40906 , \40612_40912 );
and \U$32767 ( \40911_41211 , \40606_40906 , \40619_40919 );
and \U$32768 ( \40912_41212 , \40612_40912 , \40619_40919 );
or \U$32769 ( \40913_41213 , \40910_41210 , \40911_41211 , \40912_41212 );
buf \U$32770 ( \40914_41214 , \40913_41213 );
xor \U$32771 ( \40915_41215 , \40909_41209 , \40914_41214 );
and \U$32772 ( \40916_41216 , \23495_23201 , \33994_34294_nG9ba5 );
and \U$32773 ( \40917_41217 , \22899_23198 , \34343_34643_nG9ba2 );
or \U$32774 ( \40918_41218 , \40916_41216 , \40917_41217 );
xor \U$32775 ( \40919_41219 , \22898_23197 , \40918_41218 );
buf \U$32776 ( \40920_41220 , \40919_41219 );
buf \U$32778 ( \40921_41221 , \40920_41220 );
and \U$32779 ( \40922_41222 , \21908_21658 , \34794_35094_nG9b9f );
and \U$32780 ( \40923_41223 , \21356_21655 , \35270_35570_nG9b9c );
or \U$32781 ( \40924_41224 , \40922_41222 , \40923_41223 );
xor \U$32782 ( \40925_41225 , \21355_21654 , \40924_41224 );
buf \U$32783 ( \40926_41226 , \40925_41225 );
buf \U$32785 ( \40927_41227 , \40926_41226 );
xor \U$32786 ( \40928_41228 , \40921_41221 , \40927_41227 );
and \U$32787 ( \40929_41229 , \20353_20155 , \35501_35801_nG9b99 );
and \U$32788 ( \40930_41230 , \19853_20152 , \35872_36172_nG9b96 );
or \U$32789 ( \40931_41231 , \40929_41229 , \40930_41230 );
xor \U$32790 ( \40932_41232 , \19852_20151 , \40931_41231 );
buf \U$32791 ( \40933_41233 , \40932_41232 );
buf \U$32793 ( \40934_41234 , \40933_41233 );
xor \U$32794 ( \40935_41235 , \40928_41228 , \40934_41234 );
buf \U$32795 ( \40936_41236 , \40935_41235 );
xor \U$32796 ( \40937_41237 , \40915_41215 , \40936_41236 );
buf \U$32797 ( \40938_41238 , \40937_41237 );
xor \U$32798 ( \40939_41239 , \40888_41188 , \40938_41238 );
and \U$32799 ( \40940_41240 , \40621_40921 , \40642_40942 );
and \U$32800 ( \40941_41241 , \40621_40921 , \40648_40948 );
and \U$32801 ( \40942_41242 , \40642_40942 , \40648_40948 );
or \U$32802 ( \40943_41243 , \40940_41240 , \40941_41241 , \40942_41242 );
buf \U$32803 ( \40944_41244 , \40943_41243 );
xor \U$32804 ( \40945_41245 , \40939_41239 , \40944_41244 );
buf \U$32805 ( \40946_41246 , \40945_41245 );
xor \U$32806 ( \40947_41247 , \40883_41183 , \40946_41246 );
and \U$32807 ( \40948_41248 , \40600_40900 , \40650_40950 );
and \U$32808 ( \40949_41249 , \40600_40900 , \40656_40956 );
and \U$32809 ( \40950_41250 , \40650_40950 , \40656_40956 );
or \U$32810 ( \40951_41251 , \40948_41248 , \40949_41249 , \40950_41250 );
buf \U$32811 ( \40952_41252 , \40951_41251 );
xor \U$32812 ( \40953_41253 , \40947_41247 , \40952_41252 );
buf \U$32813 ( \40954_41254 , \40953_41253 );
and \U$32814 ( \40955_41255 , \40595_40895 , \40658_40958 );
and \U$32815 ( \40956_41256 , \40595_40895 , \40664_40964 );
and \U$32816 ( \40957_41257 , \40658_40958 , \40664_40964 );
or \U$32817 ( \40958_41258 , \40955_41255 , \40956_41256 , \40957_41257 );
buf \U$32818 ( \40959_41259 , \40958_41258 );
xor \U$32819 ( \40960_41260 , \40954_41254 , \40959_41259 );
and \U$32820 ( \40961_41261 , \40823_41123 , \40828_41128 );
and \U$32821 ( \40962_41262 , \40823_41123 , \40859_41159 );
and \U$32822 ( \40963_41263 , \40828_41128 , \40859_41159 );
or \U$32823 ( \40964_41264 , \40961_41261 , \40962_41262 , \40963_41263 );
buf \U$32824 ( \40965_41265 , \40964_41264 );
and \U$32825 ( \40966_41266 , \40798_41098 , \40804_41104 );
buf \U$32826 ( \40967_41267 , \40966_41266 );
and \U$32827 ( \40968_41268 , \30670_29853 , \28877_29179_nG9bbd );
and \U$32828 ( \40969_41269 , \29551_29850 , \30064_30366_nG9bba );
or \U$32829 ( \40970_41270 , \40968_41268 , \40969_41269 );
xor \U$32830 ( \40971_41271 , \29550_29849 , \40970_41270 );
buf \U$32831 ( \40972_41272 , \40971_41271 );
buf \U$32833 ( \40973_41273 , \40972_41272 );
xor \U$32834 ( \40974_41274 , \40967_41267 , \40973_41273 );
and \U$32835 ( \40975_41275 , \28946_28118 , \30638_30940_nG9bb7 );
and \U$32836 ( \40976_41276 , \27816_28115 , \31877_32179_nG9bb4 );
or \U$32837 ( \40977_41277 , \40975_41275 , \40976_41276 );
xor \U$32838 ( \40978_41278 , \27815_28114 , \40977_41277 );
buf \U$32839 ( \40979_41279 , \40978_41278 );
buf \U$32841 ( \40980_41280 , \40979_41279 );
xor \U$32842 ( \40981_41281 , \40974_41274 , \40980_41280 );
buf \U$32843 ( \40982_41282 , \40981_41281 );
and \U$32844 ( \40983_41283 , \40627_40927 , \40633_40933 );
and \U$32845 ( \40984_41284 , \40627_40927 , \40640_40940 );
and \U$32846 ( \40985_41285 , \40633_40933 , \40640_40940 );
or \U$32847 ( \40986_41286 , \40983_41283 , \40984_41284 , \40985_41285 );
buf \U$32848 ( \40987_41287 , \40986_41286 );
xor \U$32849 ( \40988_41288 , \40982_41282 , \40987_41287 );
and \U$32850 ( \40989_41289 , \40806_41106 , \40812_41112 );
and \U$32851 ( \40990_41290 , \40806_41106 , \40819_41119 );
and \U$32852 ( \40991_41291 , \40812_41112 , \40819_41119 );
or \U$32853 ( \40992_41292 , \40989_41289 , \40990_41290 , \40991_41291 );
buf \U$32854 ( \40993_41293 , \40992_41292 );
xor \U$32855 ( \40994_41294 , \40988_41288 , \40993_41293 );
buf \U$32856 ( \40995_41295 , \40994_41294 );
and \U$32857 ( \40996_41296 , \40842_41142 , \40848_41148 );
and \U$32858 ( \40997_41297 , \40842_41142 , \40855_41155 );
and \U$32859 ( \40998_41298 , \40848_41148 , \40855_41155 );
or \U$32860 ( \40999_41299 , \40996_41296 , \40997_41297 , \40998_41298 );
buf \U$32861 ( \41000_41300 , \40999_41299 );
and \U$32862 ( \41001_41301 , \17437_17297 , \36950_37250_nG9b8d );
and \U$32863 ( \41002_41302 , \16995_17294 , \37307_37607_nG9b8a );
or \U$32864 ( \41003_41303 , \41001_41301 , \41002_41302 );
xor \U$32865 ( \41004_41304 , \16994_17293 , \41003_41303 );
buf \U$32866 ( \41005_41305 , \41004_41304 );
buf \U$32868 ( \41006_41306 , \41005_41305 );
xor \U$32869 ( \41007_41307 , \41000_41300 , \41006_41306 );
and \U$32870 ( \41008_41308 , \12183_12157 , \39663_39963_nG9b75 );
and \U$32871 ( \41009_41309 , \11855_12154 , \39904_40204_nG9b72 );
or \U$32872 ( \41010_41310 , \41008_41308 , \41009_41309 );
xor \U$32873 ( \41011_41311 , \11854_12153 , \41010_41310 );
buf \U$32874 ( \41012_41312 , \41011_41311 );
buf \U$32876 ( \41013_41313 , \41012_41312 );
xor \U$32877 ( \41014_41314 , \41007_41307 , \41013_41313 );
buf \U$32878 ( \41015_41315 , \41014_41314 );
xor \U$32879 ( \41016_41316 , \40995_41295 , \41015_41315 );
and \U$32880 ( \41017_41317 , \16405_15940 , \37674_37974_nG9b87 );
and \U$32881 ( \41018_41318 , \15638_15937 , \38037_38337_nG9b84 );
or \U$32882 ( \41019_41319 , \41017_41317 , \41018_41318 );
xor \U$32883 ( \41020_41320 , \15637_15936 , \41019_41319 );
buf \U$32884 ( \41021_41321 , \41020_41320 );
buf \U$32886 ( \41022_41322 , \41021_41321 );
and \U$32887 ( \41023_41323 , \14710_14631 , \38363_38663_nG9b81 );
and \U$32888 ( \41024_41324 , \14329_14628 , \38668_38968_nG9b7e );
or \U$32889 ( \41025_41325 , \41023_41323 , \41024_41324 );
xor \U$32890 ( \41026_41326 , \14328_14627 , \41025_41325 );
buf \U$32891 ( \41027_41327 , \41026_41326 );
buf \U$32893 ( \41028_41328 , \41027_41327 );
xor \U$32894 ( \41029_41329 , \41022_41322 , \41028_41328 );
and \U$32895 ( \41030_41330 , \10411_10707 , \40740_41040_nG9b69 );
and \U$32896 ( \41031_41331 , \40714_41014 , \40715_41015 );
and \U$32897 ( \41032_41332 , \40715_41015 , \40727_41027 );
and \U$32898 ( \41033_41333 , \40714_41014 , \40727_41027 );
or \U$32899 ( \41034_41334 , \41031_41331 , \41032_41332 , \41033_41333 );
and \U$32900 ( \41035_41335 , \40698_40998 , \40709_41009 );
and \U$32901 ( \41036_41336 , \40709_41009 , \40728_41028 );
and \U$32902 ( \41037_41337 , \40698_40998 , \40728_41028 );
or \U$32903 ( \41038_41338 , \41035_41335 , \41036_41336 , \41037_41337 );
xor \U$32904 ( \41039_41339 , \41034_41334 , \41038_41338 );
and \U$32905 ( \41040_41340 , \40699_40999 , \40703_41003 );
and \U$32906 ( \41041_41341 , \40703_41003 , \40708_41008 );
and \U$32907 ( \41042_41342 , \40699_40999 , \40708_41008 );
or \U$32908 ( \41043_41343 , \41040_41340 , \41041_41341 , \41042_41342 );
and \U$32909 ( \41044_41344 , \32495_32794 , \27095_27397 );
not \U$32910 ( \41045_41345 , \41044_41344 );
xnor \U$32911 ( \41046_41346 , \41045_41345 , \26993_27295 );
and \U$32912 ( \41047_41347 , \27011_27313 , \32555_32854 );
and \U$32913 ( \41048_41348 , \28232_28534 , \31765_32067 );
nor \U$32914 ( \41049_41349 , \41047_41347 , \41048_41348 );
xnor \U$32915 ( \41050_41350 , \41049_41349 , \32506_32805 );
xor \U$32916 ( \41051_41351 , \41046_41346 , \41050_41350 );
and \U$32917 ( \41052_41352 , \26527_26829 , \32503_32802 );
xor \U$32918 ( \41053_41353 , \41051_41351 , \41052_41352 );
xor \U$32919 ( \41054_41354 , \41043_41343 , \41053_41353 );
and \U$32920 ( \41055_41355 , \40720_41020 , \40724_41024 );
and \U$32921 ( \41056_41356 , \40724_41024 , \40726_41026 );
and \U$32922 ( \41057_41357 , \40720_41020 , \40726_41026 );
or \U$32923 ( \41058_41358 , \41055_41355 , \41056_41356 , \41057_41357 );
and \U$32924 ( \41059_41359 , \30500_30802 , \28768_29070 );
and \U$32925 ( \41060_41360 , \31752_32054 , \28224_28526 );
nor \U$32926 ( \41061_41361 , \41059_41359 , \41060_41360 );
xnor \U$32927 ( \41062_41362 , \41061_41361 , \28774_29076 );
not \U$32928 ( \41063_41363 , \41062_41362 );
xor \U$32929 ( \41064_41364 , \41058_41358 , \41063_41363 );
and \U$32930 ( \41065_41365 , \28782_29084 , \30521_30823 );
and \U$32931 ( \41066_41366 , \29966_30268 , \29944_30246 );
nor \U$32932 ( \41067_41367 , \41065_41365 , \41066_41366 );
xnor \U$32933 ( \41068_41368 , \41067_41367 , \30511_30813 );
xor \U$32934 ( \41069_41369 , \41064_41364 , \41068_41368 );
xor \U$32935 ( \41070_41370 , \41054_41354 , \41069_41369 );
xor \U$32936 ( \41071_41371 , \41039_41339 , \41070_41370 );
and \U$32937 ( \41072_41372 , \40689_40989 , \40693_40993 );
and \U$32938 ( \41073_41373 , \40693_40993 , \40729_41029 );
and \U$32939 ( \41074_41374 , \40689_40989 , \40729_41029 );
or \U$32940 ( \41075_41375 , \41072_41372 , \41073_41373 , \41074_41374 );
xor \U$32941 ( \41076_41376 , \41071_41371 , \41075_41375 );
and \U$32942 ( \41077_41377 , \40730_41030 , \40734_41034 );
and \U$32943 ( \41078_41378 , \40735_41035 , \40738_41038 );
or \U$32944 ( \41079_41379 , \41077_41377 , \41078_41378 );
xor \U$32945 ( \41080_41380 , \41076_41376 , \41079_41379 );
buf g9b66_GF_PartitionCandidate( \41081_41381_nG9b66 , \41080_41380 );
and \U$32946 ( \41082_41382 , \10402_10704 , \41081_41381_nG9b66 );
or \U$32947 ( \41083_41383 , \41030_41330 , \41082_41382 );
xor \U$32948 ( \41084_41384 , \10399_10703 , \41083_41383 );
buf \U$32949 ( \41085_41385 , \41084_41384 );
buf \U$32951 ( \41086_41386 , \41085_41385 );
xor \U$32952 ( \41087_41387 , \41029_41329 , \41086_41386 );
buf \U$32953 ( \41088_41388 , \41087_41387 );
xor \U$32954 ( \41089_41389 , \41016_41316 , \41088_41388 );
buf \U$32955 ( \41090_41390 , \41089_41389 );
xor \U$32956 ( \41091_41391 , \40965_41265 , \41090_41390 );
and \U$32957 ( \41092_41392 , \40787_41087 , \40792_41092 );
and \U$32958 ( \41093_41393 , \40787_41087 , \40821_41121 );
and \U$32959 ( \41094_41394 , \40792_41092 , \40821_41121 );
or \U$32960 ( \41095_41395 , \41092_41392 , \41093_41393 , \41094_41394 );
buf \U$32961 ( \41096_41396 , \41095_41395 );
and \U$32962 ( \41097_41397 , \40834_41134 , \40839_41139 );
and \U$32963 ( \41098_41398 , \40834_41134 , \40857_41157 );
and \U$32964 ( \41099_41399 , \40839_41139 , \40857_41157 );
or \U$32965 ( \41100_41400 , \41097_41397 , \41098_41398 , \41099_41399 );
buf \U$32966 ( \41101_41401 , \41100_41400 );
xor \U$32967 ( \41102_41402 , \41096_41396 , \41101_41401 );
and \U$32968 ( \41103_41403 , \40677_40977 , \40683_40983 );
and \U$32969 ( \41104_41404 , \40677_40977 , \40745_41045 );
and \U$32970 ( \41105_41405 , \40683_40983 , \40745_41045 );
or \U$32971 ( \41106_41406 , \41103_41403 , \41104_41404 , \41105_41405 );
buf \U$32972 ( \41107_41407 , \41106_41406 );
and \U$32973 ( \41108_41408 , \40759_41059 , \40765_41065 );
and \U$32974 ( \41109_41409 , \40759_41059 , \40772_41072 );
and \U$32975 ( \41110_41410 , \40765_41065 , \40772_41072 );
or \U$32976 ( \41111_41411 , \41108_41408 , \41109_41409 , \41110_41410 );
buf \U$32977 ( \41112_41412 , \41111_41411 );
xor \U$32978 ( \41113_41413 , \41107_41407 , \41112_41412 );
and \U$32980 ( \41114_41414 , \32617_32916 , \26585_26887_nG9bc6 );
or \U$32981 ( \41115_41415 , 1'b0 , \41114_41414 );
xor \U$32982 ( \41116_41416 , 1'b0 , \41115_41415 );
buf \U$32983 ( \41117_41417 , \41116_41416 );
buf \U$32985 ( \41118_41418 , \41117_41417 );
and \U$32986 ( \41119_41419 , \31989_31636 , \27114_27416_nG9bc3 );
and \U$32987 ( \41120_41420 , \31334_31633 , \28300_28602_nG9bc0 );
or \U$32988 ( \41121_41421 , \41119_41419 , \41120_41420 );
xor \U$32989 ( \41122_41422 , \31333_31632 , \41121_41421 );
buf \U$32990 ( \41123_41423 , \41122_41422 );
buf \U$32992 ( \41124_41424 , \41123_41423 );
xor \U$32993 ( \41125_41425 , \41118_41418 , \41124_41424 );
buf \U$32994 ( \41126_41426 , \41125_41425 );
and \U$32995 ( \41127_41427 , \27141_26431 , \32589_32888_nG9bb1 );
and \U$32996 ( \41128_41428 , \26129_26428 , \32881_33181_nG9bae );
or \U$32997 ( \41129_41429 , \41127_41427 , \41128_41428 );
xor \U$32998 ( \41130_41430 , \26128_26427 , \41129_41429 );
buf \U$32999 ( \41131_41431 , \41130_41430 );
buf \U$33001 ( \41132_41432 , \41131_41431 );
xor \U$33002 ( \41133_41433 , \41126_41426 , \41132_41432 );
and \U$33003 ( \41134_41434 , \25044_24792 , \33313_33613_nG9bab );
and \U$33004 ( \41135_41435 , \24490_24789 , \33741_34041_nG9ba8 );
or \U$33005 ( \41136_41436 , \41134_41434 , \41135_41435 );
xor \U$33006 ( \41137_41437 , \24489_24788 , \41136_41436 );
buf \U$33007 ( \41138_41438 , \41137_41437 );
buf \U$33009 ( \41139_41439 , \41138_41438 );
xor \U$33010 ( \41140_41440 , \41133_41433 , \41139_41439 );
buf \U$33011 ( \41141_41441 , \41140_41440 );
xor \U$33012 ( \41142_41442 , \41113_41413 , \41141_41441 );
buf \U$33013 ( \41143_41443 , \41142_41442 );
xor \U$33014 ( \41144_41444 , \41102_41402 , \41143_41443 );
buf \U$33015 ( \41145_41445 , \41144_41444 );
xor \U$33016 ( \41146_41446 , \41091_41391 , \41145_41445 );
buf \U$33017 ( \41147_41447 , \41146_41446 );
xor \U$33018 ( \41148_41448 , \40960_41260 , \41147_41447 );
and \U$33019 ( \41149_41449 , \40878_41178 , \41148_41448 );
and \U$33021 ( \41150_41450 , \40872_41172 , \40877_41177 );
or \U$33023 ( \41151_41451 , 1'b0 , \41150_41450 , 1'b0 );
xor \U$33024 ( \41152_41452 , \41149_41449 , \41151_41451 );
and \U$33026 ( \41153_41453 , \40865_41165 , \40871_41171 );
and \U$33027 ( \41154_41454 , \40867_41167 , \40871_41171 );
or \U$33028 ( \41155_41455 , 1'b0 , \41153_41453 , \41154_41454 );
xor \U$33029 ( \41156_41456 , \41152_41452 , \41155_41455 );
xor \U$33036 ( \41157_41457 , \41156_41456 , 1'b0 );
and \U$33037 ( \41158_41458 , \40954_41254 , \40959_41259 );
and \U$33038 ( \41159_41459 , \40954_41254 , \41147_41447 );
and \U$33039 ( \41160_41460 , \40959_41259 , \41147_41447 );
or \U$33040 ( \41161_41461 , \41158_41458 , \41159_41459 , \41160_41460 );
xor \U$33041 ( \41162_41462 , \41157_41457 , \41161_41461 );
and \U$33042 ( \41163_41463 , \40965_41265 , \41090_41390 );
and \U$33043 ( \41164_41464 , \40965_41265 , \41145_41445 );
and \U$33044 ( \41165_41465 , \41090_41390 , \41145_41445 );
or \U$33045 ( \41166_41466 , \41163_41463 , \41164_41464 , \41165_41465 );
buf \U$33046 ( \41167_41467 , \41166_41466 );
and \U$33047 ( \41168_41468 , \40888_41188 , \40938_41238 );
and \U$33048 ( \41169_41469 , \40888_41188 , \40944_41244 );
and \U$33049 ( \41170_41470 , \40938_41238 , \40944_41244 );
or \U$33050 ( \41171_41471 , \41168_41468 , \41169_41469 , \41170_41470 );
buf \U$33051 ( \41172_41472 , \41171_41471 );
xor \U$33052 ( \41173_41473 , \41167_41467 , \41172_41472 );
and \U$33053 ( \41174_41474 , \40995_41295 , \41015_41315 );
and \U$33054 ( \41175_41475 , \40995_41295 , \41088_41388 );
and \U$33055 ( \41176_41476 , \41015_41315 , \41088_41388 );
or \U$33056 ( \41177_41477 , \41174_41474 , \41175_41475 , \41176_41476 );
buf \U$33057 ( \41178_41478 , \41177_41477 );
and \U$33058 ( \41179_41479 , \16405_15940 , \38037_38337_nG9b84 );
and \U$33059 ( \41180_41480 , \15638_15937 , \38363_38663_nG9b81 );
or \U$33060 ( \41181_41481 , \41179_41479 , \41180_41480 );
xor \U$33061 ( \41182_41482 , \15637_15936 , \41181_41481 );
buf \U$33062 ( \41183_41483 , \41182_41482 );
buf \U$33064 ( \41184_41484 , \41183_41483 );
and \U$33065 ( \41185_41485 , \14710_14631 , \38668_38968_nG9b7e );
and \U$33066 ( \41186_41486 , \14329_14628 , \39034_39334_nG9b7b );
or \U$33067 ( \41187_41487 , \41185_41485 , \41186_41486 );
xor \U$33068 ( \41188_41488 , \14328_14627 , \41187_41487 );
buf \U$33069 ( \41189_41489 , \41188_41488 );
buf \U$33071 ( \41190_41490 , \41189_41489 );
xor \U$33072 ( \41191_41491 , \41184_41484 , \41190_41490 );
and \U$33073 ( \41192_41492 , \10996_10421 , \40543_40843_nG9b6c );
and \U$33074 ( \41193_41493 , \10119_10418 , \40740_41040_nG9b69 );
or \U$33075 ( \41194_41494 , \41192_41492 , \41193_41493 );
xor \U$33076 ( \41195_41495 , \10118_10417 , \41194_41494 );
buf \U$33077 ( \41196_41496 , \41195_41495 );
buf \U$33079 ( \41197_41497 , \41196_41496 );
xor \U$33080 ( \41198_41498 , \41191_41491 , \41197_41497 );
buf \U$33081 ( \41199_41499 , \41198_41498 );
and \U$33082 ( \41200_41500 , \40982_41282 , \40987_41287 );
and \U$33083 ( \41201_41501 , \40982_41282 , \40993_41293 );
and \U$33084 ( \41202_41502 , \40987_41287 , \40993_41293 );
or \U$33085 ( \41203_41503 , \41200_41500 , \41201_41501 , \41202_41502 );
buf \U$33086 ( \41204_41504 , \41203_41503 );
xor \U$33087 ( \41205_41505 , \41199_41499 , \41204_41504 );
and \U$33088 ( \41206_41506 , \41000_41300 , \41006_41306 );
and \U$33089 ( \41207_41507 , \41000_41300 , \41013_41313 );
and \U$33090 ( \41208_41508 , \41006_41306 , \41013_41313 );
or \U$33091 ( \41209_41509 , \41206_41506 , \41207_41507 , \41208_41508 );
buf \U$33092 ( \41210_41510 , \41209_41509 );
xor \U$33093 ( \41211_41511 , \41205_41505 , \41210_41510 );
buf \U$33094 ( \41212_41512 , \41211_41511 );
xor \U$33095 ( \41213_41513 , \41178_41478 , \41212_41512 );
and \U$33096 ( \41214_41514 , \40909_41209 , \40914_41214 );
and \U$33097 ( \41215_41515 , \40909_41209 , \40936_41236 );
and \U$33098 ( \41216_41516 , \40914_41214 , \40936_41236 );
or \U$33099 ( \41217_41517 , \41214_41514 , \41215_41515 , \41216_41516 );
buf \U$33100 ( \41218_41518 , \41217_41517 );
xor \U$33101 ( \41219_41519 , \41213_41513 , \41218_41518 );
buf \U$33102 ( \41220_41520 , \41219_41519 );
xor \U$33103 ( \41221_41521 , \41173_41473 , \41220_41520 );
buf \U$33104 ( \41222_41522 , \41221_41521 );
and \U$33105 ( \41223_41523 , \40883_41183 , \40946_41246 );
and \U$33106 ( \41224_41524 , \40883_41183 , \40952_41252 );
and \U$33107 ( \41225_41525 , \40946_41246 , \40952_41252 );
or \U$33108 ( \41226_41526 , \41223_41523 , \41224_41524 , \41225_41525 );
buf \U$33109 ( \41227_41527 , \41226_41526 );
xor \U$33110 ( \41228_41528 , \41222_41522 , \41227_41527 );
and \U$33111 ( \41229_41529 , \25044_24792 , \33741_34041_nG9ba8 );
and \U$33112 ( \41230_41530 , \24490_24789 , \33994_34294_nG9ba5 );
or \U$33113 ( \41231_41531 , \41229_41529 , \41230_41530 );
xor \U$33114 ( \41232_41532 , \24489_24788 , \41231_41531 );
buf \U$33115 ( \41233_41533 , \41232_41532 );
buf \U$33117 ( \41234_41534 , \41233_41533 );
and \U$33118 ( \41235_41535 , \21908_21658 , \35270_35570_nG9b9c );
and \U$33119 ( \41236_41536 , \21356_21655 , \35501_35801_nG9b99 );
or \U$33120 ( \41237_41537 , \41235_41535 , \41236_41536 );
xor \U$33121 ( \41238_41538 , \21355_21654 , \41237_41537 );
buf \U$33122 ( \41239_41539 , \41238_41538 );
buf \U$33124 ( \41240_41540 , \41239_41539 );
xor \U$33125 ( \41241_41541 , \41234_41534 , \41240_41540 );
and \U$33126 ( \41242_41542 , \18908_18702 , \36686_36986_nG9b90 );
and \U$33127 ( \41243_41543 , \18400_18699 , \36950_37250_nG9b8d );
or \U$33128 ( \41244_41544 , \41242_41542 , \41243_41543 );
xor \U$33129 ( \41245_41545 , \18399_18698 , \41244_41544 );
buf \U$33130 ( \41246_41546 , \41245_41545 );
buf \U$33132 ( \41247_41547 , \41246_41546 );
xor \U$33133 ( \41248_41548 , \41241_41541 , \41247_41547 );
buf \U$33134 ( \41249_41549 , \41248_41548 );
and \U$33135 ( \41250_41550 , \40894_41194 , \40900_41200 );
and \U$33136 ( \41251_41551 , \40894_41194 , \40907_41207 );
and \U$33137 ( \41252_41552 , \40900_41200 , \40907_41207 );
or \U$33138 ( \41253_41553 , \41250_41550 , \41251_41551 , \41252_41552 );
buf \U$33139 ( \41254_41554 , \41253_41553 );
xor \U$33140 ( \41255_41555 , \41249_41549 , \41254_41554 );
and \U$33141 ( \41256_41556 , \41022_41322 , \41028_41328 );
and \U$33142 ( \41257_41557 , \41022_41322 , \41086_41386 );
and \U$33143 ( \41258_41558 , \41028_41328 , \41086_41386 );
or \U$33144 ( \41259_41559 , \41256_41556 , \41257_41557 , \41258_41558 );
buf \U$33145 ( \41260_41560 , \41259_41559 );
xor \U$33146 ( \41261_41561 , \41255_41555 , \41260_41560 );
buf \U$33147 ( \41262_41562 , \41261_41561 );
and \U$33148 ( \41263_41563 , \41107_41407 , \41112_41412 );
and \U$33149 ( \41264_41564 , \41107_41407 , \41141_41441 );
and \U$33150 ( \41265_41565 , \41112_41412 , \41141_41441 );
or \U$33151 ( \41266_41566 , \41263_41563 , \41264_41564 , \41265_41565 );
buf \U$33152 ( \41267_41567 , \41266_41566 );
xor \U$33153 ( \41268_41568 , \41262_41562 , \41267_41567 );
and \U$33154 ( \41269_41569 , \41118_41418 , \41124_41424 );
buf \U$33155 ( \41270_41570 , \41269_41569 );
and \U$33156 ( \41271_41571 , \31989_31636 , \28300_28602_nG9bc0 );
and \U$33157 ( \41272_41572 , \31334_31633 , \28877_29179_nG9bbd );
or \U$33158 ( \41273_41573 , \41271_41571 , \41272_41572 );
xor \U$33159 ( \41274_41574 , \31333_31632 , \41273_41573 );
buf \U$33160 ( \41275_41575 , \41274_41574 );
buf \U$33162 ( \41276_41576 , \41275_41575 );
xor \U$33163 ( \41277_41577 , \41270_41570 , \41276_41576 );
and \U$33164 ( \41278_41578 , \27141_26431 , \32881_33181_nG9bae );
and \U$33165 ( \41279_41579 , \26129_26428 , \33313_33613_nG9bab );
or \U$33166 ( \41280_41580 , \41278_41578 , \41279_41579 );
xor \U$33167 ( \41281_41581 , \26128_26427 , \41280_41580 );
buf \U$33168 ( \41282_41582 , \41281_41581 );
buf \U$33170 ( \41283_41583 , \41282_41582 );
xor \U$33171 ( \41284_41584 , \41277_41577 , \41283_41583 );
buf \U$33172 ( \41285_41585 , \41284_41584 );
and \U$33173 ( \41286_41586 , \41126_41426 , \41132_41432 );
and \U$33174 ( \41287_41587 , \41126_41426 , \41139_41439 );
and \U$33175 ( \41288_41588 , \41132_41432 , \41139_41439 );
or \U$33176 ( \41289_41589 , \41286_41586 , \41287_41587 , \41288_41588 );
buf \U$33177 ( \41290_41590 , \41289_41589 );
xor \U$33178 ( \41291_41591 , \41285_41585 , \41290_41590 );
and \U$33179 ( \41292_41592 , \40921_41221 , \40927_41227 );
and \U$33180 ( \41293_41593 , \40921_41221 , \40934_41234 );
and \U$33181 ( \41294_41594 , \40927_41227 , \40934_41234 );
or \U$33182 ( \41295_41595 , \41292_41592 , \41293_41593 , \41294_41594 );
buf \U$33183 ( \41296_41596 , \41295_41595 );
xor \U$33184 ( \41297_41597 , \41291_41591 , \41296_41596 );
buf \U$33185 ( \41298_41598 , \41297_41597 );
xor \U$33186 ( \41299_41599 , \41268_41568 , \41298_41598 );
buf \U$33187 ( \41300_41600 , \41299_41599 );
and \U$33188 ( \41301_41601 , \41096_41396 , \41101_41401 );
and \U$33189 ( \41302_41602 , \41096_41396 , \41143_41443 );
and \U$33190 ( \41303_41603 , \41101_41401 , \41143_41443 );
or \U$33191 ( \41304_41604 , \41301_41601 , \41302_41602 , \41303_41603 );
buf \U$33192 ( \41305_41605 , \41304_41604 );
xor \U$33193 ( \41306_41606 , \41300_41600 , \41305_41605 );
and \U$33194 ( \41307_41607 , \40967_41267 , \40973_41273 );
and \U$33195 ( \41308_41608 , \40967_41267 , \40980_41280 );
and \U$33196 ( \41309_41609 , \40973_41273 , \40980_41280 );
or \U$33197 ( \41310_41610 , \41307_41607 , \41308_41608 , \41309_41609 );
buf \U$33198 ( \41311_41611 , \41310_41610 );
and \U$33199 ( \41312_41612 , \17437_17297 , \37307_37607_nG9b8a );
and \U$33200 ( \41313_41613 , \16995_17294 , \37674_37974_nG9b87 );
or \U$33201 ( \41314_41614 , \41312_41612 , \41313_41613 );
xor \U$33202 ( \41315_41615 , \16994_17293 , \41314_41614 );
buf \U$33203 ( \41316_41616 , \41315_41615 );
buf \U$33205 ( \41317_41617 , \41316_41616 );
xor \U$33206 ( \41318_41618 , \41311_41611 , \41317_41617 );
and \U$33207 ( \41319_41619 , \12183_12157 , \39904_40204_nG9b72 );
and \U$33208 ( \41320_41620 , \11855_12154 , \40152_40452_nG9b6f );
or \U$33209 ( \41321_41621 , \41319_41619 , \41320_41620 );
xor \U$33210 ( \41322_41622 , \11854_12153 , \41321_41621 );
buf \U$33211 ( \41323_41623 , \41322_41622 );
buf \U$33213 ( \41324_41624 , \41323_41623 );
xor \U$33214 ( \41325_41625 , \41318_41618 , \41324_41624 );
buf \U$33215 ( \41326_41626 , \41325_41625 );
and \U$33216 ( \41327_41627 , \20353_20155 , \35872_36172_nG9b96 );
and \U$33217 ( \41328_41628 , \19853_20152 , \36289_36589_nG9b93 );
or \U$33218 ( \41329_41629 , \41327_41627 , \41328_41628 );
xor \U$33219 ( \41330_41630 , \19852_20151 , \41329_41629 );
buf \U$33220 ( \41331_41631 , \41330_41630 );
buf \U$33222 ( \41332_41632 , \41331_41631 );
and \U$33223 ( \41333_41633 , \13431_13370 , \39291_39591_nG9b78 );
and \U$33224 ( \41334_41634 , \13068_13367 , \39663_39963_nG9b75 );
or \U$33225 ( \41335_41635 , \41333_41633 , \41334_41634 );
xor \U$33226 ( \41336_41636 , \13067_13366 , \41335_41635 );
buf \U$33227 ( \41337_41637 , \41336_41636 );
buf \U$33229 ( \41338_41638 , \41337_41637 );
xor \U$33230 ( \41339_41639 , \41332_41632 , \41338_41638 );
and \U$33231 ( \41340_41640 , \10411_10707 , \41081_41381_nG9b66 );
and \U$33232 ( \41341_41641 , \41034_41334 , \41038_41338 );
and \U$33233 ( \41342_41642 , \41038_41338 , \41070_41370 );
and \U$33234 ( \41343_41643 , \41034_41334 , \41070_41370 );
or \U$33235 ( \41344_41644 , \41341_41641 , \41342_41642 , \41343_41643 );
and \U$33236 ( \41345_41645 , \41058_41358 , \41063_41363 );
and \U$33237 ( \41346_41646 , \41063_41363 , \41068_41368 );
and \U$33238 ( \41347_41647 , \41058_41358 , \41068_41368 );
or \U$33239 ( \41348_41648 , \41345_41645 , \41346_41646 , \41347_41647 );
and \U$33240 ( \41349_41649 , \41043_41343 , \41053_41353 );
and \U$33241 ( \41350_41650 , \41053_41353 , \41069_41369 );
and \U$33242 ( \41351_41651 , \41043_41343 , \41069_41369 );
or \U$33243 ( \41352_41652 , \41349_41649 , \41350_41650 , \41351_41651 );
xor \U$33244 ( \41353_41653 , \41348_41648 , \41352_41652 );
and \U$33245 ( \41354_41654 , \41046_41346 , \41050_41350 );
and \U$33246 ( \41355_41655 , \41050_41350 , \41052_41352 );
and \U$33247 ( \41356_41656 , \41046_41346 , \41052_41352 );
or \U$33248 ( \41357_41657 , \41354_41654 , \41355_41655 , \41356_41656 );
not \U$33249 ( \41358_41658 , \26993_27295 );
and \U$33250 ( \41359_41659 , \31752_32054 , \28768_29070 );
and \U$33251 ( \41360_41660 , \32495_32794 , \28224_28526 );
nor \U$33252 ( \41361_41661 , \41359_41659 , \41360_41660 );
xnor \U$33253 ( \41362_41662 , \41361_41661 , \28774_29076 );
xor \U$33254 ( \41363_41663 , \41358_41658 , \41362_41662 );
and \U$33255 ( \41364_41664 , \28232_28534 , \32555_32854 );
and \U$33256 ( \41365_41665 , \28782_29084 , \31765_32067 );
nor \U$33257 ( \41366_41666 , \41364_41664 , \41365_41665 );
xnor \U$33258 ( \41367_41667 , \41366_41666 , \32506_32805 );
xor \U$33259 ( \41368_41668 , \41363_41663 , \41367_41667 );
xor \U$33260 ( \41369_41669 , \41357_41657 , \41368_41668 );
buf \U$33261 ( \41370_41670 , \41062_41362 );
and \U$33262 ( \41371_41671 , \29966_30268 , \30521_30823 );
and \U$33263 ( \41372_41672 , \30500_30802 , \29944_30246 );
nor \U$33264 ( \41373_41673 , \41371_41671 , \41372_41672 );
xnor \U$33265 ( \41374_41674 , \41373_41673 , \30511_30813 );
xor \U$33266 ( \41375_41675 , \41370_41670 , \41374_41674 );
and \U$33267 ( \41376_41676 , \27011_27313 , \32503_32802 );
xor \U$33268 ( \41377_41677 , \41375_41675 , \41376_41676 );
xor \U$33269 ( \41378_41678 , \41369_41669 , \41377_41677 );
xor \U$33270 ( \41379_41679 , \41353_41653 , \41378_41678 );
xor \U$33271 ( \41380_41680 , \41344_41644 , \41379_41679 );
and \U$33272 ( \41381_41681 , \41071_41371 , \41075_41375 );
and \U$33273 ( \41382_41682 , \41076_41376 , \41079_41379 );
or \U$33274 ( \41383_41683 , \41381_41681 , \41382_41682 );
xor \U$33275 ( \41384_41684 , \41380_41680 , \41383_41683 );
buf g9b63_GF_PartitionCandidate( \41385_41685_nG9b63 , \41384_41684 );
and \U$33276 ( \41386_41686 , \10402_10704 , \41385_41685_nG9b63 );
or \U$33277 ( \41387_41687 , \41340_41640 , \41386_41686 );
xor \U$33278 ( \41388_41688 , \10399_10703 , \41387_41687 );
buf \U$33279 ( \41389_41689 , \41388_41688 );
buf \U$33281 ( \41390_41690 , \41389_41689 );
xor \U$33282 ( \41391_41691 , \41339_41639 , \41390_41690 );
buf \U$33283 ( \41392_41692 , \41391_41691 );
xor \U$33284 ( \41393_41693 , \41326_41626 , \41392_41692 );
and \U$33286 ( \41394_41694 , \32617_32916 , \27114_27416_nG9bc3 );
or \U$33287 ( \41395_41695 , 1'b0 , \41394_41694 );
xor \U$33288 ( \41396_41696 , 1'b0 , \41395_41695 );
buf \U$33289 ( \41397_41697 , \41396_41696 );
buf \U$33291 ( \41398_41698 , \41397_41697 );
and \U$33292 ( \41399_41699 , \30670_29853 , \30064_30366_nG9bba );
and \U$33293 ( \41400_41700 , \29551_29850 , \30638_30940_nG9bb7 );
or \U$33294 ( \41401_41701 , \41399_41699 , \41400_41700 );
xor \U$33295 ( \41402_41702 , \29550_29849 , \41401_41701 );
buf \U$33296 ( \41403_41703 , \41402_41702 );
buf \U$33298 ( \41404_41704 , \41403_41703 );
xor \U$33299 ( \41405_41705 , \41398_41698 , \41404_41704 );
buf \U$33300 ( \41406_41706 , \41405_41705 );
and \U$33301 ( \41407_41707 , \28946_28118 , \31877_32179_nG9bb4 );
and \U$33302 ( \41408_41708 , \27816_28115 , \32589_32888_nG9bb1 );
or \U$33303 ( \41409_41709 , \41407_41707 , \41408_41708 );
xor \U$33304 ( \41410_41710 , \27815_28114 , \41409_41709 );
buf \U$33305 ( \41411_41711 , \41410_41710 );
buf \U$33307 ( \41412_41712 , \41411_41711 );
xor \U$33308 ( \41413_41713 , \41406_41706 , \41412_41712 );
and \U$33309 ( \41414_41714 , \23495_23201 , \34343_34643_nG9ba2 );
and \U$33310 ( \41415_41715 , \22899_23198 , \34794_35094_nG9b9f );
or \U$33311 ( \41416_41716 , \41414_41714 , \41415_41715 );
xor \U$33312 ( \41417_41717 , \22898_23197 , \41416_41716 );
buf \U$33313 ( \41418_41718 , \41417_41717 );
buf \U$33315 ( \41419_41719 , \41418_41718 );
xor \U$33316 ( \41420_41720 , \41413_41713 , \41419_41719 );
buf \U$33317 ( \41421_41721 , \41420_41720 );
xor \U$33318 ( \41422_41722 , \41393_41693 , \41421_41721 );
buf \U$33319 ( \41423_41723 , \41422_41722 );
xor \U$33320 ( \41424_41724 , \41306_41606 , \41423_41723 );
buf \U$33321 ( \41425_41725 , \41424_41724 );
xor \U$33322 ( \41426_41726 , \41228_41528 , \41425_41725 );
and \U$33323 ( \41427_41727 , \41162_41462 , \41426_41726 );
and \U$33325 ( \41428_41728 , \41156_41456 , \41161_41461 );
or \U$33327 ( \41429_41729 , 1'b0 , \41428_41728 , 1'b0 );
xor \U$33328 ( \41430_41730 , \41427_41727 , \41429_41729 );
and \U$33330 ( \41431_41731 , \41149_41449 , \41155_41455 );
and \U$33331 ( \41432_41732 , \41151_41451 , \41155_41455 );
or \U$33332 ( \41433_41733 , 1'b0 , \41431_41731 , \41432_41732 );
xor \U$33333 ( \41434_41734 , \41430_41730 , \41433_41733 );
xor \U$33340 ( \41435_41735 , \41434_41734 , 1'b0 );
and \U$33341 ( \41436_41736 , \41222_41522 , \41227_41527 );
and \U$33342 ( \41437_41737 , \41222_41522 , \41425_41725 );
and \U$33343 ( \41438_41738 , \41227_41527 , \41425_41725 );
or \U$33344 ( \41439_41739 , \41436_41736 , \41437_41737 , \41438_41738 );
xor \U$33345 ( \41440_41740 , \41435_41735 , \41439_41739 );
and \U$33346 ( \41441_41741 , \41167_41467 , \41172_41472 );
and \U$33347 ( \41442_41742 , \41167_41467 , \41220_41520 );
and \U$33348 ( \41443_41743 , \41172_41472 , \41220_41520 );
or \U$33349 ( \41444_41744 , \41441_41741 , \41442_41742 , \41443_41743 );
buf \U$33350 ( \41445_41745 , \41444_41744 );
and \U$33351 ( \41446_41746 , \41300_41600 , \41305_41605 );
and \U$33352 ( \41447_41747 , \41300_41600 , \41423_41723 );
and \U$33353 ( \41448_41748 , \41305_41605 , \41423_41723 );
or \U$33354 ( \41449_41749 , \41446_41746 , \41447_41747 , \41448_41748 );
buf \U$33355 ( \41450_41750 , \41449_41749 );
and \U$33356 ( \41451_41751 , \41285_41585 , \41290_41590 );
and \U$33357 ( \41452_41752 , \41285_41585 , \41296_41596 );
and \U$33358 ( \41453_41753 , \41290_41590 , \41296_41596 );
or \U$33359 ( \41454_41754 , \41451_41751 , \41452_41752 , \41453_41753 );
buf \U$33360 ( \41455_41755 , \41454_41754 );
and \U$33361 ( \41456_41756 , \16405_15940 , \38363_38663_nG9b81 );
and \U$33362 ( \41457_41757 , \15638_15937 , \38668_38968_nG9b7e );
or \U$33363 ( \41458_41758 , \41456_41756 , \41457_41757 );
xor \U$33364 ( \41459_41759 , \15637_15936 , \41458_41758 );
buf \U$33365 ( \41460_41760 , \41459_41759 );
buf \U$33367 ( \41461_41761 , \41460_41760 );
and \U$33368 ( \41462_41762 , \14710_14631 , \39034_39334_nG9b7b );
and \U$33369 ( \41463_41763 , \14329_14628 , \39291_39591_nG9b78 );
or \U$33370 ( \41464_41764 , \41462_41762 , \41463_41763 );
xor \U$33371 ( \41465_41765 , \14328_14627 , \41464_41764 );
buf \U$33372 ( \41466_41766 , \41465_41765 );
buf \U$33374 ( \41467_41767 , \41466_41766 );
xor \U$33375 ( \41468_41768 , \41461_41761 , \41467_41767 );
and \U$33376 ( \41469_41769 , \10996_10421 , \40740_41040_nG9b69 );
and \U$33377 ( \41470_41770 , \10119_10418 , \41081_41381_nG9b66 );
or \U$33378 ( \41471_41771 , \41469_41769 , \41470_41770 );
xor \U$33379 ( \41472_41772 , \10118_10417 , \41471_41771 );
buf \U$33380 ( \41473_41773 , \41472_41772 );
buf \U$33382 ( \41474_41774 , \41473_41773 );
xor \U$33383 ( \41475_41775 , \41468_41768 , \41474_41774 );
buf \U$33384 ( \41476_41776 , \41475_41775 );
xor \U$33385 ( \41477_41777 , \41455_41755 , \41476_41776 );
and \U$33386 ( \41478_41778 , \41311_41611 , \41317_41617 );
and \U$33387 ( \41479_41779 , \41311_41611 , \41324_41624 );
and \U$33388 ( \41480_41780 , \41317_41617 , \41324_41624 );
or \U$33389 ( \41481_41781 , \41478_41778 , \41479_41779 , \41480_41780 );
buf \U$33390 ( \41482_41782 , \41481_41781 );
xor \U$33391 ( \41483_41783 , \41477_41777 , \41482_41782 );
buf \U$33392 ( \41484_41784 , \41483_41783 );
and \U$33393 ( \41485_41785 , \41199_41499 , \41204_41504 );
and \U$33394 ( \41486_41786 , \41199_41499 , \41210_41510 );
and \U$33395 ( \41487_41787 , \41204_41504 , \41210_41510 );
or \U$33396 ( \41488_41788 , \41485_41785 , \41486_41786 , \41487_41787 );
buf \U$33397 ( \41489_41789 , \41488_41788 );
xor \U$33398 ( \41490_41790 , \41484_41784 , \41489_41789 );
and \U$33399 ( \41491_41791 , \41326_41626 , \41392_41692 );
and \U$33400 ( \41492_41792 , \41326_41626 , \41421_41721 );
and \U$33401 ( \41493_41793 , \41392_41692 , \41421_41721 );
or \U$33402 ( \41494_41794 , \41491_41791 , \41492_41792 , \41493_41793 );
buf \U$33403 ( \41495_41795 , \41494_41794 );
xor \U$33404 ( \41496_41796 , \41490_41790 , \41495_41795 );
buf \U$33405 ( \41497_41797 , \41496_41796 );
xor \U$33406 ( \41498_41798 , \41450_41750 , \41497_41797 );
and \U$33407 ( \41499_41799 , \41178_41478 , \41212_41512 );
and \U$33408 ( \41500_41800 , \41178_41478 , \41218_41518 );
and \U$33409 ( \41501_41801 , \41212_41512 , \41218_41518 );
or \U$33410 ( \41502_41802 , \41499_41799 , \41500_41800 , \41501_41801 );
buf \U$33411 ( \41503_41803 , \41502_41802 );
xor \U$33412 ( \41504_41804 , \41498_41798 , \41503_41803 );
buf \U$33413 ( \41505_41805 , \41504_41804 );
xor \U$33414 ( \41506_41806 , \41445_41745 , \41505_41805 );
and \U$33415 ( \41507_41807 , \41262_41562 , \41267_41567 );
and \U$33416 ( \41508_41808 , \41262_41562 , \41298_41598 );
and \U$33417 ( \41509_41809 , \41267_41567 , \41298_41598 );
or \U$33418 ( \41510_41810 , \41507_41807 , \41508_41808 , \41509_41809 );
buf \U$33419 ( \41511_41811 , \41510_41810 );
and \U$33420 ( \41512_41812 , \41249_41549 , \41254_41554 );
and \U$33421 ( \41513_41813 , \41249_41549 , \41260_41560 );
and \U$33422 ( \41514_41814 , \41254_41554 , \41260_41560 );
or \U$33423 ( \41515_41815 , \41512_41812 , \41513_41813 , \41514_41814 );
buf \U$33424 ( \41516_41816 , \41515_41815 );
and \U$33425 ( \41517_41817 , \41234_41534 , \41240_41540 );
and \U$33426 ( \41518_41818 , \41234_41534 , \41247_41547 );
and \U$33427 ( \41519_41819 , \41240_41540 , \41247_41547 );
or \U$33428 ( \41520_41820 , \41517_41817 , \41518_41818 , \41519_41819 );
buf \U$33429 ( \41521_41821 , \41520_41820 );
and \U$33430 ( \41522_41822 , \41406_41706 , \41412_41712 );
and \U$33431 ( \41523_41823 , \41406_41706 , \41419_41719 );
and \U$33432 ( \41524_41824 , \41412_41712 , \41419_41719 );
or \U$33433 ( \41525_41825 , \41522_41822 , \41523_41823 , \41524_41824 );
buf \U$33434 ( \41526_41826 , \41525_41825 );
xor \U$33435 ( \41527_41827 , \41521_41821 , \41526_41826 );
and \U$33436 ( \41528_41828 , \31989_31636 , \28877_29179_nG9bbd );
and \U$33437 ( \41529_41829 , \31334_31633 , \30064_30366_nG9bba );
or \U$33438 ( \41530_41830 , \41528_41828 , \41529_41829 );
xor \U$33439 ( \41531_41831 , \31333_31632 , \41530_41830 );
buf \U$33440 ( \41532_41832 , \41531_41831 );
buf \U$33442 ( \41533_41833 , \41532_41832 );
and \U$33443 ( \41534_41834 , \28946_28118 , \32589_32888_nG9bb1 );
and \U$33444 ( \41535_41835 , \27816_28115 , \32881_33181_nG9bae );
or \U$33445 ( \41536_41836 , \41534_41834 , \41535_41835 );
xor \U$33446 ( \41537_41837 , \27815_28114 , \41536_41836 );
buf \U$33447 ( \41538_41838 , \41537_41837 );
buf \U$33449 ( \41539_41839 , \41538_41838 );
xor \U$33450 ( \41540_41840 , \41533_41833 , \41539_41839 );
and \U$33451 ( \41541_41841 , \27141_26431 , \33313_33613_nG9bab );
and \U$33452 ( \41542_41842 , \26129_26428 , \33741_34041_nG9ba8 );
or \U$33453 ( \41543_41843 , \41541_41841 , \41542_41842 );
xor \U$33454 ( \41544_41844 , \26128_26427 , \41543_41843 );
buf \U$33455 ( \41545_41845 , \41544_41844 );
buf \U$33457 ( \41546_41846 , \41545_41845 );
xor \U$33458 ( \41547_41847 , \41540_41840 , \41546_41846 );
buf \U$33459 ( \41548_41848 , \41547_41847 );
xor \U$33460 ( \41549_41849 , \41527_41827 , \41548_41848 );
buf \U$33461 ( \41550_41850 , \41549_41849 );
xor \U$33462 ( \41551_41851 , \41516_41816 , \41550_41850 );
and \U$33463 ( \41552_41852 , \41332_41632 , \41338_41638 );
and \U$33464 ( \41553_41853 , \41332_41632 , \41390_41690 );
and \U$33465 ( \41554_41854 , \41338_41638 , \41390_41690 );
or \U$33466 ( \41555_41855 , \41552_41852 , \41553_41853 , \41554_41854 );
buf \U$33467 ( \41556_41856 , \41555_41855 );
and \U$33468 ( \41557_41857 , \41184_41484 , \41190_41490 );
and \U$33469 ( \41558_41858 , \41184_41484 , \41197_41497 );
and \U$33470 ( \41559_41859 , \41190_41490 , \41197_41497 );
or \U$33471 ( \41560_41860 , \41557_41857 , \41558_41858 , \41559_41859 );
buf \U$33472 ( \41561_41861 , \41560_41860 );
xor \U$33473 ( \41562_41862 , \41556_41856 , \41561_41861 );
and \U$33474 ( \41563_41863 , \25044_24792 , \33994_34294_nG9ba5 );
and \U$33475 ( \41564_41864 , \24490_24789 , \34343_34643_nG9ba2 );
or \U$33476 ( \41565_41865 , \41563_41863 , \41564_41864 );
xor \U$33477 ( \41566_41866 , \24489_24788 , \41565_41865 );
buf \U$33478 ( \41567_41867 , \41566_41866 );
buf \U$33480 ( \41568_41868 , \41567_41867 );
and \U$33481 ( \41569_41869 , \21908_21658 , \35501_35801_nG9b99 );
and \U$33482 ( \41570_41870 , \21356_21655 , \35872_36172_nG9b96 );
or \U$33483 ( \41571_41871 , \41569_41869 , \41570_41870 );
xor \U$33484 ( \41572_41872 , \21355_21654 , \41571_41871 );
buf \U$33485 ( \41573_41873 , \41572_41872 );
buf \U$33487 ( \41574_41874 , \41573_41873 );
xor \U$33488 ( \41575_41875 , \41568_41868 , \41574_41874 );
and \U$33489 ( \41576_41876 , \18908_18702 , \36950_37250_nG9b8d );
and \U$33490 ( \41577_41877 , \18400_18699 , \37307_37607_nG9b8a );
or \U$33491 ( \41578_41878 , \41576_41876 , \41577_41877 );
xor \U$33492 ( \41579_41879 , \18399_18698 , \41578_41878 );
buf \U$33493 ( \41580_41880 , \41579_41879 );
buf \U$33495 ( \41581_41881 , \41580_41880 );
xor \U$33496 ( \41582_41882 , \41575_41875 , \41581_41881 );
buf \U$33497 ( \41583_41883 , \41582_41882 );
xor \U$33498 ( \41584_41884 , \41562_41862 , \41583_41883 );
buf \U$33499 ( \41585_41885 , \41584_41884 );
xor \U$33500 ( \41586_41886 , \41551_41851 , \41585_41885 );
buf \U$33501 ( \41587_41887 , \41586_41886 );
xor \U$33502 ( \41588_41888 , \41511_41811 , \41587_41887 );
and \U$33503 ( \41589_41889 , \41270_41570 , \41276_41576 );
and \U$33504 ( \41590_41890 , \41270_41570 , \41283_41583 );
and \U$33505 ( \41591_41891 , \41276_41576 , \41283_41583 );
or \U$33506 ( \41592_41892 , \41589_41889 , \41590_41890 , \41591_41891 );
buf \U$33507 ( \41593_41893 , \41592_41892 );
and \U$33508 ( \41594_41894 , \17437_17297 , \37674_37974_nG9b87 );
and \U$33509 ( \41595_41895 , \16995_17294 , \38037_38337_nG9b84 );
or \U$33510 ( \41596_41896 , \41594_41894 , \41595_41895 );
xor \U$33511 ( \41597_41897 , \16994_17293 , \41596_41896 );
buf \U$33512 ( \41598_41898 , \41597_41897 );
buf \U$33514 ( \41599_41899 , \41598_41898 );
xor \U$33515 ( \41600_41900 , \41593_41893 , \41599_41899 );
and \U$33516 ( \41601_41901 , \12183_12157 , \40152_40452_nG9b6f );
and \U$33517 ( \41602_41902 , \11855_12154 , \40543_40843_nG9b6c );
or \U$33518 ( \41603_41903 , \41601_41901 , \41602_41902 );
xor \U$33519 ( \41604_41904 , \11854_12153 , \41603_41903 );
buf \U$33520 ( \41605_41905 , \41604_41904 );
buf \U$33522 ( \41606_41906 , \41605_41905 );
xor \U$33523 ( \41607_41907 , \41600_41900 , \41606_41906 );
buf \U$33524 ( \41608_41908 , \41607_41907 );
and \U$33525 ( \41609_41909 , \20353_20155 , \36289_36589_nG9b93 );
and \U$33526 ( \41610_41910 , \19853_20152 , \36686_36986_nG9b90 );
or \U$33527 ( \41611_41911 , \41609_41909 , \41610_41910 );
xor \U$33528 ( \41612_41912 , \19852_20151 , \41611_41911 );
buf \U$33529 ( \41613_41913 , \41612_41912 );
buf \U$33531 ( \41614_41914 , \41613_41913 );
and \U$33532 ( \41615_41915 , \13431_13370 , \39663_39963_nG9b75 );
and \U$33533 ( \41616_41916 , \13068_13367 , \39904_40204_nG9b72 );
or \U$33534 ( \41617_41917 , \41615_41915 , \41616_41916 );
xor \U$33535 ( \41618_41918 , \13067_13366 , \41617_41917 );
buf \U$33536 ( \41619_41919 , \41618_41918 );
buf \U$33538 ( \41620_41920 , \41619_41919 );
xor \U$33539 ( \41621_41921 , \41614_41914 , \41620_41920 );
and \U$33540 ( \41622_41922 , \10411_10707 , \41385_41685_nG9b63 );
and \U$33541 ( \41623_41923 , \41370_41670 , \41374_41674 );
and \U$33542 ( \41624_41924 , \41374_41674 , \41376_41676 );
and \U$33543 ( \41625_41925 , \41370_41670 , \41376_41676 );
or \U$33544 ( \41626_41926 , \41623_41923 , \41624_41924 , \41625_41925 );
and \U$33545 ( \41627_41927 , \41357_41657 , \41368_41668 );
and \U$33546 ( \41628_41928 , \41368_41668 , \41377_41677 );
and \U$33547 ( \41629_41929 , \41357_41657 , \41377_41677 );
or \U$33548 ( \41630_41930 , \41627_41927 , \41628_41928 , \41629_41929 );
xor \U$33549 ( \41631_41931 , \41626_41926 , \41630_41930 );
and \U$33550 ( \41632_41932 , \41358_41658 , \41362_41662 );
and \U$33551 ( \41633_41933 , \41362_41662 , \41367_41667 );
and \U$33552 ( \41634_41934 , \41358_41658 , \41367_41667 );
or \U$33553 ( \41635_41935 , \41632_41932 , \41633_41933 , \41634_41934 );
and \U$33554 ( \41636_41936 , \32495_32794 , \28768_29070 );
not \U$33555 ( \41637_41937 , \41636_41936 );
xnor \U$33556 ( \41638_41938 , \41637_41937 , \28774_29076 );
not \U$33557 ( \41639_41939 , \41638_41938 );
xor \U$33558 ( \41640_41940 , \41635_41935 , \41639_41939 );
and \U$33559 ( \41641_41941 , \30500_30802 , \30521_30823 );
and \U$33560 ( \41642_41942 , \31752_32054 , \29944_30246 );
nor \U$33561 ( \41643_41943 , \41641_41941 , \41642_41942 );
xnor \U$33562 ( \41644_41944 , \41643_41943 , \30511_30813 );
and \U$33563 ( \41645_41945 , \28782_29084 , \32555_32854 );
and \U$33564 ( \41646_41946 , \29966_30268 , \31765_32067 );
nor \U$33565 ( \41647_41947 , \41645_41945 , \41646_41946 );
xnor \U$33566 ( \41648_41948 , \41647_41947 , \32506_32805 );
xor \U$33567 ( \41649_41949 , \41644_41944 , \41648_41948 );
and \U$33568 ( \41650_41950 , \28232_28534 , \32503_32802 );
xor \U$33569 ( \41651_41951 , \41649_41949 , \41650_41950 );
xor \U$33570 ( \41652_41952 , \41640_41940 , \41651_41951 );
xor \U$33571 ( \41653_41953 , \41631_41931 , \41652_41952 );
and \U$33572 ( \41654_41954 , \41348_41648 , \41352_41652 );
and \U$33573 ( \41655_41955 , \41352_41652 , \41378_41678 );
and \U$33574 ( \41656_41956 , \41348_41648 , \41378_41678 );
or \U$33575 ( \41657_41957 , \41654_41954 , \41655_41955 , \41656_41956 );
xor \U$33576 ( \41658_41958 , \41653_41953 , \41657_41957 );
and \U$33577 ( \41659_41959 , \41344_41644 , \41379_41679 );
and \U$33578 ( \41660_41960 , \41380_41680 , \41383_41683 );
or \U$33579 ( \41661_41961 , \41659_41959 , \41660_41960 );
xor \U$33580 ( \41662_41962 , \41658_41958 , \41661_41961 );
buf g9b60_GF_PartitionCandidate( \41663_41963_nG9b60 , \41662_41962 );
and \U$33581 ( \41664_41964 , \10402_10704 , \41663_41963_nG9b60 );
or \U$33582 ( \41665_41965 , \41622_41922 , \41664_41964 );
xor \U$33583 ( \41666_41966 , \10399_10703 , \41665_41965 );
buf \U$33584 ( \41667_41967 , \41666_41966 );
buf \U$33586 ( \41668_41968 , \41667_41967 );
xor \U$33587 ( \41669_41969 , \41621_41921 , \41668_41968 );
buf \U$33588 ( \41670_41970 , \41669_41969 );
xor \U$33589 ( \41671_41971 , \41608_41908 , \41670_41970 );
and \U$33591 ( \41672_41972 , \32617_32916 , \28300_28602_nG9bc0 );
or \U$33592 ( \41673_41973 , 1'b0 , \41672_41972 );
xor \U$33593 ( \41674_41974 , 1'b0 , \41673_41973 );
buf \U$33594 ( \41675_41975 , \41674_41974 );
buf \U$33596 ( \41676_41976 , \41675_41975 );
and \U$33597 ( \41677_41977 , \30670_29853 , \30638_30940_nG9bb7 );
and \U$33598 ( \41678_41978 , \29551_29850 , \31877_32179_nG9bb4 );
or \U$33599 ( \41679_41979 , \41677_41977 , \41678_41978 );
xor \U$33600 ( \41680_41980 , \29550_29849 , \41679_41979 );
buf \U$33601 ( \41681_41981 , \41680_41980 );
buf \U$33603 ( \41682_41982 , \41681_41981 );
xor \U$33604 ( \41683_41983 , \41676_41976 , \41682_41982 );
buf \U$33605 ( \41684_41984 , \41683_41983 );
and \U$33606 ( \41685_41985 , \41398_41698 , \41404_41704 );
buf \U$33607 ( \41686_41986 , \41685_41985 );
xor \U$33608 ( \41687_41987 , \41684_41984 , \41686_41986 );
and \U$33609 ( \41688_41988 , \23495_23201 , \34794_35094_nG9b9f );
and \U$33610 ( \41689_41989 , \22899_23198 , \35270_35570_nG9b9c );
or \U$33611 ( \41690_41990 , \41688_41988 , \41689_41989 );
xor \U$33612 ( \41691_41991 , \22898_23197 , \41690_41990 );
buf \U$33613 ( \41692_41992 , \41691_41991 );
buf \U$33615 ( \41693_41993 , \41692_41992 );
xor \U$33616 ( \41694_41994 , \41687_41987 , \41693_41993 );
buf \U$33617 ( \41695_41995 , \41694_41994 );
xor \U$33618 ( \41696_41996 , \41671_41971 , \41695_41995 );
buf \U$33619 ( \41697_41997 , \41696_41996 );
xor \U$33620 ( \41698_41998 , \41588_41888 , \41697_41997 );
buf \U$33621 ( \41699_41999 , \41698_41998 );
xor \U$33622 ( \41700_42000 , \41506_41806 , \41699_41999 );
and \U$33623 ( \41701_42001 , \41440_41740 , \41700_42000 );
and \U$33625 ( \41702_42002 , \41434_41734 , \41439_41739 );
or \U$33627 ( \41703_42003 , 1'b0 , \41702_42002 , 1'b0 );
xor \U$33628 ( \41704_42004 , \41701_42001 , \41703_42003 );
and \U$33630 ( \41705_42005 , \41427_41727 , \41433_41733 );
and \U$33631 ( \41706_42006 , \41429_41729 , \41433_41733 );
or \U$33632 ( \41707_42007 , 1'b0 , \41705_42005 , \41706_42006 );
xor \U$33633 ( \41708_42008 , \41704_42004 , \41707_42007 );
xor \U$33640 ( \41709_42009 , \41708_42008 , 1'b0 );
and \U$33641 ( \41710_42010 , \41445_41745 , \41505_41805 );
and \U$33642 ( \41711_42011 , \41445_41745 , \41699_41999 );
and \U$33643 ( \41712_42012 , \41505_41805 , \41699_41999 );
or \U$33644 ( \41713_42013 , \41710_42010 , \41711_42011 , \41712_42012 );
xor \U$33645 ( \41714_42014 , \41709_42009 , \41713_42013 );
and \U$33646 ( \41715_42015 , \41511_41811 , \41587_41887 );
and \U$33647 ( \41716_42016 , \41511_41811 , \41697_41997 );
and \U$33648 ( \41717_42017 , \41587_41887 , \41697_41997 );
or \U$33649 ( \41718_42018 , \41715_42015 , \41716_42016 , \41717_42017 );
buf \U$33650 ( \41719_42019 , \41718_42018 );
and \U$33651 ( \41720_42020 , \41533_41833 , \41539_41839 );
and \U$33652 ( \41721_42021 , \41533_41833 , \41546_41846 );
and \U$33653 ( \41722_42022 , \41539_41839 , \41546_41846 );
or \U$33654 ( \41723_42023 , \41720_42020 , \41721_42021 , \41722_42022 );
buf \U$33655 ( \41724_42024 , \41723_42023 );
and \U$33656 ( \41725_42025 , \17437_17297 , \38037_38337_nG9b84 );
and \U$33657 ( \41726_42026 , \16995_17294 , \38363_38663_nG9b81 );
or \U$33658 ( \41727_42027 , \41725_42025 , \41726_42026 );
xor \U$33659 ( \41728_42028 , \16994_17293 , \41727_42027 );
buf \U$33660 ( \41729_42029 , \41728_42028 );
buf \U$33662 ( \41730_42030 , \41729_42029 );
xor \U$33663 ( \41731_42031 , \41724_42024 , \41730_42030 );
and \U$33664 ( \41732_42032 , \12183_12157 , \40543_40843_nG9b6c );
and \U$33665 ( \41733_42033 , \11855_12154 , \40740_41040_nG9b69 );
or \U$33666 ( \41734_42034 , \41732_42032 , \41733_42033 );
xor \U$33667 ( \41735_42035 , \11854_12153 , \41734_42034 );
buf \U$33668 ( \41736_42036 , \41735_42035 );
buf \U$33670 ( \41737_42037 , \41736_42036 );
xor \U$33671 ( \41738_42038 , \41731_42031 , \41737_42037 );
buf \U$33672 ( \41739_42039 , \41738_42038 );
and \U$33673 ( \41740_42040 , \41593_41893 , \41599_41899 );
and \U$33674 ( \41741_42041 , \41593_41893 , \41606_41906 );
and \U$33675 ( \41742_42042 , \41599_41899 , \41606_41906 );
or \U$33676 ( \41743_42043 , \41740_42040 , \41741_42041 , \41742_42042 );
buf \U$33677 ( \41744_42044 , \41743_42043 );
xor \U$33678 ( \41745_42045 , \41739_42039 , \41744_42044 );
and \U$33679 ( \41746_42046 , \20353_20155 , \36686_36986_nG9b90 );
and \U$33680 ( \41747_42047 , \19853_20152 , \36950_37250_nG9b8d );
or \U$33681 ( \41748_42048 , \41746_42046 , \41747_42047 );
xor \U$33682 ( \41749_42049 , \19852_20151 , \41748_42048 );
buf \U$33683 ( \41750_42050 , \41749_42049 );
buf \U$33685 ( \41751_42051 , \41750_42050 );
and \U$33686 ( \41752_42052 , \13431_13370 , \39904_40204_nG9b72 );
and \U$33687 ( \41753_42053 , \13068_13367 , \40152_40452_nG9b6f );
or \U$33688 ( \41754_42054 , \41752_42052 , \41753_42053 );
xor \U$33689 ( \41755_42055 , \13067_13366 , \41754_42054 );
buf \U$33690 ( \41756_42056 , \41755_42055 );
buf \U$33692 ( \41757_42057 , \41756_42056 );
xor \U$33693 ( \41758_42058 , \41751_42051 , \41757_42057 );
and \U$33694 ( \41759_42059 , \10996_10421 , \41081_41381_nG9b66 );
and \U$33695 ( \41760_42060 , \10119_10418 , \41385_41685_nG9b63 );
or \U$33696 ( \41761_42061 , \41759_42059 , \41760_42060 );
xor \U$33697 ( \41762_42062 , \10118_10417 , \41761_42061 );
buf \U$33698 ( \41763_42063 , \41762_42062 );
buf \U$33700 ( \41764_42064 , \41763_42063 );
xor \U$33701 ( \41765_42065 , \41758_42058 , \41764_42064 );
buf \U$33702 ( \41766_42066 , \41765_42065 );
xor \U$33703 ( \41767_42067 , \41745_42045 , \41766_42066 );
buf \U$33704 ( \41768_42068 , \41767_42067 );
and \U$33705 ( \41769_42069 , \41455_41755 , \41476_41776 );
and \U$33706 ( \41770_42070 , \41455_41755 , \41482_41782 );
and \U$33707 ( \41771_42071 , \41476_41776 , \41482_41782 );
or \U$33708 ( \41772_42072 , \41769_42069 , \41770_42070 , \41771_42071 );
buf \U$33709 ( \41773_42073 , \41772_42072 );
xor \U$33710 ( \41774_42074 , \41768_42068 , \41773_42073 );
and \U$33711 ( \41775_42075 , \41608_41908 , \41670_41970 );
and \U$33712 ( \41776_42076 , \41608_41908 , \41695_41995 );
and \U$33713 ( \41777_42077 , \41670_41970 , \41695_41995 );
or \U$33714 ( \41778_42078 , \41775_42075 , \41776_42076 , \41777_42077 );
buf \U$33715 ( \41779_42079 , \41778_42078 );
xor \U$33716 ( \41780_42080 , \41774_42074 , \41779_42079 );
buf \U$33717 ( \41781_42081 , \41780_42080 );
xor \U$33718 ( \41782_42082 , \41719_42019 , \41781_42081 );
and \U$33719 ( \41783_42083 , \41484_41784 , \41489_41789 );
and \U$33720 ( \41784_42084 , \41484_41784 , \41495_41795 );
and \U$33721 ( \41785_42085 , \41489_41789 , \41495_41795 );
or \U$33722 ( \41786_42086 , \41783_42083 , \41784_42084 , \41785_42085 );
buf \U$33723 ( \41787_42087 , \41786_42086 );
xor \U$33724 ( \41788_42088 , \41782_42082 , \41787_42087 );
buf \U$33725 ( \41789_42089 , \41788_42088 );
and \U$33726 ( \41790_42090 , \41450_41750 , \41497_41797 );
and \U$33727 ( \41791_42091 , \41450_41750 , \41503_41803 );
and \U$33728 ( \41792_42092 , \41497_41797 , \41503_41803 );
or \U$33729 ( \41793_42093 , \41790_42090 , \41791_42091 , \41792_42092 );
buf \U$33730 ( \41794_42094 , \41793_42093 );
xor \U$33731 ( \41795_42095 , \41789_42089 , \41794_42094 );
and \U$33732 ( \41796_42096 , \41516_41816 , \41550_41850 );
and \U$33733 ( \41797_42097 , \41516_41816 , \41585_41885 );
and \U$33734 ( \41798_42098 , \41550_41850 , \41585_41885 );
or \U$33735 ( \41799_42099 , \41796_42096 , \41797_42097 , \41798_42098 );
buf \U$33736 ( \41800_42100 , \41799_42099 );
and \U$33737 ( \41801_42101 , \41568_41868 , \41574_41874 );
and \U$33738 ( \41802_42102 , \41568_41868 , \41581_41881 );
and \U$33739 ( \41803_42103 , \41574_41874 , \41581_41881 );
or \U$33740 ( \41804_42104 , \41801_42101 , \41802_42102 , \41803_42103 );
buf \U$33741 ( \41805_42105 , \41804_42104 );
and \U$33742 ( \41806_42106 , \41684_41984 , \41686_41986 );
and \U$33743 ( \41807_42107 , \41684_41984 , \41693_41993 );
and \U$33744 ( \41808_42108 , \41686_41986 , \41693_41993 );
or \U$33745 ( \41809_42109 , \41806_42106 , \41807_42107 , \41808_42108 );
buf \U$33746 ( \41810_42110 , \41809_42109 );
xor \U$33747 ( \41811_42111 , \41805_42105 , \41810_42110 );
and \U$33748 ( \41812_42112 , \41676_41976 , \41682_41982 );
buf \U$33749 ( \41813_42113 , \41812_42112 );
and \U$33750 ( \41814_42114 , \30670_29853 , \31877_32179_nG9bb4 );
and \U$33751 ( \41815_42115 , \29551_29850 , \32589_32888_nG9bb1 );
or \U$33752 ( \41816_42116 , \41814_42114 , \41815_42115 );
xor \U$33753 ( \41817_42117 , \29550_29849 , \41816_42116 );
buf \U$33754 ( \41818_42118 , \41817_42117 );
buf \U$33756 ( \41819_42119 , \41818_42118 );
xor \U$33757 ( \41820_42120 , \41813_42113 , \41819_42119 );
and \U$33758 ( \41821_42121 , \28946_28118 , \32881_33181_nG9bae );
and \U$33759 ( \41822_42122 , \27816_28115 , \33313_33613_nG9bab );
or \U$33760 ( \41823_42123 , \41821_42121 , \41822_42122 );
xor \U$33761 ( \41824_42124 , \27815_28114 , \41823_42123 );
buf \U$33762 ( \41825_42125 , \41824_42124 );
buf \U$33764 ( \41826_42126 , \41825_42125 );
xor \U$33765 ( \41827_42127 , \41820_42120 , \41826_42126 );
buf \U$33766 ( \41828_42128 , \41827_42127 );
xor \U$33767 ( \41829_42129 , \41811_42111 , \41828_42128 );
buf \U$33768 ( \41830_42130 , \41829_42129 );
and \U$33769 ( \41831_42131 , \21908_21658 , \35872_36172_nG9b96 );
and \U$33770 ( \41832_42132 , \21356_21655 , \36289_36589_nG9b93 );
or \U$33771 ( \41833_42133 , \41831_42131 , \41832_42132 );
xor \U$33772 ( \41834_42134 , \21355_21654 , \41833_42133 );
buf \U$33773 ( \41835_42135 , \41834_42134 );
buf \U$33775 ( \41836_42136 , \41835_42135 );
and \U$33776 ( \41837_42137 , \16405_15940 , \38668_38968_nG9b7e );
and \U$33777 ( \41838_42138 , \15638_15937 , \39034_39334_nG9b7b );
or \U$33778 ( \41839_42139 , \41837_42137 , \41838_42138 );
xor \U$33779 ( \41840_42140 , \15637_15936 , \41839_42139 );
buf \U$33780 ( \41841_42141 , \41840_42140 );
buf \U$33782 ( \41842_42142 , \41841_42141 );
xor \U$33783 ( \41843_42143 , \41836_42136 , \41842_42142 );
and \U$33784 ( \41844_42144 , \14710_14631 , \39291_39591_nG9b78 );
and \U$33785 ( \41845_42145 , \14329_14628 , \39663_39963_nG9b75 );
or \U$33786 ( \41846_42146 , \41844_42144 , \41845_42145 );
xor \U$33787 ( \41847_42147 , \14328_14627 , \41846_42146 );
buf \U$33788 ( \41848_42148 , \41847_42147 );
buf \U$33790 ( \41849_42149 , \41848_42148 );
xor \U$33791 ( \41850_42150 , \41843_42143 , \41849_42149 );
buf \U$33792 ( \41851_42151 , \41850_42150 );
xor \U$33793 ( \41852_42152 , \41830_42130 , \41851_42151 );
and \U$33794 ( \41853_42153 , \25044_24792 , \34343_34643_nG9ba2 );
and \U$33795 ( \41854_42154 , \24490_24789 , \34794_35094_nG9b9f );
or \U$33796 ( \41855_42155 , \41853_42153 , \41854_42154 );
xor \U$33797 ( \41856_42156 , \24489_24788 , \41855_42155 );
buf \U$33798 ( \41857_42157 , \41856_42156 );
buf \U$33800 ( \41858_42158 , \41857_42157 );
and \U$33801 ( \41859_42159 , \18908_18702 , \37307_37607_nG9b8a );
and \U$33802 ( \41860_42160 , \18400_18699 , \37674_37974_nG9b87 );
or \U$33803 ( \41861_42161 , \41859_42159 , \41860_42160 );
xor \U$33804 ( \41862_42162 , \18399_18698 , \41861_42161 );
buf \U$33805 ( \41863_42163 , \41862_42162 );
buf \U$33807 ( \41864_42164 , \41863_42163 );
xor \U$33808 ( \41865_42165 , \41858_42158 , \41864_42164 );
and \U$33809 ( \41866_42166 , \10411_10707 , \41663_41963_nG9b60 );
and \U$33810 ( \41867_42167 , \41635_41935 , \41639_41939 );
and \U$33811 ( \41868_42168 , \41639_41939 , \41651_41951 );
and \U$33812 ( \41869_42169 , \41635_41935 , \41651_41951 );
or \U$33813 ( \41870_42170 , \41867_42167 , \41868_42168 , \41869_42169 );
not \U$33814 ( \41871_42171 , \28774_29076 );
and \U$33815 ( \41872_42172 , \31752_32054 , \30521_30823 );
and \U$33816 ( \41873_42173 , \32495_32794 , \29944_30246 );
nor \U$33817 ( \41874_42174 , \41872_42172 , \41873_42173 );
xnor \U$33818 ( \41875_42175 , \41874_42174 , \30511_30813 );
xor \U$33819 ( \41876_42176 , \41871_42171 , \41875_42175 );
and \U$33820 ( \41877_42177 , \28782_29084 , \32503_32802 );
xor \U$33821 ( \41878_42178 , \41876_42176 , \41877_42177 );
xor \U$33822 ( \41879_42179 , \41870_42170 , \41878_42178 );
and \U$33823 ( \41880_42180 , \41644_41944 , \41648_41948 );
and \U$33824 ( \41881_42181 , \41648_41948 , \41650_41950 );
and \U$33825 ( \41882_42182 , \41644_41944 , \41650_41950 );
or \U$33826 ( \41883_42183 , \41880_42180 , \41881_42181 , \41882_42182 );
buf \U$33827 ( \41884_42184 , \41638_41938 );
xor \U$33828 ( \41885_42185 , \41883_42183 , \41884_42184 );
and \U$33829 ( \41886_42186 , \29966_30268 , \32555_32854 );
and \U$33830 ( \41887_42187 , \30500_30802 , \31765_32067 );
nor \U$33831 ( \41888_42188 , \41886_42186 , \41887_42187 );
xnor \U$33832 ( \41889_42189 , \41888_42188 , \32506_32805 );
xor \U$33833 ( \41890_42190 , \41885_42185 , \41889_42189 );
xor \U$33834 ( \41891_42191 , \41879_42179 , \41890_42190 );
and \U$33835 ( \41892_42192 , \41626_41926 , \41630_41930 );
and \U$33836 ( \41893_42193 , \41630_41930 , \41652_41952 );
and \U$33837 ( \41894_42194 , \41626_41926 , \41652_41952 );
or \U$33838 ( \41895_42195 , \41892_42192 , \41893_42193 , \41894_42194 );
xor \U$33839 ( \41896_42196 , \41891_42191 , \41895_42195 );
and \U$33840 ( \41897_42197 , \41653_41953 , \41657_41957 );
and \U$33841 ( \41898_42198 , \41658_41958 , \41661_41961 );
or \U$33842 ( \41899_42199 , \41897_42197 , \41898_42198 );
xor \U$33843 ( \41900_42200 , \41896_42196 , \41899_42199 );
buf g9b5d_GF_PartitionCandidate( \41901_42201_nG9b5d , \41900_42200 );
and \U$33844 ( \41902_42202 , \10402_10704 , \41901_42201_nG9b5d );
or \U$33845 ( \41903_42203 , \41866_42166 , \41902_42202 );
xor \U$33846 ( \41904_42204 , \10399_10703 , \41903_42203 );
buf \U$33847 ( \41905_42205 , \41904_42204 );
buf \U$33849 ( \41906_42206 , \41905_42205 );
xor \U$33850 ( \41907_42207 , \41865_42165 , \41906_42206 );
buf \U$33851 ( \41908_42208 , \41907_42207 );
xor \U$33852 ( \41909_42209 , \41852_42152 , \41908_42208 );
buf \U$33853 ( \41910_42210 , \41909_42209 );
xor \U$33854 ( \41911_42211 , \41800_42100 , \41910_42210 );
and \U$33855 ( \41912_42212 , \41556_41856 , \41561_41861 );
and \U$33856 ( \41913_42213 , \41556_41856 , \41583_41883 );
and \U$33857 ( \41914_42214 , \41561_41861 , \41583_41883 );
or \U$33858 ( \41915_42215 , \41912_42212 , \41913_42213 , \41914_42214 );
buf \U$33859 ( \41916_42216 , \41915_42215 );
and \U$33861 ( \41917_42217 , \32617_32916 , \28877_29179_nG9bbd );
or \U$33862 ( \41918_42218 , 1'b0 , \41917_42217 );
xor \U$33863 ( \41919_42219 , 1'b0 , \41918_42218 );
buf \U$33864 ( \41920_42220 , \41919_42219 );
buf \U$33866 ( \41921_42221 , \41920_42220 );
and \U$33867 ( \41922_42222 , \31989_31636 , \30064_30366_nG9bba );
and \U$33868 ( \41923_42223 , \31334_31633 , \30638_30940_nG9bb7 );
or \U$33869 ( \41924_42224 , \41922_42222 , \41923_42223 );
xor \U$33870 ( \41925_42225 , \31333_31632 , \41924_42224 );
buf \U$33871 ( \41926_42226 , \41925_42225 );
buf \U$33873 ( \41927_42227 , \41926_42226 );
xor \U$33874 ( \41928_42228 , \41921_42221 , \41927_42227 );
buf \U$33875 ( \41929_42229 , \41928_42228 );
and \U$33876 ( \41930_42230 , \27141_26431 , \33741_34041_nG9ba8 );
and \U$33877 ( \41931_42231 , \26129_26428 , \33994_34294_nG9ba5 );
or \U$33878 ( \41932_42232 , \41930_42230 , \41931_42231 );
xor \U$33879 ( \41933_42233 , \26128_26427 , \41932_42232 );
buf \U$33880 ( \41934_42234 , \41933_42233 );
buf \U$33882 ( \41935_42235 , \41934_42234 );
xor \U$33883 ( \41936_42236 , \41929_42229 , \41935_42235 );
and \U$33884 ( \41937_42237 , \23495_23201 , \35270_35570_nG9b9c );
and \U$33885 ( \41938_42238 , \22899_23198 , \35501_35801_nG9b99 );
or \U$33886 ( \41939_42239 , \41937_42237 , \41938_42238 );
xor \U$33887 ( \41940_42240 , \22898_23197 , \41939_42239 );
buf \U$33888 ( \41941_42241 , \41940_42240 );
buf \U$33890 ( \41942_42242 , \41941_42241 );
xor \U$33891 ( \41943_42243 , \41936_42236 , \41942_42242 );
buf \U$33892 ( \41944_42244 , \41943_42243 );
and \U$33893 ( \41945_42245 , \41614_41914 , \41620_41920 );
and \U$33894 ( \41946_42246 , \41614_41914 , \41668_41968 );
and \U$33895 ( \41947_42247 , \41620_41920 , \41668_41968 );
or \U$33896 ( \41948_42248 , \41945_42245 , \41946_42246 , \41947_42247 );
buf \U$33897 ( \41949_42249 , \41948_42248 );
xor \U$33898 ( \41950_42250 , \41944_42244 , \41949_42249 );
and \U$33899 ( \41951_42251 , \41461_41761 , \41467_41767 );
and \U$33900 ( \41952_42252 , \41461_41761 , \41474_41774 );
and \U$33901 ( \41953_42253 , \41467_41767 , \41474_41774 );
or \U$33902 ( \41954_42254 , \41951_42251 , \41952_42252 , \41953_42253 );
buf \U$33903 ( \41955_42255 , \41954_42254 );
xor \U$33904 ( \41956_42256 , \41950_42250 , \41955_42255 );
buf \U$33905 ( \41957_42257 , \41956_42256 );
xor \U$33906 ( \41958_42258 , \41916_42216 , \41957_42257 );
and \U$33907 ( \41959_42259 , \41521_41821 , \41526_41826 );
and \U$33908 ( \41960_42260 , \41521_41821 , \41548_41848 );
and \U$33909 ( \41961_42261 , \41526_41826 , \41548_41848 );
or \U$33910 ( \41962_42262 , \41959_42259 , \41960_42260 , \41961_42261 );
buf \U$33911 ( \41963_42263 , \41962_42262 );
xor \U$33912 ( \41964_42264 , \41958_42258 , \41963_42263 );
buf \U$33913 ( \41965_42265 , \41964_42264 );
xor \U$33914 ( \41966_42266 , \41911_42211 , \41965_42265 );
buf \U$33915 ( \41967_42267 , \41966_42266 );
xor \U$33916 ( \41968_42268 , \41795_42095 , \41967_42267 );
and \U$33917 ( \41969_42269 , \41714_42014 , \41968_42268 );
and \U$33919 ( \41970_42270 , \41708_42008 , \41713_42013 );
or \U$33921 ( \41971_42271 , 1'b0 , \41970_42270 , 1'b0 );
xor \U$33922 ( \41972_42272 , \41969_42269 , \41971_42271 );
and \U$33924 ( \41973_42273 , \41701_42001 , \41707_42007 );
and \U$33925 ( \41974_42274 , \41703_42003 , \41707_42007 );
or \U$33926 ( \41975_42275 , 1'b0 , \41973_42273 , \41974_42274 );
xor \U$33927 ( \41976_42276 , \41972_42272 , \41975_42275 );
xor \U$33934 ( \41977_42277 , \41976_42276 , 1'b0 );
and \U$33935 ( \41978_42278 , \41789_42089 , \41794_42094 );
and \U$33936 ( \41979_42279 , \41789_42089 , \41967_42267 );
and \U$33937 ( \41980_42280 , \41794_42094 , \41967_42267 );
or \U$33938 ( \41981_42281 , \41978_42278 , \41979_42279 , \41980_42280 );
xor \U$33939 ( \41982_42282 , \41977_42277 , \41981_42281 );
and \U$33940 ( \41983_42283 , \41800_42100 , \41910_42210 );
and \U$33941 ( \41984_42284 , \41800_42100 , \41965_42265 );
and \U$33942 ( \41985_42285 , \41910_42210 , \41965_42265 );
or \U$33943 ( \41986_42286 , \41983_42283 , \41984_42284 , \41985_42285 );
buf \U$33944 ( \41987_42287 , \41986_42286 );
and \U$33945 ( \41988_42288 , \41921_42221 , \41927_42227 );
buf \U$33946 ( \41989_42289 , \41988_42288 );
and \U$33947 ( \41990_42290 , \30670_29853 , \32589_32888_nG9bb1 );
and \U$33948 ( \41991_42291 , \29551_29850 , \32881_33181_nG9bae );
or \U$33949 ( \41992_42292 , \41990_42290 , \41991_42291 );
xor \U$33950 ( \41993_42293 , \29550_29849 , \41992_42292 );
buf \U$33951 ( \41994_42294 , \41993_42293 );
buf \U$33953 ( \41995_42295 , \41994_42294 );
xor \U$33954 ( \41996_42296 , \41989_42289 , \41995_42295 );
and \U$33955 ( \41997_42297 , \28946_28118 , \33313_33613_nG9bab );
and \U$33956 ( \41998_42298 , \27816_28115 , \33741_34041_nG9ba8 );
or \U$33957 ( \41999_42299 , \41997_42297 , \41998_42298 );
xor \U$33958 ( \42000_42300 , \27815_28114 , \41999_42299 );
buf \U$33959 ( \42001_42301 , \42000_42300 );
buf \U$33961 ( \42002_42302 , \42001_42301 );
xor \U$33962 ( \42003_42303 , \41996_42296 , \42002_42302 );
buf \U$33963 ( \42004_42304 , \42003_42303 );
and \U$33964 ( \42005_42305 , \41929_42229 , \41935_42235 );
and \U$33965 ( \42006_42306 , \41929_42229 , \41942_42242 );
and \U$33966 ( \42007_42307 , \41935_42235 , \41942_42242 );
or \U$33967 ( \42008_42308 , \42005_42305 , \42006_42306 , \42007_42307 );
buf \U$33968 ( \42009_42309 , \42008_42308 );
xor \U$33969 ( \42010_42310 , \42004_42304 , \42009_42309 );
and \U$33970 ( \42011_42311 , \41858_42158 , \41864_42164 );
and \U$33971 ( \42012_42312 , \41858_42158 , \41906_42206 );
and \U$33972 ( \42013_42313 , \41864_42164 , \41906_42206 );
or \U$33973 ( \42014_42314 , \42011_42311 , \42012_42312 , \42013_42313 );
buf \U$33974 ( \42015_42315 , \42014_42314 );
xor \U$33975 ( \42016_42316 , \42010_42310 , \42015_42315 );
buf \U$33976 ( \42017_42317 , \42016_42316 );
and \U$33977 ( \42018_42318 , \41813_42113 , \41819_42119 );
and \U$33978 ( \42019_42319 , \41813_42113 , \41826_42126 );
and \U$33979 ( \42020_42320 , \41819_42119 , \41826_42126 );
or \U$33980 ( \42021_42321 , \42018_42318 , \42019_42319 , \42020_42320 );
buf \U$33981 ( \42022_42322 , \42021_42321 );
and \U$33982 ( \42023_42323 , \17437_17297 , \38363_38663_nG9b81 );
and \U$33983 ( \42024_42324 , \16995_17294 , \38668_38968_nG9b7e );
or \U$33984 ( \42025_42325 , \42023_42323 , \42024_42324 );
xor \U$33985 ( \42026_42326 , \16994_17293 , \42025_42325 );
buf \U$33986 ( \42027_42327 , \42026_42326 );
buf \U$33988 ( \42028_42328 , \42027_42327 );
xor \U$33989 ( \42029_42329 , \42022_42322 , \42028_42328 );
and \U$33990 ( \42030_42330 , \12183_12157 , \40740_41040_nG9b69 );
and \U$33991 ( \42031_42331 , \11855_12154 , \41081_41381_nG9b66 );
or \U$33992 ( \42032_42332 , \42030_42330 , \42031_42331 );
xor \U$33993 ( \42033_42333 , \11854_12153 , \42032_42332 );
buf \U$33994 ( \42034_42334 , \42033_42333 );
buf \U$33996 ( \42035_42335 , \42034_42334 );
xor \U$33997 ( \42036_42336 , \42029_42329 , \42035_42335 );
buf \U$33998 ( \42037_42337 , \42036_42336 );
xor \U$33999 ( \42038_42338 , \42017_42317 , \42037_42337 );
and \U$34000 ( \42039_42339 , \21908_21658 , \36289_36589_nG9b93 );
and \U$34001 ( \42040_42340 , \21356_21655 , \36686_36986_nG9b90 );
or \U$34002 ( \42041_42341 , \42039_42339 , \42040_42340 );
xor \U$34003 ( \42042_42342 , \21355_21654 , \42041_42341 );
buf \U$34004 ( \42043_42343 , \42042_42342 );
buf \U$34006 ( \42044_42344 , \42043_42343 );
and \U$34007 ( \42045_42345 , \16405_15940 , \39034_39334_nG9b7b );
and \U$34008 ( \42046_42346 , \15638_15937 , \39291_39591_nG9b78 );
or \U$34009 ( \42047_42347 , \42045_42345 , \42046_42346 );
xor \U$34010 ( \42048_42348 , \15637_15936 , \42047_42347 );
buf \U$34011 ( \42049_42349 , \42048_42348 );
buf \U$34013 ( \42050_42350 , \42049_42349 );
xor \U$34014 ( \42051_42351 , \42044_42344 , \42050_42350 );
and \U$34015 ( \42052_42352 , \14710_14631 , \39663_39963_nG9b75 );
and \U$34016 ( \42053_42353 , \14329_14628 , \39904_40204_nG9b72 );
or \U$34017 ( \42054_42354 , \42052_42352 , \42053_42353 );
xor \U$34018 ( \42055_42355 , \14328_14627 , \42054_42354 );
buf \U$34019 ( \42056_42356 , \42055_42355 );
buf \U$34021 ( \42057_42357 , \42056_42356 );
xor \U$34022 ( \42058_42358 , \42051_42351 , \42057_42357 );
buf \U$34023 ( \42059_42359 , \42058_42358 );
xor \U$34024 ( \42060_42360 , \42038_42338 , \42059_42359 );
buf \U$34025 ( \42061_42361 , \42060_42360 );
and \U$34026 ( \42062_42362 , \41724_42024 , \41730_42030 );
and \U$34027 ( \42063_42363 , \41724_42024 , \41737_42037 );
and \U$34028 ( \42064_42364 , \41730_42030 , \41737_42037 );
or \U$34029 ( \42065_42365 , \42062_42362 , \42063_42363 , \42064_42364 );
buf \U$34030 ( \42066_42366 , \42065_42365 );
and \U$34031 ( \42067_42367 , \20353_20155 , \36950_37250_nG9b8d );
and \U$34032 ( \42068_42368 , \19853_20152 , \37307_37607_nG9b8a );
or \U$34033 ( \42069_42369 , \42067_42367 , \42068_42368 );
xor \U$34034 ( \42070_42370 , \19852_20151 , \42069_42369 );
buf \U$34035 ( \42071_42371 , \42070_42370 );
buf \U$34037 ( \42072_42372 , \42071_42371 );
and \U$34038 ( \42073_42373 , \13431_13370 , \40152_40452_nG9b6f );
and \U$34039 ( \42074_42374 , \13068_13367 , \40543_40843_nG9b6c );
or \U$34040 ( \42075_42375 , \42073_42373 , \42074_42374 );
xor \U$34041 ( \42076_42376 , \13067_13366 , \42075_42375 );
buf \U$34042 ( \42077_42377 , \42076_42376 );
buf \U$34044 ( \42078_42378 , \42077_42377 );
xor \U$34045 ( \42079_42379 , \42072_42372 , \42078_42378 );
and \U$34046 ( \42080_42380 , \10996_10421 , \41385_41685_nG9b63 );
and \U$34047 ( \42081_42381 , \10119_10418 , \41663_41963_nG9b60 );
or \U$34048 ( \42082_42382 , \42080_42380 , \42081_42381 );
xor \U$34049 ( \42083_42383 , \10118_10417 , \42082_42382 );
buf \U$34050 ( \42084_42384 , \42083_42383 );
buf \U$34052 ( \42085_42385 , \42084_42384 );
xor \U$34053 ( \42086_42386 , \42079_42379 , \42085_42385 );
buf \U$34054 ( \42087_42387 , \42086_42386 );
xor \U$34055 ( \42088_42388 , \42066_42366 , \42087_42387 );
and \U$34056 ( \42089_42389 , \25044_24792 , \34794_35094_nG9b9f );
and \U$34057 ( \42090_42390 , \24490_24789 , \35270_35570_nG9b9c );
or \U$34058 ( \42091_42391 , \42089_42389 , \42090_42390 );
xor \U$34059 ( \42092_42392 , \24489_24788 , \42091_42391 );
buf \U$34060 ( \42093_42393 , \42092_42392 );
buf \U$34062 ( \42094_42394 , \42093_42393 );
and \U$34063 ( \42095_42395 , \18908_18702 , \37674_37974_nG9b87 );
and \U$34064 ( \42096_42396 , \18400_18699 , \38037_38337_nG9b84 );
or \U$34065 ( \42097_42397 , \42095_42395 , \42096_42396 );
xor \U$34066 ( \42098_42398 , \18399_18698 , \42097_42397 );
buf \U$34067 ( \42099_42399 , \42098_42398 );
buf \U$34069 ( \42100_42400 , \42099_42399 );
xor \U$34070 ( \42101_42401 , \42094_42394 , \42100_42400 );
and \U$34071 ( \42102_42402 , \10411_10707 , \41901_42201_nG9b5d );
and \U$34072 ( \42103_42403 , \41871_42171 , \41875_42175 );
and \U$34073 ( \42104_42404 , \41875_42175 , \41877_42177 );
and \U$34074 ( \42105_42405 , \41871_42171 , \41877_42177 );
or \U$34075 ( \42106_42406 , \42103_42403 , \42104_42404 , \42105_42405 );
and \U$34076 ( \42107_42407 , \41883_42183 , \41884_42184 );
and \U$34077 ( \42108_42408 , \41884_42184 , \41889_42189 );
and \U$34078 ( \42109_42409 , \41883_42183 , \41889_42189 );
or \U$34079 ( \42110_42410 , \42107_42407 , \42108_42408 , \42109_42409 );
xor \U$34080 ( \42111_42411 , \42106_42406 , \42110_42410 );
and \U$34081 ( \42112_42412 , \32495_32794 , \30521_30823 );
not \U$34082 ( \42113_42413 , \42112_42412 );
xnor \U$34083 ( \42114_42414 , \42113_42413 , \30511_30813 );
not \U$34084 ( \42115_42415 , \42114_42414 );
and \U$34085 ( \42116_42416 , \30500_30802 , \32555_32854 );
and \U$34086 ( \42117_42417 , \31752_32054 , \31765_32067 );
nor \U$34087 ( \42118_42418 , \42116_42416 , \42117_42417 );
xnor \U$34088 ( \42119_42419 , \42118_42418 , \32506_32805 );
xor \U$34089 ( \42120_42420 , \42115_42415 , \42119_42419 );
and \U$34090 ( \42121_42421 , \29966_30268 , \32503_32802 );
xor \U$34091 ( \42122_42422 , \42120_42420 , \42121_42421 );
xor \U$34092 ( \42123_42423 , \42111_42411 , \42122_42422 );
and \U$34093 ( \42124_42424 , \41870_42170 , \41878_42178 );
and \U$34094 ( \42125_42425 , \41878_42178 , \41890_42190 );
and \U$34095 ( \42126_42426 , \41870_42170 , \41890_42190 );
or \U$34096 ( \42127_42427 , \42124_42424 , \42125_42425 , \42126_42426 );
xor \U$34097 ( \42128_42428 , \42123_42423 , \42127_42427 );
and \U$34098 ( \42129_42429 , \41891_42191 , \41895_42195 );
and \U$34099 ( \42130_42430 , \41896_42196 , \41899_42199 );
or \U$34100 ( \42131_42431 , \42129_42429 , \42130_42430 );
xor \U$34101 ( \42132_42432 , \42128_42428 , \42131_42431 );
buf g9b5a_GF_PartitionCandidate( \42133_42433_nG9b5a , \42132_42432 );
and \U$34102 ( \42134_42434 , \10402_10704 , \42133_42433_nG9b5a );
or \U$34103 ( \42135_42435 , \42102_42402 , \42134_42434 );
xor \U$34104 ( \42136_42436 , \10399_10703 , \42135_42435 );
buf \U$34105 ( \42137_42437 , \42136_42436 );
buf \U$34107 ( \42138_42438 , \42137_42437 );
xor \U$34108 ( \42139_42439 , \42101_42401 , \42138_42438 );
buf \U$34109 ( \42140_42440 , \42139_42439 );
xor \U$34110 ( \42141_42441 , \42088_42388 , \42140_42440 );
buf \U$34111 ( \42142_42442 , \42141_42441 );
xor \U$34112 ( \42143_42443 , \42061_42361 , \42142_42442 );
and \U$34113 ( \42144_42444 , \41739_42039 , \41744_42044 );
and \U$34114 ( \42145_42445 , \41739_42039 , \41766_42066 );
and \U$34115 ( \42146_42446 , \41744_42044 , \41766_42066 );
or \U$34116 ( \42147_42447 , \42144_42444 , \42145_42445 , \42146_42446 );
buf \U$34117 ( \42148_42448 , \42147_42447 );
xor \U$34118 ( \42149_42449 , \42143_42443 , \42148_42448 );
buf \U$34119 ( \42150_42450 , \42149_42449 );
xor \U$34120 ( \42151_42451 , \41987_42287 , \42150_42450 );
and \U$34121 ( \42152_42452 , \41768_42068 , \41773_42073 );
and \U$34122 ( \42153_42453 , \41768_42068 , \41779_42079 );
and \U$34123 ( \42154_42454 , \41773_42073 , \41779_42079 );
or \U$34124 ( \42155_42455 , \42152_42452 , \42153_42453 , \42154_42454 );
buf \U$34125 ( \42156_42456 , \42155_42455 );
xor \U$34126 ( \42157_42457 , \42151_42451 , \42156_42456 );
buf \U$34127 ( \42158_42458 , \42157_42457 );
and \U$34128 ( \42159_42459 , \41719_42019 , \41781_42081 );
and \U$34129 ( \42160_42460 , \41719_42019 , \41787_42087 );
and \U$34130 ( \42161_42461 , \41781_42081 , \41787_42087 );
or \U$34131 ( \42162_42462 , \42159_42459 , \42160_42460 , \42161_42461 );
buf \U$34132 ( \42163_42463 , \42162_42462 );
xor \U$34133 ( \42164_42464 , \42158_42458 , \42163_42463 );
and \U$34134 ( \42165_42465 , \41916_42216 , \41957_42257 );
and \U$34135 ( \42166_42466 , \41916_42216 , \41963_42263 );
and \U$34136 ( \42167_42467 , \41957_42257 , \41963_42263 );
or \U$34137 ( \42168_42468 , \42165_42465 , \42166_42466 , \42167_42467 );
buf \U$34138 ( \42169_42469 , \42168_42468 );
and \U$34140 ( \42170_42470 , \32617_32916 , \30064_30366_nG9bba );
or \U$34141 ( \42171_42471 , 1'b0 , \42170_42470 );
xor \U$34142 ( \42172_42472 , 1'b0 , \42171_42471 );
buf \U$34143 ( \42173_42473 , \42172_42472 );
buf \U$34145 ( \42174_42474 , \42173_42473 );
and \U$34146 ( \42175_42475 , \31989_31636 , \30638_30940_nG9bb7 );
and \U$34147 ( \42176_42476 , \31334_31633 , \31877_32179_nG9bb4 );
or \U$34148 ( \42177_42477 , \42175_42475 , \42176_42476 );
xor \U$34149 ( \42178_42478 , \31333_31632 , \42177_42477 );
buf \U$34150 ( \42179_42479 , \42178_42478 );
buf \U$34152 ( \42180_42480 , \42179_42479 );
xor \U$34153 ( \42181_42481 , \42174_42474 , \42180_42480 );
buf \U$34154 ( \42182_42482 , \42181_42481 );
and \U$34155 ( \42183_42483 , \27141_26431 , \33994_34294_nG9ba5 );
and \U$34156 ( \42184_42484 , \26129_26428 , \34343_34643_nG9ba2 );
or \U$34157 ( \42185_42485 , \42183_42483 , \42184_42484 );
xor \U$34158 ( \42186_42486 , \26128_26427 , \42185_42485 );
buf \U$34159 ( \42187_42487 , \42186_42486 );
buf \U$34161 ( \42188_42488 , \42187_42487 );
xor \U$34162 ( \42189_42489 , \42182_42482 , \42188_42488 );
and \U$34163 ( \42190_42490 , \23495_23201 , \35501_35801_nG9b99 );
and \U$34164 ( \42191_42491 , \22899_23198 , \35872_36172_nG9b96 );
or \U$34165 ( \42192_42492 , \42190_42490 , \42191_42491 );
xor \U$34166 ( \42193_42493 , \22898_23197 , \42192_42492 );
buf \U$34167 ( \42194_42494 , \42193_42493 );
buf \U$34169 ( \42195_42495 , \42194_42494 );
xor \U$34170 ( \42196_42496 , \42189_42489 , \42195_42495 );
buf \U$34171 ( \42197_42497 , \42196_42496 );
and \U$34172 ( \42198_42498 , \41751_42051 , \41757_42057 );
and \U$34173 ( \42199_42499 , \41751_42051 , \41764_42064 );
and \U$34174 ( \42200_42500 , \41757_42057 , \41764_42064 );
or \U$34175 ( \42201_42501 , \42198_42498 , \42199_42499 , \42200_42500 );
buf \U$34176 ( \42202_42502 , \42201_42501 );
xor \U$34177 ( \42203_42503 , \42197_42497 , \42202_42502 );
and \U$34178 ( \42204_42504 , \41836_42136 , \41842_42142 );
and \U$34179 ( \42205_42505 , \41836_42136 , \41849_42149 );
and \U$34180 ( \42206_42506 , \41842_42142 , \41849_42149 );
or \U$34181 ( \42207_42507 , \42204_42504 , \42205_42505 , \42206_42506 );
buf \U$34182 ( \42208_42508 , \42207_42507 );
xor \U$34183 ( \42209_42509 , \42203_42503 , \42208_42508 );
buf \U$34184 ( \42210_42510 , \42209_42509 );
and \U$34185 ( \42211_42511 , \41944_42244 , \41949_42249 );
and \U$34186 ( \42212_42512 , \41944_42244 , \41955_42255 );
and \U$34187 ( \42213_42513 , \41949_42249 , \41955_42255 );
or \U$34188 ( \42214_42514 , \42211_42511 , \42212_42512 , \42213_42513 );
buf \U$34189 ( \42215_42515 , \42214_42514 );
xor \U$34190 ( \42216_42516 , \42210_42510 , \42215_42515 );
and \U$34191 ( \42217_42517 , \41805_42105 , \41810_42110 );
and \U$34192 ( \42218_42518 , \41805_42105 , \41828_42128 );
and \U$34193 ( \42219_42519 , \41810_42110 , \41828_42128 );
or \U$34194 ( \42220_42520 , \42217_42517 , \42218_42518 , \42219_42519 );
buf \U$34195 ( \42221_42521 , \42220_42520 );
xor \U$34196 ( \42222_42522 , \42216_42516 , \42221_42521 );
buf \U$34197 ( \42223_42523 , \42222_42522 );
xor \U$34198 ( \42224_42524 , \42169_42469 , \42223_42523 );
and \U$34199 ( \42225_42525 , \41830_42130 , \41851_42151 );
and \U$34200 ( \42226_42526 , \41830_42130 , \41908_42208 );
and \U$34201 ( \42227_42527 , \41851_42151 , \41908_42208 );
or \U$34202 ( \42228_42528 , \42225_42525 , \42226_42526 , \42227_42527 );
buf \U$34203 ( \42229_42529 , \42228_42528 );
xor \U$34204 ( \42230_42530 , \42224_42524 , \42229_42529 );
buf \U$34205 ( \42231_42531 , \42230_42530 );
xor \U$34206 ( \42232_42532 , \42164_42464 , \42231_42531 );
and \U$34207 ( \42233_42533 , \41982_42282 , \42232_42532 );
and \U$34209 ( \42234_42534 , \41976_42276 , \41981_42281 );
or \U$34211 ( \42235_42535 , 1'b0 , \42234_42534 , 1'b0 );
xor \U$34212 ( \42236_42536 , \42233_42533 , \42235_42535 );
and \U$34214 ( \42237_42537 , \41969_42269 , \41975_42275 );
and \U$34215 ( \42238_42538 , \41971_42271 , \41975_42275 );
or \U$34216 ( \42239_42539 , 1'b0 , \42237_42537 , \42238_42538 );
xor \U$34217 ( \42240_42540 , \42236_42536 , \42239_42539 );
xor \U$34224 ( \42241_42541 , \42240_42540 , 1'b0 );
and \U$34225 ( \42242_42542 , \42158_42458 , \42163_42463 );
and \U$34226 ( \42243_42543 , \42158_42458 , \42231_42531 );
and \U$34227 ( \42244_42544 , \42163_42463 , \42231_42531 );
or \U$34228 ( \42245_42545 , \42242_42542 , \42243_42543 , \42244_42544 );
xor \U$34229 ( \42246_42546 , \42241_42541 , \42245_42545 );
and \U$34230 ( \42247_42547 , \42169_42469 , \42223_42523 );
and \U$34231 ( \42248_42548 , \42169_42469 , \42229_42529 );
and \U$34232 ( \42249_42549 , \42223_42523 , \42229_42529 );
or \U$34233 ( \42250_42550 , \42247_42547 , \42248_42548 , \42249_42549 );
buf \U$34234 ( \42251_42551 , \42250_42550 );
and \U$34235 ( \42252_42552 , \42061_42361 , \42142_42442 );
and \U$34236 ( \42253_42553 , \42061_42361 , \42148_42448 );
and \U$34237 ( \42254_42554 , \42142_42442 , \42148_42448 );
or \U$34238 ( \42255_42555 , \42252_42552 , \42253_42553 , \42254_42554 );
buf \U$34239 ( \42256_42556 , \42255_42555 );
xor \U$34240 ( \42257_42557 , \42251_42551 , \42256_42556 );
and \U$34241 ( \42258_42558 , \42017_42317 , \42037_42337 );
and \U$34242 ( \42259_42559 , \42017_42317 , \42059_42359 );
and \U$34243 ( \42260_42560 , \42037_42337 , \42059_42359 );
or \U$34244 ( \42261_42561 , \42258_42558 , \42259_42559 , \42260_42560 );
buf \U$34245 ( \42262_42562 , \42261_42561 );
and \U$34247 ( \42263_42563 , \32617_32916 , \30638_30940_nG9bb7 );
or \U$34248 ( \42264_42564 , 1'b0 , \42263_42563 );
xor \U$34249 ( \42265_42565 , 1'b0 , \42264_42564 );
buf \U$34250 ( \42266_42566 , \42265_42565 );
buf \U$34252 ( \42267_42567 , \42266_42566 );
and \U$34253 ( \42268_42568 , \30670_29853 , \32881_33181_nG9bae );
and \U$34254 ( \42269_42569 , \29551_29850 , \33313_33613_nG9bab );
or \U$34255 ( \42270_42570 , \42268_42568 , \42269_42569 );
xor \U$34256 ( \42271_42571 , \29550_29849 , \42270_42570 );
buf \U$34257 ( \42272_42572 , \42271_42571 );
buf \U$34259 ( \42273_42573 , \42272_42572 );
xor \U$34260 ( \42274_42574 , \42267_42567 , \42273_42573 );
buf \U$34261 ( \42275_42575 , \42274_42574 );
and \U$34262 ( \42276_42576 , \20353_20155 , \37307_37607_nG9b8a );
and \U$34263 ( \42277_42577 , \19853_20152 , \37674_37974_nG9b87 );
or \U$34264 ( \42278_42578 , \42276_42576 , \42277_42577 );
xor \U$34265 ( \42279_42579 , \19852_20151 , \42278_42578 );
buf \U$34266 ( \42280_42580 , \42279_42579 );
buf \U$34268 ( \42281_42581 , \42280_42580 );
xor \U$34269 ( \42282_42582 , \42275_42575 , \42281_42581 );
and \U$34270 ( \42283_42583 , \18908_18702 , \38037_38337_nG9b84 );
and \U$34271 ( \42284_42584 , \18400_18699 , \38363_38663_nG9b81 );
or \U$34272 ( \42285_42585 , \42283_42583 , \42284_42584 );
xor \U$34273 ( \42286_42586 , \18399_18698 , \42285_42585 );
buf \U$34274 ( \42287_42587 , \42286_42586 );
buf \U$34276 ( \42288_42588 , \42287_42587 );
xor \U$34277 ( \42289_42589 , \42282_42582 , \42288_42588 );
buf \U$34278 ( \42290_42590 , \42289_42589 );
and \U$34279 ( \42291_42591 , \23495_23201 , \35872_36172_nG9b96 );
and \U$34280 ( \42292_42592 , \22899_23198 , \36289_36589_nG9b93 );
or \U$34281 ( \42293_42593 , \42291_42591 , \42292_42592 );
xor \U$34282 ( \42294_42594 , \22898_23197 , \42293_42593 );
buf \U$34283 ( \42295_42595 , \42294_42594 );
buf \U$34285 ( \42296_42596 , \42295_42595 );
and \U$34286 ( \42297_42597 , \21908_21658 , \36686_36986_nG9b90 );
and \U$34287 ( \42298_42598 , \21356_21655 , \36950_37250_nG9b8d );
or \U$34288 ( \42299_42599 , \42297_42597 , \42298_42598 );
xor \U$34289 ( \42300_42600 , \21355_21654 , \42299_42599 );
buf \U$34290 ( \42301_42601 , \42300_42600 );
buf \U$34292 ( \42302_42602 , \42301_42601 );
xor \U$34293 ( \42303_42603 , \42296_42596 , \42302_42602 );
and \U$34294 ( \42304_42604 , \14710_14631 , \39904_40204_nG9b72 );
and \U$34295 ( \42305_42605 , \14329_14628 , \40152_40452_nG9b6f );
or \U$34296 ( \42306_42606 , \42304_42604 , \42305_42605 );
xor \U$34297 ( \42307_42607 , \14328_14627 , \42306_42606 );
buf \U$34298 ( \42308_42608 , \42307_42607 );
buf \U$34300 ( \42309_42609 , \42308_42608 );
xor \U$34301 ( \42310_42610 , \42303_42603 , \42309_42609 );
buf \U$34302 ( \42311_42611 , \42310_42610 );
xor \U$34303 ( \42312_42612 , \42290_42590 , \42311_42611 );
and \U$34304 ( \42313_42613 , \16405_15940 , \39291_39591_nG9b78 );
and \U$34305 ( \42314_42614 , \15638_15937 , \39663_39963_nG9b75 );
or \U$34306 ( \42315_42615 , \42313_42613 , \42314_42614 );
xor \U$34307 ( \42316_42616 , \15637_15936 , \42315_42615 );
buf \U$34308 ( \42317_42617 , \42316_42616 );
buf \U$34310 ( \42318_42618 , \42317_42617 );
and \U$34311 ( \42319_42619 , \12183_12157 , \41081_41381_nG9b66 );
and \U$34312 ( \42320_42620 , \11855_12154 , \41385_41685_nG9b63 );
or \U$34313 ( \42321_42621 , \42319_42619 , \42320_42620 );
xor \U$34314 ( \42322_42622 , \11854_12153 , \42321_42621 );
buf \U$34315 ( \42323_42623 , \42322_42622 );
buf \U$34317 ( \42324_42624 , \42323_42623 );
xor \U$34318 ( \42325_42625 , \42318_42618 , \42324_42624 );
and \U$34319 ( \42326_42626 , \10996_10421 , \41663_41963_nG9b60 );
and \U$34320 ( \42327_42627 , \10119_10418 , \41901_42201_nG9b5d );
or \U$34321 ( \42328_42628 , \42326_42626 , \42327_42627 );
xor \U$34322 ( \42329_42629 , \10118_10417 , \42328_42628 );
buf \U$34323 ( \42330_42630 , \42329_42629 );
buf \U$34325 ( \42331_42631 , \42330_42630 );
xor \U$34326 ( \42332_42632 , \42325_42625 , \42331_42631 );
buf \U$34327 ( \42333_42633 , \42332_42632 );
xor \U$34328 ( \42334_42634 , \42312_42612 , \42333_42633 );
buf \U$34329 ( \42335_42635 , \42334_42634 );
xor \U$34330 ( \42336_42636 , \42262_42562 , \42335_42635 );
and \U$34331 ( \42337_42637 , \42066_42366 , \42087_42387 );
and \U$34332 ( \42338_42638 , \42066_42366 , \42140_42440 );
and \U$34333 ( \42339_42639 , \42087_42387 , \42140_42440 );
or \U$34334 ( \42340_42640 , \42337_42637 , \42338_42638 , \42339_42639 );
buf \U$34335 ( \42341_42641 , \42340_42640 );
xor \U$34336 ( \42342_42642 , \42336_42636 , \42341_42641 );
buf \U$34337 ( \42343_42643 , \42342_42642 );
xor \U$34338 ( \42344_42644 , \42257_42557 , \42343_42643 );
buf \U$34339 ( \42345_42645 , \42344_42644 );
and \U$34340 ( \42346_42646 , \41987_42287 , \42150_42450 );
and \U$34341 ( \42347_42647 , \41987_42287 , \42156_42456 );
and \U$34342 ( \42348_42648 , \42150_42450 , \42156_42456 );
or \U$34343 ( \42349_42649 , \42346_42646 , \42347_42647 , \42348_42648 );
buf \U$34344 ( \42350_42650 , \42349_42649 );
xor \U$34345 ( \42351_42651 , \42345_42645 , \42350_42650 );
and \U$34346 ( \42352_42652 , \42044_42344 , \42050_42350 );
and \U$34347 ( \42353_42653 , \42044_42344 , \42057_42357 );
and \U$34348 ( \42354_42654 , \42050_42350 , \42057_42357 );
or \U$34349 ( \42355_42655 , \42352_42652 , \42353_42653 , \42354_42654 );
buf \U$34350 ( \42356_42656 , \42355_42655 );
and \U$34351 ( \42357_42657 , \28946_28118 , \33741_34041_nG9ba8 );
and \U$34352 ( \42358_42658 , \27816_28115 , \33994_34294_nG9ba5 );
or \U$34353 ( \42359_42659 , \42357_42657 , \42358_42658 );
xor \U$34354 ( \42360_42660 , \27815_28114 , \42359_42659 );
buf \U$34355 ( \42361_42661 , \42360_42660 );
buf \U$34357 ( \42362_42662 , \42361_42661 );
and \U$34358 ( \42363_42663 , \27141_26431 , \34343_34643_nG9ba2 );
and \U$34359 ( \42364_42664 , \26129_26428 , \34794_35094_nG9b9f );
or \U$34360 ( \42365_42665 , \42363_42663 , \42364_42664 );
xor \U$34361 ( \42366_42666 , \26128_26427 , \42365_42665 );
buf \U$34362 ( \42367_42667 , \42366_42666 );
buf \U$34364 ( \42368_42668 , \42367_42667 );
xor \U$34365 ( \42369_42669 , \42362_42662 , \42368_42668 );
and \U$34366 ( \42370_42670 , \13431_13370 , \40543_40843_nG9b6c );
and \U$34367 ( \42371_42671 , \13068_13367 , \40740_41040_nG9b69 );
or \U$34368 ( \42372_42672 , \42370_42670 , \42371_42671 );
xor \U$34369 ( \42373_42673 , \13067_13366 , \42372_42672 );
buf \U$34370 ( \42374_42674 , \42373_42673 );
buf \U$34372 ( \42375_42675 , \42374_42674 );
xor \U$34373 ( \42376_42676 , \42369_42669 , \42375_42675 );
buf \U$34374 ( \42377_42677 , \42376_42676 );
xor \U$34375 ( \42378_42678 , \42356_42656 , \42377_42677 );
and \U$34376 ( \42379_42679 , \42174_42474 , \42180_42480 );
buf \U$34377 ( \42380_42680 , \42379_42679 );
and \U$34378 ( \42381_42681 , \31989_31636 , \31877_32179_nG9bb4 );
and \U$34379 ( \42382_42682 , \31334_31633 , \32589_32888_nG9bb1 );
or \U$34380 ( \42383_42683 , \42381_42681 , \42382_42682 );
xor \U$34381 ( \42384_42684 , \31333_31632 , \42383_42683 );
buf \U$34382 ( \42385_42685 , \42384_42684 );
buf \U$34384 ( \42386_42686 , \42385_42685 );
xor \U$34385 ( \42387_42687 , \42380_42680 , \42386_42686 );
and \U$34386 ( \42388_42688 , \25044_24792 , \35270_35570_nG9b9c );
and \U$34387 ( \42389_42689 , \24490_24789 , \35501_35801_nG9b99 );
or \U$34388 ( \42390_42690 , \42388_42688 , \42389_42689 );
xor \U$34389 ( \42391_42691 , \24489_24788 , \42390_42690 );
buf \U$34390 ( \42392_42692 , \42391_42691 );
buf \U$34392 ( \42393_42693 , \42392_42692 );
xor \U$34393 ( \42394_42694 , \42387_42687 , \42393_42693 );
buf \U$34394 ( \42395_42695 , \42394_42694 );
xor \U$34395 ( \42396_42696 , \42378_42678 , \42395_42695 );
buf \U$34396 ( \42397_42697 , \42396_42696 );
and \U$34397 ( \42398_42698 , \42094_42394 , \42100_42400 );
and \U$34398 ( \42399_42699 , \42094_42394 , \42138_42438 );
and \U$34399 ( \42400_42700 , \42100_42400 , \42138_42438 );
or \U$34400 ( \42401_42701 , \42398_42698 , \42399_42699 , \42400_42700 );
buf \U$34401 ( \42402_42702 , \42401_42701 );
and \U$34402 ( \42403_42703 , \42072_42372 , \42078_42378 );
and \U$34403 ( \42404_42704 , \42072_42372 , \42085_42385 );
and \U$34404 ( \42405_42705 , \42078_42378 , \42085_42385 );
or \U$34405 ( \42406_42706 , \42403_42703 , \42404_42704 , \42405_42705 );
buf \U$34406 ( \42407_42707 , \42406_42706 );
xor \U$34407 ( \42408_42708 , \42402_42702 , \42407_42707 );
and \U$34408 ( \42409_42709 , \42182_42482 , \42188_42488 );
and \U$34409 ( \42410_42710 , \42182_42482 , \42195_42495 );
and \U$34410 ( \42411_42711 , \42188_42488 , \42195_42495 );
or \U$34411 ( \42412_42712 , \42409_42709 , \42410_42710 , \42411_42711 );
buf \U$34412 ( \42413_42713 , \42412_42712 );
xor \U$34413 ( \42414_42714 , \42408_42708 , \42413_42713 );
buf \U$34414 ( \42415_42715 , \42414_42714 );
xor \U$34415 ( \42416_42716 , \42397_42697 , \42415_42715 );
and \U$34416 ( \42417_42717 , \42197_42497 , \42202_42502 );
and \U$34417 ( \42418_42718 , \42197_42497 , \42208_42508 );
and \U$34418 ( \42419_42719 , \42202_42502 , \42208_42508 );
or \U$34419 ( \42420_42720 , \42417_42717 , \42418_42718 , \42419_42719 );
buf \U$34420 ( \42421_42721 , \42420_42720 );
xor \U$34421 ( \42422_42722 , \42416_42716 , \42421_42721 );
buf \U$34422 ( \42423_42723 , \42422_42722 );
and \U$34423 ( \42424_42724 , \42004_42304 , \42009_42309 );
and \U$34424 ( \42425_42725 , \42004_42304 , \42015_42315 );
and \U$34425 ( \42426_42726 , \42009_42309 , \42015_42315 );
or \U$34426 ( \42427_42727 , \42424_42724 , \42425_42725 , \42426_42726 );
buf \U$34427 ( \42428_42728 , \42427_42727 );
and \U$34428 ( \42429_42729 , \41989_42289 , \41995_42295 );
and \U$34429 ( \42430_42730 , \41989_42289 , \42002_42302 );
and \U$34430 ( \42431_42731 , \41995_42295 , \42002_42302 );
or \U$34431 ( \42432_42732 , \42429_42729 , \42430_42730 , \42431_42731 );
buf \U$34432 ( \42433_42733 , \42432_42732 );
and \U$34433 ( \42434_42734 , \17437_17297 , \38668_38968_nG9b7e );
and \U$34434 ( \42435_42735 , \16995_17294 , \39034_39334_nG9b7b );
or \U$34435 ( \42436_42736 , \42434_42734 , \42435_42735 );
xor \U$34436 ( \42437_42737 , \16994_17293 , \42436_42736 );
buf \U$34437 ( \42438_42738 , \42437_42737 );
buf \U$34439 ( \42439_42739 , \42438_42738 );
xor \U$34440 ( \42440_42740 , \42433_42733 , \42439_42739 );
and \U$34441 ( \42441_42741 , \10411_10707 , \42133_42433_nG9b5a );
and \U$34442 ( \42442_42742 , \42115_42415 , \42119_42419 );
and \U$34443 ( \42443_42743 , \42119_42419 , \42121_42421 );
and \U$34444 ( \42444_42744 , \42115_42415 , \42121_42421 );
or \U$34445 ( \42445_42745 , \42442_42742 , \42443_42743 , \42444_42744 );
buf \U$34446 ( \42446_42746 , \42114_42414 );
xor \U$34447 ( \42447_42747 , \42445_42745 , \42446_42746 );
not \U$34448 ( \42448_42748 , \30511_30813 );
and \U$34449 ( \42449_42749 , \31752_32054 , \32555_32854 );
and \U$34450 ( \42450_42750 , \32495_32794 , \31765_32067 );
nor \U$34451 ( \42451_42751 , \42449_42749 , \42450_42750 );
xnor \U$34452 ( \42452_42752 , \42451_42751 , \32506_32805 );
xor \U$34453 ( \42453_42753 , \42448_42748 , \42452_42752 );
and \U$34454 ( \42454_42754 , \30500_30802 , \32503_32802 );
xor \U$34455 ( \42455_42755 , \42453_42753 , \42454_42754 );
xor \U$34456 ( \42456_42756 , \42447_42747 , \42455_42755 );
and \U$34457 ( \42457_42757 , \42106_42406 , \42110_42410 );
and \U$34458 ( \42458_42758 , \42110_42410 , \42122_42422 );
and \U$34459 ( \42459_42759 , \42106_42406 , \42122_42422 );
or \U$34460 ( \42460_42760 , \42457_42757 , \42458_42758 , \42459_42759 );
xor \U$34461 ( \42461_42761 , \42456_42756 , \42460_42760 );
and \U$34462 ( \42462_42762 , \42123_42423 , \42127_42427 );
and \U$34463 ( \42463_42763 , \42128_42428 , \42131_42431 );
or \U$34464 ( \42464_42764 , \42462_42762 , \42463_42763 );
xor \U$34465 ( \42465_42765 , \42461_42761 , \42464_42764 );
buf g9b57_GF_PartitionCandidate( \42466_42766_nG9b57 , \42465_42765 );
and \U$34466 ( \42467_42767 , \10402_10704 , \42466_42766_nG9b57 );
or \U$34467 ( \42468_42768 , \42441_42741 , \42467_42767 );
xor \U$34468 ( \42469_42769 , \10399_10703 , \42468_42768 );
buf \U$34469 ( \42470_42770 , \42469_42769 );
buf \U$34471 ( \42471_42771 , \42470_42770 );
xor \U$34472 ( \42472_42772 , \42440_42740 , \42471_42771 );
buf \U$34473 ( \42473_42773 , \42472_42772 );
xor \U$34474 ( \42474_42774 , \42428_42728 , \42473_42773 );
and \U$34475 ( \42475_42775 , \42022_42322 , \42028_42328 );
and \U$34476 ( \42476_42776 , \42022_42322 , \42035_42335 );
and \U$34477 ( \42477_42777 , \42028_42328 , \42035_42335 );
or \U$34478 ( \42478_42778 , \42475_42775 , \42476_42776 , \42477_42777 );
buf \U$34479 ( \42479_42779 , \42478_42778 );
xor \U$34480 ( \42480_42780 , \42474_42774 , \42479_42779 );
buf \U$34481 ( \42481_42781 , \42480_42780 );
xor \U$34482 ( \42482_42782 , \42423_42723 , \42481_42781 );
and \U$34483 ( \42483_42783 , \42210_42510 , \42215_42515 );
and \U$34484 ( \42484_42784 , \42210_42510 , \42221_42521 );
and \U$34485 ( \42485_42785 , \42215_42515 , \42221_42521 );
or \U$34486 ( \42486_42786 , \42483_42783 , \42484_42784 , \42485_42785 );
buf \U$34487 ( \42487_42787 , \42486_42786 );
xor \U$34488 ( \42488_42788 , \42482_42782 , \42487_42787 );
buf \U$34489 ( \42489_42789 , \42488_42788 );
xor \U$34490 ( \42490_42790 , \42351_42651 , \42489_42789 );
and \U$34491 ( \42491_42791 , \42246_42546 , \42490_42790 );
and \U$34493 ( \42492_42792 , \42240_42540 , \42245_42545 );
or \U$34495 ( \42493_42793 , 1'b0 , \42492_42792 , 1'b0 );
xor \U$34496 ( \42494_42794 , \42491_42791 , \42493_42793 );
and \U$34498 ( \42495_42795 , \42233_42533 , \42239_42539 );
and \U$34499 ( \42496_42796 , \42235_42535 , \42239_42539 );
or \U$34500 ( \42497_42797 , 1'b0 , \42495_42795 , \42496_42796 );
xor \U$34501 ( \42498_42798 , \42494_42794 , \42497_42797 );
xor \U$34508 ( \42499_42799 , \42498_42798 , 1'b0 );
and \U$34509 ( \42500_42800 , \42345_42645 , \42350_42650 );
and \U$34510 ( \42501_42801 , \42345_42645 , \42489_42789 );
and \U$34511 ( \42502_42802 , \42350_42650 , \42489_42789 );
or \U$34512 ( \42503_42803 , \42500_42800 , \42501_42801 , \42502_42802 );
xor \U$34513 ( \42504_42804 , \42499_42799 , \42503_42803 );
and \U$34514 ( \42505_42805 , \42251_42551 , \42256_42556 );
and \U$34515 ( \42506_42806 , \42251_42551 , \42343_42643 );
and \U$34516 ( \42507_42807 , \42256_42556 , \42343_42643 );
or \U$34517 ( \42508_42808 , \42505_42805 , \42506_42806 , \42507_42807 );
buf \U$34518 ( \42509_42809 , \42508_42808 );
and \U$34519 ( \42510_42810 , \42262_42562 , \42335_42635 );
and \U$34520 ( \42511_42811 , \42262_42562 , \42341_42641 );
and \U$34521 ( \42512_42812 , \42335_42635 , \42341_42641 );
or \U$34522 ( \42513_42813 , \42510_42810 , \42511_42811 , \42512_42812 );
buf \U$34523 ( \42514_42814 , \42513_42813 );
and \U$34524 ( \42515_42815 , \42380_42680 , \42386_42686 );
and \U$34525 ( \42516_42816 , \42380_42680 , \42393_42693 );
and \U$34526 ( \42517_42817 , \42386_42686 , \42393_42693 );
or \U$34527 ( \42518_42818 , \42515_42815 , \42516_42816 , \42517_42817 );
buf \U$34528 ( \42519_42819 , \42518_42818 );
and \U$34529 ( \42520_42820 , \17437_17297 , \39034_39334_nG9b7b );
and \U$34530 ( \42521_42821 , \16995_17294 , \39291_39591_nG9b78 );
or \U$34531 ( \42522_42822 , \42520_42820 , \42521_42821 );
xor \U$34532 ( \42523_42823 , \16994_17293 , \42522_42822 );
buf \U$34533 ( \42524_42824 , \42523_42823 );
buf \U$34535 ( \42525_42825 , \42524_42824 );
xor \U$34536 ( \42526_42826 , \42519_42819 , \42525_42825 );
and \U$34537 ( \42527_42827 , \10411_10707 , \42466_42766_nG9b57 );
and \U$34538 ( \42528_42828 , \42448_42748 , \42452_42752 );
and \U$34539 ( \42529_42829 , \42452_42752 , \42454_42754 );
and \U$34540 ( \42530_42830 , \42448_42748 , \42454_42754 );
or \U$34541 ( \42531_42831 , \42528_42828 , \42529_42829 , \42530_42830 );
and \U$34542 ( \42532_42832 , \32495_32794 , \32555_32854 );
not \U$34543 ( \42533_42833 , \42532_42832 );
xnor \U$34544 ( \42534_42834 , \42533_42833 , \32506_32805 );
xor \U$34545 ( \42535_42835 , \42531_42831 , \42534_42834 );
and \U$34546 ( \42536_42836 , \31752_32054 , \32503_32802 );
not \U$34547 ( \42537_42837 , \42536_42836 );
xor \U$34548 ( \42538_42838 , \42535_42835 , \42537_42837 );
and \U$34549 ( \42539_42839 , \42445_42745 , \42446_42746 );
and \U$34550 ( \42540_42840 , \42446_42746 , \42455_42755 );
and \U$34551 ( \42541_42841 , \42445_42745 , \42455_42755 );
or \U$34552 ( \42542_42842 , \42539_42839 , \42540_42840 , \42541_42841 );
xor \U$34553 ( \42543_42843 , \42538_42838 , \42542_42842 );
and \U$34554 ( \42544_42844 , \42456_42756 , \42460_42760 );
and \U$34555 ( \42545_42845 , \42461_42761 , \42464_42764 );
or \U$34556 ( \42546_42846 , \42544_42844 , \42545_42845 );
xor \U$34557 ( \42547_42847 , \42543_42843 , \42546_42846 );
buf g9b54_GF_PartitionCandidate( \42548_42848_nG9b54 , \42547_42847 );
and \U$34558 ( \42549_42849 , \10402_10704 , \42548_42848_nG9b54 );
or \U$34559 ( \42550_42850 , \42527_42827 , \42549_42849 );
xor \U$34560 ( \42551_42851 , \10399_10703 , \42550_42850 );
buf \U$34561 ( \42552_42852 , \42551_42851 );
buf \U$34563 ( \42553_42853 , \42552_42852 );
xor \U$34564 ( \42554_42854 , \42526_42826 , \42553_42853 );
buf \U$34565 ( \42555_42855 , \42554_42854 );
and \U$34566 ( \42556_42856 , \42433_42733 , \42439_42739 );
and \U$34567 ( \42557_42857 , \42433_42733 , \42471_42771 );
and \U$34568 ( \42558_42858 , \42439_42739 , \42471_42771 );
or \U$34569 ( \42559_42859 , \42556_42856 , \42557_42857 , \42558_42858 );
buf \U$34570 ( \42560_42860 , \42559_42859 );
xor \U$34571 ( \42561_42861 , \42555_42855 , \42560_42860 );
and \U$34572 ( \42562_42862 , \42402_42702 , \42407_42707 );
and \U$34573 ( \42563_42863 , \42402_42702 , \42413_42713 );
and \U$34574 ( \42564_42864 , \42407_42707 , \42413_42713 );
or \U$34575 ( \42565_42865 , \42562_42862 , \42563_42863 , \42564_42864 );
buf \U$34576 ( \42566_42866 , \42565_42865 );
xor \U$34577 ( \42567_42867 , \42561_42861 , \42566_42866 );
buf \U$34578 ( \42568_42868 , \42567_42867 );
and \U$34579 ( \42569_42869 , \28946_28118 , \33994_34294_nG9ba5 );
and \U$34580 ( \42570_42870 , \27816_28115 , \34343_34643_nG9ba2 );
or \U$34581 ( \42571_42871 , \42569_42869 , \42570_42870 );
xor \U$34582 ( \42572_42872 , \27815_28114 , \42571_42871 );
buf \U$34583 ( \42573_42873 , \42572_42872 );
buf \U$34585 ( \42574_42874 , \42573_42873 );
and \U$34586 ( \42575_42875 , \18908_18702 , \38363_38663_nG9b81 );
and \U$34587 ( \42576_42876 , \18400_18699 , \38668_38968_nG9b7e );
or \U$34588 ( \42577_42877 , \42575_42875 , \42576_42876 );
xor \U$34589 ( \42578_42878 , \18399_18698 , \42577_42877 );
buf \U$34590 ( \42579_42879 , \42578_42878 );
buf \U$34592 ( \42580_42880 , \42579_42879 );
xor \U$34593 ( \42581_42881 , \42574_42874 , \42580_42880 );
and \U$34594 ( \42582_42882 , \13431_13370 , \40740_41040_nG9b69 );
and \U$34595 ( \42583_42883 , \13068_13367 , \41081_41381_nG9b66 );
or \U$34596 ( \42584_42884 , \42582_42882 , \42583_42883 );
xor \U$34597 ( \42585_42885 , \13067_13366 , \42584_42884 );
buf \U$34598 ( \42586_42886 , \42585_42885 );
buf \U$34600 ( \42587_42887 , \42586_42886 );
xor \U$34601 ( \42588_42888 , \42581_42881 , \42587_42887 );
buf \U$34602 ( \42589_42889 , \42588_42888 );
and \U$34603 ( \42590_42890 , \42267_42567 , \42273_42573 );
buf \U$34604 ( \42591_42891 , \42590_42890 );
and \U$34606 ( \42592_42892 , \32617_32916 , \31877_32179_nG9bb4 );
or \U$34607 ( \42593_42893 , 1'b0 , \42592_42892 );
xor \U$34608 ( \42594_42894 , 1'b0 , \42593_42893 );
buf \U$34609 ( \42595_42895 , \42594_42894 );
buf \U$34611 ( \42596_42896 , \42595_42895 );
and \U$34612 ( \42597_42897 , \30670_29853 , \33313_33613_nG9bab );
and \U$34613 ( \42598_42898 , \29551_29850 , \33741_34041_nG9ba8 );
or \U$34614 ( \42599_42899 , \42597_42897 , \42598_42898 );
xor \U$34615 ( \42600_42900 , \29550_29849 , \42599_42899 );
buf \U$34616 ( \42601_42901 , \42600_42900 );
buf \U$34618 ( \42602_42902 , \42601_42901 );
xor \U$34619 ( \42603_42903 , \42596_42896 , \42602_42902 );
buf \U$34620 ( \42604_42904 , \42603_42903 );
xor \U$34621 ( \42605_42905 , \42591_42891 , \42604_42904 );
and \U$34622 ( \42606_42906 , \20353_20155 , \37674_37974_nG9b87 );
and \U$34623 ( \42607_42907 , \19853_20152 , \38037_38337_nG9b84 );
or \U$34624 ( \42608_42908 , \42606_42906 , \42607_42907 );
xor \U$34625 ( \42609_42909 , \19852_20151 , \42608_42908 );
buf \U$34626 ( \42610_42910 , \42609_42909 );
buf \U$34628 ( \42611_42911 , \42610_42910 );
xor \U$34629 ( \42612_42912 , \42605_42905 , \42611_42911 );
buf \U$34630 ( \42613_42913 , \42612_42912 );
xor \U$34631 ( \42614_42914 , \42589_42889 , \42613_42913 );
and \U$34632 ( \42615_42915 , \23495_23201 , \36289_36589_nG9b93 );
and \U$34633 ( \42616_42916 , \22899_23198 , \36686_36986_nG9b90 );
or \U$34634 ( \42617_42917 , \42615_42915 , \42616_42916 );
xor \U$34635 ( \42618_42918 , \22898_23197 , \42617_42917 );
buf \U$34636 ( \42619_42919 , \42618_42918 );
buf \U$34638 ( \42620_42920 , \42619_42919 );
and \U$34639 ( \42621_42921 , \21908_21658 , \36950_37250_nG9b8d );
and \U$34640 ( \42622_42922 , \21356_21655 , \37307_37607_nG9b8a );
or \U$34641 ( \42623_42923 , \42621_42921 , \42622_42922 );
xor \U$34642 ( \42624_42924 , \21355_21654 , \42623_42923 );
buf \U$34643 ( \42625_42925 , \42624_42924 );
buf \U$34645 ( \42626_42926 , \42625_42925 );
xor \U$34646 ( \42627_42927 , \42620_42920 , \42626_42926 );
and \U$34647 ( \42628_42928 , \14710_14631 , \40152_40452_nG9b6f );
and \U$34648 ( \42629_42929 , \14329_14628 , \40543_40843_nG9b6c );
or \U$34649 ( \42630_42930 , \42628_42928 , \42629_42929 );
xor \U$34650 ( \42631_42931 , \14328_14627 , \42630_42930 );
buf \U$34651 ( \42632_42932 , \42631_42931 );
buf \U$34653 ( \42633_42933 , \42632_42932 );
xor \U$34654 ( \42634_42934 , \42627_42927 , \42633_42933 );
buf \U$34655 ( \42635_42935 , \42634_42934 );
xor \U$34656 ( \42636_42936 , \42614_42914 , \42635_42935 );
buf \U$34657 ( \42637_42937 , \42636_42936 );
xor \U$34658 ( \42638_42938 , \42568_42868 , \42637_42937 );
and \U$34659 ( \42639_42939 , \42290_42590 , \42311_42611 );
and \U$34660 ( \42640_42940 , \42290_42590 , \42333_42633 );
and \U$34661 ( \42641_42941 , \42311_42611 , \42333_42633 );
or \U$34662 ( \42642_42942 , \42639_42939 , \42640_42940 , \42641_42941 );
buf \U$34663 ( \42643_42943 , \42642_42942 );
xor \U$34664 ( \42644_42944 , \42638_42938 , \42643_42943 );
buf \U$34665 ( \42645_42945 , \42644_42944 );
xor \U$34666 ( \42646_42946 , \42514_42814 , \42645_42945 );
and \U$34667 ( \42647_42947 , \42423_42723 , \42481_42781 );
and \U$34668 ( \42648_42948 , \42423_42723 , \42487_42787 );
and \U$34669 ( \42649_42949 , \42481_42781 , \42487_42787 );
or \U$34670 ( \42650_42950 , \42647_42947 , \42648_42948 , \42649_42949 );
buf \U$34671 ( \42651_42951 , \42650_42950 );
xor \U$34672 ( \42652_42952 , \42646_42946 , \42651_42951 );
buf \U$34673 ( \42653_42953 , \42652_42952 );
xor \U$34674 ( \42654_42954 , \42509_42809 , \42653_42953 );
and \U$34675 ( \42655_42955 , \42275_42575 , \42281_42581 );
and \U$34676 ( \42656_42956 , \42275_42575 , \42288_42588 );
and \U$34677 ( \42657_42957 , \42281_42581 , \42288_42588 );
or \U$34678 ( \42658_42958 , \42655_42955 , \42656_42956 , \42657_42957 );
buf \U$34679 ( \42659_42959 , \42658_42958 );
and \U$34680 ( \42660_42960 , \42296_42596 , \42302_42602 );
and \U$34681 ( \42661_42961 , \42296_42596 , \42309_42609 );
and \U$34682 ( \42662_42962 , \42302_42602 , \42309_42609 );
or \U$34683 ( \42663_42963 , \42660_42960 , \42661_42961 , \42662_42962 );
buf \U$34684 ( \42664_42964 , \42663_42963 );
xor \U$34685 ( \42665_42965 , \42659_42959 , \42664_42964 );
and \U$34686 ( \42666_42966 , \42362_42662 , \42368_42668 );
and \U$34687 ( \42667_42967 , \42362_42662 , \42375_42675 );
and \U$34688 ( \42668_42968 , \42368_42668 , \42375_42675 );
or \U$34689 ( \42669_42969 , \42666_42966 , \42667_42967 , \42668_42968 );
buf \U$34690 ( \42670_42970 , \42669_42969 );
xor \U$34691 ( \42671_42971 , \42665_42965 , \42670_42970 );
buf \U$34692 ( \42672_42972 , \42671_42971 );
and \U$34693 ( \42673_42973 , \42356_42656 , \42377_42677 );
and \U$34694 ( \42674_42974 , \42356_42656 , \42395_42695 );
and \U$34695 ( \42675_42975 , \42377_42677 , \42395_42695 );
or \U$34696 ( \42676_42976 , \42673_42973 , \42674_42974 , \42675_42975 );
buf \U$34697 ( \42677_42977 , \42676_42976 );
xor \U$34698 ( \42678_42978 , \42672_42972 , \42677_42977 );
and \U$34699 ( \42679_42979 , \16405_15940 , \39663_39963_nG9b75 );
and \U$34700 ( \42680_42980 , \15638_15937 , \39904_40204_nG9b72 );
or \U$34701 ( \42681_42981 , \42679_42979 , \42680_42980 );
xor \U$34702 ( \42682_42982 , \15637_15936 , \42681_42981 );
buf \U$34703 ( \42683_42983 , \42682_42982 );
buf \U$34705 ( \42684_42984 , \42683_42983 );
and \U$34706 ( \42685_42985 , \12183_12157 , \41385_41685_nG9b63 );
and \U$34707 ( \42686_42986 , \11855_12154 , \41663_41963_nG9b60 );
or \U$34708 ( \42687_42987 , \42685_42985 , \42686_42986 );
xor \U$34709 ( \42688_42988 , \11854_12153 , \42687_42987 );
buf \U$34710 ( \42689_42989 , \42688_42988 );
buf \U$34712 ( \42690_42990 , \42689_42989 );
xor \U$34713 ( \42691_42991 , \42684_42984 , \42690_42990 );
and \U$34714 ( \42692_42992 , \10996_10421 , \41901_42201_nG9b5d );
and \U$34715 ( \42693_42993 , \10119_10418 , \42133_42433_nG9b5a );
or \U$34716 ( \42694_42994 , \42692_42992 , \42693_42993 );
xor \U$34717 ( \42695_42995 , \10118_10417 , \42694_42994 );
buf \U$34718 ( \42696_42996 , \42695_42995 );
buf \U$34720 ( \42697_42997 , \42696_42996 );
xor \U$34721 ( \42698_42998 , \42691_42991 , \42697_42997 );
buf \U$34722 ( \42699_42999 , \42698_42998 );
and \U$34723 ( \42700_43000 , \31989_31636 , \32589_32888_nG9bb1 );
and \U$34724 ( \42701_43001 , \31334_31633 , \32881_33181_nG9bae );
or \U$34725 ( \42702_43002 , \42700_43000 , \42701_43001 );
xor \U$34726 ( \42703_43003 , \31333_31632 , \42702_43002 );
buf \U$34727 ( \42704_43004 , \42703_43003 );
buf \U$34729 ( \42705_43005 , \42704_43004 );
and \U$34730 ( \42706_43006 , \27141_26431 , \34794_35094_nG9b9f );
and \U$34731 ( \42707_43007 , \26129_26428 , \35270_35570_nG9b9c );
or \U$34732 ( \42708_43008 , \42706_43006 , \42707_43007 );
xor \U$34733 ( \42709_43009 , \26128_26427 , \42708_43008 );
buf \U$34734 ( \42710_43010 , \42709_43009 );
buf \U$34736 ( \42711_43011 , \42710_43010 );
xor \U$34737 ( \42712_43012 , \42705_43005 , \42711_43011 );
and \U$34738 ( \42713_43013 , \25044_24792 , \35501_35801_nG9b99 );
and \U$34739 ( \42714_43014 , \24490_24789 , \35872_36172_nG9b96 );
or \U$34740 ( \42715_43015 , \42713_43013 , \42714_43014 );
xor \U$34741 ( \42716_43016 , \24489_24788 , \42715_43015 );
buf \U$34742 ( \42717_43017 , \42716_43016 );
buf \U$34744 ( \42718_43018 , \42717_43017 );
xor \U$34745 ( \42719_43019 , \42712_43012 , \42718_43018 );
buf \U$34746 ( \42720_43020 , \42719_43019 );
xor \U$34747 ( \42721_43021 , \42699_42999 , \42720_43020 );
and \U$34748 ( \42722_43022 , \42318_42618 , \42324_42624 );
and \U$34749 ( \42723_43023 , \42318_42618 , \42331_42631 );
and \U$34750 ( \42724_43024 , \42324_42624 , \42331_42631 );
or \U$34751 ( \42725_43025 , \42722_43022 , \42723_43023 , \42724_43024 );
buf \U$34752 ( \42726_43026 , \42725_43025 );
xor \U$34753 ( \42727_43027 , \42721_43021 , \42726_43026 );
buf \U$34754 ( \42728_43028 , \42727_43027 );
xor \U$34755 ( \42729_43029 , \42678_42978 , \42728_43028 );
buf \U$34756 ( \42730_43030 , \42729_43029 );
and \U$34757 ( \42731_43031 , \42397_42697 , \42415_42715 );
and \U$34758 ( \42732_43032 , \42397_42697 , \42421_42721 );
and \U$34759 ( \42733_43033 , \42415_42715 , \42421_42721 );
or \U$34760 ( \42734_43034 , \42731_43031 , \42732_43032 , \42733_43033 );
buf \U$34761 ( \42735_43035 , \42734_43034 );
xor \U$34762 ( \42736_43036 , \42730_43030 , \42735_43035 );
and \U$34763 ( \42737_43037 , \42428_42728 , \42473_42773 );
and \U$34764 ( \42738_43038 , \42428_42728 , \42479_42779 );
and \U$34765 ( \42739_43039 , \42473_42773 , \42479_42779 );
or \U$34766 ( \42740_43040 , \42737_43037 , \42738_43038 , \42739_43039 );
buf \U$34767 ( \42741_43041 , \42740_43040 );
xor \U$34768 ( \42742_43042 , \42736_43036 , \42741_43041 );
buf \U$34769 ( \42743_43043 , \42742_43042 );
xor \U$34770 ( \42744_43044 , \42654_42954 , \42743_43043 );
and \U$34771 ( \42745_43045 , \42504_42804 , \42744_43044 );
and \U$34773 ( \42746_43046 , \42498_42798 , \42503_42803 );
or \U$34775 ( \42747_43047 , 1'b0 , \42746_43046 , 1'b0 );
xor \U$34776 ( \42748_43048 , \42745_43045 , \42747_43047 );
and \U$34778 ( \42749_43049 , \42491_42791 , \42497_42797 );
and \U$34779 ( \42750_43050 , \42493_42793 , \42497_42797 );
or \U$34780 ( \42751_43051 , 1'b0 , \42749_43049 , \42750_43050 );
xor \U$34781 ( \42752_43052 , \42748_43048 , \42751_43051 );
xor \U$34788 ( \42753_43053 , \42752_43052 , 1'b0 );
and \U$34789 ( \42754_43054 , \42509_42809 , \42653_42953 );
and \U$34790 ( \42755_43055 , \42509_42809 , \42743_43043 );
and \U$34791 ( \42756_43056 , \42653_42953 , \42743_43043 );
or \U$34792 ( \42757_43057 , \42754_43054 , \42755_43055 , \42756_43056 );
xor \U$34793 ( \42758_43058 , \42753_43053 , \42757_43057 );
and \U$34794 ( \42759_43059 , \42699_42999 , \42720_43020 );
and \U$34795 ( \42760_43060 , \42699_42999 , \42726_43026 );
and \U$34796 ( \42761_43061 , \42720_43020 , \42726_43026 );
or \U$34797 ( \42762_43062 , \42759_43059 , \42760_43060 , \42761_43061 );
buf \U$34798 ( \42763_43063 , \42762_43062 );
and \U$34799 ( \42764_43064 , \42591_42891 , \42604_42904 );
and \U$34800 ( \42765_43065 , \42591_42891 , \42611_42911 );
and \U$34801 ( \42766_43066 , \42604_42904 , \42611_42911 );
or \U$34802 ( \42767_43067 , \42764_43064 , \42765_43065 , \42766_43066 );
buf \U$34803 ( \42768_43068 , \42767_43067 );
and \U$34804 ( \42769_43069 , \42574_42874 , \42580_42880 );
and \U$34805 ( \42770_43070 , \42574_42874 , \42587_42887 );
and \U$34806 ( \42771_43071 , \42580_42880 , \42587_42887 );
or \U$34807 ( \42772_43072 , \42769_43069 , \42770_43070 , \42771_43071 );
buf \U$34808 ( \42773_43073 , \42772_43072 );
xor \U$34809 ( \42774_43074 , \42768_43068 , \42773_43073 );
and \U$34810 ( \42775_43075 , \30670_29853 , \33741_34041_nG9ba8 );
and \U$34811 ( \42776_43076 , \29551_29850 , \33994_34294_nG9ba5 );
or \U$34812 ( \42777_43077 , \42775_43075 , \42776_43076 );
xor \U$34813 ( \42778_43078 , \29550_29849 , \42777_43077 );
buf \U$34814 ( \42779_43079 , \42778_43078 );
buf \U$34816 ( \42780_43080 , \42779_43079 );
and \U$34817 ( \42781_43081 , \28946_28118 , \34343_34643_nG9ba2 );
and \U$34818 ( \42782_43082 , \27816_28115 , \34794_35094_nG9b9f );
or \U$34819 ( \42783_43083 , \42781_43081 , \42782_43082 );
xor \U$34820 ( \42784_43084 , \27815_28114 , \42783_43083 );
buf \U$34821 ( \42785_43085 , \42784_43084 );
buf \U$34823 ( \42786_43086 , \42785_43085 );
xor \U$34824 ( \42787_43087 , \42780_43080 , \42786_43086 );
and \U$34825 ( \42788_43088 , \27141_26431 , \35270_35570_nG9b9c );
and \U$34826 ( \42789_43089 , \26129_26428 , \35501_35801_nG9b99 );
or \U$34827 ( \42790_43090 , \42788_43088 , \42789_43089 );
xor \U$34828 ( \42791_43091 , \26128_26427 , \42790_43090 );
buf \U$34829 ( \42792_43092 , \42791_43091 );
buf \U$34831 ( \42793_43093 , \42792_43092 );
xor \U$34832 ( \42794_43094 , \42787_43087 , \42793_43093 );
buf \U$34833 ( \42795_43095 , \42794_43094 );
xor \U$34834 ( \42796_43096 , \42774_43074 , \42795_43095 );
buf \U$34835 ( \42797_43097 , \42796_43096 );
xor \U$34836 ( \42798_43098 , \42763_43063 , \42797_43097 );
and \U$34837 ( \42799_43099 , \25044_24792 , \35872_36172_nG9b96 );
and \U$34838 ( \42800_43100 , \24490_24789 , \36289_36589_nG9b93 );
or \U$34839 ( \42801_43101 , \42799_43099 , \42800_43100 );
xor \U$34840 ( \42802_43102 , \24489_24788 , \42801_43101 );
buf \U$34841 ( \42803_43103 , \42802_43102 );
buf \U$34843 ( \42804_43104 , \42803_43103 );
and \U$34844 ( \42805_43105 , \17437_17297 , \39291_39591_nG9b78 );
and \U$34845 ( \42806_43106 , \16995_17294 , \39663_39963_nG9b75 );
or \U$34846 ( \42807_43107 , \42805_43105 , \42806_43106 );
xor \U$34847 ( \42808_43108 , \16994_17293 , \42807_43107 );
buf \U$34848 ( \42809_43109 , \42808_43108 );
buf \U$34850 ( \42810_43110 , \42809_43109 );
xor \U$34851 ( \42811_43111 , \42804_43104 , \42810_43110 );
and \U$34852 ( \42812_43112 , \16405_15940 , \39904_40204_nG9b72 );
and \U$34853 ( \42813_43113 , \15638_15937 , \40152_40452_nG9b6f );
or \U$34854 ( \42814_43114 , \42812_43112 , \42813_43113 );
xor \U$34855 ( \42815_43115 , \15637_15936 , \42814_43114 );
buf \U$34856 ( \42816_43116 , \42815_43115 );
buf \U$34858 ( \42817_43117 , \42816_43116 );
xor \U$34859 ( \42818_43118 , \42811_43111 , \42817_43117 );
buf \U$34860 ( \42819_43119 , \42818_43118 );
and \U$34861 ( \42820_43120 , \42684_42984 , \42690_42990 );
and \U$34862 ( \42821_43121 , \42684_42984 , \42697_42997 );
and \U$34863 ( \42822_43122 , \42690_42990 , \42697_42997 );
or \U$34864 ( \42823_43123 , \42820_43120 , \42821_43121 , \42822_43122 );
buf \U$34865 ( \42824_43124 , \42823_43123 );
xor \U$34866 ( \42825_43125 , \42819_43119 , \42824_43124 );
and \U$34867 ( \42826_43126 , \42620_42920 , \42626_42926 );
and \U$34868 ( \42827_43127 , \42620_42920 , \42633_42933 );
and \U$34869 ( \42828_43128 , \42626_42926 , \42633_42933 );
or \U$34870 ( \42829_43129 , \42826_43126 , \42827_43127 , \42828_43128 );
buf \U$34871 ( \42830_43130 , \42829_43129 );
xor \U$34872 ( \42831_43131 , \42825_43125 , \42830_43130 );
buf \U$34873 ( \42832_43132 , \42831_43131 );
xor \U$34874 ( \42833_43133 , \42798_43098 , \42832_43132 );
buf \U$34875 ( \42834_43134 , \42833_43133 );
and \U$34876 ( \42835_43135 , \42672_42972 , \42677_42977 );
and \U$34877 ( \42836_43136 , \42672_42972 , \42728_43028 );
and \U$34878 ( \42837_43137 , \42677_42977 , \42728_43028 );
or \U$34879 ( \42838_43138 , \42835_43135 , \42836_43136 , \42837_43137 );
buf \U$34880 ( \42839_43139 , \42838_43138 );
xor \U$34881 ( \42840_43140 , \42834_43134 , \42839_43139 );
and \U$34882 ( \42841_43141 , \42555_42855 , \42560_42860 );
and \U$34883 ( \42842_43142 , \42555_42855 , \42566_42866 );
and \U$34884 ( \42843_43143 , \42560_42860 , \42566_42866 );
or \U$34885 ( \42844_43144 , \42841_43141 , \42842_43142 , \42843_43143 );
buf \U$34886 ( \42845_43145 , \42844_43144 );
xor \U$34887 ( \42846_43146 , \42840_43140 , \42845_43145 );
buf \U$34888 ( \42847_43147 , \42846_43146 );
and \U$34889 ( \42848_43148 , \42568_42868 , \42637_42937 );
and \U$34890 ( \42849_43149 , \42568_42868 , \42643_42943 );
and \U$34891 ( \42850_43150 , \42637_42937 , \42643_42943 );
or \U$34892 ( \42851_43151 , \42848_43148 , \42849_43149 , \42850_43150 );
buf \U$34893 ( \42852_43152 , \42851_43151 );
xor \U$34894 ( \42853_43153 , \42847_43147 , \42852_43152 );
and \U$34895 ( \42854_43154 , \42659_42959 , \42664_42964 );
and \U$34896 ( \42855_43155 , \42659_42959 , \42670_42970 );
and \U$34897 ( \42856_43156 , \42664_42964 , \42670_42970 );
or \U$34898 ( \42857_43157 , \42854_43154 , \42855_43155 , \42856_43156 );
buf \U$34899 ( \42858_43158 , \42857_43157 );
and \U$34900 ( \42859_43159 , \42705_43005 , \42711_43011 );
and \U$34901 ( \42860_43160 , \42705_43005 , \42718_43018 );
and \U$34902 ( \42861_43161 , \42711_43011 , \42718_43018 );
or \U$34903 ( \42862_43162 , \42859_43159 , \42860_43160 , \42861_43161 );
buf \U$34904 ( \42863_43163 , \42862_43162 );
and \U$34905 ( \42864_43164 , \10411_10707 , \42548_42848_nG9b54 );
and \U$34906 ( \42865_43165 , \42531_42831 , \42534_42834 );
and \U$34907 ( \42866_43166 , \42534_42834 , \42537_42837 );
and \U$34908 ( \42867_43167 , \42531_42831 , \42537_42837 );
or \U$34909 ( \42868_43168 , \42865_43165 , \42866_43166 , \42867_43167 );
buf \U$34910 ( \42869_43169 , \42536_42836 );
not \U$34911 ( \42870_43170 , \32506_32805 );
xor \U$34912 ( \42871_43171 , \42869_43169 , \42870_43170 );
and \U$34913 ( \42872_43172 , \32495_32794 , \32503_32802 );
xor \U$34914 ( \42873_43173 , \42871_43171 , \42872_43172 );
xor \U$34915 ( \42874_43174 , \42868_43168 , \42873_43173 );
and \U$34916 ( \42875_43175 , \42538_42838 , \42542_42842 );
and \U$34917 ( \42876_43176 , \42543_42843 , \42546_42846 );
or \U$34918 ( \42877_43177 , \42875_43175 , \42876_43176 );
xor \U$34919 ( \42878_43178 , \42874_43174 , \42877_43177 );
buf g9b51_GF_PartitionCandidate( \42879_43179_nG9b51 , \42878_43178 );
and \U$34920 ( \42880_43180 , \10402_10704 , \42879_43179_nG9b51 );
or \U$34921 ( \42881_43181 , \42864_43164 , \42880_43180 );
xor \U$34922 ( \42882_43182 , \10399_10703 , \42881_43181 );
buf \U$34923 ( \42883_43183 , \42882_43182 );
buf \U$34925 ( \42884_43184 , \42883_43183 );
xor \U$34926 ( \42885_43185 , \42863_43163 , \42884_43184 );
and \U$34927 ( \42886_43186 , \10996_10421 , \42133_42433_nG9b5a );
and \U$34928 ( \42887_43187 , \10119_10418 , \42466_42766_nG9b57 );
or \U$34929 ( \42888_43188 , \42886_43186 , \42887_43187 );
xor \U$34930 ( \42889_43189 , \10118_10417 , \42888_43188 );
buf \U$34931 ( \42890_43190 , \42889_43189 );
buf \U$34933 ( \42891_43191 , \42890_43190 );
xor \U$34934 ( \42892_43192 , \42885_43185 , \42891_43191 );
buf \U$34935 ( \42893_43193 , \42892_43192 );
xor \U$34936 ( \42894_43194 , \42858_43158 , \42893_43193 );
and \U$34937 ( \42895_43195 , \42519_42819 , \42525_42825 );
and \U$34938 ( \42896_43196 , \42519_42819 , \42553_42853 );
and \U$34939 ( \42897_43197 , \42525_42825 , \42553_42853 );
or \U$34940 ( \42898_43198 , \42895_43195 , \42896_43196 , \42897_43197 );
buf \U$34941 ( \42899_43199 , \42898_43198 );
xor \U$34942 ( \42900_43200 , \42894_43194 , \42899_43199 );
buf \U$34943 ( \42901_43201 , \42900_43200 );
and \U$34944 ( \42902_43202 , \42589_42889 , \42613_42913 );
and \U$34945 ( \42903_43203 , \42589_42889 , \42635_42935 );
and \U$34946 ( \42904_43204 , \42613_42913 , \42635_42935 );
or \U$34947 ( \42905_43205 , \42902_43202 , \42903_43203 , \42904_43204 );
buf \U$34948 ( \42906_43206 , \42905_43205 );
xor \U$34949 ( \42907_43207 , \42901_43201 , \42906_43206 );
and \U$34951 ( \42908_43208 , \32617_32916 , \32589_32888_nG9bb1 );
or \U$34952 ( \42909_43209 , 1'b0 , \42908_43208 );
xor \U$34953 ( \42910_43210 , 1'b0 , \42909_43209 );
buf \U$34954 ( \42911_43211 , \42910_43210 );
buf \U$34956 ( \42912_43212 , \42911_43211 );
and \U$34957 ( \42913_43213 , \31989_31636 , \32881_33181_nG9bae );
and \U$34958 ( \42914_43214 , \31334_31633 , \33313_33613_nG9bab );
or \U$34959 ( \42915_43215 , \42913_43213 , \42914_43214 );
xor \U$34960 ( \42916_43216 , \31333_31632 , \42915_43215 );
buf \U$34961 ( \42917_43217 , \42916_43216 );
buf \U$34963 ( \42918_43218 , \42917_43217 );
xor \U$34964 ( \42919_43219 , \42912_43212 , \42918_43218 );
buf \U$34965 ( \42920_43220 , \42919_43219 );
and \U$34966 ( \42921_43221 , \18908_18702 , \38668_38968_nG9b7e );
and \U$34967 ( \42922_43222 , \18400_18699 , \39034_39334_nG9b7b );
or \U$34968 ( \42923_43223 , \42921_43221 , \42922_43222 );
xor \U$34969 ( \42924_43224 , \18399_18698 , \42923_43223 );
buf \U$34970 ( \42925_43225 , \42924_43224 );
buf \U$34972 ( \42926_43226 , \42925_43225 );
xor \U$34973 ( \42927_43227 , \42920_43220 , \42926_43226 );
and \U$34974 ( \42928_43228 , \13431_13370 , \41081_41381_nG9b66 );
and \U$34975 ( \42929_43229 , \13068_13367 , \41385_41685_nG9b63 );
or \U$34976 ( \42930_43230 , \42928_43228 , \42929_43229 );
xor \U$34977 ( \42931_43231 , \13067_13366 , \42930_43230 );
buf \U$34978 ( \42932_43232 , \42931_43231 );
buf \U$34980 ( \42933_43233 , \42932_43232 );
xor \U$34981 ( \42934_43234 , \42927_43227 , \42933_43233 );
buf \U$34982 ( \42935_43235 , \42934_43234 );
and \U$34983 ( \42936_43236 , \23495_23201 , \36686_36986_nG9b90 );
and \U$34984 ( \42937_43237 , \22899_23198 , \36950_37250_nG9b8d );
or \U$34985 ( \42938_43238 , \42936_43236 , \42937_43237 );
xor \U$34986 ( \42939_43239 , \22898_23197 , \42938_43238 );
buf \U$34987 ( \42940_43240 , \42939_43239 );
buf \U$34989 ( \42941_43241 , \42940_43240 );
and \U$34990 ( \42942_43242 , \21908_21658 , \37307_37607_nG9b8a );
and \U$34991 ( \42943_43243 , \21356_21655 , \37674_37974_nG9b87 );
or \U$34992 ( \42944_43244 , \42942_43242 , \42943_43243 );
xor \U$34993 ( \42945_43245 , \21355_21654 , \42944_43244 );
buf \U$34994 ( \42946_43246 , \42945_43245 );
buf \U$34996 ( \42947_43247 , \42946_43246 );
xor \U$34997 ( \42948_43248 , \42941_43241 , \42947_43247 );
and \U$34998 ( \42949_43249 , \12183_12157 , \41663_41963_nG9b60 );
and \U$34999 ( \42950_43250 , \11855_12154 , \41901_42201_nG9b5d );
or \U$35000 ( \42951_43251 , \42949_43249 , \42950_43250 );
xor \U$35001 ( \42952_43252 , \11854_12153 , \42951_43251 );
buf \U$35002 ( \42953_43253 , \42952_43252 );
buf \U$35004 ( \42954_43254 , \42953_43253 );
xor \U$35005 ( \42955_43255 , \42948_43248 , \42954_43254 );
buf \U$35006 ( \42956_43256 , \42955_43255 );
xor \U$35007 ( \42957_43257 , \42935_43235 , \42956_43256 );
and \U$35008 ( \42958_43258 , \42596_42896 , \42602_42902 );
buf \U$35009 ( \42959_43259 , \42958_43258 );
and \U$35010 ( \42960_43260 , \20353_20155 , \38037_38337_nG9b84 );
and \U$35011 ( \42961_43261 , \19853_20152 , \38363_38663_nG9b81 );
or \U$35012 ( \42962_43262 , \42960_43260 , \42961_43261 );
xor \U$35013 ( \42963_43263 , \19852_20151 , \42962_43262 );
buf \U$35014 ( \42964_43264 , \42963_43263 );
buf \U$35016 ( \42965_43265 , \42964_43264 );
xor \U$35017 ( \42966_43266 , \42959_43259 , \42965_43265 );
and \U$35018 ( \42967_43267 , \14710_14631 , \40543_40843_nG9b6c );
and \U$35019 ( \42968_43268 , \14329_14628 , \40740_41040_nG9b69 );
or \U$35020 ( \42969_43269 , \42967_43267 , \42968_43268 );
xor \U$35021 ( \42970_43270 , \14328_14627 , \42969_43269 );
buf \U$35022 ( \42971_43271 , \42970_43270 );
buf \U$35024 ( \42972_43272 , \42971_43271 );
xor \U$35025 ( \42973_43273 , \42966_43266 , \42972_43272 );
buf \U$35026 ( \42974_43274 , \42973_43273 );
xor \U$35027 ( \42975_43275 , \42957_43257 , \42974_43274 );
buf \U$35028 ( \42976_43276 , \42975_43275 );
xor \U$35029 ( \42977_43277 , \42907_43207 , \42976_43276 );
buf \U$35030 ( \42978_43278 , \42977_43277 );
xor \U$35031 ( \42979_43279 , \42853_43153 , \42978_43278 );
buf \U$35032 ( \42980_43280 , \42979_43279 );
and \U$35033 ( \42981_43281 , \42514_42814 , \42645_42945 );
and \U$35034 ( \42982_43282 , \42514_42814 , \42651_42951 );
and \U$35035 ( \42983_43283 , \42645_42945 , \42651_42951 );
or \U$35036 ( \42984_43284 , \42981_43281 , \42982_43282 , \42983_43283 );
buf \U$35037 ( \42985_43285 , \42984_43284 );
xor \U$35038 ( \42986_43286 , \42980_43280 , \42985_43285 );
and \U$35039 ( \42987_43287 , \42730_43030 , \42735_43035 );
and \U$35040 ( \42988_43288 , \42730_43030 , \42741_43041 );
and \U$35041 ( \42989_43289 , \42735_43035 , \42741_43041 );
or \U$35042 ( \42990_43290 , \42987_43287 , \42988_43288 , \42989_43289 );
buf \U$35043 ( \42991_43291 , \42990_43290 );
xor \U$35044 ( \42992_43292 , \42986_43286 , \42991_43291 );
and \U$35045 ( \42993_43293 , \42758_43058 , \42992_43292 );
and \U$35047 ( \42994_43294 , \42752_43052 , \42757_43057 );
or \U$35049 ( \42995_43295 , 1'b0 , \42994_43294 , 1'b0 );
xor \U$35050 ( \42996_43296 , \42993_43293 , \42995_43295 );
and \U$35052 ( \42997_43297 , \42745_43045 , \42751_43051 );
and \U$35053 ( \42998_43298 , \42747_43047 , \42751_43051 );
or \U$35054 ( \42999_43299 , 1'b0 , \42997_43297 , \42998_43298 );
xor \U$35055 ( \43000_43300 , \42996_43296 , \42999_43299 );
xor \U$35062 ( \43001_43301 , \43000_43300 , 1'b0 );
and \U$35063 ( \43002_43302 , \42980_43280 , \42985_43285 );
and \U$35064 ( \43003_43303 , \42980_43280 , \42991_43291 );
and \U$35065 ( \43004_43304 , \42985_43285 , \42991_43291 );
or \U$35066 ( \43005_43305 , \43002_43302 , \43003_43303 , \43004_43304 );
xor \U$35067 ( \43006_43306 , \43001_43301 , \43005_43305 );
and \U$35068 ( \43007_43307 , \42847_43147 , \42852_43152 );
and \U$35069 ( \43008_43308 , \42847_43147 , \42978_43278 );
and \U$35070 ( \43009_43309 , \42852_43152 , \42978_43278 );
or \U$35071 ( \43010_43310 , \43007_43307 , \43008_43308 , \43009_43309 );
buf \U$35072 ( \43011_43311 , \43010_43310 );
and \U$35073 ( \43012_43312 , \42834_43134 , \42839_43139 );
and \U$35074 ( \43013_43313 , \42834_43134 , \42845_43145 );
and \U$35075 ( \43014_43314 , \42839_43139 , \42845_43145 );
or \U$35076 ( \43015_43315 , \43012_43312 , \43013_43313 , \43014_43314 );
buf \U$35077 ( \43016_43316 , \43015_43315 );
xor \U$35078 ( \43017_43317 , \43011_43311 , \43016_43316 );
and \U$35079 ( \43018_43318 , \42901_43201 , \42906_43206 );
and \U$35080 ( \43019_43319 , \42901_43201 , \42976_43276 );
and \U$35081 ( \43020_43320 , \42906_43206 , \42976_43276 );
or \U$35082 ( \43021_43321 , \43018_43318 , \43019_43319 , \43020_43320 );
buf \U$35083 ( \43022_43322 , \43021_43321 );
and \U$35085 ( \43023_43323 , \32617_32916 , \32881_33181_nG9bae );
or \U$35086 ( \43024_43324 , 1'b0 , \43023_43323 );
xor \U$35087 ( \43025_43325 , 1'b0 , \43024_43324 );
buf \U$35088 ( \43026_43326 , \43025_43325 );
buf \U$35090 ( \43027_43327 , \43026_43326 );
and \U$35091 ( \43028_43328 , \31989_31636 , \33313_33613_nG9bab );
and \U$35092 ( \43029_43329 , \31334_31633 , \33741_34041_nG9ba8 );
or \U$35093 ( \43030_43330 , \43028_43328 , \43029_43329 );
xor \U$35094 ( \43031_43331 , \31333_31632 , \43030_43330 );
buf \U$35095 ( \43032_43332 , \43031_43331 );
buf \U$35097 ( \43033_43333 , \43032_43332 );
xor \U$35098 ( \43034_43334 , \43027_43327 , \43033_43333 );
buf \U$35099 ( \43035_43335 , \43034_43334 );
and \U$35100 ( \43036_43336 , \18908_18702 , \39034_39334_nG9b7b );
and \U$35101 ( \43037_43337 , \18400_18699 , \39291_39591_nG9b78 );
or \U$35102 ( \43038_43338 , \43036_43336 , \43037_43337 );
xor \U$35103 ( \43039_43339 , \18399_18698 , \43038_43338 );
buf \U$35104 ( \43040_43340 , \43039_43339 );
buf \U$35106 ( \43041_43341 , \43040_43340 );
xor \U$35107 ( \43042_43342 , \43035_43335 , \43041_43341 );
and \U$35108 ( \43043_43343 , \13431_13370 , \41385_41685_nG9b63 );
and \U$35109 ( \43044_43344 , \13068_13367 , \41663_41963_nG9b60 );
or \U$35110 ( \43045_43345 , \43043_43343 , \43044_43344 );
xor \U$35111 ( \43046_43346 , \13067_13366 , \43045_43345 );
buf \U$35112 ( \43047_43347 , \43046_43346 );
buf \U$35114 ( \43048_43348 , \43047_43347 );
xor \U$35115 ( \43049_43349 , \43042_43342 , \43048_43348 );
buf \U$35116 ( \43050_43350 , \43049_43349 );
and \U$35117 ( \43051_43351 , \23495_23201 , \36950_37250_nG9b8d );
and \U$35118 ( \43052_43352 , \22899_23198 , \37307_37607_nG9b8a );
or \U$35119 ( \43053_43353 , \43051_43351 , \43052_43352 );
xor \U$35120 ( \43054_43354 , \22898_23197 , \43053_43353 );
buf \U$35121 ( \43055_43355 , \43054_43354 );
buf \U$35123 ( \43056_43356 , \43055_43355 );
and \U$35124 ( \43057_43357 , \21908_21658 , \37674_37974_nG9b87 );
and \U$35125 ( \43058_43358 , \21356_21655 , \38037_38337_nG9b84 );
or \U$35126 ( \43059_43359 , \43057_43357 , \43058_43358 );
xor \U$35127 ( \43060_43360 , \21355_21654 , \43059_43359 );
buf \U$35128 ( \43061_43361 , \43060_43360 );
buf \U$35130 ( \43062_43362 , \43061_43361 );
xor \U$35131 ( \43063_43363 , \43056_43356 , \43062_43362 );
and \U$35132 ( \43064_43364 , \12183_12157 , \41901_42201_nG9b5d );
and \U$35133 ( \43065_43365 , \11855_12154 , \42133_42433_nG9b5a );
or \U$35134 ( \43066_43366 , \43064_43364 , \43065_43365 );
xor \U$35135 ( \43067_43367 , \11854_12153 , \43066_43366 );
buf \U$35136 ( \43068_43368 , \43067_43367 );
buf \U$35138 ( \43069_43369 , \43068_43368 );
xor \U$35139 ( \43070_43370 , \43063_43363 , \43069_43369 );
buf \U$35140 ( \43071_43371 , \43070_43370 );
xor \U$35141 ( \43072_43372 , \43050_43350 , \43071_43371 );
and \U$35142 ( \43073_43373 , \42912_43212 , \42918_43218 );
buf \U$35143 ( \43074_43374 , \43073_43373 );
and \U$35144 ( \43075_43375 , \20353_20155 , \38363_38663_nG9b81 );
and \U$35145 ( \43076_43376 , \19853_20152 , \38668_38968_nG9b7e );
or \U$35146 ( \43077_43377 , \43075_43375 , \43076_43376 );
xor \U$35147 ( \43078_43378 , \19852_20151 , \43077_43377 );
buf \U$35148 ( \43079_43379 , \43078_43378 );
buf \U$35150 ( \43080_43380 , \43079_43379 );
xor \U$35151 ( \43081_43381 , \43074_43374 , \43080_43380 );
and \U$35152 ( \43082_43382 , \14710_14631 , \40740_41040_nG9b69 );
and \U$35153 ( \43083_43383 , \14329_14628 , \41081_41381_nG9b66 );
or \U$35154 ( \43084_43384 , \43082_43382 , \43083_43383 );
xor \U$35155 ( \43085_43385 , \14328_14627 , \43084_43384 );
buf \U$35156 ( \43086_43386 , \43085_43385 );
buf \U$35158 ( \43087_43387 , \43086_43386 );
xor \U$35159 ( \43088_43388 , \43081_43381 , \43087_43387 );
buf \U$35160 ( \43089_43389 , \43088_43388 );
xor \U$35161 ( \43090_43390 , \43072_43372 , \43089_43389 );
buf \U$35162 ( \43091_43391 , \43090_43390 );
and \U$35163 ( \43092_43392 , \42768_43068 , \42773_43073 );
and \U$35164 ( \43093_43393 , \42768_43068 , \42795_43095 );
and \U$35165 ( \43094_43394 , \42773_43073 , \42795_43095 );
or \U$35166 ( \43095_43395 , \43092_43392 , \43093_43393 , \43094_43394 );
buf \U$35167 ( \43096_43396 , \43095_43395 );
and \U$35168 ( \43097_43397 , \42780_43080 , \42786_43086 );
and \U$35169 ( \43098_43398 , \42780_43080 , \42793_43093 );
and \U$35170 ( \43099_43399 , \42786_43086 , \42793_43093 );
or \U$35171 ( \43100_43400 , \43097_43397 , \43098_43398 , \43099_43399 );
buf \U$35172 ( \43101_43401 , \43100_43400 );
and \U$35173 ( \43102_43402 , \10411_10707 , \42879_43179_nG9b51 );
or \U$35176 ( \43103_43403 , \43102_43402 , 1'b0 );
xor \U$35177 ( \43104_43404 , \10399_10703 , \43103_43403 );
buf \U$35178 ( \43105_43405 , \43104_43404 );
buf \U$35180 ( \43106_43406 , \43105_43405 );
xor \U$35181 ( \43107_43407 , \43101_43401 , \43106_43406 );
and \U$35182 ( \43108_43408 , \10996_10421 , \42466_42766_nG9b57 );
and \U$35183 ( \43109_43409 , \10119_10418 , \42548_42848_nG9b54 );
or \U$35184 ( \43110_43410 , \43108_43408 , \43109_43409 );
xor \U$35185 ( \43111_43411 , \10118_10417 , \43110_43410 );
buf \U$35186 ( \43112_43412 , \43111_43411 );
buf \U$35188 ( \43113_43413 , \43112_43412 );
xor \U$35189 ( \43114_43414 , \43107_43407 , \43113_43413 );
buf \U$35190 ( \43115_43415 , \43114_43414 );
xor \U$35191 ( \43116_43416 , \43096_43396 , \43115_43415 );
and \U$35192 ( \43117_43417 , \42863_43163 , \42884_43184 );
and \U$35193 ( \43118_43418 , \42863_43163 , \42891_43191 );
and \U$35194 ( \43119_43419 , \42884_43184 , \42891_43191 );
or \U$35195 ( \43120_43420 , \43117_43417 , \43118_43418 , \43119_43419 );
buf \U$35196 ( \43121_43421 , \43120_43420 );
xor \U$35197 ( \43122_43422 , \43116_43416 , \43121_43421 );
buf \U$35198 ( \43123_43423 , \43122_43422 );
xor \U$35199 ( \43124_43424 , \43091_43391 , \43123_43423 );
and \U$35200 ( \43125_43425 , \42935_43235 , \42956_43256 );
and \U$35201 ( \43126_43426 , \42935_43235 , \42974_43274 );
and \U$35202 ( \43127_43427 , \42956_43256 , \42974_43274 );
or \U$35203 ( \43128_43428 , \43125_43425 , \43126_43426 , \43127_43427 );
buf \U$35204 ( \43129_43429 , \43128_43428 );
xor \U$35205 ( \43130_43430 , \43124_43424 , \43129_43429 );
buf \U$35206 ( \43131_43431 , \43130_43430 );
xor \U$35207 ( \43132_43432 , \43022_43322 , \43131_43431 );
and \U$35208 ( \43133_43433 , \42858_43158 , \42893_43193 );
and \U$35209 ( \43134_43434 , \42858_43158 , \42899_43199 );
and \U$35210 ( \43135_43435 , \42893_43193 , \42899_43199 );
or \U$35211 ( \43136_43436 , \43133_43433 , \43134_43434 , \43135_43435 );
buf \U$35212 ( \43137_43437 , \43136_43436 );
and \U$35213 ( \43138_43438 , \42763_43063 , \42797_43097 );
and \U$35214 ( \43139_43439 , \42763_43063 , \42832_43132 );
and \U$35215 ( \43140_43440 , \42797_43097 , \42832_43132 );
or \U$35216 ( \43141_43441 , \43138_43438 , \43139_43439 , \43140_43440 );
buf \U$35217 ( \43142_43442 , \43141_43441 );
xor \U$35218 ( \43143_43443 , \43137_43437 , \43142_43442 );
and \U$35219 ( \43144_43444 , \42819_43119 , \42824_43124 );
and \U$35220 ( \43145_43445 , \42819_43119 , \42830_43130 );
and \U$35221 ( \43146_43446 , \42824_43124 , \42830_43130 );
or \U$35222 ( \43147_43447 , \43144_43444 , \43145_43445 , \43146_43446 );
buf \U$35223 ( \43148_43448 , \43147_43447 );
and \U$35224 ( \43149_43449 , \42959_43259 , \42965_43265 );
and \U$35225 ( \43150_43450 , \42959_43259 , \42972_43272 );
and \U$35226 ( \43151_43451 , \42965_43265 , \42972_43272 );
or \U$35227 ( \43152_43452 , \43149_43449 , \43150_43450 , \43151_43451 );
buf \U$35228 ( \43153_43453 , \43152_43452 );
and \U$35229 ( \43154_43454 , \30670_29853 , \33994_34294_nG9ba5 );
and \U$35230 ( \43155_43455 , \29551_29850 , \34343_34643_nG9ba2 );
or \U$35231 ( \43156_43456 , \43154_43454 , \43155_43455 );
xor \U$35232 ( \43157_43457 , \29550_29849 , \43156_43456 );
buf \U$35233 ( \43158_43458 , \43157_43457 );
buf \U$35235 ( \43159_43459 , \43158_43458 );
and \U$35236 ( \43160_43460 , \28946_28118 , \34794_35094_nG9b9f );
and \U$35237 ( \43161_43461 , \27816_28115 , \35270_35570_nG9b9c );
or \U$35238 ( \43162_43462 , \43160_43460 , \43161_43461 );
xor \U$35239 ( \43163_43463 , \27815_28114 , \43162_43462 );
buf \U$35240 ( \43164_43464 , \43163_43463 );
buf \U$35242 ( \43165_43465 , \43164_43464 );
xor \U$35243 ( \43166_43466 , \43159_43459 , \43165_43465 );
and \U$35244 ( \43167_43467 , \27141_26431 , \35501_35801_nG9b99 );
and \U$35245 ( \43168_43468 , \26129_26428 , \35872_36172_nG9b96 );
or \U$35246 ( \43169_43469 , \43167_43467 , \43168_43468 );
xor \U$35247 ( \43170_43470 , \26128_26427 , \43169_43469 );
buf \U$35248 ( \43171_43471 , \43170_43470 );
buf \U$35250 ( \43172_43472 , \43171_43471 );
xor \U$35251 ( \43173_43473 , \43166_43466 , \43172_43472 );
buf \U$35252 ( \43174_43474 , \43173_43473 );
xor \U$35253 ( \43175_43475 , \43153_43453 , \43174_43474 );
and \U$35254 ( \43176_43476 , \42920_43220 , \42926_43226 );
and \U$35255 ( \43177_43477 , \42920_43220 , \42933_43233 );
and \U$35256 ( \43178_43478 , \42926_43226 , \42933_43233 );
or \U$35257 ( \43179_43479 , \43176_43476 , \43177_43477 , \43178_43478 );
buf \U$35258 ( \43180_43480 , \43179_43479 );
xor \U$35259 ( \43181_43481 , \43175_43475 , \43180_43480 );
buf \U$35260 ( \43182_43482 , \43181_43481 );
xor \U$35261 ( \43183_43483 , \43148_43448 , \43182_43482 );
and \U$35262 ( \43184_43484 , \42804_43104 , \42810_43110 );
and \U$35263 ( \43185_43485 , \42804_43104 , \42817_43117 );
and \U$35264 ( \43186_43486 , \42810_43110 , \42817_43117 );
or \U$35265 ( \43187_43487 , \43184_43484 , \43185_43485 , \43186_43486 );
buf \U$35266 ( \43188_43488 , \43187_43487 );
and \U$35267 ( \43189_43489 , \25044_24792 , \36289_36589_nG9b93 );
and \U$35268 ( \43190_43490 , \24490_24789 , \36686_36986_nG9b90 );
or \U$35269 ( \43191_43491 , \43189_43489 , \43190_43490 );
xor \U$35270 ( \43192_43492 , \24489_24788 , \43191_43491 );
buf \U$35271 ( \43193_43493 , \43192_43492 );
buf \U$35273 ( \43194_43494 , \43193_43493 );
and \U$35274 ( \43195_43495 , \17437_17297 , \39663_39963_nG9b75 );
and \U$35275 ( \43196_43496 , \16995_17294 , \39904_40204_nG9b72 );
or \U$35276 ( \43197_43497 , \43195_43495 , \43196_43496 );
xor \U$35277 ( \43198_43498 , \16994_17293 , \43197_43497 );
buf \U$35278 ( \43199_43499 , \43198_43498 );
buf \U$35280 ( \43200_43500 , \43199_43499 );
xor \U$35281 ( \43201_43501 , \43194_43494 , \43200_43500 );
and \U$35282 ( \43202_43502 , \16405_15940 , \40152_40452_nG9b6f );
and \U$35283 ( \43203_43503 , \15638_15937 , \40543_40843_nG9b6c );
or \U$35284 ( \43204_43504 , \43202_43502 , \43203_43503 );
xor \U$35285 ( \43205_43505 , \15637_15936 , \43204_43504 );
buf \U$35286 ( \43206_43506 , \43205_43505 );
buf \U$35288 ( \43207_43507 , \43206_43506 );
xor \U$35289 ( \43208_43508 , \43201_43501 , \43207_43507 );
buf \U$35290 ( \43209_43509 , \43208_43508 );
xor \U$35291 ( \43210_43510 , \43188_43488 , \43209_43509 );
and \U$35292 ( \43211_43511 , \42941_43241 , \42947_43247 );
and \U$35293 ( \43212_43512 , \42941_43241 , \42954_43254 );
and \U$35294 ( \43213_43513 , \42947_43247 , \42954_43254 );
or \U$35295 ( \43214_43514 , \43211_43511 , \43212_43512 , \43213_43513 );
buf \U$35296 ( \43215_43515 , \43214_43514 );
xor \U$35297 ( \43216_43516 , \43210_43510 , \43215_43515 );
buf \U$35298 ( \43217_43517 , \43216_43516 );
xor \U$35299 ( \43218_43518 , \43183_43483 , \43217_43517 );
buf \U$35300 ( \43219_43519 , \43218_43518 );
xor \U$35301 ( \43220_43520 , \43143_43443 , \43219_43519 );
buf \U$35302 ( \43221_43521 , \43220_43520 );
xor \U$35303 ( \43222_43522 , \43132_43432 , \43221_43521 );
buf \U$35304 ( \43223_43523 , \43222_43522 );
xor \U$35305 ( \43224_43524 , \43017_43317 , \43223_43523 );
and \U$35306 ( \43225_43525 , \43006_43306 , \43224_43524 );
and \U$35308 ( \43226_43526 , \43000_43300 , \43005_43305 );
or \U$35310 ( \43227_43527 , 1'b0 , \43226_43526 , 1'b0 );
xor \U$35311 ( \43228_43528 , \43225_43525 , \43227_43527 );
and \U$35313 ( \43229_43529 , \42993_43293 , \42999_43299 );
and \U$35314 ( \43230_43530 , \42995_43295 , \42999_43299 );
or \U$35315 ( \43231_43531 , 1'b0 , \43229_43529 , \43230_43530 );
xor \U$35316 ( \43232_43532 , \43228_43528 , \43231_43531 );
xor \U$35323 ( \43233_43533 , \43232_43532 , 1'b0 );
and \U$35324 ( \43234_43534 , \43011_43311 , \43016_43316 );
and \U$35325 ( \43235_43535 , \43011_43311 , \43223_43523 );
and \U$35326 ( \43236_43536 , \43016_43316 , \43223_43523 );
or \U$35327 ( \43237_43537 , \43234_43534 , \43235_43535 , \43236_43536 );
xor \U$35328 ( \43238_43538 , \43233_43533 , \43237_43537 );
and \U$35329 ( \43239_43539 , \43022_43322 , \43131_43431 );
and \U$35330 ( \43240_43540 , \43022_43322 , \43221_43521 );
and \U$35331 ( \43241_43541 , \43131_43431 , \43221_43521 );
or \U$35332 ( \43242_43542 , \43239_43539 , \43240_43540 , \43241_43541 );
buf \U$35333 ( \43243_43543 , \43242_43542 );
and \U$35334 ( \43244_43544 , \43137_43437 , \43142_43442 );
and \U$35335 ( \43245_43545 , \43137_43437 , \43219_43519 );
and \U$35336 ( \43246_43546 , \43142_43442 , \43219_43519 );
or \U$35337 ( \43247_43547 , \43244_43544 , \43245_43545 , \43246_43546 );
buf \U$35338 ( \43248_43548 , \43247_43547 );
and \U$35339 ( \43249_43549 , \43050_43350 , \43071_43371 );
and \U$35340 ( \43250_43550 , \43050_43350 , \43089_43389 );
and \U$35341 ( \43251_43551 , \43071_43371 , \43089_43389 );
or \U$35342 ( \43252_43552 , \43249_43549 , \43250_43550 , \43251_43551 );
buf \U$35343 ( \43253_43553 , \43252_43552 );
and \U$35344 ( \43254_43554 , \43153_43453 , \43174_43474 );
and \U$35345 ( \43255_43555 , \43153_43453 , \43180_43480 );
and \U$35346 ( \43256_43556 , \43174_43474 , \43180_43480 );
or \U$35347 ( \43257_43557 , \43254_43554 , \43255_43555 , \43256_43556 );
buf \U$35348 ( \43258_43558 , \43257_43557 );
and \U$35349 ( \43259_43559 , \43159_43459 , \43165_43465 );
and \U$35350 ( \43260_43560 , \43159_43459 , \43172_43472 );
and \U$35351 ( \43261_43561 , \43165_43465 , \43172_43472 );
or \U$35352 ( \43262_43562 , \43259_43559 , \43260_43560 , \43261_43561 );
buf \U$35353 ( \43263_43563 , \43262_43562 );
xor \U$35358 ( \43264_43564 , \10399_10703 , 1'b0 );
not \U$35359 ( \43265_43565 , \43264_43564 );
buf \U$35360 ( \43266_43566 , \43265_43565 );
buf \U$35362 ( \43267_43567 , \43266_43566 );
xor \U$35363 ( \43268_43568 , 1'b1 , \43267_43567 );
and \U$35365 ( \43269_43569 , \32617_32916 , \33313_33613_nG9bab );
or \U$35366 ( \43270_43570 , 1'b0 , \43269_43569 );
xor \U$35367 ( \43271_43571 , 1'b0 , \43270_43570 );
buf \U$35368 ( \43272_43572 , \43271_43571 );
buf \U$35370 ( \43273_43573 , \43272_43572 );
xor \U$35371 ( \43274_43574 , \43268_43568 , \43273_43573 );
buf \U$35372 ( \43275_43575 , \43274_43574 );
xor \U$35373 ( \43276_43576 , \43263_43563 , \43275_43575 );
and \U$35374 ( \43277_43577 , \12183_12157 , \42133_42433_nG9b5a );
and \U$35375 ( \43278_43578 , \11855_12154 , \42466_42766_nG9b57 );
or \U$35376 ( \43279_43579 , \43277_43577 , \43278_43578 );
xor \U$35377 ( \43280_43580 , \11854_12153 , \43279_43579 );
buf \U$35378 ( \43281_43581 , \43280_43580 );
buf \U$35380 ( \43282_43582 , \43281_43581 );
xor \U$35381 ( \43283_43583 , \43276_43576 , \43282_43582 );
buf \U$35382 ( \43284_43584 , \43283_43583 );
xor \U$35383 ( \43285_43585 , \43258_43558 , \43284_43584 );
and \U$35384 ( \43286_43586 , \43101_43401 , \43106_43406 );
and \U$35385 ( \43287_43587 , \43101_43401 , \43113_43413 );
and \U$35386 ( \43288_43588 , \43106_43406 , \43113_43413 );
or \U$35387 ( \43289_43589 , \43286_43586 , \43287_43587 , \43288_43588 );
buf \U$35388 ( \43290_43590 , \43289_43589 );
xor \U$35389 ( \43291_43591 , \43285_43585 , \43290_43590 );
buf \U$35390 ( \43292_43592 , \43291_43591 );
xor \U$35391 ( \43293_43593 , \43253_43553 , \43292_43592 );
and \U$35392 ( \43294_43594 , \43027_43327 , \43033_43333 );
buf \U$35393 ( \43295_43595 , \43294_43594 );
and \U$35394 ( \43296_43596 , \20353_20155 , \38668_38968_nG9b7e );
and \U$35395 ( \43297_43597 , \19853_20152 , \39034_39334_nG9b7b );
or \U$35396 ( \43298_43598 , \43296_43596 , \43297_43597 );
xor \U$35397 ( \43299_43599 , \19852_20151 , \43298_43598 );
buf \U$35398 ( \43300_43600 , \43299_43599 );
buf \U$35400 ( \43301_43601 , \43300_43600 );
xor \U$35401 ( \43302_43602 , \43295_43595 , \43301_43601 );
and \U$35402 ( \43303_43603 , \14710_14631 , \41081_41381_nG9b66 );
and \U$35403 ( \43304_43604 , \14329_14628 , \41385_41685_nG9b63 );
or \U$35404 ( \43305_43605 , \43303_43603 , \43304_43604 );
xor \U$35405 ( \43306_43606 , \14328_14627 , \43305_43605 );
buf \U$35406 ( \43307_43607 , \43306_43606 );
buf \U$35408 ( \43308_43608 , \43307_43607 );
xor \U$35409 ( \43309_43609 , \43302_43602 , \43308_43608 );
buf \U$35410 ( \43310_43610 , \43309_43609 );
and \U$35411 ( \43311_43611 , \10996_10421 , \42548_42848_nG9b54 );
and \U$35412 ( \43312_43612 , \10119_10418 , \42879_43179_nG9b51 );
or \U$35413 ( \43313_43613 , \43311_43611 , \43312_43612 );
xor \U$35414 ( \43314_43614 , \10118_10417 , \43313_43613 );
buf \U$35415 ( \43315_43615 , \43314_43614 );
buf \U$35417 ( \43316_43616 , \43315_43615 );
and \U$35418 ( \43317_43617 , \18908_18702 , \39291_39591_nG9b78 );
and \U$35419 ( \43318_43618 , \18400_18699 , \39663_39963_nG9b75 );
or \U$35420 ( \43319_43619 , \43317_43617 , \43318_43618 );
xor \U$35421 ( \43320_43620 , \18399_18698 , \43319_43619 );
buf \U$35422 ( \43321_43621 , \43320_43620 );
buf \U$35424 ( \43322_43622 , \43321_43621 );
xor \U$35425 ( \43323_43623 , \43316_43616 , \43322_43622 );
and \U$35426 ( \43324_43624 , \13431_13370 , \41663_41963_nG9b60 );
and \U$35427 ( \43325_43625 , \13068_13367 , \41901_42201_nG9b5d );
or \U$35428 ( \43326_43626 , \43324_43624 , \43325_43625 );
xor \U$35429 ( \43327_43627 , \13067_13366 , \43326_43626 );
buf \U$35430 ( \43328_43628 , \43327_43627 );
buf \U$35432 ( \43329_43629 , \43328_43628 );
xor \U$35433 ( \43330_43630 , \43323_43623 , \43329_43629 );
buf \U$35434 ( \43331_43631 , \43330_43630 );
xor \U$35435 ( \43332_43632 , \43310_43610 , \43331_43631 );
and \U$35436 ( \43333_43633 , \25044_24792 , \36686_36986_nG9b90 );
and \U$35437 ( \43334_43634 , \24490_24789 , \36950_37250_nG9b8d );
or \U$35438 ( \43335_43635 , \43333_43633 , \43334_43634 );
xor \U$35439 ( \43336_43636 , \24489_24788 , \43335_43635 );
buf \U$35440 ( \43337_43637 , \43336_43636 );
buf \U$35442 ( \43338_43638 , \43337_43637 );
and \U$35443 ( \43339_43639 , \23495_23201 , \37307_37607_nG9b8a );
and \U$35444 ( \43340_43640 , \22899_23198 , \37674_37974_nG9b87 );
or \U$35445 ( \43341_43641 , \43339_43639 , \43340_43640 );
xor \U$35446 ( \43342_43642 , \22898_23197 , \43341_43641 );
buf \U$35447 ( \43343_43643 , \43342_43642 );
buf \U$35449 ( \43344_43644 , \43343_43643 );
xor \U$35450 ( \43345_43645 , \43338_43638 , \43344_43644 );
and \U$35451 ( \43346_43646 , \21908_21658 , \38037_38337_nG9b84 );
and \U$35452 ( \43347_43647 , \21356_21655 , \38363_38663_nG9b81 );
or \U$35453 ( \43348_43648 , \43346_43646 , \43347_43647 );
xor \U$35454 ( \43349_43649 , \21355_21654 , \43348_43648 );
buf \U$35455 ( \43350_43650 , \43349_43649 );
buf \U$35457 ( \43351_43651 , \43350_43650 );
xor \U$35458 ( \43352_43652 , \43345_43645 , \43351_43651 );
buf \U$35459 ( \43353_43653 , \43352_43652 );
xor \U$35460 ( \43354_43654 , \43332_43632 , \43353_43653 );
buf \U$35461 ( \43355_43655 , \43354_43654 );
xor \U$35462 ( \43356_43656 , \43293_43593 , \43355_43655 );
buf \U$35463 ( \43357_43657 , \43356_43656 );
xor \U$35464 ( \43358_43658 , \43248_43548 , \43357_43657 );
and \U$35465 ( \43359_43659 , \43091_43391 , \43123_43423 );
and \U$35466 ( \43360_43660 , \43091_43391 , \43129_43429 );
and \U$35467 ( \43361_43661 , \43123_43423 , \43129_43429 );
or \U$35468 ( \43362_43662 , \43359_43659 , \43360_43660 , \43361_43661 );
buf \U$35469 ( \43363_43663 , \43362_43662 );
xor \U$35470 ( \43364_43664 , \43358_43658 , \43363_43663 );
buf \U$35471 ( \43365_43665 , \43364_43664 );
xor \U$35472 ( \43366_43666 , \43243_43543 , \43365_43665 );
and \U$35473 ( \43367_43667 , \43148_43448 , \43182_43482 );
and \U$35474 ( \43368_43668 , \43148_43448 , \43217_43517 );
and \U$35475 ( \43369_43669 , \43182_43482 , \43217_43517 );
or \U$35476 ( \43370_43670 , \43367_43667 , \43368_43668 , \43369_43669 );
buf \U$35477 ( \43371_43671 , \43370_43670 );
and \U$35478 ( \43372_43672 , \43096_43396 , \43115_43415 );
and \U$35479 ( \43373_43673 , \43096_43396 , \43121_43421 );
and \U$35480 ( \43374_43674 , \43115_43415 , \43121_43421 );
or \U$35481 ( \43375_43675 , \43372_43672 , \43373_43673 , \43374_43674 );
buf \U$35482 ( \43376_43676 , \43375_43675 );
xor \U$35483 ( \43377_43677 , \43371_43671 , \43376_43676 );
and \U$35484 ( \43378_43678 , \43188_43488 , \43209_43509 );
and \U$35485 ( \43379_43679 , \43188_43488 , \43215_43515 );
and \U$35486 ( \43380_43680 , \43209_43509 , \43215_43515 );
or \U$35487 ( \43381_43681 , \43378_43678 , \43379_43679 , \43380_43680 );
buf \U$35488 ( \43382_43682 , \43381_43681 );
and \U$35489 ( \43383_43683 , \27141_26431 , \35872_36172_nG9b96 );
and \U$35490 ( \43384_43684 , \26129_26428 , \36289_36589_nG9b93 );
or \U$35491 ( \43385_43685 , \43383_43683 , \43384_43684 );
xor \U$35492 ( \43386_43686 , \26128_26427 , \43385_43685 );
buf \U$35493 ( \43387_43687 , \43386_43686 );
buf \U$35495 ( \43388_43688 , \43387_43687 );
and \U$35496 ( \43389_43689 , \17437_17297 , \39904_40204_nG9b72 );
and \U$35497 ( \43390_43690 , \16995_17294 , \40152_40452_nG9b6f );
or \U$35498 ( \43391_43691 , \43389_43689 , \43390_43690 );
xor \U$35499 ( \43392_43692 , \16994_17293 , \43391_43691 );
buf \U$35500 ( \43393_43693 , \43392_43692 );
buf \U$35502 ( \43394_43694 , \43393_43693 );
xor \U$35503 ( \43395_43695 , \43388_43688 , \43394_43694 );
and \U$35504 ( \43396_43696 , \16405_15940 , \40543_40843_nG9b6c );
and \U$35505 ( \43397_43697 , \15638_15937 , \40740_41040_nG9b69 );
or \U$35506 ( \43398_43698 , \43396_43696 , \43397_43697 );
xor \U$35507 ( \43399_43699 , \15637_15936 , \43398_43698 );
buf \U$35508 ( \43400_43700 , \43399_43699 );
buf \U$35510 ( \43401_43701 , \43400_43700 );
xor \U$35511 ( \43402_43702 , \43395_43695 , \43401_43701 );
buf \U$35512 ( \43403_43703 , \43402_43702 );
and \U$35513 ( \43404_43704 , \43194_43494 , \43200_43500 );
and \U$35514 ( \43405_43705 , \43194_43494 , \43207_43507 );
and \U$35515 ( \43406_43706 , \43200_43500 , \43207_43507 );
or \U$35516 ( \43407_43707 , \43404_43704 , \43405_43705 , \43406_43706 );
buf \U$35517 ( \43408_43708 , \43407_43707 );
xor \U$35518 ( \43409_43709 , \43403_43703 , \43408_43708 );
and \U$35519 ( \43410_43710 , \43056_43356 , \43062_43362 );
and \U$35520 ( \43411_43711 , \43056_43356 , \43069_43369 );
and \U$35521 ( \43412_43712 , \43062_43362 , \43069_43369 );
or \U$35522 ( \43413_43713 , \43410_43710 , \43411_43711 , \43412_43712 );
buf \U$35523 ( \43414_43714 , \43413_43713 );
xor \U$35524 ( \43415_43715 , \43409_43709 , \43414_43714 );
buf \U$35525 ( \43416_43716 , \43415_43715 );
xor \U$35526 ( \43417_43717 , \43382_43682 , \43416_43716 );
and \U$35527 ( \43418_43718 , \43035_43335 , \43041_43341 );
and \U$35528 ( \43419_43719 , \43035_43335 , \43048_43348 );
and \U$35529 ( \43420_43720 , \43041_43341 , \43048_43348 );
or \U$35530 ( \43421_43721 , \43418_43718 , \43419_43719 , \43420_43720 );
buf \U$35531 ( \43422_43722 , \43421_43721 );
and \U$35532 ( \43423_43723 , \31989_31636 , \33741_34041_nG9ba8 );
and \U$35533 ( \43424_43724 , \31334_31633 , \33994_34294_nG9ba5 );
or \U$35534 ( \43425_43725 , \43423_43723 , \43424_43724 );
xor \U$35535 ( \43426_43726 , \31333_31632 , \43425_43725 );
buf \U$35536 ( \43427_43727 , \43426_43726 );
buf \U$35538 ( \43428_43728 , \43427_43727 );
and \U$35539 ( \43429_43729 , \30670_29853 , \34343_34643_nG9ba2 );
and \U$35540 ( \43430_43730 , \29551_29850 , \34794_35094_nG9b9f );
or \U$35541 ( \43431_43731 , \43429_43729 , \43430_43730 );
xor \U$35542 ( \43432_43732 , \29550_29849 , \43431_43731 );
buf \U$35543 ( \43433_43733 , \43432_43732 );
buf \U$35545 ( \43434_43734 , \43433_43733 );
xor \U$35546 ( \43435_43735 , \43428_43728 , \43434_43734 );
and \U$35547 ( \43436_43736 , \28946_28118 , \35270_35570_nG9b9c );
and \U$35548 ( \43437_43737 , \27816_28115 , \35501_35801_nG9b99 );
or \U$35549 ( \43438_43738 , \43436_43736 , \43437_43737 );
xor \U$35550 ( \43439_43739 , \27815_28114 , \43438_43738 );
buf \U$35551 ( \43440_43740 , \43439_43739 );
buf \U$35553 ( \43441_43741 , \43440_43740 );
xor \U$35554 ( \43442_43742 , \43435_43735 , \43441_43741 );
buf \U$35555 ( \43443_43743 , \43442_43742 );
xor \U$35556 ( \43444_43744 , \43422_43722 , \43443_43743 );
and \U$35557 ( \43445_43745 , \43074_43374 , \43080_43380 );
and \U$35558 ( \43446_43746 , \43074_43374 , \43087_43387 );
and \U$35559 ( \43447_43747 , \43080_43380 , \43087_43387 );
or \U$35560 ( \43448_43748 , \43445_43745 , \43446_43746 , \43447_43747 );
buf \U$35561 ( \43449_43749 , \43448_43748 );
xor \U$35562 ( \43450_43750 , \43444_43744 , \43449_43749 );
buf \U$35563 ( \43451_43751 , \43450_43750 );
xor \U$35564 ( \43452_43752 , \43417_43717 , \43451_43751 );
buf \U$35565 ( \43453_43753 , \43452_43752 );
xor \U$35566 ( \43454_43754 , \43377_43677 , \43453_43753 );
buf \U$35567 ( \43455_43755 , \43454_43754 );
xor \U$35568 ( \43456_43756 , \43366_43666 , \43455_43755 );
and \U$35569 ( \43457_43757 , \43238_43538 , \43456_43756 );
and \U$35571 ( \43458_43758 , \43232_43532 , \43237_43537 );
or \U$35573 ( \43459_43759 , 1'b0 , \43458_43758 , 1'b0 );
xor \U$35574 ( \43460_43760 , \43457_43757 , \43459_43759 );
and \U$35576 ( \43461_43761 , \43225_43525 , \43231_43531 );
and \U$35577 ( \43462_43762 , \43227_43527 , \43231_43531 );
or \U$35578 ( \43463_43763 , 1'b0 , \43461_43761 , \43462_43762 );
xor \U$35579 ( \43464_43764 , \43460_43760 , \43463_43763 );
xor \U$35586 ( \43465_43765 , \43464_43764 , 1'b0 );
and \U$35587 ( \43466_43766 , \43243_43543 , \43365_43665 );
and \U$35588 ( \43467_43767 , \43243_43543 , \43455_43755 );
and \U$35589 ( \43468_43768 , \43365_43665 , \43455_43755 );
or \U$35590 ( \43469_43769 , \43466_43766 , \43467_43767 , \43468_43768 );
xor \U$35591 ( \43470_43770 , \43465_43765 , \43469_43769 );
and \U$35592 ( \43471_43771 , \43371_43671 , \43376_43676 );
and \U$35593 ( \43472_43772 , \43371_43671 , \43453_43753 );
and \U$35594 ( \43473_43773 , \43376_43676 , \43453_43753 );
or \U$35595 ( \43474_43774 , \43471_43771 , \43472_43772 , \43473_43773 );
buf \U$35596 ( \43475_43775 , \43474_43774 );
and \U$35597 ( \43476_43776 , \43253_43553 , \43292_43592 );
and \U$35598 ( \43477_43777 , \43253_43553 , \43355_43655 );
and \U$35599 ( \43478_43778 , \43292_43592 , \43355_43655 );
or \U$35600 ( \43479_43779 , \43476_43776 , \43477_43777 , \43478_43778 );
buf \U$35601 ( \43480_43780 , \43479_43779 );
xor \U$35602 ( \43481_43781 , \43475_43775 , \43480_43780 );
and \U$35603 ( \43482_43782 , \43403_43703 , \43408_43708 );
and \U$35604 ( \43483_43783 , \43403_43703 , \43414_43714 );
and \U$35605 ( \43484_43784 , \43408_43708 , \43414_43714 );
or \U$35606 ( \43485_43785 , \43482_43782 , \43483_43783 , \43484_43784 );
buf \U$35607 ( \43486_43786 , \43485_43785 );
and \U$35608 ( \43487_43787 , \43422_43722 , \43443_43743 );
and \U$35609 ( \43488_43788 , \43422_43722 , \43449_43749 );
and \U$35610 ( \43489_43789 , \43443_43743 , \43449_43749 );
or \U$35611 ( \43490_43790 , \43487_43787 , \43488_43788 , \43489_43789 );
buf \U$35612 ( \43491_43791 , \43490_43790 );
and \U$35613 ( \43492_43792 , \43428_43728 , \43434_43734 );
and \U$35614 ( \43493_43793 , \43428_43728 , \43441_43741 );
and \U$35615 ( \43494_43794 , \43434_43734 , \43441_43741 );
or \U$35616 ( \43495_43795 , \43492_43792 , \43493_43793 , \43494_43794 );
buf \U$35617 ( \43496_43796 , \43495_43795 );
and \U$35618 ( \43497_43797 , 1'b1 , \43267_43567 );
and \U$35619 ( \43498_43798 , 1'b1 , \43273_43573 );
and \U$35620 ( \43499_43799 , \43267_43567 , \43273_43573 );
or \U$35621 ( \43500_43800 , \43497_43797 , \43498_43798 , \43499_43799 );
buf \U$35622 ( \43501_43801 , \43500_43800 );
xor \U$35623 ( \43502_43802 , \43496_43796 , \43501_43801 );
and \U$35624 ( \43503_43803 , \12183_12157 , \42466_42766_nG9b57 );
and \U$35625 ( \43504_43804 , \11855_12154 , \42548_42848_nG9b54 );
or \U$35626 ( \43505_43805 , \43503_43803 , \43504_43804 );
xor \U$35627 ( \43506_43806 , \11854_12153 , \43505_43805 );
buf \U$35628 ( \43507_43807 , \43506_43806 );
buf \U$35630 ( \43508_43808 , \43507_43807 );
xor \U$35631 ( \43509_43809 , \43502_43802 , \43508_43808 );
buf \U$35632 ( \43510_43810 , \43509_43809 );
xor \U$35633 ( \43511_43811 , \43491_43791 , \43510_43810 );
and \U$35634 ( \43512_43812 , \43263_43563 , \43275_43575 );
and \U$35635 ( \43513_43813 , \43263_43563 , \43282_43582 );
and \U$35636 ( \43514_43814 , \43275_43575 , \43282_43582 );
or \U$35637 ( \43515_43815 , \43512_43812 , \43513_43813 , \43514_43814 );
buf \U$35638 ( \43516_43816 , \43515_43815 );
xor \U$35639 ( \43517_43817 , \43511_43811 , \43516_43816 );
buf \U$35640 ( \43518_43818 , \43517_43817 );
xor \U$35641 ( \43519_43819 , \43486_43786 , \43518_43818 );
and \U$35642 ( \43520_43820 , \23495_23201 , \37674_37974_nG9b87 );
and \U$35643 ( \43521_43821 , \22899_23198 , \38037_38337_nG9b84 );
or \U$35644 ( \43522_43822 , \43520_43820 , \43521_43821 );
xor \U$35645 ( \43523_43823 , \22898_23197 , \43522_43822 );
buf \U$35646 ( \43524_43824 , \43523_43823 );
buf \U$35648 ( \43525_43825 , \43524_43824 );
and \U$35649 ( \43526_43826 , \21908_21658 , \38363_38663_nG9b81 );
and \U$35650 ( \43527_43827 , \21356_21655 , \38668_38968_nG9b7e );
or \U$35651 ( \43528_43828 , \43526_43826 , \43527_43827 );
xor \U$35652 ( \43529_43829 , \21355_21654 , \43528_43828 );
buf \U$35653 ( \43530_43830 , \43529_43829 );
buf \U$35655 ( \43531_43831 , \43530_43830 );
xor \U$35656 ( \43532_43832 , \43525_43825 , \43531_43831 );
and \U$35657 ( \43533_43833 , \16405_15940 , \40740_41040_nG9b69 );
and \U$35658 ( \43534_43834 , \15638_15937 , \41081_41381_nG9b66 );
or \U$35659 ( \43535_43835 , \43533_43833 , \43534_43834 );
xor \U$35660 ( \43536_43836 , \15637_15936 , \43535_43835 );
buf \U$35661 ( \43537_43837 , \43536_43836 );
buf \U$35663 ( \43538_43838 , \43537_43837 );
xor \U$35664 ( \43539_43839 , \43532_43832 , \43538_43838 );
buf \U$35665 ( \43540_43840 , \43539_43839 );
and \U$35666 ( \43541_43841 , \27141_26431 , \36289_36589_nG9b93 );
and \U$35667 ( \43542_43842 , \26129_26428 , \36686_36986_nG9b90 );
or \U$35668 ( \43543_43843 , \43541_43841 , \43542_43842 );
xor \U$35669 ( \43544_43844 , \26128_26427 , \43543_43843 );
buf \U$35670 ( \43545_43845 , \43544_43844 );
buf \U$35672 ( \43546_43846 , \43545_43845 );
and \U$35673 ( \43547_43847 , \25044_24792 , \36950_37250_nG9b8d );
and \U$35674 ( \43548_43848 , \24490_24789 , \37307_37607_nG9b8a );
or \U$35675 ( \43549_43849 , \43547_43847 , \43548_43848 );
xor \U$35676 ( \43550_43850 , \24489_24788 , \43549_43849 );
buf \U$35677 ( \43551_43851 , \43550_43850 );
buf \U$35679 ( \43552_43852 , \43551_43851 );
xor \U$35680 ( \43553_43853 , \43546_43846 , \43552_43852 );
and \U$35681 ( \43554_43854 , \13431_13370 , \41901_42201_nG9b5d );
and \U$35682 ( \43555_43855 , \13068_13367 , \42133_42433_nG9b5a );
or \U$35683 ( \43556_43856 , \43554_43854 , \43555_43855 );
xor \U$35684 ( \43557_43857 , \13067_13366 , \43556_43856 );
buf \U$35685 ( \43558_43858 , \43557_43857 );
buf \U$35687 ( \43559_43859 , \43558_43858 );
xor \U$35688 ( \43560_43860 , \43553_43853 , \43559_43859 );
buf \U$35689 ( \43561_43861 , \43560_43860 );
xor \U$35690 ( \43562_43862 , \43540_43840 , \43561_43861 );
and \U$35692 ( \43563_43863 , \32617_32916 , \33741_34041_nG9ba8 );
or \U$35693 ( \43564_43864 , 1'b0 , \43563_43863 );
xor \U$35694 ( \43565_43865 , 1'b0 , \43564_43864 );
buf \U$35695 ( \43566_43866 , \43565_43865 );
buf \U$35696 ( \43567_43867 , \43566_43866 );
not \U$35697 ( \43568_43868 , \43567_43867 );
and \U$35698 ( \43569_43869 , \20353_20155 , \39034_39334_nG9b7b );
and \U$35699 ( \43570_43870 , \19853_20152 , \39291_39591_nG9b78 );
or \U$35700 ( \43571_43871 , \43569_43869 , \43570_43870 );
xor \U$35701 ( \43572_43872 , \19852_20151 , \43571_43871 );
buf \U$35702 ( \43573_43873 , \43572_43872 );
buf \U$35704 ( \43574_43874 , \43573_43873 );
xor \U$35705 ( \43575_43875 , \43568_43868 , \43574_43874 );
and \U$35706 ( \43576_43876 , \14710_14631 , \41385_41685_nG9b63 );
and \U$35707 ( \43577_43877 , \14329_14628 , \41663_41963_nG9b60 );
or \U$35708 ( \43578_43878 , \43576_43876 , \43577_43877 );
xor \U$35709 ( \43579_43879 , \14328_14627 , \43578_43878 );
buf \U$35710 ( \43580_43880 , \43579_43879 );
buf \U$35712 ( \43581_43881 , \43580_43880 );
xor \U$35713 ( \43582_43882 , \43575_43875 , \43581_43881 );
buf \U$35714 ( \43583_43883 , \43582_43882 );
xor \U$35715 ( \43584_43884 , \43562_43862 , \43583_43883 );
buf \U$35716 ( \43585_43885 , \43584_43884 );
xor \U$35717 ( \43586_43886 , \43519_43819 , \43585_43885 );
buf \U$35718 ( \43587_43887 , \43586_43886 );
xor \U$35719 ( \43588_43888 , \43481_43781 , \43587_43887 );
buf \U$35720 ( \43589_43889 , \43588_43888 );
and \U$35721 ( \43590_43890 , \43248_43548 , \43357_43657 );
and \U$35722 ( \43591_43891 , \43248_43548 , \43363_43663 );
and \U$35723 ( \43592_43892 , \43357_43657 , \43363_43663 );
or \U$35724 ( \43593_43893 , \43590_43890 , \43591_43891 , \43592_43892 );
buf \U$35725 ( \43594_43894 , \43593_43893 );
xor \U$35726 ( \43595_43895 , \43589_43889 , \43594_43894 );
and \U$35727 ( \43596_43896 , \43310_43610 , \43331_43631 );
and \U$35728 ( \43597_43897 , \43310_43610 , \43353_43653 );
and \U$35729 ( \43598_43898 , \43331_43631 , \43353_43653 );
or \U$35730 ( \43599_43899 , \43596_43896 , \43597_43897 , \43598_43898 );
buf \U$35731 ( \43600_43900 , \43599_43899 );
and \U$35732 ( \43601_43901 , \10996_10421 , \42879_43179_nG9b51 );
or \U$35734 ( \43602_43902 , \43601_43901 , 1'b0 );
xor \U$35735 ( \43603_43903 , \10118_10417 , \43602_43902 );
buf \U$35736 ( \43604_43904 , \43603_43903 );
buf \U$35738 ( \43605_43905 , \43604_43904 );
and \U$35739 ( \43606_43906 , \18908_18702 , \39663_39963_nG9b75 );
and \U$35740 ( \43607_43907 , \18400_18699 , \39904_40204_nG9b72 );
or \U$35741 ( \43608_43908 , \43606_43906 , \43607_43907 );
xor \U$35742 ( \43609_43909 , \18399_18698 , \43608_43908 );
buf \U$35743 ( \43610_43910 , \43609_43909 );
buf \U$35745 ( \43611_43911 , \43610_43910 );
xor \U$35746 ( \43612_43912 , \43605_43905 , \43611_43911 );
and \U$35747 ( \43613_43913 , \17437_17297 , \40152_40452_nG9b6f );
and \U$35748 ( \43614_43914 , \16995_17294 , \40543_40843_nG9b6c );
or \U$35749 ( \43615_43915 , \43613_43913 , \43614_43914 );
xor \U$35750 ( \43616_43916 , \16994_17293 , \43615_43915 );
buf \U$35751 ( \43617_43917 , \43616_43916 );
buf \U$35753 ( \43618_43918 , \43617_43917 );
xor \U$35754 ( \43619_43919 , \43612_43912 , \43618_43918 );
buf \U$35755 ( \43620_43920 , \43619_43919 );
and \U$35756 ( \43621_43921 , \43388_43688 , \43394_43694 );
and \U$35757 ( \43622_43922 , \43388_43688 , \43401_43701 );
and \U$35758 ( \43623_43923 , \43394_43694 , \43401_43701 );
or \U$35759 ( \43624_43924 , \43621_43921 , \43622_43922 , \43623_43923 );
buf \U$35760 ( \43625_43925 , \43624_43924 );
xor \U$35761 ( \43626_43926 , \43620_43920 , \43625_43925 );
and \U$35762 ( \43627_43927 , \43338_43638 , \43344_43644 );
and \U$35763 ( \43628_43928 , \43338_43638 , \43351_43651 );
and \U$35764 ( \43629_43929 , \43344_43644 , \43351_43651 );
or \U$35765 ( \43630_43930 , \43627_43927 , \43628_43928 , \43629_43929 );
buf \U$35766 ( \43631_43931 , \43630_43930 );
xor \U$35767 ( \43632_43932 , \43626_43926 , \43631_43931 );
buf \U$35768 ( \43633_43933 , \43632_43932 );
xor \U$35769 ( \43634_43934 , \43600_43900 , \43633_43933 );
and \U$35770 ( \43635_43935 , \43295_43595 , \43301_43601 );
and \U$35771 ( \43636_43936 , \43295_43595 , \43308_43608 );
and \U$35772 ( \43637_43937 , \43301_43601 , \43308_43608 );
or \U$35773 ( \43638_43938 , \43635_43935 , \43636_43936 , \43637_43937 );
buf \U$35774 ( \43639_43939 , \43638_43938 );
and \U$35775 ( \43640_43940 , \31989_31636 , \33994_34294_nG9ba5 );
and \U$35776 ( \43641_43941 , \31334_31633 , \34343_34643_nG9ba2 );
or \U$35777 ( \43642_43942 , \43640_43940 , \43641_43941 );
xor \U$35778 ( \43643_43943 , \31333_31632 , \43642_43942 );
buf \U$35779 ( \43644_43944 , \43643_43943 );
buf \U$35781 ( \43645_43945 , \43644_43944 );
and \U$35782 ( \43646_43946 , \30670_29853 , \34794_35094_nG9b9f );
and \U$35783 ( \43647_43947 , \29551_29850 , \35270_35570_nG9b9c );
or \U$35784 ( \43648_43948 , \43646_43946 , \43647_43947 );
xor \U$35785 ( \43649_43949 , \29550_29849 , \43648_43948 );
buf \U$35786 ( \43650_43950 , \43649_43949 );
buf \U$35788 ( \43651_43951 , \43650_43950 );
xor \U$35789 ( \43652_43952 , \43645_43945 , \43651_43951 );
and \U$35790 ( \43653_43953 , \28946_28118 , \35501_35801_nG9b99 );
and \U$35791 ( \43654_43954 , \27816_28115 , \35872_36172_nG9b96 );
or \U$35792 ( \43655_43955 , \43653_43953 , \43654_43954 );
xor \U$35793 ( \43656_43956 , \27815_28114 , \43655_43955 );
buf \U$35794 ( \43657_43957 , \43656_43956 );
buf \U$35796 ( \43658_43958 , \43657_43957 );
xor \U$35797 ( \43659_43959 , \43652_43952 , \43658_43958 );
buf \U$35798 ( \43660_43960 , \43659_43959 );
xor \U$35799 ( \43661_43961 , \43639_43939 , \43660_43960 );
and \U$35800 ( \43662_43962 , \43316_43616 , \43322_43622 );
and \U$35801 ( \43663_43963 , \43316_43616 , \43329_43629 );
and \U$35802 ( \43664_43964 , \43322_43622 , \43329_43629 );
or \U$35803 ( \43665_43965 , \43662_43962 , \43663_43963 , \43664_43964 );
buf \U$35804 ( \43666_43966 , \43665_43965 );
xor \U$35805 ( \43667_43967 , \43661_43961 , \43666_43966 );
buf \U$35806 ( \43668_43968 , \43667_43967 );
xor \U$35807 ( \43669_43969 , \43634_43934 , \43668_43968 );
buf \U$35808 ( \43670_43970 , \43669_43969 );
and \U$35809 ( \43671_43971 , \43258_43558 , \43284_43584 );
and \U$35810 ( \43672_43972 , \43258_43558 , \43290_43590 );
and \U$35811 ( \43673_43973 , \43284_43584 , \43290_43590 );
or \U$35812 ( \43674_43974 , \43671_43971 , \43672_43972 , \43673_43973 );
buf \U$35813 ( \43675_43975 , \43674_43974 );
xor \U$35814 ( \43676_43976 , \43670_43970 , \43675_43975 );
and \U$35815 ( \43677_43977 , \43382_43682 , \43416_43716 );
and \U$35816 ( \43678_43978 , \43382_43682 , \43451_43751 );
and \U$35817 ( \43679_43979 , \43416_43716 , \43451_43751 );
or \U$35818 ( \43680_43980 , \43677_43977 , \43678_43978 , \43679_43979 );
buf \U$35819 ( \43681_43981 , \43680_43980 );
xor \U$35820 ( \43682_43982 , \43676_43976 , \43681_43981 );
buf \U$35821 ( \43683_43983 , \43682_43982 );
xor \U$35822 ( \43684_43984 , \43595_43895 , \43683_43983 );
and \U$35823 ( \43685_43985 , \43470_43770 , \43684_43984 );
and \U$35825 ( \43686_43986 , \43464_43764 , \43469_43769 );
or \U$35827 ( \43687_43987 , 1'b0 , \43686_43986 , 1'b0 );
xor \U$35828 ( \43688_43988 , \43685_43985 , \43687_43987 );
and \U$35830 ( \43689_43989 , \43457_43757 , \43463_43763 );
and \U$35831 ( \43690_43990 , \43459_43759 , \43463_43763 );
or \U$35832 ( \43691_43991 , 1'b0 , \43689_43989 , \43690_43990 );
xor \U$35833 ( \43692_43992 , \43688_43988 , \43691_43991 );
xor \U$35840 ( \43693_43993 , \43692_43992 , 1'b0 );
and \U$35841 ( \43694_43994 , \43589_43889 , \43594_43894 );
and \U$35842 ( \43695_43995 , \43589_43889 , \43683_43983 );
and \U$35843 ( \43696_43996 , \43594_43894 , \43683_43983 );
or \U$35844 ( \43697_43997 , \43694_43994 , \43695_43995 , \43696_43996 );
xor \U$35845 ( \43698_43998 , \43693_43993 , \43697_43997 );
and \U$35846 ( \43699_43999 , \43475_43775 , \43480_43780 );
and \U$35847 ( \43700_44000 , \43475_43775 , \43587_43887 );
and \U$35848 ( \43701_44001 , \43480_43780 , \43587_43887 );
or \U$35849 ( \43702_44002 , \43699_43999 , \43700_44000 , \43701_44001 );
buf \U$35850 ( \43703_44003 , \43702_44002 );
and \U$35851 ( \43704_44004 , \43639_43939 , \43660_43960 );
and \U$35852 ( \43705_44005 , \43639_43939 , \43666_43966 );
and \U$35853 ( \43706_44006 , \43660_43960 , \43666_43966 );
or \U$35854 ( \43707_44007 , \43704_44004 , \43705_44005 , \43706_44006 );
buf \U$35855 ( \43708_44008 , \43707_44007 );
and \U$35856 ( \43709_44009 , \43496_43796 , \43501_43801 );
and \U$35857 ( \43710_44010 , \43496_43796 , \43508_43808 );
and \U$35858 ( \43711_44011 , \43501_43801 , \43508_43808 );
or \U$35859 ( \43712_44012 , \43709_44009 , \43710_44010 , \43711_44011 );
buf \U$35860 ( \43713_44013 , \43712_44012 );
xor \U$35861 ( \43714_44014 , \43708_44008 , \43713_44013 );
and \U$35862 ( \43715_44015 , \43645_43945 , \43651_43951 );
and \U$35863 ( \43716_44016 , \43645_43945 , \43658_43958 );
and \U$35864 ( \43717_44017 , \43651_43951 , \43658_43958 );
or \U$35865 ( \43718_44018 , \43715_44015 , \43716_44016 , \43717_44017 );
buf \U$35866 ( \43719_44019 , \43718_44018 );
and \U$35867 ( \43720_44020 , \17437_17297 , \40543_40843_nG9b6c );
and \U$35868 ( \43721_44021 , \16995_17294 , \40740_41040_nG9b69 );
or \U$35869 ( \43722_44022 , \43720_44020 , \43721_44021 );
xor \U$35870 ( \43723_44023 , \16994_17293 , \43722_44022 );
buf \U$35871 ( \43724_44024 , \43723_44023 );
buf \U$35873 ( \43725_44025 , \43724_44024 );
xor \U$35874 ( \43726_44026 , \43719_44019 , \43725_44025 );
and \U$35875 ( \43727_44027 , \13431_13370 , \42133_42433_nG9b5a );
and \U$35876 ( \43728_44028 , \13068_13367 , \42466_42766_nG9b57 );
or \U$35877 ( \43729_44029 , \43727_44027 , \43728_44028 );
xor \U$35878 ( \43730_44030 , \13067_13366 , \43729_44029 );
buf \U$35879 ( \43731_44031 , \43730_44030 );
buf \U$35881 ( \43732_44032 , \43731_44031 );
xor \U$35882 ( \43733_44033 , \43726_44026 , \43732_44032 );
buf \U$35883 ( \43734_44034 , \43733_44033 );
xor \U$35884 ( \43735_44035 , \43714_44014 , \43734_44034 );
buf \U$35885 ( \43736_44036 , \43735_44035 );
and \U$35886 ( \43737_44037 , \43540_43840 , \43561_43861 );
and \U$35887 ( \43738_44038 , \43540_43840 , \43583_43883 );
and \U$35888 ( \43739_44039 , \43561_43861 , \43583_43883 );
or \U$35889 ( \43740_44040 , \43737_44037 , \43738_44038 , \43739_44039 );
buf \U$35890 ( \43741_44041 , \43740_44040 );
and \U$35891 ( \43742_44042 , \28946_28118 , \35872_36172_nG9b96 );
and \U$35892 ( \43743_44043 , \27816_28115 , \36289_36589_nG9b93 );
or \U$35893 ( \43744_44044 , \43742_44042 , \43743_44043 );
xor \U$35894 ( \43745_44045 , \27815_28114 , \43744_44044 );
buf \U$35895 ( \43746_44046 , \43745_44045 );
buf \U$35897 ( \43747_44047 , \43746_44046 );
and \U$35898 ( \43748_44048 , \27141_26431 , \36686_36986_nG9b90 );
and \U$35899 ( \43749_44049 , \26129_26428 , \36950_37250_nG9b8d );
or \U$35900 ( \43750_44050 , \43748_44048 , \43749_44049 );
xor \U$35901 ( \43751_44051 , \26128_26427 , \43750_44050 );
buf \U$35902 ( \43752_44052 , \43751_44051 );
buf \U$35904 ( \43753_44053 , \43752_44052 );
xor \U$35905 ( \43754_44054 , \43747_44047 , \43753_44053 );
and \U$35906 ( \43755_44055 , \18908_18702 , \39904_40204_nG9b72 );
and \U$35907 ( \43756_44056 , \18400_18699 , \40152_40452_nG9b6f );
or \U$35908 ( \43757_44057 , \43755_44055 , \43756_44056 );
xor \U$35909 ( \43758_44058 , \18399_18698 , \43757_44057 );
buf \U$35910 ( \43759_44059 , \43758_44058 );
buf \U$35912 ( \43760_44060 , \43759_44059 );
xor \U$35913 ( \43761_44061 , \43754_44054 , \43760_44060 );
buf \U$35914 ( \43762_44062 , \43761_44061 );
and \U$35915 ( \43763_44063 , \43605_43905 , \43611_43911 );
and \U$35916 ( \43764_44064 , \43605_43905 , \43618_43918 );
and \U$35917 ( \43765_44065 , \43611_43911 , \43618_43918 );
or \U$35918 ( \43766_44066 , \43763_44063 , \43764_44064 , \43765_44065 );
buf \U$35919 ( \43767_44067 , \43766_44066 );
xor \U$35920 ( \43768_44068 , \43762_44062 , \43767_44067 );
and \U$35921 ( \43769_44069 , \43546_43846 , \43552_43852 );
and \U$35922 ( \43770_44070 , \43546_43846 , \43559_43859 );
and \U$35923 ( \43771_44071 , \43552_43852 , \43559_43859 );
or \U$35924 ( \43772_44072 , \43769_44069 , \43770_44070 , \43771_44071 );
buf \U$35925 ( \43773_44073 , \43772_44072 );
xor \U$35926 ( \43774_44074 , \43768_44068 , \43773_44073 );
buf \U$35927 ( \43775_44075 , \43774_44074 );
xor \U$35928 ( \43776_44076 , \43741_44041 , \43775_44075 );
and \U$35929 ( \43777_44077 , \43620_43920 , \43625_43925 );
and \U$35930 ( \43778_44078 , \43620_43920 , \43631_43931 );
and \U$35931 ( \43779_44079 , \43625_43925 , \43631_43931 );
or \U$35932 ( \43780_44080 , \43777_44077 , \43778_44078 , \43779_44079 );
buf \U$35933 ( \43781_44081 , \43780_44080 );
xor \U$35934 ( \43782_44082 , \43776_44076 , \43781_44081 );
buf \U$35935 ( \43783_44083 , \43782_44082 );
xor \U$35936 ( \43784_44084 , \43736_44036 , \43783_44083 );
and \U$35937 ( \43785_44085 , \43600_43900 , \43633_43933 );
and \U$35938 ( \43786_44086 , \43600_43900 , \43668_43968 );
and \U$35939 ( \43787_44087 , \43633_43933 , \43668_43968 );
or \U$35940 ( \43788_44088 , \43785_44085 , \43786_44086 , \43787_44087 );
buf \U$35941 ( \43789_44089 , \43788_44088 );
xor \U$35942 ( \43790_44090 , \43784_44084 , \43789_44089 );
buf \U$35943 ( \43791_44091 , \43790_44090 );
xor \U$35944 ( \43792_44092 , \43703_44003 , \43791_44091 );
and \U$35945 ( \43793_44093 , \43670_43970 , \43675_43975 );
and \U$35946 ( \43794_44094 , \43670_43970 , \43681_43981 );
and \U$35947 ( \43795_44095 , \43675_43975 , \43681_43981 );
or \U$35948 ( \43796_44096 , \43793_44093 , \43794_44094 , \43795_44095 );
buf \U$35949 ( \43797_44097 , \43796_44096 );
and \U$35950 ( \43798_44098 , \43491_43791 , \43510_43810 );
and \U$35951 ( \43799_44099 , \43491_43791 , \43516_43816 );
and \U$35952 ( \43800_44100 , \43510_43810 , \43516_43816 );
or \U$35953 ( \43801_44101 , \43798_44098 , \43799_44099 , \43800_44100 );
buf \U$35954 ( \43802_44102 , \43801_44101 );
buf \U$35955 ( \43803_44103 , \43567_43867 );
and \U$35956 ( \43804_44104 , \21908_21658 , \38668_38968_nG9b7e );
and \U$35957 ( \43805_44105 , \21356_21655 , \39034_39334_nG9b7b );
or \U$35958 ( \43806_44106 , \43804_44104 , \43805_44105 );
xor \U$35959 ( \43807_44107 , \21355_21654 , \43806_44106 );
buf \U$35960 ( \43808_44108 , \43807_44107 );
buf \U$35962 ( \43809_44109 , \43808_44108 );
xor \U$35963 ( \43810_44110 , \43803_44103 , \43809_44109 );
and \U$35964 ( \43811_44111 , \20353_20155 , \39291_39591_nG9b78 );
and \U$35965 ( \43812_44112 , \19853_20152 , \39663_39963_nG9b75 );
or \U$35966 ( \43813_44113 , \43811_44111 , \43812_44112 );
xor \U$35967 ( \43814_44114 , \19852_20151 , \43813_44113 );
buf \U$35968 ( \43815_44115 , \43814_44114 );
buf \U$35970 ( \43816_44116 , \43815_44115 );
xor \U$35971 ( \43817_44117 , \43810_44110 , \43816_44116 );
buf \U$35972 ( \43818_44118 , \43817_44117 );
and \U$35973 ( \43819_44119 , \12183_12157 , \42548_42848_nG9b54 );
and \U$35974 ( \43820_44120 , \11855_12154 , \42879_43179_nG9b51 );
or \U$35975 ( \43821_44121 , \43819_44119 , \43820_44120 );
xor \U$35976 ( \43822_44122 , \11854_12153 , \43821_44121 );
buf \U$35977 ( \43823_44123 , \43822_44122 );
buf \U$35979 ( \43824_44124 , \43823_44123 );
and \U$35980 ( \43825_44125 , \31989_31636 , \34343_34643_nG9ba2 );
and \U$35981 ( \43826_44126 , \31334_31633 , \34794_35094_nG9b9f );
or \U$35982 ( \43827_44127 , \43825_44125 , \43826_44126 );
xor \U$35983 ( \43828_44128 , \31333_31632 , \43827_44127 );
buf \U$35984 ( \43829_44129 , \43828_44128 );
buf \U$35986 ( \43830_44130 , \43829_44129 );
xor \U$35987 ( \43831_44131 , \43824_44124 , \43830_44130 );
and \U$35988 ( \43832_44132 , \14710_14631 , \41663_41963_nG9b60 );
and \U$35989 ( \43833_44133 , \14329_14628 , \41901_42201_nG9b5d );
or \U$35990 ( \43834_44134 , \43832_44132 , \43833_44133 );
xor \U$35991 ( \43835_44135 , \14328_14627 , \43834_44134 );
buf \U$35992 ( \43836_44136 , \43835_44135 );
buf \U$35994 ( \43837_44137 , \43836_44136 );
xor \U$35995 ( \43838_44138 , \43831_44131 , \43837_44137 );
buf \U$35996 ( \43839_44139 , \43838_44138 );
xor \U$35997 ( \43840_44140 , \43818_44118 , \43839_44139 );
and \U$35998 ( \43841_44141 , \25044_24792 , \37307_37607_nG9b8a );
and \U$35999 ( \43842_44142 , \24490_24789 , \37674_37974_nG9b87 );
or \U$36000 ( \43843_44143 , \43841_44141 , \43842_44142 );
xor \U$36001 ( \43844_44144 , \24489_24788 , \43843_44143 );
buf \U$36002 ( \43845_44145 , \43844_44144 );
buf \U$36004 ( \43846_44146 , \43845_44145 );
and \U$36005 ( \43847_44147 , \23495_23201 , \38037_38337_nG9b84 );
and \U$36006 ( \43848_44148 , \22899_23198 , \38363_38663_nG9b81 );
or \U$36007 ( \43849_44149 , \43847_44147 , \43848_44148 );
xor \U$36008 ( \43850_44150 , \22898_23197 , \43849_44149 );
buf \U$36009 ( \43851_44151 , \43850_44150 );
buf \U$36011 ( \43852_44152 , \43851_44151 );
xor \U$36012 ( \43853_44153 , \43846_44146 , \43852_44152 );
and \U$36013 ( \43854_44154 , \16405_15940 , \41081_41381_nG9b66 );
and \U$36014 ( \43855_44155 , \15638_15937 , \41385_41685_nG9b63 );
or \U$36015 ( \43856_44156 , \43854_44154 , \43855_44155 );
xor \U$36016 ( \43857_44157 , \15637_15936 , \43856_44156 );
buf \U$36017 ( \43858_44158 , \43857_44157 );
buf \U$36019 ( \43859_44159 , \43858_44158 );
xor \U$36020 ( \43860_44160 , \43853_44153 , \43859_44159 );
buf \U$36021 ( \43861_44161 , \43860_44160 );
xor \U$36022 ( \43862_44162 , \43840_44140 , \43861_44161 );
buf \U$36023 ( \43863_44163 , \43862_44162 );
xor \U$36024 ( \43864_44164 , \43802_44102 , \43863_44163 );
and \U$36025 ( \43865_44165 , \43525_43825 , \43531_43831 );
and \U$36026 ( \43866_44166 , \43525_43825 , \43538_43838 );
and \U$36027 ( \43867_44167 , \43531_43831 , \43538_43838 );
or \U$36028 ( \43868_44168 , \43865_44165 , \43866_44166 , \43867_44167 );
buf \U$36029 ( \43869_44169 , \43868_44168 );
and \U$36030 ( \43870_44170 , \43568_43868 , \43574_43874 );
and \U$36031 ( \43871_44171 , \43568_43868 , \43581_43881 );
and \U$36032 ( \43872_44172 , \43574_43874 , \43581_43881 );
or \U$36033 ( \43873_44173 , \43870_44170 , \43871_44171 , \43872_44172 );
buf \U$36034 ( \43874_44174 , \43873_44173 );
xor \U$36035 ( \43875_44175 , \43869_44169 , \43874_44174 );
xor \U$36039 ( \43876_44176 , \10118_10417 , 1'b0 );
not \U$36040 ( \43877_44177 , \43876_44176 );
buf \U$36041 ( \43878_44178 , \43877_44177 );
buf \U$36043 ( \43879_44179 , \43878_44178 );
and \U$36045 ( \43880_44180 , \32617_32916 , \33994_34294_nG9ba5 );
or \U$36046 ( \43881_44181 , 1'b0 , \43880_44180 );
xor \U$36047 ( \43882_44182 , 1'b0 , \43881_44181 );
buf \U$36048 ( \43883_44183 , \43882_44182 );
buf \U$36050 ( \43884_44184 , \43883_44183 );
xor \U$36051 ( \43885_44185 , \43879_44179 , \43884_44184 );
and \U$36052 ( \43886_44186 , \30670_29853 , \35270_35570_nG9b9c );
and \U$36053 ( \43887_44187 , \29551_29850 , \35501_35801_nG9b99 );
or \U$36054 ( \43888_44188 , \43886_44186 , \43887_44187 );
xor \U$36055 ( \43889_44189 , \29550_29849 , \43888_44188 );
buf \U$36056 ( \43890_44190 , \43889_44189 );
buf \U$36058 ( \43891_44191 , \43890_44190 );
xor \U$36059 ( \43892_44192 , \43885_44185 , \43891_44191 );
buf \U$36060 ( \43893_44193 , \43892_44192 );
xor \U$36061 ( \43894_44194 , \43875_44175 , \43893_44193 );
buf \U$36062 ( \43895_44195 , \43894_44194 );
xor \U$36063 ( \43896_44196 , \43864_44164 , \43895_44195 );
buf \U$36064 ( \43897_44197 , \43896_44196 );
xor \U$36065 ( \43898_44198 , \43797_44097 , \43897_44197 );
and \U$36066 ( \43899_44199 , \43486_43786 , \43518_43818 );
and \U$36067 ( \43900_44200 , \43486_43786 , \43585_43885 );
and \U$36068 ( \43901_44201 , \43518_43818 , \43585_43885 );
or \U$36069 ( \43902_44202 , \43899_44199 , \43900_44200 , \43901_44201 );
buf \U$36070 ( \43903_44203 , \43902_44202 );
xor \U$36071 ( \43904_44204 , \43898_44198 , \43903_44203 );
buf \U$36072 ( \43905_44205 , \43904_44204 );
xor \U$36073 ( \43906_44206 , \43792_44092 , \43905_44205 );
and \U$36074 ( \43907_44207 , \43698_43998 , \43906_44206 );
and \U$36076 ( \43908_44208 , \43692_43992 , \43697_43997 );
or \U$36078 ( \43909_44209 , 1'b0 , \43908_44208 , 1'b0 );
xor \U$36079 ( \43910_44210 , \43907_44207 , \43909_44209 );
and \U$36081 ( \43911_44211 , \43685_43985 , \43691_43991 );
and \U$36082 ( \43912_44212 , \43687_43987 , \43691_43991 );
or \U$36083 ( \43913_44213 , 1'b0 , \43911_44211 , \43912_44212 );
xor \U$36084 ( \43914_44214 , \43910_44210 , \43913_44213 );
xor \U$36091 ( \43915_44215 , \43914_44214 , 1'b0 );
and \U$36092 ( \43916_44216 , \43703_44003 , \43791_44091 );
and \U$36093 ( \43917_44217 , \43703_44003 , \43905_44205 );
and \U$36094 ( \43918_44218 , \43791_44091 , \43905_44205 );
or \U$36095 ( \43919_44219 , \43916_44216 , \43917_44217 , \43918_44218 );
xor \U$36096 ( \43920_44220 , \43915_44215 , \43919_44219 );
and \U$36097 ( \43921_44221 , \43797_44097 , \43897_44197 );
and \U$36098 ( \43922_44222 , \43797_44097 , \43903_44203 );
and \U$36099 ( \43923_44223 , \43897_44197 , \43903_44203 );
or \U$36100 ( \43924_44224 , \43921_44221 , \43922_44222 , \43923_44223 );
buf \U$36101 ( \43925_44225 , \43924_44224 );
and \U$36102 ( \43926_44226 , \43741_44041 , \43775_44075 );
and \U$36103 ( \43927_44227 , \43741_44041 , \43781_44081 );
and \U$36104 ( \43928_44228 , \43775_44075 , \43781_44081 );
or \U$36105 ( \43929_44229 , \43926_44226 , \43927_44227 , \43928_44228 );
buf \U$36106 ( \43930_44230 , \43929_44229 );
and \U$36107 ( \43931_44231 , \43818_44118 , \43839_44139 );
and \U$36108 ( \43932_44232 , \43818_44118 , \43861_44161 );
and \U$36109 ( \43933_44233 , \43839_44139 , \43861_44161 );
or \U$36110 ( \43934_44234 , \43931_44231 , \43932_44232 , \43933_44233 );
buf \U$36111 ( \43935_44235 , \43934_44234 );
and \U$36113 ( \43936_44236 , \32617_32916 , \34343_34643_nG9ba2 );
or \U$36114 ( \43937_44237 , 1'b0 , \43936_44236 );
xor \U$36115 ( \43938_44238 , 1'b0 , \43937_44237 );
buf \U$36116 ( \43939_44239 , \43938_44238 );
buf \U$36118 ( \43940_44240 , \43939_44239 );
and \U$36119 ( \43941_44241 , \31989_31636 , \34794_35094_nG9b9f );
and \U$36120 ( \43942_44242 , \31334_31633 , \35270_35570_nG9b9c );
or \U$36121 ( \43943_44243 , \43941_44241 , \43942_44242 );
xor \U$36122 ( \43944_44244 , \31333_31632 , \43943_44243 );
buf \U$36123 ( \43945_44245 , \43944_44244 );
buf \U$36125 ( \43946_44246 , \43945_44245 );
xor \U$36126 ( \43947_44247 , \43940_44240 , \43946_44246 );
and \U$36127 ( \43948_44248 , \16405_15940 , \41385_41685_nG9b63 );
and \U$36128 ( \43949_44249 , \15638_15937 , \41663_41963_nG9b60 );
or \U$36129 ( \43950_44250 , \43948_44248 , \43949_44249 );
xor \U$36130 ( \43951_44251 , \15637_15936 , \43950_44250 );
buf \U$36131 ( \43952_44252 , \43951_44251 );
buf \U$36133 ( \43953_44253 , \43952_44252 );
xor \U$36134 ( \43954_44254 , \43947_44247 , \43953_44253 );
buf \U$36135 ( \43955_44255 , \43954_44254 );
and \U$36136 ( \43956_44256 , \43846_44146 , \43852_44152 );
and \U$36137 ( \43957_44257 , \43846_44146 , \43859_44159 );
and \U$36138 ( \43958_44258 , \43852_44152 , \43859_44159 );
or \U$36139 ( \43959_44259 , \43956_44256 , \43957_44257 , \43958_44258 );
buf \U$36140 ( \43960_44260 , \43959_44259 );
xor \U$36141 ( \43961_44261 , \43955_44255 , \43960_44260 );
and \U$36142 ( \43962_44262 , \43747_44047 , \43753_44053 );
and \U$36143 ( \43963_44263 , \43747_44047 , \43760_44060 );
and \U$36144 ( \43964_44264 , \43753_44053 , \43760_44060 );
or \U$36145 ( \43965_44265 , \43962_44262 , \43963_44263 , \43964_44264 );
buf \U$36146 ( \43966_44266 , \43965_44265 );
xor \U$36147 ( \43967_44267 , \43961_44261 , \43966_44266 );
buf \U$36148 ( \43968_44268 , \43967_44267 );
xor \U$36149 ( \43969_44269 , \43935_44235 , \43968_44268 );
and \U$36150 ( \43970_44270 , \43824_44124 , \43830_44130 );
and \U$36151 ( \43971_44271 , \43824_44124 , \43837_44137 );
and \U$36152 ( \43972_44272 , \43830_44130 , \43837_44137 );
or \U$36153 ( \43973_44273 , \43970_44270 , \43971_44271 , \43972_44272 );
buf \U$36154 ( \43974_44274 , \43973_44273 );
and \U$36155 ( \43975_44275 , \43879_44179 , \43884_44184 );
and \U$36156 ( \43976_44276 , \43879_44179 , \43891_44191 );
and \U$36157 ( \43977_44277 , \43884_44184 , \43891_44191 );
or \U$36158 ( \43978_44278 , \43975_44275 , \43976_44276 , \43977_44277 );
buf \U$36159 ( \43979_44279 , \43978_44278 );
xor \U$36160 ( \43980_44280 , \43974_44274 , \43979_44279 );
and \U$36161 ( \43981_44281 , \43803_44103 , \43809_44109 );
and \U$36162 ( \43982_44282 , \43803_44103 , \43816_44116 );
and \U$36163 ( \43983_44283 , \43809_44109 , \43816_44116 );
or \U$36164 ( \43984_44284 , \43981_44281 , \43982_44282 , \43983_44283 );
buf \U$36165 ( \43985_44285 , \43984_44284 );
xor \U$36166 ( \43986_44286 , \43980_44280 , \43985_44285 );
buf \U$36167 ( \43987_44287 , \43986_44286 );
xor \U$36168 ( \43988_44288 , \43969_44269 , \43987_44287 );
buf \U$36169 ( \43989_44289 , \43988_44288 );
xor \U$36170 ( \43990_44290 , \43930_44230 , \43989_44289 );
and \U$36171 ( \43991_44291 , \12183_12157 , \42879_43179_nG9b51 );
or \U$36173 ( \43992_44292 , \43991_44291 , 1'b0 );
xor \U$36174 ( \43993_44293 , \11854_12153 , \43992_44292 );
buf \U$36175 ( \43994_44294 , \43993_44293 );
buf \U$36177 ( \43995_44295 , \43994_44294 );
and \U$36178 ( \43996_44296 , \30670_29853 , \35501_35801_nG9b99 );
and \U$36179 ( \43997_44297 , \29551_29850 , \35872_36172_nG9b96 );
or \U$36180 ( \43998_44298 , \43996_44296 , \43997_44297 );
xor \U$36181 ( \43999_44299 , \29550_29849 , \43998_44298 );
buf \U$36182 ( \44000_44300 , \43999_44299 );
buf \U$36183 ( \44001_44301 , \44000_44300 );
not \U$36184 ( \44002_44302 , \44001_44301 );
xor \U$36185 ( \44003_44303 , \43995_44295 , \44002_44302 );
and \U$36186 ( \44004_44304 , \13431_13370 , \42466_42766_nG9b57 );
and \U$36187 ( \44005_44305 , \13068_13367 , \42548_42848_nG9b54 );
or \U$36188 ( \44006_44306 , \44004_44304 , \44005_44305 );
xor \U$36189 ( \44007_44307 , \13067_13366 , \44006_44306 );
buf \U$36190 ( \44008_44308 , \44007_44307 );
buf \U$36192 ( \44009_44309 , \44008_44308 );
xor \U$36193 ( \44010_44310 , \44003_44303 , \44009_44309 );
buf \U$36194 ( \44011_44311 , \44010_44310 );
and \U$36195 ( \44012_44312 , \43719_44019 , \43725_44025 );
and \U$36196 ( \44013_44313 , \43719_44019 , \43732_44032 );
and \U$36197 ( \44014_44314 , \43725_44025 , \43732_44032 );
or \U$36198 ( \44015_44315 , \44012_44312 , \44013_44313 , \44014_44314 );
buf \U$36199 ( \44016_44316 , \44015_44315 );
xor \U$36200 ( \44017_44317 , \44011_44311 , \44016_44316 );
and \U$36201 ( \44018_44318 , \43869_44169 , \43874_44174 );
and \U$36202 ( \44019_44319 , \43869_44169 , \43893_44193 );
and \U$36203 ( \44020_44320 , \43874_44174 , \43893_44193 );
or \U$36204 ( \44021_44321 , \44018_44318 , \44019_44319 , \44020_44320 );
buf \U$36205 ( \44022_44322 , \44021_44321 );
xor \U$36206 ( \44023_44323 , \44017_44317 , \44022_44322 );
buf \U$36207 ( \44024_44324 , \44023_44323 );
xor \U$36208 ( \44025_44325 , \43990_44290 , \44024_44324 );
buf \U$36209 ( \44026_44326 , \44025_44325 );
and \U$36210 ( \44027_44327 , \43802_44102 , \43863_44163 );
and \U$36211 ( \44028_44328 , \43802_44102 , \43895_44195 );
and \U$36212 ( \44029_44329 , \43863_44163 , \43895_44195 );
or \U$36213 ( \44030_44330 , \44027_44327 , \44028_44328 , \44029_44329 );
buf \U$36214 ( \44031_44331 , \44030_44330 );
xor \U$36215 ( \44032_44332 , \44026_44326 , \44031_44331 );
and \U$36216 ( \44033_44333 , \43708_44008 , \43713_44013 );
and \U$36217 ( \44034_44334 , \43708_44008 , \43734_44034 );
and \U$36218 ( \44035_44335 , \43713_44013 , \43734_44034 );
or \U$36219 ( \44036_44336 , \44033_44333 , \44034_44334 , \44035_44335 );
buf \U$36220 ( \44037_44337 , \44036_44336 );
and \U$36221 ( \44038_44338 , \28946_28118 , \36289_36589_nG9b93 );
and \U$36222 ( \44039_44339 , \27816_28115 , \36686_36986_nG9b90 );
or \U$36223 ( \44040_44340 , \44038_44338 , \44039_44339 );
xor \U$36224 ( \44041_44341 , \27815_28114 , \44040_44340 );
buf \U$36225 ( \44042_44342 , \44041_44341 );
buf \U$36227 ( \44043_44343 , \44042_44342 );
and \U$36228 ( \44044_44344 , \20353_20155 , \39663_39963_nG9b75 );
and \U$36229 ( \44045_44345 , \19853_20152 , \39904_40204_nG9b72 );
or \U$36230 ( \44046_44346 , \44044_44344 , \44045_44345 );
xor \U$36231 ( \44047_44347 , \19852_20151 , \44046_44346 );
buf \U$36232 ( \44048_44348 , \44047_44347 );
buf \U$36234 ( \44049_44349 , \44048_44348 );
xor \U$36235 ( \44050_44350 , \44043_44343 , \44049_44349 );
and \U$36236 ( \44051_44351 , \18908_18702 , \40152_40452_nG9b6f );
and \U$36237 ( \44052_44352 , \18400_18699 , \40543_40843_nG9b6c );
or \U$36238 ( \44053_44353 , \44051_44351 , \44052_44352 );
xor \U$36239 ( \44054_44354 , \18399_18698 , \44053_44353 );
buf \U$36240 ( \44055_44355 , \44054_44354 );
buf \U$36242 ( \44056_44356 , \44055_44355 );
xor \U$36243 ( \44057_44357 , \44050_44350 , \44056_44356 );
buf \U$36244 ( \44058_44358 , \44057_44357 );
and \U$36245 ( \44059_44359 , \23495_23201 , \38363_38663_nG9b81 );
and \U$36246 ( \44060_44360 , \22899_23198 , \38668_38968_nG9b7e );
or \U$36247 ( \44061_44361 , \44059_44359 , \44060_44360 );
xor \U$36248 ( \44062_44362 , \22898_23197 , \44061_44361 );
buf \U$36249 ( \44063_44363 , \44062_44362 );
buf \U$36251 ( \44064_44364 , \44063_44363 );
and \U$36252 ( \44065_44365 , \21908_21658 , \39034_39334_nG9b7b );
and \U$36253 ( \44066_44366 , \21356_21655 , \39291_39591_nG9b78 );
or \U$36254 ( \44067_44367 , \44065_44365 , \44066_44366 );
xor \U$36255 ( \44068_44368 , \21355_21654 , \44067_44367 );
buf \U$36256 ( \44069_44369 , \44068_44368 );
buf \U$36258 ( \44070_44370 , \44069_44369 );
xor \U$36259 ( \44071_44371 , \44064_44364 , \44070_44370 );
and \U$36260 ( \44072_44372 , \17437_17297 , \40740_41040_nG9b69 );
and \U$36261 ( \44073_44373 , \16995_17294 , \41081_41381_nG9b66 );
or \U$36262 ( \44074_44374 , \44072_44372 , \44073_44373 );
xor \U$36263 ( \44075_44375 , \16994_17293 , \44074_44374 );
buf \U$36264 ( \44076_44376 , \44075_44375 );
buf \U$36266 ( \44077_44377 , \44076_44376 );
xor \U$36267 ( \44078_44378 , \44071_44371 , \44077_44377 );
buf \U$36268 ( \44079_44379 , \44078_44378 );
xor \U$36269 ( \44080_44380 , \44058_44358 , \44079_44379 );
and \U$36270 ( \44081_44381 , \27141_26431 , \36950_37250_nG9b8d );
and \U$36271 ( \44082_44382 , \26129_26428 , \37307_37607_nG9b8a );
or \U$36272 ( \44083_44383 , \44081_44381 , \44082_44382 );
xor \U$36273 ( \44084_44384 , \26128_26427 , \44083_44383 );
buf \U$36274 ( \44085_44385 , \44084_44384 );
buf \U$36276 ( \44086_44386 , \44085_44385 );
and \U$36277 ( \44087_44387 , \25044_24792 , \37674_37974_nG9b87 );
and \U$36278 ( \44088_44388 , \24490_24789 , \38037_38337_nG9b84 );
or \U$36279 ( \44089_44389 , \44087_44387 , \44088_44388 );
xor \U$36280 ( \44090_44390 , \24489_24788 , \44089_44389 );
buf \U$36281 ( \44091_44391 , \44090_44390 );
buf \U$36283 ( \44092_44392 , \44091_44391 );
xor \U$36284 ( \44093_44393 , \44086_44386 , \44092_44392 );
and \U$36285 ( \44094_44394 , \14710_14631 , \41901_42201_nG9b5d );
and \U$36286 ( \44095_44395 , \14329_14628 , \42133_42433_nG9b5a );
or \U$36287 ( \44096_44396 , \44094_44394 , \44095_44395 );
xor \U$36288 ( \44097_44397 , \14328_14627 , \44096_44396 );
buf \U$36289 ( \44098_44398 , \44097_44397 );
buf \U$36291 ( \44099_44399 , \44098_44398 );
xor \U$36292 ( \44100_44400 , \44093_44393 , \44099_44399 );
buf \U$36293 ( \44101_44401 , \44100_44400 );
xor \U$36294 ( \44102_44402 , \44080_44380 , \44101_44401 );
buf \U$36295 ( \44103_44403 , \44102_44402 );
xor \U$36296 ( \44104_44404 , \44037_44337 , \44103_44403 );
and \U$36297 ( \44105_44405 , \43762_44062 , \43767_44067 );
and \U$36298 ( \44106_44406 , \43762_44062 , \43773_44073 );
and \U$36299 ( \44107_44407 , \43767_44067 , \43773_44073 );
or \U$36300 ( \44108_44408 , \44105_44405 , \44106_44406 , \44107_44407 );
buf \U$36301 ( \44109_44409 , \44108_44408 );
xor \U$36302 ( \44110_44410 , \44104_44404 , \44109_44409 );
buf \U$36303 ( \44111_44411 , \44110_44410 );
xor \U$36304 ( \44112_44412 , \44032_44332 , \44111_44411 );
buf \U$36305 ( \44113_44413 , \44112_44412 );
xor \U$36306 ( \44114_44414 , \43925_44225 , \44113_44413 );
and \U$36307 ( \44115_44415 , \43736_44036 , \43783_44083 );
and \U$36308 ( \44116_44416 , \43736_44036 , \43789_44089 );
and \U$36309 ( \44117_44417 , \43783_44083 , \43789_44089 );
or \U$36310 ( \44118_44418 , \44115_44415 , \44116_44416 , \44117_44417 );
buf \U$36311 ( \44119_44419 , \44118_44418 );
xor \U$36312 ( \44120_44420 , \44114_44414 , \44119_44419 );
and \U$36313 ( \44121_44421 , \43920_44220 , \44120_44420 );
and \U$36315 ( \44122_44422 , \43914_44214 , \43919_44219 );
or \U$36317 ( \44123_44423 , 1'b0 , \44122_44422 , 1'b0 );
xor \U$36318 ( \44124_44424 , \44121_44421 , \44123_44423 );
and \U$36320 ( \44125_44425 , \43907_44207 , \43913_44213 );
and \U$36321 ( \44126_44426 , \43909_44209 , \43913_44213 );
or \U$36322 ( \44127_44427 , 1'b0 , \44125_44425 , \44126_44426 );
xor \U$36323 ( \44128_44428 , \44124_44424 , \44127_44427 );
xor \U$36330 ( \44129_44429 , \44128_44428 , 1'b0 );
and \U$36331 ( \44130_44430 , \43925_44225 , \44113_44413 );
and \U$36332 ( \44131_44431 , \43925_44225 , \44119_44419 );
and \U$36333 ( \44132_44432 , \44113_44413 , \44119_44419 );
or \U$36334 ( \44133_44433 , \44130_44430 , \44131_44431 , \44132_44432 );
xor \U$36335 ( \44134_44434 , \44129_44429 , \44133_44433 );
and \U$36336 ( \44135_44435 , \44026_44326 , \44031_44331 );
and \U$36337 ( \44136_44436 , \44026_44326 , \44111_44411 );
and \U$36338 ( \44137_44437 , \44031_44331 , \44111_44411 );
or \U$36339 ( \44138_44438 , \44135_44435 , \44136_44436 , \44137_44437 );
buf \U$36340 ( \44139_44439 , \44138_44438 );
and \U$36341 ( \44140_44440 , \44011_44311 , \44016_44316 );
and \U$36342 ( \44141_44441 , \44011_44311 , \44022_44322 );
and \U$36343 ( \44142_44442 , \44016_44316 , \44022_44322 );
or \U$36344 ( \44143_44443 , \44140_44440 , \44141_44441 , \44142_44442 );
buf \U$36345 ( \44144_44444 , \44143_44443 );
and \U$36346 ( \44145_44445 , \43940_44240 , \43946_44246 );
and \U$36347 ( \44146_44446 , \43940_44240 , \43953_44253 );
and \U$36348 ( \44147_44447 , \43946_44246 , \43953_44253 );
or \U$36349 ( \44148_44448 , \44145_44445 , \44146_44446 , \44147_44447 );
buf \U$36350 ( \44149_44449 , \44148_44448 );
and \U$36351 ( \44150_44450 , \44064_44364 , \44070_44370 );
and \U$36352 ( \44151_44451 , \44064_44364 , \44077_44377 );
and \U$36353 ( \44152_44452 , \44070_44370 , \44077_44377 );
or \U$36354 ( \44153_44453 , \44150_44450 , \44151_44451 , \44152_44452 );
buf \U$36355 ( \44154_44454 , \44153_44453 );
xor \U$36356 ( \44155_44455 , \44149_44449 , \44154_44454 );
and \U$36357 ( \44156_44456 , \14710_14631 , \42133_42433_nG9b5a );
and \U$36358 ( \44157_44457 , \14329_14628 , \42466_42766_nG9b57 );
or \U$36359 ( \44158_44458 , \44156_44456 , \44157_44457 );
xor \U$36360 ( \44159_44459 , \14328_14627 , \44158_44458 );
buf \U$36361 ( \44160_44460 , \44159_44459 );
buf \U$36363 ( \44161_44461 , \44160_44460 );
xor \U$36364 ( \44162_44462 , \44155_44455 , \44161_44461 );
buf \U$36365 ( \44163_44463 , \44162_44462 );
xor \U$36366 ( \44164_44464 , \44144_44444 , \44163_44463 );
and \U$36367 ( \44165_44465 , \30670_29853 , \35872_36172_nG9b96 );
and \U$36368 ( \44166_44466 , \29551_29850 , \36289_36589_nG9b93 );
or \U$36369 ( \44167_44467 , \44165_44465 , \44166_44466 );
xor \U$36370 ( \44168_44468 , \29550_29849 , \44167_44467 );
buf \U$36371 ( \44169_44469 , \44168_44468 );
buf \U$36373 ( \44170_44470 , \44169_44469 );
and \U$36374 ( \44171_44471 , \28946_28118 , \36686_36986_nG9b90 );
and \U$36375 ( \44172_44472 , \27816_28115 , \36950_37250_nG9b8d );
or \U$36376 ( \44173_44473 , \44171_44471 , \44172_44472 );
xor \U$36377 ( \44174_44474 , \27815_28114 , \44173_44473 );
buf \U$36378 ( \44175_44475 , \44174_44474 );
buf \U$36380 ( \44176_44476 , \44175_44475 );
xor \U$36381 ( \44177_44477 , \44170_44470 , \44176_44476 );
and \U$36382 ( \44178_44478 , \27141_26431 , \37307_37607_nG9b8a );
and \U$36383 ( \44179_44479 , \26129_26428 , \37674_37974_nG9b87 );
or \U$36384 ( \44180_44480 , \44178_44478 , \44179_44479 );
xor \U$36385 ( \44181_44481 , \26128_26427 , \44180_44480 );
buf \U$36386 ( \44182_44482 , \44181_44481 );
buf \U$36388 ( \44183_44483 , \44182_44482 );
xor \U$36389 ( \44184_44484 , \44177_44477 , \44183_44483 );
buf \U$36390 ( \44185_44485 , \44184_44484 );
buf \U$36391 ( \44186_44486 , \44001_44301 );
and \U$36392 ( \44187_44487 , \20353_20155 , \39904_40204_nG9b72 );
and \U$36393 ( \44188_44488 , \19853_20152 , \40152_40452_nG9b6f );
or \U$36394 ( \44189_44489 , \44187_44487 , \44188_44488 );
xor \U$36395 ( \44190_44490 , \19852_20151 , \44189_44489 );
buf \U$36396 ( \44191_44491 , \44190_44490 );
buf \U$36398 ( \44192_44492 , \44191_44491 );
xor \U$36399 ( \44193_44493 , \44186_44486 , \44192_44492 );
and \U$36400 ( \44194_44494 , \18908_18702 , \40543_40843_nG9b6c );
and \U$36401 ( \44195_44495 , \18400_18699 , \40740_41040_nG9b69 );
or \U$36402 ( \44196_44496 , \44194_44494 , \44195_44495 );
xor \U$36403 ( \44197_44497 , \18399_18698 , \44196_44496 );
buf \U$36404 ( \44198_44498 , \44197_44497 );
buf \U$36406 ( \44199_44499 , \44198_44498 );
xor \U$36407 ( \44200_44500 , \44193_44493 , \44199_44499 );
buf \U$36408 ( \44201_44501 , \44200_44500 );
xor \U$36409 ( \44202_44502 , \44185_44485 , \44201_44501 );
and \U$36410 ( \44203_44503 , \43995_44295 , \44002_44302 );
and \U$36411 ( \44204_44504 , \43995_44295 , \44009_44309 );
and \U$36412 ( \44205_44505 , \44002_44302 , \44009_44309 );
or \U$36413 ( \44206_44506 , \44203_44503 , \44204_44504 , \44205_44505 );
buf \U$36414 ( \44207_44507 , \44206_44506 );
xor \U$36415 ( \44208_44508 , \44202_44502 , \44207_44507 );
buf \U$36416 ( \44209_44509 , \44208_44508 );
xor \U$36417 ( \44210_44510 , \44164_44464 , \44209_44509 );
buf \U$36418 ( \44211_44511 , \44210_44510 );
and \U$36419 ( \44212_44512 , \44037_44337 , \44103_44403 );
and \U$36420 ( \44213_44513 , \44037_44337 , \44109_44409 );
and \U$36421 ( \44214_44514 , \44103_44403 , \44109_44409 );
or \U$36422 ( \44215_44515 , \44212_44512 , \44213_44513 , \44214_44514 );
buf \U$36423 ( \44216_44516 , \44215_44515 );
xor \U$36424 ( \44217_44517 , \44211_44511 , \44216_44516 );
and \U$36425 ( \44218_44518 , \43930_44230 , \43989_44289 );
and \U$36426 ( \44219_44519 , \43930_44230 , \44024_44324 );
and \U$36427 ( \44220_44520 , \43989_44289 , \44024_44324 );
or \U$36428 ( \44221_44521 , \44218_44518 , \44219_44519 , \44220_44520 );
buf \U$36429 ( \44222_44522 , \44221_44521 );
xor \U$36430 ( \44223_44523 , \44217_44517 , \44222_44522 );
buf \U$36431 ( \44224_44524 , \44223_44523 );
xor \U$36432 ( \44225_44525 , \44139_44439 , \44224_44524 );
and \U$36433 ( \44226_44526 , \43935_44235 , \43968_44268 );
and \U$36434 ( \44227_44527 , \43935_44235 , \43987_44287 );
and \U$36435 ( \44228_44528 , \43968_44268 , \43987_44287 );
or \U$36436 ( \44229_44529 , \44226_44526 , \44227_44527 , \44228_44528 );
buf \U$36437 ( \44230_44530 , \44229_44529 );
and \U$36438 ( \44231_44531 , \44058_44358 , \44079_44379 );
and \U$36439 ( \44232_44532 , \44058_44358 , \44101_44401 );
and \U$36440 ( \44233_44533 , \44079_44379 , \44101_44401 );
or \U$36441 ( \44234_44534 , \44231_44531 , \44232_44532 , \44233_44533 );
buf \U$36442 ( \44235_44535 , \44234_44534 );
and \U$36443 ( \44236_44536 , \44043_44343 , \44049_44349 );
and \U$36444 ( \44237_44537 , \44043_44343 , \44056_44356 );
and \U$36445 ( \44238_44538 , \44049_44349 , \44056_44356 );
or \U$36446 ( \44239_44539 , \44236_44536 , \44237_44537 , \44238_44538 );
buf \U$36447 ( \44240_44540 , \44239_44539 );
and \U$36448 ( \44241_44541 , \44086_44386 , \44092_44392 );
and \U$36449 ( \44242_44542 , \44086_44386 , \44099_44399 );
and \U$36450 ( \44243_44543 , \44092_44392 , \44099_44399 );
or \U$36451 ( \44244_44544 , \44241_44541 , \44242_44542 , \44243_44543 );
buf \U$36452 ( \44245_44545 , \44244_44544 );
xor \U$36453 ( \44246_44546 , \44240_44540 , \44245_44545 );
xor \U$36457 ( \44247_44547 , \11854_12153 , 1'b0 );
not \U$36458 ( \44248_44548 , \44247_44547 );
buf \U$36459 ( \44249_44549 , \44248_44548 );
buf \U$36461 ( \44250_44550 , \44249_44549 );
and \U$36463 ( \44251_44551 , \32617_32916 , \34794_35094_nG9b9f );
or \U$36464 ( \44252_44552 , 1'b0 , \44251_44551 );
xor \U$36465 ( \44253_44553 , 1'b0 , \44252_44552 );
buf \U$36466 ( \44254_44554 , \44253_44553 );
buf \U$36468 ( \44255_44555 , \44254_44554 );
xor \U$36469 ( \44256_44556 , \44250_44550 , \44255_44555 );
and \U$36470 ( \44257_44557 , \31989_31636 , \35270_35570_nG9b9c );
and \U$36471 ( \44258_44558 , \31334_31633 , \35501_35801_nG9b99 );
or \U$36472 ( \44259_44559 , \44257_44557 , \44258_44558 );
xor \U$36473 ( \44260_44560 , \31333_31632 , \44259_44559 );
buf \U$36474 ( \44261_44561 , \44260_44560 );
buf \U$36476 ( \44262_44562 , \44261_44561 );
xor \U$36477 ( \44263_44563 , \44256_44556 , \44262_44562 );
buf \U$36478 ( \44264_44564 , \44263_44563 );
xor \U$36479 ( \44265_44565 , \44246_44546 , \44264_44564 );
buf \U$36480 ( \44266_44566 , \44265_44565 );
xor \U$36481 ( \44267_44567 , \44235_44535 , \44266_44566 );
and \U$36482 ( \44268_44568 , \43955_44255 , \43960_44260 );
and \U$36483 ( \44269_44569 , \43955_44255 , \43966_44266 );
and \U$36484 ( \44270_44570 , \43960_44260 , \43966_44266 );
or \U$36485 ( \44271_44571 , \44268_44568 , \44269_44569 , \44270_44570 );
buf \U$36486 ( \44272_44572 , \44271_44571 );
xor \U$36487 ( \44273_44573 , \44267_44567 , \44272_44572 );
buf \U$36488 ( \44274_44574 , \44273_44573 );
xor \U$36489 ( \44275_44575 , \44230_44530 , \44274_44574 );
and \U$36490 ( \44276_44576 , \43974_44274 , \43979_44279 );
and \U$36491 ( \44277_44577 , \43974_44274 , \43985_44285 );
and \U$36492 ( \44278_44578 , \43979_44279 , \43985_44285 );
or \U$36493 ( \44279_44579 , \44276_44576 , \44277_44577 , \44278_44578 );
buf \U$36494 ( \44280_44580 , \44279_44579 );
and \U$36495 ( \44281_44581 , \25044_24792 , \38037_38337_nG9b84 );
and \U$36496 ( \44282_44582 , \24490_24789 , \38363_38663_nG9b81 );
or \U$36497 ( \44283_44583 , \44281_44581 , \44282_44582 );
xor \U$36498 ( \44284_44584 , \24489_24788 , \44283_44583 );
buf \U$36499 ( \44285_44585 , \44284_44584 );
buf \U$36501 ( \44286_44586 , \44285_44585 );
and \U$36502 ( \44287_44587 , \23495_23201 , \38668_38968_nG9b7e );
and \U$36503 ( \44288_44588 , \22899_23198 , \39034_39334_nG9b7b );
or \U$36504 ( \44289_44589 , \44287_44587 , \44288_44588 );
xor \U$36505 ( \44290_44590 , \22898_23197 , \44289_44589 );
buf \U$36506 ( \44291_44591 , \44290_44590 );
buf \U$36508 ( \44292_44592 , \44291_44591 );
xor \U$36509 ( \44293_44593 , \44286_44586 , \44292_44592 );
and \U$36510 ( \44294_44594 , \17437_17297 , \41081_41381_nG9b66 );
and \U$36511 ( \44295_44595 , \16995_17294 , \41385_41685_nG9b63 );
or \U$36512 ( \44296_44596 , \44294_44594 , \44295_44595 );
xor \U$36513 ( \44297_44597 , \16994_17293 , \44296_44596 );
buf \U$36514 ( \44298_44598 , \44297_44597 );
buf \U$36516 ( \44299_44599 , \44298_44598 );
xor \U$36517 ( \44300_44600 , \44293_44593 , \44299_44599 );
buf \U$36518 ( \44301_44601 , \44300_44600 );
xor \U$36519 ( \44302_44602 , \44280_44580 , \44301_44601 );
and \U$36520 ( \44303_44603 , \13431_13370 , \42548_42848_nG9b54 );
and \U$36521 ( \44304_44604 , \13068_13367 , \42879_43179_nG9b51 );
or \U$36522 ( \44305_44605 , \44303_44603 , \44304_44604 );
xor \U$36523 ( \44306_44606 , \13067_13366 , \44305_44605 );
buf \U$36524 ( \44307_44607 , \44306_44606 );
buf \U$36526 ( \44308_44608 , \44307_44607 );
and \U$36527 ( \44309_44609 , \21908_21658 , \39291_39591_nG9b78 );
and \U$36528 ( \44310_44610 , \21356_21655 , \39663_39963_nG9b75 );
or \U$36529 ( \44311_44611 , \44309_44609 , \44310_44610 );
xor \U$36530 ( \44312_44612 , \21355_21654 , \44311_44611 );
buf \U$36531 ( \44313_44613 , \44312_44612 );
buf \U$36533 ( \44314_44614 , \44313_44613 );
xor \U$36534 ( \44315_44615 , \44308_44608 , \44314_44614 );
and \U$36535 ( \44316_44616 , \16405_15940 , \41663_41963_nG9b60 );
and \U$36536 ( \44317_44617 , \15638_15937 , \41901_42201_nG9b5d );
or \U$36537 ( \44318_44618 , \44316_44616 , \44317_44617 );
xor \U$36538 ( \44319_44619 , \15637_15936 , \44318_44618 );
buf \U$36539 ( \44320_44620 , \44319_44619 );
buf \U$36541 ( \44321_44621 , \44320_44620 );
xor \U$36542 ( \44322_44622 , \44315_44615 , \44321_44621 );
buf \U$36543 ( \44323_44623 , \44322_44622 );
xor \U$36544 ( \44324_44624 , \44302_44602 , \44323_44623 );
buf \U$36545 ( \44325_44625 , \44324_44624 );
xor \U$36546 ( \44326_44626 , \44275_44575 , \44325_44625 );
buf \U$36547 ( \44327_44627 , \44326_44626 );
xor \U$36548 ( \44328_44628 , \44225_44525 , \44327_44627 );
and \U$36549 ( \44329_44629 , \44134_44434 , \44328_44628 );
and \U$36551 ( \44330_44630 , \44128_44428 , \44133_44433 );
or \U$36553 ( \44331_44631 , 1'b0 , \44330_44630 , 1'b0 );
xor \U$36554 ( \44332_44632 , \44329_44629 , \44331_44631 );
and \U$36556 ( \44333_44633 , \44121_44421 , \44127_44427 );
and \U$36557 ( \44334_44634 , \44123_44423 , \44127_44427 );
or \U$36558 ( \44335_44635 , 1'b0 , \44333_44633 , \44334_44634 );
xor \U$36559 ( \44336_44636 , \44332_44632 , \44335_44635 );
xor \U$36566 ( \44337_44637 , \44336_44636 , 1'b0 );
and \U$36567 ( \44338_44638 , \44139_44439 , \44224_44524 );
and \U$36568 ( \44339_44639 , \44139_44439 , \44327_44627 );
and \U$36569 ( \44340_44640 , \44224_44524 , \44327_44627 );
or \U$36570 ( \44341_44641 , \44338_44638 , \44339_44639 , \44340_44640 );
xor \U$36571 ( \44342_44642 , \44337_44637 , \44341_44641 );
and \U$36572 ( \44343_44643 , \44211_44511 , \44216_44516 );
and \U$36573 ( \44344_44644 , \44211_44511 , \44222_44522 );
and \U$36574 ( \44345_44645 , \44216_44516 , \44222_44522 );
or \U$36575 ( \44346_44646 , \44343_44643 , \44344_44644 , \44345_44645 );
buf \U$36576 ( \44347_44647 , \44346_44646 );
and \U$36577 ( \44348_44648 , \44230_44530 , \44274_44574 );
and \U$36578 ( \44349_44649 , \44230_44530 , \44325_44625 );
and \U$36579 ( \44350_44650 , \44274_44574 , \44325_44625 );
or \U$36580 ( \44351_44651 , \44348_44648 , \44349_44649 , \44350_44650 );
buf \U$36581 ( \44352_44652 , \44351_44651 );
and \U$36582 ( \44353_44653 , \44144_44444 , \44163_44463 );
and \U$36583 ( \44354_44654 , \44144_44444 , \44209_44509 );
and \U$36584 ( \44355_44655 , \44163_44463 , \44209_44509 );
or \U$36585 ( \44356_44656 , \44353_44653 , \44354_44654 , \44355_44655 );
buf \U$36586 ( \44357_44657 , \44356_44656 );
xor \U$36587 ( \44358_44658 , \44352_44652 , \44357_44657 );
and \U$36588 ( \44359_44659 , \44250_44550 , \44255_44555 );
and \U$36589 ( \44360_44660 , \44250_44550 , \44262_44562 );
and \U$36590 ( \44361_44661 , \44255_44555 , \44262_44562 );
or \U$36591 ( \44362_44662 , \44359_44659 , \44360_44660 , \44361_44661 );
buf \U$36592 ( \44363_44663 , \44362_44662 );
and \U$36593 ( \44364_44664 , \31989_31636 , \35501_35801_nG9b99 );
and \U$36594 ( \44365_44665 , \31334_31633 , \35872_36172_nG9b96 );
or \U$36595 ( \44366_44666 , \44364_44664 , \44365_44665 );
xor \U$36596 ( \44367_44667 , \31333_31632 , \44366_44666 );
buf \U$36597 ( \44368_44668 , \44367_44667 );
buf \U$36598 ( \44369_44669 , \44368_44668 );
not \U$36599 ( \44370_44670 , \44369_44669 );
xor \U$36600 ( \44371_44671 , \44363_44663 , \44370_44670 );
and \U$36601 ( \44372_44672 , \14710_14631 , \42466_42766_nG9b57 );
and \U$36602 ( \44373_44673 , \14329_14628 , \42548_42848_nG9b54 );
or \U$36603 ( \44374_44674 , \44372_44672 , \44373_44673 );
xor \U$36604 ( \44375_44675 , \14328_14627 , \44374_44674 );
buf \U$36605 ( \44376_44676 , \44375_44675 );
buf \U$36607 ( \44377_44677 , \44376_44676 );
xor \U$36608 ( \44378_44678 , \44371_44671 , \44377_44677 );
buf \U$36609 ( \44379_44679 , \44378_44678 );
and \U$36610 ( \44380_44680 , \27141_26431 , \37674_37974_nG9b87 );
and \U$36611 ( \44381_44681 , \26129_26428 , \38037_38337_nG9b84 );
or \U$36612 ( \44382_44682 , \44380_44680 , \44381_44681 );
xor \U$36613 ( \44383_44683 , \26128_26427 , \44382_44682 );
buf \U$36614 ( \44384_44684 , \44383_44683 );
buf \U$36616 ( \44385_44685 , \44384_44684 );
and \U$36617 ( \44386_44686 , \25044_24792 , \38363_38663_nG9b81 );
and \U$36618 ( \44387_44687 , \24490_24789 , \38668_38968_nG9b7e );
or \U$36619 ( \44388_44688 , \44386_44686 , \44387_44687 );
xor \U$36620 ( \44389_44689 , \24489_24788 , \44388_44688 );
buf \U$36621 ( \44390_44690 , \44389_44689 );
buf \U$36623 ( \44391_44691 , \44390_44690 );
xor \U$36624 ( \44392_44692 , \44385_44685 , \44391_44691 );
and \U$36625 ( \44393_44693 , \18908_18702 , \40740_41040_nG9b69 );
and \U$36626 ( \44394_44694 , \18400_18699 , \41081_41381_nG9b66 );
or \U$36627 ( \44395_44695 , \44393_44693 , \44394_44694 );
xor \U$36628 ( \44396_44696 , \18399_18698 , \44395_44695 );
buf \U$36629 ( \44397_44697 , \44396_44696 );
buf \U$36631 ( \44398_44698 , \44397_44697 );
xor \U$36632 ( \44399_44699 , \44392_44692 , \44398_44698 );
buf \U$36633 ( \44400_44700 , \44399_44699 );
xor \U$36634 ( \44401_44701 , \44379_44679 , \44400_44700 );
and \U$36635 ( \44402_44702 , \30670_29853 , \36289_36589_nG9b93 );
and \U$36636 ( \44403_44703 , \29551_29850 , \36686_36986_nG9b90 );
or \U$36637 ( \44404_44704 , \44402_44702 , \44403_44703 );
xor \U$36638 ( \44405_44705 , \29550_29849 , \44404_44704 );
buf \U$36639 ( \44406_44706 , \44405_44705 );
buf \U$36641 ( \44407_44707 , \44406_44706 );
and \U$36642 ( \44408_44708 , \28946_28118 , \36950_37250_nG9b8d );
and \U$36643 ( \44409_44709 , \27816_28115 , \37307_37607_nG9b8a );
or \U$36644 ( \44410_44710 , \44408_44708 , \44409_44709 );
xor \U$36645 ( \44411_44711 , \27815_28114 , \44410_44710 );
buf \U$36646 ( \44412_44712 , \44411_44711 );
buf \U$36648 ( \44413_44713 , \44412_44712 );
xor \U$36649 ( \44414_44714 , \44407_44707 , \44413_44713 );
and \U$36650 ( \44415_44715 , \16405_15940 , \41901_42201_nG9b5d );
and \U$36651 ( \44416_44716 , \15638_15937 , \42133_42433_nG9b5a );
or \U$36652 ( \44417_44717 , \44415_44715 , \44416_44716 );
xor \U$36653 ( \44418_44718 , \15637_15936 , \44417_44717 );
buf \U$36654 ( \44419_44719 , \44418_44718 );
buf \U$36656 ( \44420_44720 , \44419_44719 );
xor \U$36657 ( \44421_44721 , \44414_44714 , \44420_44720 );
buf \U$36658 ( \44422_44722 , \44421_44721 );
xor \U$36659 ( \44423_44723 , \44401_44701 , \44422_44722 );
buf \U$36660 ( \44424_44724 , \44423_44723 );
and \U$36661 ( \44425_44725 , \13431_13370 , \42879_43179_nG9b51 );
or \U$36663 ( \44426_44726 , \44425_44725 , 1'b0 );
xor \U$36664 ( \44427_44727 , \13067_13366 , \44426_44726 );
buf \U$36665 ( \44428_44728 , \44427_44727 );
buf \U$36667 ( \44429_44729 , \44428_44728 );
and \U$36668 ( \44430_44730 , \21908_21658 , \39663_39963_nG9b75 );
and \U$36669 ( \44431_44731 , \21356_21655 , \39904_40204_nG9b72 );
or \U$36670 ( \44432_44732 , \44430_44730 , \44431_44731 );
xor \U$36671 ( \44433_44733 , \21355_21654 , \44432_44732 );
buf \U$36672 ( \44434_44734 , \44433_44733 );
buf \U$36674 ( \44435_44735 , \44434_44734 );
xor \U$36675 ( \44436_44736 , \44429_44729 , \44435_44735 );
and \U$36676 ( \44437_44737 , \20353_20155 , \40152_40452_nG9b6f );
and \U$36677 ( \44438_44738 , \19853_20152 , \40543_40843_nG9b6c );
or \U$36678 ( \44439_44739 , \44437_44737 , \44438_44738 );
xor \U$36679 ( \44440_44740 , \19852_20151 , \44439_44739 );
buf \U$36680 ( \44441_44741 , \44440_44740 );
buf \U$36682 ( \44442_44742 , \44441_44741 );
xor \U$36683 ( \44443_44743 , \44436_44736 , \44442_44742 );
buf \U$36684 ( \44444_44744 , \44443_44743 );
and \U$36685 ( \44445_44745 , \44186_44486 , \44192_44492 );
and \U$36686 ( \44446_44746 , \44186_44486 , \44199_44499 );
and \U$36687 ( \44447_44747 , \44192_44492 , \44199_44499 );
or \U$36688 ( \44448_44748 , \44445_44745 , \44446_44746 , \44447_44747 );
buf \U$36689 ( \44449_44749 , \44448_44748 );
xor \U$36690 ( \44450_44750 , \44444_44744 , \44449_44749 );
and \U$36692 ( \44451_44751 , \32617_32916 , \35270_35570_nG9b9c );
or \U$36693 ( \44452_44752 , 1'b0 , \44451_44751 );
xor \U$36694 ( \44453_44753 , 1'b0 , \44452_44752 );
buf \U$36695 ( \44454_44754 , \44453_44753 );
buf \U$36697 ( \44455_44755 , \44454_44754 );
and \U$36698 ( \44456_44756 , \23495_23201 , \39034_39334_nG9b7b );
and \U$36699 ( \44457_44757 , \22899_23198 , \39291_39591_nG9b78 );
or \U$36700 ( \44458_44758 , \44456_44756 , \44457_44757 );
xor \U$36701 ( \44459_44759 , \22898_23197 , \44458_44758 );
buf \U$36702 ( \44460_44760 , \44459_44759 );
buf \U$36704 ( \44461_44761 , \44460_44760 );
xor \U$36705 ( \44462_44762 , \44455_44755 , \44461_44761 );
and \U$36706 ( \44463_44763 , \17437_17297 , \41385_41685_nG9b63 );
and \U$36707 ( \44464_44764 , \16995_17294 , \41663_41963_nG9b60 );
or \U$36708 ( \44465_44765 , \44463_44763 , \44464_44764 );
xor \U$36709 ( \44466_44766 , \16994_17293 , \44465_44765 );
buf \U$36710 ( \44467_44767 , \44466_44766 );
buf \U$36712 ( \44468_44768 , \44467_44767 );
xor \U$36713 ( \44469_44769 , \44462_44762 , \44468_44768 );
buf \U$36714 ( \44470_44770 , \44469_44769 );
xor \U$36715 ( \44471_44771 , \44450_44750 , \44470_44770 );
buf \U$36716 ( \44472_44772 , \44471_44771 );
xor \U$36717 ( \44473_44773 , \44424_44724 , \44472_44772 );
and \U$36718 ( \44474_44774 , \44185_44485 , \44201_44501 );
and \U$36719 ( \44475_44775 , \44185_44485 , \44207_44507 );
and \U$36720 ( \44476_44776 , \44201_44501 , \44207_44507 );
or \U$36721 ( \44477_44777 , \44474_44774 , \44475_44775 , \44476_44776 );
buf \U$36722 ( \44478_44778 , \44477_44777 );
xor \U$36723 ( \44479_44779 , \44473_44773 , \44478_44778 );
buf \U$36724 ( \44480_44780 , \44479_44779 );
xor \U$36725 ( \44481_44781 , \44358_44658 , \44480_44780 );
buf \U$36726 ( \44482_44782 , \44481_44781 );
xor \U$36727 ( \44483_44783 , \44347_44647 , \44482_44782 );
and \U$36728 ( \44484_44784 , \44235_44535 , \44266_44566 );
and \U$36729 ( \44485_44785 , \44235_44535 , \44272_44572 );
and \U$36730 ( \44486_44786 , \44266_44566 , \44272_44572 );
or \U$36731 ( \44487_44787 , \44484_44784 , \44485_44785 , \44486_44786 );
buf \U$36732 ( \44488_44788 , \44487_44787 );
and \U$36733 ( \44489_44789 , \44280_44580 , \44301_44601 );
and \U$36734 ( \44490_44790 , \44280_44580 , \44323_44623 );
and \U$36735 ( \44491_44791 , \44301_44601 , \44323_44623 );
or \U$36736 ( \44492_44792 , \44489_44789 , \44490_44790 , \44491_44791 );
buf \U$36737 ( \44493_44793 , \44492_44792 );
xor \U$36738 ( \44494_44794 , \44488_44788 , \44493_44793 );
and \U$36739 ( \44495_44795 , \44240_44540 , \44245_44545 );
and \U$36740 ( \44496_44796 , \44240_44540 , \44264_44564 );
and \U$36741 ( \44497_44797 , \44245_44545 , \44264_44564 );
or \U$36742 ( \44498_44798 , \44495_44795 , \44496_44796 , \44497_44797 );
buf \U$36743 ( \44499_44799 , \44498_44798 );
and \U$36744 ( \44500_44800 , \44149_44449 , \44154_44454 );
and \U$36745 ( \44501_44801 , \44149_44449 , \44161_44461 );
and \U$36746 ( \44502_44802 , \44154_44454 , \44161_44461 );
or \U$36747 ( \44503_44803 , \44500_44800 , \44501_44801 , \44502_44802 );
buf \U$36748 ( \44504_44804 , \44503_44803 );
xor \U$36749 ( \44505_44805 , \44499_44799 , \44504_44804 );
and \U$36750 ( \44506_44806 , \44308_44608 , \44314_44614 );
and \U$36751 ( \44507_44807 , \44308_44608 , \44321_44621 );
and \U$36752 ( \44508_44808 , \44314_44614 , \44321_44621 );
or \U$36753 ( \44509_44809 , \44506_44806 , \44507_44807 , \44508_44808 );
buf \U$36754 ( \44510_44810 , \44509_44809 );
and \U$36755 ( \44511_44811 , \44170_44470 , \44176_44476 );
and \U$36756 ( \44512_44812 , \44170_44470 , \44183_44483 );
and \U$36757 ( \44513_44813 , \44176_44476 , \44183_44483 );
or \U$36758 ( \44514_44814 , \44511_44811 , \44512_44812 , \44513_44813 );
buf \U$36759 ( \44515_44815 , \44514_44814 );
xor \U$36760 ( \44516_44816 , \44510_44810 , \44515_44815 );
and \U$36761 ( \44517_44817 , \44286_44586 , \44292_44592 );
and \U$36762 ( \44518_44818 , \44286_44586 , \44299_44599 );
and \U$36763 ( \44519_44819 , \44292_44592 , \44299_44599 );
or \U$36764 ( \44520_44820 , \44517_44817 , \44518_44818 , \44519_44819 );
buf \U$36765 ( \44521_44821 , \44520_44820 );
xor \U$36766 ( \44522_44822 , \44516_44816 , \44521_44821 );
buf \U$36767 ( \44523_44823 , \44522_44822 );
xor \U$36768 ( \44524_44824 , \44505_44805 , \44523_44823 );
buf \U$36769 ( \44525_44825 , \44524_44824 );
xor \U$36770 ( \44526_44826 , \44494_44794 , \44525_44825 );
buf \U$36771 ( \44527_44827 , \44526_44826 );
xor \U$36772 ( \44528_44828 , \44483_44783 , \44527_44827 );
and \U$36773 ( \44529_44829 , \44342_44642 , \44528_44828 );
and \U$36775 ( \44530_44830 , \44336_44636 , \44341_44641 );
or \U$36777 ( \44531_44831 , 1'b0 , \44530_44830 , 1'b0 );
xor \U$36778 ( \44532_44832 , \44529_44829 , \44531_44831 );
and \U$36780 ( \44533_44833 , \44329_44629 , \44335_44635 );
and \U$36781 ( \44534_44834 , \44331_44631 , \44335_44635 );
or \U$36782 ( \44535_44835 , 1'b0 , \44533_44833 , \44534_44834 );
xor \U$36783 ( \44536_44836 , \44532_44832 , \44535_44835 );
xor \U$36790 ( \44537_44837 , \44536_44836 , 1'b0 );
and \U$36791 ( \44538_44838 , \44352_44652 , \44357_44657 );
and \U$36792 ( \44539_44839 , \44352_44652 , \44480_44780 );
and \U$36793 ( \44540_44840 , \44357_44657 , \44480_44780 );
or \U$36794 ( \44541_44841 , \44538_44838 , \44539_44839 , \44540_44840 );
buf \U$36795 ( \44542_44842 , \44541_44841 );
and \U$36796 ( \44543_44843 , \44510_44810 , \44515_44815 );
and \U$36797 ( \44544_44844 , \44510_44810 , \44521_44821 );
and \U$36798 ( \44545_44845 , \44515_44815 , \44521_44821 );
or \U$36799 ( \44546_44846 , \44543_44843 , \44544_44844 , \44545_44845 );
buf \U$36800 ( \44547_44847 , \44546_44846 );
and \U$36801 ( \44548_44848 , \25044_24792 , \38668_38968_nG9b7e );
and \U$36802 ( \44549_44849 , \24490_24789 , \39034_39334_nG9b7b );
or \U$36803 ( \44550_44850 , \44548_44848 , \44549_44849 );
xor \U$36804 ( \44551_44851 , \24489_24788 , \44550_44850 );
buf \U$36805 ( \44552_44852 , \44551_44851 );
buf \U$36807 ( \44553_44853 , \44552_44852 );
and \U$36808 ( \44554_44854 , \23495_23201 , \39291_39591_nG9b78 );
and \U$36809 ( \44555_44855 , \22899_23198 , \39663_39963_nG9b75 );
or \U$36810 ( \44556_44856 , \44554_44854 , \44555_44855 );
xor \U$36811 ( \44557_44857 , \22898_23197 , \44556_44856 );
buf \U$36812 ( \44558_44858 , \44557_44857 );
buf \U$36814 ( \44559_44859 , \44558_44858 );
xor \U$36815 ( \44560_44860 , \44553_44853 , \44559_44859 );
and \U$36816 ( \44561_44861 , \17437_17297 , \41663_41963_nG9b60 );
and \U$36817 ( \44562_44862 , \16995_17294 , \41901_42201_nG9b5d );
or \U$36818 ( \44563_44863 , \44561_44861 , \44562_44862 );
xor \U$36819 ( \44564_44864 , \16994_17293 , \44563_44863 );
buf \U$36820 ( \44565_44865 , \44564_44864 );
buf \U$36822 ( \44566_44866 , \44565_44865 );
xor \U$36823 ( \44567_44867 , \44560_44860 , \44566_44866 );
buf \U$36824 ( \44568_44868 , \44567_44867 );
and \U$36825 ( \44569_44869 , \44429_44729 , \44435_44735 );
and \U$36826 ( \44570_44870 , \44429_44729 , \44442_44742 );
and \U$36827 ( \44571_44871 , \44435_44735 , \44442_44742 );
or \U$36828 ( \44572_44872 , \44569_44869 , \44570_44870 , \44571_44871 );
buf \U$36829 ( \44573_44873 , \44572_44872 );
xor \U$36830 ( \44574_44874 , \44568_44868 , \44573_44873 );
and \U$36831 ( \44575_44875 , \14710_14631 , \42548_42848_nG9b54 );
and \U$36832 ( \44576_44876 , \14329_14628 , \42879_43179_nG9b51 );
or \U$36833 ( \44577_44877 , \44575_44875 , \44576_44876 );
xor \U$36834 ( \44578_44878 , \14328_14627 , \44577_44877 );
buf \U$36835 ( \44579_44879 , \44578_44878 );
buf \U$36837 ( \44580_44880 , \44579_44879 );
xor \U$36841 ( \44581_44881 , \13067_13366 , 1'b0 );
not \U$36842 ( \44582_44882 , \44581_44881 );
buf \U$36843 ( \44583_44883 , \44582_44882 );
buf \U$36845 ( \44584_44884 , \44583_44883 );
xor \U$36846 ( \44585_44885 , \44580_44880 , \44584_44884 );
and \U$36848 ( \44586_44886 , \32617_32916 , \35501_35801_nG9b99 );
or \U$36849 ( \44587_44887 , 1'b0 , \44586_44886 );
xor \U$36850 ( \44588_44888 , 1'b0 , \44587_44887 );
buf \U$36851 ( \44589_44889 , \44588_44888 );
buf \U$36853 ( \44590_44890 , \44589_44889 );
xor \U$36854 ( \44591_44891 , \44585_44885 , \44590_44890 );
buf \U$36855 ( \44592_44892 , \44591_44891 );
xor \U$36856 ( \44593_44893 , \44574_44874 , \44592_44892 );
buf \U$36857 ( \44594_44894 , \44593_44893 );
xor \U$36858 ( \44595_44895 , \44547_44847 , \44594_44894 );
and \U$36859 ( \44596_44896 , \44363_44663 , \44370_44670 );
and \U$36860 ( \44597_44897 , \44363_44663 , \44377_44677 );
and \U$36861 ( \44598_44898 , \44370_44670 , \44377_44677 );
or \U$36862 ( \44599_44899 , \44596_44896 , \44597_44897 , \44598_44898 );
buf \U$36863 ( \44600_44900 , \44599_44899 );
xor \U$36864 ( \44601_44901 , \44595_44895 , \44600_44900 );
buf \U$36865 ( \44602_44902 , \44601_44901 );
and \U$36866 ( \44603_44903 , \44499_44799 , \44504_44804 );
and \U$36867 ( \44604_44904 , \44499_44799 , \44523_44823 );
and \U$36868 ( \44605_44905 , \44504_44804 , \44523_44823 );
or \U$36869 ( \44606_44906 , \44603_44903 , \44604_44904 , \44605_44905 );
buf \U$36870 ( \44607_44907 , \44606_44906 );
xor \U$36871 ( \44608_44908 , \44602_44902 , \44607_44907 );
and \U$36872 ( \44609_44909 , \28946_28118 , \37307_37607_nG9b8a );
and \U$36873 ( \44610_44910 , \27816_28115 , \37674_37974_nG9b87 );
or \U$36874 ( \44611_44911 , \44609_44909 , \44610_44910 );
xor \U$36875 ( \44612_44912 , \27815_28114 , \44611_44911 );
buf \U$36876 ( \44613_44913 , \44612_44912 );
buf \U$36878 ( \44614_44914 , \44613_44913 );
and \U$36879 ( \44615_44915 , \27141_26431 , \38037_38337_nG9b84 );
and \U$36880 ( \44616_44916 , \26129_26428 , \38363_38663_nG9b81 );
or \U$36881 ( \44617_44917 , \44615_44915 , \44616_44916 );
xor \U$36882 ( \44618_44918 , \26128_26427 , \44617_44917 );
buf \U$36883 ( \44619_44919 , \44618_44918 );
buf \U$36885 ( \44620_44920 , \44619_44919 );
xor \U$36886 ( \44621_44921 , \44614_44914 , \44620_44920 );
and \U$36887 ( \44622_44922 , \18908_18702 , \41081_41381_nG9b66 );
and \U$36888 ( \44623_44923 , \18400_18699 , \41385_41685_nG9b63 );
or \U$36889 ( \44624_44924 , \44622_44922 , \44623_44923 );
xor \U$36890 ( \44625_44925 , \18399_18698 , \44624_44924 );
buf \U$36891 ( \44626_44926 , \44625_44925 );
buf \U$36893 ( \44627_44927 , \44626_44926 );
xor \U$36894 ( \44628_44928 , \44621_44921 , \44627_44927 );
buf \U$36895 ( \44629_44929 , \44628_44928 );
buf \U$36896 ( \44630_44930 , \44369_44669 );
and \U$36897 ( \44631_44931 , \21908_21658 , \39904_40204_nG9b72 );
and \U$36898 ( \44632_44932 , \21356_21655 , \40152_40452_nG9b6f );
or \U$36899 ( \44633_44933 , \44631_44931 , \44632_44932 );
xor \U$36900 ( \44634_44934 , \21355_21654 , \44633_44933 );
buf \U$36901 ( \44635_44935 , \44634_44934 );
buf \U$36903 ( \44636_44936 , \44635_44935 );
xor \U$36904 ( \44637_44937 , \44630_44930 , \44636_44936 );
and \U$36905 ( \44638_44938 , \16405_15940 , \42133_42433_nG9b5a );
and \U$36906 ( \44639_44939 , \15638_15937 , \42466_42766_nG9b57 );
or \U$36907 ( \44640_44940 , \44638_44938 , \44639_44939 );
xor \U$36908 ( \44641_44941 , \15637_15936 , \44640_44940 );
buf \U$36909 ( \44642_44942 , \44641_44941 );
buf \U$36911 ( \44643_44943 , \44642_44942 );
xor \U$36912 ( \44644_44944 , \44637_44937 , \44643_44943 );
buf \U$36913 ( \44645_44945 , \44644_44944 );
xor \U$36914 ( \44646_44946 , \44629_44929 , \44645_44945 );
and \U$36915 ( \44647_44947 , \31989_31636 , \35872_36172_nG9b96 );
and \U$36916 ( \44648_44948 , \31334_31633 , \36289_36589_nG9b93 );
or \U$36917 ( \44649_44949 , \44647_44947 , \44648_44948 );
xor \U$36918 ( \44650_44950 , \31333_31632 , \44649_44949 );
buf \U$36919 ( \44651_44951 , \44650_44950 );
buf \U$36921 ( \44652_44952 , \44651_44951 );
and \U$36922 ( \44653_44953 , \30670_29853 , \36686_36986_nG9b90 );
and \U$36923 ( \44654_44954 , \29551_29850 , \36950_37250_nG9b8d );
or \U$36924 ( \44655_44955 , \44653_44953 , \44654_44954 );
xor \U$36925 ( \44656_44956 , \29550_29849 , \44655_44955 );
buf \U$36926 ( \44657_44957 , \44656_44956 );
buf \U$36928 ( \44658_44958 , \44657_44957 );
xor \U$36929 ( \44659_44959 , \44652_44952 , \44658_44958 );
and \U$36930 ( \44660_44960 , \20353_20155 , \40543_40843_nG9b6c );
and \U$36931 ( \44661_44961 , \19853_20152 , \40740_41040_nG9b69 );
or \U$36932 ( \44662_44962 , \44660_44960 , \44661_44961 );
xor \U$36933 ( \44663_44963 , \19852_20151 , \44662_44962 );
buf \U$36934 ( \44664_44964 , \44663_44963 );
buf \U$36936 ( \44665_44965 , \44664_44964 );
xor \U$36937 ( \44666_44966 , \44659_44959 , \44665_44965 );
buf \U$36938 ( \44667_44967 , \44666_44966 );
xor \U$36939 ( \44668_44968 , \44646_44946 , \44667_44967 );
buf \U$36940 ( \44669_44969 , \44668_44968 );
xor \U$36941 ( \44670_44970 , \44608_44908 , \44669_44969 );
buf \U$36942 ( \44671_44971 , \44670_44970 );
xor \U$36943 ( \44672_44972 , \44542_44842 , \44671_44971 );
and \U$36944 ( \44673_44973 , \44488_44788 , \44493_44793 );
and \U$36945 ( \44674_44974 , \44488_44788 , \44525_44825 );
and \U$36946 ( \44675_44975 , \44493_44793 , \44525_44825 );
or \U$36947 ( \44676_44976 , \44673_44973 , \44674_44974 , \44675_44975 );
buf \U$36948 ( \44677_44977 , \44676_44976 );
and \U$36949 ( \44678_44978 , \44424_44724 , \44472_44772 );
and \U$36950 ( \44679_44979 , \44424_44724 , \44478_44778 );
and \U$36951 ( \44680_44980 , \44472_44772 , \44478_44778 );
or \U$36952 ( \44681_44981 , \44678_44978 , \44679_44979 , \44680_44980 );
buf \U$36953 ( \44682_44982 , \44681_44981 );
xor \U$36954 ( \44683_44983 , \44677_44977 , \44682_44982 );
and \U$36955 ( \44684_44984 , \44444_44744 , \44449_44749 );
and \U$36956 ( \44685_44985 , \44444_44744 , \44470_44770 );
and \U$36957 ( \44686_44986 , \44449_44749 , \44470_44770 );
or \U$36958 ( \44687_44987 , \44684_44984 , \44685_44985 , \44686_44986 );
buf \U$36959 ( \44688_44988 , \44687_44987 );
and \U$36960 ( \44689_44989 , \44385_44685 , \44391_44691 );
and \U$36961 ( \44690_44990 , \44385_44685 , \44398_44698 );
and \U$36962 ( \44691_44991 , \44391_44691 , \44398_44698 );
or \U$36963 ( \44692_44992 , \44689_44989 , \44690_44990 , \44691_44991 );
buf \U$36964 ( \44693_44993 , \44692_44992 );
and \U$36965 ( \44694_44994 , \44455_44755 , \44461_44761 );
and \U$36966 ( \44695_44995 , \44455_44755 , \44468_44768 );
and \U$36967 ( \44696_44996 , \44461_44761 , \44468_44768 );
or \U$36968 ( \44697_44997 , \44694_44994 , \44695_44995 , \44696_44996 );
buf \U$36969 ( \44698_44998 , \44697_44997 );
xor \U$36970 ( \44699_44999 , \44693_44993 , \44698_44998 );
and \U$36971 ( \44700_45000 , \44407_44707 , \44413_44713 );
and \U$36972 ( \44701_45001 , \44407_44707 , \44420_44720 );
and \U$36973 ( \44702_45002 , \44413_44713 , \44420_44720 );
or \U$36974 ( \44703_45003 , \44700_45000 , \44701_45001 , \44702_45002 );
buf \U$36975 ( \44704_45004 , \44703_45003 );
xor \U$36976 ( \44705_45005 , \44699_44999 , \44704_45004 );
buf \U$36977 ( \44706_45006 , \44705_45005 );
xor \U$36978 ( \44707_45007 , \44688_44988 , \44706_45006 );
and \U$36979 ( \44708_45008 , \44379_44679 , \44400_44700 );
and \U$36980 ( \44709_45009 , \44379_44679 , \44422_44722 );
and \U$36981 ( \44710_45010 , \44400_44700 , \44422_44722 );
or \U$36982 ( \44711_45011 , \44708_45008 , \44709_45009 , \44710_45010 );
buf \U$36983 ( \44712_45012 , \44711_45011 );
xor \U$36984 ( \44713_45013 , \44707_45007 , \44712_45012 );
buf \U$36985 ( \44714_45014 , \44713_45013 );
xor \U$36986 ( \44715_45015 , \44683_44983 , \44714_45014 );
buf \U$36987 ( \44716_45016 , \44715_45015 );
xor \U$36988 ( \44717_45017 , \44672_44972 , \44716_45016 );
xor \U$36989 ( \44718_45018 , \44537_44837 , \44717_45017 );
and \U$36990 ( \44719_45019 , \44347_44647 , \44482_44782 );
and \U$36991 ( \44720_45020 , \44347_44647 , \44527_44827 );
and \U$36992 ( \44721_45021 , \44482_44782 , \44527_44827 );
or \U$36993 ( \44722_45022 , \44719_45019 , \44720_45020 , \44721_45021 );
and \U$36994 ( \44723_45023 , \44718_45018 , \44722_45022 );
and \U$36996 ( \44724_45024 , \44536_44836 , \44717_45017 );
or \U$36998 ( \44725_45025 , 1'b0 , \44724_45024 , 1'b0 );
xor \U$36999 ( \44726_45026 , \44723_45023 , \44725_45025 );
and \U$37001 ( \44727_45027 , \44529_44829 , \44535_44835 );
and \U$37002 ( \44728_45028 , \44531_44831 , \44535_44835 );
or \U$37003 ( \44729_45029 , 1'b0 , \44727_45027 , \44728_45028 );
xor \U$37004 ( \44730_45030 , \44726_45026 , \44729_45029 );
xor \U$37011 ( \44731_45031 , \44730_45030 , 1'b0 );
and \U$37012 ( \44732_45032 , \44542_44842 , \44671_44971 );
and \U$37013 ( \44733_45033 , \44542_44842 , \44716_45016 );
and \U$37014 ( \44734_45034 , \44671_44971 , \44716_45016 );
or \U$37015 ( \44735_45035 , \44732_45032 , \44733_45033 , \44734_45034 );
xor \U$37016 ( \44736_45036 , \44731_45031 , \44735_45035 );
and \U$37017 ( \44737_45037 , \44677_44977 , \44682_44982 );
and \U$37018 ( \44738_45038 , \44677_44977 , \44714_45014 );
and \U$37019 ( \44739_45039 , \44682_44982 , \44714_45014 );
or \U$37020 ( \44740_45040 , \44737_45037 , \44738_45038 , \44739_45039 );
buf \U$37021 ( \44741_45041 , \44740_45040 );
and \U$37022 ( \44742_45042 , \44602_44902 , \44607_44907 );
and \U$37023 ( \44743_45043 , \44602_44902 , \44669_44969 );
and \U$37024 ( \44744_45044 , \44607_44907 , \44669_44969 );
or \U$37025 ( \44745_45045 , \44742_45042 , \44743_45043 , \44744_45044 );
buf \U$37026 ( \44746_45046 , \44745_45045 );
and \U$37027 ( \44747_45047 , \31989_31636 , \36289_36589_nG9b93 );
and \U$37028 ( \44748_45048 , \31334_31633 , \36686_36986_nG9b90 );
or \U$37029 ( \44749_45049 , \44747_45047 , \44748_45048 );
xor \U$37030 ( \44750_45050 , \31333_31632 , \44749_45049 );
buf \U$37031 ( \44751_45051 , \44750_45050 );
buf \U$37033 ( \44752_45052 , \44751_45051 );
and \U$37034 ( \44753_45053 , \21908_21658 , \40152_40452_nG9b6f );
and \U$37035 ( \44754_45054 , \21356_21655 , \40543_40843_nG9b6c );
or \U$37036 ( \44755_45055 , \44753_45053 , \44754_45054 );
xor \U$37037 ( \44756_45056 , \21355_21654 , \44755_45055 );
buf \U$37038 ( \44757_45057 , \44756_45056 );
buf \U$37040 ( \44758_45058 , \44757_45057 );
xor \U$37041 ( \44759_45059 , \44752_45052 , \44758_45058 );
and \U$37042 ( \44760_45060 , \17437_17297 , \41901_42201_nG9b5d );
and \U$37043 ( \44761_45061 , \16995_17294 , \42133_42433_nG9b5a );
or \U$37044 ( \44762_45062 , \44760_45060 , \44761_45061 );
xor \U$37045 ( \44763_45063 , \16994_17293 , \44762_45062 );
buf \U$37046 ( \44764_45064 , \44763_45063 );
buf \U$37048 ( \44765_45065 , \44764_45064 );
xor \U$37049 ( \44766_45066 , \44759_45059 , \44765_45065 );
buf \U$37050 ( \44767_45067 , \44766_45066 );
and \U$37051 ( \44768_45068 , \30670_29853 , \36950_37250_nG9b8d );
and \U$37052 ( \44769_45069 , \29551_29850 , \37307_37607_nG9b8a );
or \U$37053 ( \44770_45070 , \44768_45068 , \44769_45069 );
xor \U$37054 ( \44771_45071 , \29550_29849 , \44770_45070 );
buf \U$37055 ( \44772_45072 , \44771_45071 );
buf \U$37057 ( \44773_45073 , \44772_45072 );
and \U$37058 ( \44774_45074 , \28946_28118 , \37674_37974_nG9b87 );
and \U$37059 ( \44775_45075 , \27816_28115 , \38037_38337_nG9b84 );
or \U$37060 ( \44776_45076 , \44774_45074 , \44775_45075 );
xor \U$37061 ( \44777_45077 , \27815_28114 , \44776_45076 );
buf \U$37062 ( \44778_45078 , \44777_45077 );
buf \U$37064 ( \44779_45079 , \44778_45078 );
xor \U$37065 ( \44780_45080 , \44773_45073 , \44779_45079 );
and \U$37066 ( \44781_45081 , \20353_20155 , \40740_41040_nG9b69 );
and \U$37067 ( \44782_45082 , \19853_20152 , \41081_41381_nG9b66 );
or \U$37068 ( \44783_45083 , \44781_45081 , \44782_45082 );
xor \U$37069 ( \44784_45084 , \19852_20151 , \44783_45083 );
buf \U$37070 ( \44785_45085 , \44784_45084 );
buf \U$37072 ( \44786_45086 , \44785_45085 );
xor \U$37073 ( \44787_45087 , \44780_45080 , \44786_45086 );
buf \U$37074 ( \44788_45088 , \44787_45087 );
xor \U$37075 ( \44789_45089 , \44767_45067 , \44788_45088 );
and \U$37076 ( \44790_45090 , \14710_14631 , \42879_43179_nG9b51 );
or \U$37078 ( \44791_45091 , \44790_45090 , 1'b0 );
xor \U$37079 ( \44792_45092 , \14328_14627 , \44791_45091 );
buf \U$37080 ( \44793_45093 , \44792_45092 );
buf \U$37082 ( \44794_45094 , \44793_45093 );
and \U$37084 ( \44795_45095 , \32617_32916 , \35872_36172_nG9b96 );
or \U$37085 ( \44796_45096 , 1'b0 , \44795_45095 );
xor \U$37086 ( \44797_45097 , 1'b0 , \44796_45096 );
buf \U$37087 ( \44798_45098 , \44797_45097 );
buf \U$37088 ( \44799_45099 , \44798_45098 );
not \U$37089 ( \44800_45100 , \44799_45099 );
xor \U$37090 ( \44801_45101 , \44794_45094 , \44800_45100 );
and \U$37091 ( \44802_45102 , \23495_23201 , \39663_39963_nG9b75 );
and \U$37092 ( \44803_45103 , \22899_23198 , \39904_40204_nG9b72 );
or \U$37093 ( \44804_45104 , \44802_45102 , \44803_45103 );
xor \U$37094 ( \44805_45105 , \22898_23197 , \44804_45104 );
buf \U$37095 ( \44806_45106 , \44805_45105 );
buf \U$37097 ( \44807_45107 , \44806_45106 );
xor \U$37098 ( \44808_45108 , \44801_45101 , \44807_45107 );
buf \U$37099 ( \44809_45109 , \44808_45108 );
xor \U$37100 ( \44810_45110 , \44789_45089 , \44809_45109 );
buf \U$37101 ( \44811_45111 , \44810_45110 );
and \U$37102 ( \44812_45112 , \44568_44868 , \44573_44873 );
and \U$37103 ( \44813_45113 , \44568_44868 , \44592_44892 );
and \U$37104 ( \44814_45114 , \44573_44873 , \44592_44892 );
or \U$37105 ( \44815_45115 , \44812_45112 , \44813_45113 , \44814_45114 );
buf \U$37106 ( \44816_45116 , \44815_45115 );
xor \U$37107 ( \44817_45117 , \44811_45111 , \44816_45116 );
and \U$37108 ( \44818_45118 , \44630_44930 , \44636_44936 );
and \U$37109 ( \44819_45119 , \44630_44930 , \44643_44943 );
and \U$37110 ( \44820_45120 , \44636_44936 , \44643_44943 );
or \U$37111 ( \44821_45121 , \44818_45118 , \44819_45119 , \44820_45120 );
buf \U$37112 ( \44822_45122 , \44821_45121 );
and \U$37113 ( \44823_45123 , \44580_44880 , \44584_44884 );
and \U$37114 ( \44824_45124 , \44580_44880 , \44590_44890 );
and \U$37115 ( \44825_45125 , \44584_44884 , \44590_44890 );
or \U$37116 ( \44826_45126 , \44823_45123 , \44824_45124 , \44825_45125 );
buf \U$37117 ( \44827_45127 , \44826_45126 );
xor \U$37118 ( \44828_45128 , \44822_45122 , \44827_45127 );
and \U$37119 ( \44829_45129 , \44652_44952 , \44658_44958 );
and \U$37120 ( \44830_45130 , \44652_44952 , \44665_44965 );
and \U$37121 ( \44831_45131 , \44658_44958 , \44665_44965 );
or \U$37122 ( \44832_45132 , \44829_45129 , \44830_45130 , \44831_45131 );
buf \U$37123 ( \44833_45133 , \44832_45132 );
xor \U$37124 ( \44834_45134 , \44828_45128 , \44833_45133 );
buf \U$37125 ( \44835_45135 , \44834_45134 );
xor \U$37126 ( \44836_45136 , \44817_45117 , \44835_45135 );
buf \U$37127 ( \44837_45137 , \44836_45136 );
xor \U$37128 ( \44838_45138 , \44746_45046 , \44837_45137 );
and \U$37129 ( \44839_45139 , \44688_44988 , \44706_45006 );
and \U$37130 ( \44840_45140 , \44688_44988 , \44712_45012 );
and \U$37131 ( \44841_45141 , \44706_45006 , \44712_45012 );
or \U$37132 ( \44842_45142 , \44839_45139 , \44840_45140 , \44841_45141 );
buf \U$37133 ( \44843_45143 , \44842_45142 );
xor \U$37134 ( \44844_45144 , \44838_45138 , \44843_45143 );
buf \U$37135 ( \44845_45145 , \44844_45144 );
xor \U$37136 ( \44846_45146 , \44741_45041 , \44845_45145 );
and \U$37137 ( \44847_45147 , \44547_44847 , \44594_44894 );
and \U$37138 ( \44848_45148 , \44547_44847 , \44600_44900 );
and \U$37139 ( \44849_45149 , \44594_44894 , \44600_44900 );
or \U$37140 ( \44850_45150 , \44847_45147 , \44848_45148 , \44849_45149 );
buf \U$37141 ( \44851_45151 , \44850_45150 );
and \U$37142 ( \44852_45152 , \44553_44853 , \44559_44859 );
and \U$37143 ( \44853_45153 , \44553_44853 , \44566_44866 );
and \U$37144 ( \44854_45154 , \44559_44859 , \44566_44866 );
or \U$37145 ( \44855_45155 , \44852_45152 , \44853_45153 , \44854_45154 );
buf \U$37146 ( \44856_45156 , \44855_45155 );
and \U$37147 ( \44857_45157 , \44614_44914 , \44620_44920 );
and \U$37148 ( \44858_45158 , \44614_44914 , \44627_44927 );
and \U$37149 ( \44859_45159 , \44620_44920 , \44627_44927 );
or \U$37150 ( \44860_45160 , \44857_45157 , \44858_45158 , \44859_45159 );
buf \U$37151 ( \44861_45161 , \44860_45160 );
xor \U$37152 ( \44862_45162 , \44856_45156 , \44861_45161 );
and \U$37153 ( \44863_45163 , \16405_15940 , \42466_42766_nG9b57 );
and \U$37154 ( \44864_45164 , \15638_15937 , \42548_42848_nG9b54 );
or \U$37155 ( \44865_45165 , \44863_45163 , \44864_45164 );
xor \U$37156 ( \44866_45166 , \15637_15936 , \44865_45165 );
buf \U$37157 ( \44867_45167 , \44866_45166 );
buf \U$37159 ( \44868_45168 , \44867_45167 );
xor \U$37160 ( \44869_45169 , \44862_45162 , \44868_45168 );
buf \U$37161 ( \44870_45170 , \44869_45169 );
and \U$37162 ( \44871_45171 , \44693_44993 , \44698_44998 );
and \U$37163 ( \44872_45172 , \44693_44993 , \44704_45004 );
and \U$37164 ( \44873_45173 , \44698_44998 , \44704_45004 );
or \U$37165 ( \44874_45174 , \44871_45171 , \44872_45172 , \44873_45173 );
buf \U$37166 ( \44875_45175 , \44874_45174 );
xor \U$37167 ( \44876_45176 , \44870_45170 , \44875_45175 );
and \U$37168 ( \44877_45177 , \27141_26431 , \38363_38663_nG9b81 );
and \U$37169 ( \44878_45178 , \26129_26428 , \38668_38968_nG9b7e );
or \U$37170 ( \44879_45179 , \44877_45177 , \44878_45178 );
xor \U$37171 ( \44880_45180 , \26128_26427 , \44879_45179 );
buf \U$37172 ( \44881_45181 , \44880_45180 );
buf \U$37174 ( \44882_45182 , \44881_45181 );
and \U$37175 ( \44883_45183 , \25044_24792 , \39034_39334_nG9b7b );
and \U$37176 ( \44884_45184 , \24490_24789 , \39291_39591_nG9b78 );
or \U$37177 ( \44885_45185 , \44883_45183 , \44884_45184 );
xor \U$37178 ( \44886_45186 , \24489_24788 , \44885_45185 );
buf \U$37179 ( \44887_45187 , \44886_45186 );
buf \U$37181 ( \44888_45188 , \44887_45187 );
xor \U$37182 ( \44889_45189 , \44882_45182 , \44888_45188 );
and \U$37183 ( \44890_45190 , \18908_18702 , \41385_41685_nG9b63 );
and \U$37184 ( \44891_45191 , \18400_18699 , \41663_41963_nG9b60 );
or \U$37185 ( \44892_45192 , \44890_45190 , \44891_45191 );
xor \U$37186 ( \44893_45193 , \18399_18698 , \44892_45192 );
buf \U$37187 ( \44894_45194 , \44893_45193 );
buf \U$37189 ( \44895_45195 , \44894_45194 );
xor \U$37190 ( \44896_45196 , \44889_45189 , \44895_45195 );
buf \U$37191 ( \44897_45197 , \44896_45196 );
xor \U$37192 ( \44898_45198 , \44876_45176 , \44897_45197 );
buf \U$37193 ( \44899_45199 , \44898_45198 );
xor \U$37194 ( \44900_45200 , \44851_45151 , \44899_45199 );
and \U$37195 ( \44901_45201 , \44629_44929 , \44645_44945 );
and \U$37196 ( \44902_45202 , \44629_44929 , \44667_44967 );
and \U$37197 ( \44903_45203 , \44645_44945 , \44667_44967 );
or \U$37198 ( \44904_45204 , \44901_45201 , \44902_45202 , \44903_45203 );
buf \U$37199 ( \44905_45205 , \44904_45204 );
xor \U$37200 ( \44906_45206 , \44900_45200 , \44905_45205 );
buf \U$37201 ( \44907_45207 , \44906_45206 );
xor \U$37202 ( \44908_45208 , \44846_45146 , \44907_45207 );
and \U$37203 ( \44909_45209 , \44736_45036 , \44908_45208 );
and \U$37205 ( \44910_45210 , \44730_45030 , \44735_45035 );
or \U$37207 ( \44911_45211 , 1'b0 , \44910_45210 , 1'b0 );
xor \U$37208 ( \44912_45212 , \44909_45209 , \44911_45211 );
and \U$37210 ( \44913_45213 , \44723_45023 , \44729_45029 );
and \U$37211 ( \44914_45214 , \44725_45025 , \44729_45029 );
or \U$37212 ( \44915_45215 , 1'b0 , \44913_45213 , \44914_45214 );
xor \U$37213 ( \44916_45216 , \44912_45212 , \44915_45215 );
xor \U$37220 ( \44917_45217 , \44916_45216 , 1'b0 );
and \U$37221 ( \44918_45218 , \44741_45041 , \44845_45145 );
and \U$37222 ( \44919_45219 , \44741_45041 , \44907_45207 );
and \U$37223 ( \44920_45220 , \44845_45145 , \44907_45207 );
or \U$37224 ( \44921_45221 , \44918_45218 , \44919_45219 , \44920_45220 );
xor \U$37225 ( \44922_45222 , \44917_45217 , \44921_45221 );
and \U$37226 ( \44923_45223 , \44767_45067 , \44788_45088 );
and \U$37227 ( \44924_45224 , \44767_45067 , \44809_45109 );
and \U$37228 ( \44925_45225 , \44788_45088 , \44809_45109 );
or \U$37229 ( \44926_45226 , \44923_45223 , \44924_45224 , \44925_45225 );
buf \U$37230 ( \44927_45227 , \44926_45226 );
and \U$37231 ( \44928_45228 , \44752_45052 , \44758_45058 );
and \U$37232 ( \44929_45229 , \44752_45052 , \44765_45065 );
and \U$37233 ( \44930_45230 , \44758_45058 , \44765_45065 );
or \U$37234 ( \44931_45231 , \44928_45228 , \44929_45229 , \44930_45230 );
buf \U$37235 ( \44932_45232 , \44931_45231 );
and \U$37236 ( \44933_45233 , \44794_45094 , \44800_45100 );
and \U$37237 ( \44934_45234 , \44794_45094 , \44807_45107 );
and \U$37238 ( \44935_45235 , \44800_45100 , \44807_45107 );
or \U$37239 ( \44936_45236 , \44933_45233 , \44934_45234 , \44935_45235 );
buf \U$37240 ( \44937_45237 , \44936_45236 );
xor \U$37241 ( \44938_45238 , \44932_45232 , \44937_45237 );
and \U$37242 ( \44939_45239 , \44882_45182 , \44888_45188 );
and \U$37243 ( \44940_45240 , \44882_45182 , \44895_45195 );
and \U$37244 ( \44941_45241 , \44888_45188 , \44895_45195 );
or \U$37245 ( \44942_45242 , \44939_45239 , \44940_45240 , \44941_45241 );
buf \U$37246 ( \44943_45243 , \44942_45242 );
xor \U$37247 ( \44944_45244 , \44938_45238 , \44943_45243 );
buf \U$37248 ( \44945_45245 , \44944_45244 );
xor \U$37249 ( \44946_45246 , \44927_45227 , \44945_45245 );
and \U$37250 ( \44947_45247 , \44822_45122 , \44827_45127 );
and \U$37251 ( \44948_45248 , \44822_45122 , \44833_45133 );
and \U$37252 ( \44949_45249 , \44827_45127 , \44833_45133 );
or \U$37253 ( \44950_45250 , \44947_45247 , \44948_45248 , \44949_45249 );
buf \U$37254 ( \44951_45251 , \44950_45250 );
xor \U$37255 ( \44952_45252 , \44946_45246 , \44951_45251 );
buf \U$37256 ( \44953_45253 , \44952_45252 );
and \U$37257 ( \44954_45254 , \44811_45111 , \44816_45116 );
and \U$37258 ( \44955_45255 , \44811_45111 , \44835_45135 );
and \U$37259 ( \44956_45256 , \44816_45116 , \44835_45135 );
or \U$37260 ( \44957_45257 , \44954_45254 , \44955_45255 , \44956_45256 );
buf \U$37261 ( \44958_45258 , \44957_45257 );
xor \U$37262 ( \44959_45259 , \44953_45253 , \44958_45258 );
and \U$37263 ( \44960_45260 , \44851_45151 , \44899_45199 );
and \U$37264 ( \44961_45261 , \44851_45151 , \44905_45205 );
and \U$37265 ( \44962_45262 , \44899_45199 , \44905_45205 );
or \U$37266 ( \44963_45263 , \44960_45260 , \44961_45261 , \44962_45262 );
buf \U$37267 ( \44964_45264 , \44963_45263 );
xor \U$37268 ( \44965_45265 , \44959_45259 , \44964_45264 );
buf \U$37269 ( \44966_45266 , \44965_45265 );
and \U$37270 ( \44967_45267 , \44746_45046 , \44837_45137 );
and \U$37271 ( \44968_45268 , \44746_45046 , \44843_45143 );
and \U$37272 ( \44969_45269 , \44837_45137 , \44843_45143 );
or \U$37273 ( \44970_45270 , \44967_45267 , \44968_45268 , \44969_45269 );
buf \U$37274 ( \44971_45271 , \44970_45270 );
xor \U$37275 ( \44972_45272 , \44966_45266 , \44971_45271 );
and \U$37276 ( \44973_45273 , \44773_45073 , \44779_45079 );
and \U$37277 ( \44974_45274 , \44773_45073 , \44786_45086 );
and \U$37278 ( \44975_45275 , \44779_45079 , \44786_45086 );
or \U$37279 ( \44976_45276 , \44973_45273 , \44974_45274 , \44975_45275 );
buf \U$37280 ( \44977_45277 , \44976_45276 );
buf \U$37281 ( \44978_45278 , \44799_45099 );
xor \U$37282 ( \44979_45279 , \44977_45277 , \44978_45278 );
and \U$37283 ( \44980_45280 , \17437_17297 , \42133_42433_nG9b5a );
and \U$37284 ( \44981_45281 , \16995_17294 , \42466_42766_nG9b57 );
or \U$37285 ( \44982_45282 , \44980_45280 , \44981_45281 );
xor \U$37286 ( \44983_45283 , \16994_17293 , \44982_45282 );
buf \U$37287 ( \44984_45284 , \44983_45283 );
buf \U$37289 ( \44985_45285 , \44984_45284 );
xor \U$37290 ( \44986_45286 , \44979_45279 , \44985_45285 );
buf \U$37291 ( \44987_45287 , \44986_45286 );
and \U$37292 ( \44988_45288 , \44856_45156 , \44861_45161 );
and \U$37293 ( \44989_45289 , \44856_45156 , \44868_45168 );
and \U$37294 ( \44990_45290 , \44861_45161 , \44868_45168 );
or \U$37295 ( \44991_45291 , \44988_45288 , \44989_45289 , \44990_45290 );
buf \U$37296 ( \44992_45292 , \44991_45291 );
xor \U$37297 ( \44993_45293 , \44987_45287 , \44992_45292 );
and \U$37299 ( \44994_45294 , \32617_32916 , \36289_36589_nG9b93 );
or \U$37300 ( \44995_45295 , 1'b0 , \44994_45294 );
xor \U$37301 ( \44996_45296 , 1'b0 , \44995_45295 );
buf \U$37302 ( \44997_45297 , \44996_45296 );
buf \U$37304 ( \44998_45298 , \44997_45297 );
and \U$37305 ( \44999_45299 , \31989_31636 , \36686_36986_nG9b90 );
and \U$37306 ( \45000_45300 , \31334_31633 , \36950_37250_nG9b8d );
or \U$37307 ( \45001_45301 , \44999_45299 , \45000_45300 );
xor \U$37308 ( \45002_45302 , \31333_31632 , \45001_45301 );
buf \U$37309 ( \45003_45303 , \45002_45302 );
buf \U$37311 ( \45004_45304 , \45003_45303 );
xor \U$37312 ( \45005_45305 , \44998_45298 , \45004_45304 );
and \U$37313 ( \45006_45306 , \23495_23201 , \39904_40204_nG9b72 );
and \U$37314 ( \45007_45307 , \22899_23198 , \40152_40452_nG9b6f );
or \U$37315 ( \45008_45308 , \45006_45306 , \45007_45307 );
xor \U$37316 ( \45009_45309 , \22898_23197 , \45008_45308 );
buf \U$37317 ( \45010_45310 , \45009_45309 );
buf \U$37319 ( \45011_45311 , \45010_45310 );
xor \U$37320 ( \45012_45312 , \45005_45305 , \45011_45311 );
buf \U$37321 ( \45013_45313 , \45012_45312 );
xor \U$37322 ( \45014_45314 , \44993_45293 , \45013_45313 );
buf \U$37323 ( \45015_45315 , \45014_45314 );
and \U$37324 ( \45016_45316 , \44870_45170 , \44875_45175 );
and \U$37325 ( \45017_45317 , \44870_45170 , \44897_45197 );
and \U$37326 ( \45018_45318 , \44875_45175 , \44897_45197 );
or \U$37327 ( \45019_45319 , \45016_45316 , \45017_45317 , \45018_45318 );
buf \U$37328 ( \45020_45320 , \45019_45319 );
xor \U$37329 ( \45021_45321 , \45015_45315 , \45020_45320 );
and \U$37330 ( \45022_45322 , \27141_26431 , \38668_38968_nG9b7e );
and \U$37331 ( \45023_45323 , \26129_26428 , \39034_39334_nG9b7b );
or \U$37332 ( \45024_45324 , \45022_45322 , \45023_45323 );
xor \U$37333 ( \45025_45325 , \26128_26427 , \45024_45324 );
buf \U$37334 ( \45026_45326 , \45025_45325 );
buf \U$37336 ( \45027_45327 , \45026_45326 );
and \U$37337 ( \45028_45328 , \25044_24792 , \39291_39591_nG9b78 );
and \U$37338 ( \45029_45329 , \24490_24789 , \39663_39963_nG9b75 );
or \U$37339 ( \45030_45330 , \45028_45328 , \45029_45329 );
xor \U$37340 ( \45031_45331 , \24489_24788 , \45030_45330 );
buf \U$37341 ( \45032_45332 , \45031_45331 );
buf \U$37343 ( \45033_45333 , \45032_45332 );
xor \U$37344 ( \45034_45334 , \45027_45327 , \45033_45333 );
and \U$37345 ( \45035_45335 , \20353_20155 , \41081_41381_nG9b66 );
and \U$37346 ( \45036_45336 , \19853_20152 , \41385_41685_nG9b63 );
or \U$37347 ( \45037_45337 , \45035_45335 , \45036_45336 );
xor \U$37348 ( \45038_45338 , \19852_20151 , \45037_45337 );
buf \U$37349 ( \45039_45339 , \45038_45338 );
buf \U$37351 ( \45040_45340 , \45039_45339 );
xor \U$37352 ( \45041_45341 , \45034_45334 , \45040_45340 );
buf \U$37353 ( \45042_45342 , \45041_45341 );
and \U$37354 ( \45043_45343 , \16405_15940 , \42548_42848_nG9b54 );
and \U$37355 ( \45044_45344 , \15638_15937 , \42879_43179_nG9b51 );
or \U$37356 ( \45045_45345 , \45043_45343 , \45044_45344 );
xor \U$37357 ( \45046_45346 , \15637_15936 , \45045_45345 );
buf \U$37358 ( \45047_45347 , \45046_45346 );
buf \U$37360 ( \45048_45348 , \45047_45347 );
xor \U$37364 ( \45049_45349 , \14328_14627 , 1'b0 );
not \U$37365 ( \45050_45350 , \45049_45349 );
buf \U$37366 ( \45051_45351 , \45050_45350 );
buf \U$37368 ( \45052_45352 , \45051_45351 );
xor \U$37369 ( \45053_45353 , \45048_45348 , \45052_45352 );
and \U$37370 ( \45054_45354 , \18908_18702 , \41663_41963_nG9b60 );
and \U$37371 ( \45055_45355 , \18400_18699 , \41901_42201_nG9b5d );
or \U$37372 ( \45056_45356 , \45054_45354 , \45055_45355 );
xor \U$37373 ( \45057_45357 , \18399_18698 , \45056_45356 );
buf \U$37374 ( \45058_45358 , \45057_45357 );
buf \U$37376 ( \45059_45359 , \45058_45358 );
xor \U$37377 ( \45060_45360 , \45053_45353 , \45059_45359 );
buf \U$37378 ( \45061_45361 , \45060_45360 );
xor \U$37379 ( \45062_45362 , \45042_45342 , \45061_45361 );
and \U$37380 ( \45063_45363 , \30670_29853 , \37307_37607_nG9b8a );
and \U$37381 ( \45064_45364 , \29551_29850 , \37674_37974_nG9b87 );
or \U$37382 ( \45065_45365 , \45063_45363 , \45064_45364 );
xor \U$37383 ( \45066_45366 , \29550_29849 , \45065_45365 );
buf \U$37384 ( \45067_45367 , \45066_45366 );
buf \U$37386 ( \45068_45368 , \45067_45367 );
and \U$37387 ( \45069_45369 , \28946_28118 , \38037_38337_nG9b84 );
and \U$37388 ( \45070_45370 , \27816_28115 , \38363_38663_nG9b81 );
or \U$37389 ( \45071_45371 , \45069_45369 , \45070_45370 );
xor \U$37390 ( \45072_45372 , \27815_28114 , \45071_45371 );
buf \U$37391 ( \45073_45373 , \45072_45372 );
buf \U$37393 ( \45074_45374 , \45073_45373 );
xor \U$37394 ( \45075_45375 , \45068_45368 , \45074_45374 );
and \U$37395 ( \45076_45376 , \21908_21658 , \40543_40843_nG9b6c );
and \U$37396 ( \45077_45377 , \21356_21655 , \40740_41040_nG9b69 );
or \U$37397 ( \45078_45378 , \45076_45376 , \45077_45377 );
xor \U$37398 ( \45079_45379 , \21355_21654 , \45078_45378 );
buf \U$37399 ( \45080_45380 , \45079_45379 );
buf \U$37401 ( \45081_45381 , \45080_45380 );
xor \U$37402 ( \45082_45382 , \45075_45375 , \45081_45381 );
buf \U$37403 ( \45083_45383 , \45082_45382 );
xor \U$37404 ( \45084_45384 , \45062_45362 , \45083_45383 );
buf \U$37405 ( \45085_45385 , \45084_45384 );
xor \U$37406 ( \45086_45386 , \45021_45321 , \45085_45385 );
buf \U$37407 ( \45087_45387 , \45086_45386 );
xor \U$37408 ( \45088_45388 , \44972_45272 , \45087_45387 );
and \U$37409 ( \45089_45389 , \44922_45222 , \45088_45388 );
and \U$37411 ( \45090_45390 , \44916_45216 , \44921_45221 );
or \U$37413 ( \45091_45391 , 1'b0 , \45090_45390 , 1'b0 );
xor \U$37414 ( \45092_45392 , \45089_45389 , \45091_45391 );
and \U$37416 ( \45093_45393 , \44909_45209 , \44915_45215 );
and \U$37417 ( \45094_45394 , \44911_45211 , \44915_45215 );
or \U$37418 ( \45095_45395 , 1'b0 , \45093_45393 , \45094_45394 );
xor \U$37419 ( \45096_45396 , \45092_45392 , \45095_45395 );
xor \U$37426 ( \45097_45397 , \45096_45396 , 1'b0 );
and \U$37427 ( \45098_45398 , \44966_45266 , \44971_45271 );
and \U$37428 ( \45099_45399 , \44966_45266 , \45087_45387 );
and \U$37429 ( \45100_45400 , \44971_45271 , \45087_45387 );
or \U$37430 ( \45101_45401 , \45098_45398 , \45099_45399 , \45100_45400 );
xor \U$37431 ( \45102_45402 , \45097_45397 , \45101_45401 );
and \U$37432 ( \45103_45403 , \44977_45277 , \44978_45278 );
and \U$37433 ( \45104_45404 , \44977_45277 , \44985_45285 );
and \U$37434 ( \45105_45405 , \44978_45278 , \44985_45285 );
or \U$37435 ( \45106_45406 , \45103_45403 , \45104_45404 , \45105_45405 );
buf \U$37436 ( \45107_45407 , \45106_45406 );
and \U$37437 ( \45108_45408 , \25044_24792 , \39663_39963_nG9b75 );
and \U$37438 ( \45109_45409 , \24490_24789 , \39904_40204_nG9b72 );
or \U$37439 ( \45110_45410 , \45108_45408 , \45109_45409 );
xor \U$37440 ( \45111_45411 , \24489_24788 , \45110_45410 );
buf \U$37441 ( \45112_45412 , \45111_45411 );
buf \U$37443 ( \45113_45413 , \45112_45412 );
and \U$37444 ( \45114_45414 , \20353_20155 , \41385_41685_nG9b63 );
and \U$37445 ( \45115_45415 , \19853_20152 , \41663_41963_nG9b60 );
or \U$37446 ( \45116_45416 , \45114_45414 , \45115_45415 );
xor \U$37447 ( \45117_45417 , \19852_20151 , \45116_45416 );
buf \U$37448 ( \45118_45418 , \45117_45417 );
buf \U$37449 ( \45119_45419 , \45118_45418 );
not \U$37450 ( \45120_45420 , \45119_45419 );
xor \U$37451 ( \45121_45421 , \45113_45413 , \45120_45420 );
and \U$37452 ( \45122_45422 , \17437_17297 , \42466_42766_nG9b57 );
and \U$37453 ( \45123_45423 , \16995_17294 , \42548_42848_nG9b54 );
or \U$37454 ( \45124_45424 , \45122_45422 , \45123_45423 );
xor \U$37455 ( \45125_45425 , \16994_17293 , \45124_45424 );
buf \U$37456 ( \45126_45426 , \45125_45425 );
buf \U$37458 ( \45127_45427 , \45126_45426 );
xor \U$37459 ( \45128_45428 , \45121_45421 , \45127_45427 );
buf \U$37460 ( \45129_45429 , \45128_45428 );
xor \U$37461 ( \45130_45430 , \45107_45407 , \45129_45429 );
and \U$37462 ( \45131_45431 , \28946_28118 , \38363_38663_nG9b81 );
and \U$37463 ( \45132_45432 , \27816_28115 , \38668_38968_nG9b7e );
or \U$37464 ( \45133_45433 , \45131_45431 , \45132_45432 );
xor \U$37465 ( \45134_45434 , \27815_28114 , \45133_45433 );
buf \U$37466 ( \45135_45435 , \45134_45434 );
buf \U$37468 ( \45136_45436 , \45135_45435 );
and \U$37469 ( \45137_45437 , \27141_26431 , \39034_39334_nG9b7b );
and \U$37470 ( \45138_45438 , \26129_26428 , \39291_39591_nG9b78 );
or \U$37471 ( \45139_45439 , \45137_45437 , \45138_45438 );
xor \U$37472 ( \45140_45440 , \26128_26427 , \45139_45439 );
buf \U$37473 ( \45141_45441 , \45140_45440 );
buf \U$37475 ( \45142_45442 , \45141_45441 );
xor \U$37476 ( \45143_45443 , \45136_45436 , \45142_45442 );
and \U$37477 ( \45144_45444 , \21908_21658 , \40740_41040_nG9b69 );
and \U$37478 ( \45145_45445 , \21356_21655 , \41081_41381_nG9b66 );
or \U$37479 ( \45146_45446 , \45144_45444 , \45145_45445 );
xor \U$37480 ( \45147_45447 , \21355_21654 , \45146_45446 );
buf \U$37481 ( \45148_45448 , \45147_45447 );
buf \U$37483 ( \45149_45449 , \45148_45448 );
xor \U$37484 ( \45150_45450 , \45143_45443 , \45149_45449 );
buf \U$37485 ( \45151_45451 , \45150_45450 );
xor \U$37486 ( \45152_45452 , \45130_45430 , \45151_45451 );
buf \U$37487 ( \45153_45453 , \45152_45452 );
and \U$37488 ( \45154_45454 , \44987_45287 , \44992_45292 );
and \U$37489 ( \45155_45455 , \44987_45287 , \45013_45313 );
and \U$37490 ( \45156_45456 , \44992_45292 , \45013_45313 );
or \U$37491 ( \45157_45457 , \45154_45454 , \45155_45455 , \45156_45456 );
buf \U$37492 ( \45158_45458 , \45157_45457 );
xor \U$37493 ( \45159_45459 , \45153_45453 , \45158_45458 );
and \U$37494 ( \45160_45460 , \16405_15940 , \42879_43179_nG9b51 );
or \U$37496 ( \45161_45461 , \45160_45460 , 1'b0 );
xor \U$37497 ( \45162_45462 , \15637_15936 , \45161_45461 );
buf \U$37498 ( \45163_45463 , \45162_45462 );
buf \U$37500 ( \45164_45464 , \45163_45463 );
and \U$37501 ( \45165_45465 , \31989_31636 , \36950_37250_nG9b8d );
and \U$37502 ( \45166_45466 , \31334_31633 , \37307_37607_nG9b8a );
or \U$37503 ( \45167_45467 , \45165_45465 , \45166_45466 );
xor \U$37504 ( \45168_45468 , \31333_31632 , \45167_45467 );
buf \U$37505 ( \45169_45469 , \45168_45468 );
buf \U$37507 ( \45170_45470 , \45169_45469 );
xor \U$37508 ( \45171_45471 , \45164_45464 , \45170_45470 );
and \U$37509 ( \45172_45472 , \30670_29853 , \37674_37974_nG9b87 );
and \U$37510 ( \45173_45473 , \29551_29850 , \38037_38337_nG9b84 );
or \U$37511 ( \45174_45474 , \45172_45472 , \45173_45473 );
xor \U$37512 ( \45175_45475 , \29550_29849 , \45174_45474 );
buf \U$37513 ( \45176_45476 , \45175_45475 );
buf \U$37515 ( \45177_45477 , \45176_45476 );
xor \U$37516 ( \45178_45478 , \45171_45471 , \45177_45477 );
buf \U$37517 ( \45179_45479 , \45178_45478 );
and \U$37519 ( \45180_45480 , \32617_32916 , \36686_36986_nG9b90 );
or \U$37520 ( \45181_45481 , 1'b0 , \45180_45480 );
xor \U$37521 ( \45182_45482 , 1'b0 , \45181_45481 );
buf \U$37522 ( \45183_45483 , \45182_45482 );
buf \U$37524 ( \45184_45484 , \45183_45483 );
and \U$37525 ( \45185_45485 , \23495_23201 , \40152_40452_nG9b6f );
and \U$37526 ( \45186_45486 , \22899_23198 , \40543_40843_nG9b6c );
or \U$37527 ( \45187_45487 , \45185_45485 , \45186_45486 );
xor \U$37528 ( \45188_45488 , \22898_23197 , \45187_45487 );
buf \U$37529 ( \45189_45489 , \45188_45488 );
buf \U$37531 ( \45190_45490 , \45189_45489 );
xor \U$37532 ( \45191_45491 , \45184_45484 , \45190_45490 );
and \U$37533 ( \45192_45492 , \18908_18702 , \41901_42201_nG9b5d );
and \U$37534 ( \45193_45493 , \18400_18699 , \42133_42433_nG9b5a );
or \U$37535 ( \45194_45494 , \45192_45492 , \45193_45493 );
xor \U$37536 ( \45195_45495 , \18399_18698 , \45194_45494 );
buf \U$37537 ( \45196_45496 , \45195_45495 );
buf \U$37539 ( \45197_45497 , \45196_45496 );
xor \U$37540 ( \45198_45498 , \45191_45491 , \45197_45497 );
buf \U$37541 ( \45199_45499 , \45198_45498 );
xor \U$37542 ( \45200_45500 , \45179_45479 , \45199_45499 );
and \U$37543 ( \45201_45501 , \45027_45327 , \45033_45333 );
and \U$37544 ( \45202_45502 , \45027_45327 , \45040_45340 );
and \U$37545 ( \45203_45503 , \45033_45333 , \45040_45340 );
or \U$37546 ( \45204_45504 , \45201_45501 , \45202_45502 , \45203_45503 );
buf \U$37547 ( \45205_45505 , \45204_45504 );
xor \U$37548 ( \45206_45506 , \45200_45500 , \45205_45505 );
buf \U$37549 ( \45207_45507 , \45206_45506 );
xor \U$37550 ( \45208_45508 , \45159_45459 , \45207_45507 );
buf \U$37551 ( \45209_45509 , \45208_45508 );
and \U$37552 ( \45210_45510 , \45042_45342 , \45061_45361 );
and \U$37553 ( \45211_45511 , \45042_45342 , \45083_45383 );
and \U$37554 ( \45212_45512 , \45061_45361 , \45083_45383 );
or \U$37555 ( \45213_45513 , \45210_45510 , \45211_45511 , \45212_45512 );
buf \U$37556 ( \45214_45514 , \45213_45513 );
and \U$37557 ( \45215_45515 , \45048_45348 , \45052_45352 );
and \U$37558 ( \45216_45516 , \45048_45348 , \45059_45359 );
and \U$37559 ( \45217_45517 , \45052_45352 , \45059_45359 );
or \U$37560 ( \45218_45518 , \45215_45515 , \45216_45516 , \45217_45517 );
buf \U$37561 ( \45219_45519 , \45218_45518 );
and \U$37562 ( \45220_45520 , \45068_45368 , \45074_45374 );
and \U$37563 ( \45221_45521 , \45068_45368 , \45081_45381 );
and \U$37564 ( \45222_45522 , \45074_45374 , \45081_45381 );
or \U$37565 ( \45223_45523 , \45220_45520 , \45221_45521 , \45222_45522 );
buf \U$37566 ( \45224_45524 , \45223_45523 );
xor \U$37567 ( \45225_45525 , \45219_45519 , \45224_45524 );
and \U$37568 ( \45226_45526 , \44998_45298 , \45004_45304 );
and \U$37569 ( \45227_45527 , \44998_45298 , \45011_45311 );
and \U$37570 ( \45228_45528 , \45004_45304 , \45011_45311 );
or \U$37571 ( \45229_45529 , \45226_45526 , \45227_45527 , \45228_45528 );
buf \U$37572 ( \45230_45530 , \45229_45529 );
xor \U$37573 ( \45231_45531 , \45225_45525 , \45230_45530 );
buf \U$37574 ( \45232_45532 , \45231_45531 );
xor \U$37575 ( \45233_45533 , \45214_45514 , \45232_45532 );
and \U$37576 ( \45234_45534 , \44932_45232 , \44937_45237 );
and \U$37577 ( \45235_45535 , \44932_45232 , \44943_45243 );
and \U$37578 ( \45236_45536 , \44937_45237 , \44943_45243 );
or \U$37579 ( \45237_45537 , \45234_45534 , \45235_45535 , \45236_45536 );
buf \U$37580 ( \45238_45538 , \45237_45537 );
xor \U$37581 ( \45239_45539 , \45233_45533 , \45238_45538 );
buf \U$37582 ( \45240_45540 , \45239_45539 );
xor \U$37583 ( \45241_45541 , \45209_45509 , \45240_45540 );
and \U$37584 ( \45242_45542 , \44927_45227 , \44945_45245 );
and \U$37585 ( \45243_45543 , \44927_45227 , \44951_45251 );
and \U$37586 ( \45244_45544 , \44945_45245 , \44951_45251 );
or \U$37587 ( \45245_45545 , \45242_45542 , \45243_45543 , \45244_45544 );
buf \U$37588 ( \45246_45546 , \45245_45545 );
xor \U$37589 ( \45247_45547 , \45241_45541 , \45246_45546 );
buf \U$37590 ( \45248_45548 , \45247_45547 );
and \U$37591 ( \45249_45549 , \44953_45253 , \44958_45258 );
and \U$37592 ( \45250_45550 , \44953_45253 , \44964_45264 );
and \U$37593 ( \45251_45551 , \44958_45258 , \44964_45264 );
or \U$37594 ( \45252_45552 , \45249_45549 , \45250_45550 , \45251_45551 );
buf \U$37595 ( \45253_45553 , \45252_45552 );
xor \U$37596 ( \45254_45554 , \45248_45548 , \45253_45553 );
and \U$37597 ( \45255_45555 , \45015_45315 , \45020_45320 );
and \U$37598 ( \45256_45556 , \45015_45315 , \45085_45385 );
and \U$37599 ( \45257_45557 , \45020_45320 , \45085_45385 );
or \U$37600 ( \45258_45558 , \45255_45555 , \45256_45556 , \45257_45557 );
buf \U$37601 ( \45259_45559 , \45258_45558 );
xor \U$37602 ( \45260_45560 , \45254_45554 , \45259_45559 );
and \U$37603 ( \45261_45561 , \45102_45402 , \45260_45560 );
and \U$37605 ( \45262_45562 , \45096_45396 , \45101_45401 );
or \U$37607 ( \45263_45563 , 1'b0 , \45262_45562 , 1'b0 );
xor \U$37608 ( \45264_45564 , \45261_45561 , \45263_45563 );
and \U$37610 ( \45265_45565 , \45089_45389 , \45095_45395 );
and \U$37611 ( \45266_45566 , \45091_45391 , \45095_45395 );
or \U$37612 ( \45267_45567 , 1'b0 , \45265_45565 , \45266_45566 );
xor \U$37613 ( \45268_45568 , \45264_45564 , \45267_45567 );
xor \U$37620 ( \45269_45569 , \45268_45568 , 1'b0 );
and \U$37621 ( \45270_45570 , \45248_45548 , \45253_45553 );
and \U$37622 ( \45271_45571 , \45248_45548 , \45259_45559 );
and \U$37623 ( \45272_45572 , \45253_45553 , \45259_45559 );
or \U$37624 ( \45273_45573 , \45270_45570 , \45271_45571 , \45272_45572 );
xor \U$37625 ( \45274_45574 , \45269_45569 , \45273_45573 );
and \U$37626 ( \45275_45575 , \45107_45407 , \45129_45429 );
and \U$37627 ( \45276_45576 , \45107_45407 , \45151_45451 );
and \U$37628 ( \45277_45577 , \45129_45429 , \45151_45451 );
or \U$37629 ( \45278_45578 , \45275_45575 , \45276_45576 , \45277_45577 );
buf \U$37630 ( \45279_45579 , \45278_45578 );
and \U$37631 ( \45280_45580 , \45113_45413 , \45120_45420 );
and \U$37632 ( \45281_45581 , \45113_45413 , \45127_45427 );
and \U$37633 ( \45282_45582 , \45120_45420 , \45127_45427 );
or \U$37634 ( \45283_45583 , \45280_45580 , \45281_45581 , \45282_45582 );
buf \U$37635 ( \45284_45584 , \45283_45583 );
and \U$37636 ( \45285_45585 , \28946_28118 , \38668_38968_nG9b7e );
and \U$37637 ( \45286_45586 , \27816_28115 , \39034_39334_nG9b7b );
or \U$37638 ( \45287_45587 , \45285_45585 , \45286_45586 );
xor \U$37639 ( \45288_45588 , \27815_28114 , \45287_45587 );
buf \U$37640 ( \45289_45589 , \45288_45588 );
buf \U$37642 ( \45290_45590 , \45289_45589 );
and \U$37643 ( \45291_45591 , \27141_26431 , \39291_39591_nG9b78 );
and \U$37644 ( \45292_45592 , \26129_26428 , \39663_39963_nG9b75 );
or \U$37645 ( \45293_45593 , \45291_45591 , \45292_45592 );
xor \U$37646 ( \45294_45594 , \26128_26427 , \45293_45593 );
buf \U$37647 ( \45295_45595 , \45294_45594 );
buf \U$37649 ( \45296_45596 , \45295_45595 );
xor \U$37650 ( \45297_45597 , \45290_45590 , \45296_45596 );
and \U$37651 ( \45298_45598 , \21908_21658 , \41081_41381_nG9b66 );
and \U$37652 ( \45299_45599 , \21356_21655 , \41385_41685_nG9b63 );
or \U$37653 ( \45300_45600 , \45298_45598 , \45299_45599 );
xor \U$37654 ( \45301_45601 , \21355_21654 , \45300_45600 );
buf \U$37655 ( \45302_45602 , \45301_45601 );
buf \U$37657 ( \45303_45603 , \45302_45602 );
xor \U$37658 ( \45304_45604 , \45297_45597 , \45303_45603 );
buf \U$37659 ( \45305_45605 , \45304_45604 );
xor \U$37660 ( \45306_45606 , \45284_45584 , \45305_45605 );
and \U$37661 ( \45307_45607 , \17437_17297 , \42548_42848_nG9b54 );
and \U$37662 ( \45308_45608 , \16995_17294 , \42879_43179_nG9b51 );
or \U$37663 ( \45309_45609 , \45307_45607 , \45308_45608 );
xor \U$37664 ( \45310_45610 , \16994_17293 , \45309_45609 );
buf \U$37665 ( \45311_45611 , \45310_45610 );
buf \U$37667 ( \45312_45612 , \45311_45611 );
xor \U$37671 ( \45313_45613 , \15637_15936 , 1'b0 );
not \U$37672 ( \45314_45614 , \45313_45613 );
buf \U$37673 ( \45315_45615 , \45314_45614 );
buf \U$37675 ( \45316_45616 , \45315_45615 );
xor \U$37676 ( \45317_45617 , \45312_45612 , \45316_45616 );
and \U$37677 ( \45318_45618 , \20353_20155 , \41663_41963_nG9b60 );
and \U$37678 ( \45319_45619 , \19853_20152 , \41901_42201_nG9b5d );
or \U$37679 ( \45320_45620 , \45318_45618 , \45319_45619 );
xor \U$37680 ( \45321_45621 , \19852_20151 , \45320_45620 );
buf \U$37681 ( \45322_45622 , \45321_45621 );
buf \U$37683 ( \45323_45623 , \45322_45622 );
xor \U$37684 ( \45324_45624 , \45317_45617 , \45323_45623 );
buf \U$37685 ( \45325_45625 , \45324_45624 );
xor \U$37686 ( \45326_45626 , \45306_45606 , \45325_45625 );
buf \U$37687 ( \45327_45627 , \45326_45626 );
xor \U$37688 ( \45328_45628 , \45279_45579 , \45327_45627 );
and \U$37690 ( \45329_45629 , \32617_32916 , \36950_37250_nG9b8d );
or \U$37691 ( \45330_45630 , 1'b0 , \45329_45629 );
xor \U$37692 ( \45331_45631 , 1'b0 , \45330_45630 );
buf \U$37693 ( \45332_45632 , \45331_45631 );
buf \U$37695 ( \45333_45633 , \45332_45632 );
and \U$37696 ( \45334_45634 , \25044_24792 , \39904_40204_nG9b72 );
and \U$37697 ( \45335_45635 , \24490_24789 , \40152_40452_nG9b6f );
or \U$37698 ( \45336_45636 , \45334_45634 , \45335_45635 );
xor \U$37699 ( \45337_45637 , \24489_24788 , \45336_45636 );
buf \U$37700 ( \45338_45638 , \45337_45637 );
buf \U$37702 ( \45339_45639 , \45338_45638 );
xor \U$37703 ( \45340_45640 , \45333_45633 , \45339_45639 );
and \U$37704 ( \45341_45641 , \18908_18702 , \42133_42433_nG9b5a );
and \U$37705 ( \45342_45642 , \18400_18699 , \42466_42766_nG9b57 );
or \U$37706 ( \45343_45643 , \45341_45641 , \45342_45642 );
xor \U$37707 ( \45344_45644 , \18399_18698 , \45343_45643 );
buf \U$37708 ( \45345_45645 , \45344_45644 );
buf \U$37710 ( \45346_45646 , \45345_45645 );
xor \U$37711 ( \45347_45647 , \45340_45640 , \45346_45646 );
buf \U$37712 ( \45348_45648 , \45347_45647 );
and \U$37713 ( \45349_45649 , \31989_31636 , \37307_37607_nG9b8a );
and \U$37714 ( \45350_45650 , \31334_31633 , \37674_37974_nG9b87 );
or \U$37715 ( \45351_45651 , \45349_45649 , \45350_45650 );
xor \U$37716 ( \45352_45652 , \31333_31632 , \45351_45651 );
buf \U$37717 ( \45353_45653 , \45352_45652 );
buf \U$37719 ( \45354_45654 , \45353_45653 );
and \U$37720 ( \45355_45655 , \30670_29853 , \38037_38337_nG9b84 );
and \U$37721 ( \45356_45656 , \29551_29850 , \38363_38663_nG9b81 );
or \U$37722 ( \45357_45657 , \45355_45655 , \45356_45656 );
xor \U$37723 ( \45358_45658 , \29550_29849 , \45357_45657 );
buf \U$37724 ( \45359_45659 , \45358_45658 );
buf \U$37726 ( \45360_45660 , \45359_45659 );
xor \U$37727 ( \45361_45661 , \45354_45654 , \45360_45660 );
and \U$37728 ( \45362_45662 , \23495_23201 , \40543_40843_nG9b6c );
and \U$37729 ( \45363_45663 , \22899_23198 , \40740_41040_nG9b69 );
or \U$37730 ( \45364_45664 , \45362_45662 , \45363_45663 );
xor \U$37731 ( \45365_45665 , \22898_23197 , \45364_45664 );
buf \U$37732 ( \45366_45666 , \45365_45665 );
buf \U$37734 ( \45367_45667 , \45366_45666 );
xor \U$37735 ( \45368_45668 , \45361_45661 , \45367_45667 );
buf \U$37736 ( \45369_45669 , \45368_45668 );
xor \U$37737 ( \45370_45670 , \45348_45648 , \45369_45669 );
and \U$37738 ( \45371_45671 , \45164_45464 , \45170_45470 );
and \U$37739 ( \45372_45672 , \45164_45464 , \45177_45477 );
and \U$37740 ( \45373_45673 , \45170_45470 , \45177_45477 );
or \U$37741 ( \45374_45674 , \45371_45671 , \45372_45672 , \45373_45673 );
buf \U$37742 ( \45375_45675 , \45374_45674 );
xor \U$37743 ( \45376_45676 , \45370_45670 , \45375_45675 );
buf \U$37744 ( \45377_45677 , \45376_45676 );
xor \U$37745 ( \45378_45678 , \45328_45628 , \45377_45677 );
buf \U$37746 ( \45379_45679 , \45378_45678 );
and \U$37747 ( \45380_45680 , \45179_45479 , \45199_45499 );
and \U$37748 ( \45381_45681 , \45179_45479 , \45205_45505 );
and \U$37749 ( \45382_45682 , \45199_45499 , \45205_45505 );
or \U$37750 ( \45383_45683 , \45380_45680 , \45381_45681 , \45382_45682 );
buf \U$37751 ( \45384_45684 , \45383_45683 );
and \U$37752 ( \45385_45685 , \45219_45519 , \45224_45524 );
and \U$37753 ( \45386_45686 , \45219_45519 , \45230_45530 );
and \U$37754 ( \45387_45687 , \45224_45524 , \45230_45530 );
or \U$37755 ( \45388_45688 , \45385_45685 , \45386_45686 , \45387_45687 );
buf \U$37756 ( \45389_45689 , \45388_45688 );
xor \U$37757 ( \45390_45690 , \45384_45684 , \45389_45689 );
and \U$37758 ( \45391_45691 , \45184_45484 , \45190_45490 );
and \U$37759 ( \45392_45692 , \45184_45484 , \45197_45497 );
and \U$37760 ( \45393_45693 , \45190_45490 , \45197_45497 );
or \U$37761 ( \45394_45694 , \45391_45691 , \45392_45692 , \45393_45693 );
buf \U$37762 ( \45395_45695 , \45394_45694 );
and \U$37763 ( \45396_45696 , \45136_45436 , \45142_45442 );
and \U$37764 ( \45397_45697 , \45136_45436 , \45149_45449 );
and \U$37765 ( \45398_45698 , \45142_45442 , \45149_45449 );
or \U$37766 ( \45399_45699 , \45396_45696 , \45397_45697 , \45398_45698 );
buf \U$37767 ( \45400_45700 , \45399_45699 );
xor \U$37768 ( \45401_45701 , \45395_45695 , \45400_45700 );
buf \U$37769 ( \45402_45702 , \45119_45419 );
xor \U$37770 ( \45403_45703 , \45401_45701 , \45402_45702 );
buf \U$37771 ( \45404_45704 , \45403_45703 );
xor \U$37772 ( \45405_45705 , \45390_45690 , \45404_45704 );
buf \U$37773 ( \45406_45706 , \45405_45705 );
xor \U$37774 ( \45407_45707 , \45379_45679 , \45406_45706 );
and \U$37775 ( \45408_45708 , \45214_45514 , \45232_45532 );
and \U$37776 ( \45409_45709 , \45214_45514 , \45238_45538 );
and \U$37777 ( \45410_45710 , \45232_45532 , \45238_45538 );
or \U$37778 ( \45411_45711 , \45408_45708 , \45409_45709 , \45410_45710 );
buf \U$37779 ( \45412_45712 , \45411_45711 );
xor \U$37780 ( \45413_45713 , \45407_45707 , \45412_45712 );
buf \U$37781 ( \45414_45714 , \45413_45713 );
and \U$37782 ( \45415_45715 , \45209_45509 , \45240_45540 );
and \U$37783 ( \45416_45716 , \45209_45509 , \45246_45546 );
and \U$37784 ( \45417_45717 , \45240_45540 , \45246_45546 );
or \U$37785 ( \45418_45718 , \45415_45715 , \45416_45716 , \45417_45717 );
buf \U$37786 ( \45419_45719 , \45418_45718 );
xor \U$37787 ( \45420_45720 , \45414_45714 , \45419_45719 );
and \U$37788 ( \45421_45721 , \45153_45453 , \45158_45458 );
and \U$37789 ( \45422_45722 , \45153_45453 , \45207_45507 );
and \U$37790 ( \45423_45723 , \45158_45458 , \45207_45507 );
or \U$37791 ( \45424_45724 , \45421_45721 , \45422_45722 , \45423_45723 );
buf \U$37792 ( \45425_45725 , \45424_45724 );
xor \U$37793 ( \45426_45726 , \45420_45720 , \45425_45725 );
and \U$37794 ( \45427_45727 , \45274_45574 , \45426_45726 );
and \U$37796 ( \45428_45728 , \45268_45568 , \45273_45573 );
or \U$37798 ( \45429_45729 , 1'b0 , \45428_45728 , 1'b0 );
xor \U$37799 ( \45430_45730 , \45427_45727 , \45429_45729 );
and \U$37801 ( \45431_45731 , \45261_45561 , \45267_45567 );
and \U$37802 ( \45432_45732 , \45263_45563 , \45267_45567 );
or \U$37803 ( \45433_45733 , 1'b0 , \45431_45731 , \45432_45732 );
xor \U$37804 ( \45434_45734 , \45430_45730 , \45433_45733 );
xor \U$37811 ( \45435_45735 , \45434_45734 , 1'b0 );
and \U$37812 ( \45436_45736 , \45414_45714 , \45419_45719 );
and \U$37813 ( \45437_45737 , \45414_45714 , \45425_45725 );
and \U$37814 ( \45438_45738 , \45419_45719 , \45425_45725 );
or \U$37815 ( \45439_45739 , \45436_45736 , \45437_45737 , \45438_45738 );
xor \U$37816 ( \45440_45740 , \45435_45735 , \45439_45739 );
and \U$37817 ( \45441_45741 , \45379_45679 , \45406_45706 );
and \U$37818 ( \45442_45742 , \45379_45679 , \45412_45712 );
and \U$37819 ( \45443_45743 , \45406_45706 , \45412_45712 );
or \U$37820 ( \45444_45744 , \45441_45741 , \45442_45742 , \45443_45743 );
buf \U$37821 ( \45445_45745 , \45444_45744 );
and \U$37822 ( \45446_45746 , \27141_26431 , \39663_39963_nG9b75 );
and \U$37823 ( \45447_45747 , \26129_26428 , \39904_40204_nG9b72 );
or \U$37824 ( \45448_45748 , \45446_45746 , \45447_45747 );
xor \U$37825 ( \45449_45749 , \26128_26427 , \45448_45748 );
buf \U$37826 ( \45450_45750 , \45449_45749 );
buf \U$37828 ( \45451_45751 , \45450_45750 );
and \U$37829 ( \45452_45752 , \25044_24792 , \40152_40452_nG9b6f );
and \U$37830 ( \45453_45753 , \24490_24789 , \40543_40843_nG9b6c );
or \U$37831 ( \45454_45754 , \45452_45752 , \45453_45753 );
xor \U$37832 ( \45455_45755 , \24489_24788 , \45454_45754 );
buf \U$37833 ( \45456_45756 , \45455_45755 );
buf \U$37835 ( \45457_45757 , \45456_45756 );
xor \U$37836 ( \45458_45758 , \45451_45751 , \45457_45757 );
and \U$37837 ( \45459_45759 , \20353_20155 , \41901_42201_nG9b5d );
and \U$37838 ( \45460_45760 , \19853_20152 , \42133_42433_nG9b5a );
or \U$37839 ( \45461_45761 , \45459_45759 , \45460_45760 );
xor \U$37840 ( \45462_45762 , \19852_20151 , \45461_45761 );
buf \U$37841 ( \45463_45763 , \45462_45762 );
buf \U$37843 ( \45464_45764 , \45463_45763 );
xor \U$37844 ( \45465_45765 , \45458_45758 , \45464_45764 );
buf \U$37845 ( \45466_45766 , \45465_45765 );
and \U$37846 ( \45467_45767 , \30670_29853 , \38363_38663_nG9b81 );
and \U$37847 ( \45468_45768 , \29551_29850 , \38668_38968_nG9b7e );
or \U$37848 ( \45469_45769 , \45467_45767 , \45468_45768 );
xor \U$37849 ( \45470_45770 , \29550_29849 , \45469_45769 );
buf \U$37850 ( \45471_45771 , \45470_45770 );
buf \U$37852 ( \45472_45772 , \45471_45771 );
and \U$37853 ( \45473_45773 , \28946_28118 , \39034_39334_nG9b7b );
and \U$37854 ( \45474_45774 , \27816_28115 , \39291_39591_nG9b78 );
or \U$37855 ( \45475_45775 , \45473_45773 , \45474_45774 );
xor \U$37856 ( \45476_45776 , \27815_28114 , \45475_45775 );
buf \U$37857 ( \45477_45777 , \45476_45776 );
buf \U$37859 ( \45478_45778 , \45477_45777 );
xor \U$37860 ( \45479_45779 , \45472_45772 , \45478_45778 );
and \U$37861 ( \45480_45780 , \23495_23201 , \40740_41040_nG9b69 );
and \U$37862 ( \45481_45781 , \22899_23198 , \41081_41381_nG9b66 );
or \U$37863 ( \45482_45782 , \45480_45780 , \45481_45781 );
xor \U$37864 ( \45483_45783 , \22898_23197 , \45482_45782 );
buf \U$37865 ( \45484_45784 , \45483_45783 );
buf \U$37867 ( \45485_45785 , \45484_45784 );
xor \U$37868 ( \45486_45786 , \45479_45779 , \45485_45785 );
buf \U$37869 ( \45487_45787 , \45486_45786 );
xor \U$37870 ( \45488_45788 , \45466_45766 , \45487_45787 );
and \U$37871 ( \45489_45789 , \17437_17297 , \42879_43179_nG9b51 );
or \U$37873 ( \45490_45790 , \45489_45789 , 1'b0 );
xor \U$37874 ( \45491_45791 , \16994_17293 , \45490_45790 );
buf \U$37875 ( \45492_45792 , \45491_45791 );
buf \U$37877 ( \45493_45793 , \45492_45792 );
and \U$37879 ( \45494_45794 , \32617_32916 , \37307_37607_nG9b8a );
or \U$37880 ( \45495_45795 , 1'b0 , \45494_45794 );
xor \U$37881 ( \45496_45796 , 1'b0 , \45495_45795 );
buf \U$37882 ( \45497_45797 , \45496_45796 );
buf \U$37884 ( \45498_45798 , \45497_45797 );
xor \U$37885 ( \45499_45799 , \45493_45793 , \45498_45798 );
and \U$37886 ( \45500_45800 , \31989_31636 , \37674_37974_nG9b87 );
and \U$37887 ( \45501_45801 , \31334_31633 , \38037_38337_nG9b84 );
or \U$37888 ( \45502_45802 , \45500_45800 , \45501_45801 );
xor \U$37889 ( \45503_45803 , \31333_31632 , \45502_45802 );
buf \U$37890 ( \45504_45804 , \45503_45803 );
buf \U$37892 ( \45505_45805 , \45504_45804 );
xor \U$37893 ( \45506_45806 , \45499_45799 , \45505_45805 );
buf \U$37894 ( \45507_45807 , \45506_45806 );
xor \U$37895 ( \45508_45808 , \45488_45788 , \45507_45807 );
buf \U$37896 ( \45509_45809 , \45508_45808 );
and \U$37897 ( \45510_45810 , \45348_45648 , \45369_45669 );
and \U$37898 ( \45511_45811 , \45348_45648 , \45375_45675 );
and \U$37899 ( \45512_45812 , \45369_45669 , \45375_45675 );
or \U$37900 ( \45513_45813 , \45510_45810 , \45511_45811 , \45512_45812 );
buf \U$37901 ( \45514_45814 , \45513_45813 );
xor \U$37902 ( \45515_45815 , \45509_45809 , \45514_45814 );
and \U$37903 ( \45516_45816 , \45284_45584 , \45305_45605 );
and \U$37904 ( \45517_45817 , \45284_45584 , \45325_45625 );
and \U$37905 ( \45518_45818 , \45305_45605 , \45325_45625 );
or \U$37906 ( \45519_45819 , \45516_45816 , \45517_45817 , \45518_45818 );
buf \U$37907 ( \45520_45820 , \45519_45819 );
xor \U$37908 ( \45521_45821 , \45515_45815 , \45520_45820 );
buf \U$37909 ( \45522_45822 , \45521_45821 );
and \U$37910 ( \45523_45823 , \45333_45633 , \45339_45639 );
and \U$37911 ( \45524_45824 , \45333_45633 , \45346_45646 );
and \U$37912 ( \45525_45825 , \45339_45639 , \45346_45646 );
or \U$37913 ( \45526_45826 , \45523_45823 , \45524_45824 , \45525_45825 );
buf \U$37914 ( \45527_45827 , \45526_45826 );
and \U$37915 ( \45528_45828 , \45312_45612 , \45316_45616 );
and \U$37916 ( \45529_45829 , \45312_45612 , \45323_45623 );
and \U$37917 ( \45530_45830 , \45316_45616 , \45323_45623 );
or \U$37918 ( \45531_45831 , \45528_45828 , \45529_45829 , \45530_45830 );
buf \U$37919 ( \45532_45832 , \45531_45831 );
xor \U$37920 ( \45533_45833 , \45527_45827 , \45532_45832 );
and \U$37921 ( \45534_45834 , \45290_45590 , \45296_45596 );
and \U$37922 ( \45535_45835 , \45290_45590 , \45303_45603 );
and \U$37923 ( \45536_45836 , \45296_45596 , \45303_45603 );
or \U$37924 ( \45537_45837 , \45534_45834 , \45535_45835 , \45536_45836 );
buf \U$37925 ( \45538_45838 , \45537_45837 );
xor \U$37926 ( \45539_45839 , \45533_45833 , \45538_45838 );
buf \U$37927 ( \45540_45840 , \45539_45839 );
and \U$37928 ( \45541_45841 , \45395_45695 , \45400_45700 );
and \U$37929 ( \45542_45842 , \45395_45695 , \45402_45702 );
and \U$37930 ( \45543_45843 , \45400_45700 , \45402_45702 );
or \U$37931 ( \45544_45844 , \45541_45841 , \45542_45842 , \45543_45843 );
buf \U$37932 ( \45545_45845 , \45544_45844 );
xor \U$37933 ( \45546_45846 , \45540_45840 , \45545_45845 );
and \U$37934 ( \45547_45847 , \45354_45654 , \45360_45660 );
and \U$37935 ( \45548_45848 , \45354_45654 , \45367_45667 );
and \U$37936 ( \45549_45849 , \45360_45660 , \45367_45667 );
or \U$37937 ( \45550_45850 , \45547_45847 , \45548_45848 , \45549_45849 );
buf \U$37938 ( \45551_45851 , \45550_45850 );
and \U$37939 ( \45552_45852 , \21908_21658 , \41385_41685_nG9b63 );
and \U$37940 ( \45553_45853 , \21356_21655 , \41663_41963_nG9b60 );
or \U$37941 ( \45554_45854 , \45552_45852 , \45553_45853 );
xor \U$37942 ( \45555_45855 , \21355_21654 , \45554_45854 );
buf \U$37943 ( \45556_45856 , \45555_45855 );
buf \U$37944 ( \45557_45857 , \45556_45856 );
not \U$37945 ( \45558_45858 , \45557_45857 );
xor \U$37946 ( \45559_45859 , \45551_45851 , \45558_45858 );
and \U$37947 ( \45560_45860 , \18908_18702 , \42466_42766_nG9b57 );
and \U$37948 ( \45561_45861 , \18400_18699 , \42548_42848_nG9b54 );
or \U$37949 ( \45562_45862 , \45560_45860 , \45561_45861 );
xor \U$37950 ( \45563_45863 , \18399_18698 , \45562_45862 );
buf \U$37951 ( \45564_45864 , \45563_45863 );
buf \U$37953 ( \45565_45865 , \45564_45864 );
xor \U$37954 ( \45566_45866 , \45559_45859 , \45565_45865 );
buf \U$37955 ( \45567_45867 , \45566_45866 );
xor \U$37956 ( \45568_45868 , \45546_45846 , \45567_45867 );
buf \U$37957 ( \45569_45869 , \45568_45868 );
xor \U$37958 ( \45570_45870 , \45522_45822 , \45569_45869 );
and \U$37959 ( \45571_45871 , \45384_45684 , \45389_45689 );
and \U$37960 ( \45572_45872 , \45384_45684 , \45404_45704 );
and \U$37961 ( \45573_45873 , \45389_45689 , \45404_45704 );
or \U$37962 ( \45574_45874 , \45571_45871 , \45572_45872 , \45573_45873 );
buf \U$37963 ( \45575_45875 , \45574_45874 );
xor \U$37964 ( \45576_45876 , \45570_45870 , \45575_45875 );
buf \U$37965 ( \45577_45877 , \45576_45876 );
xor \U$37966 ( \45578_45878 , \45445_45745 , \45577_45877 );
and \U$37967 ( \45579_45879 , \45279_45579 , \45327_45627 );
and \U$37968 ( \45580_45880 , \45279_45579 , \45377_45677 );
and \U$37969 ( \45581_45881 , \45327_45627 , \45377_45677 );
or \U$37970 ( \45582_45882 , \45579_45879 , \45580_45880 , \45581_45881 );
buf \U$37971 ( \45583_45883 , \45582_45882 );
xor \U$37972 ( \45584_45884 , \45578_45878 , \45583_45883 );
and \U$37973 ( \45585_45885 , \45440_45740 , \45584_45884 );
and \U$37975 ( \45586_45886 , \45434_45734 , \45439_45739 );
or \U$37977 ( \45587_45887 , 1'b0 , \45586_45886 , 1'b0 );
xor \U$37978 ( \45588_45888 , \45585_45885 , \45587_45887 );
and \U$37980 ( \45589_45889 , \45427_45727 , \45433_45733 );
and \U$37981 ( \45590_45890 , \45429_45729 , \45433_45733 );
or \U$37982 ( \45591_45891 , 1'b0 , \45589_45889 , \45590_45890 );
xor \U$37983 ( \45592_45892 , \45588_45888 , \45591_45891 );
xor \U$37990 ( \45593_45893 , \45592_45892 , 1'b0 );
and \U$37991 ( \45594_45894 , \45445_45745 , \45577_45877 );
and \U$37992 ( \45595_45895 , \45445_45745 , \45583_45883 );
and \U$37993 ( \45596_45896 , \45577_45877 , \45583_45883 );
or \U$37994 ( \45597_45897 , \45594_45894 , \45595_45895 , \45596_45896 );
xor \U$37995 ( \45598_45898 , \45593_45893 , \45597_45897 );
and \U$37996 ( \45599_45899 , \45522_45822 , \45569_45869 );
and \U$37997 ( \45600_45900 , \45522_45822 , \45575_45875 );
and \U$37998 ( \45601_45901 , \45569_45869 , \45575_45875 );
or \U$37999 ( \45602_45902 , \45599_45899 , \45600_45900 , \45601_45901 );
buf \U$38000 ( \45603_45903 , \45602_45902 );
and \U$38001 ( \45604_45904 , \18908_18702 , \42548_42848_nG9b54 );
and \U$38002 ( \45605_45905 , \18400_18699 , \42879_43179_nG9b51 );
or \U$38003 ( \45606_45906 , \45604_45904 , \45605_45905 );
xor \U$38004 ( \45607_45907 , \18399_18698 , \45606_45906 );
buf \U$38005 ( \45608_45908 , \45607_45907 );
buf \U$38007 ( \45609_45909 , \45608_45908 );
xor \U$38011 ( \45610_45910 , \16994_17293 , 1'b0 );
not \U$38012 ( \45611_45911 , \45610_45910 );
buf \U$38013 ( \45612_45912 , \45611_45911 );
buf \U$38015 ( \45613_45913 , \45612_45912 );
xor \U$38016 ( \45614_45914 , \45609_45909 , \45613_45913 );
and \U$38017 ( \45615_45915 , \21908_21658 , \41663_41963_nG9b60 );
and \U$38018 ( \45616_45916 , \21356_21655 , \41901_42201_nG9b5d );
or \U$38019 ( \45617_45917 , \45615_45915 , \45616_45916 );
xor \U$38020 ( \45618_45918 , \21355_21654 , \45617_45917 );
buf \U$38021 ( \45619_45919 , \45618_45918 );
buf \U$38023 ( \45620_45920 , \45619_45919 );
xor \U$38024 ( \45621_45921 , \45614_45914 , \45620_45920 );
buf \U$38025 ( \45622_45922 , \45621_45921 );
and \U$38026 ( \45623_45923 , \30670_29853 , \38668_38968_nG9b7e );
and \U$38027 ( \45624_45924 , \29551_29850 , \39034_39334_nG9b7b );
or \U$38028 ( \45625_45925 , \45623_45923 , \45624_45924 );
xor \U$38029 ( \45626_45926 , \29550_29849 , \45625_45925 );
buf \U$38030 ( \45627_45927 , \45626_45926 );
buf \U$38032 ( \45628_45928 , \45627_45927 );
and \U$38033 ( \45629_45929 , \28946_28118 , \39291_39591_nG9b78 );
and \U$38034 ( \45630_45930 , \27816_28115 , \39663_39963_nG9b75 );
or \U$38035 ( \45631_45931 , \45629_45929 , \45630_45930 );
xor \U$38036 ( \45632_45932 , \27815_28114 , \45631_45931 );
buf \U$38037 ( \45633_45933 , \45632_45932 );
buf \U$38039 ( \45634_45934 , \45633_45933 );
xor \U$38040 ( \45635_45935 , \45628_45928 , \45634_45934 );
and \U$38041 ( \45636_45936 , \23495_23201 , \41081_41381_nG9b66 );
and \U$38042 ( \45637_45937 , \22899_23198 , \41385_41685_nG9b63 );
or \U$38043 ( \45638_45938 , \45636_45936 , \45637_45937 );
xor \U$38044 ( \45639_45939 , \22898_23197 , \45638_45938 );
buf \U$38045 ( \45640_45940 , \45639_45939 );
buf \U$38047 ( \45641_45941 , \45640_45940 );
xor \U$38048 ( \45642_45942 , \45635_45935 , \45641_45941 );
buf \U$38049 ( \45643_45943 , \45642_45942 );
xor \U$38050 ( \45644_45944 , \45622_45922 , \45643_45943 );
and \U$38052 ( \45645_45945 , \32617_32916 , \37674_37974_nG9b87 );
or \U$38053 ( \45646_45946 , 1'b0 , \45645_45945 );
xor \U$38054 ( \45647_45947 , 1'b0 , \45646_45946 );
buf \U$38055 ( \45648_45948 , \45647_45947 );
buf \U$38057 ( \45649_45949 , \45648_45948 );
and \U$38058 ( \45650_45950 , \31989_31636 , \38037_38337_nG9b84 );
and \U$38059 ( \45651_45951 , \31334_31633 , \38363_38663_nG9b81 );
or \U$38060 ( \45652_45952 , \45650_45950 , \45651_45951 );
xor \U$38061 ( \45653_45953 , \31333_31632 , \45652_45952 );
buf \U$38062 ( \45654_45954 , \45653_45953 );
buf \U$38064 ( \45655_45955 , \45654_45954 );
xor \U$38065 ( \45656_45956 , \45649_45949 , \45655_45955 );
and \U$38066 ( \45657_45957 , \25044_24792 , \40543_40843_nG9b6c );
and \U$38067 ( \45658_45958 , \24490_24789 , \40740_41040_nG9b69 );
or \U$38068 ( \45659_45959 , \45657_45957 , \45658_45958 );
xor \U$38069 ( \45660_45960 , \24489_24788 , \45659_45959 );
buf \U$38070 ( \45661_45961 , \45660_45960 );
buf \U$38072 ( \45662_45962 , \45661_45961 );
xor \U$38073 ( \45663_45963 , \45656_45956 , \45662_45962 );
buf \U$38074 ( \45664_45964 , \45663_45963 );
xor \U$38075 ( \45665_45965 , \45644_45944 , \45664_45964 );
buf \U$38076 ( \45666_45966 , \45665_45965 );
and \U$38077 ( \45667_45967 , \45451_45751 , \45457_45757 );
and \U$38078 ( \45668_45968 , \45451_45751 , \45464_45764 );
and \U$38079 ( \45669_45969 , \45457_45757 , \45464_45764 );
or \U$38080 ( \45670_45970 , \45667_45967 , \45668_45968 , \45669_45969 );
buf \U$38081 ( \45671_45971 , \45670_45970 );
and \U$38082 ( \45672_45972 , \45493_45793 , \45498_45798 );
and \U$38083 ( \45673_45973 , \45493_45793 , \45505_45805 );
and \U$38084 ( \45674_45974 , \45498_45798 , \45505_45805 );
or \U$38085 ( \45675_45975 , \45672_45972 , \45673_45973 , \45674_45974 );
buf \U$38086 ( \45676_45976 , \45675_45975 );
xor \U$38087 ( \45677_45977 , \45671_45971 , \45676_45976 );
and \U$38088 ( \45678_45978 , \45472_45772 , \45478_45778 );
and \U$38089 ( \45679_45979 , \45472_45772 , \45485_45785 );
and \U$38090 ( \45680_45980 , \45478_45778 , \45485_45785 );
or \U$38091 ( \45681_45981 , \45678_45978 , \45679_45979 , \45680_45980 );
buf \U$38092 ( \45682_45982 , \45681_45981 );
xor \U$38093 ( \45683_45983 , \45677_45977 , \45682_45982 );
buf \U$38094 ( \45684_45984 , \45683_45983 );
xor \U$38095 ( \45685_45985 , \45666_45966 , \45684_45984 );
and \U$38096 ( \45686_45986 , \45527_45827 , \45532_45832 );
and \U$38097 ( \45687_45987 , \45527_45827 , \45538_45838 );
and \U$38098 ( \45688_45988 , \45532_45832 , \45538_45838 );
or \U$38099 ( \45689_45989 , \45686_45986 , \45687_45987 , \45688_45988 );
buf \U$38100 ( \45690_45990 , \45689_45989 );
xor \U$38101 ( \45691_45991 , \45685_45985 , \45690_45990 );
buf \U$38102 ( \45692_45992 , \45691_45991 );
and \U$38103 ( \45693_45993 , \45540_45840 , \45545_45845 );
and \U$38104 ( \45694_45994 , \45540_45840 , \45567_45867 );
and \U$38105 ( \45695_45995 , \45545_45845 , \45567_45867 );
or \U$38106 ( \45696_45996 , \45693_45993 , \45694_45994 , \45695_45995 );
buf \U$38107 ( \45697_45997 , \45696_45996 );
xor \U$38108 ( \45698_45998 , \45692_45992 , \45697_45997 );
and \U$38109 ( \45699_45999 , \45466_45766 , \45487_45787 );
and \U$38110 ( \45700_46000 , \45466_45766 , \45507_45807 );
and \U$38111 ( \45701_46001 , \45487_45787 , \45507_45807 );
or \U$38112 ( \45702_46002 , \45699_45999 , \45700_46000 , \45701_46001 );
buf \U$38113 ( \45703_46003 , \45702_46002 );
and \U$38114 ( \45704_46004 , \27141_26431 , \39904_40204_nG9b72 );
and \U$38115 ( \45705_46005 , \26129_26428 , \40152_40452_nG9b6f );
or \U$38116 ( \45706_46006 , \45704_46004 , \45705_46005 );
xor \U$38117 ( \45707_46007 , \26128_26427 , \45706_46006 );
buf \U$38118 ( \45708_46008 , \45707_46007 );
buf \U$38120 ( \45709_46009 , \45708_46008 );
buf \U$38121 ( \45710_46010 , \45557_45857 );
xor \U$38122 ( \45711_46011 , \45709_46009 , \45710_46010 );
and \U$38123 ( \45712_46012 , \20353_20155 , \42133_42433_nG9b5a );
and \U$38124 ( \45713_46013 , \19853_20152 , \42466_42766_nG9b57 );
or \U$38125 ( \45714_46014 , \45712_46012 , \45713_46013 );
xor \U$38126 ( \45715_46015 , \19852_20151 , \45714_46014 );
buf \U$38127 ( \45716_46016 , \45715_46015 );
buf \U$38129 ( \45717_46017 , \45716_46016 );
xor \U$38130 ( \45718_46018 , \45711_46011 , \45717_46017 );
buf \U$38131 ( \45719_46019 , \45718_46018 );
xor \U$38132 ( \45720_46020 , \45703_46003 , \45719_46019 );
and \U$38133 ( \45721_46021 , \45551_45851 , \45558_45858 );
and \U$38134 ( \45722_46022 , \45551_45851 , \45565_45865 );
and \U$38135 ( \45723_46023 , \45558_45858 , \45565_45865 );
or \U$38136 ( \45724_46024 , \45721_46021 , \45722_46022 , \45723_46023 );
buf \U$38137 ( \45725_46025 , \45724_46024 );
xor \U$38138 ( \45726_46026 , \45720_46020 , \45725_46025 );
buf \U$38139 ( \45727_46027 , \45726_46026 );
xor \U$38140 ( \45728_46028 , \45698_45998 , \45727_46027 );
buf \U$38141 ( \45729_46029 , \45728_46028 );
xor \U$38142 ( \45730_46030 , \45603_45903 , \45729_46029 );
and \U$38143 ( \45731_46031 , \45509_45809 , \45514_45814 );
and \U$38144 ( \45732_46032 , \45509_45809 , \45520_45820 );
and \U$38145 ( \45733_46033 , \45514_45814 , \45520_45820 );
or \U$38146 ( \45734_46034 , \45731_46031 , \45732_46032 , \45733_46033 );
buf \U$38147 ( \45735_46035 , \45734_46034 );
xor \U$38148 ( \45736_46036 , \45730_46030 , \45735_46035 );
and \U$38149 ( \45737_46037 , \45598_45898 , \45736_46036 );
and \U$38151 ( \45738_46038 , \45592_45892 , \45597_45897 );
or \U$38153 ( \45739_46039 , 1'b0 , \45738_46038 , 1'b0 );
xor \U$38154 ( \45740_46040 , \45737_46037 , \45739_46039 );
and \U$38156 ( \45741_46041 , \45585_45885 , \45591_45891 );
and \U$38157 ( \45742_46042 , \45587_45887 , \45591_45891 );
or \U$38158 ( \45743_46043 , 1'b0 , \45741_46041 , \45742_46042 );
xor \U$38159 ( \45744_46044 , \45740_46040 , \45743_46043 );
xor \U$38166 ( \45745_46045 , \45744_46044 , 1'b0 );
and \U$38167 ( \45746_46046 , \45692_45992 , \45697_45997 );
and \U$38168 ( \45747_46047 , \45692_45992 , \45727_46027 );
and \U$38169 ( \45748_46048 , \45697_45997 , \45727_46027 );
or \U$38170 ( \45749_46049 , \45746_46046 , \45747_46047 , \45748_46048 );
buf \U$38171 ( \45750_46050 , \45749_46049 );
and \U$38172 ( \45751_46051 , \45671_45971 , \45676_45976 );
and \U$38173 ( \45752_46052 , \45671_45971 , \45682_45982 );
and \U$38174 ( \45753_46053 , \45676_45976 , \45682_45982 );
or \U$38175 ( \45754_46054 , \45751_46051 , \45752_46052 , \45753_46053 );
buf \U$38176 ( \45755_46055 , \45754_46054 );
and \U$38177 ( \45756_46056 , \45709_46009 , \45710_46010 );
and \U$38178 ( \45757_46057 , \45709_46009 , \45717_46017 );
and \U$38179 ( \45758_46058 , \45710_46010 , \45717_46017 );
or \U$38180 ( \45759_46059 , \45756_46056 , \45757_46057 , \45758_46058 );
buf \U$38181 ( \45760_46060 , \45759_46059 );
xor \U$38182 ( \45761_46061 , \45755_46055 , \45760_46060 );
and \U$38183 ( \45762_46062 , \28946_28118 , \39663_39963_nG9b75 );
and \U$38184 ( \45763_46063 , \27816_28115 , \39904_40204_nG9b72 );
or \U$38185 ( \45764_46064 , \45762_46062 , \45763_46063 );
xor \U$38186 ( \45765_46065 , \27815_28114 , \45764_46064 );
buf \U$38187 ( \45766_46066 , \45765_46065 );
buf \U$38189 ( \45767_46067 , \45766_46066 );
and \U$38190 ( \45768_46068 , \27141_26431 , \40152_40452_nG9b6f );
and \U$38191 ( \45769_46069 , \26129_26428 , \40543_40843_nG9b6c );
or \U$38192 ( \45770_46070 , \45768_46068 , \45769_46069 );
xor \U$38193 ( \45771_46071 , \26128_26427 , \45770_46070 );
buf \U$38194 ( \45772_46072 , \45771_46071 );
buf \U$38196 ( \45773_46073 , \45772_46072 );
xor \U$38197 ( \45774_46074 , \45767_46067 , \45773_46073 );
and \U$38198 ( \45775_46075 , \20353_20155 , \42466_42766_nG9b57 );
and \U$38199 ( \45776_46076 , \19853_20152 , \42548_42848_nG9b54 );
or \U$38200 ( \45777_46077 , \45775_46075 , \45776_46076 );
xor \U$38201 ( \45778_46078 , \19852_20151 , \45777_46077 );
buf \U$38202 ( \45779_46079 , \45778_46078 );
buf \U$38204 ( \45780_46080 , \45779_46079 );
xor \U$38205 ( \45781_46081 , \45774_46074 , \45780_46080 );
buf \U$38206 ( \45782_46082 , \45781_46081 );
xor \U$38207 ( \45783_46083 , \45761_46061 , \45782_46082 );
buf \U$38208 ( \45784_46084 , \45783_46083 );
and \U$38209 ( \45785_46085 , \45703_46003 , \45719_46019 );
and \U$38210 ( \45786_46086 , \45703_46003 , \45725_46025 );
and \U$38211 ( \45787_46087 , \45719_46019 , \45725_46025 );
or \U$38212 ( \45788_46088 , \45785_46085 , \45786_46086 , \45787_46087 );
buf \U$38213 ( \45789_46089 , \45788_46088 );
xor \U$38214 ( \45790_46090 , \45784_46084 , \45789_46089 );
and \U$38215 ( \45791_46091 , \45666_45966 , \45684_45984 );
and \U$38216 ( \45792_46092 , \45666_45966 , \45690_45990 );
and \U$38217 ( \45793_46093 , \45684_45984 , \45690_45990 );
or \U$38218 ( \45794_46094 , \45791_46091 , \45792_46092 , \45793_46093 );
buf \U$38219 ( \45795_46095 , \45794_46094 );
xor \U$38220 ( \45796_46096 , \45790_46090 , \45795_46095 );
buf \U$38221 ( \45797_46097 , \45796_46096 );
xor \U$38222 ( \45798_46098 , \45750_46050 , \45797_46097 );
and \U$38223 ( \45799_46099 , \31989_31636 , \38363_38663_nG9b81 );
and \U$38224 ( \45800_46100 , \31334_31633 , \38668_38968_nG9b7e );
or \U$38225 ( \45801_46101 , \45799_46099 , \45800_46100 );
xor \U$38226 ( \45802_46102 , \31333_31632 , \45801_46101 );
buf \U$38227 ( \45803_46103 , \45802_46102 );
buf \U$38229 ( \45804_46104 , \45803_46103 );
and \U$38230 ( \45805_46105 , \30670_29853 , \39034_39334_nG9b7b );
and \U$38231 ( \45806_46106 , \29551_29850 , \39291_39591_nG9b78 );
or \U$38232 ( \45807_46107 , \45805_46105 , \45806_46106 );
xor \U$38233 ( \45808_46108 , \29550_29849 , \45807_46107 );
buf \U$38234 ( \45809_46109 , \45808_46108 );
buf \U$38236 ( \45810_46110 , \45809_46109 );
xor \U$38237 ( \45811_46111 , \45804_46104 , \45810_46110 );
and \U$38238 ( \45812_46112 , \23495_23201 , \41385_41685_nG9b63 );
and \U$38239 ( \45813_46113 , \22899_23198 , \41663_41963_nG9b60 );
or \U$38240 ( \45814_46114 , \45812_46112 , \45813_46113 );
xor \U$38241 ( \45815_46115 , \22898_23197 , \45814_46114 );
buf \U$38242 ( \45816_46116 , \45815_46115 );
buf \U$38244 ( \45817_46117 , \45816_46116 );
xor \U$38245 ( \45818_46118 , \45811_46111 , \45817_46117 );
buf \U$38246 ( \45819_46119 , \45818_46118 );
and \U$38248 ( \45820_46120 , \32617_32916 , \38037_38337_nG9b84 );
or \U$38249 ( \45821_46121 , 1'b0 , \45820_46120 );
xor \U$38250 ( \45822_46122 , 1'b0 , \45821_46121 );
buf \U$38251 ( \45823_46123 , \45822_46122 );
buf \U$38253 ( \45824_46124 , \45823_46123 );
and \U$38254 ( \45825_46125 , \25044_24792 , \40740_41040_nG9b69 );
and \U$38255 ( \45826_46126 , \24490_24789 , \41081_41381_nG9b66 );
or \U$38256 ( \45827_46127 , \45825_46125 , \45826_46126 );
xor \U$38257 ( \45828_46128 , \24489_24788 , \45827_46127 );
buf \U$38258 ( \45829_46129 , \45828_46128 );
buf \U$38260 ( \45830_46130 , \45829_46129 );
xor \U$38261 ( \45831_46131 , \45824_46124 , \45830_46130 );
and \U$38262 ( \45832_46132 , \21908_21658 , \41901_42201_nG9b5d );
and \U$38263 ( \45833_46133 , \21356_21655 , \42133_42433_nG9b5a );
or \U$38264 ( \45834_46134 , \45832_46132 , \45833_46133 );
xor \U$38265 ( \45835_46135 , \21355_21654 , \45834_46134 );
buf \U$38266 ( \45836_46136 , \45835_46135 );
buf \U$38268 ( \45837_46137 , \45836_46136 );
xor \U$38269 ( \45838_46138 , \45831_46131 , \45837_46137 );
buf \U$38270 ( \45839_46139 , \45838_46138 );
xor \U$38271 ( \45840_46140 , \45819_46119 , \45839_46139 );
and \U$38272 ( \45841_46141 , \45649_45949 , \45655_45955 );
and \U$38273 ( \45842_46142 , \45649_45949 , \45662_45962 );
and \U$38274 ( \45843_46143 , \45655_45955 , \45662_45962 );
or \U$38275 ( \45844_46144 , \45841_46141 , \45842_46142 , \45843_46143 );
buf \U$38276 ( \45845_46145 , \45844_46144 );
xor \U$38277 ( \45846_46146 , \45840_46140 , \45845_46145 );
buf \U$38278 ( \45847_46147 , \45846_46146 );
and \U$38279 ( \45848_46148 , \45622_45922 , \45643_45943 );
and \U$38280 ( \45849_46149 , \45622_45922 , \45664_45964 );
and \U$38281 ( \45850_46150 , \45643_45943 , \45664_45964 );
or \U$38282 ( \45851_46151 , \45848_46148 , \45849_46149 , \45850_46150 );
buf \U$38283 ( \45852_46152 , \45851_46151 );
xor \U$38284 ( \45853_46153 , \45847_46147 , \45852_46152 );
and \U$38285 ( \45854_46154 , \45609_45909 , \45613_45913 );
and \U$38286 ( \45855_46155 , \45609_45909 , \45620_45920 );
and \U$38287 ( \45856_46156 , \45613_45913 , \45620_45920 );
or \U$38288 ( \45857_46157 , \45854_46154 , \45855_46155 , \45856_46156 );
buf \U$38289 ( \45858_46158 , \45857_46157 );
and \U$38290 ( \45859_46159 , \45628_45928 , \45634_45934 );
and \U$38291 ( \45860_46160 , \45628_45928 , \45641_45941 );
and \U$38292 ( \45861_46161 , \45634_45934 , \45641_45941 );
or \U$38293 ( \45862_46162 , \45859_46159 , \45860_46160 , \45861_46161 );
buf \U$38294 ( \45863_46163 , \45862_46162 );
xor \U$38295 ( \45864_46164 , \45858_46158 , \45863_46163 );
and \U$38296 ( \45865_46165 , \18908_18702 , \42879_43179_nG9b51 );
or \U$38298 ( \45866_46166 , \45865_46165 , 1'b0 );
xor \U$38299 ( \45867_46167 , \18399_18698 , \45866_46166 );
buf \U$38300 ( \45868_46168 , \45867_46167 );
buf \U$38301 ( \45869_46169 , \45868_46168 );
not \U$38302 ( \45870_46170 , \45869_46169 );
xor \U$38303 ( \45871_46171 , \45864_46164 , \45870_46170 );
buf \U$38304 ( \45872_46172 , \45871_46171 );
xor \U$38305 ( \45873_46173 , \45853_46153 , \45872_46172 );
buf \U$38306 ( \45874_46174 , \45873_46173 );
xor \U$38307 ( \45875_46175 , \45798_46098 , \45874_46174 );
xor \U$38308 ( \45876_46176 , \45745_46045 , \45875_46175 );
and \U$38309 ( \45877_46177 , \45603_45903 , \45729_46029 );
and \U$38310 ( \45878_46178 , \45603_45903 , \45735_46035 );
and \U$38311 ( \45879_46179 , \45729_46029 , \45735_46035 );
or \U$38312 ( \45880_46180 , \45877_46177 , \45878_46178 , \45879_46179 );
and \U$38313 ( \45881_46181 , \45876_46176 , \45880_46180 );
and \U$38315 ( \45882_46182 , \45744_46044 , \45875_46175 );
or \U$38317 ( \45883_46183 , 1'b0 , \45882_46182 , 1'b0 );
xor \U$38318 ( \45884_46184 , \45881_46181 , \45883_46183 );
and \U$38320 ( \45885_46185 , \45737_46037 , \45743_46043 );
and \U$38321 ( \45886_46186 , \45739_46039 , \45743_46043 );
or \U$38322 ( \45887_46187 , 1'b0 , \45885_46185 , \45886_46186 );
xor \U$38323 ( \45888_46188 , \45884_46184 , \45887_46187 );
xor \U$38330 ( \45889_46189 , \45888_46188 , 1'b0 );
and \U$38331 ( \45890_46190 , \45784_46084 , \45789_46089 );
and \U$38332 ( \45891_46191 , \45784_46084 , \45795_46095 );
and \U$38333 ( \45892_46192 , \45789_46089 , \45795_46095 );
or \U$38334 ( \45893_46193 , \45890_46190 , \45891_46191 , \45892_46192 );
buf \U$38335 ( \45894_46194 , \45893_46193 );
and \U$38336 ( \45895_46195 , \20353_20155 , \42548_42848_nG9b54 );
and \U$38337 ( \45896_46196 , \19853_20152 , \42879_43179_nG9b51 );
or \U$38338 ( \45897_46197 , \45895_46195 , \45896_46196 );
xor \U$38339 ( \45898_46198 , \19852_20151 , \45897_46197 );
buf \U$38340 ( \45899_46199 , \45898_46198 );
buf \U$38342 ( \45900_46200 , \45899_46199 );
xor \U$38346 ( \45901_46201 , \18399_18698 , 1'b0 );
not \U$38347 ( \45902_46202 , \45901_46201 );
buf \U$38348 ( \45903_46203 , \45902_46202 );
buf \U$38350 ( \45904_46204 , \45903_46203 );
xor \U$38351 ( \45905_46205 , \45900_46200 , \45904_46204 );
and \U$38352 ( \45906_46206 , \23495_23201 , \41663_41963_nG9b60 );
and \U$38353 ( \45907_46207 , \22899_23198 , \41901_42201_nG9b5d );
or \U$38354 ( \45908_46208 , \45906_46206 , \45907_46207 );
xor \U$38355 ( \45909_46209 , \22898_23197 , \45908_46208 );
buf \U$38356 ( \45910_46210 , \45909_46209 );
buf \U$38358 ( \45911_46211 , \45910_46210 );
xor \U$38359 ( \45912_46212 , \45905_46205 , \45911_46211 );
buf \U$38360 ( \45913_46213 , \45912_46212 );
and \U$38362 ( \45914_46214 , \32617_32916 , \38363_38663_nG9b81 );
or \U$38363 ( \45915_46215 , 1'b0 , \45914_46214 );
xor \U$38364 ( \45916_46216 , 1'b0 , \45915_46215 );
buf \U$38365 ( \45917_46217 , \45916_46216 );
buf \U$38367 ( \45918_46218 , \45917_46217 );
and \U$38368 ( \45919_46219 , \28946_28118 , \39904_40204_nG9b72 );
and \U$38369 ( \45920_46220 , \27816_28115 , \40152_40452_nG9b6f );
or \U$38370 ( \45921_46221 , \45919_46219 , \45920_46220 );
xor \U$38371 ( \45922_46222 , \27815_28114 , \45921_46221 );
buf \U$38372 ( \45923_46223 , \45922_46222 );
buf \U$38374 ( \45924_46224 , \45923_46223 );
xor \U$38375 ( \45925_46225 , \45918_46218 , \45924_46224 );
and \U$38376 ( \45926_46226 , \27141_26431 , \40543_40843_nG9b6c );
and \U$38377 ( \45927_46227 , \26129_26428 , \40740_41040_nG9b69 );
or \U$38378 ( \45928_46228 , \45926_46226 , \45927_46227 );
xor \U$38379 ( \45929_46229 , \26128_26427 , \45928_46228 );
buf \U$38380 ( \45930_46230 , \45929_46229 );
buf \U$38382 ( \45931_46231 , \45930_46230 );
xor \U$38383 ( \45932_46232 , \45925_46225 , \45931_46231 );
buf \U$38384 ( \45933_46233 , \45932_46232 );
xor \U$38385 ( \45934_46234 , \45913_46213 , \45933_46233 );
and \U$38386 ( \45935_46235 , \45824_46124 , \45830_46130 );
and \U$38387 ( \45936_46236 , \45824_46124 , \45837_46137 );
and \U$38388 ( \45937_46237 , \45830_46130 , \45837_46137 );
or \U$38389 ( \45938_46238 , \45935_46235 , \45936_46236 , \45937_46237 );
buf \U$38390 ( \45939_46239 , \45938_46238 );
xor \U$38391 ( \45940_46240 , \45934_46234 , \45939_46239 );
buf \U$38392 ( \45941_46241 , \45940_46240 );
and \U$38393 ( \45942_46242 , \45858_46158 , \45863_46163 );
and \U$38394 ( \45943_46243 , \45858_46158 , \45870_46170 );
and \U$38395 ( \45944_46244 , \45863_46163 , \45870_46170 );
or \U$38396 ( \45945_46245 , \45942_46242 , \45943_46243 , \45944_46244 );
buf \U$38397 ( \45946_46246 , \45945_46245 );
xor \U$38398 ( \45947_46247 , \45941_46241 , \45946_46246 );
and \U$38399 ( \45948_46248 , \45819_46119 , \45839_46139 );
and \U$38400 ( \45949_46249 , \45819_46119 , \45845_46145 );
and \U$38401 ( \45950_46250 , \45839_46139 , \45845_46145 );
or \U$38402 ( \45951_46251 , \45948_46248 , \45949_46249 , \45950_46250 );
buf \U$38403 ( \45952_46252 , \45951_46251 );
xor \U$38404 ( \45953_46253 , \45947_46247 , \45952_46252 );
buf \U$38405 ( \45954_46254 , \45953_46253 );
xor \U$38406 ( \45955_46255 , \45894_46194 , \45954_46254 );
and \U$38407 ( \45956_46256 , \45755_46055 , \45760_46060 );
and \U$38408 ( \45957_46257 , \45755_46055 , \45782_46082 );
and \U$38409 ( \45958_46258 , \45760_46060 , \45782_46082 );
or \U$38410 ( \45959_46259 , \45956_46256 , \45957_46257 , \45958_46258 );
buf \U$38411 ( \45960_46260 , \45959_46259 );
and \U$38412 ( \45961_46261 , \45804_46104 , \45810_46110 );
and \U$38413 ( \45962_46262 , \45804_46104 , \45817_46117 );
and \U$38414 ( \45963_46263 , \45810_46110 , \45817_46117 );
or \U$38415 ( \45964_46264 , \45961_46261 , \45962_46262 , \45963_46263 );
buf \U$38416 ( \45965_46265 , \45964_46264 );
buf \U$38417 ( \45966_46266 , \45869_46169 );
xor \U$38418 ( \45967_46267 , \45965_46265 , \45966_46266 );
and \U$38419 ( \45968_46268 , \21908_21658 , \42133_42433_nG9b5a );
and \U$38420 ( \45969_46269 , \21356_21655 , \42466_42766_nG9b57 );
or \U$38421 ( \45970_46270 , \45968_46268 , \45969_46269 );
xor \U$38422 ( \45971_46271 , \21355_21654 , \45970_46270 );
buf \U$38423 ( \45972_46272 , \45971_46271 );
buf \U$38425 ( \45973_46273 , \45972_46272 );
xor \U$38426 ( \45974_46274 , \45967_46267 , \45973_46273 );
buf \U$38427 ( \45975_46275 , \45974_46274 );
and \U$38428 ( \45976_46276 , \31989_31636 , \38668_38968_nG9b7e );
and \U$38429 ( \45977_46277 , \31334_31633 , \39034_39334_nG9b7b );
or \U$38430 ( \45978_46278 , \45976_46276 , \45977_46277 );
xor \U$38431 ( \45979_46279 , \31333_31632 , \45978_46278 );
buf \U$38432 ( \45980_46280 , \45979_46279 );
buf \U$38434 ( \45981_46281 , \45980_46280 );
and \U$38435 ( \45982_46282 , \30670_29853 , \39291_39591_nG9b78 );
and \U$38436 ( \45983_46283 , \29551_29850 , \39663_39963_nG9b75 );
or \U$38437 ( \45984_46284 , \45982_46282 , \45983_46283 );
xor \U$38438 ( \45985_46285 , \29550_29849 , \45984_46284 );
buf \U$38439 ( \45986_46286 , \45985_46285 );
buf \U$38441 ( \45987_46287 , \45986_46286 );
xor \U$38442 ( \45988_46288 , \45981_46281 , \45987_46287 );
and \U$38443 ( \45989_46289 , \25044_24792 , \41081_41381_nG9b66 );
and \U$38444 ( \45990_46290 , \24490_24789 , \41385_41685_nG9b63 );
or \U$38445 ( \45991_46291 , \45989_46289 , \45990_46290 );
xor \U$38446 ( \45992_46292 , \24489_24788 , \45991_46291 );
buf \U$38447 ( \45993_46293 , \45992_46292 );
buf \U$38449 ( \45994_46294 , \45993_46293 );
xor \U$38450 ( \45995_46295 , \45988_46288 , \45994_46294 );
buf \U$38451 ( \45996_46296 , \45995_46295 );
xor \U$38452 ( \45997_46297 , \45975_46275 , \45996_46296 );
and \U$38453 ( \45998_46298 , \45767_46067 , \45773_46073 );
and \U$38454 ( \45999_46299 , \45767_46067 , \45780_46080 );
and \U$38455 ( \46000_46300 , \45773_46073 , \45780_46080 );
or \U$38456 ( \46001_46301 , \45998_46298 , \45999_46299 , \46000_46300 );
buf \U$38457 ( \46002_46302 , \46001_46301 );
xor \U$38458 ( \46003_46303 , \45997_46297 , \46002_46302 );
buf \U$38459 ( \46004_46304 , \46003_46303 );
xor \U$38460 ( \46005_46305 , \45960_46260 , \46004_46304 );
and \U$38461 ( \46006_46306 , \45847_46147 , \45852_46152 );
and \U$38462 ( \46007_46307 , \45847_46147 , \45872_46172 );
and \U$38463 ( \46008_46308 , \45852_46152 , \45872_46172 );
or \U$38464 ( \46009_46309 , \46006_46306 , \46007_46307 , \46008_46308 );
buf \U$38465 ( \46010_46310 , \46009_46309 );
xor \U$38466 ( \46011_46311 , \46005_46305 , \46010_46310 );
buf \U$38467 ( \46012_46312 , \46011_46311 );
xor \U$38468 ( \46013_46313 , \45955_46255 , \46012_46312 );
xor \U$38469 ( \46014_46314 , \45889_46189 , \46013_46313 );
and \U$38470 ( \46015_46315 , \45750_46050 , \45797_46097 );
and \U$38471 ( \46016_46316 , \45750_46050 , \45874_46174 );
and \U$38472 ( \46017_46317 , \45797_46097 , \45874_46174 );
or \U$38473 ( \46018_46318 , \46015_46315 , \46016_46316 , \46017_46317 );
and \U$38474 ( \46019_46319 , \46014_46314 , \46018_46318 );
and \U$38476 ( \46020_46320 , \45888_46188 , \46013_46313 );
or \U$38478 ( \46021_46321 , 1'b0 , \46020_46320 , 1'b0 );
xor \U$38479 ( \46022_46322 , \46019_46319 , \46021_46321 );
and \U$38481 ( \46023_46323 , \45881_46181 , \45887_46187 );
and \U$38482 ( \46024_46324 , \45883_46183 , \45887_46187 );
or \U$38483 ( \46025_46325 , 1'b0 , \46023_46323 , \46024_46324 );
xor \U$38484 ( \46026_46326 , \46022_46322 , \46025_46325 );
xor \U$38491 ( \46027_46327 , \46026_46326 , 1'b0 );
and \U$38492 ( \46028_46328 , \45894_46194 , \45954_46254 );
and \U$38493 ( \46029_46329 , \45894_46194 , \46012_46312 );
and \U$38494 ( \46030_46330 , \45954_46254 , \46012_46312 );
or \U$38495 ( \46031_46331 , \46028_46328 , \46029_46329 , \46030_46330 );
xor \U$38496 ( \46032_46332 , \46027_46327 , \46031_46331 );
and \U$38497 ( \46033_46333 , \28946_28118 , \40152_40452_nG9b6f );
and \U$38498 ( \46034_46334 , \27816_28115 , \40543_40843_nG9b6c );
or \U$38499 ( \46035_46335 , \46033_46333 , \46034_46334 );
xor \U$38500 ( \46036_46336 , \27815_28114 , \46035_46335 );
buf \U$38501 ( \46037_46337 , \46036_46336 );
buf \U$38503 ( \46038_46338 , \46037_46337 );
and \U$38504 ( \46039_46339 , \27141_26431 , \40740_41040_nG9b69 );
and \U$38505 ( \46040_46340 , \26129_26428 , \41081_41381_nG9b66 );
or \U$38506 ( \46041_46341 , \46039_46339 , \46040_46340 );
xor \U$38507 ( \46042_46342 , \26128_26427 , \46041_46341 );
buf \U$38508 ( \46043_46343 , \46042_46342 );
buf \U$38510 ( \46044_46344 , \46043_46343 );
xor \U$38511 ( \46045_46345 , \46038_46338 , \46044_46344 );
and \U$38512 ( \46046_46346 , \23495_23201 , \41901_42201_nG9b5d );
and \U$38513 ( \46047_46347 , \22899_23198 , \42133_42433_nG9b5a );
or \U$38514 ( \46048_46348 , \46046_46346 , \46047_46347 );
xor \U$38515 ( \46049_46349 , \22898_23197 , \46048_46348 );
buf \U$38516 ( \46050_46350 , \46049_46349 );
buf \U$38518 ( \46051_46351 , \46050_46350 );
xor \U$38519 ( \46052_46352 , \46045_46345 , \46051_46351 );
buf \U$38520 ( \46053_46353 , \46052_46352 );
and \U$38521 ( \46054_46354 , \20353_20155 , \42879_43179_nG9b51 );
or \U$38523 ( \46055_46355 , \46054_46354 , 1'b0 );
xor \U$38524 ( \46056_46356 , \19852_20151 , \46055_46355 );
buf \U$38525 ( \46057_46357 , \46056_46356 );
buf \U$38526 ( \46058_46358 , \46057_46357 );
not \U$38527 ( \46059_46359 , \46058_46358 );
and \U$38528 ( \46060_46360 , \30670_29853 , \39663_39963_nG9b75 );
and \U$38529 ( \46061_46361 , \29551_29850 , \39904_40204_nG9b72 );
or \U$38530 ( \46062_46362 , \46060_46360 , \46061_46361 );
xor \U$38531 ( \46063_46363 , \29550_29849 , \46062_46362 );
buf \U$38532 ( \46064_46364 , \46063_46363 );
buf \U$38534 ( \46065_46365 , \46064_46364 );
xor \U$38535 ( \46066_46366 , \46059_46359 , \46065_46365 );
and \U$38536 ( \46067_46367 , \21908_21658 , \42466_42766_nG9b57 );
and \U$38537 ( \46068_46368 , \21356_21655 , \42548_42848_nG9b54 );
or \U$38538 ( \46069_46369 , \46067_46367 , \46068_46368 );
xor \U$38539 ( \46070_46370 , \21355_21654 , \46069_46369 );
buf \U$38540 ( \46071_46371 , \46070_46370 );
buf \U$38542 ( \46072_46372 , \46071_46371 );
xor \U$38543 ( \46073_46373 , \46066_46366 , \46072_46372 );
buf \U$38544 ( \46074_46374 , \46073_46373 );
xor \U$38545 ( \46075_46375 , \46053_46353 , \46074_46374 );
and \U$38547 ( \46076_46376 , \32617_32916 , \38668_38968_nG9b7e );
or \U$38548 ( \46077_46377 , 1'b0 , \46076_46376 );
xor \U$38549 ( \46078_46378 , 1'b0 , \46077_46377 );
buf \U$38550 ( \46079_46379 , \46078_46378 );
buf \U$38552 ( \46080_46380 , \46079_46379 );
and \U$38553 ( \46081_46381 , \31989_31636 , \39034_39334_nG9b7b );
and \U$38554 ( \46082_46382 , \31334_31633 , \39291_39591_nG9b78 );
or \U$38555 ( \46083_46383 , \46081_46381 , \46082_46382 );
xor \U$38556 ( \46084_46384 , \31333_31632 , \46083_46383 );
buf \U$38557 ( \46085_46385 , \46084_46384 );
buf \U$38559 ( \46086_46386 , \46085_46385 );
xor \U$38560 ( \46087_46387 , \46080_46380 , \46086_46386 );
and \U$38561 ( \46088_46388 , \25044_24792 , \41385_41685_nG9b63 );
and \U$38562 ( \46089_46389 , \24490_24789 , \41663_41963_nG9b60 );
or \U$38563 ( \46090_46390 , \46088_46388 , \46089_46389 );
xor \U$38564 ( \46091_46391 , \24489_24788 , \46090_46390 );
buf \U$38565 ( \46092_46392 , \46091_46391 );
buf \U$38567 ( \46093_46393 , \46092_46392 );
xor \U$38568 ( \46094_46394 , \46087_46387 , \46093_46393 );
buf \U$38569 ( \46095_46395 , \46094_46394 );
xor \U$38570 ( \46096_46396 , \46075_46375 , \46095_46395 );
buf \U$38571 ( \46097_46397 , \46096_46396 );
and \U$38572 ( \46098_46398 , \45975_46275 , \45996_46296 );
and \U$38573 ( \46099_46399 , \45975_46275 , \46002_46302 );
and \U$38574 ( \46100_46400 , \45996_46296 , \46002_46302 );
or \U$38575 ( \46101_46401 , \46098_46398 , \46099_46399 , \46100_46400 );
buf \U$38576 ( \46102_46402 , \46101_46401 );
xor \U$38577 ( \46103_46403 , \46097_46397 , \46102_46402 );
and \U$38578 ( \46104_46404 , \45913_46213 , \45933_46233 );
and \U$38579 ( \46105_46405 , \45913_46213 , \45939_46239 );
and \U$38580 ( \46106_46406 , \45933_46233 , \45939_46239 );
or \U$38581 ( \46107_46407 , \46104_46404 , \46105_46405 , \46106_46406 );
buf \U$38582 ( \46108_46408 , \46107_46407 );
and \U$38583 ( \46109_46409 , \45900_46200 , \45904_46204 );
and \U$38584 ( \46110_46410 , \45900_46200 , \45911_46211 );
and \U$38585 ( \46111_46411 , \45904_46204 , \45911_46211 );
or \U$38586 ( \46112_46412 , \46109_46409 , \46110_46410 , \46111_46411 );
buf \U$38587 ( \46113_46413 , \46112_46412 );
and \U$38588 ( \46114_46414 , \45918_46218 , \45924_46224 );
and \U$38589 ( \46115_46415 , \45918_46218 , \45931_46231 );
and \U$38590 ( \46116_46416 , \45924_46224 , \45931_46231 );
or \U$38591 ( \46117_46417 , \46114_46414 , \46115_46415 , \46116_46416 );
buf \U$38592 ( \46118_46418 , \46117_46417 );
xor \U$38593 ( \46119_46419 , \46113_46413 , \46118_46418 );
and \U$38594 ( \46120_46420 , \45981_46281 , \45987_46287 );
and \U$38595 ( \46121_46421 , \45981_46281 , \45994_46294 );
and \U$38596 ( \46122_46422 , \45987_46287 , \45994_46294 );
or \U$38597 ( \46123_46423 , \46120_46420 , \46121_46421 , \46122_46422 );
buf \U$38598 ( \46124_46424 , \46123_46423 );
xor \U$38599 ( \46125_46425 , \46119_46419 , \46124_46424 );
buf \U$38600 ( \46126_46426 , \46125_46425 );
xor \U$38601 ( \46127_46427 , \46108_46408 , \46126_46426 );
and \U$38602 ( \46128_46428 , \45965_46265 , \45966_46266 );
and \U$38603 ( \46129_46429 , \45965_46265 , \45973_46273 );
and \U$38604 ( \46130_46430 , \45966_46266 , \45973_46273 );
or \U$38605 ( \46131_46431 , \46128_46428 , \46129_46429 , \46130_46430 );
buf \U$38606 ( \46132_46432 , \46131_46431 );
xor \U$38607 ( \46133_46433 , \46127_46427 , \46132_46432 );
buf \U$38608 ( \46134_46434 , \46133_46433 );
xor \U$38609 ( \46135_46435 , \46103_46403 , \46134_46434 );
buf \U$38610 ( \46136_46436 , \46135_46435 );
and \U$38611 ( \46137_46437 , \45960_46260 , \46004_46304 );
and \U$38612 ( \46138_46438 , \45960_46260 , \46010_46310 );
and \U$38613 ( \46139_46439 , \46004_46304 , \46010_46310 );
or \U$38614 ( \46140_46440 , \46137_46437 , \46138_46438 , \46139_46439 );
buf \U$38615 ( \46141_46441 , \46140_46440 );
xor \U$38616 ( \46142_46442 , \46136_46436 , \46141_46441 );
and \U$38617 ( \46143_46443 , \45941_46241 , \45946_46246 );
and \U$38618 ( \46144_46444 , \45941_46241 , \45952_46252 );
and \U$38619 ( \46145_46445 , \45946_46246 , \45952_46252 );
or \U$38620 ( \46146_46446 , \46143_46443 , \46144_46444 , \46145_46445 );
buf \U$38621 ( \46147_46447 , \46146_46446 );
xor \U$38622 ( \46148_46448 , \46142_46442 , \46147_46447 );
and \U$38623 ( \46149_46449 , \46032_46332 , \46148_46448 );
and \U$38625 ( \46150_46450 , \46026_46326 , \46031_46331 );
or \U$38627 ( \46151_46451 , 1'b0 , \46150_46450 , 1'b0 );
xor \U$38628 ( \46152_46452 , \46149_46449 , \46151_46451 );
and \U$38630 ( \46153_46453 , \46019_46319 , \46025_46325 );
and \U$38631 ( \46154_46454 , \46021_46321 , \46025_46325 );
or \U$38632 ( \46155_46455 , 1'b0 , \46153_46453 , \46154_46454 );
xor \U$38633 ( \46156_46456 , \46152_46452 , \46155_46455 );
xor \U$38640 ( \46157_46457 , \46156_46456 , 1'b0 );
and \U$38641 ( \46158_46458 , \46136_46436 , \46141_46441 );
and \U$38642 ( \46159_46459 , \46136_46436 , \46147_46447 );
and \U$38643 ( \46160_46460 , \46141_46441 , \46147_46447 );
or \U$38644 ( \46161_46461 , \46158_46458 , \46159_46459 , \46160_46460 );
xor \U$38645 ( \46162_46462 , \46157_46457 , \46161_46461 );
and \U$38646 ( \46163_46463 , \46097_46397 , \46102_46402 );
and \U$38647 ( \46164_46464 , \46097_46397 , \46134_46434 );
and \U$38648 ( \46165_46465 , \46102_46402 , \46134_46434 );
or \U$38649 ( \46166_46466 , \46163_46463 , \46164_46464 , \46165_46465 );
buf \U$38650 ( \46167_46467 , \46166_46466 );
and \U$38651 ( \46168_46468 , \30670_29853 , \39904_40204_nG9b72 );
and \U$38652 ( \46169_46469 , \29551_29850 , \40152_40452_nG9b6f );
or \U$38653 ( \46170_46470 , \46168_46468 , \46169_46469 );
xor \U$38654 ( \46171_46471 , \29550_29849 , \46170_46470 );
buf \U$38655 ( \46172_46472 , \46171_46471 );
buf \U$38657 ( \46173_46473 , \46172_46472 );
and \U$38658 ( \46174_46474 , \28946_28118 , \40543_40843_nG9b6c );
and \U$38659 ( \46175_46475 , \27816_28115 , \40740_41040_nG9b69 );
or \U$38660 ( \46176_46476 , \46174_46474 , \46175_46475 );
xor \U$38661 ( \46177_46477 , \27815_28114 , \46176_46476 );
buf \U$38662 ( \46178_46478 , \46177_46477 );
buf \U$38664 ( \46179_46479 , \46178_46478 );
xor \U$38665 ( \46180_46480 , \46173_46473 , \46179_46479 );
and \U$38666 ( \46181_46481 , \23495_23201 , \42133_42433_nG9b5a );
and \U$38667 ( \46182_46482 , \22899_23198 , \42466_42766_nG9b57 );
or \U$38668 ( \46183_46483 , \46181_46481 , \46182_46482 );
xor \U$38669 ( \46184_46484 , \22898_23197 , \46183_46483 );
buf \U$38670 ( \46185_46485 , \46184_46484 );
buf \U$38672 ( \46186_46486 , \46185_46485 );
xor \U$38673 ( \46187_46487 , \46180_46480 , \46186_46486 );
buf \U$38674 ( \46188_46488 , \46187_46487 );
and \U$38676 ( \46189_46489 , \32617_32916 , \39034_39334_nG9b7b );
or \U$38677 ( \46190_46490 , 1'b0 , \46189_46489 );
xor \U$38678 ( \46191_46491 , 1'b0 , \46190_46490 );
buf \U$38679 ( \46192_46492 , \46191_46491 );
buf \U$38681 ( \46193_46493 , \46192_46492 );
and \U$38682 ( \46194_46494 , \31989_31636 , \39291_39591_nG9b78 );
and \U$38683 ( \46195_46495 , \31334_31633 , \39663_39963_nG9b75 );
or \U$38684 ( \46196_46496 , \46194_46494 , \46195_46495 );
xor \U$38685 ( \46197_46497 , \31333_31632 , \46196_46496 );
buf \U$38686 ( \46198_46498 , \46197_46497 );
buf \U$38688 ( \46199_46499 , \46198_46498 );
xor \U$38689 ( \46200_46500 , \46193_46493 , \46199_46499 );
and \U$38690 ( \46201_46501 , \27141_26431 , \41081_41381_nG9b66 );
and \U$38691 ( \46202_46502 , \26129_26428 , \41385_41685_nG9b63 );
or \U$38692 ( \46203_46503 , \46201_46501 , \46202_46502 );
xor \U$38693 ( \46204_46504 , \26128_26427 , \46203_46503 );
buf \U$38694 ( \46205_46505 , \46204_46504 );
buf \U$38696 ( \46206_46506 , \46205_46505 );
xor \U$38697 ( \46207_46507 , \46200_46500 , \46206_46506 );
buf \U$38698 ( \46208_46508 , \46207_46507 );
xor \U$38699 ( \46209_46509 , \46188_46488 , \46208_46508 );
and \U$38700 ( \46210_46510 , \21908_21658 , \42548_42848_nG9b54 );
and \U$38701 ( \46211_46511 , \21356_21655 , \42879_43179_nG9b51 );
or \U$38702 ( \46212_46512 , \46210_46510 , \46211_46511 );
xor \U$38703 ( \46213_46513 , \21355_21654 , \46212_46512 );
buf \U$38704 ( \46214_46514 , \46213_46513 );
buf \U$38706 ( \46215_46515 , \46214_46514 );
xor \U$38710 ( \46216_46516 , \19852_20151 , 1'b0 );
not \U$38711 ( \46217_46517 , \46216_46516 );
buf \U$38712 ( \46218_46518 , \46217_46517 );
buf \U$38714 ( \46219_46519 , \46218_46518 );
xor \U$38715 ( \46220_46520 , \46215_46515 , \46219_46519 );
and \U$38716 ( \46221_46521 , \25044_24792 , \41663_41963_nG9b60 );
and \U$38717 ( \46222_46522 , \24490_24789 , \41901_42201_nG9b5d );
or \U$38718 ( \46223_46523 , \46221_46521 , \46222_46522 );
xor \U$38719 ( \46224_46524 , \24489_24788 , \46223_46523 );
buf \U$38720 ( \46225_46525 , \46224_46524 );
buf \U$38722 ( \46226_46526 , \46225_46525 );
xor \U$38723 ( \46227_46527 , \46220_46520 , \46226_46526 );
buf \U$38724 ( \46228_46528 , \46227_46527 );
xor \U$38725 ( \46229_46529 , \46209_46509 , \46228_46528 );
buf \U$38726 ( \46230_46530 , \46229_46529 );
and \U$38727 ( \46231_46531 , \46053_46353 , \46074_46374 );
and \U$38728 ( \46232_46532 , \46053_46353 , \46095_46395 );
and \U$38729 ( \46233_46533 , \46074_46374 , \46095_46395 );
or \U$38730 ( \46234_46534 , \46231_46531 , \46232_46532 , \46233_46533 );
buf \U$38731 ( \46235_46535 , \46234_46534 );
xor \U$38732 ( \46236_46536 , \46230_46530 , \46235_46535 );
and \U$38733 ( \46237_46537 , \46108_46408 , \46126_46426 );
and \U$38734 ( \46238_46538 , \46108_46408 , \46132_46432 );
and \U$38735 ( \46239_46539 , \46126_46426 , \46132_46432 );
or \U$38736 ( \46240_46540 , \46237_46537 , \46238_46538 , \46239_46539 );
buf \U$38737 ( \46241_46541 , \46240_46540 );
xor \U$38738 ( \46242_46542 , \46236_46536 , \46241_46541 );
buf \U$38739 ( \46243_46543 , \46242_46542 );
xor \U$38740 ( \46244_46544 , \46167_46467 , \46243_46543 );
and \U$38741 ( \46245_46545 , \46113_46413 , \46118_46418 );
and \U$38742 ( \46246_46546 , \46113_46413 , \46124_46424 );
and \U$38743 ( \46247_46547 , \46118_46418 , \46124_46424 );
or \U$38744 ( \46248_46548 , \46245_46545 , \46246_46546 , \46247_46547 );
buf \U$38745 ( \46249_46549 , \46248_46548 );
and \U$38746 ( \46250_46550 , \46080_46380 , \46086_46386 );
and \U$38747 ( \46251_46551 , \46080_46380 , \46093_46393 );
and \U$38748 ( \46252_46552 , \46086_46386 , \46093_46393 );
or \U$38749 ( \46253_46553 , \46250_46550 , \46251_46551 , \46252_46552 );
buf \U$38750 ( \46254_46554 , \46253_46553 );
and \U$38751 ( \46255_46555 , \46038_46338 , \46044_46344 );
and \U$38752 ( \46256_46556 , \46038_46338 , \46051_46351 );
and \U$38753 ( \46257_46557 , \46044_46344 , \46051_46351 );
or \U$38754 ( \46258_46558 , \46255_46555 , \46256_46556 , \46257_46557 );
buf \U$38755 ( \46259_46559 , \46258_46558 );
xor \U$38756 ( \46260_46560 , \46254_46554 , \46259_46559 );
buf \U$38757 ( \46261_46561 , \46058_46358 );
xor \U$38758 ( \46262_46562 , \46260_46560 , \46261_46561 );
buf \U$38759 ( \46263_46563 , \46262_46562 );
xor \U$38760 ( \46264_46564 , \46249_46549 , \46263_46563 );
and \U$38761 ( \46265_46565 , \46059_46359 , \46065_46365 );
and \U$38762 ( \46266_46566 , \46059_46359 , \46072_46372 );
and \U$38763 ( \46267_46567 , \46065_46365 , \46072_46372 );
or \U$38764 ( \46268_46568 , \46265_46565 , \46266_46566 , \46267_46567 );
buf \U$38765 ( \46269_46569 , \46268_46568 );
xor \U$38766 ( \46270_46570 , \46264_46564 , \46269_46569 );
buf \U$38767 ( \46271_46571 , \46270_46570 );
xor \U$38768 ( \46272_46572 , \46244_46544 , \46271_46571 );
and \U$38769 ( \46273_46573 , \46162_46462 , \46272_46572 );
and \U$38771 ( \46274_46574 , \46156_46456 , \46161_46461 );
or \U$38773 ( \46275_46575 , 1'b0 , \46274_46574 , 1'b0 );
xor \U$38774 ( \46276_46576 , \46273_46573 , \46275_46575 );
and \U$38776 ( \46277_46577 , \46149_46449 , \46155_46455 );
and \U$38777 ( \46278_46578 , \46151_46451 , \46155_46455 );
or \U$38778 ( \46279_46579 , 1'b0 , \46277_46577 , \46278_46578 );
xor \U$38779 ( \46280_46580 , \46276_46576 , \46279_46579 );
xor \U$38786 ( \46281_46581 , \46280_46580 , 1'b0 );
and \U$38787 ( \46282_46582 , \46167_46467 , \46243_46543 );
and \U$38788 ( \46283_46583 , \46167_46467 , \46271_46571 );
and \U$38789 ( \46284_46584 , \46243_46543 , \46271_46571 );
or \U$38790 ( \46285_46585 , \46282_46582 , \46283_46583 , \46284_46584 );
xor \U$38791 ( \46286_46586 , \46281_46581 , \46285_46585 );
and \U$38792 ( \46287_46587 , \46230_46530 , \46235_46535 );
and \U$38793 ( \46288_46588 , \46230_46530 , \46241_46541 );
and \U$38794 ( \46289_46589 , \46235_46535 , \46241_46541 );
or \U$38795 ( \46290_46590 , \46287_46587 , \46288_46588 , \46289_46589 );
buf \U$38796 ( \46291_46591 , \46290_46590 );
and \U$38797 ( \46292_46592 , \46188_46488 , \46208_46508 );
and \U$38798 ( \46293_46593 , \46188_46488 , \46228_46528 );
and \U$38799 ( \46294_46594 , \46208_46508 , \46228_46528 );
or \U$38800 ( \46295_46595 , \46292_46592 , \46293_46593 , \46294_46594 );
buf \U$38801 ( \46296_46596 , \46295_46595 );
and \U$38802 ( \46297_46597 , \46254_46554 , \46259_46559 );
and \U$38803 ( \46298_46598 , \46254_46554 , \46261_46561 );
and \U$38804 ( \46299_46599 , \46259_46559 , \46261_46561 );
or \U$38805 ( \46300_46600 , \46297_46597 , \46298_46598 , \46299_46599 );
buf \U$38806 ( \46301_46601 , \46300_46600 );
and \U$38807 ( \46302_46602 , \46215_46515 , \46219_46519 );
and \U$38808 ( \46303_46603 , \46215_46515 , \46226_46526 );
and \U$38809 ( \46304_46604 , \46219_46519 , \46226_46526 );
or \U$38810 ( \46305_46605 , \46302_46602 , \46303_46603 , \46304_46604 );
buf \U$38811 ( \46306_46606 , \46305_46605 );
and \U$38812 ( \46307_46607 , \21908_21658 , \42879_43179_nG9b51 );
or \U$38814 ( \46308_46608 , \46307_46607 , 1'b0 );
xor \U$38815 ( \46309_46609 , \21355_21654 , \46308_46608 );
buf \U$38816 ( \46310_46610 , \46309_46609 );
buf \U$38817 ( \46311_46611 , \46310_46610 );
not \U$38818 ( \46312_46612 , \46311_46611 );
xor \U$38819 ( \46313_46613 , \46306_46606 , \46312_46612 );
and \U$38820 ( \46314_46614 , \23495_23201 , \42466_42766_nG9b57 );
and \U$38821 ( \46315_46615 , \22899_23198 , \42548_42848_nG9b54 );
or \U$38822 ( \46316_46616 , \46314_46614 , \46315_46615 );
xor \U$38823 ( \46317_46617 , \22898_23197 , \46316_46616 );
buf \U$38824 ( \46318_46618 , \46317_46617 );
buf \U$38826 ( \46319_46619 , \46318_46618 );
xor \U$38827 ( \46320_46620 , \46313_46613 , \46319_46619 );
buf \U$38828 ( \46321_46621 , \46320_46620 );
xor \U$38829 ( \46322_46622 , \46301_46601 , \46321_46621 );
and \U$38831 ( \46323_46623 , \32617_32916 , \39291_39591_nG9b78 );
or \U$38832 ( \46324_46624 , 1'b0 , \46323_46623 );
xor \U$38833 ( \46325_46625 , 1'b0 , \46324_46624 );
buf \U$38834 ( \46326_46626 , \46325_46625 );
buf \U$38836 ( \46327_46627 , \46326_46626 );
and \U$38837 ( \46328_46628 , \28946_28118 , \40740_41040_nG9b69 );
and \U$38838 ( \46329_46629 , \27816_28115 , \41081_41381_nG9b66 );
or \U$38839 ( \46330_46630 , \46328_46628 , \46329_46629 );
xor \U$38840 ( \46331_46631 , \27815_28114 , \46330_46630 );
buf \U$38841 ( \46332_46632 , \46331_46631 );
buf \U$38843 ( \46333_46633 , \46332_46632 );
xor \U$38844 ( \46334_46634 , \46327_46627 , \46333_46633 );
and \U$38845 ( \46335_46635 , \27141_26431 , \41385_41685_nG9b63 );
and \U$38846 ( \46336_46636 , \26129_26428 , \41663_41963_nG9b60 );
or \U$38847 ( \46337_46637 , \46335_46635 , \46336_46636 );
xor \U$38848 ( \46338_46638 , \26128_26427 , \46337_46637 );
buf \U$38849 ( \46339_46639 , \46338_46638 );
buf \U$38851 ( \46340_46640 , \46339_46639 );
xor \U$38852 ( \46341_46641 , \46334_46634 , \46340_46640 );
buf \U$38853 ( \46342_46642 , \46341_46641 );
xor \U$38854 ( \46343_46643 , \46322_46622 , \46342_46642 );
buf \U$38855 ( \46344_46644 , \46343_46643 );
xor \U$38856 ( \46345_46645 , \46296_46596 , \46344_46644 );
and \U$38857 ( \46346_46646 , \46193_46493 , \46199_46499 );
and \U$38858 ( \46347_46647 , \46193_46493 , \46206_46506 );
and \U$38859 ( \46348_46648 , \46199_46499 , \46206_46506 );
or \U$38860 ( \46349_46649 , \46346_46646 , \46347_46647 , \46348_46648 );
buf \U$38861 ( \46350_46650 , \46349_46649 );
and \U$38862 ( \46351_46651 , \31989_31636 , \39663_39963_nG9b75 );
and \U$38863 ( \46352_46652 , \31334_31633 , \39904_40204_nG9b72 );
or \U$38864 ( \46353_46653 , \46351_46651 , \46352_46652 );
xor \U$38865 ( \46354_46654 , \31333_31632 , \46353_46653 );
buf \U$38866 ( \46355_46655 , \46354_46654 );
buf \U$38868 ( \46356_46656 , \46355_46655 );
and \U$38869 ( \46357_46657 , \30670_29853 , \40152_40452_nG9b6f );
and \U$38870 ( \46358_46658 , \29551_29850 , \40543_40843_nG9b6c );
or \U$38871 ( \46359_46659 , \46357_46657 , \46358_46658 );
xor \U$38872 ( \46360_46660 , \29550_29849 , \46359_46659 );
buf \U$38873 ( \46361_46661 , \46360_46660 );
buf \U$38875 ( \46362_46662 , \46361_46661 );
xor \U$38876 ( \46363_46663 , \46356_46656 , \46362_46662 );
and \U$38877 ( \46364_46664 , \25044_24792 , \41901_42201_nG9b5d );
and \U$38878 ( \46365_46665 , \24490_24789 , \42133_42433_nG9b5a );
or \U$38879 ( \46366_46666 , \46364_46664 , \46365_46665 );
xor \U$38880 ( \46367_46667 , \24489_24788 , \46366_46666 );
buf \U$38881 ( \46368_46668 , \46367_46667 );
buf \U$38883 ( \46369_46669 , \46368_46668 );
xor \U$38884 ( \46370_46670 , \46363_46663 , \46369_46669 );
buf \U$38885 ( \46371_46671 , \46370_46670 );
xor \U$38886 ( \46372_46672 , \46350_46650 , \46371_46671 );
and \U$38887 ( \46373_46673 , \46173_46473 , \46179_46479 );
and \U$38888 ( \46374_46674 , \46173_46473 , \46186_46486 );
and \U$38889 ( \46375_46675 , \46179_46479 , \46186_46486 );
or \U$38890 ( \46376_46676 , \46373_46673 , \46374_46674 , \46375_46675 );
buf \U$38891 ( \46377_46677 , \46376_46676 );
xor \U$38892 ( \46378_46678 , \46372_46672 , \46377_46677 );
buf \U$38893 ( \46379_46679 , \46378_46678 );
xor \U$38894 ( \46380_46680 , \46345_46645 , \46379_46679 );
buf \U$38895 ( \46381_46681 , \46380_46680 );
xor \U$38896 ( \46382_46682 , \46291_46591 , \46381_46681 );
and \U$38897 ( \46383_46683 , \46249_46549 , \46263_46563 );
and \U$38898 ( \46384_46684 , \46249_46549 , \46269_46569 );
and \U$38899 ( \46385_46685 , \46263_46563 , \46269_46569 );
or \U$38900 ( \46386_46686 , \46383_46683 , \46384_46684 , \46385_46685 );
buf \U$38901 ( \46387_46687 , \46386_46686 );
xor \U$38902 ( \46388_46688 , \46382_46682 , \46387_46687 );
and \U$38903 ( \46389_46689 , \46286_46586 , \46388_46688 );
and \U$38905 ( \46390_46690 , \46280_46580 , \46285_46585 );
or \U$38907 ( \46391_46691 , 1'b0 , \46390_46690 , 1'b0 );
xor \U$38908 ( \46392_46692 , \46389_46689 , \46391_46691 );
and \U$38910 ( \46393_46693 , \46273_46573 , \46279_46579 );
and \U$38911 ( \46394_46694 , \46275_46575 , \46279_46579 );
or \U$38912 ( \46395_46695 , 1'b0 , \46393_46693 , \46394_46694 );
xor \U$38913 ( \46396_46696 , \46392_46692 , \46395_46695 );
xor \U$38920 ( \46397_46697 , \46396_46696 , 1'b0 );
and \U$38921 ( \46398_46698 , \46291_46591 , \46381_46681 );
and \U$38922 ( \46399_46699 , \46291_46591 , \46387_46687 );
and \U$38923 ( \46400_46700 , \46381_46681 , \46387_46687 );
or \U$38924 ( \46401_46701 , \46398_46698 , \46399_46699 , \46400_46700 );
xor \U$38925 ( \46402_46702 , \46397_46697 , \46401_46701 );
and \U$38926 ( \46403_46703 , \46296_46596 , \46344_46644 );
and \U$38927 ( \46404_46704 , \46296_46596 , \46379_46679 );
and \U$38928 ( \46405_46705 , \46344_46644 , \46379_46679 );
or \U$38929 ( \46406_46706 , \46403_46703 , \46404_46704 , \46405_46705 );
buf \U$38930 ( \46407_46707 , \46406_46706 );
and \U$38931 ( \46408_46708 , \46301_46601 , \46321_46621 );
and \U$38932 ( \46409_46709 , \46301_46601 , \46342_46642 );
and \U$38933 ( \46410_46710 , \46321_46621 , \46342_46642 );
or \U$38934 ( \46411_46711 , \46408_46708 , \46409_46709 , \46410_46710 );
buf \U$38935 ( \46412_46712 , \46411_46711 );
and \U$38936 ( \46413_46713 , \23495_23201 , \42548_42848_nG9b54 );
and \U$38937 ( \46414_46714 , \22899_23198 , \42879_43179_nG9b51 );
or \U$38938 ( \46415_46715 , \46413_46713 , \46414_46714 );
xor \U$38939 ( \46416_46716 , \22898_23197 , \46415_46715 );
buf \U$38940 ( \46417_46717 , \46416_46716 );
buf \U$38942 ( \46418_46718 , \46417_46717 );
xor \U$38946 ( \46419_46719 , \21355_21654 , 1'b0 );
not \U$38947 ( \46420_46720 , \46419_46719 );
buf \U$38948 ( \46421_46721 , \46420_46720 );
buf \U$38950 ( \46422_46722 , \46421_46721 );
xor \U$38951 ( \46423_46723 , \46418_46718 , \46422_46722 );
and \U$38952 ( \46424_46724 , \27141_26431 , \41663_41963_nG9b60 );
and \U$38953 ( \46425_46725 , \26129_26428 , \41901_42201_nG9b5d );
or \U$38954 ( \46426_46726 , \46424_46724 , \46425_46725 );
xor \U$38955 ( \46427_46727 , \26128_26427 , \46426_46726 );
buf \U$38956 ( \46428_46728 , \46427_46727 );
buf \U$38958 ( \46429_46729 , \46428_46728 );
xor \U$38959 ( \46430_46730 , \46423_46723 , \46429_46729 );
buf \U$38960 ( \46431_46731 , \46430_46730 );
and \U$38961 ( \46432_46732 , \46356_46656 , \46362_46662 );
and \U$38962 ( \46433_46733 , \46356_46656 , \46369_46669 );
and \U$38963 ( \46434_46734 , \46362_46662 , \46369_46669 );
or \U$38964 ( \46435_46735 , \46432_46732 , \46433_46733 , \46434_46734 );
buf \U$38965 ( \46436_46736 , \46435_46735 );
xor \U$38966 ( \46437_46737 , \46431_46731 , \46436_46736 );
and \U$38967 ( \46438_46738 , \46327_46627 , \46333_46633 );
and \U$38968 ( \46439_46739 , \46327_46627 , \46340_46640 );
and \U$38969 ( \46440_46740 , \46333_46633 , \46340_46640 );
or \U$38970 ( \46441_46741 , \46438_46738 , \46439_46739 , \46440_46740 );
buf \U$38971 ( \46442_46742 , \46441_46741 );
xor \U$38972 ( \46443_46743 , \46437_46737 , \46442_46742 );
buf \U$38973 ( \46444_46744 , \46443_46743 );
xor \U$38974 ( \46445_46745 , \46412_46712 , \46444_46744 );
and \U$38975 ( \46446_46746 , \46350_46650 , \46371_46671 );
and \U$38976 ( \46447_46747 , \46350_46650 , \46377_46677 );
and \U$38977 ( \46448_46748 , \46371_46671 , \46377_46677 );
or \U$38978 ( \46449_46749 , \46446_46746 , \46447_46747 , \46448_46748 );
buf \U$38979 ( \46450_46750 , \46449_46749 );
xor \U$38980 ( \46451_46751 , \46445_46745 , \46450_46750 );
buf \U$38981 ( \46452_46752 , \46451_46751 );
xor \U$38982 ( \46453_46753 , \46407_46707 , \46452_46752 );
and \U$38983 ( \46454_46754 , \46306_46606 , \46312_46612 );
and \U$38984 ( \46455_46755 , \46306_46606 , \46319_46619 );
and \U$38985 ( \46456_46756 , \46312_46612 , \46319_46619 );
or \U$38986 ( \46457_46757 , \46454_46754 , \46455_46755 , \46456_46756 );
buf \U$38987 ( \46458_46758 , \46457_46757 );
buf \U$38988 ( \46459_46759 , \46311_46611 );
and \U$38989 ( \46460_46760 , \31989_31636 , \39904_40204_nG9b72 );
and \U$38990 ( \46461_46761 , \31334_31633 , \40152_40452_nG9b6f );
or \U$38991 ( \46462_46762 , \46460_46760 , \46461_46761 );
xor \U$38992 ( \46463_46763 , \31333_31632 , \46462_46762 );
buf \U$38993 ( \46464_46764 , \46463_46763 );
buf \U$38995 ( \46465_46765 , \46464_46764 );
xor \U$38996 ( \46466_46766 , \46459_46759 , \46465_46765 );
and \U$38997 ( \46467_46767 , \25044_24792 , \42133_42433_nG9b5a );
and \U$38998 ( \46468_46768 , \24490_24789 , \42466_42766_nG9b57 );
or \U$38999 ( \46469_46769 , \46467_46767 , \46468_46768 );
xor \U$39000 ( \46470_46770 , \24489_24788 , \46469_46769 );
buf \U$39001 ( \46471_46771 , \46470_46770 );
buf \U$39003 ( \46472_46772 , \46471_46771 );
xor \U$39004 ( \46473_46773 , \46466_46766 , \46472_46772 );
buf \U$39005 ( \46474_46774 , \46473_46773 );
xor \U$39006 ( \46475_46775 , \46458_46758 , \46474_46774 );
and \U$39008 ( \46476_46776 , \32617_32916 , \39663_39963_nG9b75 );
or \U$39009 ( \46477_46777 , 1'b0 , \46476_46776 );
xor \U$39010 ( \46478_46778 , 1'b0 , \46477_46777 );
buf \U$39011 ( \46479_46779 , \46478_46778 );
buf \U$39013 ( \46480_46780 , \46479_46779 );
and \U$39014 ( \46481_46781 , \30670_29853 , \40543_40843_nG9b6c );
and \U$39015 ( \46482_46782 , \29551_29850 , \40740_41040_nG9b69 );
or \U$39016 ( \46483_46783 , \46481_46781 , \46482_46782 );
xor \U$39017 ( \46484_46784 , \29550_29849 , \46483_46783 );
buf \U$39018 ( \46485_46785 , \46484_46784 );
buf \U$39020 ( \46486_46786 , \46485_46785 );
xor \U$39021 ( \46487_46787 , \46480_46780 , \46486_46786 );
and \U$39022 ( \46488_46788 , \28946_28118 , \41081_41381_nG9b66 );
and \U$39023 ( \46489_46789 , \27816_28115 , \41385_41685_nG9b63 );
or \U$39024 ( \46490_46790 , \46488_46788 , \46489_46789 );
xor \U$39025 ( \46491_46791 , \27815_28114 , \46490_46790 );
buf \U$39026 ( \46492_46792 , \46491_46791 );
buf \U$39028 ( \46493_46793 , \46492_46792 );
xor \U$39029 ( \46494_46794 , \46487_46787 , \46493_46793 );
buf \U$39030 ( \46495_46795 , \46494_46794 );
xor \U$39031 ( \46496_46796 , \46475_46775 , \46495_46795 );
buf \U$39032 ( \46497_46797 , \46496_46796 );
xor \U$39033 ( \46498_46798 , \46453_46753 , \46497_46797 );
and \U$39034 ( \46499_46799 , \46402_46702 , \46498_46798 );
and \U$39036 ( \46500_46800 , \46396_46696 , \46401_46701 );
or \U$39038 ( \46501_46801 , 1'b0 , \46500_46800 , 1'b0 );
xor \U$39039 ( \46502_46802 , \46499_46799 , \46501_46801 );
and \U$39041 ( \46503_46803 , \46389_46689 , \46395_46695 );
and \U$39042 ( \46504_46804 , \46391_46691 , \46395_46695 );
or \U$39043 ( \46505_46805 , 1'b0 , \46503_46803 , \46504_46804 );
xor \U$39044 ( \46506_46806 , \46502_46802 , \46505_46805 );
xor \U$39051 ( \46507_46807 , \46506_46806 , 1'b0 );
and \U$39052 ( \46508_46808 , \46407_46707 , \46452_46752 );
and \U$39053 ( \46509_46809 , \46407_46707 , \46497_46797 );
and \U$39054 ( \46510_46810 , \46452_46752 , \46497_46797 );
or \U$39055 ( \46511_46811 , \46508_46808 , \46509_46809 , \46510_46810 );
xor \U$39056 ( \46512_46812 , \46507_46807 , \46511_46811 );
and \U$39057 ( \46513_46813 , \46412_46712 , \46444_46744 );
and \U$39058 ( \46514_46814 , \46412_46712 , \46450_46750 );
and \U$39059 ( \46515_46815 , \46444_46744 , \46450_46750 );
or \U$39060 ( \46516_46816 , \46513_46813 , \46514_46814 , \46515_46815 );
buf \U$39061 ( \46517_46817 , \46516_46816 );
and \U$39062 ( \46518_46818 , \30670_29853 , \40740_41040_nG9b69 );
and \U$39063 ( \46519_46819 , \29551_29850 , \41081_41381_nG9b66 );
or \U$39064 ( \46520_46820 , \46518_46818 , \46519_46819 );
xor \U$39065 ( \46521_46821 , \29550_29849 , \46520_46820 );
buf \U$39066 ( \46522_46822 , \46521_46821 );
buf \U$39068 ( \46523_46823 , \46522_46822 );
and \U$39069 ( \46524_46824 , \28946_28118 , \41385_41685_nG9b63 );
and \U$39070 ( \46525_46825 , \27816_28115 , \41663_41963_nG9b60 );
or \U$39071 ( \46526_46826 , \46524_46824 , \46525_46825 );
xor \U$39072 ( \46527_46827 , \27815_28114 , \46526_46826 );
buf \U$39073 ( \46528_46828 , \46527_46827 );
buf \U$39075 ( \46529_46829 , \46528_46828 );
xor \U$39076 ( \46530_46830 , \46523_46823 , \46529_46829 );
and \U$39077 ( \46531_46831 , \27141_26431 , \41901_42201_nG9b5d );
and \U$39078 ( \46532_46832 , \26129_26428 , \42133_42433_nG9b5a );
or \U$39079 ( \46533_46833 , \46531_46831 , \46532_46832 );
xor \U$39080 ( \46534_46834 , \26128_26427 , \46533_46833 );
buf \U$39081 ( \46535_46835 , \46534_46834 );
buf \U$39083 ( \46536_46836 , \46535_46835 );
xor \U$39084 ( \46537_46837 , \46530_46830 , \46536_46836 );
buf \U$39085 ( \46538_46838 , \46537_46837 );
and \U$39087 ( \46539_46839 , \32617_32916 , \39904_40204_nG9b72 );
or \U$39088 ( \46540_46840 , 1'b0 , \46539_46839 );
xor \U$39089 ( \46541_46841 , 1'b0 , \46540_46840 );
buf \U$39090 ( \46542_46842 , \46541_46841 );
buf \U$39092 ( \46543_46843 , \46542_46842 );
and \U$39093 ( \46544_46844 , \31989_31636 , \40152_40452_nG9b6f );
and \U$39094 ( \46545_46845 , \31334_31633 , \40543_40843_nG9b6c );
or \U$39095 ( \46546_46846 , \46544_46844 , \46545_46845 );
xor \U$39096 ( \46547_46847 , \31333_31632 , \46546_46846 );
buf \U$39097 ( \46548_46848 , \46547_46847 );
buf \U$39099 ( \46549_46849 , \46548_46848 );
xor \U$39100 ( \46550_46850 , \46543_46843 , \46549_46849 );
and \U$39101 ( \46551_46851 , \25044_24792 , \42466_42766_nG9b57 );
and \U$39102 ( \46552_46852 , \24490_24789 , \42548_42848_nG9b54 );
or \U$39103 ( \46553_46853 , \46551_46851 , \46552_46852 );
xor \U$39104 ( \46554_46854 , \24489_24788 , \46553_46853 );
buf \U$39105 ( \46555_46855 , \46554_46854 );
buf \U$39107 ( \46556_46856 , \46555_46855 );
xor \U$39108 ( \46557_46857 , \46550_46850 , \46556_46856 );
buf \U$39109 ( \46558_46858 , \46557_46857 );
xor \U$39110 ( \46559_46859 , \46538_46838 , \46558_46858 );
and \U$39111 ( \46560_46860 , \46459_46759 , \46465_46765 );
and \U$39112 ( \46561_46861 , \46459_46759 , \46472_46772 );
and \U$39113 ( \46562_46862 , \46465_46765 , \46472_46772 );
or \U$39114 ( \46563_46863 , \46560_46860 , \46561_46861 , \46562_46862 );
buf \U$39115 ( \46564_46864 , \46563_46863 );
xor \U$39116 ( \46565_46865 , \46559_46859 , \46564_46864 );
buf \U$39117 ( \46566_46866 , \46565_46865 );
and \U$39118 ( \46567_46867 , \46431_46731 , \46436_46736 );
and \U$39119 ( \46568_46868 , \46431_46731 , \46442_46742 );
and \U$39120 ( \46569_46869 , \46436_46736 , \46442_46742 );
or \U$39121 ( \46570_46870 , \46567_46867 , \46568_46868 , \46569_46869 );
buf \U$39122 ( \46571_46871 , \46570_46870 );
xor \U$39123 ( \46572_46872 , \46566_46866 , \46571_46871 );
and \U$39124 ( \46573_46873 , \46418_46718 , \46422_46722 );
and \U$39125 ( \46574_46874 , \46418_46718 , \46429_46729 );
and \U$39126 ( \46575_46875 , \46422_46722 , \46429_46729 );
or \U$39127 ( \46576_46876 , \46573_46873 , \46574_46874 , \46575_46875 );
buf \U$39128 ( \46577_46877 , \46576_46876 );
and \U$39129 ( \46578_46878 , \46480_46780 , \46486_46786 );
and \U$39130 ( \46579_46879 , \46480_46780 , \46493_46793 );
and \U$39131 ( \46580_46880 , \46486_46786 , \46493_46793 );
or \U$39132 ( \46581_46881 , \46578_46878 , \46579_46879 , \46580_46880 );
buf \U$39133 ( \46582_46882 , \46581_46881 );
xor \U$39134 ( \46583_46883 , \46577_46877 , \46582_46882 );
and \U$39135 ( \46584_46884 , \23495_23201 , \42879_43179_nG9b51 );
or \U$39137 ( \46585_46885 , \46584_46884 , 1'b0 );
xor \U$39138 ( \46586_46886 , \22898_23197 , \46585_46885 );
buf \U$39139 ( \46587_46887 , \46586_46886 );
buf \U$39140 ( \46588_46888 , \46587_46887 );
not \U$39141 ( \46589_46889 , \46588_46888 );
xor \U$39142 ( \46590_46890 , \46583_46883 , \46589_46889 );
buf \U$39143 ( \46591_46891 , \46590_46890 );
xor \U$39144 ( \46592_46892 , \46572_46872 , \46591_46891 );
buf \U$39145 ( \46593_46893 , \46592_46892 );
xor \U$39146 ( \46594_46894 , \46517_46817 , \46593_46893 );
and \U$39147 ( \46595_46895 , \46458_46758 , \46474_46774 );
and \U$39148 ( \46596_46896 , \46458_46758 , \46495_46795 );
and \U$39149 ( \46597_46897 , \46474_46774 , \46495_46795 );
or \U$39150 ( \46598_46898 , \46595_46895 , \46596_46896 , \46597_46897 );
buf \U$39151 ( \46599_46899 , \46598_46898 );
xor \U$39152 ( \46600_46900 , \46594_46894 , \46599_46899 );
and \U$39153 ( \46601_46901 , \46512_46812 , \46600_46900 );
and \U$39155 ( \46602_46902 , \46506_46806 , \46511_46811 );
or \U$39157 ( \46603_46903 , 1'b0 , \46602_46902 , 1'b0 );
xor \U$39158 ( \46604_46904 , \46601_46901 , \46603_46903 );
and \U$39160 ( \46605_46905 , \46499_46799 , \46505_46805 );
and \U$39161 ( \46606_46906 , \46501_46801 , \46505_46805 );
or \U$39162 ( \46607_46907 , 1'b0 , \46605_46905 , \46606_46906 );
xor \U$39163 ( \46608_46908 , \46604_46904 , \46607_46907 );
xor \U$39170 ( \46609_46909 , \46608_46908 , 1'b0 );
and \U$39171 ( \46610_46910 , \46517_46817 , \46593_46893 );
and \U$39172 ( \46611_46911 , \46517_46817 , \46599_46899 );
and \U$39173 ( \46612_46912 , \46593_46893 , \46599_46899 );
or \U$39174 ( \46613_46913 , \46610_46910 , \46611_46911 , \46612_46912 );
xor \U$39175 ( \46614_46914 , \46609_46909 , \46613_46913 );
and \U$39176 ( \46615_46915 , \46566_46866 , \46571_46871 );
and \U$39177 ( \46616_46916 , \46566_46866 , \46591_46891 );
and \U$39178 ( \46617_46917 , \46571_46871 , \46591_46891 );
or \U$39179 ( \46618_46918 , \46615_46915 , \46616_46916 , \46617_46917 );
buf \U$39180 ( \46619_46919 , \46618_46918 );
and \U$39181 ( \46620_46920 , \46538_46838 , \46558_46858 );
and \U$39182 ( \46621_46921 , \46538_46838 , \46564_46864 );
and \U$39183 ( \46622_46922 , \46558_46858 , \46564_46864 );
or \U$39184 ( \46623_46923 , \46620_46920 , \46621_46921 , \46622_46922 );
buf \U$39185 ( \46624_46924 , \46623_46923 );
and \U$39186 ( \46625_46925 , \46577_46877 , \46582_46882 );
and \U$39187 ( \46626_46926 , \46577_46877 , \46589_46889 );
and \U$39188 ( \46627_46927 , \46582_46882 , \46589_46889 );
or \U$39189 ( \46628_46928 , \46625_46925 , \46626_46926 , \46627_46927 );
buf \U$39190 ( \46629_46929 , \46628_46928 );
xor \U$39191 ( \46630_46930 , \46624_46924 , \46629_46929 );
and \U$39192 ( \46631_46931 , \46523_46823 , \46529_46829 );
and \U$39193 ( \46632_46932 , \46523_46823 , \46536_46836 );
and \U$39194 ( \46633_46933 , \46529_46829 , \46536_46836 );
or \U$39195 ( \46634_46934 , \46631_46931 , \46632_46932 , \46633_46933 );
buf \U$39196 ( \46635_46935 , \46634_46934 );
buf \U$39197 ( \46636_46936 , \46588_46888 );
xor \U$39198 ( \46637_46937 , \46635_46935 , \46636_46936 );
and \U$39199 ( \46638_46938 , \27141_26431 , \42133_42433_nG9b5a );
and \U$39200 ( \46639_46939 , \26129_26428 , \42466_42766_nG9b57 );
or \U$39201 ( \46640_46940 , \46638_46938 , \46639_46939 );
xor \U$39202 ( \46641_46941 , \26128_26427 , \46640_46940 );
buf \U$39203 ( \46642_46942 , \46641_46941 );
buf \U$39205 ( \46643_46943 , \46642_46942 );
xor \U$39206 ( \46644_46944 , \46637_46937 , \46643_46943 );
buf \U$39207 ( \46645_46945 , \46644_46944 );
xor \U$39208 ( \46646_46946 , \46630_46930 , \46645_46945 );
buf \U$39209 ( \46647_46947 , \46646_46946 );
xor \U$39210 ( \46648_46948 , \46619_46919 , \46647_46947 );
and \U$39212 ( \46649_46949 , \32617_32916 , \40152_40452_nG9b6f );
or \U$39213 ( \46650_46950 , 1'b0 , \46649_46949 );
xor \U$39214 ( \46651_46951 , 1'b0 , \46650_46950 );
buf \U$39215 ( \46652_46952 , \46651_46951 );
buf \U$39217 ( \46653_46953 , \46652_46952 );
and \U$39218 ( \46654_46954 , \31989_31636 , \40543_40843_nG9b6c );
and \U$39219 ( \46655_46955 , \31334_31633 , \40740_41040_nG9b69 );
or \U$39220 ( \46656_46956 , \46654_46954 , \46655_46955 );
xor \U$39221 ( \46657_46957 , \31333_31632 , \46656_46956 );
buf \U$39222 ( \46658_46958 , \46657_46957 );
buf \U$39224 ( \46659_46959 , \46658_46958 );
xor \U$39225 ( \46660_46960 , \46653_46953 , \46659_46959 );
and \U$39226 ( \46661_46961 , \30670_29853 , \41081_41381_nG9b66 );
and \U$39227 ( \46662_46962 , \29551_29850 , \41385_41685_nG9b63 );
or \U$39228 ( \46663_46963 , \46661_46961 , \46662_46962 );
xor \U$39229 ( \46664_46964 , \29550_29849 , \46663_46963 );
buf \U$39230 ( \46665_46965 , \46664_46964 );
buf \U$39232 ( \46666_46966 , \46665_46965 );
xor \U$39233 ( \46667_46967 , \46660_46960 , \46666_46966 );
buf \U$39234 ( \46668_46968 , \46667_46967 );
and \U$39235 ( \46669_46969 , \25044_24792 , \42548_42848_nG9b54 );
and \U$39236 ( \46670_46970 , \24490_24789 , \42879_43179_nG9b51 );
or \U$39237 ( \46671_46971 , \46669_46969 , \46670_46970 );
xor \U$39238 ( \46672_46972 , \24489_24788 , \46671_46971 );
buf \U$39239 ( \46673_46973 , \46672_46972 );
buf \U$39241 ( \46674_46974 , \46673_46973 );
xor \U$39245 ( \46675_46975 , \22898_23197 , 1'b0 );
not \U$39246 ( \46676_46976 , \46675_46975 );
buf \U$39247 ( \46677_46977 , \46676_46976 );
buf \U$39249 ( \46678_46978 , \46677_46977 );
xor \U$39250 ( \46679_46979 , \46674_46974 , \46678_46978 );
and \U$39251 ( \46680_46980 , \28946_28118 , \41663_41963_nG9b60 );
and \U$39252 ( \46681_46981 , \27816_28115 , \41901_42201_nG9b5d );
or \U$39253 ( \46682_46982 , \46680_46980 , \46681_46981 );
xor \U$39254 ( \46683_46983 , \27815_28114 , \46682_46982 );
buf \U$39255 ( \46684_46984 , \46683_46983 );
buf \U$39257 ( \46685_46985 , \46684_46984 );
xor \U$39258 ( \46686_46986 , \46679_46979 , \46685_46985 );
buf \U$39259 ( \46687_46987 , \46686_46986 );
xor \U$39260 ( \46688_46988 , \46668_46968 , \46687_46987 );
and \U$39261 ( \46689_46989 , \46543_46843 , \46549_46849 );
and \U$39262 ( \46690_46990 , \46543_46843 , \46556_46856 );
and \U$39263 ( \46691_46991 , \46549_46849 , \46556_46856 );
or \U$39264 ( \46692_46992 , \46689_46989 , \46690_46990 , \46691_46991 );
buf \U$39265 ( \46693_46993 , \46692_46992 );
xor \U$39266 ( \46694_46994 , \46688_46988 , \46693_46993 );
buf \U$39267 ( \46695_46995 , \46694_46994 );
xor \U$39268 ( \46696_46996 , \46648_46948 , \46695_46995 );
and \U$39269 ( \46697_46997 , \46614_46914 , \46696_46996 );
and \U$39271 ( \46698_46998 , \46608_46908 , \46613_46913 );
or \U$39273 ( \46699_46999 , 1'b0 , \46698_46998 , 1'b0 );
xor \U$39274 ( \46700_47000 , \46697_46997 , \46699_46999 );
and \U$39276 ( \46701_47001 , \46601_46901 , \46607_46907 );
and \U$39277 ( \46702_47002 , \46603_46903 , \46607_46907 );
or \U$39278 ( \46703_47003 , 1'b0 , \46701_47001 , \46702_47002 );
xor \U$39279 ( \46704_47004 , \46700_47000 , \46703_47003 );
xor \U$39286 ( \46705_47005 , \46704_47004 , 1'b0 );
and \U$39287 ( \46706_47006 , \46619_46919 , \46647_46947 );
and \U$39288 ( \46707_47007 , \46619_46919 , \46695_46995 );
and \U$39289 ( \46708_47008 , \46647_46947 , \46695_46995 );
or \U$39290 ( \46709_47009 , \46706_47006 , \46707_47007 , \46708_47008 );
xor \U$39291 ( \46710_47010 , \46705_47005 , \46709_47009 );
and \U$39292 ( \46711_47011 , \46624_46924 , \46629_46929 );
and \U$39293 ( \46712_47012 , \46624_46924 , \46645_46945 );
and \U$39294 ( \46713_47013 , \46629_46929 , \46645_46945 );
or \U$39295 ( \46714_47014 , \46711_47011 , \46712_47012 , \46713_47013 );
buf \U$39296 ( \46715_47015 , \46714_47014 );
and \U$39297 ( \46716_47016 , \46668_46968 , \46687_46987 );
and \U$39298 ( \46717_47017 , \46668_46968 , \46693_46993 );
and \U$39299 ( \46718_47018 , \46687_46987 , \46693_46993 );
or \U$39300 ( \46719_47019 , \46716_47016 , \46717_47017 , \46718_47018 );
buf \U$39301 ( \46720_47020 , \46719_47019 );
and \U$39302 ( \46721_47021 , \46635_46935 , \46636_46936 );
and \U$39303 ( \46722_47022 , \46635_46935 , \46643_46943 );
and \U$39304 ( \46723_47023 , \46636_46936 , \46643_46943 );
or \U$39305 ( \46724_47024 , \46721_47021 , \46722_47022 , \46723_47023 );
buf \U$39306 ( \46725_47025 , \46724_47024 );
xor \U$39307 ( \46726_47026 , \46720_47020 , \46725_47025 );
and \U$39308 ( \46727_47027 , \30670_29853 , \41385_41685_nG9b63 );
and \U$39309 ( \46728_47028 , \29551_29850 , \41663_41963_nG9b60 );
or \U$39310 ( \46729_47029 , \46727_47027 , \46728_47028 );
xor \U$39311 ( \46730_47030 , \29550_29849 , \46729_47029 );
buf \U$39312 ( \46731_47031 , \46730_47030 );
buf \U$39313 ( \46732_47032 , \46731_47031 );
not \U$39314 ( \46733_47033 , \46732_47032 );
and \U$39315 ( \46734_47034 , \28946_28118 , \41901_42201_nG9b5d );
and \U$39316 ( \46735_47035 , \27816_28115 , \42133_42433_nG9b5a );
or \U$39317 ( \46736_47036 , \46734_47034 , \46735_47035 );
xor \U$39318 ( \46737_47037 , \27815_28114 , \46736_47036 );
buf \U$39319 ( \46738_47038 , \46737_47037 );
buf \U$39321 ( \46739_47039 , \46738_47038 );
xor \U$39322 ( \46740_47040 , \46733_47033 , \46739_47039 );
and \U$39323 ( \46741_47041 , \27141_26431 , \42466_42766_nG9b57 );
and \U$39324 ( \46742_47042 , \26129_26428 , \42548_42848_nG9b54 );
or \U$39325 ( \46743_47043 , \46741_47041 , \46742_47042 );
xor \U$39326 ( \46744_47044 , \26128_26427 , \46743_47043 );
buf \U$39327 ( \46745_47045 , \46744_47044 );
buf \U$39329 ( \46746_47046 , \46745_47045 );
xor \U$39330 ( \46747_47047 , \46740_47040 , \46746_47046 );
buf \U$39331 ( \46748_47048 , \46747_47047 );
xor \U$39332 ( \46749_47049 , \46726_47026 , \46748_47048 );
buf \U$39333 ( \46750_47050 , \46749_47049 );
xor \U$39334 ( \46751_47051 , \46715_47015 , \46750_47050 );
and \U$39335 ( \46752_47052 , \46674_46974 , \46678_46978 );
and \U$39336 ( \46753_47053 , \46674_46974 , \46685_46985 );
and \U$39337 ( \46754_47054 , \46678_46978 , \46685_46985 );
or \U$39338 ( \46755_47055 , \46752_47052 , \46753_47053 , \46754_47054 );
buf \U$39339 ( \46756_47056 , \46755_47055 );
and \U$39340 ( \46757_47057 , \25044_24792 , \42879_43179_nG9b51 );
or \U$39342 ( \46758_47058 , \46757_47057 , 1'b0 );
xor \U$39343 ( \46759_47059 , \24489_24788 , \46758_47058 );
buf \U$39344 ( \46760_47060 , \46759_47059 );
buf \U$39346 ( \46761_47061 , \46760_47060 );
and \U$39348 ( \46762_47062 , \32617_32916 , \40543_40843_nG9b6c );
or \U$39349 ( \46763_47063 , 1'b0 , \46762_47062 );
xor \U$39350 ( \46764_47064 , 1'b0 , \46763_47063 );
buf \U$39351 ( \46765_47065 , \46764_47064 );
buf \U$39353 ( \46766_47066 , \46765_47065 );
xor \U$39354 ( \46767_47067 , \46761_47061 , \46766_47066 );
and \U$39355 ( \46768_47068 , \31989_31636 , \40740_41040_nG9b69 );
and \U$39356 ( \46769_47069 , \31334_31633 , \41081_41381_nG9b66 );
or \U$39357 ( \46770_47070 , \46768_47068 , \46769_47069 );
xor \U$39358 ( \46771_47071 , \31333_31632 , \46770_47070 );
buf \U$39359 ( \46772_47072 , \46771_47071 );
buf \U$39361 ( \46773_47073 , \46772_47072 );
xor \U$39362 ( \46774_47074 , \46767_47067 , \46773_47073 );
buf \U$39363 ( \46775_47075 , \46774_47074 );
xor \U$39364 ( \46776_47076 , \46756_47056 , \46775_47075 );
and \U$39365 ( \46777_47077 , \46653_46953 , \46659_46959 );
and \U$39366 ( \46778_47078 , \46653_46953 , \46666_46966 );
and \U$39367 ( \46779_47079 , \46659_46959 , \46666_46966 );
or \U$39368 ( \46780_47080 , \46777_47077 , \46778_47078 , \46779_47079 );
buf \U$39369 ( \46781_47081 , \46780_47080 );
xor \U$39370 ( \46782_47082 , \46776_47076 , \46781_47081 );
buf \U$39371 ( \46783_47083 , \46782_47082 );
xor \U$39372 ( \46784_47084 , \46751_47051 , \46783_47083 );
and \U$39373 ( \46785_47085 , \46710_47010 , \46784_47084 );
and \U$39375 ( \46786_47086 , \46704_47004 , \46709_47009 );
or \U$39377 ( \46787_47087 , 1'b0 , \46786_47086 , 1'b0 );
xor \U$39378 ( \46788_47088 , \46785_47085 , \46787_47087 );
and \U$39380 ( \46789_47089 , \46697_46997 , \46703_47003 );
and \U$39381 ( \46790_47090 , \46699_46999 , \46703_47003 );
or \U$39382 ( \46791_47091 , 1'b0 , \46789_47089 , \46790_47090 );
xor \U$39383 ( \46792_47092 , \46788_47088 , \46791_47091 );
xor \U$39390 ( \46793_47093 , \46792_47092 , 1'b0 );
and \U$39391 ( \46794_47094 , \27141_26431 , \42548_42848_nG9b54 );
and \U$39392 ( \46795_47095 , \26129_26428 , \42879_43179_nG9b51 );
or \U$39393 ( \46796_47096 , \46794_47094 , \46795_47095 );
xor \U$39394 ( \46797_47097 , \26128_26427 , \46796_47096 );
buf \U$39395 ( \46798_47098 , \46797_47097 );
buf \U$39397 ( \46799_47099 , \46798_47098 );
xor \U$39401 ( \46800_47100 , \24489_24788 , 1'b0 );
not \U$39402 ( \46801_47101 , \46800_47100 );
buf \U$39403 ( \46802_47102 , \46801_47101 );
buf \U$39405 ( \46803_47103 , \46802_47102 );
xor \U$39406 ( \46804_47104 , \46799_47099 , \46803_47103 );
and \U$39407 ( \46805_47105 , \30670_29853 , \41663_41963_nG9b60 );
and \U$39408 ( \46806_47106 , \29551_29850 , \41901_42201_nG9b5d );
or \U$39409 ( \46807_47107 , \46805_47105 , \46806_47106 );
xor \U$39410 ( \46808_47108 , \29550_29849 , \46807_47107 );
buf \U$39411 ( \46809_47109 , \46808_47108 );
buf \U$39413 ( \46810_47110 , \46809_47109 );
xor \U$39414 ( \46811_47111 , \46804_47104 , \46810_47110 );
buf \U$39415 ( \46812_47112 , \46811_47111 );
and \U$39416 ( \46813_47113 , \46733_47033 , \46739_47039 );
and \U$39417 ( \46814_47114 , \46733_47033 , \46746_47046 );
and \U$39418 ( \46815_47115 , \46739_47039 , \46746_47046 );
or \U$39419 ( \46816_47116 , \46813_47113 , \46814_47114 , \46815_47115 );
buf \U$39420 ( \46817_47117 , \46816_47116 );
xor \U$39421 ( \46818_47118 , \46812_47112 , \46817_47117 );
and \U$39422 ( \46819_47119 , \46761_47061 , \46766_47066 );
and \U$39423 ( \46820_47120 , \46761_47061 , \46773_47073 );
and \U$39424 ( \46821_47121 , \46766_47066 , \46773_47073 );
or \U$39425 ( \46822_47122 , \46819_47119 , \46820_47120 , \46821_47121 );
buf \U$39426 ( \46823_47123 , \46822_47122 );
and \U$39428 ( \46824_47124 , \32617_32916 , \40740_41040_nG9b69 );
or \U$39429 ( \46825_47125 , 1'b0 , \46824_47124 );
xor \U$39430 ( \46826_47126 , 1'b0 , \46825_47125 );
buf \U$39431 ( \46827_47127 , \46826_47126 );
buf \U$39433 ( \46828_47128 , \46827_47127 );
and \U$39434 ( \46829_47129 , \31989_31636 , \41081_41381_nG9b66 );
and \U$39435 ( \46830_47130 , \31334_31633 , \41385_41685_nG9b63 );
or \U$39436 ( \46831_47131 , \46829_47129 , \46830_47130 );
xor \U$39437 ( \46832_47132 , \31333_31632 , \46831_47131 );
buf \U$39438 ( \46833_47133 , \46832_47132 );
buf \U$39440 ( \46834_47134 , \46833_47133 );
xor \U$39441 ( \46835_47135 , \46828_47128 , \46834_47134 );
and \U$39442 ( \46836_47136 , \28946_28118 , \42133_42433_nG9b5a );
and \U$39443 ( \46837_47137 , \27816_28115 , \42466_42766_nG9b57 );
or \U$39444 ( \46838_47138 , \46836_47136 , \46837_47137 );
xor \U$39445 ( \46839_47139 , \27815_28114 , \46838_47138 );
buf \U$39446 ( \46840_47140 , \46839_47139 );
buf \U$39448 ( \46841_47141 , \46840_47140 );
xor \U$39449 ( \46842_47142 , \46835_47135 , \46841_47141 );
buf \U$39450 ( \46843_47143 , \46842_47142 );
xor \U$39451 ( \46844_47144 , \46823_47123 , \46843_47143 );
buf \U$39452 ( \46845_47145 , \46732_47032 );
xor \U$39453 ( \46846_47146 , \46844_47144 , \46845_47145 );
buf \U$39454 ( \46847_47147 , \46846_47146 );
xor \U$39455 ( \46848_47148 , \46818_47118 , \46847_47147 );
buf \U$39456 ( \46849_47149 , \46848_47148 );
and \U$39457 ( \46850_47150 , \46720_47020 , \46725_47025 );
and \U$39458 ( \46851_47151 , \46720_47020 , \46748_47048 );
and \U$39459 ( \46852_47152 , \46725_47025 , \46748_47048 );
or \U$39460 ( \46853_47153 , \46850_47150 , \46851_47151 , \46852_47152 );
buf \U$39461 ( \46854_47154 , \46853_47153 );
xor \U$39462 ( \46855_47155 , \46849_47149 , \46854_47154 );
and \U$39463 ( \46856_47156 , \46756_47056 , \46775_47075 );
and \U$39464 ( \46857_47157 , \46756_47056 , \46781_47081 );
and \U$39465 ( \46858_47158 , \46775_47075 , \46781_47081 );
or \U$39466 ( \46859_47159 , \46856_47156 , \46857_47157 , \46858_47158 );
buf \U$39467 ( \46860_47160 , \46859_47159 );
xor \U$39468 ( \46861_47161 , \46855_47155 , \46860_47160 );
xor \U$39469 ( \46862_47162 , \46793_47093 , \46861_47161 );
and \U$39470 ( \46863_47163 , \46715_47015 , \46750_47050 );
and \U$39471 ( \46864_47164 , \46715_47015 , \46783_47083 );
and \U$39472 ( \46865_47165 , \46750_47050 , \46783_47083 );
or \U$39473 ( \46866_47166 , \46863_47163 , \46864_47164 , \46865_47165 );
and \U$39474 ( \46867_47167 , \46862_47162 , \46866_47166 );
and \U$39476 ( \46868_47168 , \46792_47092 , \46861_47161 );
or \U$39478 ( \46869_47169 , 1'b0 , \46868_47168 , 1'b0 );
xor \U$39479 ( \46870_47170 , \46867_47167 , \46869_47169 );
and \U$39481 ( \46871_47171 , \46785_47085 , \46791_47091 );
and \U$39482 ( \46872_47172 , \46787_47087 , \46791_47091 );
or \U$39483 ( \46873_47173 , 1'b0 , \46871_47171 , \46872_47172 );
xor \U$39484 ( \46874_47174 , \46870_47170 , \46873_47173 );
xor \U$39491 ( \46875_47175 , \46874_47174 , 1'b0 );
and \U$39492 ( \46876_47176 , \46812_47112 , \46817_47117 );
and \U$39493 ( \46877_47177 , \46812_47112 , \46847_47147 );
and \U$39494 ( \46878_47178 , \46817_47117 , \46847_47147 );
or \U$39495 ( \46879_47179 , \46876_47176 , \46877_47177 , \46878_47178 );
buf \U$39496 ( \46880_47180 , \46879_47179 );
and \U$39497 ( \46881_47181 , \46799_47099 , \46803_47103 );
and \U$39498 ( \46882_47182 , \46799_47099 , \46810_47110 );
and \U$39499 ( \46883_47183 , \46803_47103 , \46810_47110 );
or \U$39500 ( \46884_47184 , \46881_47181 , \46882_47182 , \46883_47183 );
buf \U$39501 ( \46885_47185 , \46884_47184 );
and \U$39502 ( \46886_47186 , \31989_31636 , \41385_41685_nG9b63 );
and \U$39503 ( \46887_47187 , \31334_31633 , \41663_41963_nG9b60 );
or \U$39504 ( \46888_47188 , \46886_47186 , \46887_47187 );
xor \U$39505 ( \46889_47189 , \31333_31632 , \46888_47188 );
buf \U$39506 ( \46890_47190 , \46889_47189 );
buf \U$39507 ( \46891_47191 , \46890_47190 );
not \U$39508 ( \46892_47192 , \46891_47191 );
xor \U$39509 ( \46893_47193 , \46885_47185 , \46892_47192 );
and \U$39510 ( \46894_47194 , \28946_28118 , \42466_42766_nG9b57 );
and \U$39511 ( \46895_47195 , \27816_28115 , \42548_42848_nG9b54 );
or \U$39512 ( \46896_47196 , \46894_47194 , \46895_47195 );
xor \U$39513 ( \46897_47197 , \27815_28114 , \46896_47196 );
buf \U$39514 ( \46898_47198 , \46897_47197 );
buf \U$39516 ( \46899_47199 , \46898_47198 );
xor \U$39517 ( \46900_47200 , \46893_47193 , \46899_47199 );
buf \U$39518 ( \46901_47201 , \46900_47200 );
and \U$39519 ( \46902_47202 , \27141_26431 , \42879_43179_nG9b51 );
or \U$39521 ( \46903_47203 , \46902_47202 , 1'b0 );
xor \U$39522 ( \46904_47204 , \26128_26427 , \46903_47203 );
buf \U$39523 ( \46905_47205 , \46904_47204 );
buf \U$39525 ( \46906_47206 , \46905_47205 );
and \U$39527 ( \46907_47207 , \32617_32916 , \41081_41381_nG9b66 );
or \U$39528 ( \46908_47208 , 1'b0 , \46907_47207 );
xor \U$39529 ( \46909_47209 , 1'b0 , \46908_47208 );
buf \U$39530 ( \46910_47210 , \46909_47209 );
buf \U$39532 ( \46911_47211 , \46910_47210 );
xor \U$39533 ( \46912_47212 , \46906_47206 , \46911_47211 );
and \U$39534 ( \46913_47213 , \30670_29853 , \41901_42201_nG9b5d );
and \U$39535 ( \46914_47214 , \29551_29850 , \42133_42433_nG9b5a );
or \U$39536 ( \46915_47215 , \46913_47213 , \46914_47214 );
xor \U$39537 ( \46916_47216 , \29550_29849 , \46915_47215 );
buf \U$39538 ( \46917_47217 , \46916_47216 );
buf \U$39540 ( \46918_47218 , \46917_47217 );
xor \U$39541 ( \46919_47219 , \46912_47212 , \46918_47218 );
buf \U$39542 ( \46920_47220 , \46919_47219 );
xor \U$39543 ( \46921_47221 , \46901_47201 , \46920_47220 );
and \U$39544 ( \46922_47222 , \46828_47128 , \46834_47134 );
and \U$39545 ( \46923_47223 , \46828_47128 , \46841_47141 );
and \U$39546 ( \46924_47224 , \46834_47134 , \46841_47141 );
or \U$39547 ( \46925_47225 , \46922_47222 , \46923_47223 , \46924_47224 );
buf \U$39548 ( \46926_47226 , \46925_47225 );
xor \U$39549 ( \46927_47227 , \46921_47221 , \46926_47226 );
buf \U$39550 ( \46928_47228 , \46927_47227 );
xor \U$39551 ( \46929_47229 , \46880_47180 , \46928_47228 );
and \U$39552 ( \46930_47230 , \46823_47123 , \46843_47143 );
and \U$39553 ( \46931_47231 , \46823_47123 , \46845_47145 );
and \U$39554 ( \46932_47232 , \46843_47143 , \46845_47145 );
or \U$39555 ( \46933_47233 , \46930_47230 , \46931_47231 , \46932_47232 );
buf \U$39556 ( \46934_47234 , \46933_47233 );
xor \U$39557 ( \46935_47235 , \46929_47229 , \46934_47234 );
xor \U$39558 ( \46936_47236 , \46875_47175 , \46935_47235 );
and \U$39559 ( \46937_47237 , \46849_47149 , \46854_47154 );
and \U$39560 ( \46938_47238 , \46849_47149 , \46860_47160 );
and \U$39561 ( \46939_47239 , \46854_47154 , \46860_47160 );
or \U$39562 ( \46940_47240 , \46937_47237 , \46938_47238 , \46939_47239 );
and \U$39563 ( \46941_47241 , \46936_47236 , \46940_47240 );
and \U$39565 ( \46942_47242 , \46874_47174 , \46935_47235 );
or \U$39567 ( \46943_47243 , 1'b0 , \46942_47242 , 1'b0 );
xor \U$39568 ( \46944_47244 , \46941_47241 , \46943_47243 );
and \U$39570 ( \46945_47245 , \46867_47167 , \46873_47173 );
and \U$39571 ( \46946_47246 , \46869_47169 , \46873_47173 );
or \U$39572 ( \46947_47247 , 1'b0 , \46945_47245 , \46946_47246 );
xor \U$39573 ( \46948_47248 , \46944_47244 , \46947_47247 );
xor \U$39580 ( \46949_47249 , \46948_47248 , 1'b0 );
and \U$39581 ( \46950_47250 , \46880_47180 , \46928_47228 );
and \U$39582 ( \46951_47251 , \46880_47180 , \46934_47234 );
and \U$39583 ( \46952_47252 , \46928_47228 , \46934_47234 );
or \U$39584 ( \46953_47253 , \46950_47250 , \46951_47251 , \46952_47252 );
xor \U$39585 ( \46954_47254 , \46949_47249 , \46953_47253 );
and \U$39586 ( \46955_47255 , \46885_47185 , \46892_47192 );
and \U$39587 ( \46956_47256 , \46885_47185 , \46899_47199 );
and \U$39588 ( \46957_47257 , \46892_47192 , \46899_47199 );
or \U$39589 ( \46958_47258 , \46955_47255 , \46956_47256 , \46957_47257 );
buf \U$39590 ( \46959_47259 , \46958_47258 );
and \U$39592 ( \46960_47260 , \32617_32916 , \41385_41685_nG9b63 );
or \U$39593 ( \46961_47261 , 1'b0 , \46960_47260 );
xor \U$39594 ( \46962_47262 , 1'b0 , \46961_47261 );
buf \U$39595 ( \46963_47263 , \46962_47262 );
buf \U$39597 ( \46964_47264 , \46963_47263 );
buf \U$39598 ( \46965_47265 , \46891_47191 );
xor \U$39599 ( \46966_47266 , \46964_47264 , \46965_47265 );
and \U$39600 ( \46967_47267 , \30670_29853 , \42133_42433_nG9b5a );
and \U$39601 ( \46968_47268 , \29551_29850 , \42466_42766_nG9b57 );
or \U$39602 ( \46969_47269 , \46967_47267 , \46968_47268 );
xor \U$39603 ( \46970_47270 , \29550_29849 , \46969_47269 );
buf \U$39604 ( \46971_47271 , \46970_47270 );
buf \U$39606 ( \46972_47272 , \46971_47271 );
xor \U$39607 ( \46973_47273 , \46966_47266 , \46972_47272 );
buf \U$39608 ( \46974_47274 , \46973_47273 );
and \U$39609 ( \46975_47275 , \28946_28118 , \42548_42848_nG9b54 );
and \U$39610 ( \46976_47276 , \27816_28115 , \42879_43179_nG9b51 );
or \U$39611 ( \46977_47277 , \46975_47275 , \46976_47276 );
xor \U$39612 ( \46978_47278 , \27815_28114 , \46977_47277 );
buf \U$39613 ( \46979_47279 , \46978_47278 );
buf \U$39615 ( \46980_47280 , \46979_47279 );
xor \U$39619 ( \46981_47281 , \26128_26427 , 1'b0 );
not \U$39620 ( \46982_47282 , \46981_47281 );
buf \U$39621 ( \46983_47283 , \46982_47282 );
buf \U$39623 ( \46984_47284 , \46983_47283 );
xor \U$39624 ( \46985_47285 , \46980_47280 , \46984_47284 );
and \U$39625 ( \46986_47286 , \31989_31636 , \41663_41963_nG9b60 );
and \U$39626 ( \46987_47287 , \31334_31633 , \41901_42201_nG9b5d );
or \U$39627 ( \46988_47288 , \46986_47286 , \46987_47287 );
xor \U$39628 ( \46989_47289 , \31333_31632 , \46988_47288 );
buf \U$39629 ( \46990_47290 , \46989_47289 );
buf \U$39631 ( \46991_47291 , \46990_47290 );
xor \U$39632 ( \46992_47292 , \46985_47285 , \46991_47291 );
buf \U$39633 ( \46993_47293 , \46992_47292 );
xor \U$39634 ( \46994_47294 , \46974_47274 , \46993_47293 );
and \U$39635 ( \46995_47295 , \46906_47206 , \46911_47211 );
and \U$39636 ( \46996_47296 , \46906_47206 , \46918_47218 );
and \U$39637 ( \46997_47297 , \46911_47211 , \46918_47218 );
or \U$39638 ( \46998_47298 , \46995_47295 , \46996_47296 , \46997_47297 );
buf \U$39639 ( \46999_47299 , \46998_47298 );
xor \U$39640 ( \47000_47300 , \46994_47294 , \46999_47299 );
buf \U$39641 ( \47001_47301 , \47000_47300 );
xor \U$39642 ( \47002_47302 , \46959_47259 , \47001_47301 );
and \U$39643 ( \47003_47303 , \46901_47201 , \46920_47220 );
and \U$39644 ( \47004_47304 , \46901_47201 , \46926_47226 );
and \U$39645 ( \47005_47305 , \46920_47220 , \46926_47226 );
or \U$39646 ( \47006_47306 , \47003_47303 , \47004_47304 , \47005_47305 );
buf \U$39647 ( \47007_47307 , \47006_47306 );
xor \U$39648 ( \47008_47308 , \47002_47302 , \47007_47307 );
and \U$39649 ( \47009_47309 , \46954_47254 , \47008_47308 );
and \U$39651 ( \47010_47310 , \46948_47248 , \46953_47253 );
or \U$39653 ( \47011_47311 , 1'b0 , \47010_47310 , 1'b0 );
xor \U$39654 ( \47012_47312 , \47009_47309 , \47011_47311 );
and \U$39656 ( \47013_47313 , \46941_47241 , \46947_47247 );
and \U$39657 ( \47014_47314 , \46943_47243 , \46947_47247 );
or \U$39658 ( \47015_47315 , 1'b0 , \47013_47313 , \47014_47314 );
xor \U$39659 ( \47016_47316 , \47012_47312 , \47015_47315 );
xor \U$39666 ( \47017_47317 , \47016_47316 , 1'b0 );
and \U$39667 ( \47018_47318 , \46974_47274 , \46993_47293 );
and \U$39668 ( \47019_47319 , \46974_47274 , \46999_47299 );
and \U$39669 ( \47020_47320 , \46993_47293 , \46999_47299 );
or \U$39670 ( \47021_47321 , \47018_47318 , \47019_47319 , \47020_47320 );
buf \U$39671 ( \47022_47322 , \47021_47321 );
and \U$39672 ( \47023_47323 , \46980_47280 , \46984_47284 );
and \U$39673 ( \47024_47324 , \46980_47280 , \46991_47291 );
and \U$39674 ( \47025_47325 , \46984_47284 , \46991_47291 );
or \U$39675 ( \47026_47326 , \47023_47323 , \47024_47324 , \47025_47325 );
buf \U$39676 ( \47027_47327 , \47026_47326 );
and \U$39678 ( \47028_47328 , \32617_32916 , \41663_41963_nG9b60 );
or \U$39679 ( \47029_47329 , 1'b0 , \47028_47328 );
xor \U$39680 ( \47030_47330 , 1'b0 , \47029_47329 );
buf \U$39681 ( \47031_47331 , \47030_47330 );
buf \U$39683 ( \47032_47332 , \47031_47331 );
and \U$39684 ( \47033_47333 , \31989_31636 , \41901_42201_nG9b5d );
and \U$39685 ( \47034_47334 , \31334_31633 , \42133_42433_nG9b5a );
or \U$39686 ( \47035_47335 , \47033_47333 , \47034_47334 );
xor \U$39687 ( \47036_47336 , \31333_31632 , \47035_47335 );
buf \U$39688 ( \47037_47337 , \47036_47336 );
buf \U$39690 ( \47038_47338 , \47037_47337 );
xor \U$39691 ( \47039_47339 , \47032_47332 , \47038_47338 );
and \U$39692 ( \47040_47340 , \30670_29853 , \42466_42766_nG9b57 );
and \U$39693 ( \47041_47341 , \29551_29850 , \42548_42848_nG9b54 );
or \U$39694 ( \47042_47342 , \47040_47340 , \47041_47341 );
xor \U$39695 ( \47043_47343 , \29550_29849 , \47042_47342 );
buf \U$39696 ( \47044_47344 , \47043_47343 );
buf \U$39698 ( \47045_47345 , \47044_47344 );
xor \U$39699 ( \47046_47346 , \47039_47339 , \47045_47345 );
buf \U$39700 ( \47047_47347 , \47046_47346 );
xor \U$39701 ( \47048_47348 , \47027_47327 , \47047_47347 );
and \U$39702 ( \47049_47349 , \28946_28118 , \42879_43179_nG9b51 );
or \U$39704 ( \47050_47350 , \47049_47349 , 1'b0 );
xor \U$39705 ( \47051_47351 , \27815_28114 , \47050_47350 );
buf \U$39706 ( \47052_47352 , \47051_47351 );
buf \U$39707 ( \47053_47353 , \47052_47352 );
not \U$39708 ( \47054_47354 , \47053_47353 );
xor \U$39709 ( \47055_47355 , \47048_47348 , \47054_47354 );
buf \U$39710 ( \47056_47356 , \47055_47355 );
xor \U$39711 ( \47057_47357 , \47022_47322 , \47056_47356 );
and \U$39712 ( \47058_47358 , \46964_47264 , \46965_47265 );
and \U$39713 ( \47059_47359 , \46964_47264 , \46972_47272 );
and \U$39714 ( \47060_47360 , \46965_47265 , \46972_47272 );
or \U$39715 ( \47061_47361 , \47058_47358 , \47059_47359 , \47060_47360 );
buf \U$39716 ( \47062_47362 , \47061_47361 );
xor \U$39717 ( \47063_47363 , \47057_47357 , \47062_47362 );
xor \U$39718 ( \47064_47364 , \47017_47317 , \47063_47363 );
and \U$39719 ( \47065_47365 , \46959_47259 , \47001_47301 );
and \U$39720 ( \47066_47366 , \46959_47259 , \47007_47307 );
and \U$39721 ( \47067_47367 , \47001_47301 , \47007_47307 );
or \U$39722 ( \47068_47368 , \47065_47365 , \47066_47366 , \47067_47367 );
and \U$39723 ( \47069_47369 , \47064_47364 , \47068_47368 );
and \U$39725 ( \47070_47370 , \47016_47316 , \47063_47363 );
or \U$39727 ( \47071_47371 , 1'b0 , \47070_47370 , 1'b0 );
xor \U$39728 ( \47072_47372 , \47069_47369 , \47071_47371 );
and \U$39730 ( \47073_47373 , \47009_47309 , \47015_47315 );
and \U$39731 ( \47074_47374 , \47011_47311 , \47015_47315 );
or \U$39732 ( \47075_47375 , 1'b0 , \47073_47373 , \47074_47374 );
xor \U$39733 ( \47076_47376 , \47072_47372 , \47075_47375 );
xor \U$39740 ( \47077_47377 , \47076_47376 , 1'b0 );
and \U$39741 ( \47078_47378 , \47022_47322 , \47056_47356 );
and \U$39742 ( \47079_47379 , \47022_47322 , \47062_47362 );
and \U$39743 ( \47080_47380 , \47056_47356 , \47062_47362 );
or \U$39744 ( \47081_47381 , \47078_47378 , \47079_47379 , \47080_47380 );
xor \U$39745 ( \47082_47382 , \47077_47377 , \47081_47381 );
and \U$39746 ( \47083_47383 , \47027_47327 , \47047_47347 );
and \U$39747 ( \47084_47384 , \47027_47327 , \47054_47354 );
and \U$39748 ( \47085_47385 , \47047_47347 , \47054_47354 );
or \U$39749 ( \47086_47386 , \47083_47383 , \47084_47384 , \47085_47385 );
buf \U$39750 ( \47087_47387 , \47086_47386 );
and \U$39751 ( \47088_47388 , \30670_29853 , \42548_42848_nG9b54 );
and \U$39752 ( \47089_47389 , \29551_29850 , \42879_43179_nG9b51 );
or \U$39753 ( \47090_47390 , \47088_47388 , \47089_47389 );
xor \U$39754 ( \47091_47391 , \29550_29849 , \47090_47390 );
buf \U$39755 ( \47092_47392 , \47091_47391 );
buf \U$39757 ( \47093_47393 , \47092_47392 );
xor \U$39761 ( \47094_47394 , \27815_28114 , 1'b0 );
not \U$39762 ( \47095_47395 , \47094_47394 );
buf \U$39763 ( \47096_47396 , \47095_47395 );
buf \U$39765 ( \47097_47397 , \47096_47396 );
xor \U$39766 ( \47098_47398 , \47093_47393 , \47097_47397 );
and \U$39768 ( \47099_47399 , \32617_32916 , \41901_42201_nG9b5d );
or \U$39769 ( \47100_47400 , 1'b0 , \47099_47399 );
xor \U$39770 ( \47101_47401 , 1'b0 , \47100_47400 );
buf \U$39771 ( \47102_47402 , \47101_47401 );
buf \U$39773 ( \47103_47403 , \47102_47402 );
xor \U$39774 ( \47104_47404 , \47098_47398 , \47103_47403 );
buf \U$39775 ( \47105_47405 , \47104_47404 );
buf \U$39776 ( \47106_47406 , \47053_47353 );
xor \U$39777 ( \47107_47407 , \47105_47405 , \47106_47406 );
and \U$39778 ( \47108_47408 , \31989_31636 , \42133_42433_nG9b5a );
and \U$39779 ( \47109_47409 , \31334_31633 , \42466_42766_nG9b57 );
or \U$39780 ( \47110_47410 , \47108_47408 , \47109_47409 );
xor \U$39781 ( \47111_47411 , \31333_31632 , \47110_47410 );
buf \U$39782 ( \47112_47412 , \47111_47411 );
buf \U$39784 ( \47113_47413 , \47112_47412 );
xor \U$39785 ( \47114_47414 , \47107_47407 , \47113_47413 );
buf \U$39786 ( \47115_47415 , \47114_47414 );
xor \U$39787 ( \47116_47416 , \47087_47387 , \47115_47415 );
and \U$39788 ( \47117_47417 , \47032_47332 , \47038_47338 );
and \U$39789 ( \47118_47418 , \47032_47332 , \47045_47345 );
and \U$39790 ( \47119_47419 , \47038_47338 , \47045_47345 );
or \U$39791 ( \47120_47420 , \47117_47417 , \47118_47418 , \47119_47419 );
buf \U$39792 ( \47121_47421 , \47120_47420 );
xor \U$39793 ( \47122_47422 , \47116_47416 , \47121_47421 );
and \U$39794 ( \47123_47423 , \47082_47382 , \47122_47422 );
and \U$39796 ( \47124_47424 , \47076_47376 , \47081_47381 );
or \U$39798 ( \47125_47425 , 1'b0 , \47124_47424 , 1'b0 );
xor \U$39799 ( \47126_47426 , \47123_47423 , \47125_47425 );
and \U$39801 ( \47127_47427 , \47069_47369 , \47075_47375 );
and \U$39802 ( \47128_47428 , \47071_47371 , \47075_47375 );
or \U$39803 ( \47129_47429 , 1'b0 , \47127_47427 , \47128_47428 );
xor \U$39804 ( \47130_47430 , \47126_47426 , \47129_47429 );
xor \U$39811 ( \47131_47431 , \47130_47430 , 1'b0 );
and \U$39812 ( \47132_47432 , \47105_47405 , \47106_47406 );
and \U$39813 ( \47133_47433 , \47105_47405 , \47113_47413 );
and \U$39814 ( \47134_47434 , \47106_47406 , \47113_47413 );
or \U$39815 ( \47135_47435 , \47132_47432 , \47133_47433 , \47134_47434 );
buf \U$39816 ( \47136_47436 , \47135_47435 );
and \U$39817 ( \47137_47437 , \30670_29853 , \42879_43179_nG9b51 );
or \U$39819 ( \47138_47438 , \47137_47437 , 1'b0 );
xor \U$39820 ( \47139_47439 , \29550_29849 , \47138_47438 );
buf \U$39821 ( \47140_47440 , \47139_47439 );
buf \U$39822 ( \47141_47441 , \47140_47440 );
not \U$39823 ( \47142_47442 , \47141_47441 );
and \U$39825 ( \47143_47443 , \32617_32916 , \42133_42433_nG9b5a );
or \U$39826 ( \47144_47444 , 1'b0 , \47143_47443 );
xor \U$39827 ( \47145_47445 , 1'b0 , \47144_47444 );
buf \U$39828 ( \47146_47446 , \47145_47445 );
buf \U$39830 ( \47147_47447 , \47146_47446 );
xor \U$39831 ( \47148_47448 , \47142_47442 , \47147_47447 );
and \U$39832 ( \47149_47449 , \31989_31636 , \42466_42766_nG9b57 );
and \U$39833 ( \47150_47450 , \31334_31633 , \42548_42848_nG9b54 );
or \U$39834 ( \47151_47451 , \47149_47449 , \47150_47450 );
xor \U$39835 ( \47152_47452 , \31333_31632 , \47151_47451 );
buf \U$39836 ( \47153_47453 , \47152_47452 );
buf \U$39838 ( \47154_47454 , \47153_47453 );
xor \U$39839 ( \47155_47455 , \47148_47448 , \47154_47454 );
buf \U$39840 ( \47156_47456 , \47155_47455 );
xor \U$39841 ( \47157_47457 , \47136_47436 , \47156_47456 );
and \U$39842 ( \47158_47458 , \47093_47393 , \47097_47397 );
and \U$39843 ( \47159_47459 , \47093_47393 , \47103_47403 );
and \U$39844 ( \47160_47460 , \47097_47397 , \47103_47403 );
or \U$39845 ( \47161_47461 , \47158_47458 , \47159_47459 , \47160_47460 );
buf \U$39846 ( \47162_47462 , \47161_47461 );
xor \U$39847 ( \47163_47463 , \47157_47457 , \47162_47462 );
xor \U$39848 ( \47164_47464 , \47131_47431 , \47163_47463 );
and \U$39849 ( \47165_47465 , \47087_47387 , \47115_47415 );
and \U$39850 ( \47166_47466 , \47087_47387 , \47121_47421 );
and \U$39851 ( \47167_47467 , \47115_47415 , \47121_47421 );
or \U$39852 ( \47168_47468 , \47165_47465 , \47166_47466 , \47167_47467 );
and \U$39853 ( \47169_47469 , \47164_47464 , \47168_47468 );
and \U$39855 ( \47170_47470 , \47130_47430 , \47163_47463 );
or \U$39857 ( \47171_47471 , 1'b0 , \47170_47470 , 1'b0 );
xor \U$39858 ( \47172_47472 , \47169_47469 , \47171_47471 );
and \U$39860 ( \47173_47473 , \47123_47423 , \47129_47429 );
and \U$39861 ( \47174_47474 , \47125_47425 , \47129_47429 );
or \U$39862 ( \47175_47475 , 1'b0 , \47173_47473 , \47174_47474 );
xor \U$39863 ( \47176_47476 , \47172_47472 , \47175_47475 );
xor \U$39865 ( \47177_47477 , \47176_47476 , 1'b1 );
buf \U$39867 ( \47178_47478 , \47141_47441 );
xor \U$39868 ( \47179_47479 , 1'b1 , \47178_47478 );
and \U$39870 ( \47180_47480 , \32617_32916 , \42466_42766_nG9b57 );
or \U$39871 ( \47181_47481 , 1'b0 , \47180_47480 );
xor \U$39872 ( \47182_47482 , 1'b0 , \47181_47481 );
buf \U$39873 ( \47183_47483 , \47182_47482 );
buf \U$39874 ( \47184_47484 , \47183_47483 );
not \U$39875 ( \47185_47485 , \47184_47484 );
xor \U$39876 ( \47186_47486 , \47179_47479 , \47185_47485 );
buf \U$39877 ( \47187_47487 , \47186_47486 );
xor \U$39881 ( \47188_47488 , \29550_29849 , 1'b0 );
not \U$39882 ( \47189_47489 , \47188_47488 );
buf \U$39883 ( \47190_47490 , \47189_47489 );
buf \U$39885 ( \47191_47491 , \47190_47490 );
buf \U$39886 ( \47192_47492 , \47184_47484 );
xor \U$39887 ( \47193_47493 , \47191_47491 , \47192_47492 );
buf \U$39888 ( \47194_47494 , \47193_47493 );
xor \U$39889 ( \47195_47495 , \47187_47487 , \47194_47494 );
xor \U$39890 ( \47196_47496 , \47177_47477 , \47195_47495 );
xor \U$39897 ( \47197_47497 , \47196_47496 , 1'b0 );
and \U$39898 ( \47198_47498 , \47142_47442 , \47147_47447 );
and \U$39899 ( \47199_47499 , \47142_47442 , \47154_47454 );
and \U$39900 ( \47200_47500 , \47147_47447 , \47154_47454 );
or \U$39901 ( \47201_47501 , \47198_47498 , \47199_47499 , \47200_47500 );
buf \U$39902 ( \47202_47502 , \47201_47501 );
and \U$39903 ( \47203_47503 , \31989_31636 , \42548_42848_nG9b54 );
and \U$39904 ( \47204_47504 , \31334_31633 , \42879_43179_nG9b51 );
or \U$39905 ( \47205_47505 , \47203_47503 , \47204_47504 );
xor \U$39906 ( \47206_47506 , \31333_31632 , \47205_47505 );
buf \U$39907 ( \47207_47507 , \47206_47506 );
buf \U$39909 ( \47208_47508 , \47207_47507 );
not \U$39910 ( \47209_47509 , \47141_47441 );
xor \U$39911 ( \47210_47510 , \47208_47508 , \47209_47509 );
buf \U$39912 ( \47211_47511 , \47184_47484 );
xor \U$39913 ( \47212_47512 , \47210_47510 , \47211_47511 );
buf \U$39914 ( \47213_47513 , \47212_47512 );
xor \U$39915 ( \47214_47514 , \47202_47502 , \47213_47513 );
buf \U$39916 ( \47215_47515 , \47141_47441 );
xor \U$39917 ( \47216_47516 , \47214_47514 , \47215_47515 );
xor \U$39918 ( \47217_47517 , \47197_47497 , \47216_47516 );
and \U$39919 ( \47218_47518 , \47136_47436 , \47156_47456 );
and \U$39920 ( \47219_47519 , \47136_47436 , \47162_47462 );
and \U$39921 ( \47220_47520 , \47156_47456 , \47162_47462 );
or \U$39922 ( \47221_47521 , \47218_47518 , \47219_47519 , \47220_47520 );
and \U$39923 ( \47222_47522 , \47217_47517 , \47221_47521 );
and \U$39925 ( \47223_47523 , \47196_47496 , \47216_47516 );
or \U$39927 ( \47224_47524 , 1'b0 , \47223_47523 , 1'b0 );
xor \U$39928 ( \47225_47525 , \47222_47522 , \47224_47524 );
and \U$39929 ( \47226_47526 , \47176_47476 , 1'b1 );
and \U$39930 ( \47227_47527 , \47176_47476 , \47195_47495 );
and \U$39931 ( \47228_47528 , 1'b1 , \47195_47495 );
or \U$39932 ( \47229_47529 , \47226_47526 , \47227_47527 , \47228_47528 );
xor \U$39933 ( \47230_47530 , \47225_47525 , \47229_47529 );
and \U$39935 ( \47231_47531 , \47169_47469 , \47175_47475 );
and \U$39936 ( \47232_47532 , \47171_47471 , \47175_47475 );
or \U$39937 ( \47233_47533 , 1'b0 , \47231_47531 , \47232_47532 );
xor \U$39938 ( \47234_47534 , \47230_47530 , \47233_47533 );
and \U$39939 ( \47235_47535 , \47187_47487 , \47194_47494 );
xor \U$39940 ( \47236_47536 , \47234_47534 , \47235_47535 );
xor \U$39947 ( \47237_47537 , \47236_47536 , 1'b0 );
and \U$39949 ( \47238_47538 , \32617_32916 , \42548_42848_nG9b54 );
or \U$39950 ( \47239_47539 , 1'b0 , \47238_47538 );
xor \U$39951 ( \47240_47540 , 1'b0 , \47239_47539 );
buf \U$39952 ( \47241_47541 , \47240_47540 );
buf \U$39953 ( \47242_47542 , \47241_47541 );
xor \U$39954 ( \47243_47543 , \47237_47537 , \47242_47542 );
and \U$39955 ( \47244_47544 , \47208_47508 , \47209_47509 );
and \U$39956 ( \47245_47545 , \47208_47508 , \47211_47511 );
and \U$39957 ( \47246_47546 , \47209_47509 , \47211_47511 );
or \U$39958 ( \47247_47547 , \47244_47544 , \47245_47545 , \47246_47546 );
buf \U$39959 ( \47248_47548 , \47247_47547 );
and \U$39960 ( \47249_47549 , 1'b1 , \47178_47478 );
and \U$39961 ( \47250_47550 , 1'b1 , \47185_47485 );
and \U$39962 ( \47251_47551 , \47178_47478 , \47185_47485 );
or \U$39963 ( \47252_47552 , \47249_47549 , \47250_47550 , \47251_47551 );
buf \U$39964 ( \47253_47553 , \47252_47552 );
xor \U$39965 ( \47254_47554 , \47248_47548 , \47253_47553 );
and \U$39967 ( \47255_47555 , \47191_47491 , \47192_47492 );
buf \U$39968 ( \47256_47556 , \47255_47555 );
xor \U$39969 ( \47257_47557 , 1'b1 , \47256_47556 );
and \U$39970 ( \47258_47558 , \31989_31636 , \42879_43179_nG9b51 );
or \U$39972 ( \47259_47559 , \47258_47558 , 1'b0 );
xor \U$39973 ( \47260_47560 , \31333_31632 , \47259_47559 );
buf \U$39974 ( \47261_47561 , \47260_47560 );
buf \U$39976 ( \47262_47562 , \47261_47561 );
xor \U$39977 ( \47263_47563 , \47257_47557 , \47262_47562 );
xor \U$39978 ( \47264_47564 , \47254_47554 , \47263_47563 );
and \U$39979 ( \47265_47565 , \47243_47543 , \47264_47564 );
and \U$39980 ( \47266_47566 , \47202_47502 , \47213_47513 );
and \U$39981 ( \47267_47567 , \47202_47502 , \47215_47515 );
and \U$39982 ( \47268_47568 , \47213_47513 , \47215_47515 );
or \U$39983 ( \47269_47569 , \47266_47566 , \47267_47567 , \47268_47568 );
and \U$39984 ( \47270_47570 , \47243_47543 , \47269_47569 );
and \U$39985 ( \47271_47571 , \47264_47564 , \47269_47569 );
or \U$39986 ( \47272_47572 , \47265_47565 , \47270_47570 , \47271_47571 );
and \U$39988 ( \47273_47573 , \47236_47536 , \47242_47542 );
or \U$39990 ( \47274_47574 , 1'b0 , \47273_47573 , 1'b0 );
xor \U$39991 ( \47275_47575 , \47272_47572 , \47274_47574 );
and \U$39992 ( \47276_47576 , \47230_47530 , \47233_47533 );
and \U$39993 ( \47277_47577 , \47230_47530 , \47235_47535 );
and \U$39994 ( \47278_47578 , \47233_47533 , \47235_47535 );
or \U$39995 ( \47279_47579 , \47276_47576 , \47277_47577 , \47278_47578 );
xor \U$39996 ( \47280_47580 , \47275_47575 , \47279_47579 );
and \U$39998 ( \47281_47581 , \47222_47522 , \47229_47529 );
and \U$39999 ( \47282_47582 , \47224_47524 , \47229_47529 );
or \U$40000 ( \47283_47583 , 1'b0 , \47281_47581 , \47282_47582 );
xor \U$40001 ( \47284_47584 , \47280_47580 , \47283_47583 );
xor \U$40003 ( \47285_47585 , \47284_47584 , 1'b1 );
xor \U$40010 ( \47286_47586 , \47285_47585 , 1'b0 );
and \U$40012 ( \47287_47587 , \32617_32916 , \42879_43179_nG9b51 );
or \U$40013 ( \47288_47588 , 1'b0 , \47287_47587 );
xor \U$40014 ( \47289_47589 , 1'b0 , \47288_47588 );
buf \U$40015 ( \47290_47590 , \47289_47589 );
buf \U$40016 ( \47291_47591 , \47290_47590 );
xor \U$40017 ( \47292_47592 , \47286_47586 , \47291_47591 );
and \U$40018 ( \47293_47593 , \47248_47548 , \47253_47553 );
and \U$40019 ( \47294_47594 , \47248_47548 , \47263_47563 );
and \U$40020 ( \47295_47595 , \47253_47553 , \47263_47563 );
or \U$40021 ( \47296_47596 , \47293_47593 , \47294_47594 , \47295_47595 );
xor \U$40022 ( \47297_47597 , \47292_47592 , \47296_47596 );
and \U$40023 ( \47298_47598 , 1'b1 , \47256_47556 );
and \U$40024 ( \47299_47599 , 1'b1 , \47262_47562 );
and \U$40025 ( \47300_47600 , \47256_47556 , \47262_47562 );
or \U$40026 ( \47301_47601 , \47298_47598 , \47299_47599 , \47300_47600 );
xor \U$40027 ( \47302_47602 , \47297_47597 , \47301_47601 );
xor \U$40031 ( \47303_47603 , \31333_31632 , 1'b0 );
not \U$40032 ( \47304_47604 , \47303_47603 );
buf \U$40033 ( \47305_47605 , \47304_47604 );
buf \U$40034 ( \47306_47606 , \47305_47605 );
xor \U$40035 ( \47307_47607 , \47302_47602 , \47306_47606 );
buf gdf4e_GF_PartitionCandidate( \47308_47608_nGdf4e , \47307_47607 );
buf \U$labaj5628 ( \47309_R_58_102f1b78 , \47308_47608_nGdf4e );
xor \U$40037 ( \47310_47610 , \47243_47543 , \47264_47564 );
xor \U$40038 ( \47311_47611 , \47310_47610 , \47269_47569 );
buf gdf51_GF_PartitionCandidate( \47312_47612_nGdf51 , \47311_47611 );
buf \U$labaj5629 ( \47313_R_59_be1fc68 , \47312_47612_nGdf51 );
xor \U$40040 ( \47314_47614 , \47217_47517 , \47221_47521 );
buf gdf53_GF_PartitionCandidate( \47315_47615_nGdf53 , \47314_47614 );
buf \U$labaj5630 ( \47316_R_5a_10279198 , \47315_47615_nGdf53 );
xor \U$40042 ( \47317_47617 , \47164_47464 , \47168_47468 );
buf gdf55_GF_PartitionCandidate( \47318_47618_nGdf55 , \47317_47617 );
buf \U$labaj5631 ( \47319_R_5b_102299e8 , \47318_47618_nGdf55 );
xor \U$40044 ( \47320_47620 , \47082_47382 , \47122_47422 );
buf gdf57_GF_PartitionCandidate( \47321_47621_nGdf57 , \47320_47620 );
buf \U$labaj5632 ( \47322_R_5c_101d0448 , \47321_47621_nGdf57 );
xor \U$40046 ( \47323_47623 , \47064_47364 , \47068_47368 );
buf gdf59_GF_PartitionCandidate( \47324_47624_nGdf59 , \47323_47623 );
buf \U$labaj5633 ( \47325_R_5d_f7f82f0 , \47324_47624_nGdf59 );
xor \U$40048 ( \47326_47626 , \46954_47254 , \47008_47308 );
buf gdf5b_GF_PartitionCandidate( \47327_47627_nGdf5b , \47326_47626 );
buf \U$labaj5634 ( \47328_R_5e_be21600 , \47327_47627_nGdf5b );
xor \U$40050 ( \47329_47629 , \46936_47236 , \46940_47240 );
buf gdf5d_GF_PartitionCandidate( \47330_47630_nGdf5d , \47329_47629 );
buf \U$labaj5635 ( \47331_R_5f_f7fa5b8 , \47330_47630_nGdf5d );
xor \U$40052 ( \47332_47632 , \46862_47162 , \46866_47166 );
buf gdf5f_GF_PartitionCandidate( \47333_47633_nGdf5f , \47332_47632 );
buf \U$labaj5636 ( \47334_R_60_1027d530 , \47333_47633_nGdf5f );
xor \U$40054 ( \47335_47635 , \46710_47010 , \46784_47084 );
buf gdf61_GF_PartitionCandidate( \47336_47636_nGdf61 , \47335_47635 );
buf \U$labaj5637 ( \47337_R_61_10205ae8 , \47336_47636_nGdf61 );
xor \U$40056 ( \47338_47638 , \46614_46914 , \46696_46996 );
buf gdf63_GF_PartitionCandidate( \47339_47639_nGdf63 , \47338_47638 );
buf \U$labaj5638 ( \47340_R_62_10283510 , \47339_47639_nGdf63 );
xor \U$40058 ( \47341_47641 , \46512_46812 , \46600_46900 );
buf gdf65_GF_PartitionCandidate( \47342_47642_nGdf65 , \47341_47641 );
buf \U$labaj5639 ( \47343_R_63_f82b578 , \47342_47642_nGdf65 );
xor \U$40060 ( \47344_47644 , \46402_46702 , \46498_46798 );
buf gdf67_GF_PartitionCandidate( \47345_47645_nGdf67 , \47344_47644 );
buf \U$labaj5640 ( \47346_R_64_ace4e68 , \47345_47645_nGdf67 );
xor \U$40062 ( \47347_47647 , \46286_46586 , \46388_46688 );
buf gdf69_GF_PartitionCandidate( \47348_47648_nGdf69 , \47347_47647 );
buf \U$labaj5641 ( \47349_R_65_f8204e0 , \47348_47648_nGdf69 );
xor \U$40064 ( \47350_47650 , \46162_46462 , \46272_46572 );
buf gdf6b_GF_PartitionCandidate( \47351_47651_nGdf6b , \47350_47650 );
buf \U$labaj5642 ( \47352_R_66_1027a0b0 , \47351_47651_nGdf6b );
xor \U$40066 ( \47353_47653 , \46032_46332 , \46148_46448 );
buf gdf6d_GF_PartitionCandidate( \47354_47654_nGdf6d , \47353_47653 );
buf \U$labaj5643 ( \47355_R_67_1022dc30 , \47354_47654_nGdf6d );
xor \U$40068 ( \47356_47656 , \46014_46314 , \46018_46318 );
buf gdf6f_GF_PartitionCandidate( \47357_47657_nGdf6f , \47356_47656 );
buf \U$labaj5644 ( \47358_R_68_102478a8 , \47357_47657_nGdf6f );
xor \U$40070 ( \47359_47659 , \45876_46176 , \45880_46180 );
buf gdf71_GF_PartitionCandidate( \47360_47660_nGdf71 , \47359_47659 );
buf \U$labaj5645 ( \47361_R_69_10286f78 , \47360_47660_nGdf71 );
xor \U$40072 ( \47362_47662 , \45598_45898 , \45736_46036 );
buf gdf73_GF_PartitionCandidate( \47363_47663_nGdf73 , \47362_47662 );
buf \U$labaj5646 ( \47364_R_6a_f7edd80 , \47363_47663_nGdf73 );
xor \U$40074 ( \47365_47665 , \45440_45740 , \45584_45884 );
buf gdf75_GF_PartitionCandidate( \47366_47666_nGdf75 , \47365_47665 );
buf \U$labaj5647 ( \47367_R_6b_101c3628 , \47366_47666_nGdf75 );
xor \U$40076 ( \47368_47668 , \45274_45574 , \45426_45726 );
buf gdf77_GF_PartitionCandidate( \47369_47669_nGdf77 , \47368_47668 );
buf \U$labaj5648 ( \47370_R_6c_f7fbe00 , \47369_47669_nGdf77 );
xor \U$40078 ( \47371_47671 , \45102_45402 , \45260_45560 );
buf gdf79_GF_PartitionCandidate( \47372_47672_nGdf79 , \47371_47671 );
buf \U$labaj5649 ( \47373_R_6d_f7ce9f8 , \47372_47672_nGdf79 );
xor \U$40080 ( \47374_47674 , \44922_45222 , \45088_45388 );
buf gdf7b_GF_PartitionCandidate( \47375_47675_nGdf7b , \47374_47674 );
buf \U$labaj5650 ( \47376_R_6e_f7c8830 , \47375_47675_nGdf7b );
xor \U$40082 ( \47377_47677 , \44736_45036 , \44908_45208 );
buf gdf7d_GF_PartitionCandidate( \47378_47678_nGdf7d , \47377_47677 );
buf \U$labaj5651 ( \47379_R_6f_101ffc68 , \47378_47678_nGdf7d );
xor \U$40084 ( \47380_47680 , \44718_45018 , \44722_45022 );
buf gdf7f_GF_PartitionCandidate( \47381_47681_nGdf7f , \47380_47680 );
buf \U$labaj5652 ( \47382_R_70_f7d4000 , \47381_47681_nGdf7f );
xor \U$40086 ( \47383_47683 , \44342_44642 , \44528_44828 );
buf gdf81_GF_PartitionCandidate( \47384_47684_nGdf81 , \47383_47683 );
buf \U$labaj5653 ( \47385_R_71_acee958 , \47384_47684_nGdf81 );
xor \U$40088 ( \47386_47686 , \44134_44434 , \44328_44628 );
buf gdf83_GF_PartitionCandidate( \47387_47687_nGdf83 , \47386_47686 );
buf \U$labaj5654 ( \47388_R_72_94046c0 , \47387_47687_nGdf83 );
xor \U$40090 ( \47389_47689 , \43920_44220 , \44120_44420 );
buf gdf85_GF_PartitionCandidate( \47390_47690_nGdf85 , \47389_47689 );
buf \U$labaj5655 ( \47391_R_73_101ee420 , \47390_47690_nGdf85 );
xor \U$40092 ( \47392_47692 , \43698_43998 , \43906_44206 );
buf gdf87_GF_PartitionCandidate( \47393_47693_nGdf87 , \47392_47692 );
buf \U$labaj5656 ( \47394_R_74_102eb268 , \47393_47693_nGdf87 );
xor \U$40094 ( \47395_47695 , \43470_43770 , \43684_43984 );
buf gdf89_GF_PartitionCandidate( \47396_47696_nGdf89 , \47395_47695 );
buf \U$labaj5657 ( \47397_R_75_b320c50 , \47396_47696_nGdf89 );
xor \U$40096 ( \47398_47698 , \43238_43538 , \43456_43756 );
buf gdf8b_GF_PartitionCandidate( \47399_47699_nGdf8b , \47398_47698 );
buf \U$labaj5658 ( \47400_R_76_ad80a90 , \47399_47699_nGdf8b );
xor \U$40098 ( \47401_47701 , \43006_43306 , \43224_43524 );
buf gdf8d_GF_PartitionCandidate( \47402_47702_nGdf8d , \47401_47701 );
buf \U$labaj5659 ( \47403_R_77_1027fd48 , \47402_47702_nGdf8d );
xor \U$40100 ( \47404_47704 , \42758_43058 , \42992_43292 );
buf gdf8f_GF_PartitionCandidate( \47405_47705_nGdf8f , \47404_47704 );
buf \U$labaj5660 ( \47406_R_78_f7ce4b8 , \47405_47705_nGdf8f );
xor \U$40102 ( \47407_47707 , \42504_42804 , \42744_43044 );
buf gdf91_GF_PartitionCandidate( \47408_47708_nGdf91 , \47407_47707 );
buf \U$labaj5661 ( \47409_R_79_ad77048 , \47408_47708_nGdf91 );
xor \U$40104 ( \47410_47710 , \42246_42546 , \42490_42790 );
buf gdf93_GF_PartitionCandidate( \47411_47711_nGdf93 , \47410_47710 );
buf \U$labaj5662 ( \47412_R_7a_102a6ae0 , \47411_47711_nGdf93 );
xor \U$40106 ( \47413_47713 , \41982_42282 , \42232_42532 );
buf gdf95_GF_PartitionCandidate( \47414_47714_nGdf95 , \47413_47713 );
buf \U$labaj5663 ( \47415_R_7b_f7e4c78 , \47414_47714_nGdf95 );
xor \U$40108 ( \47416_47716 , \41714_42014 , \41968_42268 );
buf gdf97_GF_PartitionCandidate( \47417_47717_nGdf97 , \47416_47716 );
buf \U$labaj5664 ( \47418_R_7c_e2a6ce0 , \47417_47717_nGdf97 );
xor \U$40110 ( \47419_47719 , \41440_41740 , \41700_42000 );
buf gdf99_GF_PartitionCandidate( \47420_47720_nGdf99 , \47419_47719 );
buf \U$labaj5665 ( \47421_R_7d_101e86e0 , \47420_47720_nGdf99 );
xor \U$40112 ( \47422_47722 , \41162_41462 , \41426_41726 );
buf gdf9b_GF_PartitionCandidate( \47423_47723_nGdf9b , \47422_47722 );
buf \U$labaj5666 ( \47424_R_7e_e2a9cc8 , \47423_47723_nGdf9b );
xor \U$40114 ( \47425_47725 , \40878_41178 , \41148_41448 );
buf gdf9d_GF_PartitionCandidate( \47426_47726_nGdf9d , \47425_47725 );
buf \U$labaj5667 ( \47427_R_7f_10292be0 , \47426_47726_nGdf9d );
xor \U$40116 ( \47428_47728 , \40590_40890 , \40864_41164 );
buf gdf9f_GF_PartitionCandidate( \47429_47729_nGdf9f , \47428_47728 );
buf \U$labaj5668 ( \47430_R_80_b33cde8 , \47429_47729_nGdf9f );
xor \U$40118 ( \47431_47731 , \40296_40596 , \40576_40876 );
buf gdfa1_GF_PartitionCandidate( \47432_47732_nGdfa1 , \47431_47731 );
buf \U$labaj5669 ( \47433_R_81_101e2908 , \47432_47732_nGdfa1 );
xor \U$40120 ( \47434_47734 , \39998_40298 , \40282_40582 );
buf gdfa3_GF_PartitionCandidate( \47435_47735_nGdfa3 , \47434_47734 );
buf \U$labaj5670 ( \47436_R_82_102e9780 , \47435_47735_nGdfa3 );
xor \U$40122 ( \47437_47737 , \39694_39994 , \39984_40284 );
buf gdfa5_GF_PartitionCandidate( \47438_47738_nGdfa5 , \47437_47737 );
buf \U$labaj5671 ( \47439_R_83_f8157a0 , \47438_47738_nGdfa5 );
xor \U$40124 ( \47440_47740 , \39676_39976 , \39680_39980 );
buf gdfa7_GF_PartitionCandidate( \47441_47741_nGdfa7 , \47440_47740 );
buf \U$labaj5672 ( \47442_R_84_f819358 , \47441_47741_nGdfa7 );
xor \U$40126 ( \47443_47743 , \39072_39372 , \39372_39672 );
buf gdfa9_GF_PartitionCandidate( \47444_47744_nGdfa9 , \47443_47743 );
buf \U$labaj5673 ( \47445_R_85_ace8b70 , \47444_47744_nGdfa9 );
xor \U$40128 ( \47446_47746 , \38754_39054 , \39058_39358 );
buf gdfab_GF_PartitionCandidate( \47447_47747_nGdfab , \47446_47746 );
buf \U$labaj5674 ( \47448_R_86_be142b0 , \47447_47747_nGdfab );
xor \U$40130 ( \47449_47749 , \38430_38730 , \38740_39040 );
buf gdfad_GF_PartitionCandidate( \47450_47750_nGdfad , \47449_47749 );
buf \U$labaj5675 ( \47451_R_87_f81b770 , \47450_47750_nGdfad );
xor \U$40132 ( \47452_47752 , \38412_38712 , \38416_38716 );
buf gdfaf_GF_PartitionCandidate( \47453_47753_nGdfaf , \47452_47752 );
buf \U$labaj5676 ( \47454_R_88_b330278 , \47453_47753_nGdfaf );
xor \U$40134 ( \47455_47755 , \37768_38068 , \38088_38388 );
buf gdfb1_GF_PartitionCandidate( \47456_47756_nGdfb1 , \47455_47755 );
buf \U$labaj5677 ( \47457_R_89_f7fe9f8 , \47456_47756_nGdfb1 );
xor \U$40136 ( \47458_47758 , \37430_37730 , \37754_38054 );
buf gdfb3_GF_PartitionCandidate( \47459_47759_nGdfb3 , \47458_47758 );
buf \U$labaj5678 ( \47460_R_8a_101cf488 , \47459_47759_nGdfb3 );
xor \U$40138 ( \47461_47761 , \37086_37386 , \37416_37716 );
buf gdfb5_GF_PartitionCandidate( \47462_47762_nGdfb5 , \47461_47761 );
buf \U$labaj5679 ( \47463_R_8b_f8225c0 , \47462_47762_nGdfb5 );
xor \U$40140 ( \47464_47764 , \36738_37038 , \37072_37372 );
buf gdfb7_GF_PartitionCandidate( \47465_47765_nGdfb7 , \47464_47764 );
buf \U$labaj5680 ( \47466_R_8c_101d4738 , \47465_47765_nGdfb7 );
xor \U$40142 ( \47467_47767 , \36384_36684 , \36724_37024 );
buf gdfb9_GF_PartitionCandidate( \47468_47768_nGdfb9 , \47467_47767 );
buf \U$labaj5681 ( \47469_R_8d_101c4000 , \47468_47768_nGdfb9 );
xor \U$40144 ( \47470_47770 , \36026_36326 , \36370_36670 );
buf gdfbb_GF_PartitionCandidate( \47471_47771_nGdfbb , \47470_47770 );
buf \U$labaj5682 ( \47472_R_8e_101fe960 , \47471_47771_nGdfbb );
xor \U$40146 ( \47473_47773 , \35662_35962 , \36012_36312 );
buf gdfbd_GF_PartitionCandidate( \47474_47774_nGdfbd , \47473_47773 );
buf \U$labaj5683 ( \47475_R_8f_102a0330 , \47474_47774_nGdfbd );
xor \U$40148 ( \47476_47776 , \35294_35594 , \35648_35948 );
buf gdfbf_GF_PartitionCandidate( \47477_47777_nGdfbf , \47476_47776 );
buf \U$labaj5684 ( \47478_R_90_f7f4bd0 , \47477_47777_nGdfbf );
xor \U$40150 ( \47479_47779 , \34920_35220 , \35280_35580 );
buf gdfc1_GF_PartitionCandidate( \47480_47780_nGdfc1 , \47479_47779 );
buf \U$labaj5685 ( \47481_R_91_1023e5a8 , \47480_47780_nGdfc1 );
xor \U$40152 ( \47482_47782 , \34542_34842 , \34906_35206 );
buf gdfc3_GF_PartitionCandidate( \47483_47783_nGdfc3 , \47482_47782 );
buf \U$labaj5686 ( \47484_R_92_10248da8 , \47483_47783_nGdfc3 );
xor \U$40154 ( \47485_47785 , \34159_34459 , \34529_34829 );
buf gdfc5_GF_PartitionCandidate( \47486_47786_nGdfc5 , \47485_47785 );
buf \U$labaj5687 ( \47487_R_93_be2c938 , \47486_47786_nGdfc5 );
xor \U$40156 ( \47488_47788 , \33775_34075 , \34146_34446 );
buf gdfc7_GF_PartitionCandidate( \47489_47789_nGdfc7 , \47488_47788 );
buf \U$labaj5688 ( \47490_R_94_f7f5458 , \47489_47789_nGdfc7 );
xor \U$40158 ( \47491_47791 , \33382_33682 , \33386_33686 );
xor \U$40159 ( \47492_47792 , \47491_47791 , \33762_34062 );
buf gdfca_GF_PartitionCandidate( \47493_47793_nGdfca , \47492_47792 );
buf \U$labaj5689 ( \47494_R_95_f7c6808 , \47493_47793_nGdfca );
xor \U$40161 ( \47495_47795 , \33001_33301 , \33370_33670 );
xor \U$40162 ( \47496_47796 , \47495_47795 , \33375_33675 );
buf gdfcd_GF_PartitionCandidate( \47497_47797_nGdfcd , \47496_47796 );
buf \U$labaj5690 ( \47498_R_96_be316a8 , \47497_47797_nGdfcd );
xor \U$40164 ( \47499_47799 , \32624_32924 , \32628_32928 );
xor \U$40165 ( \47500_47800 , \47499_47799 , \32992_33292 );
buf gdfd0_GF_PartitionCandidate( \47501_47801_nGdfd0 , \47500_47800 );
buf \U$labaj5691 ( \47502_R_97_e2a0328 , \47501_47801_nGdfd0 );
xor \U$40167 ( \47503_47803 , \32606_32905 , \32610_32909 );
buf gdfd2_GF_PartitionCandidate( \47504_47804_nGdfd2 , \47503_47803 );
buf \U$labaj5692 ( \47505_R_98_be2d850 , \47504_47804_nGdfd2 );
xor \U$40169 ( \47506_47806 , \31341_31643 , \31345_31647 );
xor \U$40170 ( \47507_47807 , \47506_47806 , \31957_32259 );
buf gdfd5_GF_PartitionCandidate( \47508_47808_nGdfd5 , \47507_47807 );
buf \U$labaj5693 ( \47509_R_99_10217db0 , \47508_47808_nGdfd5 );
xor \U$40172 ( \47510_47810 , \30163_30465 , \30779_31078 );
buf gdfd7_GF_PartitionCandidate( \47511_47811_nGdfd7 , \47510_47810 );
buf \U$labaj5694 ( \47512_R_9a_f7ec340 , \47511_47811_nGdfd7 );
xor \U$40174 ( \47513_47813 , \29558_29860 , \29562_29864 );
xor \U$40175 ( \47514_47814 , \47513_47813 , \30150_30452 );
buf gdfda_GF_PartitionCandidate( \47515_47815_nGdfda , \47514_47814 );
buf \U$labaj5695 ( \47516_R_9b_be23ec0 , \47515_47815_nGdfda );
xor \U$40177 ( \47517_47817 , \28404_28706 , \28996_29295 );
buf gdfdc_GF_PartitionCandidate( \47518_47818_nGdfdc , \47517_47817 );
buf \U$labaj5696 ( \47519_R_9c_101d4540 , \47518_47818_nGdfdc );
xor \U$40179 ( \47520_47820 , \27823_28125 , \27827_28129 );
xor \U$40180 ( \47521_47821 , \47520_47820 , \28391_28693 );
buf gdfdf_GF_PartitionCandidate( \47522_47822_nGdfdf , \47521_47821 );
buf \U$labaj5697 ( \47523_R_9d_f800828 , \47522_47822_nGdfdf );
xor \U$40182 ( \47524_47824 , \26693_26995 , \27261_27560 );
buf gdfe1_GF_PartitionCandidate( \47525_47825_nGdfe1 , \47524_47824 );
buf \U$labaj5698 ( \47526_R_9e_102970c8 , \47525_47825_nGdfe1 );
xor \U$40184 ( \47527_47827 , \26136_26438 , \26140_26442 );
xor \U$40185 ( \47528_47828 , \47527_47827 , \26680_26982 );
buf gdfe4_GF_PartitionCandidate( \47529_47829_nGdfe4 , \47528_47828 );
buf \U$labaj5699 ( \47530_R_9f_10221de0 , \47529_47829_nGdfe4 );
xor \U$40187 ( \47531_47831 , \25570_25869 , \25574_25873 );
buf gdfe6_GF_PartitionCandidate( \47532_47832_nGdfe6 , \47531_47831 );
buf \U$labaj5700 ( \47533_R_a0_ad8d568 , \47532_47832_nGdfe6 );
xor \U$40189 ( \47534_47834 , \24497_24799 , \25012_25314 );
xor \U$40190 ( \47535_47835 , \47534_47834 , \25017_25319 );
buf gdfe9_GF_PartitionCandidate( \47536_47836_nGdfe9 , \47535_47835 );
buf \U$labaj5701 ( \47537_R_a1_be4eb58 , \47536_47836_nGdfe9 );
xor \U$40192 ( \47538_47838 , \23415_23717 , \23935_24234 );
buf gdfeb_GF_PartitionCandidate( \47539_47839_nGdfeb , \47538_47838 );
buf \U$labaj5702 ( \47540_R_a2_f7c5500 , \47539_47839_nGdfeb );
xor \U$40194 ( \47541_47841 , \22906_23208 , \22910_23212 );
xor \U$40195 ( \47542_47842 , \47541_47841 , \23402_23704 );
buf gdfee_GF_PartitionCandidate( \47543_47843_nGdfee , \47542_47842 );
buf \U$labaj5703 ( \47544_R_a3_ad88f30 , \47543_47843_nGdfee );
xor \U$40197 ( \47545_47845 , \21848_22150 , \22344_22643 );
buf gdff0_GF_PartitionCandidate( \47546_47846_nGdff0 , \47545_47845 );
buf \U$labaj5704 ( \47547_R_a4_f82f088 , \47546_47846_nGdff0 );
xor \U$40199 ( \47548_47848 , \21363_21665 , \21367_21669 );
xor \U$40200 ( \47549_47849 , \47548_47848 , \21835_22137 );
buf gdff3_GF_PartitionCandidate( \47550_47850_nGdff3 , \47549_47849 );
buf \U$labaj5705 ( \47551_R_a5_f7dcbc8 , \47550_47850_nGdff3 );
xor \U$40202 ( \47552_47852 , \20329_20631 , \20801_21100 );
buf gdff5_GF_PartitionCandidate( \47553_47853_nGdff5 , \47552_47852 );
buf \U$labaj5706 ( \47554_R_a6_10292940 , \47553_47853_nGdff5 );
xor \U$40204 ( \47555_47855 , \19304_19603 , \19859_20161 );
xor \U$40205 ( \47556_47856 , \47555_47855 , \20316_20618 );
buf gdff8_GF_PartitionCandidate( \47557_47857_nGdff8 , \47556_47856 );
buf \U$labaj5707 ( \47558_R_a7_be138d8 , \47557_47857_nGdff8 );
xor \U$40207 ( \47559_47859 , \18842_19144 , \19303_19602 );
buf gdffa_GF_PartitionCandidate( \47560_47860_nGdffa , \47559_47859 );
buf \U$labaj5708 ( \47561_R_a8_acee418 , \47560_47860_nGdffa );
xor \U$40209 ( \47562_47862 , \17851_18150 , \18406_18708 );
xor \U$40210 ( \47563_47863 , \47562_47862 , \18839_19141 );
buf gdffd_GF_PartitionCandidate( \47564_47864_nGdffd , \47563_47863 );
buf \U$labaj5709 ( \47565_R_a9_ad84450 , \47564_47864_nGdffd );
xor \U$40212 ( \47566_47866 , \17413_17715 , \17850_18149 );
buf gdfff_GF_PartitionCandidate( \47567_47867_nGdfff , \47566_47866 );
buf \U$labaj5710 ( \47568_R_aa_be10838 , \47567_47867_nGdfff );
xor \U$40214 ( \47569_47869 , \16446_16745 , \17001_17303 );
xor \U$40215 ( \47570_47870 , \47569_47869 , \17410_17712 );
buf ge002_GF_PartitionCandidate( \47571_47871_nGe002 , \47570_47870 );
buf \U$labaj5711 ( \47572_R_ab_be31fd8 , \47571_47871_nGe002 );
xor \U$40217 ( \47573_47873 , \16032_16334 , \16445_16744 );
buf ge004_GF_PartitionCandidate( \47574_47874_nGe004 , \47573_47873 );
buf \U$labaj5712 ( \47575_R_ac_acdaef0 , \47574_47874_nGe004 );
xor \U$40219 ( \47576_47876 , \15089_15388 , \15644_15946 );
xor \U$40220 ( \47577_47877 , \47576_47876 , \16029_16331 );
buf ge007_GF_PartitionCandidate( \47578_47878_nGe007 , \47577_47877 );
buf \U$labaj5713 ( \47579_R_ad_acea908 , \47578_47878_nGe007 );
xor \U$40222 ( \47580_47880 , \14699_15001 , \15088_15387 );
buf ge009_GF_PartitionCandidate( \47581_47881_nGe009 , \47580_47880 );
buf \U$labaj5714 ( \47582_R_ae_101f8830 , \47581_47881_nGe009 );
xor \U$40224 ( \47583_47883 , \13780_14079 , \14335_14637 );
xor \U$40225 ( \47584_47884 , \47583_47883 , \14696_14998 );
buf ge00c_GF_PartitionCandidate( \47585_47885_nGe00c , \47584_47884 );
buf \U$labaj5715 ( \47586_R_af_f7dec98 , \47585_47885_nGe00c );
xor \U$40227 ( \47587_47887 , \13414_13716 , \13779_14078 );
buf ge00e_GF_PartitionCandidate( \47588_47888_nGe00e , \47587_47887 );
buf \U$labaj5716 ( \47589_R_b0_101e2c50 , \47588_47888_nGe00e );
xor \U$40229 ( \47590_47890 , \12519_12818 , \13074_13376 );
xor \U$40230 ( \47591_47891 , \47590_47890 , \13411_13713 );
buf ge011_GF_PartitionCandidate( \47592_47892_nGe011 , \47591_47891 );
buf \U$labaj5717 ( \47593_R_b1_f801b30 , \47592_47892_nGe011 );
xor \U$40232 ( \47594_47894 , \12177_12479 , \12518_12817 );
buf ge013_GF_PartitionCandidate( \47595_47895_nGe013 , \47594_47894 );
buf \U$labaj5718 ( \47596_R_b2_be16e00 , \47595_47895_nGe013 );
xor \U$40234 ( \47597_47897 , \11306_11605 , \11861_12163 );
xor \U$40235 ( \47598_47898 , \47597_47897 , \12174_12476 );
buf ge016_GF_PartitionCandidate( \47599_47899_nGe016 , \47598_47898 );
buf \U$labaj5719 ( \47600_R_b3_102e3cf0 , \47599_47899_nGe016 );
xor \U$40237 ( \47601_47901 , \10988_11290 , \11305_11604 );
buf ge018_GF_PartitionCandidate( \47602_47902_nGe018 , \47601_47901 );
buf \U$labaj5720 ( \47603_R_b4_10291788 , \47602_47902_nGe018 );
endmodule

