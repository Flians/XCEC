//
// Conformal-LEC Version 20.10-d215 (04-Sep-2020)
//
module top(RIa148a08_33,RIa147bf8_3,RIa148e40_42,RIa148eb8_43,RIa148dc8_41,RIa148fa8_45,RIa148f30_44,RIa149020_46,RIa149098_47,
        RIa149110_48,RIa1480a8_13,RIa148558_23,RIa148a80_34,RIa148030_12,RIa147b80_2,RIa1484e0_22,RIa148af8_35,RIa147fb8_11,RIa147b08_1,
        RIa148468_21,RIa148b70_36,RIa148c60_38,RIa148cd8_39,RIa148d50_40,RIa1485d0_24,RIa147c70_4,RIa148120_14,RIa148198_15,RIa147ce8_5,
        RIa148648_25,RIa148210_16,RIa147d60_6,RIa1486c0_26,RIa1487b0_28,RIa147e50_8,RIa148300_18,RIa1483f0_20,RIa147f40_10,RIa1488a0_30,
        RIa148378_19,RIa147ec8_9,RIa148828_29,RIa148288_17,RIa147dd8_7,RIa148738_27,RIa148be8_37,RIa148990_32,RIa148918_31,R_31_942fc58,
        R_32_942fd00,R_33_942fda8,R_34_942fe50,R_35_942fef8,R_36_942ffa0,R_37_9430048,R_38_94300f0,R_39_9430198,R_3a_9430240,R_3b_94302e8,
        R_3c_9430390);
input RIa148a08_33,RIa147bf8_3,RIa148e40_42,RIa148eb8_43,RIa148dc8_41,RIa148fa8_45,RIa148f30_44,RIa149020_46,RIa149098_47,
        RIa149110_48,RIa1480a8_13,RIa148558_23,RIa148a80_34,RIa148030_12,RIa147b80_2,RIa1484e0_22,RIa148af8_35,RIa147fb8_11,RIa147b08_1,
        RIa148468_21,RIa148b70_36,RIa148c60_38,RIa148cd8_39,RIa148d50_40,RIa1485d0_24,RIa147c70_4,RIa148120_14,RIa148198_15,RIa147ce8_5,
        RIa148648_25,RIa148210_16,RIa147d60_6,RIa1486c0_26,RIa1487b0_28,RIa147e50_8,RIa148300_18,RIa1483f0_20,RIa147f40_10,RIa1488a0_30,
        RIa148378_19,RIa147ec8_9,RIa148828_29,RIa148288_17,RIa147dd8_7,RIa148738_27,RIa148be8_37,RIa148990_32,RIa148918_31;
output R_31_942fc58,R_32_942fd00,R_33_942fda8,R_34_942fe50,R_35_942fef8,R_36_942ffa0,R_37_9430048,R_38_94300f0,R_39_9430198,
        R_3a_9430240,R_3b_94302e8,R_3c_9430390;

wire \61_ZERO , \62_ONE , \63 , \64 , \65 , \66 , \67 , \68 , \69 ,
         \70 , \71 , \72 , \73 , \74 , \75 , \76 , \77 , \78 , \79 ,
         \80 , \81 , \82 , \83_nG93 , \84 , \85 , \86 , \87 , \88 , \89 ,
         \90 , \91 , \92_nG9b , \93 , \94 , \95 , \96 , \97 , \98 , \99 ,
         \100 , \101_nGa3 , \102 , \103 , \104 , \105 , \106 , \107 , \108 , \109 ,
         \110 , \111 , \112 , \113 , \114 , \115 , \116 , \117 , \118 , \119 ,
         \120 , \121 , \122 , \123_nG8b , \124 , \125 , \126 , \127 , \128 , \129 ,
         \130 , \131 , \132 , \133 , \134_nG83 , \135 , \136 , \137 , \138 , \139 ,
         \140 , \141 , \142 , \143_nG7b , \144 , \145 , \146 , \147 , \148 , \149 ,
         \150 , \151 , \152 , \153 , \154_nG6b , \155 , \156 , \157 , \158 , \159 ,
         \160 , \161 , \162_nG5b , \163 , \164 , \165 , \166 , \167 , \168 , \169 ,
         \170 , \171_nG63 , \172 , \173 , \174 , \175 , \176 , \177 , \178 , \179 ,
         \180_nG73 , \181 , \182 , \183 , \184 , \185 , \186 , \187 , \188 , \189 ,
         \190 , \191 , \192 , \193 , \194 , \195 , \196 , \197 , \198 , \199 ,
         \200 , \201 , \202 , \203 , \204 , \205 , \206 , \207 , \208 , \209 ,
         \210 , \211 , \212 , \213 , \214 , \215 , \216 , \217 , \218 , \219 ,
         \220 , \221 , \222 , \223 , \224 , \225 , \226 , \227 , \228 , \229 ,
         \230 , \231 , \232 , \233 , \234 , \235 , \236 , \237 , \238 , \239 ,
         \240 , \241 , \242 , \243 , \244 , \245 , \246 , \247 , \248 , \249 ,
         \250 , \251 , \252 , \253 , \254 , \255 , \256 , \257 , \258 , \259 ,
         \260 , \261 , \262 , \263 , \264 , \265 , \266 , \267 , \268 , \269 ,
         \270 , \271 , \272 , \273 , \274 , \275 , \276 , \277 , \278 , \279 ,
         \280 , \281 , \282 , \283 , \284 , \285 , \286 , \287 , \288 , \289 ,
         \290 , \291 , \292 , \293 , \294 , \295 , \296 , \297 , \298 , \299 ,
         \300 , \301 , \302 , \303 , \304 , \305 , \306 , \307 , \308 , \309 ,
         \310 , \311 , \312 , \313 , \314 , \315 , \316 , \317 , \318 , \319 ,
         \320 , \321 , \322 , \323 , \324 , \325 , \326 , \327 , \328 , \329 ,
         \330 , \331 , \332 , \333 , \334 , \335 , \336 , \337 , \338 , \339 ,
         \340 , \341 , \342 , \343 , \344 , \345 , \346 , \347 , \348 , \349 ,
         \350 , \351 , \352 , \353 , \354 , \355 , \356 , \357 , \358 , \359 ,
         \360 , \361 , \362 , \363 , \364 , \365 , \366 , \367 , \368 , \369 ,
         \370 , \371 , \372 , \373 , \374 , \375 , \376 , \377 , \378 , \379 ,
         \380 , \381 , \382 , \383 , \384 , \385 , \386 , \387 , \388 , \389 ,
         \390 , \391 , \392 , \393 , \394 , \395 , \396 , \397 , \398 , \399 ,
         \400 , \401 , \402 , \403 , \404 , \405 , \406 , \407 , \408 , \409 ,
         \410 , \411 , \412 , \413 , \414 , \415 , \416 , \417 , \418 , \419 ,
         \420 , \421 , \422 , \423 , \424 , \425 , \426 , \427 , \428 , \429 ,
         \430 , \431 , \432 , \433 , \434 , \435 , \436 , \437 , \438 , \439 ,
         \440 , \441 , \442 , \443 , \444 , \445 , \446 , \447 , \448 , \449 ,
         \450 , \451 , \452 , \453 , \454 , \455 , \456 , \457 , \458 , \459 ,
         \460 , \461 , \462 , \463 , \464 , \465 , \466 , \467 , \468 , \469 ,
         \470 , \471 , \472 , \473 , \474 , \475 , \476 , \477 , \478 , \479 ,
         \480 , \481 , \482 , \483 , \484 , \485 , \486 , \487 , \488 , \489 ,
         \490 , \491 , \492 , \493 , \494 , \495 , \496 , \497 , \498 , \499 ,
         \500 , \501 , \502 , \503 , \504 , \505 , \506 , \507 , \508 , \509 ,
         \510 , \511 , \512 , \513 , \514 , \515 , \516 , \517 , \518 , \519 ,
         \520 , \521 , \522 , \523 , \524 , \525 , \526 , \527 , \528 , \529 ,
         \530 , \531 , \532 , \533 , \534 , \535 , \536 , \537 , \538 , \539 ,
         \540 , \541 , \542 , \543 , \544 , \545 , \546 , \547 , \548 , \549 ,
         \550 , \551 , \552 , \553 , \554 , \555 , \556 , \557 , \558 , \559 ,
         \560 , \561 , \562 , \563 , \564 , \565 , \566 , \567 , \568 , \569 ,
         \570 , \571 , \572 , \573 , \574 , \575 , \576 , \577 , \578 , \579 ,
         \580 , \581 , \582 , \583 , \584 , \585 , \586 , \587 , \588 , \589 ,
         \590 , \591 , \592 , \593 , \594 , \595 , \596 , \597 , \598 , \599 ,
         \600 , \601 , \602 , \603 , \604 , \605 , \606 , \607 , \608 , \609 ,
         \610 , \611 , \612 , \613 , \614 , \615 , \616 , \617 , \618 , \619 ,
         \620 , \621 , \622 , \623 , \624 , \625 , \626 , \627 , \628 , \629 ,
         \630 , \631 , \632 , \633 , \634 , \635 , \636 , \637 , \638 , \639 ,
         \640 , \641 , \642 , \643 , \644 , \645 , \646 , \647 , \648 , \649 ,
         \650 , \651 , \652 , \653 , \654 , \655 , \656 , \657 , \658 , \659 ,
         \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 , \668 , \669 ,
         \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677 , \678 , \679 ,
         \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 , \688 , \689 ,
         \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 ,
         \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 ,
         \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 ,
         \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 ,
         \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 ,
         \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 ,
         \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 ,
         \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 ,
         \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 ,
         \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 ,
         \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 ,
         \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 ,
         \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 ,
         \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 ,
         \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 ,
         \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 ,
         \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 ,
         \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 ,
         \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 ,
         \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 ,
         \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 ,
         \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 ,
         \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 ,
         \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 ,
         \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 ,
         \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 ,
         \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 ,
         \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 ,
         \970 , \971 , \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 ,
         \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 ,
         \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 , \998 , \999 ,
         \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 ,
         \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 ,
         \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 ,
         \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 ,
         \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 ,
         \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 ,
         \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 ,
         \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 ,
         \1080 , \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 ,
         \1090 , \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 ,
         \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 ,
         \1110 , \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 ,
         \1120 , \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 ,
         \1130 , \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 ,
         \1140 , \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 ,
         \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 ,
         \1160 , \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 ,
         \1170 , \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 ,
         \1180 , \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 ,
         \1190 , \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 ,
         \1200 , \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 ;
buf \U$labajz134 ( R_31_942fc58, \1177 );
buf \U$labajz135 ( R_32_942fd00, \1183 );
buf \U$labajz136 ( R_33_942fda8, \1185 );
buf \U$labajz137 ( R_34_942fe50, \1187 );
buf \U$labajz138 ( R_35_942fef8, \1189 );
buf \U$labajz139 ( R_36_942ffa0, \1191 );
buf \U$labajz140 ( R_37_9430048, \1193 );
buf \U$labajz141 ( R_38_94300f0, \1195 );
buf \U$labajz142 ( R_39_9430198, \1200 );
buf \U$labajz143 ( R_3a_9430240, \1203 );
buf \U$labajz144 ( R_3b_94302e8, \1205 );
buf \U$labajz145 ( R_3c_9430390, \1207 );
not \U$1 ( \63 , RIa147bf8_3);
or \U$2 ( \64 , RIa148e40_42, RIa148eb8_43, RIa148dc8_41, RIa148fa8_45);
nor \U$3 ( \65 , \64 , RIa148f30_44, RIa149020_46);
not \U$4 ( \66 , \65 );
nor \U$5 ( \67 , \66 , RIa149098_47, RIa149110_48);
not \U$6 ( \68 , \67 );
or \U$7 ( \69 , \63 , \68 );
not \U$8 ( \70 , RIa149110_48);
nor \U$9 ( \71 , \70 , \66 , RIa149098_47);
and \U$10 ( \72 , \71 , RIa1480a8_13);
not \U$11 ( \73 , \66 );
nand \U$12 ( \74 , \73 , RIa149098_47);
nor \U$13 ( \75 , \74 , RIa149110_48);
and \U$14 ( \76 , RIa148558_23, \75 );
nor \U$15 ( \77 , \72 , \76 );
nand \U$16 ( \78 , \69 , \77 );
not \U$17 ( \79 , RIa149110_48);
not \U$18 ( \80 , RIa149098_47);
or \U$19 ( \81 , \79 , \80 );
nand \U$20 ( \82 , \81 , \65 );
_DC g93 ( \83_nG93 , \78 , \82 );
nand \U$21 ( \84 , RIa148a08_33, \83_nG93 );
not \U$22 ( \85 , RIa148030_12);
not \U$23 ( \86 , \71 );
or \U$24 ( \87 , \85 , \86 );
and \U$25 ( \88 , \67 , RIa147b80_2);
and \U$26 ( \89 , RIa1484e0_22, \75 );
nor \U$27 ( \90 , \88 , \89 );
nand \U$28 ( \91 , \87 , \90 );
_DC g9b ( \92_nG9b , \91 , \82 );
nand \U$29 ( \93 , RIa148a80_34, \92_nG9b );
not \U$30 ( \94 , RIa147fb8_11);
not \U$31 ( \95 , \71 );
or \U$32 ( \96 , \94 , \95 );
and \U$33 ( \97 , \67 , RIa147b08_1);
and \U$34 ( \98 , RIa148468_21, \75 );
nor \U$35 ( \99 , \97 , \98 );
nand \U$36 ( \100 , \96 , \99 );
_DC ga3 ( \101_nGa3 , \100 , \82 );
nand \U$37 ( \102 , RIa148af8_35, \101_nGa3 );
not \U$38 ( \103 , \101_nGa3 );
not \U$39 ( \104 , RIa148b70_36);
nor \U$40 ( \105 , \103 , \104 );
nand \U$41 ( \106 , RIa148c60_38, \101_nGa3 );
nand \U$42 ( \107 , RIa148cd8_39, \92_nG9b );
nand \U$43 ( \108 , RIa148d50_40, \101_nGa3 );
xor \U$44 ( \109 , \107 , \108 );
not \U$45 ( \110 , \109 );
nand \U$46 ( \111 , RIa148d50_40, \92_nG9b );
nand \U$47 ( \112 , RIa148cd8_39, \83_nG93 );
xor \U$48 ( \113 , \111 , \112 );
not \U$49 ( \114 , \113 );
nand \U$50 ( \115 , RIa148d50_40, \83_nG93 );
not \U$51 ( \116 , RIa1485d0_24);
not \U$52 ( \117 , \75 );
or \U$53 ( \118 , \116 , \117 );
and \U$54 ( \119 , \67 , RIa147c70_4);
and \U$55 ( \120 , RIa148120_14, \71 );
nor \U$56 ( \121 , \119 , \120 );
nand \U$57 ( \122 , \118 , \121 );
_DC g8b ( \123_nG8b , \122 , \82 );
nand \U$58 ( \124 , RIa148cd8_39, \123_nG8b );
xor \U$59 ( \125 , \115 , \124 );
not \U$60 ( \126 , \125 );
not \U$61 ( \127 , RIa148198_15);
not \U$62 ( \128 , \71 );
or \U$63 ( \129 , \127 , \128 );
and \U$64 ( \130 , \67 , RIa147ce8_5);
and \U$65 ( \131 , RIa148648_25, \75 );
nor \U$66 ( \132 , \130 , \131 );
nand \U$67 ( \133 , \129 , \132 );
_DC g83 ( \134_nG83 , \133 , \82 );
nand \U$68 ( \135 , RIa148d50_40, \134_nG83 );
not \U$69 ( \136 , RIa148210_16);
not \U$70 ( \137 , \71 );
or \U$71 ( \138 , \136 , \137 );
and \U$72 ( \139 , \67 , RIa147d60_6);
and \U$73 ( \140 , RIa1486c0_26, \75 );
nor \U$74 ( \141 , \139 , \140 );
nand \U$75 ( \142 , \138 , \141 );
_DC g7b ( \143_nG7b , \142 , \82 );
nand \U$76 ( \144 , RIa148cd8_39, \143_nG7b );
xor \U$77 ( \145 , \135 , \144 );
not \U$78 ( \146 , \145 );
not \U$79 ( \147 , RIa1487b0_28);
not \U$80 ( \148 , \75 );
or \U$81 ( \149 , \147 , \148 );
and \U$82 ( \150 , \67 , RIa147e50_8);
and \U$83 ( \151 , RIa148300_18, \71 );
nor \U$84 ( \152 , \150 , \151 );
nand \U$85 ( \153 , \149 , \152 );
_DC g6b ( \154_nG6b , \153 , \82 );
not \U$86 ( \155 , RIa1483f0_20);
not \U$87 ( \156 , \71 );
or \U$88 ( \157 , \155 , \156 );
and \U$89 ( \158 , \67 , RIa147f40_10);
and \U$90 ( \159 , RIa1488a0_30, \75 );
nor \U$91 ( \160 , \158 , \159 );
nand \U$92 ( \161 , \157 , \160 );
_DC g5b ( \162_nG5b , \161 , \82 );
or \U$93 ( \163 , \154_nG6b , \162_nG5b );
not \U$94 ( \164 , RIa148378_19);
not \U$95 ( \165 , \71 );
or \U$96 ( \166 , \164 , \165 );
and \U$97 ( \167 , \67 , RIa147ec8_9);
and \U$98 ( \168 , RIa148828_29, \75 );
nor \U$99 ( \169 , \167 , \168 );
nand \U$100 ( \170 , \166 , \169 );
_DC g63 ( \171_nG63 , \170 , \82 );
nand \U$101 ( \172 , \163 , \171_nG63 );
not \U$102 ( \173 , RIa148288_17);
not \U$103 ( \174 , \71 );
or \U$104 ( \175 , \173 , \174 );
and \U$105 ( \176 , \67 , RIa147dd8_7);
and \U$106 ( \177 , RIa148738_27, \75 );
nor \U$107 ( \178 , \176 , \177 );
nand \U$108 ( \179 , \175 , \178 );
_DC g73 ( \180_nG73 , \179 , \82 );
nand \U$109 ( \181 , \154_nG6b , \180_nG73 );
and \U$110 ( \182 , \172 , \181 );
not \U$111 ( \183 , \154_nG6b );
not \U$112 ( \184 , \180_nG73 );
and \U$113 ( \185 , \183 , \184 );
nor \U$114 ( \186 , \182 , \185 );
nand \U$115 ( \187 , \186 , RIa148d50_40, RIa148cd8_39);
not \U$116 ( \188 , \187 );
not \U$117 ( \189 , \188 );
nand \U$118 ( \190 , RIa148d50_40, \143_nG7b );
not \U$119 ( \191 , \190 );
and \U$120 ( \192 , RIa148cd8_39, \180_nG73 );
not \U$121 ( \193 , \192 );
or \U$122 ( \194 , \191 , \193 );
or \U$123 ( \195 , \192 , \190 );
nand \U$124 ( \196 , \194 , \195 );
not \U$125 ( \197 , \196 );
or \U$126 ( \198 , \189 , \197 );
not \U$127 ( \199 , \190 );
nand \U$128 ( \200 , \199 , \192 );
nand \U$129 ( \201 , \198 , \200 );
not \U$130 ( \202 , \201 );
or \U$131 ( \203 , \146 , \202 );
or \U$132 ( \204 , \144 , \135 );
nand \U$133 ( \205 , \203 , \204 );
not \U$134 ( \206 , \205 );
nand \U$135 ( \207 , RIa148cd8_39, \134_nG83 );
nand \U$136 ( \208 , RIa148d50_40, \123_nG8b );
xor \U$137 ( \209 , \207 , \208 );
not \U$138 ( \210 , \209 );
or \U$139 ( \211 , \206 , \210 );
or \U$140 ( \212 , \207 , \208 );
nand \U$141 ( \213 , \211 , \212 );
not \U$142 ( \214 , \213 );
or \U$143 ( \215 , \126 , \214 );
or \U$144 ( \216 , \124 , \115 );
nand \U$145 ( \217 , \215 , \216 );
not \U$146 ( \218 , \217 );
or \U$147 ( \219 , \114 , \218 );
or \U$148 ( \220 , \112 , \111 );
nand \U$149 ( \221 , \219 , \220 );
not \U$150 ( \222 , \221 );
or \U$151 ( \223 , \110 , \222 );
or \U$152 ( \224 , \107 , \108 );
nand \U$153 ( \225 , \223 , \224 );
and \U$154 ( \226 , RIa148cd8_39, \101_nGa3 );
nand \U$155 ( \227 , \225 , \226 );
not \U$156 ( \228 , \227 );
and \U$157 ( \229 , \106 , \228 );
not \U$158 ( \230 , \106 );
and \U$159 ( \231 , \230 , \227 );
or \U$160 ( \232 , \229 , \231 );
not \U$161 ( \233 , \232 );
nand \U$162 ( \234 , RIa148c60_38, \92_nG9b );
xor \U$163 ( \235 , \234 , \226 );
xnor \U$164 ( \236 , \235 , \225 );
not \U$165 ( \237 , \236 );
nand \U$166 ( \238 , RIa148c60_38, \83_nG93 );
xor \U$167 ( \239 , \238 , \109 );
xnor \U$168 ( \240 , \239 , \221 );
not \U$169 ( \241 , \240 );
nand \U$170 ( \242 , RIa148c60_38, \123_nG8b );
xor \U$171 ( \243 , \242 , \113 );
xnor \U$172 ( \244 , \243 , \217 );
not \U$173 ( \245 , \244 );
nand \U$174 ( \246 , RIa148c60_38, \134_nG83 );
xor \U$175 ( \247 , \246 , \125 );
xnor \U$176 ( \248 , \247 , \213 );
not \U$177 ( \249 , \248 );
nand \U$178 ( \250 , RIa148c60_38, \143_nG7b );
xor \U$179 ( \251 , \250 , \209 );
xnor \U$180 ( \252 , \251 , \205 );
not \U$181 ( \253 , \252 );
and \U$182 ( \254 , RIa148c60_38, \180_nG73 );
not \U$183 ( \255 , \254 );
xor \U$184 ( \256 , \201 , \145 );
not \U$185 ( \257 , \256 );
or \U$186 ( \258 , \255 , \257 );
xor \U$187 ( \259 , \254 , \145 );
xnor \U$188 ( \260 , \259 , \201 );
not \U$189 ( \261 , \260 );
nand \U$190 ( \262 , RIa148c60_38, \154_nG6b );
xor \U$191 ( \263 , \262 , \187 );
xnor \U$192 ( \264 , \263 , \196 );
not \U$193 ( \265 , \264 );
not \U$194 ( \266 , \265 );
nand \U$195 ( \267 , RIa148d50_40, \154_nG6b );
not \U$196 ( \268 , \267 );
not \U$197 ( \269 , \268 );
nand \U$198 ( \270 , RIa148cd8_39, \171_nG63 );
not \U$199 ( \271 , \270 );
and \U$200 ( \272 , \269 , \271 );
and \U$201 ( \273 , \268 , \270 );
nor \U$202 ( \274 , \272 , \273 );
nand \U$203 ( \275 , RIa148cd8_39, RIa148d50_40, \171_nG63 , \162_nG5b );
and \U$204 ( \276 , \274 , \275 );
not \U$205 ( \277 , \274 );
nand \U$206 ( \278 , \275 , \171_nG63 );
and \U$207 ( \279 , \277 , \278 );
nor \U$208 ( \280 , \276 , \279 );
not \U$209 ( \281 , \280 );
nand \U$210 ( \282 , RIa148c60_38, \162_nG5b );
not \U$211 ( \283 , \282 );
not \U$212 ( \284 , \283 );
or \U$213 ( \285 , \281 , \284 );
nand \U$214 ( \286 , RIa148c60_38, \171_nG63 );
not \U$215 ( \287 , \286 );
nand \U$216 ( \288 , RIa148d50_40, \162_nG5b );
nor \U$217 ( \289 , \270 , \288 );
not \U$218 ( \290 , \289 );
not \U$219 ( \291 , \274 );
not \U$220 ( \292 , \291 );
or \U$221 ( \293 , \290 , \292 );
and \U$222 ( \294 , \274 , \275 );
nor \U$223 ( \295 , \294 , \282 );
nand \U$224 ( \296 , \293 , \295 );
not \U$225 ( \297 , \296 );
or \U$226 ( \298 , \287 , \297 );
nand \U$227 ( \299 , RIa148cd8_39, \154_nG6b );
nand \U$228 ( \300 , RIa148d50_40, \180_nG73 );
xor \U$229 ( \301 , \299 , \300 );
not \U$230 ( \302 , \301 );
not \U$231 ( \303 , \172 );
nand \U$232 ( \304 , \303 , RIa148d50_40, RIa148cd8_39);
not \U$233 ( \305 , \304 );
not \U$234 ( \306 , \305 );
and \U$235 ( \307 , \302 , \306 );
and \U$236 ( \308 , \301 , \305 );
nor \U$237 ( \309 , \307 , \308 );
buf \U$238 ( \310 , \309 );
nand \U$239 ( \311 , \298 , \310 );
nand \U$240 ( \312 , \285 , \311 );
not \U$241 ( \313 , \312 );
or \U$242 ( \314 , \266 , \313 );
not \U$243 ( \315 , \262 );
and \U$244 ( \316 , \196 , \188 );
not \U$245 ( \317 , \196 );
and \U$246 ( \318 , \317 , \187 );
nor \U$247 ( \319 , \316 , \318 );
nand \U$248 ( \320 , \315 , \319 );
nand \U$249 ( \321 , \314 , \320 );
nand \U$250 ( \322 , \261 , \321 );
nand \U$251 ( \323 , \258 , \322 );
not \U$252 ( \324 , \323 );
or \U$253 ( \325 , \253 , \324 );
not \U$254 ( \326 , \250 );
xor \U$255 ( \327 , \205 , \209 );
nand \U$256 ( \328 , \326 , \327 );
nand \U$257 ( \329 , \325 , \328 );
not \U$258 ( \330 , \329 );
or \U$259 ( \331 , \249 , \330 );
not \U$260 ( \332 , \246 );
xor \U$261 ( \333 , \213 , \125 );
nand \U$262 ( \334 , \332 , \333 );
nand \U$263 ( \335 , \331 , \334 );
not \U$264 ( \336 , \335 );
or \U$265 ( \337 , \245 , \336 );
not \U$266 ( \338 , \242 );
xor \U$267 ( \339 , \217 , \113 );
nand \U$268 ( \340 , \338 , \339 );
nand \U$269 ( \341 , \337 , \340 );
not \U$270 ( \342 , \341 );
or \U$271 ( \343 , \241 , \342 );
not \U$272 ( \344 , \238 );
xor \U$273 ( \345 , \221 , \109 );
nand \U$274 ( \346 , \344 , \345 );
nand \U$275 ( \347 , \343 , \346 );
not \U$276 ( \348 , \347 );
or \U$277 ( \349 , \237 , \348 );
not \U$278 ( \350 , \234 );
xor \U$279 ( \351 , \225 , \226 );
nand \U$280 ( \352 , \350 , \351 );
nand \U$281 ( \353 , \349 , \352 );
not \U$282 ( \354 , \353 );
or \U$283 ( \355 , \233 , \354 );
not \U$284 ( \356 , \106 );
nand \U$285 ( \357 , \356 , \228 );
nand \U$286 ( \358 , \355 , \357 );
nand \U$287 ( \359 , RIa148be8_37, \101_nGa3 );
xnor \U$288 ( \360 , \358 , \359 );
not \U$289 ( \361 , \360 );
nand \U$290 ( \362 , RIa148be8_37, \92_nG9b );
xor \U$291 ( \363 , \362 , \232 );
xnor \U$292 ( \364 , \363 , \353 );
not \U$293 ( \365 , \364 );
nand \U$294 ( \366 , RIa148be8_37, \83_nG93 );
xor \U$295 ( \367 , \366 , \236 );
xnor \U$296 ( \368 , \367 , \347 );
not \U$297 ( \369 , \368 );
nand \U$298 ( \370 , RIa148be8_37, \123_nG8b );
xor \U$299 ( \371 , \370 , \240 );
not \U$300 ( \372 , \341 );
xnor \U$301 ( \373 , \371 , \372 );
not \U$302 ( \374 , \373 );
not \U$303 ( \375 , \374 );
nand \U$304 ( \376 , RIa148be8_37, \134_nG83 );
xor \U$305 ( \377 , \376 , \244 );
xnor \U$306 ( \378 , \377 , \335 );
not \U$307 ( \379 , \378 );
nand \U$308 ( \380 , RIa148be8_37, \143_nG7b );
not \U$309 ( \381 , \248 );
xor \U$310 ( \382 , \380 , \381 );
xor \U$311 ( \383 , \382 , \329 );
not \U$312 ( \384 , \383 );
not \U$313 ( \385 , \312 );
not \U$314 ( \386 , \264 );
and \U$315 ( \387 , \385 , \386 );
and \U$316 ( \388 , \312 , \264 );
nor \U$317 ( \389 , \387 , \388 );
not \U$318 ( \390 , \389 );
nand \U$319 ( \391 , RIa148be8_37, \171_nG63 );
not \U$320 ( \392 , \391 );
and \U$321 ( \393 , \390 , \392 );
and \U$322 ( \394 , \389 , \391 );
buf \U$323 ( \395 , \296 );
not \U$324 ( \396 , \286 );
not \U$325 ( \397 , \309 );
or \U$326 ( \398 , \396 , \397 );
or \U$327 ( \399 , \286 , \309 );
nand \U$328 ( \400 , \398 , \399 );
xnor \U$329 ( \401 , \395 , \400 );
nand \U$330 ( \402 , RIa148be8_37, \162_nG5b );
not \U$331 ( \403 , \402 );
nand \U$332 ( \404 , \401 , \403 );
nor \U$333 ( \405 , \394 , \404 );
nor \U$334 ( \406 , \393 , \405 );
not \U$335 ( \407 , \406 );
nand \U$336 ( \408 , RIa148be8_37, \154_nG6b );
xor \U$337 ( \409 , \408 , \260 );
not \U$338 ( \410 , \321 );
xnor \U$339 ( \411 , \409 , \410 );
nand \U$340 ( \412 , \407 , \411 );
not \U$341 ( \413 , \408 );
xor \U$342 ( \414 , \410 , \260 );
nand \U$343 ( \415 , \413 , \414 );
nand \U$344 ( \416 , \412 , \415 );
not \U$345 ( \417 , \416 );
nand \U$346 ( \418 , RIa148be8_37, \180_nG73 );
xor \U$347 ( \419 , \418 , \252 );
xnor \U$348 ( \420 , \419 , \323 );
not \U$349 ( \421 , \420 );
or \U$350 ( \422 , \417 , \421 );
not \U$351 ( \423 , \418 );
xor \U$352 ( \424 , \323 , \252 );
nand \U$353 ( \425 , \423 , \424 );
nand \U$354 ( \426 , \422 , \425 );
not \U$355 ( \427 , \426 );
or \U$356 ( \428 , \384 , \427 );
not \U$357 ( \429 , \380 );
and \U$358 ( \430 , \329 , \248 );
not \U$359 ( \431 , \329 );
and \U$360 ( \432 , \431 , \381 );
nor \U$361 ( \433 , \430 , \432 );
nand \U$362 ( \434 , \429 , \433 );
nand \U$363 ( \435 , \428 , \434 );
not \U$364 ( \436 , \435 );
or \U$365 ( \437 , \379 , \436 );
not \U$366 ( \438 , \376 );
xor \U$367 ( \439 , \335 , \244 );
nand \U$368 ( \440 , \438 , \439 );
nand \U$369 ( \441 , \437 , \440 );
not \U$370 ( \442 , \441 );
or \U$371 ( \443 , \375 , \442 );
not \U$372 ( \444 , \370 );
not \U$373 ( \445 , \240 );
not \U$374 ( \446 , \372 );
or \U$375 ( \447 , \445 , \446 );
or \U$376 ( \448 , \372 , \240 );
nand \U$377 ( \449 , \447 , \448 );
nand \U$378 ( \450 , \444 , \449 );
nand \U$379 ( \451 , \443 , \450 );
not \U$380 ( \452 , \451 );
or \U$381 ( \453 , \369 , \452 );
not \U$382 ( \454 , \366 );
xor \U$383 ( \455 , \347 , \236 );
nand \U$384 ( \456 , \454 , \455 );
nand \U$385 ( \457 , \453 , \456 );
not \U$386 ( \458 , \457 );
or \U$387 ( \459 , \365 , \458 );
not \U$388 ( \460 , \362 );
not \U$389 ( \461 , \232 );
not \U$390 ( \462 , \353 );
not \U$391 ( \463 , \462 );
or \U$392 ( \464 , \461 , \463 );
or \U$393 ( \465 , \462 , \232 );
nand \U$394 ( \466 , \464 , \465 );
nand \U$395 ( \467 , \460 , \466 );
nand \U$396 ( \468 , \459 , \467 );
not \U$397 ( \469 , \468 );
or \U$398 ( \470 , \361 , \469 );
not \U$399 ( \471 , \359 );
nand \U$400 ( \472 , \471 , \358 );
nand \U$401 ( \473 , \470 , \472 );
xnor \U$402 ( \474 , \105 , \473 );
not \U$403 ( \475 , \474 );
not \U$404 ( \476 , \475 );
nand \U$405 ( \477 , RIa148b70_36, \92_nG9b );
xor \U$406 ( \478 , \477 , \360 );
xnor \U$407 ( \479 , \478 , \468 );
not \U$408 ( \480 , \479 );
nand \U$409 ( \481 , RIa148b70_36, \83_nG93 );
xor \U$410 ( \482 , \481 , \364 );
xnor \U$411 ( \483 , \482 , \457 );
not \U$412 ( \484 , \483 );
nand \U$413 ( \485 , RIa148b70_36, \134_nG83 );
xor \U$414 ( \486 , \485 , \373 );
xnor \U$415 ( \487 , \486 , \441 );
not \U$416 ( \488 , \487 );
not \U$417 ( \489 , \488 );
nand \U$418 ( \490 , RIa148b70_36, \143_nG7b );
xor \U$419 ( \491 , \490 , \378 );
xnor \U$420 ( \492 , \491 , \435 );
not \U$421 ( \493 , \492 );
nand \U$422 ( \494 , RIa148b70_36, \180_nG73 );
xor \U$423 ( \495 , \494 , \383 );
xnor \U$424 ( \496 , \495 , \426 );
not \U$425 ( \497 , \496 );
nand \U$426 ( \498 , RIa148b70_36, \154_nG6b );
xor \U$427 ( \499 , \498 , \416 );
xnor \U$428 ( \500 , \499 , \420 );
not \U$429 ( \501 , \500 );
xor \U$430 ( \502 , \391 , \404 );
xnor \U$431 ( \503 , \502 , \389 );
nand \U$432 ( \504 , RIa148b70_36, \162_nG5b );
not \U$433 ( \505 , \504 );
and \U$434 ( \506 , \503 , \505 );
not \U$435 ( \507 , \171_nG63 );
nor \U$436 ( \508 , \104 , \507 );
xor \U$437 ( \509 , \506 , \508 );
and \U$438 ( \510 , \411 , \407 );
not \U$439 ( \511 , \411 );
and \U$440 ( \512 , \511 , \406 );
nor \U$441 ( \513 , \510 , \512 );
and \U$442 ( \514 , \509 , \513 );
and \U$443 ( \515 , \506 , \508 );
or \U$444 ( \516 , \514 , \515 );
not \U$445 ( \517 , \516 );
or \U$446 ( \518 , \501 , \517 );
not \U$447 ( \519 , \498 );
xor \U$448 ( \520 , \420 , \416 );
nand \U$449 ( \521 , \519 , \520 );
nand \U$450 ( \522 , \518 , \521 );
not \U$451 ( \523 , \522 );
or \U$452 ( \524 , \497 , \523 );
not \U$453 ( \525 , \494 );
xor \U$454 ( \526 , \426 , \383 );
nand \U$455 ( \527 , \525 , \526 );
nand \U$456 ( \528 , \524 , \527 );
not \U$457 ( \529 , \528 );
or \U$458 ( \530 , \493 , \529 );
not \U$459 ( \531 , \490 );
xor \U$460 ( \532 , \378 , \435 );
nand \U$461 ( \533 , \531 , \532 );
nand \U$462 ( \534 , \530 , \533 );
not \U$463 ( \535 , \534 );
or \U$464 ( \536 , \489 , \535 );
not \U$465 ( \537 , \485 );
and \U$466 ( \538 , \441 , \373 );
not \U$467 ( \539 , \441 );
and \U$468 ( \540 , \539 , \374 );
or \U$469 ( \541 , \538 , \540 );
nand \U$470 ( \542 , \537 , \541 );
nand \U$471 ( \543 , \536 , \542 );
not \U$472 ( \544 , \543 );
nand \U$473 ( \545 , RIa148b70_36, \123_nG8b );
xor \U$474 ( \546 , \545 , \368 );
xnor \U$475 ( \547 , \546 , \451 );
not \U$476 ( \548 , \547 );
or \U$477 ( \549 , \544 , \548 );
not \U$478 ( \550 , \545 );
xor \U$479 ( \551 , \368 , \451 );
nand \U$480 ( \552 , \550 , \551 );
nand \U$481 ( \553 , \549 , \552 );
not \U$482 ( \554 , \553 );
or \U$483 ( \555 , \484 , \554 );
not \U$484 ( \556 , \481 );
xor \U$485 ( \557 , \457 , \364 );
nand \U$486 ( \558 , \556 , \557 );
nand \U$487 ( \559 , \555 , \558 );
not \U$488 ( \560 , \559 );
or \U$489 ( \561 , \480 , \560 );
not \U$490 ( \562 , \477 );
xor \U$491 ( \563 , \468 , \360 );
nand \U$492 ( \564 , \562 , \563 );
nand \U$493 ( \565 , \561 , \564 );
not \U$494 ( \566 , \565 );
or \U$495 ( \567 , \476 , \566 );
nand \U$496 ( \568 , \473 , \105 );
nand \U$497 ( \569 , \567 , \568 );
xnor \U$498 ( \570 , \102 , \569 );
xor \U$499 ( \571 , \93 , \570 );
nand \U$500 ( \572 , RIa148af8_35, \92_nG9b );
xor \U$501 ( \573 , \572 , \474 );
xnor \U$502 ( \574 , \573 , \565 );
not \U$503 ( \575 , \574 );
not \U$504 ( \576 , \575 );
nand \U$505 ( \577 , RIa148af8_35, \83_nG93 );
xor \U$506 ( \578 , \577 , \479 );
xnor \U$507 ( \579 , \578 , \559 );
not \U$508 ( \580 , \579 );
nand \U$509 ( \581 , RIa148af8_35, \123_nG8b );
xor \U$510 ( \582 , \581 , \483 );
not \U$511 ( \583 , \553 );
xnor \U$512 ( \584 , \582 , \583 );
not \U$513 ( \585 , \584 );
not \U$514 ( \586 , \585 );
nand \U$515 ( \587 , RIa148af8_35, \134_nG83 );
xor \U$516 ( \588 , \587 , \547 );
not \U$517 ( \589 , \543 );
xnor \U$518 ( \590 , \588 , \589 );
not \U$519 ( \591 , \590 );
not \U$520 ( \592 , \591 );
nand \U$521 ( \593 , RIa148af8_35, \143_nG7b );
not \U$522 ( \594 , \593 );
not \U$523 ( \595 , \488 );
not \U$524 ( \596 , \534 );
not \U$525 ( \597 , \596 );
or \U$526 ( \598 , \595 , \597 );
nand \U$527 ( \599 , \534 , \487 );
nand \U$528 ( \600 , \598 , \599 );
not \U$529 ( \601 , \600 );
or \U$530 ( \602 , \594 , \601 );
or \U$531 ( \603 , \593 , \600 );
nand \U$532 ( \604 , \602 , \603 );
not \U$533 ( \605 , \604 );
and \U$534 ( \606 , RIa148af8_35, \171_nG63 );
and \U$535 ( \607 , RIa148af8_35, \162_nG5b );
xor \U$536 ( \608 , \506 , \508 );
xor \U$537 ( \609 , \608 , \513 );
and \U$538 ( \610 , \607 , \609 );
xor \U$539 ( \611 , \606 , \610 );
xor \U$540 ( \612 , \500 , \516 );
and \U$541 ( \613 , \611 , \612 );
and \U$542 ( \614 , \606 , \610 );
or \U$543 ( \615 , \613 , \614 );
not \U$544 ( \616 , \615 );
nand \U$545 ( \617 , RIa148af8_35, \154_nG6b );
xor \U$546 ( \618 , \617 , \522 );
not \U$547 ( \619 , \496 );
xor \U$548 ( \620 , \618 , \619 );
not \U$549 ( \621 , \620 );
or \U$550 ( \622 , \616 , \621 );
not \U$551 ( \623 , \617 );
and \U$552 ( \624 , \522 , \619 );
not \U$553 ( \625 , \522 );
and \U$554 ( \626 , \625 , \496 );
or \U$555 ( \627 , \624 , \626 );
nand \U$556 ( \628 , \623 , \627 );
nand \U$557 ( \629 , \622 , \628 );
not \U$558 ( \630 , \629 );
nand \U$559 ( \631 , RIa148af8_35, \180_nG73 );
not \U$560 ( \632 , \492 );
xor \U$561 ( \633 , \631 , \632 );
not \U$562 ( \634 , \528 );
xnor \U$563 ( \635 , \633 , \634 );
not \U$564 ( \636 , \635 );
or \U$565 ( \637 , \630 , \636 );
not \U$566 ( \638 , \631 );
and \U$567 ( \639 , \634 , \492 );
not \U$568 ( \640 , \634 );
and \U$569 ( \641 , \640 , \632 );
or \U$570 ( \642 , \639 , \641 );
nand \U$571 ( \643 , \638 , \642 );
nand \U$572 ( \644 , \637 , \643 );
not \U$573 ( \645 , \644 );
or \U$574 ( \646 , \605 , \645 );
not \U$575 ( \647 , \593 );
nand \U$576 ( \648 , \647 , \600 );
nand \U$577 ( \649 , \646 , \648 );
not \U$578 ( \650 , \649 );
or \U$579 ( \651 , \592 , \650 );
not \U$580 ( \652 , \587 );
and \U$581 ( \653 , \547 , \589 );
not \U$582 ( \654 , \547 );
and \U$583 ( \655 , \654 , \543 );
or \U$584 ( \656 , \653 , \655 );
nand \U$585 ( \657 , \652 , \656 );
nand \U$586 ( \658 , \651 , \657 );
not \U$587 ( \659 , \658 );
or \U$588 ( \660 , \586 , \659 );
not \U$589 ( \661 , \581 );
and \U$590 ( \662 , \483 , \583 );
not \U$591 ( \663 , \483 );
and \U$592 ( \664 , \663 , \553 );
or \U$593 ( \665 , \662 , \664 );
nand \U$594 ( \666 , \661 , \665 );
nand \U$595 ( \667 , \660 , \666 );
not \U$596 ( \668 , \667 );
or \U$597 ( \669 , \580 , \668 );
not \U$598 ( \670 , \479 );
and \U$599 ( \671 , \559 , \670 );
nor \U$600 ( \672 , \559 , \670 );
or \U$601 ( \673 , \671 , \672 );
not \U$602 ( \674 , \577 );
nand \U$603 ( \675 , \673 , \674 );
nand \U$604 ( \676 , \669 , \675 );
not \U$605 ( \677 , \676 );
or \U$606 ( \678 , \576 , \677 );
not \U$607 ( \679 , \572 );
xnor \U$608 ( \680 , \565 , \474 );
nand \U$609 ( \681 , \679 , \680 );
nand \U$610 ( \682 , \678 , \681 );
xnor \U$611 ( \683 , \571 , \682 );
xor \U$612 ( \684 , \84 , \683 );
nand \U$613 ( \685 , RIa148a80_34, \83_nG93 );
xor \U$614 ( \686 , \685 , \574 );
xnor \U$615 ( \687 , \686 , \676 );
not \U$616 ( \688 , \687 );
not \U$617 ( \689 , \688 );
nand \U$618 ( \690 , RIa148a80_34, \123_nG8b );
xor \U$619 ( \691 , \690 , \579 );
xnor \U$620 ( \692 , \691 , \667 );
not \U$621 ( \693 , \692 );
nand \U$622 ( \694 , RIa148a80_34, \134_nG83 );
not \U$623 ( \695 , \694 );
not \U$624 ( \696 , \585 );
not \U$625 ( \697 , \658 );
not \U$626 ( \698 , \697 );
or \U$627 ( \699 , \696 , \698 );
nand \U$628 ( \700 , \658 , \584 );
nand \U$629 ( \701 , \699 , \700 );
not \U$630 ( \702 , \701 );
or \U$631 ( \703 , \695 , \702 );
or \U$632 ( \704 , \694 , \701 );
nand \U$633 ( \705 , \703 , \704 );
not \U$634 ( \706 , \705 );
not \U$635 ( \707 , RIa148a80_34);
nor \U$636 ( \708 , \507 , \707 );
xor \U$637 ( \709 , \606 , \610 );
xor \U$638 ( \710 , \709 , \612 );
not \U$639 ( \711 , \710 );
nand \U$640 ( \712 , RIa148a80_34, \162_nG5b );
nor \U$641 ( \713 , \711 , \712 );
xor \U$642 ( \714 , \708 , \713 );
xor \U$643 ( \715 , \620 , \615 );
and \U$644 ( \716 , \714 , \715 );
and \U$645 ( \717 , \708 , \713 );
or \U$646 ( \718 , \716 , \717 );
not \U$647 ( \719 , \718 );
nand \U$648 ( \720 , RIa148a80_34, \154_nG6b );
not \U$649 ( \721 , \629 );
xor \U$650 ( \722 , \720 , \721 );
not \U$651 ( \723 , \635 );
xnor \U$652 ( \724 , \722 , \723 );
not \U$653 ( \725 , \724 );
or \U$654 ( \726 , \719 , \725 );
nand \U$655 ( \727 , \635 , \721 );
not \U$656 ( \728 , \727 );
nand \U$657 ( \729 , \723 , \629 );
not \U$658 ( \730 , \729 );
or \U$659 ( \731 , \728 , \730 );
not \U$660 ( \732 , \720 );
nand \U$661 ( \733 , \731 , \732 );
nand \U$662 ( \734 , \726 , \733 );
not \U$663 ( \735 , \734 );
nor \U$664 ( \736 , \184 , \707 );
not \U$665 ( \737 , \736 );
not \U$666 ( \738 , \644 );
not \U$667 ( \739 , \738 );
not \U$668 ( \740 , \604 );
or \U$669 ( \741 , \739 , \740 );
not \U$670 ( \742 , \604 );
nand \U$671 ( \743 , \742 , \644 );
nand \U$672 ( \744 , \741 , \743 );
not \U$673 ( \745 , \744 );
not \U$674 ( \746 , \745 );
or \U$675 ( \747 , \737 , \746 );
not \U$676 ( \748 , \736 );
nand \U$677 ( \749 , \744 , \748 );
nand \U$678 ( \750 , \747 , \749 );
not \U$679 ( \751 , \750 );
or \U$680 ( \752 , \735 , \751 );
nand \U$681 ( \753 , \744 , \736 );
nand \U$682 ( \754 , \752 , \753 );
not \U$683 ( \755 , \754 );
not \U$684 ( \756 , \143_nG7b );
nor \U$685 ( \757 , \707 , \756 );
not \U$686 ( \758 , \757 );
not \U$687 ( \759 , \591 );
not \U$688 ( \760 , \649 );
not \U$689 ( \761 , \760 );
or \U$690 ( \762 , \759 , \761 );
nand \U$691 ( \763 , \649 , \590 );
nand \U$692 ( \764 , \762 , \763 );
not \U$693 ( \765 , \764 );
not \U$694 ( \766 , \765 );
or \U$695 ( \767 , \758 , \766 );
not \U$696 ( \768 , RIa148a80_34);
not \U$697 ( \769 , \143_nG7b );
or \U$698 ( \770 , \768 , \769 );
nand \U$699 ( \771 , \770 , \764 );
nand \U$700 ( \772 , \767 , \771 );
not \U$701 ( \773 , \772 );
or \U$702 ( \774 , \755 , \773 );
nand \U$703 ( \775 , \764 , \757 );
nand \U$704 ( \776 , \774 , \775 );
not \U$705 ( \777 , \776 );
or \U$706 ( \778 , \706 , \777 );
not \U$707 ( \779 , \694 );
not \U$708 ( \780 , \585 );
not \U$709 ( \781 , \697 );
or \U$710 ( \782 , \780 , \781 );
nand \U$711 ( \783 , \782 , \700 );
nand \U$712 ( \784 , \779 , \783 );
nand \U$713 ( \785 , \778 , \784 );
not \U$714 ( \786 , \785 );
or \U$715 ( \787 , \693 , \786 );
not \U$716 ( \788 , \690 );
xor \U$717 ( \789 , \579 , \667 );
nand \U$718 ( \790 , \788 , \789 );
nand \U$719 ( \791 , \787 , \790 );
not \U$720 ( \792 , \791 );
or \U$721 ( \793 , \689 , \792 );
not \U$722 ( \794 , \575 );
nand \U$723 ( \795 , \794 , \676 );
not \U$724 ( \796 , \795 );
not \U$725 ( \797 , \676 );
nand \U$726 ( \798 , \797 , \575 );
not \U$727 ( \799 , \798 );
or \U$728 ( \800 , \796 , \799 );
not \U$729 ( \801 , \685 );
nand \U$730 ( \802 , \800 , \801 );
nand \U$731 ( \803 , \793 , \802 );
xnor \U$732 ( \804 , \684 , \803 );
not \U$733 ( \805 , \804 );
nand \U$734 ( \806 , RIa148a08_33, \134_nG83 );
not \U$735 ( \807 , \692 );
xor \U$736 ( \808 , \806 , \807 );
buf \U$737 ( \809 , \785 );
not \U$738 ( \810 , \809 );
xnor \U$739 ( \811 , \808 , \810 );
not \U$740 ( \812 , \811 );
nand \U$741 ( \813 , RIa148a08_33, \154_nG6b );
xor \U$742 ( \814 , \813 , \734 );
xnor \U$743 ( \815 , \814 , \750 );
not \U$744 ( \816 , \815 );
nand \U$745 ( \817 , RIa148a08_33, \171_nG63 );
not \U$746 ( \818 , \817 );
xnor \U$747 ( \819 , \724 , \718 );
not \U$748 ( \820 , \819 );
or \U$749 ( \821 , \818 , \820 );
xor \U$750 ( \822 , \708 , \713 );
xor \U$751 ( \823 , \822 , \715 );
nand \U$752 ( \824 , RIa148a08_33, \162_nG5b );
not \U$753 ( \825 , \824 );
and \U$754 ( \826 , \823 , \825 );
nand \U$755 ( \827 , \821 , \826 );
or \U$756 ( \828 , \817 , \819 );
nand \U$757 ( \829 , \827 , \828 );
not \U$758 ( \830 , \829 );
or \U$759 ( \831 , \816 , \830 );
not \U$760 ( \832 , \750 );
nand \U$761 ( \833 , \832 , \734 );
not \U$762 ( \834 , \833 );
not \U$763 ( \835 , \734 );
nand \U$764 ( \836 , \835 , \750 );
not \U$765 ( \837 , \836 );
or \U$766 ( \838 , \834 , \837 );
not \U$767 ( \839 , \813 );
nand \U$768 ( \840 , \838 , \839 );
nand \U$769 ( \841 , \831 , \840 );
not \U$770 ( \842 , \841 );
nand \U$771 ( \843 , RIa148a08_33, \180_nG73 );
xor \U$772 ( \844 , \843 , \772 );
xnor \U$773 ( \845 , \844 , \754 );
not \U$774 ( \846 , \845 );
or \U$775 ( \847 , \842 , \846 );
not \U$776 ( \848 , \843 );
not \U$777 ( \849 , \757 );
not \U$778 ( \850 , \765 );
or \U$779 ( \851 , \849 , \850 );
nand \U$780 ( \852 , \851 , \771 );
xor \U$781 ( \853 , \852 , \754 );
nand \U$782 ( \854 , \848 , \853 );
nand \U$783 ( \855 , \847 , \854 );
not \U$784 ( \856 , \855 );
not \U$785 ( \857 , RIa148a08_33);
nor \U$786 ( \858 , \857 , \756 );
not \U$787 ( \859 , \858 );
not \U$788 ( \860 , \705 );
not \U$789 ( \861 , \776 );
not \U$790 ( \862 , \861 );
or \U$791 ( \863 , \860 , \862 );
not \U$792 ( \864 , \705 );
nand \U$793 ( \865 , \864 , \776 );
nand \U$794 ( \866 , \863 , \865 );
not \U$795 ( \867 , \866 );
not \U$796 ( \868 , \867 );
or \U$797 ( \869 , \859 , \868 );
not \U$798 ( \870 , \858 );
nand \U$799 ( \871 , \870 , \866 );
nand \U$800 ( \872 , \869 , \871 );
not \U$801 ( \873 , \872 );
or \U$802 ( \874 , \856 , \873 );
nand \U$803 ( \875 , \866 , \858 );
nand \U$804 ( \876 , \874 , \875 );
not \U$805 ( \877 , \876 );
or \U$806 ( \878 , \812 , \877 );
not \U$807 ( \879 , \806 );
not \U$808 ( \880 , \807 );
not \U$809 ( \881 , \809 );
or \U$810 ( \882 , \880 , \881 );
nand \U$811 ( \883 , \810 , \692 );
nand \U$812 ( \884 , \882 , \883 );
nand \U$813 ( \885 , \879 , \884 );
nand \U$814 ( \886 , \878 , \885 );
not \U$815 ( \887 , \886 );
not \U$816 ( \888 , \687 );
not \U$817 ( \889 , \791 );
or \U$818 ( \890 , \888 , \889 );
or \U$819 ( \891 , \687 , \791 );
nand \U$820 ( \892 , \890 , \891 );
not \U$821 ( \893 , \892 );
nand \U$822 ( \894 , RIa148a08_33, \123_nG8b );
not \U$823 ( \895 , \894 );
and \U$824 ( \896 , \893 , \895 );
and \U$825 ( \897 , \892 , \894 );
nor \U$826 ( \898 , \896 , \897 );
not \U$827 ( \899 , \898 );
not \U$828 ( \900 , \899 );
or \U$829 ( \901 , \887 , \900 );
not \U$830 ( \902 , \894 );
nand \U$831 ( \903 , \902 , \892 );
nand \U$832 ( \904 , \901 , \903 );
not \U$833 ( \905 , \904 );
or \U$834 ( \906 , \805 , \905 );
not \U$835 ( \907 , \84 );
not \U$836 ( \908 , \683 );
not \U$837 ( \909 , \908 );
not \U$838 ( \910 , \803 );
or \U$839 ( \911 , \909 , \910 );
or \U$840 ( \912 , \803 , \908 );
nand \U$841 ( \913 , \911 , \912 );
nand \U$842 ( \914 , \907 , \913 );
nand \U$843 ( \915 , \906 , \914 );
not \U$844 ( \916 , \915 );
nand \U$845 ( \917 , RIa148a08_33, \92_nG9b );
not \U$846 ( \918 , \570 );
not \U$847 ( \919 , \682 );
or \U$848 ( \920 , \918 , \919 );
not \U$849 ( \921 , \102 );
nand \U$850 ( \922 , \921 , \569 );
nand \U$851 ( \923 , \920 , \922 );
nand \U$852 ( \924 , RIa148a80_34, \101_nGa3 );
xnor \U$853 ( \925 , \923 , \924 );
xor \U$854 ( \926 , \917 , \925 );
not \U$855 ( \927 , \683 );
not \U$856 ( \928 , \803 );
or \U$857 ( \929 , \927 , \928 );
not \U$858 ( \930 , \93 );
xor \U$859 ( \931 , \682 , \570 );
nand \U$860 ( \932 , \930 , \931 );
nand \U$861 ( \933 , \929 , \932 );
xnor \U$862 ( \934 , \926 , \933 );
not \U$863 ( \935 , \934 );
or \U$864 ( \936 , \916 , \935 );
not \U$865 ( \937 , \917 );
xor \U$866 ( \938 , \933 , \925 );
nand \U$867 ( \939 , \937 , \938 );
nand \U$868 ( \940 , \936 , \939 );
not \U$869 ( \941 , \940 );
not \U$870 ( \942 , \925 );
not \U$871 ( \943 , \933 );
or \U$872 ( \944 , \942 , \943 );
not \U$873 ( \945 , \924 );
nand \U$874 ( \946 , \945 , \923 );
nand \U$875 ( \947 , \944 , \946 );
nand \U$876 ( \948 , RIa148a08_33, \101_nGa3 );
xnor \U$877 ( \949 , \947 , \948 );
not \U$878 ( \950 , \949 );
or \U$879 ( \951 , \941 , \950 );
not \U$880 ( \952 , \948 );
nand \U$881 ( \953 , \952 , \947 );
nand \U$882 ( \954 , \951 , \953 );
nand \U$883 ( \955 , RIa148990_32, \101_nGa3 );
and \U$884 ( \956 , \954 , \955 );
not \U$885 ( \957 , \954 );
not \U$886 ( \958 , \955 );
and \U$887 ( \959 , \957 , \958 );
or \U$888 ( \960 , \956 , \959 );
not \U$889 ( \961 , \960 );
nand \U$890 ( \962 , RIa148990_32, \92_nG9b );
xor \U$891 ( \963 , \962 , \949 );
xnor \U$892 ( \964 , \963 , \940 );
not \U$893 ( \965 , \964 );
nand \U$894 ( \966 , RIa148990_32, \83_nG93 );
not \U$895 ( \967 , \934 );
xor \U$896 ( \968 , \966 , \967 );
xor \U$897 ( \969 , \968 , \915 );
not \U$898 ( \970 , \969 );
xor \U$899 ( \971 , \817 , \826 );
xnor \U$900 ( \972 , \971 , \819 );
nand \U$901 ( \973 , RIa148990_32, \162_nG5b );
nor \U$902 ( \974 , \972 , \973 );
and \U$903 ( \975 , RIa148990_32, \171_nG63 );
xor \U$904 ( \976 , \974 , \975 );
xor \U$905 ( \977 , \815 , \829 );
and \U$906 ( \978 , \976 , \977 );
and \U$907 ( \979 , \974 , \975 );
or \U$908 ( \980 , \978 , \979 );
not \U$909 ( \981 , \980 );
nand \U$910 ( \982 , RIa148990_32, \154_nG6b );
xor \U$911 ( \983 , \982 , \841 );
xnor \U$912 ( \984 , \983 , \845 );
not \U$913 ( \985 , \984 );
or \U$914 ( \986 , \981 , \985 );
not \U$915 ( \987 , \845 );
nand \U$916 ( \988 , \987 , \841 );
not \U$917 ( \989 , \988 );
not \U$918 ( \990 , \841 );
nand \U$919 ( \991 , \990 , \845 );
not \U$920 ( \992 , \991 );
or \U$921 ( \993 , \989 , \992 );
not \U$922 ( \994 , \982 );
nand \U$923 ( \995 , \993 , \994 );
nand \U$924 ( \996 , \986 , \995 );
not \U$925 ( \997 , \996 );
nand \U$926 ( \998 , RIa148990_32, \180_nG73 );
not \U$927 ( \999 , \872 );
xor \U$928 ( \1000 , \998 , \999 );
not \U$929 ( \1001 , \855 );
xnor \U$930 ( \1002 , \1000 , \1001 );
not \U$931 ( \1003 , \1002 );
or \U$932 ( \1004 , \997 , \1003 );
not \U$933 ( \1005 , \1001 );
nand \U$934 ( \1006 , \1005 , \999 );
not \U$935 ( \1007 , \1006 );
not \U$936 ( \1008 , \999 );
nand \U$937 ( \1009 , \1008 , \1001 );
not \U$938 ( \1010 , \1009 );
or \U$939 ( \1011 , \1007 , \1010 );
not \U$940 ( \1012 , \998 );
nand \U$941 ( \1013 , \1011 , \1012 );
nand \U$942 ( \1014 , \1004 , \1013 );
not \U$943 ( \1015 , \1014 );
not \U$944 ( \1016 , RIa148990_32);
nor \U$945 ( \1017 , \1016 , \756 );
not \U$946 ( \1018 , \1017 );
xor \U$947 ( \1019 , \811 , \876 );
not \U$948 ( \1020 , \1019 );
not \U$949 ( \1021 , \1020 );
or \U$950 ( \1022 , \1018 , \1021 );
not \U$951 ( \1023 , \1017 );
nand \U$952 ( \1024 , \1023 , \1019 );
nand \U$953 ( \1025 , \1022 , \1024 );
not \U$954 ( \1026 , \1025 );
or \U$955 ( \1027 , \1015 , \1026 );
nand \U$956 ( \1028 , \1019 , \1017 );
nand \U$957 ( \1029 , \1027 , \1028 );
not \U$958 ( \1030 , \1029 );
not \U$959 ( \1031 , \898 );
not \U$960 ( \1032 , \886 );
or \U$961 ( \1033 , \1031 , \1032 );
or \U$962 ( \1034 , \898 , \886 );
nand \U$963 ( \1035 , \1033 , \1034 );
not \U$964 ( \1036 , \1035 );
nand \U$965 ( \1037 , RIa148990_32, \134_nG83 );
not \U$966 ( \1038 , \1037 );
and \U$967 ( \1039 , \1036 , \1038 );
and \U$968 ( \1040 , \1035 , \1037 );
nor \U$969 ( \1041 , \1039 , \1040 );
not \U$970 ( \1042 , \1041 );
not \U$971 ( \1043 , \1042 );
or \U$972 ( \1044 , \1030 , \1043 );
not \U$973 ( \1045 , \1037 );
nand \U$974 ( \1046 , \1045 , \1035 );
nand \U$975 ( \1047 , \1044 , \1046 );
nand \U$976 ( \1048 , RIa148990_32, \123_nG8b );
xor \U$977 ( \1049 , \1048 , \804 );
xnor \U$978 ( \1050 , \1049 , \904 );
nand \U$979 ( \1051 , \1047 , \1050 );
not \U$980 ( \1052 , \1048 );
xor \U$981 ( \1053 , \904 , \804 );
nand \U$982 ( \1054 , \1052 , \1053 );
nand \U$983 ( \1055 , \1051 , \1054 );
not \U$984 ( \1056 , \1055 );
or \U$985 ( \1057 , \970 , \1056 );
not \U$986 ( \1058 , \966 );
xnor \U$987 ( \1059 , \915 , \967 );
nand \U$988 ( \1060 , \1058 , \1059 );
nand \U$989 ( \1061 , \1057 , \1060 );
not \U$990 ( \1062 , \1061 );
or \U$991 ( \1063 , \965 , \1062 );
not \U$992 ( \1064 , \962 );
xor \U$993 ( \1065 , \940 , \949 );
nand \U$994 ( \1066 , \1064 , \1065 );
nand \U$995 ( \1067 , \1063 , \1066 );
not \U$996 ( \1068 , \1067 );
or \U$997 ( \1069 , \961 , \1068 );
nand \U$998 ( \1070 , \954 , \958 );
nand \U$999 ( \1071 , \1069 , \1070 );
nand \U$1000 ( \1072 , RIa148918_31, \101_nGa3 );
xor \U$1001 ( \1073 , \1071 , \1072 );
not \U$1002 ( \1074 , \1073 );
not \U$1003 ( \1075 , \1074 );
nand \U$1004 ( \1076 , RIa148918_31, \123_nG8b );
xor \U$1005 ( \1077 , \1076 , \969 );
xnor \U$1006 ( \1078 , \1077 , \1055 );
not \U$1007 ( \1079 , \1078 );
nand \U$1008 ( \1080 , RIa148918_31, \134_nG83 );
xor \U$1009 ( \1081 , \1080 , \1050 );
xnor \U$1010 ( \1082 , \1081 , \1047 );
not \U$1011 ( \1083 , \1082 );
nand \U$1012 ( \1084 , RIa148918_31, \171_nG63 );
not \U$1013 ( \1085 , \1084 );
xor \U$1014 ( \1086 , \980 , \984 );
not \U$1015 ( \1087 , \1086 );
not \U$1016 ( \1088 , \1087 );
or \U$1017 ( \1089 , \1085 , \1088 );
and \U$1018 ( \1090 , RIa148918_31, \162_nG5b );
xor \U$1019 ( \1091 , \974 , \975 );
xor \U$1020 ( \1092 , \1091 , \977 );
and \U$1021 ( \1093 , \1090 , \1092 );
nand \U$1022 ( \1094 , \1089 , \1093 );
not \U$1023 ( \1095 , \1084 );
nand \U$1024 ( \1096 , \1095 , \1086 );
and \U$1025 ( \1097 , \1094 , \1096 );
not \U$1026 ( \1098 , \1097 );
not \U$1027 ( \1099 , \1098 );
nand \U$1028 ( \1100 , RIa148918_31, \154_nG6b );
xor \U$1029 ( \1101 , \1100 , \996 );
xnor \U$1030 ( \1102 , \1101 , \1002 );
not \U$1031 ( \1103 , \1102 );
or \U$1032 ( \1104 , \1099 , \1103 );
not \U$1033 ( \1105 , \1100 );
xor \U$1034 ( \1106 , \1002 , \996 );
nand \U$1035 ( \1107 , \1105 , \1106 );
nand \U$1036 ( \1108 , \1104 , \1107 );
not \U$1037 ( \1109 , \1108 );
nand \U$1038 ( \1110 , RIa148918_31, \180_nG73 );
xor \U$1039 ( \1111 , \1110 , \1025 );
xnor \U$1040 ( \1112 , \1111 , \1014 );
not \U$1041 ( \1113 , \1112 );
or \U$1042 ( \1114 , \1109 , \1113 );
not \U$1043 ( \1115 , \1110 );
xor \U$1044 ( \1116 , \1025 , \1014 );
nand \U$1045 ( \1117 , \1115 , \1116 );
nand \U$1046 ( \1118 , \1114 , \1117 );
not \U$1047 ( \1119 , \1118 );
nand \U$1048 ( \1120 , RIa148918_31, \143_nG7b );
xor \U$1049 ( \1121 , \1120 , \1041 );
not \U$1050 ( \1122 , \1029 );
xnor \U$1051 ( \1123 , \1121 , \1122 );
not \U$1052 ( \1124 , \1123 );
or \U$1053 ( \1125 , \1119 , \1124 );
not \U$1054 ( \1126 , \1120 );
not \U$1055 ( \1127 , \1029 );
not \U$1056 ( \1128 , \1041 );
or \U$1057 ( \1129 , \1127 , \1128 );
nand \U$1058 ( \1130 , \1122 , \1042 );
nand \U$1059 ( \1131 , \1129 , \1130 );
nand \U$1060 ( \1132 , \1126 , \1131 );
nand \U$1061 ( \1133 , \1125 , \1132 );
not \U$1062 ( \1134 , \1133 );
or \U$1063 ( \1135 , \1083 , \1134 );
not \U$1064 ( \1136 , \1050 );
nand \U$1065 ( \1137 , \1136 , \1047 );
not \U$1066 ( \1138 , \1137 );
not \U$1067 ( \1139 , \1047 );
nand \U$1068 ( \1140 , \1139 , \1050 );
not \U$1069 ( \1141 , \1140 );
or \U$1070 ( \1142 , \1138 , \1141 );
not \U$1071 ( \1143 , \1080 );
nand \U$1072 ( \1144 , \1142 , \1143 );
nand \U$1073 ( \1145 , \1135 , \1144 );
not \U$1074 ( \1146 , \1145 );
or \U$1075 ( \1147 , \1079 , \1146 );
not \U$1076 ( \1148 , \1076 );
xor \U$1077 ( \1149 , \969 , \1055 );
nand \U$1078 ( \1150 , \1148 , \1149 );
nand \U$1079 ( \1151 , \1147 , \1150 );
not \U$1080 ( \1152 , \1151 );
nand \U$1081 ( \1153 , RIa148918_31, \83_nG93 );
xor \U$1082 ( \1154 , \1153 , \964 );
xnor \U$1083 ( \1155 , \1154 , \1061 );
not \U$1084 ( \1156 , \1155 );
or \U$1085 ( \1157 , \1152 , \1156 );
not \U$1086 ( \1158 , \1153 );
xor \U$1087 ( \1159 , \964 , \1061 );
nand \U$1088 ( \1160 , \1158 , \1159 );
nand \U$1089 ( \1161 , \1157 , \1160 );
not \U$1090 ( \1162 , \1161 );
nand \U$1091 ( \1163 , RIa148918_31, \92_nG9b );
xor \U$1092 ( \1164 , \1163 , \960 );
xnor \U$1093 ( \1165 , \1164 , \1067 );
not \U$1094 ( \1166 , \1165 );
or \U$1095 ( \1167 , \1162 , \1166 );
not \U$1096 ( \1168 , \1163 );
xor \U$1097 ( \1169 , \960 , \1067 );
nand \U$1098 ( \1170 , \1168 , \1169 );
nand \U$1099 ( \1171 , \1167 , \1170 );
not \U$1100 ( \1172 , \1171 );
or \U$1101 ( \1173 , \1075 , \1172 );
not \U$1102 ( \1174 , \1072 );
nand \U$1103 ( \1175 , \1174 , \1071 );
nand \U$1104 ( \1176 , \1173 , \1175 );
buf \U$1105 ( \1177 , \1176 );
not \U$1106 ( \1178 , \1073 );
not \U$1107 ( \1179 , \1171 );
or \U$1108 ( \1180 , \1178 , \1179 );
or \U$1109 ( \1181 , \1171 , \1073 );
nand \U$1110 ( \1182 , \1180 , \1181 );
buf \U$1111 ( \1183 , \1182 );
xor \U$1112 ( \1184 , \1165 , \1161 );
buf \U$1113 ( \1185 , \1184 );
xor \U$1114 ( \1186 , \1155 , \1151 );
buf \U$1115 ( \1187 , \1186 );
xor \U$1116 ( \1188 , \1078 , \1145 );
buf \U$1117 ( \1189 , \1188 );
xor \U$1118 ( \1190 , \1082 , \1133 );
buf \U$1119 ( \1191 , \1190 );
xor \U$1120 ( \1192 , \1123 , \1118 );
buf \U$1121 ( \1193 , \1192 );
xor \U$1122 ( \1194 , \1108 , \1112 );
buf \U$1123 ( \1195 , \1194 );
and \U$1124 ( \1196 , \1102 , \1098 );
not \U$1125 ( \1197 , \1102 );
and \U$1126 ( \1198 , \1197 , \1097 );
nor \U$1127 ( \1199 , \1196 , \1198 );
buf \U$1128 ( \1200 , \1199 );
xor \U$1129 ( \1201 , \1084 , \1093 );
xnor \U$1130 ( \1202 , \1201 , \1086 );
buf \U$1131 ( \1203 , \1202 );
xor \U$1132 ( \1204 , \1090 , \1092 );
buf \U$1133 ( \1205 , \1204 );
xor \U$1134 ( \1206 , \973 , \972 );
buf \U$1135 ( \1207 , \1206 );
endmodule

