//
// Conformal-LEC Version 20.10-d207 (02-Sep-2020)
//
module top(i1,i2,i3,i4,i5,i6,i7,i8,i9,
        i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
        i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
        i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
        i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
        i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
        i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
        i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
        i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
        i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
        i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
        i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
        i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
        i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
        i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
        i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
        i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
        i170,i171,i172,i173,i174,i175,i176,i177,i178,i179,
        i180,i181,i182,i183,i184,i185,i186,i187,i188,i189,
        i190,i191,i192,i193,i194,i195,i196,i197,i198,i199,
        i200,i201,i202,i203,i204,i205,i206,i207,i208,i209,
        i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,
        i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,
        i230,i231,i232,i233,i234,i235,i236,i237,i238,i239,
        i240,i241,i242,i243,i244,i245,i246,i247,i248,i249,
        i250,i251,i252,i253,i254,i255,i256,i257,i258,i259,
        i260,i261,i262,i263,i264,i265,i266,i267,i268,i269,
        i270,i271,i272,i273,i274,i275,i276,i277,i278,i279,
        i280,i281,i282,i283,i284,i285,i286,i287,i288,i289,
        i290,i291,i292,i293,i294,i295,i296,i297,i298,i299,
        i300,i301,i302,i303,i304,i305,i306,i307,i308,i309,
        i310,i311,i312,i313,i314,i315,i316,i317,i318,i319,
        i320,i321,i322,i323,i324,i325,i326,i327,i328,i329,
        i330,i331,i332,i333,i334,i335,i336,i337,i338,i339,
        i340,i341,i342,i343,i344,i345,i346,i347,i348,i349,
        i350,i351,i352,i353,i354,i355,i356,i357,i358,i359,
        i360,i361,i362,i363,i364,i365,i366,i367,i368,i369,
        i370,i371,i372,i373,i374,i375,i376,i377,i378,i379,
        i380,i381,i382,i383,i384,i385,i386,i387,i388,i389,
        i390,i391,i392,i393,i394,i395,i396,i397,i398,i399,
        i400,i401,i402,i403,i404,i405,i406,i407,i408,i409,
        i410,i411,i412,i413,i414,i415,i416,i417,i418,i419,
        i420,i421,i422,i423,i424,i425,i426,i427,i428,i429,
        i430,i431,i432,i433,i434,i435,i436,i437,i438,i439,
        i440,i441,i442,i443,i444,i445,i446,i447,i448,i449,
        i450,i451,i452,i453,i454,i455,i456,i457,i458,i459,
        i460,i461,i462,i463,i464,i465,i466,i467,i468,i469,
        i470,i471,i472,i473,i474,i475,i476,i477,i478,i479,
        i480,i481,i482,i483,i484,i485,i486,i487,i488,i489,
        i490,i491,i492,i493,i494,i495,i496,i497,i498,i499,
        i500,i501,i502,i503,i504,i505,i506,i507,i508,i509,
        i510,i511,i512,i513,i514,i515,i516,i517,i518,i519,
        i520,i521,i522,i523,i524,i525,i526,i527,i528,i529,
        i530,i531,i532,i533,i534,i535,i536,i537,i538,i539,
        i540,i541,i542,i543,i544,i545,i546,i547,i548,i549,
        i550,i551,i552,i553,i554,i555,i556,i557,i558,i559,
        i560,i561,i562,i563,i564,i565,i566,i567,i568,i569,
        i570,i571,i572,i573,i574,i575,i576,i577,i578,i579,
        i580,i581,i582,i583,i584,i585,i586,i587,i588,i589,
        i590,i591,i592,i593,i594,i595,i596,i597,i598,i599,
        i600,i601,i602,i603,i604,i605,i606,i607,i608,i609,
        i610,i611,i612,i613,i614,i615,i616,i617,i618,i619,
        i620,i621,i622,i623,i624,i625,i626,i627,i628,i629,
        i630,i631,i632,i633,i634,i635,i636,i637,i638,i639,
        i640,i641,i642,i643,i644,i645,i646,i647,i648,i649,
        i650,i651,i652,i653,i654,i655,i656,i657,i658,i659,
        i660,i661,i662,i663,i664,i665,i666,i667,i668,i669,
        i670,i671,i672,i673,i674,i675,i676,i677,i678,i679,
        i680,i681,i682,i683,i684,i685,i686,i687,i688,i689,
        i690,i691,i692,i693,i694,i695,i696,i697,i698,i699,
        i700,i701,i702,i703,i704,i705,i706,i707,i708,i709,
        i710,i711,i712,i713,i714,i715,i716,i717,i718,i719,
        i720,i721,i722,i723,i724,i725,i726,i727,i728,i729,
        i730,i731,i732,i733,i734,i735,i736,i737,i738,i739,
        i740,i741,i742,i743,i744,i745,i746,i747,i748,i749,
        i750,i751,i752,i753,i754,i755,i756,i757,i758,i759,
        i760,i761,i762,i763,i764,i765,i766,i767,i768,i769,
        i770,i771,i772,i773,i774,i775,i776,i777,i778,i779,
        i780,i781,i782,i783,i784,i785,i786,i787,i788,i789,
        i790,i791,i792,i793,i794,i795,i796,i797,i798,i799,
        i800,i801,i802,i803,i804,i805,i806,i807,i808,i809,
        i810,i811,i812,i813,i814,i815,i816,i817,i818,i819,
        i820,i821,i822,i823,i824,i825,i826,i827,i828,i829,
        i830,i831,i832,i833,i834,i835,i836,i837,i838,i839,
        i840,i841,i842,i843,i844,i845,i846,i847,i848,i849,
        i850,i851,i852,i853,i854,i855,i856,i857,i858,i859,
        i860,i861,i862,i863,i864,i865,i866,i867,i868,i869,
        i870,i871,i872,i873,i874,i875,i876,i877,i878,i879,
        i880,i881,i882,i883,i884,i885,i886,i887,i888,i889,
        i890,i891,i892,i893,i894,i895,i896,i897,i898,i899,
        i900,i901,i902,i903,i904,i905,i906,i907,i908,i909,
        i910,i911,i912,i913,i914,i915,i916,i917,i918,i919,
        i920,i921,i922,i923,i924,i925,i926,i927,i928,i929,
        i930,i931,i932,i933,i934,i935,i936,i937,i938,i939,
        i940,i941,i942,i943,i944,i945,i946,i947,i948,i949,
        i950,i951,i952,i953,i954,i955,i956,i957,i958,i959,
        i960,i961,i962,i963,i964,i965,i966,i967,i968,i969,
        i970,i971,i972,i973,i974,i975,i976,i977,i978,i979,
        i980,i981,i982,i983,i984,i985,i986,i987,i988,i989,
        i990,i991,i992,i993,i994,i995,i996,i997,i998,i999,
        i1000,i1001,i1002,i1003,i1004,i1005,i1006,i1007,i1008,i1009,
        i1010,i1011,i1012,i1013,i1014,i1015,i1016,i1017,i1018,i1019,
        i1020,i1021,i1022,i1023,i1024,i1025,i1026,i1027,i1028,i1029,
        i1030,i1031,i1032,i1033,i1034,i1035,i1036,i1037,i1038,i1039,
        i1040,i1041,i1042,i1043,i1044,i1045,i1046,i1047,i1048,i1049,
        i1050,i1051,i1052,i1053,i1054,i1055,i1056,i1057,i1058,i1059,
        i1060,i1061,i1062,i1063,i1064,i1065,i1066,i1067,i1068,i1069,
        i1070,i1071,i1072,i1073,i1074,i1075,i1076,i1077,i1078,i1079,
        i1080,i1081,i1082,i1083,i1084,i1085,o1,o2,o3,o4,
        o5,o6,o7,o8,o9);
input i1,i2,i3,i4,i5,i6,i7,i8,i9,
        i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,
        i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,
        i30,i31,i32,i33,i34,i35,i36,i37,i38,i39,
        i40,i41,i42,i43,i44,i45,i46,i47,i48,i49,
        i50,i51,i52,i53,i54,i55,i56,i57,i58,i59,
        i60,i61,i62,i63,i64,i65,i66,i67,i68,i69,
        i70,i71,i72,i73,i74,i75,i76,i77,i78,i79,
        i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,
        i90,i91,i92,i93,i94,i95,i96,i97,i98,i99,
        i100,i101,i102,i103,i104,i105,i106,i107,i108,i109,
        i110,i111,i112,i113,i114,i115,i116,i117,i118,i119,
        i120,i121,i122,i123,i124,i125,i126,i127,i128,i129,
        i130,i131,i132,i133,i134,i135,i136,i137,i138,i139,
        i140,i141,i142,i143,i144,i145,i146,i147,i148,i149,
        i150,i151,i152,i153,i154,i155,i156,i157,i158,i159,
        i160,i161,i162,i163,i164,i165,i166,i167,i168,i169,
        i170,i171,i172,i173,i174,i175,i176,i177,i178,i179,
        i180,i181,i182,i183,i184,i185,i186,i187,i188,i189,
        i190,i191,i192,i193,i194,i195,i196,i197,i198,i199,
        i200,i201,i202,i203,i204,i205,i206,i207,i208,i209,
        i210,i211,i212,i213,i214,i215,i216,i217,i218,i219,
        i220,i221,i222,i223,i224,i225,i226,i227,i228,i229,
        i230,i231,i232,i233,i234,i235,i236,i237,i238,i239,
        i240,i241,i242,i243,i244,i245,i246,i247,i248,i249,
        i250,i251,i252,i253,i254,i255,i256,i257,i258,i259,
        i260,i261,i262,i263,i264,i265,i266,i267,i268,i269,
        i270,i271,i272,i273,i274,i275,i276,i277,i278,i279,
        i280,i281,i282,i283,i284,i285,i286,i287,i288,i289,
        i290,i291,i292,i293,i294,i295,i296,i297,i298,i299,
        i300,i301,i302,i303,i304,i305,i306,i307,i308,i309,
        i310,i311,i312,i313,i314,i315,i316,i317,i318,i319,
        i320,i321,i322,i323,i324,i325,i326,i327,i328,i329,
        i330,i331,i332,i333,i334,i335,i336,i337,i338,i339,
        i340,i341,i342,i343,i344,i345,i346,i347,i348,i349,
        i350,i351,i352,i353,i354,i355,i356,i357,i358,i359,
        i360,i361,i362,i363,i364,i365,i366,i367,i368,i369,
        i370,i371,i372,i373,i374,i375,i376,i377,i378,i379,
        i380,i381,i382,i383,i384,i385,i386,i387,i388,i389,
        i390,i391,i392,i393,i394,i395,i396,i397,i398,i399,
        i400,i401,i402,i403,i404,i405,i406,i407,i408,i409,
        i410,i411,i412,i413,i414,i415,i416,i417,i418,i419,
        i420,i421,i422,i423,i424,i425,i426,i427,i428,i429,
        i430,i431,i432,i433,i434,i435,i436,i437,i438,i439,
        i440,i441,i442,i443,i444,i445,i446,i447,i448,i449,
        i450,i451,i452,i453,i454,i455,i456,i457,i458,i459,
        i460,i461,i462,i463,i464,i465,i466,i467,i468,i469,
        i470,i471,i472,i473,i474,i475,i476,i477,i478,i479,
        i480,i481,i482,i483,i484,i485,i486,i487,i488,i489,
        i490,i491,i492,i493,i494,i495,i496,i497,i498,i499,
        i500,i501,i502,i503,i504,i505,i506,i507,i508,i509,
        i510,i511,i512,i513,i514,i515,i516,i517,i518,i519,
        i520,i521,i522,i523,i524,i525,i526,i527,i528,i529,
        i530,i531,i532,i533,i534,i535,i536,i537,i538,i539,
        i540,i541,i542,i543,i544,i545,i546,i547,i548,i549,
        i550,i551,i552,i553,i554,i555,i556,i557,i558,i559,
        i560,i561,i562,i563,i564,i565,i566,i567,i568,i569,
        i570,i571,i572,i573,i574,i575,i576,i577,i578,i579,
        i580,i581,i582,i583,i584,i585,i586,i587,i588,i589,
        i590,i591,i592,i593,i594,i595,i596,i597,i598,i599,
        i600,i601,i602,i603,i604,i605,i606,i607,i608,i609,
        i610,i611,i612,i613,i614,i615,i616,i617,i618,i619,
        i620,i621,i622,i623,i624,i625,i626,i627,i628,i629,
        i630,i631,i632,i633,i634,i635,i636,i637,i638,i639,
        i640,i641,i642,i643,i644,i645,i646,i647,i648,i649,
        i650,i651,i652,i653,i654,i655,i656,i657,i658,i659,
        i660,i661,i662,i663,i664,i665,i666,i667,i668,i669,
        i670,i671,i672,i673,i674,i675,i676,i677,i678,i679,
        i680,i681,i682,i683,i684,i685,i686,i687,i688,i689,
        i690,i691,i692,i693,i694,i695,i696,i697,i698,i699,
        i700,i701,i702,i703,i704,i705,i706,i707,i708,i709,
        i710,i711,i712,i713,i714,i715,i716,i717,i718,i719,
        i720,i721,i722,i723,i724,i725,i726,i727,i728,i729,
        i730,i731,i732,i733,i734,i735,i736,i737,i738,i739,
        i740,i741,i742,i743,i744,i745,i746,i747,i748,i749,
        i750,i751,i752,i753,i754,i755,i756,i757,i758,i759,
        i760,i761,i762,i763,i764,i765,i766,i767,i768,i769,
        i770,i771,i772,i773,i774,i775,i776,i777,i778,i779,
        i780,i781,i782,i783,i784,i785,i786,i787,i788,i789,
        i790,i791,i792,i793,i794,i795,i796,i797,i798,i799,
        i800,i801,i802,i803,i804,i805,i806,i807,i808,i809,
        i810,i811,i812,i813,i814,i815,i816,i817,i818,i819,
        i820,i821,i822,i823,i824,i825,i826,i827,i828,i829,
        i830,i831,i832,i833,i834,i835,i836,i837,i838,i839,
        i840,i841,i842,i843,i844,i845,i846,i847,i848,i849,
        i850,i851,i852,i853,i854,i855,i856,i857,i858,i859,
        i860,i861,i862,i863,i864,i865,i866,i867,i868,i869,
        i870,i871,i872,i873,i874,i875,i876,i877,i878,i879,
        i880,i881,i882,i883,i884,i885,i886,i887,i888,i889,
        i890,i891,i892,i893,i894,i895,i896,i897,i898,i899,
        i900,i901,i902,i903,i904,i905,i906,i907,i908,i909,
        i910,i911,i912,i913,i914,i915,i916,i917,i918,i919,
        i920,i921,i922,i923,i924,i925,i926,i927,i928,i929,
        i930,i931,i932,i933,i934,i935,i936,i937,i938,i939,
        i940,i941,i942,i943,i944,i945,i946,i947,i948,i949,
        i950,i951,i952,i953,i954,i955,i956,i957,i958,i959,
        i960,i961,i962,i963,i964,i965,i966,i967,i968,i969,
        i970,i971,i972,i973,i974,i975,i976,i977,i978,i979,
        i980,i981,i982,i983,i984,i985,i986,i987,i988,i989,
        i990,i991,i992,i993,i994,i995,i996,i997,i998,i999,
        i1000,i1001,i1002,i1003,i1004,i1005,i1006,i1007,i1008,i1009,
        i1010,i1011,i1012,i1013,i1014,i1015,i1016,i1017,i1018,i1019,
        i1020,i1021,i1022,i1023,i1024,i1025,i1026,i1027,i1028,i1029,
        i1030,i1031,i1032,i1033,i1034,i1035,i1036,i1037,i1038,i1039,
        i1040,i1041,i1042,i1043,i1044,i1045,i1046,i1047,i1048,i1049,
        i1050,i1051,i1052,i1053,i1054,i1055,i1056,i1057,i1058,i1059,
        i1060,i1061,i1062,i1063,i1064,i1065,i1066,i1067,i1068,i1069,
        i1070,i1071,i1072,i1073,i1074,i1075,i1076,i1077,i1078,i1079,
        i1080,i1081,i1082,i1083,i1084,i1085;
output o1,o2,o3,o4,o5,o6,o7,o8,o9;

wire \1095_o1 , \1096_o2 , \1097_o3 , \1098_o4 , \1099_o5 , \1100_o6 , \1101_o7 , \1102_o8 , \1103_o9 ,
         \1104_N$1 , \1105_N$2 , \1106_N$3 , \1107_N$4 , \1108_N$5 , \1109_N$6 , \1110_N$7 , \1111_N$8 , \1112_N$9 , \1113_ZERO ,
         \1114_ONE ;
buf \U$labajz228 ( o1, 1'b0 );
buf \U$labajz229 ( o2, 1'b0 );
buf \U$labajz230 ( o3, 1'b0 );
buf \U$labajz231 ( o4, 1'b0 );
buf \U$labajz232 ( o5, 1'b0 );
buf \U$labajz233 ( o6, 1'b0 );
buf \U$labajz234 ( o7, 1'b0 );
buf \U$labajz235 ( o8, 1'b0 );
buf \U$labajz236 ( o9, 1'b0 );
endmodule

