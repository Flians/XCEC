//
// Conformal-LEC Version 20.10-d215 (04-Sep-2020)
//
module top(RIa139848_33,RIa138a38_3,RIa139c80_42,RIa139cf8_43,RIa139c08_41,RIa139de8_45,RIa139d70_44,RIa139e60_46,RIa139ed8_47,
        RIa139f50_48,RIa138ee8_13,RIa139398_23,RIa1398c0_34,RIa138e70_12,RIa1389c0_2,RIa139320_22,RIa139938_35,RIa138df8_11,RIa138948_1,
        RIa1392a8_21,RIa1399b0_36,RIa139aa0_38,RIa139b18_39,RIa139b90_40,RIa139410_24,RIa138ab0_4,RIa138f60_14,RIa138fd8_15,RIa138b28_5,
        RIa139488_25,RIa139050_16,RIa138ba0_6,RIa139500_26,RIa1395f0_28,RIa138c90_8,RIa139140_18,RIa139230_20,RIa138d80_10,RIa1396e0_30,
        RIa1391b8_19,RIa138d08_9,RIa139668_29,RIa1390c8_17,RIa138c18_7,RIa139578_27,RIa139a28_37,RIa1397d0_32,RIa139758_31,R_31_942aab8,
        R_32_942ab60,R_33_942ac08,R_34_942acb0,R_35_942ad58,R_36_942ae00,R_37_942aea8,R_38_942af50,R_39_942aff8,R_3a_942b0a0,R_3b_942b148,
        R_3c_942b1f0,R_3d_942b298,R_3e_942b340,R_3f_942b3e8,R_40_942b490,R_41_942b538,R_42_942b5e0,R_43_942b688,R_44_942b730);
input RIa139848_33,RIa138a38_3,RIa139c80_42,RIa139cf8_43,RIa139c08_41,RIa139de8_45,RIa139d70_44,RIa139e60_46,RIa139ed8_47,
        RIa139f50_48,RIa138ee8_13,RIa139398_23,RIa1398c0_34,RIa138e70_12,RIa1389c0_2,RIa139320_22,RIa139938_35,RIa138df8_11,RIa138948_1,
        RIa1392a8_21,RIa1399b0_36,RIa139aa0_38,RIa139b18_39,RIa139b90_40,RIa139410_24,RIa138ab0_4,RIa138f60_14,RIa138fd8_15,RIa138b28_5,
        RIa139488_25,RIa139050_16,RIa138ba0_6,RIa139500_26,RIa1395f0_28,RIa138c90_8,RIa139140_18,RIa139230_20,RIa138d80_10,RIa1396e0_30,
        RIa1391b8_19,RIa138d08_9,RIa139668_29,RIa1390c8_17,RIa138c18_7,RIa139578_27,RIa139a28_37,RIa1397d0_32,RIa139758_31;
output R_31_942aab8,R_32_942ab60,R_33_942ac08,R_34_942acb0,R_35_942ad58,R_36_942ae00,R_37_942aea8,R_38_942af50,R_39_942aff8,
        R_3a_942b0a0,R_3b_942b148,R_3c_942b1f0,R_3d_942b298,R_3e_942b340,R_3f_942b3e8,R_40_942b490,R_41_942b538,R_42_942b5e0,R_43_942b688,
        R_44_942b730;

wire \69_ZERO , \70_ONE , \71 , \72 , \73 , \74 , \75 , \76 , \77 ,
         \78 , \79 , \80 , \81 , \82 , \83 , \84 , \85 , \86 , \87 ,
         \88 , \89 , \90 , \91_nG93 , \92 , \93 , \94 , \95 , \96 , \97 ,
         \98 , \99 , \100_nG9b , \101 , \102 , \103 , \104 , \105 , \106 , \107 ,
         \108 , \109_nGa3 , \110 , \111 , \112 , \113 , \114 , \115 , \116 , \117 ,
         \118 , \119 , \120 , \121 , \122 , \123 , \124 , \125 , \126 , \127 ,
         \128 , \129 , \130 , \131_nG8b , \132 , \133 , \134 , \135 , \136 , \137 ,
         \138 , \139 , \140 , \141 , \142_nG83 , \143 , \144 , \145 , \146 , \147 ,
         \148 , \149 , \150 , \151_nG7b , \152 , \153 , \154 , \155 , \156 , \157 ,
         \158 , \159 , \160 , \161 , \162_nG6b , \163 , \164 , \165 , \166 , \167 ,
         \168 , \169 , \170_nG5b , \171 , \172 , \173 , \174 , \175 , \176 , \177 ,
         \178 , \179_nG63 , \180 , \181 , \182 , \183 , \184 , \185 , \186 , \187 ,
         \188_nG73 , \189 , \190 , \191 , \192 , \193 , \194 , \195 , \196 , \197 ,
         \198 , \199 , \200 , \201 , \202 , \203 , \204 , \205 , \206 , \207 ,
         \208 , \209 , \210 , \211 , \212 , \213 , \214 , \215 , \216 , \217 ,
         \218 , \219 , \220 , \221 , \222 , \223 , \224 , \225 , \226 , \227 ,
         \228 , \229 , \230 , \231 , \232 , \233 , \234 , \235 , \236 , \237 ,
         \238 , \239 , \240 , \241 , \242 , \243 , \244 , \245 , \246 , \247 ,
         \248 , \249 , \250 , \251 , \252 , \253 , \254 , \255 , \256 , \257 ,
         \258 , \259 , \260 , \261 , \262 , \263 , \264 , \265 , \266 , \267 ,
         \268 , \269 , \270 , \271 , \272 , \273 , \274 , \275 , \276 , \277 ,
         \278 , \279 , \280 , \281 , \282 , \283 , \284 , \285 , \286 , \287 ,
         \288 , \289 , \290 , \291 , \292 , \293 , \294 , \295 , \296 , \297 ,
         \298 , \299 , \300 , \301 , \302 , \303 , \304 , \305 , \306 , \307 ,
         \308 , \309 , \310 , \311 , \312 , \313 , \314 , \315 , \316 , \317 ,
         \318 , \319 , \320 , \321 , \322 , \323 , \324 , \325 , \326 , \327 ,
         \328 , \329 , \330 , \331 , \332 , \333 , \334 , \335 , \336 , \337 ,
         \338 , \339 , \340 , \341 , \342 , \343 , \344 , \345 , \346 , \347 ,
         \348 , \349 , \350 , \351 , \352 , \353 , \354 , \355 , \356 , \357 ,
         \358 , \359 , \360 , \361 , \362 , \363 , \364 , \365 , \366 , \367 ,
         \368 , \369 , \370 , \371 , \372 , \373 , \374 , \375 , \376 , \377 ,
         \378 , \379 , \380 , \381 , \382 , \383 , \384 , \385 , \386 , \387 ,
         \388 , \389 , \390 , \391 , \392 , \393 , \394 , \395 , \396 , \397 ,
         \398 , \399 , \400 , \401 , \402 , \403 , \404 , \405 , \406 , \407 ,
         \408 , \409 , \410 , \411 , \412 , \413 , \414 , \415 , \416 , \417 ,
         \418 , \419 , \420 , \421 , \422 , \423 , \424 , \425 , \426 , \427 ,
         \428 , \429 , \430 , \431 , \432 , \433 , \434 , \435 , \436 , \437 ,
         \438 , \439 , \440 , \441 , \442 , \443 , \444 , \445 , \446 , \447 ,
         \448 , \449 , \450 , \451 , \452 , \453 , \454 , \455 , \456 , \457 ,
         \458 , \459 , \460 , \461 , \462 , \463 , \464 , \465 , \466 , \467 ,
         \468 , \469 , \470 , \471 , \472 , \473 , \474 , \475 , \476 , \477 ,
         \478 , \479 , \480 , \481 , \482 , \483 , \484 , \485 , \486 , \487 ,
         \488 , \489 , \490 , \491 , \492 , \493 , \494 , \495 , \496 , \497 ,
         \498 , \499 , \500 , \501 , \502 , \503 , \504 , \505 , \506 , \507 ,
         \508 , \509 , \510 , \511 , \512 , \513 , \514 , \515 , \516 , \517 ,
         \518 , \519 , \520 , \521 , \522 , \523 , \524 , \525 , \526 , \527 ,
         \528 , \529 , \530 , \531 , \532 , \533 , \534 , \535 , \536 , \537 ,
         \538 , \539 , \540 , \541 , \542 , \543 , \544 , \545 , \546 , \547 ,
         \548 , \549 , \550 , \551 , \552 , \553 , \554 , \555 , \556 , \557 ,
         \558 , \559 , \560 , \561 , \562 , \563 , \564 , \565 , \566 , \567 ,
         \568 , \569 , \570 , \571 , \572 , \573 , \574 , \575 , \576 , \577 ,
         \578 , \579 , \580 , \581 , \582 , \583 , \584 , \585 , \586 , \587 ,
         \588 , \589 , \590 , \591 , \592 , \593 , \594 , \595 , \596 , \597 ,
         \598 , \599 , \600 , \601 , \602 , \603 , \604 , \605 , \606 , \607 ,
         \608 , \609 , \610 , \611 , \612 , \613 , \614 , \615 , \616 , \617 ,
         \618 , \619 , \620 , \621 , \622 , \623 , \624 , \625 , \626 , \627 ,
         \628 , \629 , \630 , \631 , \632 , \633 , \634 , \635 , \636 , \637 ,
         \638 , \639 , \640 , \641 , \642 , \643 , \644 , \645 , \646 , \647 ,
         \648 , \649 , \650 , \651 , \652 , \653 , \654 , \655 , \656 , \657 ,
         \658 , \659 , \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 ,
         \668 , \669 , \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677 ,
         \678 , \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 ,
         \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 ,
         \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 ,
         \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 ,
         \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 ,
         \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 ,
         \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 ,
         \748 , \749 , \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 ,
         \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 ,
         \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 ,
         \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 ,
         \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 ,
         \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 ,
         \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 ,
         \818 , \819 , \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 ,
         \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 ,
         \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 ,
         \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 ,
         \858 , \859 , \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 ,
         \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 ,
         \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 ,
         \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 ,
         \898 , \899 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 ,
         \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 ,
         \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 ,
         \928 , \929 , \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937 ,
         \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 ,
         \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 ,
         \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 ,
         \968 , \969 , \970 , \971 , \972 , \973 , \974 , \975 , \976 , \977 ,
         \978 , \979 , \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 ,
         \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 ,
         \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 ,
         \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 ,
         \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 ,
         \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 ,
         \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 ,
         \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 ,
         \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 ,
         \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 ,
         \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 ,
         \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 ,
         \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 ,
         \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 ,
         \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 ,
         \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 ,
         \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 ,
         \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 ,
         \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 ,
         \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 ,
         \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 ,
         \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 ,
         \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 ,
         \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 ,
         \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 ,
         \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 ,
         \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 ,
         \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 ,
         \1258 ;
buf \U$labajz140 ( R_31_942aab8, \1185 );
buf \U$labajz141 ( R_32_942ab60, \1191 );
buf \U$labajz142 ( R_33_942ac08, \1193 );
buf \U$labajz143 ( R_34_942acb0, \1195 );
buf \U$labajz144 ( R_35_942ad58, \1197 );
buf \U$labajz145 ( R_36_942ae00, \1199 );
buf \U$labajz146 ( R_37_942aea8, \1201 );
buf \U$labajz147 ( R_38_942af50, \1203 );
buf \U$labajz148 ( R_39_942aff8, \1208 );
buf \U$labajz149 ( R_3a_942b0a0, \1211 );
buf \U$labajz150 ( R_3b_942b148, \1213 );
buf \U$labajz151 ( R_3c_942b1f0, \1215 );
buf \U$labajz152 ( R_3d_942b298, \1217 );
buf \U$labajz153 ( R_3e_942b340, \1223 );
buf \U$labajz154 ( R_3f_942b3e8, \1225 );
buf \U$labajz155 ( R_40_942b490, \1232 );
buf \U$labajz156 ( R_41_942b538, \1239 );
buf \U$labajz157 ( R_42_942b5e0, \1248 );
buf \U$labajz158 ( R_43_942b688, \1256 );
buf \U$labajz159 ( R_44_942b730, \1258 );
not \U$1 ( \71 , RIa138a38_3);
or \U$2 ( \72 , RIa139c80_42, RIa139cf8_43, RIa139c08_41, RIa139de8_45);
nor \U$3 ( \73 , \72 , RIa139d70_44, RIa139e60_46);
not \U$4 ( \74 , \73 );
nor \U$5 ( \75 , \74 , RIa139ed8_47, RIa139f50_48);
not \U$6 ( \76 , \75 );
or \U$7 ( \77 , \71 , \76 );
not \U$8 ( \78 , RIa139f50_48);
nor \U$9 ( \79 , \78 , \74 , RIa139ed8_47);
and \U$10 ( \80 , \79 , RIa138ee8_13);
not \U$11 ( \81 , \74 );
nand \U$12 ( \82 , \81 , RIa139ed8_47);
nor \U$13 ( \83 , \82 , RIa139f50_48);
and \U$14 ( \84 , RIa139398_23, \83 );
nor \U$15 ( \85 , \80 , \84 );
nand \U$16 ( \86 , \77 , \85 );
not \U$17 ( \87 , RIa139f50_48);
not \U$18 ( \88 , RIa139ed8_47);
or \U$19 ( \89 , \87 , \88 );
nand \U$20 ( \90 , \89 , \73 );
_DC g93 ( \91_nG93 , \86 , \90 );
nand \U$21 ( \92 , RIa139848_33, \91_nG93 );
not \U$22 ( \93 , RIa138e70_12);
not \U$23 ( \94 , \79 );
or \U$24 ( \95 , \93 , \94 );
and \U$25 ( \96 , \75 , RIa1389c0_2);
and \U$26 ( \97 , RIa139320_22, \83 );
nor \U$27 ( \98 , \96 , \97 );
nand \U$28 ( \99 , \95 , \98 );
_DC g9b ( \100_nG9b , \99 , \90 );
nand \U$29 ( \101 , RIa1398c0_34, \100_nG9b );
not \U$30 ( \102 , RIa138df8_11);
not \U$31 ( \103 , \79 );
or \U$32 ( \104 , \102 , \103 );
and \U$33 ( \105 , \75 , RIa138948_1);
and \U$34 ( \106 , RIa1392a8_21, \83 );
nor \U$35 ( \107 , \105 , \106 );
nand \U$36 ( \108 , \104 , \107 );
_DC ga3 ( \109_nGa3 , \108 , \90 );
nand \U$37 ( \110 , RIa139938_35, \109_nGa3 );
not \U$38 ( \111 , \109_nGa3 );
not \U$39 ( \112 , RIa1399b0_36);
nor \U$40 ( \113 , \111 , \112 );
nand \U$41 ( \114 , RIa139aa0_38, \109_nGa3 );
nand \U$42 ( \115 , RIa139b18_39, \100_nG9b );
nand \U$43 ( \116 , RIa139b90_40, \109_nGa3 );
xor \U$44 ( \117 , \115 , \116 );
not \U$45 ( \118 , \117 );
nand \U$46 ( \119 , RIa139b90_40, \100_nG9b );
nand \U$47 ( \120 , RIa139b18_39, \91_nG93 );
xor \U$48 ( \121 , \119 , \120 );
not \U$49 ( \122 , \121 );
nand \U$50 ( \123 , RIa139b90_40, \91_nG93 );
not \U$51 ( \124 , RIa139410_24);
not \U$52 ( \125 , \83 );
or \U$53 ( \126 , \124 , \125 );
and \U$54 ( \127 , \75 , RIa138ab0_4);
and \U$55 ( \128 , RIa138f60_14, \79 );
nor \U$56 ( \129 , \127 , \128 );
nand \U$57 ( \130 , \126 , \129 );
_DC g8b ( \131_nG8b , \130 , \90 );
nand \U$58 ( \132 , RIa139b18_39, \131_nG8b );
xor \U$59 ( \133 , \123 , \132 );
not \U$60 ( \134 , \133 );
not \U$61 ( \135 , RIa138fd8_15);
not \U$62 ( \136 , \79 );
or \U$63 ( \137 , \135 , \136 );
and \U$64 ( \138 , \75 , RIa138b28_5);
and \U$65 ( \139 , RIa139488_25, \83 );
nor \U$66 ( \140 , \138 , \139 );
nand \U$67 ( \141 , \137 , \140 );
_DC g83 ( \142_nG83 , \141 , \90 );
nand \U$68 ( \143 , RIa139b90_40, \142_nG83 );
not \U$69 ( \144 , RIa139050_16);
not \U$70 ( \145 , \79 );
or \U$71 ( \146 , \144 , \145 );
and \U$72 ( \147 , \75 , RIa138ba0_6);
and \U$73 ( \148 , RIa139500_26, \83 );
nor \U$74 ( \149 , \147 , \148 );
nand \U$75 ( \150 , \146 , \149 );
_DC g7b ( \151_nG7b , \150 , \90 );
nand \U$76 ( \152 , RIa139b18_39, \151_nG7b );
xor \U$77 ( \153 , \143 , \152 );
not \U$78 ( \154 , \153 );
not \U$79 ( \155 , RIa1395f0_28);
not \U$80 ( \156 , \83 );
or \U$81 ( \157 , \155 , \156 );
and \U$82 ( \158 , \75 , RIa138c90_8);
and \U$83 ( \159 , RIa139140_18, \79 );
nor \U$84 ( \160 , \158 , \159 );
nand \U$85 ( \161 , \157 , \160 );
_DC g6b ( \162_nG6b , \161 , \90 );
not \U$86 ( \163 , RIa139230_20);
not \U$87 ( \164 , \79 );
or \U$88 ( \165 , \163 , \164 );
and \U$89 ( \166 , \75 , RIa138d80_10);
and \U$90 ( \167 , RIa1396e0_30, \83 );
nor \U$91 ( \168 , \166 , \167 );
nand \U$92 ( \169 , \165 , \168 );
_DC g5b ( \170_nG5b , \169 , \90 );
or \U$93 ( \171 , \162_nG6b , \170_nG5b );
not \U$94 ( \172 , RIa1391b8_19);
not \U$95 ( \173 , \79 );
or \U$96 ( \174 , \172 , \173 );
and \U$97 ( \175 , \75 , RIa138d08_9);
and \U$98 ( \176 , RIa139668_29, \83 );
nor \U$99 ( \177 , \175 , \176 );
nand \U$100 ( \178 , \174 , \177 );
_DC g63 ( \179_nG63 , \178 , \90 );
nand \U$101 ( \180 , \171 , \179_nG63 );
not \U$102 ( \181 , RIa1390c8_17);
not \U$103 ( \182 , \79 );
or \U$104 ( \183 , \181 , \182 );
and \U$105 ( \184 , \75 , RIa138c18_7);
and \U$106 ( \185 , RIa139578_27, \83 );
nor \U$107 ( \186 , \184 , \185 );
nand \U$108 ( \187 , \183 , \186 );
_DC g73 ( \188_nG73 , \187 , \90 );
nand \U$109 ( \189 , \162_nG6b , \188_nG73 );
and \U$110 ( \190 , \180 , \189 );
not \U$111 ( \191 , \162_nG6b );
not \U$112 ( \192 , \188_nG73 );
and \U$113 ( \193 , \191 , \192 );
nor \U$114 ( \194 , \190 , \193 );
nand \U$115 ( \195 , \194 , RIa139b90_40, RIa139b18_39);
not \U$116 ( \196 , \195 );
not \U$117 ( \197 , \196 );
nand \U$118 ( \198 , RIa139b90_40, \151_nG7b );
not \U$119 ( \199 , \198 );
and \U$120 ( \200 , RIa139b18_39, \188_nG73 );
not \U$121 ( \201 , \200 );
or \U$122 ( \202 , \199 , \201 );
or \U$123 ( \203 , \200 , \198 );
nand \U$124 ( \204 , \202 , \203 );
not \U$125 ( \205 , \204 );
or \U$126 ( \206 , \197 , \205 );
not \U$127 ( \207 , \198 );
nand \U$128 ( \208 , \207 , \200 );
nand \U$129 ( \209 , \206 , \208 );
not \U$130 ( \210 , \209 );
or \U$131 ( \211 , \154 , \210 );
or \U$132 ( \212 , \152 , \143 );
nand \U$133 ( \213 , \211 , \212 );
not \U$134 ( \214 , \213 );
nand \U$135 ( \215 , RIa139b18_39, \142_nG83 );
nand \U$136 ( \216 , RIa139b90_40, \131_nG8b );
xor \U$137 ( \217 , \215 , \216 );
not \U$138 ( \218 , \217 );
or \U$139 ( \219 , \214 , \218 );
or \U$140 ( \220 , \215 , \216 );
nand \U$141 ( \221 , \219 , \220 );
not \U$142 ( \222 , \221 );
or \U$143 ( \223 , \134 , \222 );
or \U$144 ( \224 , \132 , \123 );
nand \U$145 ( \225 , \223 , \224 );
not \U$146 ( \226 , \225 );
or \U$147 ( \227 , \122 , \226 );
or \U$148 ( \228 , \120 , \119 );
nand \U$149 ( \229 , \227 , \228 );
not \U$150 ( \230 , \229 );
or \U$151 ( \231 , \118 , \230 );
or \U$152 ( \232 , \115 , \116 );
nand \U$153 ( \233 , \231 , \232 );
and \U$154 ( \234 , RIa139b18_39, \109_nGa3 );
nand \U$155 ( \235 , \233 , \234 );
not \U$156 ( \236 , \235 );
and \U$157 ( \237 , \114 , \236 );
not \U$158 ( \238 , \114 );
and \U$159 ( \239 , \238 , \235 );
or \U$160 ( \240 , \237 , \239 );
not \U$161 ( \241 , \240 );
nand \U$162 ( \242 , RIa139aa0_38, \100_nG9b );
xor \U$163 ( \243 , \242 , \234 );
xnor \U$164 ( \244 , \243 , \233 );
not \U$165 ( \245 , \244 );
nand \U$166 ( \246 , RIa139aa0_38, \91_nG93 );
xor \U$167 ( \247 , \246 , \117 );
xnor \U$168 ( \248 , \247 , \229 );
not \U$169 ( \249 , \248 );
nand \U$170 ( \250 , RIa139aa0_38, \131_nG8b );
xor \U$171 ( \251 , \250 , \121 );
xnor \U$172 ( \252 , \251 , \225 );
not \U$173 ( \253 , \252 );
nand \U$174 ( \254 , RIa139aa0_38, \142_nG83 );
xor \U$175 ( \255 , \254 , \133 );
xnor \U$176 ( \256 , \255 , \221 );
not \U$177 ( \257 , \256 );
nand \U$178 ( \258 , RIa139aa0_38, \151_nG7b );
xor \U$179 ( \259 , \258 , \217 );
xnor \U$180 ( \260 , \259 , \213 );
not \U$181 ( \261 , \260 );
and \U$182 ( \262 , RIa139aa0_38, \188_nG73 );
not \U$183 ( \263 , \262 );
xor \U$184 ( \264 , \209 , \153 );
not \U$185 ( \265 , \264 );
or \U$186 ( \266 , \263 , \265 );
xor \U$187 ( \267 , \262 , \153 );
xnor \U$188 ( \268 , \267 , \209 );
not \U$189 ( \269 , \268 );
nand \U$190 ( \270 , RIa139aa0_38, \162_nG6b );
xor \U$191 ( \271 , \270 , \195 );
xnor \U$192 ( \272 , \271 , \204 );
not \U$193 ( \273 , \272 );
not \U$194 ( \274 , \273 );
nand \U$195 ( \275 , RIa139b90_40, \162_nG6b );
not \U$196 ( \276 , \275 );
not \U$197 ( \277 , \276 );
nand \U$198 ( \278 , RIa139b18_39, \179_nG63 );
not \U$199 ( \279 , \278 );
and \U$200 ( \280 , \277 , \279 );
and \U$201 ( \281 , \276 , \278 );
nor \U$202 ( \282 , \280 , \281 );
nand \U$203 ( \283 , RIa139b18_39, RIa139b90_40, \179_nG63 , \170_nG5b );
and \U$204 ( \284 , \282 , \283 );
not \U$205 ( \285 , \282 );
nand \U$206 ( \286 , \283 , \179_nG63 );
and \U$207 ( \287 , \285 , \286 );
nor \U$208 ( \288 , \284 , \287 );
not \U$209 ( \289 , \288 );
nand \U$210 ( \290 , RIa139aa0_38, \170_nG5b );
not \U$211 ( \291 , \290 );
not \U$212 ( \292 , \291 );
or \U$213 ( \293 , \289 , \292 );
nand \U$214 ( \294 , RIa139aa0_38, \179_nG63 );
not \U$215 ( \295 , \294 );
nand \U$216 ( \296 , RIa139b90_40, \170_nG5b );
nor \U$217 ( \297 , \278 , \296 );
not \U$218 ( \298 , \297 );
not \U$219 ( \299 , \282 );
not \U$220 ( \300 , \299 );
or \U$221 ( \301 , \298 , \300 );
and \U$222 ( \302 , \282 , \283 );
nor \U$223 ( \303 , \302 , \290 );
nand \U$224 ( \304 , \301 , \303 );
not \U$225 ( \305 , \304 );
or \U$226 ( \306 , \295 , \305 );
nand \U$227 ( \307 , RIa139b18_39, \162_nG6b );
nand \U$228 ( \308 , RIa139b90_40, \188_nG73 );
xor \U$229 ( \309 , \307 , \308 );
not \U$230 ( \310 , \309 );
not \U$231 ( \311 , \180 );
nand \U$232 ( \312 , \311 , RIa139b90_40, RIa139b18_39);
not \U$233 ( \313 , \312 );
not \U$234 ( \314 , \313 );
and \U$235 ( \315 , \310 , \314 );
and \U$236 ( \316 , \309 , \313 );
nor \U$237 ( \317 , \315 , \316 );
buf \U$238 ( \318 , \317 );
nand \U$239 ( \319 , \306 , \318 );
nand \U$240 ( \320 , \293 , \319 );
not \U$241 ( \321 , \320 );
or \U$242 ( \322 , \274 , \321 );
not \U$243 ( \323 , \270 );
and \U$244 ( \324 , \204 , \196 );
not \U$245 ( \325 , \204 );
and \U$246 ( \326 , \325 , \195 );
nor \U$247 ( \327 , \324 , \326 );
nand \U$248 ( \328 , \323 , \327 );
nand \U$249 ( \329 , \322 , \328 );
nand \U$250 ( \330 , \269 , \329 );
nand \U$251 ( \331 , \266 , \330 );
not \U$252 ( \332 , \331 );
or \U$253 ( \333 , \261 , \332 );
not \U$254 ( \334 , \258 );
xor \U$255 ( \335 , \213 , \217 );
nand \U$256 ( \336 , \334 , \335 );
nand \U$257 ( \337 , \333 , \336 );
not \U$258 ( \338 , \337 );
or \U$259 ( \339 , \257 , \338 );
not \U$260 ( \340 , \254 );
xor \U$261 ( \341 , \221 , \133 );
nand \U$262 ( \342 , \340 , \341 );
nand \U$263 ( \343 , \339 , \342 );
not \U$264 ( \344 , \343 );
or \U$265 ( \345 , \253 , \344 );
not \U$266 ( \346 , \250 );
xor \U$267 ( \347 , \225 , \121 );
nand \U$268 ( \348 , \346 , \347 );
nand \U$269 ( \349 , \345 , \348 );
not \U$270 ( \350 , \349 );
or \U$271 ( \351 , \249 , \350 );
not \U$272 ( \352 , \246 );
xor \U$273 ( \353 , \229 , \117 );
nand \U$274 ( \354 , \352 , \353 );
nand \U$275 ( \355 , \351 , \354 );
not \U$276 ( \356 , \355 );
or \U$277 ( \357 , \245 , \356 );
not \U$278 ( \358 , \242 );
xor \U$279 ( \359 , \233 , \234 );
nand \U$280 ( \360 , \358 , \359 );
nand \U$281 ( \361 , \357 , \360 );
not \U$282 ( \362 , \361 );
or \U$283 ( \363 , \241 , \362 );
not \U$284 ( \364 , \114 );
nand \U$285 ( \365 , \364 , \236 );
nand \U$286 ( \366 , \363 , \365 );
nand \U$287 ( \367 , RIa139a28_37, \109_nGa3 );
xnor \U$288 ( \368 , \366 , \367 );
not \U$289 ( \369 , \368 );
nand \U$290 ( \370 , RIa139a28_37, \100_nG9b );
xor \U$291 ( \371 , \370 , \240 );
xnor \U$292 ( \372 , \371 , \361 );
not \U$293 ( \373 , \372 );
nand \U$294 ( \374 , RIa139a28_37, \91_nG93 );
xor \U$295 ( \375 , \374 , \244 );
xnor \U$296 ( \376 , \375 , \355 );
not \U$297 ( \377 , \376 );
nand \U$298 ( \378 , RIa139a28_37, \131_nG8b );
xor \U$299 ( \379 , \378 , \248 );
not \U$300 ( \380 , \349 );
xnor \U$301 ( \381 , \379 , \380 );
not \U$302 ( \382 , \381 );
not \U$303 ( \383 , \382 );
nand \U$304 ( \384 , RIa139a28_37, \142_nG83 );
xor \U$305 ( \385 , \384 , \252 );
xnor \U$306 ( \386 , \385 , \343 );
not \U$307 ( \387 , \386 );
nand \U$308 ( \388 , RIa139a28_37, \151_nG7b );
not \U$309 ( \389 , \256 );
xor \U$310 ( \390 , \388 , \389 );
xor \U$311 ( \391 , \390 , \337 );
not \U$312 ( \392 , \391 );
not \U$313 ( \393 , \320 );
not \U$314 ( \394 , \272 );
and \U$315 ( \395 , \393 , \394 );
and \U$316 ( \396 , \320 , \272 );
nor \U$317 ( \397 , \395 , \396 );
not \U$318 ( \398 , \397 );
nand \U$319 ( \399 , RIa139a28_37, \179_nG63 );
not \U$320 ( \400 , \399 );
and \U$321 ( \401 , \398 , \400 );
and \U$322 ( \402 , \397 , \399 );
buf \U$323 ( \403 , \304 );
not \U$324 ( \404 , \294 );
not \U$325 ( \405 , \317 );
or \U$326 ( \406 , \404 , \405 );
or \U$327 ( \407 , \294 , \317 );
nand \U$328 ( \408 , \406 , \407 );
xnor \U$329 ( \409 , \403 , \408 );
nand \U$330 ( \410 , RIa139a28_37, \170_nG5b );
not \U$331 ( \411 , \410 );
nand \U$332 ( \412 , \409 , \411 );
nor \U$333 ( \413 , \402 , \412 );
nor \U$334 ( \414 , \401 , \413 );
not \U$335 ( \415 , \414 );
nand \U$336 ( \416 , RIa139a28_37, \162_nG6b );
xor \U$337 ( \417 , \416 , \268 );
not \U$338 ( \418 , \329 );
xnor \U$339 ( \419 , \417 , \418 );
nand \U$340 ( \420 , \415 , \419 );
not \U$341 ( \421 , \416 );
xor \U$342 ( \422 , \418 , \268 );
nand \U$343 ( \423 , \421 , \422 );
nand \U$344 ( \424 , \420 , \423 );
not \U$345 ( \425 , \424 );
nand \U$346 ( \426 , RIa139a28_37, \188_nG73 );
xor \U$347 ( \427 , \426 , \260 );
xnor \U$348 ( \428 , \427 , \331 );
not \U$349 ( \429 , \428 );
or \U$350 ( \430 , \425 , \429 );
not \U$351 ( \431 , \426 );
xor \U$352 ( \432 , \331 , \260 );
nand \U$353 ( \433 , \431 , \432 );
nand \U$354 ( \434 , \430 , \433 );
not \U$355 ( \435 , \434 );
or \U$356 ( \436 , \392 , \435 );
not \U$357 ( \437 , \388 );
and \U$358 ( \438 , \337 , \256 );
not \U$359 ( \439 , \337 );
and \U$360 ( \440 , \439 , \389 );
nor \U$361 ( \441 , \438 , \440 );
nand \U$362 ( \442 , \437 , \441 );
nand \U$363 ( \443 , \436 , \442 );
not \U$364 ( \444 , \443 );
or \U$365 ( \445 , \387 , \444 );
not \U$366 ( \446 , \384 );
xor \U$367 ( \447 , \343 , \252 );
nand \U$368 ( \448 , \446 , \447 );
nand \U$369 ( \449 , \445 , \448 );
not \U$370 ( \450 , \449 );
or \U$371 ( \451 , \383 , \450 );
not \U$372 ( \452 , \378 );
not \U$373 ( \453 , \248 );
not \U$374 ( \454 , \380 );
or \U$375 ( \455 , \453 , \454 );
or \U$376 ( \456 , \380 , \248 );
nand \U$377 ( \457 , \455 , \456 );
nand \U$378 ( \458 , \452 , \457 );
nand \U$379 ( \459 , \451 , \458 );
not \U$380 ( \460 , \459 );
or \U$381 ( \461 , \377 , \460 );
not \U$382 ( \462 , \374 );
xor \U$383 ( \463 , \355 , \244 );
nand \U$384 ( \464 , \462 , \463 );
nand \U$385 ( \465 , \461 , \464 );
not \U$386 ( \466 , \465 );
or \U$387 ( \467 , \373 , \466 );
not \U$388 ( \468 , \370 );
not \U$389 ( \469 , \240 );
not \U$390 ( \470 , \361 );
not \U$391 ( \471 , \470 );
or \U$392 ( \472 , \469 , \471 );
or \U$393 ( \473 , \470 , \240 );
nand \U$394 ( \474 , \472 , \473 );
nand \U$395 ( \475 , \468 , \474 );
nand \U$396 ( \476 , \467 , \475 );
not \U$397 ( \477 , \476 );
or \U$398 ( \478 , \369 , \477 );
not \U$399 ( \479 , \367 );
nand \U$400 ( \480 , \479 , \366 );
nand \U$401 ( \481 , \478 , \480 );
xnor \U$402 ( \482 , \113 , \481 );
not \U$403 ( \483 , \482 );
not \U$404 ( \484 , \483 );
nand \U$405 ( \485 , RIa1399b0_36, \100_nG9b );
xor \U$406 ( \486 , \485 , \368 );
xnor \U$407 ( \487 , \486 , \476 );
not \U$408 ( \488 , \487 );
nand \U$409 ( \489 , RIa1399b0_36, \91_nG93 );
xor \U$410 ( \490 , \489 , \372 );
xnor \U$411 ( \491 , \490 , \465 );
not \U$412 ( \492 , \491 );
nand \U$413 ( \493 , RIa1399b0_36, \142_nG83 );
xor \U$414 ( \494 , \493 , \381 );
xnor \U$415 ( \495 , \494 , \449 );
not \U$416 ( \496 , \495 );
not \U$417 ( \497 , \496 );
nand \U$418 ( \498 , RIa1399b0_36, \151_nG7b );
xor \U$419 ( \499 , \498 , \386 );
xnor \U$420 ( \500 , \499 , \443 );
not \U$421 ( \501 , \500 );
nand \U$422 ( \502 , RIa1399b0_36, \188_nG73 );
xor \U$423 ( \503 , \502 , \391 );
xnor \U$424 ( \504 , \503 , \434 );
not \U$425 ( \505 , \504 );
nand \U$426 ( \506 , RIa1399b0_36, \162_nG6b );
xor \U$427 ( \507 , \506 , \424 );
xnor \U$428 ( \508 , \507 , \428 );
not \U$429 ( \509 , \508 );
xor \U$430 ( \510 , \399 , \412 );
xnor \U$431 ( \511 , \510 , \397 );
nand \U$432 ( \512 , RIa1399b0_36, \170_nG5b );
not \U$433 ( \513 , \512 );
and \U$434 ( \514 , \511 , \513 );
not \U$435 ( \515 , \179_nG63 );
nor \U$436 ( \516 , \112 , \515 );
xor \U$437 ( \517 , \514 , \516 );
and \U$438 ( \518 , \419 , \415 );
not \U$439 ( \519 , \419 );
and \U$440 ( \520 , \519 , \414 );
nor \U$441 ( \521 , \518 , \520 );
and \U$442 ( \522 , \517 , \521 );
and \U$443 ( \523 , \514 , \516 );
or \U$444 ( \524 , \522 , \523 );
not \U$445 ( \525 , \524 );
or \U$446 ( \526 , \509 , \525 );
not \U$447 ( \527 , \506 );
xor \U$448 ( \528 , \428 , \424 );
nand \U$449 ( \529 , \527 , \528 );
nand \U$450 ( \530 , \526 , \529 );
not \U$451 ( \531 , \530 );
or \U$452 ( \532 , \505 , \531 );
not \U$453 ( \533 , \502 );
xor \U$454 ( \534 , \434 , \391 );
nand \U$455 ( \535 , \533 , \534 );
nand \U$456 ( \536 , \532 , \535 );
not \U$457 ( \537 , \536 );
or \U$458 ( \538 , \501 , \537 );
not \U$459 ( \539 , \498 );
xor \U$460 ( \540 , \386 , \443 );
nand \U$461 ( \541 , \539 , \540 );
nand \U$462 ( \542 , \538 , \541 );
not \U$463 ( \543 , \542 );
or \U$464 ( \544 , \497 , \543 );
not \U$465 ( \545 , \493 );
and \U$466 ( \546 , \449 , \381 );
not \U$467 ( \547 , \449 );
and \U$468 ( \548 , \547 , \382 );
or \U$469 ( \549 , \546 , \548 );
nand \U$470 ( \550 , \545 , \549 );
nand \U$471 ( \551 , \544 , \550 );
not \U$472 ( \552 , \551 );
nand \U$473 ( \553 , RIa1399b0_36, \131_nG8b );
xor \U$474 ( \554 , \553 , \376 );
xnor \U$475 ( \555 , \554 , \459 );
not \U$476 ( \556 , \555 );
or \U$477 ( \557 , \552 , \556 );
not \U$478 ( \558 , \553 );
xor \U$479 ( \559 , \376 , \459 );
nand \U$480 ( \560 , \558 , \559 );
nand \U$481 ( \561 , \557 , \560 );
not \U$482 ( \562 , \561 );
or \U$483 ( \563 , \492 , \562 );
not \U$484 ( \564 , \489 );
xor \U$485 ( \565 , \465 , \372 );
nand \U$486 ( \566 , \564 , \565 );
nand \U$487 ( \567 , \563 , \566 );
not \U$488 ( \568 , \567 );
or \U$489 ( \569 , \488 , \568 );
not \U$490 ( \570 , \485 );
xor \U$491 ( \571 , \476 , \368 );
nand \U$492 ( \572 , \570 , \571 );
nand \U$493 ( \573 , \569 , \572 );
not \U$494 ( \574 , \573 );
or \U$495 ( \575 , \484 , \574 );
nand \U$496 ( \576 , \481 , \113 );
nand \U$497 ( \577 , \575 , \576 );
xnor \U$498 ( \578 , \110 , \577 );
xor \U$499 ( \579 , \101 , \578 );
nand \U$500 ( \580 , RIa139938_35, \100_nG9b );
xor \U$501 ( \581 , \580 , \482 );
xnor \U$502 ( \582 , \581 , \573 );
not \U$503 ( \583 , \582 );
not \U$504 ( \584 , \583 );
nand \U$505 ( \585 , RIa139938_35, \91_nG93 );
xor \U$506 ( \586 , \585 , \487 );
xnor \U$507 ( \587 , \586 , \567 );
not \U$508 ( \588 , \587 );
nand \U$509 ( \589 , RIa139938_35, \131_nG8b );
xor \U$510 ( \590 , \589 , \491 );
not \U$511 ( \591 , \561 );
xnor \U$512 ( \592 , \590 , \591 );
not \U$513 ( \593 , \592 );
not \U$514 ( \594 , \593 );
nand \U$515 ( \595 , RIa139938_35, \142_nG83 );
xor \U$516 ( \596 , \595 , \555 );
not \U$517 ( \597 , \551 );
xnor \U$518 ( \598 , \596 , \597 );
not \U$519 ( \599 , \598 );
not \U$520 ( \600 , \599 );
nand \U$521 ( \601 , RIa139938_35, \151_nG7b );
not \U$522 ( \602 , \601 );
not \U$523 ( \603 , \496 );
not \U$524 ( \604 , \542 );
not \U$525 ( \605 , \604 );
or \U$526 ( \606 , \603 , \605 );
nand \U$527 ( \607 , \542 , \495 );
nand \U$528 ( \608 , \606 , \607 );
not \U$529 ( \609 , \608 );
or \U$530 ( \610 , \602 , \609 );
or \U$531 ( \611 , \601 , \608 );
nand \U$532 ( \612 , \610 , \611 );
not \U$533 ( \613 , \612 );
and \U$534 ( \614 , RIa139938_35, \179_nG63 );
and \U$535 ( \615 , RIa139938_35, \170_nG5b );
xor \U$536 ( \616 , \514 , \516 );
xor \U$537 ( \617 , \616 , \521 );
and \U$538 ( \618 , \615 , \617 );
xor \U$539 ( \619 , \614 , \618 );
xor \U$540 ( \620 , \508 , \524 );
and \U$541 ( \621 , \619 , \620 );
and \U$542 ( \622 , \614 , \618 );
or \U$543 ( \623 , \621 , \622 );
not \U$544 ( \624 , \623 );
nand \U$545 ( \625 , RIa139938_35, \162_nG6b );
xor \U$546 ( \626 , \625 , \530 );
not \U$547 ( \627 , \504 );
xor \U$548 ( \628 , \626 , \627 );
not \U$549 ( \629 , \628 );
or \U$550 ( \630 , \624 , \629 );
not \U$551 ( \631 , \625 );
and \U$552 ( \632 , \530 , \627 );
not \U$553 ( \633 , \530 );
and \U$554 ( \634 , \633 , \504 );
or \U$555 ( \635 , \632 , \634 );
nand \U$556 ( \636 , \631 , \635 );
nand \U$557 ( \637 , \630 , \636 );
not \U$558 ( \638 , \637 );
nand \U$559 ( \639 , RIa139938_35, \188_nG73 );
not \U$560 ( \640 , \500 );
xor \U$561 ( \641 , \639 , \640 );
not \U$562 ( \642 , \536 );
xnor \U$563 ( \643 , \641 , \642 );
not \U$564 ( \644 , \643 );
or \U$565 ( \645 , \638 , \644 );
not \U$566 ( \646 , \639 );
and \U$567 ( \647 , \642 , \500 );
not \U$568 ( \648 , \642 );
and \U$569 ( \649 , \648 , \640 );
or \U$570 ( \650 , \647 , \649 );
nand \U$571 ( \651 , \646 , \650 );
nand \U$572 ( \652 , \645 , \651 );
not \U$573 ( \653 , \652 );
or \U$574 ( \654 , \613 , \653 );
not \U$575 ( \655 , \601 );
nand \U$576 ( \656 , \655 , \608 );
nand \U$577 ( \657 , \654 , \656 );
not \U$578 ( \658 , \657 );
or \U$579 ( \659 , \600 , \658 );
not \U$580 ( \660 , \595 );
and \U$581 ( \661 , \555 , \597 );
not \U$582 ( \662 , \555 );
and \U$583 ( \663 , \662 , \551 );
or \U$584 ( \664 , \661 , \663 );
nand \U$585 ( \665 , \660 , \664 );
nand \U$586 ( \666 , \659 , \665 );
not \U$587 ( \667 , \666 );
or \U$588 ( \668 , \594 , \667 );
not \U$589 ( \669 , \589 );
and \U$590 ( \670 , \491 , \591 );
not \U$591 ( \671 , \491 );
and \U$592 ( \672 , \671 , \561 );
or \U$593 ( \673 , \670 , \672 );
nand \U$594 ( \674 , \669 , \673 );
nand \U$595 ( \675 , \668 , \674 );
not \U$596 ( \676 , \675 );
or \U$597 ( \677 , \588 , \676 );
not \U$598 ( \678 , \487 );
and \U$599 ( \679 , \567 , \678 );
nor \U$600 ( \680 , \567 , \678 );
or \U$601 ( \681 , \679 , \680 );
not \U$602 ( \682 , \585 );
nand \U$603 ( \683 , \681 , \682 );
nand \U$604 ( \684 , \677 , \683 );
not \U$605 ( \685 , \684 );
or \U$606 ( \686 , \584 , \685 );
not \U$607 ( \687 , \580 );
xnor \U$608 ( \688 , \573 , \482 );
nand \U$609 ( \689 , \687 , \688 );
nand \U$610 ( \690 , \686 , \689 );
xnor \U$611 ( \691 , \579 , \690 );
xor \U$612 ( \692 , \92 , \691 );
nand \U$613 ( \693 , RIa1398c0_34, \91_nG93 );
xor \U$614 ( \694 , \693 , \582 );
xnor \U$615 ( \695 , \694 , \684 );
not \U$616 ( \696 , \695 );
not \U$617 ( \697 , \696 );
nand \U$618 ( \698 , RIa1398c0_34, \131_nG8b );
xor \U$619 ( \699 , \698 , \587 );
xnor \U$620 ( \700 , \699 , \675 );
not \U$621 ( \701 , \700 );
nand \U$622 ( \702 , RIa1398c0_34, \142_nG83 );
not \U$623 ( \703 , \702 );
not \U$624 ( \704 , \593 );
not \U$625 ( \705 , \666 );
not \U$626 ( \706 , \705 );
or \U$627 ( \707 , \704 , \706 );
nand \U$628 ( \708 , \666 , \592 );
nand \U$629 ( \709 , \707 , \708 );
not \U$630 ( \710 , \709 );
or \U$631 ( \711 , \703 , \710 );
or \U$632 ( \712 , \702 , \709 );
nand \U$633 ( \713 , \711 , \712 );
not \U$634 ( \714 , \713 );
not \U$635 ( \715 , RIa1398c0_34);
nor \U$636 ( \716 , \515 , \715 );
xor \U$637 ( \717 , \614 , \618 );
xor \U$638 ( \718 , \717 , \620 );
not \U$639 ( \719 , \718 );
nand \U$640 ( \720 , RIa1398c0_34, \170_nG5b );
nor \U$641 ( \721 , \719 , \720 );
xor \U$642 ( \722 , \716 , \721 );
xor \U$643 ( \723 , \628 , \623 );
and \U$644 ( \724 , \722 , \723 );
and \U$645 ( \725 , \716 , \721 );
or \U$646 ( \726 , \724 , \725 );
not \U$647 ( \727 , \726 );
nand \U$648 ( \728 , RIa1398c0_34, \162_nG6b );
not \U$649 ( \729 , \637 );
xor \U$650 ( \730 , \728 , \729 );
not \U$651 ( \731 , \643 );
xnor \U$652 ( \732 , \730 , \731 );
not \U$653 ( \733 , \732 );
or \U$654 ( \734 , \727 , \733 );
nand \U$655 ( \735 , \643 , \729 );
not \U$656 ( \736 , \735 );
nand \U$657 ( \737 , \731 , \637 );
not \U$658 ( \738 , \737 );
or \U$659 ( \739 , \736 , \738 );
not \U$660 ( \740 , \728 );
nand \U$661 ( \741 , \739 , \740 );
nand \U$662 ( \742 , \734 , \741 );
not \U$663 ( \743 , \742 );
nor \U$664 ( \744 , \192 , \715 );
not \U$665 ( \745 , \744 );
not \U$666 ( \746 , \652 );
not \U$667 ( \747 , \746 );
not \U$668 ( \748 , \612 );
or \U$669 ( \749 , \747 , \748 );
not \U$670 ( \750 , \612 );
nand \U$671 ( \751 , \750 , \652 );
nand \U$672 ( \752 , \749 , \751 );
not \U$673 ( \753 , \752 );
not \U$674 ( \754 , \753 );
or \U$675 ( \755 , \745 , \754 );
not \U$676 ( \756 , \744 );
nand \U$677 ( \757 , \752 , \756 );
nand \U$678 ( \758 , \755 , \757 );
not \U$679 ( \759 , \758 );
or \U$680 ( \760 , \743 , \759 );
nand \U$681 ( \761 , \752 , \744 );
nand \U$682 ( \762 , \760 , \761 );
not \U$683 ( \763 , \762 );
not \U$684 ( \764 , \151_nG7b );
nor \U$685 ( \765 , \715 , \764 );
not \U$686 ( \766 , \765 );
not \U$687 ( \767 , \599 );
not \U$688 ( \768 , \657 );
not \U$689 ( \769 , \768 );
or \U$690 ( \770 , \767 , \769 );
nand \U$691 ( \771 , \657 , \598 );
nand \U$692 ( \772 , \770 , \771 );
not \U$693 ( \773 , \772 );
not \U$694 ( \774 , \773 );
or \U$695 ( \775 , \766 , \774 );
not \U$696 ( \776 , RIa1398c0_34);
not \U$697 ( \777 , \151_nG7b );
or \U$698 ( \778 , \776 , \777 );
nand \U$699 ( \779 , \778 , \772 );
nand \U$700 ( \780 , \775 , \779 );
not \U$701 ( \781 , \780 );
or \U$702 ( \782 , \763 , \781 );
nand \U$703 ( \783 , \772 , \765 );
nand \U$704 ( \784 , \782 , \783 );
not \U$705 ( \785 , \784 );
or \U$706 ( \786 , \714 , \785 );
not \U$707 ( \787 , \702 );
not \U$708 ( \788 , \593 );
not \U$709 ( \789 , \705 );
or \U$710 ( \790 , \788 , \789 );
nand \U$711 ( \791 , \790 , \708 );
nand \U$712 ( \792 , \787 , \791 );
nand \U$713 ( \793 , \786 , \792 );
not \U$714 ( \794 , \793 );
or \U$715 ( \795 , \701 , \794 );
not \U$716 ( \796 , \698 );
xor \U$717 ( \797 , \587 , \675 );
nand \U$718 ( \798 , \796 , \797 );
nand \U$719 ( \799 , \795 , \798 );
not \U$720 ( \800 , \799 );
or \U$721 ( \801 , \697 , \800 );
not \U$722 ( \802 , \583 );
nand \U$723 ( \803 , \802 , \684 );
not \U$724 ( \804 , \803 );
not \U$725 ( \805 , \684 );
nand \U$726 ( \806 , \805 , \583 );
not \U$727 ( \807 , \806 );
or \U$728 ( \808 , \804 , \807 );
not \U$729 ( \809 , \693 );
nand \U$730 ( \810 , \808 , \809 );
nand \U$731 ( \811 , \801 , \810 );
xnor \U$732 ( \812 , \692 , \811 );
not \U$733 ( \813 , \812 );
nand \U$734 ( \814 , RIa139848_33, \142_nG83 );
not \U$735 ( \815 , \700 );
xor \U$736 ( \816 , \814 , \815 );
buf \U$737 ( \817 , \793 );
not \U$738 ( \818 , \817 );
xnor \U$739 ( \819 , \816 , \818 );
not \U$740 ( \820 , \819 );
nand \U$741 ( \821 , RIa139848_33, \162_nG6b );
xor \U$742 ( \822 , \821 , \742 );
xnor \U$743 ( \823 , \822 , \758 );
not \U$744 ( \824 , \823 );
nand \U$745 ( \825 , RIa139848_33, \179_nG63 );
not \U$746 ( \826 , \825 );
xnor \U$747 ( \827 , \732 , \726 );
not \U$748 ( \828 , \827 );
or \U$749 ( \829 , \826 , \828 );
xor \U$750 ( \830 , \716 , \721 );
xor \U$751 ( \831 , \830 , \723 );
nand \U$752 ( \832 , RIa139848_33, \170_nG5b );
not \U$753 ( \833 , \832 );
and \U$754 ( \834 , \831 , \833 );
nand \U$755 ( \835 , \829 , \834 );
or \U$756 ( \836 , \825 , \827 );
nand \U$757 ( \837 , \835 , \836 );
not \U$758 ( \838 , \837 );
or \U$759 ( \839 , \824 , \838 );
not \U$760 ( \840 , \758 );
nand \U$761 ( \841 , \840 , \742 );
not \U$762 ( \842 , \841 );
not \U$763 ( \843 , \742 );
nand \U$764 ( \844 , \843 , \758 );
not \U$765 ( \845 , \844 );
or \U$766 ( \846 , \842 , \845 );
not \U$767 ( \847 , \821 );
nand \U$768 ( \848 , \846 , \847 );
nand \U$769 ( \849 , \839 , \848 );
not \U$770 ( \850 , \849 );
nand \U$771 ( \851 , RIa139848_33, \188_nG73 );
xor \U$772 ( \852 , \851 , \780 );
xnor \U$773 ( \853 , \852 , \762 );
not \U$774 ( \854 , \853 );
or \U$775 ( \855 , \850 , \854 );
not \U$776 ( \856 , \851 );
not \U$777 ( \857 , \765 );
not \U$778 ( \858 , \773 );
or \U$779 ( \859 , \857 , \858 );
nand \U$780 ( \860 , \859 , \779 );
xor \U$781 ( \861 , \860 , \762 );
nand \U$782 ( \862 , \856 , \861 );
nand \U$783 ( \863 , \855 , \862 );
not \U$784 ( \864 , \863 );
not \U$785 ( \865 , RIa139848_33);
nor \U$786 ( \866 , \865 , \764 );
not \U$787 ( \867 , \866 );
not \U$788 ( \868 , \713 );
not \U$789 ( \869 , \784 );
not \U$790 ( \870 , \869 );
or \U$791 ( \871 , \868 , \870 );
not \U$792 ( \872 , \713 );
nand \U$793 ( \873 , \872 , \784 );
nand \U$794 ( \874 , \871 , \873 );
not \U$795 ( \875 , \874 );
not \U$796 ( \876 , \875 );
or \U$797 ( \877 , \867 , \876 );
not \U$798 ( \878 , \866 );
nand \U$799 ( \879 , \878 , \874 );
nand \U$800 ( \880 , \877 , \879 );
not \U$801 ( \881 , \880 );
or \U$802 ( \882 , \864 , \881 );
nand \U$803 ( \883 , \874 , \866 );
nand \U$804 ( \884 , \882 , \883 );
not \U$805 ( \885 , \884 );
or \U$806 ( \886 , \820 , \885 );
not \U$807 ( \887 , \814 );
not \U$808 ( \888 , \815 );
not \U$809 ( \889 , \817 );
or \U$810 ( \890 , \888 , \889 );
nand \U$811 ( \891 , \818 , \700 );
nand \U$812 ( \892 , \890 , \891 );
nand \U$813 ( \893 , \887 , \892 );
nand \U$814 ( \894 , \886 , \893 );
not \U$815 ( \895 , \894 );
not \U$816 ( \896 , \695 );
not \U$817 ( \897 , \799 );
or \U$818 ( \898 , \896 , \897 );
or \U$819 ( \899 , \695 , \799 );
nand \U$820 ( \900 , \898 , \899 );
not \U$821 ( \901 , \900 );
nand \U$822 ( \902 , RIa139848_33, \131_nG8b );
not \U$823 ( \903 , \902 );
and \U$824 ( \904 , \901 , \903 );
and \U$825 ( \905 , \900 , \902 );
nor \U$826 ( \906 , \904 , \905 );
not \U$827 ( \907 , \906 );
not \U$828 ( \908 , \907 );
or \U$829 ( \909 , \895 , \908 );
not \U$830 ( \910 , \902 );
nand \U$831 ( \911 , \910 , \900 );
nand \U$832 ( \912 , \909 , \911 );
not \U$833 ( \913 , \912 );
or \U$834 ( \914 , \813 , \913 );
not \U$835 ( \915 , \92 );
not \U$836 ( \916 , \691 );
not \U$837 ( \917 , \916 );
not \U$838 ( \918 , \811 );
or \U$839 ( \919 , \917 , \918 );
or \U$840 ( \920 , \811 , \916 );
nand \U$841 ( \921 , \919 , \920 );
nand \U$842 ( \922 , \915 , \921 );
nand \U$843 ( \923 , \914 , \922 );
not \U$844 ( \924 , \923 );
nand \U$845 ( \925 , RIa139848_33, \100_nG9b );
not \U$846 ( \926 , \578 );
not \U$847 ( \927 , \690 );
or \U$848 ( \928 , \926 , \927 );
not \U$849 ( \929 , \110 );
nand \U$850 ( \930 , \929 , \577 );
nand \U$851 ( \931 , \928 , \930 );
nand \U$852 ( \932 , RIa1398c0_34, \109_nGa3 );
xnor \U$853 ( \933 , \931 , \932 );
xor \U$854 ( \934 , \925 , \933 );
not \U$855 ( \935 , \691 );
not \U$856 ( \936 , \811 );
or \U$857 ( \937 , \935 , \936 );
not \U$858 ( \938 , \101 );
xor \U$859 ( \939 , \690 , \578 );
nand \U$860 ( \940 , \938 , \939 );
nand \U$861 ( \941 , \937 , \940 );
xnor \U$862 ( \942 , \934 , \941 );
not \U$863 ( \943 , \942 );
or \U$864 ( \944 , \924 , \943 );
not \U$865 ( \945 , \925 );
xor \U$866 ( \946 , \941 , \933 );
nand \U$867 ( \947 , \945 , \946 );
nand \U$868 ( \948 , \944 , \947 );
not \U$869 ( \949 , \948 );
not \U$870 ( \950 , \933 );
not \U$871 ( \951 , \941 );
or \U$872 ( \952 , \950 , \951 );
not \U$873 ( \953 , \932 );
nand \U$874 ( \954 , \953 , \931 );
nand \U$875 ( \955 , \952 , \954 );
nand \U$876 ( \956 , RIa139848_33, \109_nGa3 );
xnor \U$877 ( \957 , \955 , \956 );
not \U$878 ( \958 , \957 );
or \U$879 ( \959 , \949 , \958 );
not \U$880 ( \960 , \956 );
nand \U$881 ( \961 , \960 , \955 );
nand \U$882 ( \962 , \959 , \961 );
nand \U$883 ( \963 , RIa1397d0_32, \109_nGa3 );
and \U$884 ( \964 , \962 , \963 );
not \U$885 ( \965 , \962 );
not \U$886 ( \966 , \963 );
and \U$887 ( \967 , \965 , \966 );
or \U$888 ( \968 , \964 , \967 );
not \U$889 ( \969 , \968 );
nand \U$890 ( \970 , RIa1397d0_32, \100_nG9b );
xor \U$891 ( \971 , \970 , \957 );
xnor \U$892 ( \972 , \971 , \948 );
not \U$893 ( \973 , \972 );
nand \U$894 ( \974 , RIa1397d0_32, \91_nG93 );
not \U$895 ( \975 , \942 );
xor \U$896 ( \976 , \974 , \975 );
xor \U$897 ( \977 , \976 , \923 );
not \U$898 ( \978 , \977 );
xor \U$899 ( \979 , \825 , \834 );
xnor \U$900 ( \980 , \979 , \827 );
nand \U$901 ( \981 , RIa1397d0_32, \170_nG5b );
nor \U$902 ( \982 , \980 , \981 );
and \U$903 ( \983 , RIa1397d0_32, \179_nG63 );
xor \U$904 ( \984 , \982 , \983 );
xor \U$905 ( \985 , \823 , \837 );
and \U$906 ( \986 , \984 , \985 );
and \U$907 ( \987 , \982 , \983 );
or \U$908 ( \988 , \986 , \987 );
not \U$909 ( \989 , \988 );
nand \U$910 ( \990 , RIa1397d0_32, \162_nG6b );
xor \U$911 ( \991 , \990 , \849 );
xnor \U$912 ( \992 , \991 , \853 );
not \U$913 ( \993 , \992 );
or \U$914 ( \994 , \989 , \993 );
not \U$915 ( \995 , \853 );
nand \U$916 ( \996 , \995 , \849 );
not \U$917 ( \997 , \996 );
not \U$918 ( \998 , \849 );
nand \U$919 ( \999 , \998 , \853 );
not \U$920 ( \1000 , \999 );
or \U$921 ( \1001 , \997 , \1000 );
not \U$922 ( \1002 , \990 );
nand \U$923 ( \1003 , \1001 , \1002 );
nand \U$924 ( \1004 , \994 , \1003 );
not \U$925 ( \1005 , \1004 );
nand \U$926 ( \1006 , RIa1397d0_32, \188_nG73 );
not \U$927 ( \1007 , \880 );
xor \U$928 ( \1008 , \1006 , \1007 );
not \U$929 ( \1009 , \863 );
xnor \U$930 ( \1010 , \1008 , \1009 );
not \U$931 ( \1011 , \1010 );
or \U$932 ( \1012 , \1005 , \1011 );
not \U$933 ( \1013 , \1009 );
nand \U$934 ( \1014 , \1013 , \1007 );
not \U$935 ( \1015 , \1014 );
not \U$936 ( \1016 , \1007 );
nand \U$937 ( \1017 , \1016 , \1009 );
not \U$938 ( \1018 , \1017 );
or \U$939 ( \1019 , \1015 , \1018 );
not \U$940 ( \1020 , \1006 );
nand \U$941 ( \1021 , \1019 , \1020 );
nand \U$942 ( \1022 , \1012 , \1021 );
not \U$943 ( \1023 , \1022 );
not \U$944 ( \1024 , RIa1397d0_32);
nor \U$945 ( \1025 , \1024 , \764 );
not \U$946 ( \1026 , \1025 );
xor \U$947 ( \1027 , \819 , \884 );
not \U$948 ( \1028 , \1027 );
not \U$949 ( \1029 , \1028 );
or \U$950 ( \1030 , \1026 , \1029 );
not \U$951 ( \1031 , \1025 );
nand \U$952 ( \1032 , \1031 , \1027 );
nand \U$953 ( \1033 , \1030 , \1032 );
not \U$954 ( \1034 , \1033 );
or \U$955 ( \1035 , \1023 , \1034 );
nand \U$956 ( \1036 , \1027 , \1025 );
nand \U$957 ( \1037 , \1035 , \1036 );
not \U$958 ( \1038 , \1037 );
not \U$959 ( \1039 , \906 );
not \U$960 ( \1040 , \894 );
or \U$961 ( \1041 , \1039 , \1040 );
or \U$962 ( \1042 , \906 , \894 );
nand \U$963 ( \1043 , \1041 , \1042 );
not \U$964 ( \1044 , \1043 );
nand \U$965 ( \1045 , RIa1397d0_32, \142_nG83 );
not \U$966 ( \1046 , \1045 );
and \U$967 ( \1047 , \1044 , \1046 );
and \U$968 ( \1048 , \1043 , \1045 );
nor \U$969 ( \1049 , \1047 , \1048 );
not \U$970 ( \1050 , \1049 );
not \U$971 ( \1051 , \1050 );
or \U$972 ( \1052 , \1038 , \1051 );
not \U$973 ( \1053 , \1045 );
nand \U$974 ( \1054 , \1053 , \1043 );
nand \U$975 ( \1055 , \1052 , \1054 );
nand \U$976 ( \1056 , RIa1397d0_32, \131_nG8b );
xor \U$977 ( \1057 , \1056 , \812 );
xnor \U$978 ( \1058 , \1057 , \912 );
nand \U$979 ( \1059 , \1055 , \1058 );
not \U$980 ( \1060 , \1056 );
xor \U$981 ( \1061 , \912 , \812 );
nand \U$982 ( \1062 , \1060 , \1061 );
nand \U$983 ( \1063 , \1059 , \1062 );
not \U$984 ( \1064 , \1063 );
or \U$985 ( \1065 , \978 , \1064 );
not \U$986 ( \1066 , \974 );
xnor \U$987 ( \1067 , \923 , \975 );
nand \U$988 ( \1068 , \1066 , \1067 );
nand \U$989 ( \1069 , \1065 , \1068 );
not \U$990 ( \1070 , \1069 );
or \U$991 ( \1071 , \973 , \1070 );
not \U$992 ( \1072 , \970 );
xor \U$993 ( \1073 , \948 , \957 );
nand \U$994 ( \1074 , \1072 , \1073 );
nand \U$995 ( \1075 , \1071 , \1074 );
not \U$996 ( \1076 , \1075 );
or \U$997 ( \1077 , \969 , \1076 );
nand \U$998 ( \1078 , \962 , \966 );
nand \U$999 ( \1079 , \1077 , \1078 );
nand \U$1000 ( \1080 , RIa139758_31, \109_nGa3 );
xor \U$1001 ( \1081 , \1079 , \1080 );
not \U$1002 ( \1082 , \1081 );
not \U$1003 ( \1083 , \1082 );
nand \U$1004 ( \1084 , RIa139758_31, \131_nG8b );
xor \U$1005 ( \1085 , \1084 , \977 );
xnor \U$1006 ( \1086 , \1085 , \1063 );
not \U$1007 ( \1087 , \1086 );
nand \U$1008 ( \1088 , RIa139758_31, \142_nG83 );
xor \U$1009 ( \1089 , \1088 , \1058 );
xnor \U$1010 ( \1090 , \1089 , \1055 );
not \U$1011 ( \1091 , \1090 );
nand \U$1012 ( \1092 , RIa139758_31, \179_nG63 );
not \U$1013 ( \1093 , \1092 );
xor \U$1014 ( \1094 , \988 , \992 );
not \U$1015 ( \1095 , \1094 );
not \U$1016 ( \1096 , \1095 );
or \U$1017 ( \1097 , \1093 , \1096 );
and \U$1018 ( \1098 , RIa139758_31, \170_nG5b );
xor \U$1019 ( \1099 , \982 , \983 );
xor \U$1020 ( \1100 , \1099 , \985 );
and \U$1021 ( \1101 , \1098 , \1100 );
nand \U$1022 ( \1102 , \1097 , \1101 );
not \U$1023 ( \1103 , \1092 );
nand \U$1024 ( \1104 , \1103 , \1094 );
and \U$1025 ( \1105 , \1102 , \1104 );
not \U$1026 ( \1106 , \1105 );
not \U$1027 ( \1107 , \1106 );
nand \U$1028 ( \1108 , RIa139758_31, \162_nG6b );
xor \U$1029 ( \1109 , \1108 , \1004 );
xnor \U$1030 ( \1110 , \1109 , \1010 );
not \U$1031 ( \1111 , \1110 );
or \U$1032 ( \1112 , \1107 , \1111 );
not \U$1033 ( \1113 , \1108 );
xor \U$1034 ( \1114 , \1010 , \1004 );
nand \U$1035 ( \1115 , \1113 , \1114 );
nand \U$1036 ( \1116 , \1112 , \1115 );
not \U$1037 ( \1117 , \1116 );
nand \U$1038 ( \1118 , RIa139758_31, \188_nG73 );
xor \U$1039 ( \1119 , \1118 , \1033 );
xnor \U$1040 ( \1120 , \1119 , \1022 );
not \U$1041 ( \1121 , \1120 );
or \U$1042 ( \1122 , \1117 , \1121 );
not \U$1043 ( \1123 , \1118 );
xor \U$1044 ( \1124 , \1033 , \1022 );
nand \U$1045 ( \1125 , \1123 , \1124 );
nand \U$1046 ( \1126 , \1122 , \1125 );
not \U$1047 ( \1127 , \1126 );
nand \U$1048 ( \1128 , RIa139758_31, \151_nG7b );
xor \U$1049 ( \1129 , \1128 , \1049 );
not \U$1050 ( \1130 , \1037 );
xnor \U$1051 ( \1131 , \1129 , \1130 );
not \U$1052 ( \1132 , \1131 );
or \U$1053 ( \1133 , \1127 , \1132 );
not \U$1054 ( \1134 , \1128 );
not \U$1055 ( \1135 , \1037 );
not \U$1056 ( \1136 , \1049 );
or \U$1057 ( \1137 , \1135 , \1136 );
nand \U$1058 ( \1138 , \1130 , \1050 );
nand \U$1059 ( \1139 , \1137 , \1138 );
nand \U$1060 ( \1140 , \1134 , \1139 );
nand \U$1061 ( \1141 , \1133 , \1140 );
not \U$1062 ( \1142 , \1141 );
or \U$1063 ( \1143 , \1091 , \1142 );
not \U$1064 ( \1144 , \1058 );
nand \U$1065 ( \1145 , \1144 , \1055 );
not \U$1066 ( \1146 , \1145 );
not \U$1067 ( \1147 , \1055 );
nand \U$1068 ( \1148 , \1147 , \1058 );
not \U$1069 ( \1149 , \1148 );
or \U$1070 ( \1150 , \1146 , \1149 );
not \U$1071 ( \1151 , \1088 );
nand \U$1072 ( \1152 , \1150 , \1151 );
nand \U$1073 ( \1153 , \1143 , \1152 );
not \U$1074 ( \1154 , \1153 );
or \U$1075 ( \1155 , \1087 , \1154 );
not \U$1076 ( \1156 , \1084 );
xor \U$1077 ( \1157 , \977 , \1063 );
nand \U$1078 ( \1158 , \1156 , \1157 );
nand \U$1079 ( \1159 , \1155 , \1158 );
not \U$1080 ( \1160 , \1159 );
nand \U$1081 ( \1161 , RIa139758_31, \91_nG93 );
xor \U$1082 ( \1162 , \1161 , \972 );
xnor \U$1083 ( \1163 , \1162 , \1069 );
not \U$1084 ( \1164 , \1163 );
or \U$1085 ( \1165 , \1160 , \1164 );
not \U$1086 ( \1166 , \1161 );
xor \U$1087 ( \1167 , \972 , \1069 );
nand \U$1088 ( \1168 , \1166 , \1167 );
nand \U$1089 ( \1169 , \1165 , \1168 );
not \U$1090 ( \1170 , \1169 );
nand \U$1091 ( \1171 , RIa139758_31, \100_nG9b );
xor \U$1092 ( \1172 , \1171 , \968 );
xnor \U$1093 ( \1173 , \1172 , \1075 );
not \U$1094 ( \1174 , \1173 );
or \U$1095 ( \1175 , \1170 , \1174 );
not \U$1096 ( \1176 , \1171 );
xor \U$1097 ( \1177 , \968 , \1075 );
nand \U$1098 ( \1178 , \1176 , \1177 );
nand \U$1099 ( \1179 , \1175 , \1178 );
not \U$1100 ( \1180 , \1179 );
or \U$1101 ( \1181 , \1083 , \1180 );
not \U$1102 ( \1182 , \1080 );
nand \U$1103 ( \1183 , \1182 , \1079 );
nand \U$1104 ( \1184 , \1181 , \1183 );
buf \U$1105 ( \1185 , \1184 );
not \U$1106 ( \1186 , \1081 );
not \U$1107 ( \1187 , \1179 );
or \U$1108 ( \1188 , \1186 , \1187 );
or \U$1109 ( \1189 , \1179 , \1081 );
nand \U$1110 ( \1190 , \1188 , \1189 );
buf \U$1111 ( \1191 , \1190 );
xor \U$1112 ( \1192 , \1173 , \1169 );
buf \U$1113 ( \1193 , \1192 );
xor \U$1114 ( \1194 , \1163 , \1159 );
buf \U$1115 ( \1195 , \1194 );
xor \U$1116 ( \1196 , \1086 , \1153 );
buf \U$1117 ( \1197 , \1196 );
xor \U$1118 ( \1198 , \1090 , \1141 );
buf \U$1119 ( \1199 , \1198 );
xor \U$1120 ( \1200 , \1131 , \1126 );
buf \U$1121 ( \1201 , \1200 );
xor \U$1122 ( \1202 , \1116 , \1120 );
buf \U$1123 ( \1203 , \1202 );
and \U$1124 ( \1204 , \1110 , \1106 );
not \U$1125 ( \1205 , \1110 );
and \U$1126 ( \1206 , \1205 , \1105 );
nor \U$1127 ( \1207 , \1204 , \1206 );
buf \U$1128 ( \1208 , \1207 );
xor \U$1129 ( \1209 , \1092 , \1101 );
xnor \U$1130 ( \1210 , \1209 , \1094 );
buf \U$1131 ( \1211 , \1210 );
xor \U$1132 ( \1212 , \1098 , \1100 );
buf \U$1133 ( \1213 , \1212 );
xor \U$1134 ( \1214 , \981 , \980 );
buf \U$1135 ( \1215 , \1214 );
xnor \U$1136 ( \1216 , \832 , \831 );
buf \U$1137 ( \1217 , \1216 );
not \U$1138 ( \1218 , \720 );
not \U$1139 ( \1219 , \718 );
or \U$1140 ( \1220 , \1218 , \1219 );
or \U$1141 ( \1221 , \718 , \720 );
nand \U$1142 ( \1222 , \1220 , \1221 );
buf \U$1143 ( \1223 , \1222 );
xor \U$1144 ( \1224 , \615 , \617 );
buf \U$1145 ( \1225 , \1224 );
not \U$1146 ( \1226 , \512 );
buf \U$1147 ( \1227 , \511 );
not \U$1148 ( \1228 , \1227 );
or \U$1149 ( \1229 , \1226 , \1228 );
or \U$1150 ( \1230 , \1227 , \512 );
nand \U$1151 ( \1231 , \1229 , \1230 );
buf \U$1152 ( \1232 , \1231 );
not \U$1153 ( \1233 , \410 );
not \U$1154 ( \1234 , \409 );
or \U$1155 ( \1235 , \1233 , \1234 );
xnor \U$1156 ( \1236 , \403 , \408 );
or \U$1157 ( \1237 , \1236 , \410 );
nand \U$1158 ( \1238 , \1235 , \1237 );
buf \U$1159 ( \1239 , \1238 );
and \U$1160 ( \1240 , \282 , \297 );
and \U$1161 ( \1241 , \299 , \283 );
nor \U$1162 ( \1242 , \1240 , \1241 );
not \U$1163 ( \1243 , \1242 );
not \U$1164 ( \1244 , \291 );
or \U$1165 ( \1245 , \1243 , \1244 );
or \U$1166 ( \1246 , \291 , \1242 );
nand \U$1167 ( \1247 , \1245 , \1246 );
buf \U$1168 ( \1248 , \1247 );
nand \U$1169 ( \1249 , RIa139b18_39, \170_nG5b );
not \U$1170 ( \1250 , \1249 );
and \U$1171 ( \1251 , RIa139b90_40, \179_nG63 );
not \U$1172 ( \1252 , \1251 );
or \U$1173 ( \1253 , \1250 , \1252 );
or \U$1174 ( \1254 , \1249 , \1251 );
nand \U$1175 ( \1255 , \1253 , \1254 );
buf \U$1176 ( \1256 , \1255 );
not \U$1177 ( \1257 , \296 );
buf \U$1178 ( \1258 , \1257 );
endmodule

