//
// Conformal-LEC Version 20.10-d211 (31-Aug-2020)
//
module top(RI8929640_33,RI8929dc0_49,RI89296b8_34,RI8929e38_50,RI8929730_35,RI8929eb0_51,RI89297a8_36,RI8929f28_52,RI8929820_37,
        RI8929fa0_53,RI8929898_38,RI892a018_54,RI8929910_39,RI892a090_55,RI8929988_40,RI892a108_56,RI8929a00_41,RI892a180_57,RI8929a78_42,
        RI892a1f8_58,RI8929af0_43,RI892a270_59,RI8929b68_44,RI892a2e8_60,RI8929be0_45,RI892a360_61,RI8929c58_46,RI892a3d8_62,RI8929cd0_47,
        RI892a450_63,RI8929d48_48,RI892a4c8_64,RI8928e48_16,RI89295c8_32,RI8928dd0_15,RI8929550_31,RI8928d58_14,RI89294d8_30,RI8928ce0_13,
        RI8929460_29,RI8928c68_12,RI89293e8_28,RI8928bf0_11,RI8929370_27,RI8928b78_10,RI89292f8_26,RI8928b00_9,RI8929280_25,RI8928a88_8,
        RI8929208_24,RI8928a10_7,RI8929190_23,RI8928998_6,RI8929118_22,RI8928920_5,RI89290a0_21,RI89288a8_4,RI8929028_20,RI8928830_3,
        RI8928fb0_19,RI89287b8_2,RI8928f38_18,RI8928740_1,RI8928ec0_17,R_41_7a88898,R_42_7a83a80,R_43_7a83bd0,R_44_7a87788,R_45_7a88be0,
        R_46_7a81ef0,R_47_7a889e8,R_48_7a84a40,R_49_7a882b0,R_4a_7a82c10,R_4b_7a82d60,R_4c_7a87b78,R_4d_7a84b90,R_4e_7a86f00,R_4f_7a84ce0,
        R_50_7a87440,R_51_7a88160,R_52_7a83d20,R_53_7a88c88,R_54_7a82040,R_55_7a84e30,R_56_7a876e0,R_57_7a87f68,R_58_7a82eb0,R_59_7a88dd8,
        R_5a_7a86e58,R_5b_7a83e70);
input RI8929640_33,RI8929dc0_49,RI89296b8_34,RI8929e38_50,RI8929730_35,RI8929eb0_51,RI89297a8_36,RI8929f28_52,RI8929820_37,
        RI8929fa0_53,RI8929898_38,RI892a018_54,RI8929910_39,RI892a090_55,RI8929988_40,RI892a108_56,RI8929a00_41,RI892a180_57,RI8929a78_42,
        RI892a1f8_58,RI8929af0_43,RI892a270_59,RI8929b68_44,RI892a2e8_60,RI8929be0_45,RI892a360_61,RI8929c58_46,RI892a3d8_62,RI8929cd0_47,
        RI892a450_63,RI8929d48_48,RI892a4c8_64,RI8928e48_16,RI89295c8_32,RI8928dd0_15,RI8929550_31,RI8928d58_14,RI89294d8_30,RI8928ce0_13,
        RI8929460_29,RI8928c68_12,RI89293e8_28,RI8928bf0_11,RI8929370_27,RI8928b78_10,RI89292f8_26,RI8928b00_9,RI8929280_25,RI8928a88_8,
        RI8929208_24,RI8928a10_7,RI8929190_23,RI8928998_6,RI8929118_22,RI8928920_5,RI89290a0_21,RI89288a8_4,RI8929028_20,RI8928830_3,
        RI8928fb0_19,RI89287b8_2,RI8928f38_18,RI8928740_1,RI8928ec0_17;
output R_41_7a88898,R_42_7a83a80,R_43_7a83bd0,R_44_7a87788,R_45_7a88be0,R_46_7a81ef0,R_47_7a889e8,R_48_7a84a40,R_49_7a882b0,
        R_4a_7a82c10,R_4b_7a82d60,R_4c_7a87b78,R_4d_7a84b90,R_4e_7a86f00,R_4f_7a84ce0,R_50_7a87440,R_51_7a88160,R_52_7a83d20,R_53_7a88c88,
        R_54_7a82040,R_55_7a84e30,R_56_7a876e0,R_57_7a87f68,R_58_7a82eb0,R_59_7a88dd8,R_5a_7a86e58,R_5b_7a83e70;

wire \92 , \93 , \94 , \95 , \96 , \97 , \98 , \99 , \100 ,
         \101 , \102 , \103 , \104 , \105 , \106 , \107 , \108_N$1 , \109_N$2 , \110_N$3 ,
         \111_N$4 , \112_N$5 , \113_N$6 , \114_N$7 , \115_N$8 , \116_N$9 , \117_N$10 , \118_N$11 , \119_N$12 , \120_N$13 ,
         \121_N$14 , \122_N$15 , \123_N$16 , \124_ZERO , \125_ONE , \126 , \127 , \128 , \129 , \130 ,
         \131 , \132 , \133 , \134 , \135 , \136 , \137 , \138 , \139 , \140 ,
         \141 , \142 , \143 , \144 , \145 , \146 , \147 , \148 , \149 , \150 ,
         \151 , \152 , \153 , \154 , \155 , \156 , \157 , \158 , \159 , \160 ,
         \161 , \162 , \163 , \164 , \165 , \166 , \167 , \168 , \169 , \170 ,
         \171 , \172 , \173 , \174 , \175 , \176 , \177 , \178 , \179 , \180 ,
         \181 , \182 , \183 , \184 , \185 , \186 , \187 , \188 , \189 , \190 ,
         \191 , \192 , \193 , \194 , \195 , \196 , \197 , \198 , \199 , \200 ,
         \201 , \202 , \203 , \204 , \205 , \206 , \207 , \208 , \209 , \210 ,
         \211 , \212 , \213 , \214 , \215 , \216 , \217 , \218 , \219 , \220 ,
         \221 , \222 , \223 , \224 , \225 , \226 , \227 , \228 , \229 , \230 ,
         \231 , \232 , \233 , \234 , \235 , \236 , \237 , \238 , \239 , \240 ,
         \241 , \242 , \243 , \244 , \245 , \246 , \247 , \248 , \249 , \250 ,
         \251 , \252 , \253 , \254 , \255 , \256 , \257 , \258 , \259 , \260 ,
         \261 , \262 , \263 , \264 , \265 , \266 , \267 , \268 , \269 , \270 ,
         \271 , \272 , \273 , \274 , \275 , \276 , \277 , \278 , \279 , \280 ,
         \281 , \282 , \283 , \284 , \285 , \286 , \287 , \288 , \289 , \290 ,
         \291 , \292 , \293 , \294 , \295 , \296 , \297 , \298 , \299 , \300 ,
         \301 , \302 , \303 , \304 , \305 , \306 , \307 , \308 , \309 , \310 ,
         \311 , \312 , \313 , \314 , \315 , \316 , \317 , \318 , \319 , \320 ,
         \321 , \322 , \323 , \324 , \325 , \326 , \327 , \328 , \329 , \330 ,
         \331 , \332 , \333 , \334 , \335 , \336 , \337 , \338 , \339 , \340 ,
         \341 , \342 , \343 , \344 , \345 , \346 , \347 , \348 , \349 , \350 ,
         \351 , \352 , \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 ,
         \361 , \362 , \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 ,
         \371 , \372 , \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 ,
         \381 , \382 , \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 ,
         \391 , \392 , \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 ,
         \401 , \402 , \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 ,
         \411 , \412 , \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 ,
         \421 , \422 , \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 ,
         \431 , \432 , \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 ,
         \441 , \442 , \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 ,
         \451 , \452 , \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 ,
         \461 , \462 , \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 ,
         \471 , \472 , \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 ,
         \481 , \482 , \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 ,
         \491 , \492 , \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 ,
         \501 , \502 , \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 ,
         \511 , \512 , \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 ,
         \521 , \522 , \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 ,
         \531 , \532 , \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 ,
         \541 , \542 , \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 ,
         \551 , \552 , \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 ,
         \561 , \562 , \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 ,
         \571 , \572 , \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 ,
         \581 , \582 , \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 ,
         \591 , \592 , \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 ,
         \601 , \602 , \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 ,
         \611 , \612 , \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 ,
         \621 , \622 , \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 ,
         \631 , \632 , \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 ,
         \641 , \642 , \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 ,
         \651 , \652 , \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 ,
         \661 , \662 , \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 ,
         \671 , \672 , \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 ,
         \681 , \682 , \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 ,
         \691 , \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 ,
         \701 , \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 ,
         \711 , \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 ,
         \721 , \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 ,
         \731 , \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 ,
         \741 , \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 ,
         \751 , \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 ,
         \761 , \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 ,
         \771 , \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 ,
         \781 , \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 ,
         \791 , \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 ,
         \801 , \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 ,
         \811 , \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 ,
         \821 , \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 ,
         \831 , \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 ,
         \841 , \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 ,
         \851 , \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 ,
         \861 , \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 ,
         \871 , \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 ,
         \881 , \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 ,
         \891 , \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 ,
         \901 , \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 ,
         \911 , \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 ,
         \921 , \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 ,
         \931 , \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 ,
         \941 , \942_nG3a2 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 ,
         \951 , \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 ,
         \961 , \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 ,
         \971 , \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 ,
         \981 , \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 ,
         \991 , \992 , \993 , \994_nG3d6 , \995 , \996 , \997 , \998 , \999 , \1000 ,
         \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 ,
         \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 ,
         \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 ,
         \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 ,
         \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 ,
         \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 ,
         \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 ,
         \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 ,
         \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 ,
         \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 ,
         \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 ,
         \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 ,
         \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 ,
         \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 ,
         \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 ,
         \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 ,
         \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 ,
         \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178_nG48e , \1179 , \1180 ,
         \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 ,
         \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 ,
         \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 ,
         \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 ,
         \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 ,
         \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 ,
         \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 ,
         \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 ,
         \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 ,
         \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 ,
         \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 ,
         \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 ,
         \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 ,
         \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 ,
         \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 ,
         \1331 , \1332 , \1333_nG529 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 ,
         \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 ,
         \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 ,
         \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 ,
         \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 ,
         \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 ,
         \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 ,
         \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 ,
         \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 ,
         \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 ,
         \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 ,
         \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 ,
         \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 ,
         \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 ,
         \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 ,
         \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 ,
         \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500_nG5d0 ,
         \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 ,
         \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 ,
         \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 ,
         \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 ,
         \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 ,
         \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 ,
         \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 ,
         \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 ,
         \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 ,
         \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 ,
         \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 ,
         \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 ,
         \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 ,
         \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 ,
         \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 ,
         \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 ,
         \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 ,
         \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679_nG683 , \1680 ,
         \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 ,
         \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 ,
         \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 ,
         \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 ,
         \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 ,
         \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 ,
         \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 ,
         \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 ,
         \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 ,
         \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 ,
         \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 ,
         \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 ,
         \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 ,
         \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 ,
         \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 ,
         \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 ,
         \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 ,
         \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 ,
         \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870_nG742 ,
         \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 ,
         \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 ,
         \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 ,
         \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 ,
         \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 ,
         \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 ,
         \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 ,
         \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 ,
         \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 ,
         \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 ,
         \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 ,
         \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 ,
         \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 ,
         \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 ,
         \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 ,
         \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 ,
         \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 ,
         \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 ,
         \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 ,
         \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 ,
         \2071 , \2072 , \2073_nG80d , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 ,
         \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 ,
         \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 ,
         \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 ,
         \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 ,
         \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 ,
         \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 ,
         \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 ,
         \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 ,
         \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 ,
         \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 ,
         \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 ,
         \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 ,
         \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 ,
         \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 ,
         \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 ,
         \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 ,
         \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 ,
         \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 ,
         \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 ,
         \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 ,
         \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288_nG8e4 , \2289 , \2290 ,
         \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 ,
         \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 ,
         \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 ,
         \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 ,
         \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 ,
         \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 ,
         \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 ,
         \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 ,
         \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 ,
         \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 ,
         \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 ,
         \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 ,
         \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 ,
         \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 ,
         \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 ,
         \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 ,
         \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 ,
         \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 ,
         \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 ,
         \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 ,
         \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 ,
         \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 ,
         \2511 , \2512 , \2513 , \2514 , \2515_nG9c7 , \2516 , \2517 , \2518 , \2519 , \2520 ,
         \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 ,
         \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 ,
         \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 ,
         \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 ,
         \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 ,
         \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 ,
         \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 ,
         \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 ,
         \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 ,
         \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 ,
         \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 ,
         \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 ,
         \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 ,
         \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 ,
         \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 ,
         \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 ,
         \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 ,
         \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 ,
         \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 ,
         \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 ,
         \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 ,
         \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 ,
         \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 ,
         \2751 , \2752 , \2753 , \2754_nGab6 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 ,
         \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 ,
         \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 ,
         \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 ,
         \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 ,
         \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 ,
         \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 ,
         \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 ,
         \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 ,
         \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 ,
         \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 ,
         \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 ,
         \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 ,
         \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 ,
         \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 ,
         \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 ,
         \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 ,
         \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 ,
         \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 ,
         \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 ,
         \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 ,
         \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 ,
         \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 ,
         \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 ,
         \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 ,
         \3001 , \3002 , \3003 , \3004 , \3005_nGbb1 , \3006 , \3007 , \3008 , \3009 , \3010 ,
         \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 ,
         \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 ,
         \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 ,
         \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 ,
         \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 ,
         \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 ,
         \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 ,
         \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 ,
         \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 ,
         \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 ,
         \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 ,
         \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 ,
         \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 ,
         \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 ,
         \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 ,
         \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 ,
         \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 ,
         \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 ,
         \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 ,
         \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 ,
         \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 ,
         \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 ,
         \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 ,
         \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 ,
         \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 ,
         \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268_nGcb8 , \3269 , \3270 ,
         \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 ,
         \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 ,
         \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 ,
         \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 ,
         \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 ,
         \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 ,
         \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 ,
         \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 ,
         \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 ,
         \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 ,
         \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 ,
         \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 ,
         \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 ,
         \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 ,
         \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 ,
         \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 ,
         \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 ,
         \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 ,
         \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 ,
         \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 ,
         \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 ,
         \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 ,
         \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 ,
         \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 ,
         \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 ,
         \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 ,
         \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 ,
         \3541 , \3542 , \3543_nGdcb , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 ,
         \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 ,
         \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 ,
         \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 ,
         \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 ,
         \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 ,
         \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 ,
         \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 ,
         \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 ,
         \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 ,
         \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 ,
         \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 ,
         \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 ,
         \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 ,
         \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 ,
         \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 ,
         \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 ,
         \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 ,
         \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 ,
         \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 ,
         \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 ,
         \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 ,
         \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 ,
         \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 ,
         \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 ,
         \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 ,
         \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 ,
         \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 ,
         \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830_nGeea ,
         \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 ,
         \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 ,
         \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 ,
         \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 ,
         \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 ,
         \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 ,
         \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 ,
         \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 ,
         \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 ,
         \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 ,
         \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 ,
         \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 ,
         \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 ,
         \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 ,
         \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 ,
         \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 ,
         \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 ,
         \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 ,
         \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 ,
         \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 ,
         \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 ,
         \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 ,
         \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 ,
         \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 ,
         \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 ,
         \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 ,
         \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 ,
         \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 ,
         \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 ,
         \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129_nG1015 , \4130 ,
         \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 ,
         \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 ,
         \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 ,
         \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 ,
         \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 ,
         \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 ,
         \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 ,
         \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 ,
         \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 ,
         \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 ,
         \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 ,
         \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 ,
         \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 ,
         \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 ,
         \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 ,
         \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 ,
         \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 ,
         \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 ,
         \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 ,
         \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 ,
         \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 ,
         \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 ,
         \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 ,
         \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 ,
         \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 ,
         \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 ,
         \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 ,
         \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 ,
         \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 ,
         \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 ,
         \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 ,
         \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 ,
         \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 ,
         \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 ,
         \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 ,
         \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 ,
         \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 ,
         \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 ,
         \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 ;
buf \U$labaj468 ( R_41_7a88898, \4439 );
buf \U$labaj469 ( R_42_7a83a80, \4442 );
buf \U$labaj470 ( R_43_7a83bd0, \4445 );
buf \U$labaj471 ( R_44_7a87788, \4448 );
buf \U$labaj472 ( R_45_7a88be0, \4451 );
buf \U$labaj473 ( R_46_7a81ef0, \4454 );
buf \U$labaj474 ( R_47_7a889e8, \4457 );
buf \U$labaj475 ( R_48_7a84a40, \4460 );
buf \U$labaj476 ( R_49_7a882b0, \4463 );
buf \U$labaj477 ( R_4a_7a82c10, \4466 );
buf \U$labaj478 ( R_4b_7a82d60, \4469 );
buf \U$labaj479 ( R_4c_7a87b78, \4472 );
buf \U$labaj480 ( R_4d_7a84b90, \4475 );
buf \U$labaj481 ( R_4e_7a86f00, \4478 );
buf \U$labaj482 ( R_4f_7a84ce0, \4481 );
buf \U$labaj483 ( R_50_7a87440, \4484 );
buf \U$labaj484 ( R_51_7a88160, \4487 );
buf \U$labaj485 ( R_52_7a83d20, \4490 );
buf \U$labaj486 ( R_53_7a88c88, \4493 );
buf \U$labaj487 ( R_54_7a82040, \4496 );
buf \U$labaj488 ( R_55_7a84e30, \4499 );
buf \U$labaj489 ( R_56_7a876e0, \4502 );
buf \U$labaj490 ( R_57_7a87f68, \4505 );
buf \U$labaj491 ( R_58_7a82eb0, \4508 );
buf \U$labaj492 ( R_59_7a88dd8, \4511 );
buf \U$labaj493 ( R_5a_7a86e58, \4514 );
buf \U$labaj494 ( R_5b_7a83e70, \4517 );
buf \U$1 ( \126 , RI8929640_33);
buf \U$2 ( \127 , RI8929dc0_49);
and \U$3 ( \128 , \126 , \127 );
buf \U$4 ( \129 , RI89296b8_34);
buf \U$5 ( \130 , RI8929e38_50);
and \U$6 ( \131 , \129 , \130 );
buf \U$7 ( \132 , RI8929730_35);
buf \U$8 ( \133 , RI8929eb0_51);
and \U$9 ( \134 , \132 , \133 );
buf \U$10 ( \135 , RI89297a8_36);
buf \U$11 ( \136 , RI8929f28_52);
and \U$12 ( \137 , \135 , \136 );
buf \U$13 ( \138 , RI8929820_37);
buf \U$14 ( \139 , RI8929fa0_53);
and \U$15 ( \140 , \138 , \139 );
buf \U$16 ( \141 , RI8929898_38);
buf \U$17 ( \142 , RI892a018_54);
and \U$18 ( \143 , \141 , \142 );
buf \U$19 ( \144 , RI8929910_39);
buf \U$20 ( \145 , RI892a090_55);
and \U$21 ( \146 , \144 , \145 );
buf \U$22 ( \147 , RI8929988_40);
buf \U$23 ( \148 , RI892a108_56);
and \U$24 ( \149 , \147 , \148 );
buf \U$25 ( \150 , RI8929a00_41);
buf \U$26 ( \151 , RI892a180_57);
and \U$27 ( \152 , \150 , \151 );
buf \U$28 ( \153 , RI8929a78_42);
buf \U$29 ( \154 , RI892a1f8_58);
and \U$30 ( \155 , \153 , \154 );
buf \U$31 ( \156 , RI8929af0_43);
buf \U$32 ( \157 , RI892a270_59);
and \U$33 ( \158 , \156 , \157 );
buf \U$34 ( \159 , RI8929b68_44);
buf \U$35 ( \160 , RI892a2e8_60);
and \U$36 ( \161 , \159 , \160 );
buf \U$37 ( \162 , RI8929be0_45);
buf \U$38 ( \163 , RI892a360_61);
and \U$39 ( \164 , \162 , \163 );
buf \U$40 ( \165 , RI8929c58_46);
buf \U$41 ( \166 , RI892a3d8_62);
and \U$42 ( \167 , \165 , \166 );
buf \U$43 ( \168 , RI8929cd0_47);
buf \U$44 ( \169 , RI892a450_63);
and \U$45 ( \170 , \168 , \169 );
buf \U$46 ( \171 , RI8929d48_48);
buf \U$47 ( \172 , RI892a4c8_64);
and \U$48 ( \173 , \171 , \172 );
and \U$49 ( \174 , \169 , \173 );
and \U$50 ( \175 , \168 , \173 );
or \U$51 ( \176 , \170 , \174 , \175 );
and \U$52 ( \177 , \166 , \176 );
and \U$53 ( \178 , \165 , \176 );
or \U$54 ( \179 , \167 , \177 , \178 );
and \U$55 ( \180 , \163 , \179 );
and \U$56 ( \181 , \162 , \179 );
or \U$57 ( \182 , \164 , \180 , \181 );
and \U$58 ( \183 , \160 , \182 );
and \U$59 ( \184 , \159 , \182 );
or \U$60 ( \185 , \161 , \183 , \184 );
and \U$61 ( \186 , \157 , \185 );
and \U$62 ( \187 , \156 , \185 );
or \U$63 ( \188 , \158 , \186 , \187 );
and \U$64 ( \189 , \154 , \188 );
and \U$65 ( \190 , \153 , \188 );
or \U$66 ( \191 , \155 , \189 , \190 );
and \U$67 ( \192 , \151 , \191 );
and \U$68 ( \193 , \150 , \191 );
or \U$69 ( \194 , \152 , \192 , \193 );
and \U$70 ( \195 , \148 , \194 );
and \U$71 ( \196 , \147 , \194 );
or \U$72 ( \197 , \149 , \195 , \196 );
and \U$73 ( \198 , \145 , \197 );
and \U$74 ( \199 , \144 , \197 );
or \U$75 ( \200 , \146 , \198 , \199 );
and \U$76 ( \201 , \142 , \200 );
and \U$77 ( \202 , \141 , \200 );
or \U$78 ( \203 , \143 , \201 , \202 );
and \U$79 ( \204 , \139 , \203 );
and \U$80 ( \205 , \138 , \203 );
or \U$81 ( \206 , \140 , \204 , \205 );
and \U$82 ( \207 , \136 , \206 );
and \U$83 ( \208 , \135 , \206 );
or \U$84 ( \209 , \137 , \207 , \208 );
and \U$85 ( \210 , \133 , \209 );
and \U$86 ( \211 , \132 , \209 );
or \U$87 ( \212 , \134 , \210 , \211 );
and \U$88 ( \213 , \130 , \212 );
and \U$89 ( \214 , \129 , \212 );
or \U$90 ( \215 , \131 , \213 , \214 );
and \U$91 ( \216 , \127 , \215 );
and \U$92 ( \217 , \126 , \215 );
or \U$93 ( \218 , \128 , \216 , \217 );
buf \U$94 ( \219 , \218 );
buf \U$95 ( \220 , \219 );
buf \U$97 ( \221 , RI8928e48_16);
buf \U$98 ( \222 , RI89295c8_32);
and \U$99 ( \223 , \221 , \222 );
buf \U$100 ( \224 , \223 );
not \U$101 ( \225 , \224 );
buf \U$102 ( \226 , RI8928dd0_15);
and \U$103 ( \227 , \226 , \222 );
buf \U$104 ( \228 , RI8929550_31);
and \U$105 ( \229 , \221 , \228 );
xor \U$106 ( \230 , \227 , \229 );
buf \U$107 ( \231 , \230 );
buf \U$108 ( \232 , RI8928d58_14);
and \U$109 ( \233 , \232 , \222 );
and \U$110 ( \234 , \226 , \228 );
xor \U$111 ( \235 , \233 , \234 );
and \U$112 ( \236 , \227 , \229 );
xor \U$113 ( \237 , \235 , \236 );
buf \U$114 ( \238 , RI89294d8_30);
and \U$115 ( \239 , \221 , \238 );
xor \U$116 ( \240 , \237 , \239 );
buf \U$117 ( \241 , \240 );
buf \U$118 ( \242 , RI8928ce0_13);
and \U$119 ( \243 , \242 , \222 );
and \U$120 ( \244 , \232 , \228 );
xor \U$121 ( \245 , \243 , \244 );
and \U$122 ( \246 , \233 , \234 );
and \U$123 ( \247 , \235 , \236 );
or \U$124 ( \248 , \246 , \247 );
xor \U$125 ( \249 , \245 , \248 );
and \U$126 ( \250 , \226 , \238 );
xor \U$127 ( \251 , \249 , \250 );
and \U$128 ( \252 , \237 , \239 );
xor \U$129 ( \253 , \251 , \252 );
buf \U$130 ( \254 , RI8929460_29);
and \U$131 ( \255 , \221 , \254 );
xor \U$132 ( \256 , \253 , \255 );
buf \U$133 ( \257 , \256 );
buf \U$134 ( \258 , RI8928c68_12);
and \U$135 ( \259 , \258 , \222 );
and \U$136 ( \260 , \242 , \228 );
xor \U$137 ( \261 , \259 , \260 );
and \U$138 ( \262 , \243 , \244 );
and \U$139 ( \263 , \245 , \248 );
or \U$140 ( \264 , \262 , \263 );
xor \U$141 ( \265 , \261 , \264 );
and \U$142 ( \266 , \232 , \238 );
xor \U$143 ( \267 , \265 , \266 );
and \U$144 ( \268 , \249 , \250 );
and \U$145 ( \269 , \251 , \252 );
or \U$146 ( \270 , \268 , \269 );
xor \U$147 ( \271 , \267 , \270 );
and \U$148 ( \272 , \226 , \254 );
xor \U$149 ( \273 , \271 , \272 );
and \U$150 ( \274 , \253 , \255 );
xor \U$151 ( \275 , \273 , \274 );
buf \U$152 ( \276 , RI89293e8_28);
and \U$153 ( \277 , \221 , \276 );
xor \U$154 ( \278 , \275 , \277 );
buf \U$155 ( \279 , \278 );
buf \U$156 ( \280 , RI8928bf0_11);
and \U$157 ( \281 , \280 , \222 );
and \U$158 ( \282 , \258 , \228 );
xor \U$159 ( \283 , \281 , \282 );
and \U$160 ( \284 , \259 , \260 );
and \U$161 ( \285 , \261 , \264 );
or \U$162 ( \286 , \284 , \285 );
xor \U$163 ( \287 , \283 , \286 );
and \U$164 ( \288 , \242 , \238 );
xor \U$165 ( \289 , \287 , \288 );
and \U$166 ( \290 , \265 , \266 );
and \U$167 ( \291 , \267 , \270 );
or \U$168 ( \292 , \290 , \291 );
xor \U$169 ( \293 , \289 , \292 );
and \U$170 ( \294 , \232 , \254 );
xor \U$171 ( \295 , \293 , \294 );
and \U$172 ( \296 , \271 , \272 );
and \U$173 ( \297 , \273 , \274 );
or \U$174 ( \298 , \296 , \297 );
xor \U$175 ( \299 , \295 , \298 );
and \U$176 ( \300 , \226 , \276 );
xor \U$177 ( \301 , \299 , \300 );
and \U$178 ( \302 , \275 , \277 );
xor \U$179 ( \303 , \301 , \302 );
buf \U$180 ( \304 , RI8929370_27);
and \U$181 ( \305 , \221 , \304 );
xor \U$182 ( \306 , \303 , \305 );
buf \U$183 ( \307 , \306 );
buf \U$184 ( \308 , RI8928b78_10);
and \U$185 ( \309 , \308 , \222 );
and \U$186 ( \310 , \280 , \228 );
xor \U$187 ( \311 , \309 , \310 );
and \U$188 ( \312 , \281 , \282 );
and \U$189 ( \313 , \283 , \286 );
or \U$190 ( \314 , \312 , \313 );
xor \U$191 ( \315 , \311 , \314 );
and \U$192 ( \316 , \258 , \238 );
xor \U$193 ( \317 , \315 , \316 );
and \U$194 ( \318 , \287 , \288 );
and \U$195 ( \319 , \289 , \292 );
or \U$196 ( \320 , \318 , \319 );
xor \U$197 ( \321 , \317 , \320 );
and \U$198 ( \322 , \242 , \254 );
xor \U$199 ( \323 , \321 , \322 );
and \U$200 ( \324 , \293 , \294 );
and \U$201 ( \325 , \295 , \298 );
or \U$202 ( \326 , \324 , \325 );
xor \U$203 ( \327 , \323 , \326 );
and \U$204 ( \328 , \232 , \276 );
xor \U$205 ( \329 , \327 , \328 );
and \U$206 ( \330 , \299 , \300 );
and \U$207 ( \331 , \301 , \302 );
or \U$208 ( \332 , \330 , \331 );
xor \U$209 ( \333 , \329 , \332 );
and \U$210 ( \334 , \226 , \304 );
xor \U$211 ( \335 , \333 , \334 );
and \U$212 ( \336 , \303 , \305 );
xor \U$213 ( \337 , \335 , \336 );
buf \U$214 ( \338 , RI89292f8_26);
and \U$215 ( \339 , \221 , \338 );
xor \U$216 ( \340 , \337 , \339 );
buf \U$217 ( \341 , \340 );
buf \U$218 ( \342 , RI8928b00_9);
and \U$219 ( \343 , \342 , \222 );
and \U$220 ( \344 , \308 , \228 );
xor \U$221 ( \345 , \343 , \344 );
and \U$222 ( \346 , \309 , \310 );
and \U$223 ( \347 , \311 , \314 );
or \U$224 ( \348 , \346 , \347 );
xor \U$225 ( \349 , \345 , \348 );
and \U$226 ( \350 , \280 , \238 );
xor \U$227 ( \351 , \349 , \350 );
and \U$228 ( \352 , \315 , \316 );
and \U$229 ( \353 , \317 , \320 );
or \U$230 ( \354 , \352 , \353 );
xor \U$231 ( \355 , \351 , \354 );
and \U$232 ( \356 , \258 , \254 );
xor \U$233 ( \357 , \355 , \356 );
and \U$234 ( \358 , \321 , \322 );
and \U$235 ( \359 , \323 , \326 );
or \U$236 ( \360 , \358 , \359 );
xor \U$237 ( \361 , \357 , \360 );
and \U$238 ( \362 , \242 , \276 );
xor \U$239 ( \363 , \361 , \362 );
and \U$240 ( \364 , \327 , \328 );
and \U$241 ( \365 , \329 , \332 );
or \U$242 ( \366 , \364 , \365 );
xor \U$243 ( \367 , \363 , \366 );
and \U$244 ( \368 , \232 , \304 );
xor \U$245 ( \369 , \367 , \368 );
and \U$246 ( \370 , \333 , \334 );
and \U$247 ( \371 , \335 , \336 );
or \U$248 ( \372 , \370 , \371 );
xor \U$249 ( \373 , \369 , \372 );
and \U$250 ( \374 , \226 , \338 );
xor \U$251 ( \375 , \373 , \374 );
and \U$252 ( \376 , \337 , \339 );
xor \U$253 ( \377 , \375 , \376 );
buf \U$254 ( \378 , RI8929280_25);
and \U$255 ( \379 , \221 , \378 );
xor \U$256 ( \380 , \377 , \379 );
buf \U$257 ( \381 , \380 );
buf \U$258 ( \382 , RI8928a88_8);
and \U$259 ( \383 , \382 , \222 );
and \U$260 ( \384 , \342 , \228 );
xor \U$261 ( \385 , \383 , \384 );
and \U$262 ( \386 , \343 , \344 );
and \U$263 ( \387 , \345 , \348 );
or \U$264 ( \388 , \386 , \387 );
xor \U$265 ( \389 , \385 , \388 );
and \U$266 ( \390 , \308 , \238 );
xor \U$267 ( \391 , \389 , \390 );
and \U$268 ( \392 , \349 , \350 );
and \U$269 ( \393 , \351 , \354 );
or \U$270 ( \394 , \392 , \393 );
xor \U$271 ( \395 , \391 , \394 );
and \U$272 ( \396 , \280 , \254 );
xor \U$273 ( \397 , \395 , \396 );
and \U$274 ( \398 , \355 , \356 );
and \U$275 ( \399 , \357 , \360 );
or \U$276 ( \400 , \398 , \399 );
xor \U$277 ( \401 , \397 , \400 );
and \U$278 ( \402 , \258 , \276 );
xor \U$279 ( \403 , \401 , \402 );
and \U$280 ( \404 , \361 , \362 );
and \U$281 ( \405 , \363 , \366 );
or \U$282 ( \406 , \404 , \405 );
xor \U$283 ( \407 , \403 , \406 );
and \U$284 ( \408 , \242 , \304 );
xor \U$285 ( \409 , \407 , \408 );
and \U$286 ( \410 , \367 , \368 );
and \U$287 ( \411 , \369 , \372 );
or \U$288 ( \412 , \410 , \411 );
xor \U$289 ( \413 , \409 , \412 );
and \U$290 ( \414 , \232 , \338 );
xor \U$291 ( \415 , \413 , \414 );
and \U$292 ( \416 , \373 , \374 );
and \U$293 ( \417 , \375 , \376 );
or \U$294 ( \418 , \416 , \417 );
xor \U$295 ( \419 , \415 , \418 );
and \U$296 ( \420 , \226 , \378 );
xor \U$297 ( \421 , \419 , \420 );
and \U$298 ( \422 , \377 , \379 );
xor \U$299 ( \423 , \421 , \422 );
buf \U$300 ( \424 , RI8929208_24);
and \U$301 ( \425 , \221 , \424 );
xor \U$302 ( \426 , \423 , \425 );
buf \U$303 ( \427 , \426 );
buf \U$304 ( \428 , RI8928a10_7);
and \U$305 ( \429 , \428 , \222 );
and \U$306 ( \430 , \382 , \228 );
xor \U$307 ( \431 , \429 , \430 );
and \U$308 ( \432 , \383 , \384 );
and \U$309 ( \433 , \385 , \388 );
or \U$310 ( \434 , \432 , \433 );
xor \U$311 ( \435 , \431 , \434 );
and \U$312 ( \436 , \342 , \238 );
xor \U$313 ( \437 , \435 , \436 );
and \U$314 ( \438 , \389 , \390 );
and \U$315 ( \439 , \391 , \394 );
or \U$316 ( \440 , \438 , \439 );
xor \U$317 ( \441 , \437 , \440 );
and \U$318 ( \442 , \308 , \254 );
xor \U$319 ( \443 , \441 , \442 );
and \U$320 ( \444 , \395 , \396 );
and \U$321 ( \445 , \397 , \400 );
or \U$322 ( \446 , \444 , \445 );
xor \U$323 ( \447 , \443 , \446 );
and \U$324 ( \448 , \280 , \276 );
xor \U$325 ( \449 , \447 , \448 );
and \U$326 ( \450 , \401 , \402 );
and \U$327 ( \451 , \403 , \406 );
or \U$328 ( \452 , \450 , \451 );
xor \U$329 ( \453 , \449 , \452 );
and \U$330 ( \454 , \258 , \304 );
xor \U$331 ( \455 , \453 , \454 );
and \U$332 ( \456 , \407 , \408 );
and \U$333 ( \457 , \409 , \412 );
or \U$334 ( \458 , \456 , \457 );
xor \U$335 ( \459 , \455 , \458 );
and \U$336 ( \460 , \242 , \338 );
xor \U$337 ( \461 , \459 , \460 );
and \U$338 ( \462 , \413 , \414 );
and \U$339 ( \463 , \415 , \418 );
or \U$340 ( \464 , \462 , \463 );
xor \U$341 ( \465 , \461 , \464 );
and \U$342 ( \466 , \232 , \378 );
xor \U$343 ( \467 , \465 , \466 );
and \U$344 ( \468 , \419 , \420 );
and \U$345 ( \469 , \421 , \422 );
or \U$346 ( \470 , \468 , \469 );
xor \U$347 ( \471 , \467 , \470 );
and \U$348 ( \472 , \226 , \424 );
xor \U$349 ( \473 , \471 , \472 );
and \U$350 ( \474 , \423 , \425 );
xor \U$351 ( \475 , \473 , \474 );
buf \U$352 ( \476 , RI8929190_23);
and \U$353 ( \477 , \221 , \476 );
xor \U$354 ( \478 , \475 , \477 );
buf \U$355 ( \479 , \478 );
buf \U$356 ( \480 , RI8928998_6);
and \U$357 ( \481 , \480 , \222 );
and \U$358 ( \482 , \428 , \228 );
xor \U$359 ( \483 , \481 , \482 );
and \U$360 ( \484 , \429 , \430 );
and \U$361 ( \485 , \431 , \434 );
or \U$362 ( \486 , \484 , \485 );
xor \U$363 ( \487 , \483 , \486 );
and \U$364 ( \488 , \382 , \238 );
xor \U$365 ( \489 , \487 , \488 );
and \U$366 ( \490 , \435 , \436 );
and \U$367 ( \491 , \437 , \440 );
or \U$368 ( \492 , \490 , \491 );
xor \U$369 ( \493 , \489 , \492 );
and \U$370 ( \494 , \342 , \254 );
xor \U$371 ( \495 , \493 , \494 );
and \U$372 ( \496 , \441 , \442 );
and \U$373 ( \497 , \443 , \446 );
or \U$374 ( \498 , \496 , \497 );
xor \U$375 ( \499 , \495 , \498 );
and \U$376 ( \500 , \308 , \276 );
xor \U$377 ( \501 , \499 , \500 );
and \U$378 ( \502 , \447 , \448 );
and \U$379 ( \503 , \449 , \452 );
or \U$380 ( \504 , \502 , \503 );
xor \U$381 ( \505 , \501 , \504 );
and \U$382 ( \506 , \280 , \304 );
xor \U$383 ( \507 , \505 , \506 );
and \U$384 ( \508 , \453 , \454 );
and \U$385 ( \509 , \455 , \458 );
or \U$386 ( \510 , \508 , \509 );
xor \U$387 ( \511 , \507 , \510 );
and \U$388 ( \512 , \258 , \338 );
xor \U$389 ( \513 , \511 , \512 );
and \U$390 ( \514 , \459 , \460 );
and \U$391 ( \515 , \461 , \464 );
or \U$392 ( \516 , \514 , \515 );
xor \U$393 ( \517 , \513 , \516 );
and \U$394 ( \518 , \242 , \378 );
xor \U$395 ( \519 , \517 , \518 );
and \U$396 ( \520 , \465 , \466 );
and \U$397 ( \521 , \467 , \470 );
or \U$398 ( \522 , \520 , \521 );
xor \U$399 ( \523 , \519 , \522 );
and \U$400 ( \524 , \232 , \424 );
xor \U$401 ( \525 , \523 , \524 );
and \U$402 ( \526 , \471 , \472 );
and \U$403 ( \527 , \473 , \474 );
or \U$404 ( \528 , \526 , \527 );
xor \U$405 ( \529 , \525 , \528 );
and \U$406 ( \530 , \226 , \476 );
xor \U$407 ( \531 , \529 , \530 );
and \U$408 ( \532 , \475 , \477 );
xor \U$409 ( \533 , \531 , \532 );
buf \U$410 ( \534 , RI8929118_22);
and \U$411 ( \535 , \221 , \534 );
xor \U$412 ( \536 , \533 , \535 );
buf \U$413 ( \537 , \536 );
buf \U$414 ( \538 , RI8928920_5);
and \U$415 ( \539 , \538 , \222 );
and \U$416 ( \540 , \480 , \228 );
xor \U$417 ( \541 , \539 , \540 );
and \U$418 ( \542 , \481 , \482 );
and \U$419 ( \543 , \483 , \486 );
or \U$420 ( \544 , \542 , \543 );
xor \U$421 ( \545 , \541 , \544 );
and \U$422 ( \546 , \428 , \238 );
xor \U$423 ( \547 , \545 , \546 );
and \U$424 ( \548 , \487 , \488 );
and \U$425 ( \549 , \489 , \492 );
or \U$426 ( \550 , \548 , \549 );
xor \U$427 ( \551 , \547 , \550 );
and \U$428 ( \552 , \382 , \254 );
xor \U$429 ( \553 , \551 , \552 );
and \U$430 ( \554 , \493 , \494 );
and \U$431 ( \555 , \495 , \498 );
or \U$432 ( \556 , \554 , \555 );
xor \U$433 ( \557 , \553 , \556 );
and \U$434 ( \558 , \342 , \276 );
xor \U$435 ( \559 , \557 , \558 );
and \U$436 ( \560 , \499 , \500 );
and \U$437 ( \561 , \501 , \504 );
or \U$438 ( \562 , \560 , \561 );
xor \U$439 ( \563 , \559 , \562 );
and \U$440 ( \564 , \308 , \304 );
xor \U$441 ( \565 , \563 , \564 );
and \U$442 ( \566 , \505 , \506 );
and \U$443 ( \567 , \507 , \510 );
or \U$444 ( \568 , \566 , \567 );
xor \U$445 ( \569 , \565 , \568 );
and \U$446 ( \570 , \280 , \338 );
xor \U$447 ( \571 , \569 , \570 );
and \U$448 ( \572 , \511 , \512 );
and \U$449 ( \573 , \513 , \516 );
or \U$450 ( \574 , \572 , \573 );
xor \U$451 ( \575 , \571 , \574 );
and \U$452 ( \576 , \258 , \378 );
xor \U$453 ( \577 , \575 , \576 );
and \U$454 ( \578 , \517 , \518 );
and \U$455 ( \579 , \519 , \522 );
or \U$456 ( \580 , \578 , \579 );
xor \U$457 ( \581 , \577 , \580 );
and \U$458 ( \582 , \242 , \424 );
xor \U$459 ( \583 , \581 , \582 );
and \U$460 ( \584 , \523 , \524 );
and \U$461 ( \585 , \525 , \528 );
or \U$462 ( \586 , \584 , \585 );
xor \U$463 ( \587 , \583 , \586 );
and \U$464 ( \588 , \232 , \476 );
xor \U$465 ( \589 , \587 , \588 );
and \U$466 ( \590 , \529 , \530 );
and \U$467 ( \591 , \531 , \532 );
or \U$468 ( \592 , \590 , \591 );
xor \U$469 ( \593 , \589 , \592 );
and \U$470 ( \594 , \226 , \534 );
xor \U$471 ( \595 , \593 , \594 );
and \U$472 ( \596 , \533 , \535 );
xor \U$473 ( \597 , \595 , \596 );
buf \U$474 ( \598 , RI89290a0_21);
and \U$475 ( \599 , \221 , \598 );
xor \U$476 ( \600 , \597 , \599 );
buf \U$477 ( \601 , \600 );
buf \U$478 ( \602 , RI89288a8_4);
and \U$479 ( \603 , \602 , \222 );
and \U$480 ( \604 , \538 , \228 );
xor \U$481 ( \605 , \603 , \604 );
and \U$482 ( \606 , \539 , \540 );
and \U$483 ( \607 , \541 , \544 );
or \U$484 ( \608 , \606 , \607 );
xor \U$485 ( \609 , \605 , \608 );
and \U$486 ( \610 , \480 , \238 );
xor \U$487 ( \611 , \609 , \610 );
and \U$488 ( \612 , \545 , \546 );
and \U$489 ( \613 , \547 , \550 );
or \U$490 ( \614 , \612 , \613 );
xor \U$491 ( \615 , \611 , \614 );
and \U$492 ( \616 , \428 , \254 );
xor \U$493 ( \617 , \615 , \616 );
and \U$494 ( \618 , \551 , \552 );
and \U$495 ( \619 , \553 , \556 );
or \U$496 ( \620 , \618 , \619 );
xor \U$497 ( \621 , \617 , \620 );
and \U$498 ( \622 , \382 , \276 );
xor \U$499 ( \623 , \621 , \622 );
and \U$500 ( \624 , \557 , \558 );
and \U$501 ( \625 , \559 , \562 );
or \U$502 ( \626 , \624 , \625 );
xor \U$503 ( \627 , \623 , \626 );
and \U$504 ( \628 , \342 , \304 );
xor \U$505 ( \629 , \627 , \628 );
and \U$506 ( \630 , \563 , \564 );
and \U$507 ( \631 , \565 , \568 );
or \U$508 ( \632 , \630 , \631 );
xor \U$509 ( \633 , \629 , \632 );
and \U$510 ( \634 , \308 , \338 );
xor \U$511 ( \635 , \633 , \634 );
and \U$512 ( \636 , \569 , \570 );
and \U$513 ( \637 , \571 , \574 );
or \U$514 ( \638 , \636 , \637 );
xor \U$515 ( \639 , \635 , \638 );
and \U$516 ( \640 , \280 , \378 );
xor \U$517 ( \641 , \639 , \640 );
and \U$518 ( \642 , \575 , \576 );
and \U$519 ( \643 , \577 , \580 );
or \U$520 ( \644 , \642 , \643 );
xor \U$521 ( \645 , \641 , \644 );
and \U$522 ( \646 , \258 , \424 );
xor \U$523 ( \647 , \645 , \646 );
and \U$524 ( \648 , \581 , \582 );
and \U$525 ( \649 , \583 , \586 );
or \U$526 ( \650 , \648 , \649 );
xor \U$527 ( \651 , \647 , \650 );
and \U$528 ( \652 , \242 , \476 );
xor \U$529 ( \653 , \651 , \652 );
and \U$530 ( \654 , \587 , \588 );
and \U$531 ( \655 , \589 , \592 );
or \U$532 ( \656 , \654 , \655 );
xor \U$533 ( \657 , \653 , \656 );
and \U$534 ( \658 , \232 , \534 );
xor \U$535 ( \659 , \657 , \658 );
and \U$536 ( \660 , \593 , \594 );
and \U$537 ( \661 , \595 , \596 );
or \U$538 ( \662 , \660 , \661 );
xor \U$539 ( \663 , \659 , \662 );
and \U$540 ( \664 , \226 , \598 );
xor \U$541 ( \665 , \663 , \664 );
and \U$542 ( \666 , \597 , \599 );
xor \U$543 ( \667 , \665 , \666 );
buf \U$544 ( \668 , RI8929028_20);
and \U$545 ( \669 , \221 , \668 );
xor \U$546 ( \670 , \667 , \669 );
buf \U$547 ( \671 , \670 );
buf \U$548 ( \672 , RI8928830_3);
and \U$549 ( \673 , \672 , \222 );
and \U$550 ( \674 , \602 , \228 );
xor \U$551 ( \675 , \673 , \674 );
and \U$552 ( \676 , \603 , \604 );
and \U$553 ( \677 , \605 , \608 );
or \U$554 ( \678 , \676 , \677 );
xor \U$555 ( \679 , \675 , \678 );
and \U$556 ( \680 , \538 , \238 );
xor \U$557 ( \681 , \679 , \680 );
and \U$558 ( \682 , \609 , \610 );
and \U$559 ( \683 , \611 , \614 );
or \U$560 ( \684 , \682 , \683 );
xor \U$561 ( \685 , \681 , \684 );
and \U$562 ( \686 , \480 , \254 );
xor \U$563 ( \687 , \685 , \686 );
and \U$564 ( \688 , \615 , \616 );
and \U$565 ( \689 , \617 , \620 );
or \U$566 ( \690 , \688 , \689 );
xor \U$567 ( \691 , \687 , \690 );
and \U$568 ( \692 , \428 , \276 );
xor \U$569 ( \693 , \691 , \692 );
and \U$570 ( \694 , \621 , \622 );
and \U$571 ( \695 , \623 , \626 );
or \U$572 ( \696 , \694 , \695 );
xor \U$573 ( \697 , \693 , \696 );
and \U$574 ( \698 , \382 , \304 );
xor \U$575 ( \699 , \697 , \698 );
and \U$576 ( \700 , \627 , \628 );
and \U$577 ( \701 , \629 , \632 );
or \U$578 ( \702 , \700 , \701 );
xor \U$579 ( \703 , \699 , \702 );
and \U$580 ( \704 , \342 , \338 );
xor \U$581 ( \705 , \703 , \704 );
and \U$582 ( \706 , \633 , \634 );
and \U$583 ( \707 , \635 , \638 );
or \U$584 ( \708 , \706 , \707 );
xor \U$585 ( \709 , \705 , \708 );
and \U$586 ( \710 , \308 , \378 );
xor \U$587 ( \711 , \709 , \710 );
and \U$588 ( \712 , \639 , \640 );
and \U$589 ( \713 , \641 , \644 );
or \U$590 ( \714 , \712 , \713 );
xor \U$591 ( \715 , \711 , \714 );
and \U$592 ( \716 , \280 , \424 );
xor \U$593 ( \717 , \715 , \716 );
and \U$594 ( \718 , \645 , \646 );
and \U$595 ( \719 , \647 , \650 );
or \U$596 ( \720 , \718 , \719 );
xor \U$597 ( \721 , \717 , \720 );
and \U$598 ( \722 , \258 , \476 );
xor \U$599 ( \723 , \721 , \722 );
and \U$600 ( \724 , \651 , \652 );
and \U$601 ( \725 , \653 , \656 );
or \U$602 ( \726 , \724 , \725 );
xor \U$603 ( \727 , \723 , \726 );
and \U$604 ( \728 , \242 , \534 );
xor \U$605 ( \729 , \727 , \728 );
and \U$606 ( \730 , \657 , \658 );
and \U$607 ( \731 , \659 , \662 );
or \U$608 ( \732 , \730 , \731 );
xor \U$609 ( \733 , \729 , \732 );
and \U$610 ( \734 , \232 , \598 );
xor \U$611 ( \735 , \733 , \734 );
and \U$612 ( \736 , \663 , \664 );
and \U$613 ( \737 , \665 , \666 );
or \U$614 ( \738 , \736 , \737 );
xor \U$615 ( \739 , \735 , \738 );
and \U$616 ( \740 , \226 , \668 );
xor \U$617 ( \741 , \739 , \740 );
and \U$618 ( \742 , \667 , \669 );
xor \U$619 ( \743 , \741 , \742 );
buf \U$620 ( \744 , RI8928fb0_19);
and \U$621 ( \745 , \221 , \744 );
xor \U$622 ( \746 , \743 , \745 );
buf \U$623 ( \747 , \746 );
buf \U$624 ( \748 , RI89287b8_2);
and \U$625 ( \749 , \748 , \222 );
and \U$626 ( \750 , \672 , \228 );
xor \U$627 ( \751 , \749 , \750 );
and \U$628 ( \752 , \673 , \674 );
and \U$629 ( \753 , \675 , \678 );
or \U$630 ( \754 , \752 , \753 );
xor \U$631 ( \755 , \751 , \754 );
and \U$632 ( \756 , \602 , \238 );
xor \U$633 ( \757 , \755 , \756 );
and \U$634 ( \758 , \679 , \680 );
and \U$635 ( \759 , \681 , \684 );
or \U$636 ( \760 , \758 , \759 );
xor \U$637 ( \761 , \757 , \760 );
and \U$638 ( \762 , \538 , \254 );
xor \U$639 ( \763 , \761 , \762 );
and \U$640 ( \764 , \685 , \686 );
and \U$641 ( \765 , \687 , \690 );
or \U$642 ( \766 , \764 , \765 );
xor \U$643 ( \767 , \763 , \766 );
and \U$644 ( \768 , \480 , \276 );
xor \U$645 ( \769 , \767 , \768 );
and \U$646 ( \770 , \691 , \692 );
and \U$647 ( \771 , \693 , \696 );
or \U$648 ( \772 , \770 , \771 );
xor \U$649 ( \773 , \769 , \772 );
and \U$650 ( \774 , \428 , \304 );
xor \U$651 ( \775 , \773 , \774 );
and \U$652 ( \776 , \697 , \698 );
and \U$653 ( \777 , \699 , \702 );
or \U$654 ( \778 , \776 , \777 );
xor \U$655 ( \779 , \775 , \778 );
and \U$656 ( \780 , \382 , \338 );
xor \U$657 ( \781 , \779 , \780 );
and \U$658 ( \782 , \703 , \704 );
and \U$659 ( \783 , \705 , \708 );
or \U$660 ( \784 , \782 , \783 );
xor \U$661 ( \785 , \781 , \784 );
and \U$662 ( \786 , \342 , \378 );
xor \U$663 ( \787 , \785 , \786 );
and \U$664 ( \788 , \709 , \710 );
and \U$665 ( \789 , \711 , \714 );
or \U$666 ( \790 , \788 , \789 );
xor \U$667 ( \791 , \787 , \790 );
and \U$668 ( \792 , \308 , \424 );
xor \U$669 ( \793 , \791 , \792 );
and \U$670 ( \794 , \715 , \716 );
and \U$671 ( \795 , \717 , \720 );
or \U$672 ( \796 , \794 , \795 );
xor \U$673 ( \797 , \793 , \796 );
and \U$674 ( \798 , \280 , \476 );
xor \U$675 ( \799 , \797 , \798 );
and \U$676 ( \800 , \721 , \722 );
and \U$677 ( \801 , \723 , \726 );
or \U$678 ( \802 , \800 , \801 );
xor \U$679 ( \803 , \799 , \802 );
and \U$680 ( \804 , \258 , \534 );
xor \U$681 ( \805 , \803 , \804 );
and \U$682 ( \806 , \727 , \728 );
and \U$683 ( \807 , \729 , \732 );
or \U$684 ( \808 , \806 , \807 );
xor \U$685 ( \809 , \805 , \808 );
and \U$686 ( \810 , \242 , \598 );
xor \U$687 ( \811 , \809 , \810 );
and \U$688 ( \812 , \733 , \734 );
and \U$689 ( \813 , \735 , \738 );
or \U$690 ( \814 , \812 , \813 );
xor \U$691 ( \815 , \811 , \814 );
and \U$692 ( \816 , \232 , \668 );
xor \U$693 ( \817 , \815 , \816 );
and \U$694 ( \818 , \739 , \740 );
and \U$695 ( \819 , \741 , \742 );
or \U$696 ( \820 , \818 , \819 );
xor \U$697 ( \821 , \817 , \820 );
and \U$698 ( \822 , \226 , \744 );
xor \U$699 ( \823 , \821 , \822 );
and \U$700 ( \824 , \743 , \745 );
xor \U$701 ( \825 , \823 , \824 );
buf \U$702 ( \826 , RI8928f38_18);
and \U$703 ( \827 , \221 , \826 );
xor \U$704 ( \828 , \825 , \827 );
buf \U$705 ( \829 , \828 );
buf \U$706 ( \830 , RI8928740_1);
and \U$707 ( \831 , \830 , \222 );
and \U$708 ( \832 , \748 , \228 );
xor \U$709 ( \833 , \831 , \832 );
and \U$710 ( \834 , \749 , \750 );
and \U$711 ( \835 , \751 , \754 );
or \U$712 ( \836 , \834 , \835 );
xor \U$713 ( \837 , \833 , \836 );
and \U$714 ( \838 , \672 , \238 );
xor \U$715 ( \839 , \837 , \838 );
and \U$716 ( \840 , \755 , \756 );
and \U$717 ( \841 , \757 , \760 );
or \U$718 ( \842 , \840 , \841 );
xor \U$719 ( \843 , \839 , \842 );
and \U$720 ( \844 , \602 , \254 );
xor \U$721 ( \845 , \843 , \844 );
and \U$722 ( \846 , \761 , \762 );
and \U$723 ( \847 , \763 , \766 );
or \U$724 ( \848 , \846 , \847 );
xor \U$725 ( \849 , \845 , \848 );
and \U$726 ( \850 , \538 , \276 );
xor \U$727 ( \851 , \849 , \850 );
and \U$728 ( \852 , \767 , \768 );
and \U$729 ( \853 , \769 , \772 );
or \U$730 ( \854 , \852 , \853 );
xor \U$731 ( \855 , \851 , \854 );
and \U$732 ( \856 , \480 , \304 );
xor \U$733 ( \857 , \855 , \856 );
and \U$734 ( \858 , \773 , \774 );
and \U$735 ( \859 , \775 , \778 );
or \U$736 ( \860 , \858 , \859 );
xor \U$737 ( \861 , \857 , \860 );
and \U$738 ( \862 , \428 , \338 );
xor \U$739 ( \863 , \861 , \862 );
and \U$740 ( \864 , \779 , \780 );
and \U$741 ( \865 , \781 , \784 );
or \U$742 ( \866 , \864 , \865 );
xor \U$743 ( \867 , \863 , \866 );
and \U$744 ( \868 , \382 , \378 );
xor \U$745 ( \869 , \867 , \868 );
and \U$746 ( \870 , \785 , \786 );
and \U$747 ( \871 , \787 , \790 );
or \U$748 ( \872 , \870 , \871 );
xor \U$749 ( \873 , \869 , \872 );
and \U$750 ( \874 , \342 , \424 );
xor \U$751 ( \875 , \873 , \874 );
and \U$752 ( \876 , \791 , \792 );
and \U$753 ( \877 , \793 , \796 );
or \U$754 ( \878 , \876 , \877 );
xor \U$755 ( \879 , \875 , \878 );
and \U$756 ( \880 , \308 , \476 );
xor \U$757 ( \881 , \879 , \880 );
and \U$758 ( \882 , \797 , \798 );
and \U$759 ( \883 , \799 , \802 );
or \U$760 ( \884 , \882 , \883 );
xor \U$761 ( \885 , \881 , \884 );
and \U$762 ( \886 , \280 , \534 );
xor \U$763 ( \887 , \885 , \886 );
and \U$764 ( \888 , \803 , \804 );
and \U$765 ( \889 , \805 , \808 );
or \U$766 ( \890 , \888 , \889 );
xor \U$767 ( \891 , \887 , \890 );
and \U$768 ( \892 , \258 , \598 );
xor \U$769 ( \893 , \891 , \892 );
and \U$770 ( \894 , \809 , \810 );
and \U$771 ( \895 , \811 , \814 );
or \U$772 ( \896 , \894 , \895 );
xor \U$773 ( \897 , \893 , \896 );
and \U$774 ( \898 , \242 , \668 );
xor \U$775 ( \899 , \897 , \898 );
and \U$776 ( \900 , \815 , \816 );
and \U$777 ( \901 , \817 , \820 );
or \U$778 ( \902 , \900 , \901 );
xor \U$779 ( \903 , \899 , \902 );
and \U$780 ( \904 , \232 , \744 );
xor \U$781 ( \905 , \903 , \904 );
and \U$782 ( \906 , \821 , \822 );
and \U$783 ( \907 , \823 , \824 );
or \U$784 ( \908 , \906 , \907 );
xor \U$785 ( \909 , \905 , \908 );
and \U$786 ( \910 , \226 , \826 );
xor \U$787 ( \911 , \909 , \910 );
and \U$788 ( \912 , \825 , \827 );
xor \U$789 ( \913 , \911 , \912 );
buf \U$790 ( \914 , RI8928ec0_17);
and \U$791 ( \915 , \221 , \914 );
xor \U$792 ( \916 , \913 , \915 );
buf \U$793 ( \917 , \916 );
nor \U$794 ( \918 , \225 , \231 , \241 , \257 , \279 , \307 , \341 , \381 , \427 , \479 , \537 , \601 , \671 , \747 , \829 , \917 );
not \U$795 ( \919 , \231 );
nor \U$796 ( \920 , \224 , \919 , \241 , \257 , \279 , \307 , \341 , \381 , \427 , \479 , \537 , \601 , \671 , \747 , \829 , \917 );
not \U$797 ( \921 , \241 );
nor \U$798 ( \922 , \224 , \231 , \921 , \257 , \279 , \307 , \341 , \381 , \427 , \479 , \537 , \601 , \671 , \747 , \829 , \917 );
not \U$799 ( \923 , \257 );
nor \U$800 ( \924 , \224 , \231 , \241 , \923 , \279 , \307 , \341 , \381 , \427 , \479 , \537 , \601 , \671 , \747 , \829 , \917 );
not \U$801 ( \925 , \279 );
nor \U$802 ( \926 , \224 , \231 , \241 , \257 , \925 , \307 , \341 , \381 , \427 , \479 , \537 , \601 , \671 , \747 , \829 , \917 );
not \U$803 ( \927 , \307 );
nor \U$804 ( \928 , \224 , \231 , \241 , \257 , \279 , \927 , \341 , \381 , \427 , \479 , \537 , \601 , \671 , \747 , \829 , \917 );
not \U$805 ( \929 , \341 );
nor \U$806 ( \930 , \224 , \231 , \241 , \257 , \279 , \307 , \929 , \381 , \427 , \479 , \537 , \601 , \671 , \747 , \829 , \917 );
not \U$807 ( \931 , \381 );
nor \U$808 ( \932 , \224 , \231 , \241 , \257 , \279 , \307 , \341 , \931 , \427 , \479 , \537 , \601 , \671 , \747 , \829 , \917 );
not \U$809 ( \933 , \427 );
nor \U$810 ( \934 , \224 , \231 , \241 , \257 , \279 , \307 , \341 , \381 , \933 , \479 , \537 , \601 , \671 , \747 , \829 , \917 );
not \U$811 ( \935 , \479 );
nor \U$812 ( \936 , \224 , \231 , \241 , \257 , \279 , \307 , \341 , \381 , \427 , \935 , \537 , \601 , \671 , \747 , \829 , \917 );
not \U$813 ( \937 , \537 );
nor \U$814 ( \938 , \224 , \231 , \241 , \257 , \279 , \307 , \341 , \381 , \427 , \479 , \937 , \601 , \671 , \747 , \829 , \917 );
not \U$815 ( \939 , \601 );
nor \U$816 ( \940 , \224 , \231 , \241 , \257 , \279 , \307 , \341 , \381 , \427 , \479 , \537 , \939 , \671 , \747 , \829 , \917 );
nor \U$817 ( \941 , \918 , \920 , \922 , \924 , \926 , \928 , \930 , \932 , \934 , \936 , \938 , \940 );
_DC g3a2 ( \942_nG3a2 , 1'b0 , \941 );
or \U$818 ( \943 , RI8928dd0_15, RI892a450_63);
and \U$819 ( \944 , \943 , \940 );
and \U$820 ( \945 , RI8929550_31, RI8929cd0_47);
and \U$821 ( \946 , \945 , \938 );
or \U$822 ( \947 , RI8928dd0_15, RI8929550_31);
and \U$823 ( \948 , \947 , \936 );
xor \U$824 ( \949 , RI8929cd0_47, RI892a450_63);
and \U$825 ( \950 , \949 , \934 );
buf \U$826 ( \951 , RI8929550_31);
buf \U$827 ( \952 , RI8929d48_48);
and \U$828 ( \953 , \951 , \952 );
buf \U$829 ( \954 , RI89295c8_32);
buf \U$830 ( \955 , RI8929cd0_47);
and \U$831 ( \956 , \954 , \955 );
xor \U$832 ( \957 , \953 , \956 );
buf \U$833 ( \958 , \957 );
and \U$834 ( \959 , \958 , \932 );
buf \U$835 ( \960 , RI8928dd0_15);
buf \U$836 ( \961 , RI892a4c8_64);
and \U$837 ( \962 , \960 , \961 );
buf \U$838 ( \963 , RI8928e48_16);
buf \U$839 ( \964 , RI892a450_63);
and \U$840 ( \965 , \963 , \964 );
xor \U$841 ( \966 , \962 , \965 );
buf \U$842 ( \967 , \966 );
and \U$843 ( \968 , \967 , \930 );
buf \U$844 ( \969 , RI8929550_31);
buf \U$845 ( \970 , RI892a450_63);
xor \U$846 ( \971 , \969 , \970 );
buf \U$847 ( \972 , RI89295c8_32);
buf \U$848 ( \973 , RI892a4c8_64);
and \U$849 ( \974 , \972 , \973 );
xor \U$850 ( \975 , \971 , \974 );
buf \U$851 ( \976 , \975 );
and \U$852 ( \977 , \976 , \928 );
buf \U$853 ( \978 , RI8928dd0_15);
buf \U$854 ( \979 , RI8929cd0_47);
xor \U$855 ( \980 , \978 , \979 );
buf \U$856 ( \981 , RI8928e48_16);
buf \U$857 ( \982 , RI8929d48_48);
and \U$858 ( \983 , \981 , \982 );
xor \U$859 ( \984 , \980 , \983 );
buf \U$860 ( \985 , \984 );
and \U$861 ( \986 , \985 , \926 );
and \U$862 ( \987 , RI892a450_63, \924 );
and \U$863 ( \988 , RI8929cd0_47, \922 );
and \U$864 ( \989 , RI8929550_31, \920 );
and \U$865 ( \990 , RI8928dd0_15, \918 );
or \U$866 ( \991 , \942_nG3a2 , \944 , \946 , \948 , \950 , \959 , \968 , \977 , \986 , \987 , \988 , \989 , \990 );
buf \U$867 ( \992 , \991 );
and \U$868 ( \993 , \220 , \992 );
_DC g3d6 ( \994_nG3d6 , 1'b0 , \941 );
or \U$870 ( \995 , RI8928e48_16, RI892a4c8_64);
and \U$871 ( \996 , \995 , \940 );
and \U$872 ( \997 , RI89295c8_32, RI8929d48_48);
and \U$873 ( \998 , \997 , \938 );
or \U$874 ( \999 , RI8928e48_16, RI89295c8_32);
and \U$875 ( \1000 , \999 , \936 );
xor \U$876 ( \1001 , RI8929d48_48, RI892a4c8_64);
and \U$877 ( \1002 , \1001 , \934 );
and \U$878 ( \1003 , \954 , \952 );
buf \U$879 ( \1004 , \1003 );
and \U$880 ( \1005 , \1004 , \932 );
and \U$881 ( \1006 , \963 , \961 );
buf \U$882 ( \1007 , \1006 );
and \U$883 ( \1008 , \1007 , \930 );
xor \U$884 ( \1009 , \972 , \973 );
buf \U$885 ( \1010 , \1009 );
and \U$886 ( \1011 , \1010 , \928 );
xor \U$887 ( \1012 , \981 , \982 );
buf \U$888 ( \1013 , \1012 );
and \U$889 ( \1014 , \1013 , \926 );
and \U$890 ( \1015 , RI892a4c8_64, \924 );
and \U$891 ( \1016 , RI8929d48_48, \922 );
and \U$892 ( \1017 , RI89295c8_32, \920 );
and \U$893 ( \1018 , RI8928e48_16, \918 );
or \U$894 ( \1019 , \994_nG3d6 , \996 , \998 , \1000 , \1002 , \1005 , \1008 , \1011 , \1014 , \1015 , \1016 , \1017 , \1018 );
buf \U$895 ( \1020 , \1019 );
and \U$896 ( \1021 , \220 , \1020 );
xor \U$897 ( \1022 , \126 , \127 );
xor \U$898 ( \1023 , \1022 , \215 );
buf \U$899 ( \1024 , \1023 );
buf \U$900 ( \1025 , \1024 );
and \U$901 ( \1026 , \1025 , \992 );
and \U$902 ( \1027 , \1021 , \1026 );
xor \U$903 ( \1028 , \1021 , \1026 );
and \U$904 ( \1029 , \1025 , \1020 );
xor \U$905 ( \1030 , \129 , \130 );
xor \U$906 ( \1031 , \1030 , \212 );
buf \U$907 ( \1032 , \1031 );
buf \U$908 ( \1033 , \1032 );
and \U$909 ( \1034 , \1033 , \992 );
and \U$910 ( \1035 , \1029 , \1034 );
xor \U$911 ( \1036 , \1029 , \1034 );
and \U$912 ( \1037 , \1033 , \1020 );
xor \U$913 ( \1038 , \132 , \133 );
xor \U$914 ( \1039 , \1038 , \209 );
buf \U$915 ( \1040 , \1039 );
buf \U$916 ( \1041 , \1040 );
and \U$917 ( \1042 , \1041 , \992 );
and \U$918 ( \1043 , \1037 , \1042 );
xor \U$919 ( \1044 , \1037 , \1042 );
and \U$920 ( \1045 , \1041 , \1020 );
xor \U$921 ( \1046 , \135 , \136 );
xor \U$922 ( \1047 , \1046 , \206 );
buf \U$923 ( \1048 , \1047 );
buf \U$924 ( \1049 , \1048 );
and \U$925 ( \1050 , \1049 , \992 );
and \U$926 ( \1051 , \1045 , \1050 );
xor \U$927 ( \1052 , \1045 , \1050 );
and \U$928 ( \1053 , \1049 , \1020 );
xor \U$929 ( \1054 , \138 , \139 );
xor \U$930 ( \1055 , \1054 , \203 );
buf \U$931 ( \1056 , \1055 );
buf \U$932 ( \1057 , \1056 );
and \U$933 ( \1058 , \1057 , \992 );
and \U$934 ( \1059 , \1053 , \1058 );
xor \U$935 ( \1060 , \1053 , \1058 );
and \U$936 ( \1061 , \1057 , \1020 );
xor \U$937 ( \1062 , \141 , \142 );
xor \U$938 ( \1063 , \1062 , \200 );
buf \U$939 ( \1064 , \1063 );
buf \U$940 ( \1065 , \1064 );
and \U$941 ( \1066 , \1065 , \992 );
and \U$942 ( \1067 , \1061 , \1066 );
xor \U$943 ( \1068 , \1061 , \1066 );
and \U$944 ( \1069 , \1065 , \1020 );
xor \U$945 ( \1070 , \144 , \145 );
xor \U$946 ( \1071 , \1070 , \197 );
buf \U$947 ( \1072 , \1071 );
buf \U$948 ( \1073 , \1072 );
and \U$949 ( \1074 , \1073 , \992 );
and \U$950 ( \1075 , \1069 , \1074 );
xor \U$951 ( \1076 , \1069 , \1074 );
and \U$952 ( \1077 , \1073 , \1020 );
xor \U$953 ( \1078 , \147 , \148 );
xor \U$954 ( \1079 , \1078 , \194 );
buf \U$955 ( \1080 , \1079 );
buf \U$956 ( \1081 , \1080 );
and \U$957 ( \1082 , \1081 , \992 );
and \U$958 ( \1083 , \1077 , \1082 );
xor \U$959 ( \1084 , \1077 , \1082 );
and \U$960 ( \1085 , \1081 , \1020 );
xor \U$961 ( \1086 , \150 , \151 );
xor \U$962 ( \1087 , \1086 , \191 );
buf \U$963 ( \1088 , \1087 );
buf \U$964 ( \1089 , \1088 );
and \U$965 ( \1090 , \1089 , \992 );
and \U$966 ( \1091 , \1085 , \1090 );
xor \U$967 ( \1092 , \1085 , \1090 );
and \U$968 ( \1093 , \1089 , \1020 );
xor \U$969 ( \1094 , \153 , \154 );
xor \U$970 ( \1095 , \1094 , \188 );
buf \U$971 ( \1096 , \1095 );
buf \U$972 ( \1097 , \1096 );
and \U$973 ( \1098 , \1097 , \992 );
and \U$974 ( \1099 , \1093 , \1098 );
xor \U$975 ( \1100 , \1093 , \1098 );
and \U$976 ( \1101 , \1097 , \1020 );
xor \U$977 ( \1102 , \156 , \157 );
xor \U$978 ( \1103 , \1102 , \185 );
buf \U$979 ( \1104 , \1103 );
buf \U$980 ( \1105 , \1104 );
and \U$981 ( \1106 , \1105 , \992 );
and \U$982 ( \1107 , \1101 , \1106 );
xor \U$983 ( \1108 , \1101 , \1106 );
and \U$984 ( \1109 , \1105 , \1020 );
xor \U$985 ( \1110 , \159 , \160 );
xor \U$986 ( \1111 , \1110 , \182 );
buf \U$987 ( \1112 , \1111 );
buf \U$988 ( \1113 , \1112 );
and \U$989 ( \1114 , \1113 , \992 );
and \U$990 ( \1115 , \1109 , \1114 );
xor \U$991 ( \1116 , \1109 , \1114 );
and \U$992 ( \1117 , \1113 , \1020 );
xor \U$993 ( \1118 , \162 , \163 );
xor \U$994 ( \1119 , \1118 , \179 );
buf \U$995 ( \1120 , \1119 );
buf \U$996 ( \1121 , \1120 );
and \U$997 ( \1122 , \1121 , \992 );
and \U$998 ( \1123 , \1117 , \1122 );
xor \U$999 ( \1124 , \1117 , \1122 );
and \U$1000 ( \1125 , \1121 , \1020 );
xor \U$1001 ( \1126 , \165 , \166 );
xor \U$1002 ( \1127 , \1126 , \176 );
buf \U$1003 ( \1128 , \1127 );
buf \U$1004 ( \1129 , \1128 );
and \U$1005 ( \1130 , \1129 , \992 );
and \U$1006 ( \1131 , \1125 , \1130 );
xor \U$1007 ( \1132 , \1125 , \1130 );
and \U$1008 ( \1133 , \1129 , \1020 );
xor \U$1009 ( \1134 , \168 , \169 );
xor \U$1010 ( \1135 , \1134 , \173 );
buf \U$1011 ( \1136 , \1135 );
buf \U$1012 ( \1137 , \1136 );
and \U$1013 ( \1138 , \1137 , \992 );
and \U$1014 ( \1139 , \1133 , \1138 );
xor \U$1015 ( \1140 , \1133 , \1138 );
and \U$1016 ( \1141 , \1137 , \1020 );
xor \U$1017 ( \1142 , \171 , \172 );
buf \U$1018 ( \1143 , \1142 );
buf \U$1019 ( \1144 , \1143 );
and \U$1020 ( \1145 , \1144 , \992 );
and \U$1021 ( \1146 , \1141 , \1145 );
and \U$1022 ( \1147 , \1140 , \1146 );
or \U$1023 ( \1148 , \1139 , \1147 );
and \U$1024 ( \1149 , \1132 , \1148 );
or \U$1025 ( \1150 , \1131 , \1149 );
and \U$1026 ( \1151 , \1124 , \1150 );
or \U$1027 ( \1152 , \1123 , \1151 );
and \U$1028 ( \1153 , \1116 , \1152 );
or \U$1029 ( \1154 , \1115 , \1153 );
and \U$1030 ( \1155 , \1108 , \1154 );
or \U$1031 ( \1156 , \1107 , \1155 );
and \U$1032 ( \1157 , \1100 , \1156 );
or \U$1033 ( \1158 , \1099 , \1157 );
and \U$1034 ( \1159 , \1092 , \1158 );
or \U$1035 ( \1160 , \1091 , \1159 );
and \U$1036 ( \1161 , \1084 , \1160 );
or \U$1037 ( \1162 , \1083 , \1161 );
and \U$1038 ( \1163 , \1076 , \1162 );
or \U$1039 ( \1164 , \1075 , \1163 );
and \U$1040 ( \1165 , \1068 , \1164 );
or \U$1041 ( \1166 , \1067 , \1165 );
and \U$1042 ( \1167 , \1060 , \1166 );
or \U$1043 ( \1168 , \1059 , \1167 );
and \U$1044 ( \1169 , \1052 , \1168 );
or \U$1045 ( \1170 , \1051 , \1169 );
and \U$1046 ( \1171 , \1044 , \1170 );
or \U$1047 ( \1172 , \1043 , \1171 );
and \U$1048 ( \1173 , \1036 , \1172 );
or \U$1049 ( \1174 , \1035 , \1173 );
and \U$1050 ( \1175 , \1028 , \1174 );
or \U$1051 ( \1176 , \1027 , \1175 );
and \U$1052 ( \1177 , \993 , \1176 );
_DC g48e ( \1178_nG48e , 1'b0 , \941 );
or \U$1054 ( \1179 , RI8928d58_14, RI892a3d8_62);
and \U$1055 ( \1180 , \1179 , \940 );
and \U$1056 ( \1181 , RI89294d8_30, RI8929c58_46);
and \U$1057 ( \1182 , \1181 , \938 );
or \U$1058 ( \1183 , RI8928d58_14, RI89294d8_30);
and \U$1059 ( \1184 , \1183 , \936 );
xor \U$1060 ( \1185 , RI8929c58_46, RI892a3d8_62);
and \U$1061 ( \1186 , \1185 , \934 );
buf \U$1062 ( \1187 , RI89294d8_30);
and \U$1063 ( \1188 , \1187 , \952 );
and \U$1064 ( \1189 , \951 , \955 );
xor \U$1065 ( \1190 , \1188 , \1189 );
and \U$1066 ( \1191 , \953 , \956 );
xor \U$1067 ( \1192 , \1190 , \1191 );
buf \U$1068 ( \1193 , RI8929c58_46);
and \U$1069 ( \1194 , \954 , \1193 );
xor \U$1070 ( \1195 , \1192 , \1194 );
buf \U$1071 ( \1196 , \1195 );
and \U$1072 ( \1197 , \1196 , \932 );
buf \U$1073 ( \1198 , RI8928d58_14);
and \U$1074 ( \1199 , \1198 , \961 );
and \U$1075 ( \1200 , \960 , \964 );
xor \U$1076 ( \1201 , \1199 , \1200 );
and \U$1077 ( \1202 , \962 , \965 );
xor \U$1078 ( \1203 , \1201 , \1202 );
buf \U$1079 ( \1204 , RI892a3d8_62);
and \U$1080 ( \1205 , \963 , \1204 );
xor \U$1081 ( \1206 , \1203 , \1205 );
buf \U$1082 ( \1207 , \1206 );
and \U$1083 ( \1208 , \1207 , \930 );
buf \U$1084 ( \1209 , RI89294d8_30);
buf \U$1085 ( \1210 , RI892a3d8_62);
xor \U$1086 ( \1211 , \1209 , \1210 );
and \U$1087 ( \1212 , \969 , \970 );
and \U$1088 ( \1213 , \970 , \974 );
and \U$1089 ( \1214 , \969 , \974 );
or \U$1090 ( \1215 , \1212 , \1213 , \1214 );
xor \U$1091 ( \1216 , \1211 , \1215 );
buf \U$1092 ( \1217 , \1216 );
and \U$1093 ( \1218 , \1217 , \928 );
buf \U$1094 ( \1219 , RI8928d58_14);
buf \U$1095 ( \1220 , RI8929c58_46);
xor \U$1096 ( \1221 , \1219 , \1220 );
and \U$1097 ( \1222 , \978 , \979 );
and \U$1098 ( \1223 , \979 , \983 );
and \U$1099 ( \1224 , \978 , \983 );
or \U$1100 ( \1225 , \1222 , \1223 , \1224 );
xor \U$1101 ( \1226 , \1221 , \1225 );
buf \U$1102 ( \1227 , \1226 );
and \U$1103 ( \1228 , \1227 , \926 );
and \U$1104 ( \1229 , RI892a3d8_62, \924 );
and \U$1105 ( \1230 , RI8929c58_46, \922 );
and \U$1106 ( \1231 , RI89294d8_30, \920 );
and \U$1107 ( \1232 , RI8928d58_14, \918 );
or \U$1108 ( \1233 , \1178_nG48e , \1180 , \1182 , \1184 , \1186 , \1197 , \1208 , \1218 , \1228 , \1229 , \1230 , \1231 , \1232 );
buf \U$1109 ( \1234 , \1233 );
and \U$1110 ( \1235 , \220 , \1234 );
and \U$1111 ( \1236 , \1177 , \1235 );
xor \U$1112 ( \1237 , \1177 , \1235 );
xor \U$1113 ( \1238 , \993 , \1176 );
and \U$1114 ( \1239 , \1025 , \1234 );
and \U$1115 ( \1240 , \1238 , \1239 );
xor \U$1116 ( \1241 , \1238 , \1239 );
xor \U$1117 ( \1242 , \1028 , \1174 );
and \U$1118 ( \1243 , \1033 , \1234 );
and \U$1119 ( \1244 , \1242 , \1243 );
xor \U$1120 ( \1245 , \1242 , \1243 );
xor \U$1121 ( \1246 , \1036 , \1172 );
and \U$1122 ( \1247 , \1041 , \1234 );
and \U$1123 ( \1248 , \1246 , \1247 );
xor \U$1124 ( \1249 , \1246 , \1247 );
xor \U$1125 ( \1250 , \1044 , \1170 );
and \U$1126 ( \1251 , \1049 , \1234 );
and \U$1127 ( \1252 , \1250 , \1251 );
xor \U$1128 ( \1253 , \1250 , \1251 );
xor \U$1129 ( \1254 , \1052 , \1168 );
and \U$1130 ( \1255 , \1057 , \1234 );
and \U$1131 ( \1256 , \1254 , \1255 );
xor \U$1132 ( \1257 , \1254 , \1255 );
xor \U$1133 ( \1258 , \1060 , \1166 );
and \U$1134 ( \1259 , \1065 , \1234 );
and \U$1135 ( \1260 , \1258 , \1259 );
xor \U$1136 ( \1261 , \1258 , \1259 );
xor \U$1137 ( \1262 , \1068 , \1164 );
and \U$1138 ( \1263 , \1073 , \1234 );
and \U$1139 ( \1264 , \1262 , \1263 );
xor \U$1140 ( \1265 , \1262 , \1263 );
xor \U$1141 ( \1266 , \1076 , \1162 );
and \U$1142 ( \1267 , \1081 , \1234 );
and \U$1143 ( \1268 , \1266 , \1267 );
xor \U$1144 ( \1269 , \1266 , \1267 );
xor \U$1145 ( \1270 , \1084 , \1160 );
and \U$1146 ( \1271 , \1089 , \1234 );
and \U$1147 ( \1272 , \1270 , \1271 );
xor \U$1148 ( \1273 , \1270 , \1271 );
xor \U$1149 ( \1274 , \1092 , \1158 );
and \U$1150 ( \1275 , \1097 , \1234 );
and \U$1151 ( \1276 , \1274 , \1275 );
xor \U$1152 ( \1277 , \1274 , \1275 );
xor \U$1153 ( \1278 , \1100 , \1156 );
and \U$1154 ( \1279 , \1105 , \1234 );
and \U$1155 ( \1280 , \1278 , \1279 );
xor \U$1156 ( \1281 , \1278 , \1279 );
xor \U$1157 ( \1282 , \1108 , \1154 );
and \U$1158 ( \1283 , \1113 , \1234 );
and \U$1159 ( \1284 , \1282 , \1283 );
xor \U$1160 ( \1285 , \1282 , \1283 );
xor \U$1161 ( \1286 , \1116 , \1152 );
and \U$1162 ( \1287 , \1121 , \1234 );
and \U$1163 ( \1288 , \1286 , \1287 );
xor \U$1164 ( \1289 , \1286 , \1287 );
xor \U$1165 ( \1290 , \1124 , \1150 );
and \U$1166 ( \1291 , \1129 , \1234 );
and \U$1167 ( \1292 , \1290 , \1291 );
xor \U$1168 ( \1293 , \1290 , \1291 );
xor \U$1169 ( \1294 , \1132 , \1148 );
and \U$1170 ( \1295 , \1137 , \1234 );
and \U$1171 ( \1296 , \1294 , \1295 );
xor \U$1172 ( \1297 , \1294 , \1295 );
xor \U$1173 ( \1298 , \1140 , \1146 );
and \U$1174 ( \1299 , \1144 , \1234 );
and \U$1175 ( \1300 , \1298 , \1299 );
and \U$1176 ( \1301 , \1297 , \1300 );
or \U$1177 ( \1302 , \1296 , \1301 );
and \U$1178 ( \1303 , \1293 , \1302 );
or \U$1179 ( \1304 , \1292 , \1303 );
and \U$1180 ( \1305 , \1289 , \1304 );
or \U$1181 ( \1306 , \1288 , \1305 );
and \U$1182 ( \1307 , \1285 , \1306 );
or \U$1183 ( \1308 , \1284 , \1307 );
and \U$1184 ( \1309 , \1281 , \1308 );
or \U$1185 ( \1310 , \1280 , \1309 );
and \U$1186 ( \1311 , \1277 , \1310 );
or \U$1187 ( \1312 , \1276 , \1311 );
and \U$1188 ( \1313 , \1273 , \1312 );
or \U$1189 ( \1314 , \1272 , \1313 );
and \U$1190 ( \1315 , \1269 , \1314 );
or \U$1191 ( \1316 , \1268 , \1315 );
and \U$1192 ( \1317 , \1265 , \1316 );
or \U$1193 ( \1318 , \1264 , \1317 );
and \U$1194 ( \1319 , \1261 , \1318 );
or \U$1195 ( \1320 , \1260 , \1319 );
and \U$1196 ( \1321 , \1257 , \1320 );
or \U$1197 ( \1322 , \1256 , \1321 );
and \U$1198 ( \1323 , \1253 , \1322 );
or \U$1199 ( \1324 , \1252 , \1323 );
and \U$1200 ( \1325 , \1249 , \1324 );
or \U$1201 ( \1326 , \1248 , \1325 );
and \U$1202 ( \1327 , \1245 , \1326 );
or \U$1203 ( \1328 , \1244 , \1327 );
and \U$1204 ( \1329 , \1241 , \1328 );
or \U$1205 ( \1330 , \1240 , \1329 );
and \U$1206 ( \1331 , \1237 , \1330 );
or \U$1207 ( \1332 , \1236 , \1331 );
_DC g529 ( \1333_nG529 , 1'b0 , \941 );
or \U$1209 ( \1334 , RI8928ce0_13, RI892a360_61);
and \U$1210 ( \1335 , \1334 , \940 );
and \U$1211 ( \1336 , RI8929460_29, RI8929be0_45);
and \U$1212 ( \1337 , \1336 , \938 );
or \U$1213 ( \1338 , RI8928ce0_13, RI8929460_29);
and \U$1214 ( \1339 , \1338 , \936 );
xor \U$1215 ( \1340 , RI8929be0_45, RI892a360_61);
and \U$1216 ( \1341 , \1340 , \934 );
buf \U$1217 ( \1342 , RI8929460_29);
and \U$1218 ( \1343 , \1342 , \952 );
and \U$1219 ( \1344 , \1187 , \955 );
xor \U$1220 ( \1345 , \1343 , \1344 );
and \U$1221 ( \1346 , \1188 , \1189 );
and \U$1222 ( \1347 , \1190 , \1191 );
or \U$1223 ( \1348 , \1346 , \1347 );
xor \U$1224 ( \1349 , \1345 , \1348 );
and \U$1225 ( \1350 , \951 , \1193 );
xor \U$1226 ( \1351 , \1349 , \1350 );
and \U$1227 ( \1352 , \1192 , \1194 );
xor \U$1228 ( \1353 , \1351 , \1352 );
buf \U$1229 ( \1354 , RI8929be0_45);
and \U$1230 ( \1355 , \954 , \1354 );
xor \U$1231 ( \1356 , \1353 , \1355 );
buf \U$1232 ( \1357 , \1356 );
and \U$1233 ( \1358 , \1357 , \932 );
buf \U$1234 ( \1359 , RI8928ce0_13);
and \U$1235 ( \1360 , \1359 , \961 );
and \U$1236 ( \1361 , \1198 , \964 );
xor \U$1237 ( \1362 , \1360 , \1361 );
and \U$1238 ( \1363 , \1199 , \1200 );
and \U$1239 ( \1364 , \1201 , \1202 );
or \U$1240 ( \1365 , \1363 , \1364 );
xor \U$1241 ( \1366 , \1362 , \1365 );
and \U$1242 ( \1367 , \960 , \1204 );
xor \U$1243 ( \1368 , \1366 , \1367 );
and \U$1244 ( \1369 , \1203 , \1205 );
xor \U$1245 ( \1370 , \1368 , \1369 );
buf \U$1246 ( \1371 , RI892a360_61);
and \U$1247 ( \1372 , \963 , \1371 );
xor \U$1248 ( \1373 , \1370 , \1372 );
buf \U$1249 ( \1374 , \1373 );
and \U$1250 ( \1375 , \1374 , \930 );
buf \U$1251 ( \1376 , RI8929460_29);
buf \U$1252 ( \1377 , RI892a360_61);
xor \U$1253 ( \1378 , \1376 , \1377 );
and \U$1254 ( \1379 , \1209 , \1210 );
and \U$1255 ( \1380 , \1210 , \1215 );
and \U$1256 ( \1381 , \1209 , \1215 );
or \U$1257 ( \1382 , \1379 , \1380 , \1381 );
xor \U$1258 ( \1383 , \1378 , \1382 );
buf \U$1259 ( \1384 , \1383 );
and \U$1260 ( \1385 , \1384 , \928 );
buf \U$1261 ( \1386 , RI8928ce0_13);
buf \U$1262 ( \1387 , RI8929be0_45);
xor \U$1263 ( \1388 , \1386 , \1387 );
and \U$1264 ( \1389 , \1219 , \1220 );
and \U$1265 ( \1390 , \1220 , \1225 );
and \U$1266 ( \1391 , \1219 , \1225 );
or \U$1267 ( \1392 , \1389 , \1390 , \1391 );
xor \U$1268 ( \1393 , \1388 , \1392 );
buf \U$1269 ( \1394 , \1393 );
and \U$1270 ( \1395 , \1394 , \926 );
and \U$1271 ( \1396 , RI892a360_61, \924 );
and \U$1272 ( \1397 , RI8929be0_45, \922 );
and \U$1273 ( \1398 , RI8929460_29, \920 );
and \U$1274 ( \1399 , RI8928ce0_13, \918 );
or \U$1275 ( \1400 , \1333_nG529 , \1335 , \1337 , \1339 , \1341 , \1358 , \1375 , \1385 , \1395 , \1396 , \1397 , \1398 , \1399 );
buf \U$1276 ( \1401 , \1400 );
and \U$1277 ( \1402 , \220 , \1401 );
and \U$1278 ( \1403 , \1332 , \1402 );
xor \U$1279 ( \1404 , \1332 , \1402 );
xor \U$1280 ( \1405 , \1237 , \1330 );
and \U$1281 ( \1406 , \1025 , \1401 );
and \U$1282 ( \1407 , \1405 , \1406 );
xor \U$1283 ( \1408 , \1405 , \1406 );
xor \U$1284 ( \1409 , \1241 , \1328 );
and \U$1285 ( \1410 , \1033 , \1401 );
and \U$1286 ( \1411 , \1409 , \1410 );
xor \U$1287 ( \1412 , \1409 , \1410 );
xor \U$1288 ( \1413 , \1245 , \1326 );
and \U$1289 ( \1414 , \1041 , \1401 );
and \U$1290 ( \1415 , \1413 , \1414 );
xor \U$1291 ( \1416 , \1413 , \1414 );
xor \U$1292 ( \1417 , \1249 , \1324 );
and \U$1293 ( \1418 , \1049 , \1401 );
and \U$1294 ( \1419 , \1417 , \1418 );
xor \U$1295 ( \1420 , \1417 , \1418 );
xor \U$1296 ( \1421 , \1253 , \1322 );
and \U$1297 ( \1422 , \1057 , \1401 );
and \U$1298 ( \1423 , \1421 , \1422 );
xor \U$1299 ( \1424 , \1421 , \1422 );
xor \U$1300 ( \1425 , \1257 , \1320 );
and \U$1301 ( \1426 , \1065 , \1401 );
and \U$1302 ( \1427 , \1425 , \1426 );
xor \U$1303 ( \1428 , \1425 , \1426 );
xor \U$1304 ( \1429 , \1261 , \1318 );
and \U$1305 ( \1430 , \1073 , \1401 );
and \U$1306 ( \1431 , \1429 , \1430 );
xor \U$1307 ( \1432 , \1429 , \1430 );
xor \U$1308 ( \1433 , \1265 , \1316 );
and \U$1309 ( \1434 , \1081 , \1401 );
and \U$1310 ( \1435 , \1433 , \1434 );
xor \U$1311 ( \1436 , \1433 , \1434 );
xor \U$1312 ( \1437 , \1269 , \1314 );
and \U$1313 ( \1438 , \1089 , \1401 );
and \U$1314 ( \1439 , \1437 , \1438 );
xor \U$1315 ( \1440 , \1437 , \1438 );
xor \U$1316 ( \1441 , \1273 , \1312 );
and \U$1317 ( \1442 , \1097 , \1401 );
and \U$1318 ( \1443 , \1441 , \1442 );
xor \U$1319 ( \1444 , \1441 , \1442 );
xor \U$1320 ( \1445 , \1277 , \1310 );
and \U$1321 ( \1446 , \1105 , \1401 );
and \U$1322 ( \1447 , \1445 , \1446 );
xor \U$1323 ( \1448 , \1445 , \1446 );
xor \U$1324 ( \1449 , \1281 , \1308 );
and \U$1325 ( \1450 , \1113 , \1401 );
and \U$1326 ( \1451 , \1449 , \1450 );
xor \U$1327 ( \1452 , \1449 , \1450 );
xor \U$1328 ( \1453 , \1285 , \1306 );
and \U$1329 ( \1454 , \1121 , \1401 );
and \U$1330 ( \1455 , \1453 , \1454 );
xor \U$1331 ( \1456 , \1453 , \1454 );
xor \U$1332 ( \1457 , \1289 , \1304 );
and \U$1333 ( \1458 , \1129 , \1401 );
and \U$1334 ( \1459 , \1457 , \1458 );
xor \U$1335 ( \1460 , \1457 , \1458 );
xor \U$1336 ( \1461 , \1293 , \1302 );
and \U$1337 ( \1462 , \1137 , \1401 );
and \U$1338 ( \1463 , \1461 , \1462 );
xor \U$1339 ( \1464 , \1461 , \1462 );
xor \U$1340 ( \1465 , \1297 , \1300 );
and \U$1341 ( \1466 , \1144 , \1401 );
and \U$1342 ( \1467 , \1465 , \1466 );
and \U$1343 ( \1468 , \1464 , \1467 );
or \U$1344 ( \1469 , \1463 , \1468 );
and \U$1345 ( \1470 , \1460 , \1469 );
or \U$1346 ( \1471 , \1459 , \1470 );
and \U$1347 ( \1472 , \1456 , \1471 );
or \U$1348 ( \1473 , \1455 , \1472 );
and \U$1349 ( \1474 , \1452 , \1473 );
or \U$1350 ( \1475 , \1451 , \1474 );
and \U$1351 ( \1476 , \1448 , \1475 );
or \U$1352 ( \1477 , \1447 , \1476 );
and \U$1353 ( \1478 , \1444 , \1477 );
or \U$1354 ( \1479 , \1443 , \1478 );
and \U$1355 ( \1480 , \1440 , \1479 );
or \U$1356 ( \1481 , \1439 , \1480 );
and \U$1357 ( \1482 , \1436 , \1481 );
or \U$1358 ( \1483 , \1435 , \1482 );
and \U$1359 ( \1484 , \1432 , \1483 );
or \U$1360 ( \1485 , \1431 , \1484 );
and \U$1361 ( \1486 , \1428 , \1485 );
or \U$1362 ( \1487 , \1427 , \1486 );
and \U$1363 ( \1488 , \1424 , \1487 );
or \U$1364 ( \1489 , \1423 , \1488 );
and \U$1365 ( \1490 , \1420 , \1489 );
or \U$1366 ( \1491 , \1419 , \1490 );
and \U$1367 ( \1492 , \1416 , \1491 );
or \U$1368 ( \1493 , \1415 , \1492 );
and \U$1369 ( \1494 , \1412 , \1493 );
or \U$1370 ( \1495 , \1411 , \1494 );
and \U$1371 ( \1496 , \1408 , \1495 );
or \U$1372 ( \1497 , \1407 , \1496 );
and \U$1373 ( \1498 , \1404 , \1497 );
or \U$1374 ( \1499 , \1403 , \1498 );
_DC g5d0 ( \1500_nG5d0 , 1'b0 , \941 );
or \U$1376 ( \1501 , RI8928c68_12, RI892a2e8_60);
and \U$1377 ( \1502 , \1501 , \940 );
and \U$1378 ( \1503 , RI89293e8_28, RI8929b68_44);
and \U$1379 ( \1504 , \1503 , \938 );
or \U$1380 ( \1505 , RI8928c68_12, RI89293e8_28);
and \U$1381 ( \1506 , \1505 , \936 );
xor \U$1382 ( \1507 , RI8929b68_44, RI892a2e8_60);
and \U$1383 ( \1508 , \1507 , \934 );
buf \U$1384 ( \1509 , RI89293e8_28);
and \U$1385 ( \1510 , \1509 , \952 );
and \U$1386 ( \1511 , \1342 , \955 );
xor \U$1387 ( \1512 , \1510 , \1511 );
and \U$1388 ( \1513 , \1343 , \1344 );
and \U$1389 ( \1514 , \1345 , \1348 );
or \U$1390 ( \1515 , \1513 , \1514 );
xor \U$1391 ( \1516 , \1512 , \1515 );
and \U$1392 ( \1517 , \1187 , \1193 );
xor \U$1393 ( \1518 , \1516 , \1517 );
and \U$1394 ( \1519 , \1349 , \1350 );
and \U$1395 ( \1520 , \1351 , \1352 );
or \U$1396 ( \1521 , \1519 , \1520 );
xor \U$1397 ( \1522 , \1518 , \1521 );
and \U$1398 ( \1523 , \951 , \1354 );
xor \U$1399 ( \1524 , \1522 , \1523 );
and \U$1400 ( \1525 , \1353 , \1355 );
xor \U$1401 ( \1526 , \1524 , \1525 );
buf \U$1402 ( \1527 , RI8929b68_44);
and \U$1403 ( \1528 , \954 , \1527 );
xor \U$1404 ( \1529 , \1526 , \1528 );
buf \U$1405 ( \1530 , \1529 );
and \U$1406 ( \1531 , \1530 , \932 );
buf \U$1407 ( \1532 , RI8928c68_12);
and \U$1408 ( \1533 , \1532 , \961 );
and \U$1409 ( \1534 , \1359 , \964 );
xor \U$1410 ( \1535 , \1533 , \1534 );
and \U$1411 ( \1536 , \1360 , \1361 );
and \U$1412 ( \1537 , \1362 , \1365 );
or \U$1413 ( \1538 , \1536 , \1537 );
xor \U$1414 ( \1539 , \1535 , \1538 );
and \U$1415 ( \1540 , \1198 , \1204 );
xor \U$1416 ( \1541 , \1539 , \1540 );
and \U$1417 ( \1542 , \1366 , \1367 );
and \U$1418 ( \1543 , \1368 , \1369 );
or \U$1419 ( \1544 , \1542 , \1543 );
xor \U$1420 ( \1545 , \1541 , \1544 );
and \U$1421 ( \1546 , \960 , \1371 );
xor \U$1422 ( \1547 , \1545 , \1546 );
and \U$1423 ( \1548 , \1370 , \1372 );
xor \U$1424 ( \1549 , \1547 , \1548 );
buf \U$1425 ( \1550 , RI892a2e8_60);
and \U$1426 ( \1551 , \963 , \1550 );
xor \U$1427 ( \1552 , \1549 , \1551 );
buf \U$1428 ( \1553 , \1552 );
and \U$1429 ( \1554 , \1553 , \930 );
buf \U$1430 ( \1555 , RI89293e8_28);
buf \U$1431 ( \1556 , RI892a2e8_60);
xor \U$1432 ( \1557 , \1555 , \1556 );
and \U$1433 ( \1558 , \1376 , \1377 );
and \U$1434 ( \1559 , \1377 , \1382 );
and \U$1435 ( \1560 , \1376 , \1382 );
or \U$1436 ( \1561 , \1558 , \1559 , \1560 );
xor \U$1437 ( \1562 , \1557 , \1561 );
buf \U$1438 ( \1563 , \1562 );
and \U$1439 ( \1564 , \1563 , \928 );
buf \U$1440 ( \1565 , RI8928c68_12);
buf \U$1441 ( \1566 , RI8929b68_44);
xor \U$1442 ( \1567 , \1565 , \1566 );
and \U$1443 ( \1568 , \1386 , \1387 );
and \U$1444 ( \1569 , \1387 , \1392 );
and \U$1445 ( \1570 , \1386 , \1392 );
or \U$1446 ( \1571 , \1568 , \1569 , \1570 );
xor \U$1447 ( \1572 , \1567 , \1571 );
buf \U$1448 ( \1573 , \1572 );
and \U$1449 ( \1574 , \1573 , \926 );
and \U$1450 ( \1575 , RI892a2e8_60, \924 );
and \U$1451 ( \1576 , RI8929b68_44, \922 );
and \U$1452 ( \1577 , RI89293e8_28, \920 );
and \U$1453 ( \1578 , RI8928c68_12, \918 );
or \U$1454 ( \1579 , \1500_nG5d0 , \1502 , \1504 , \1506 , \1508 , \1531 , \1554 , \1564 , \1574 , \1575 , \1576 , \1577 , \1578 );
buf \U$1455 ( \1580 , \1579 );
and \U$1456 ( \1581 , \220 , \1580 );
and \U$1457 ( \1582 , \1499 , \1581 );
xor \U$1458 ( \1583 , \1499 , \1581 );
xor \U$1459 ( \1584 , \1404 , \1497 );
and \U$1460 ( \1585 , \1025 , \1580 );
and \U$1461 ( \1586 , \1584 , \1585 );
xor \U$1462 ( \1587 , \1584 , \1585 );
xor \U$1463 ( \1588 , \1408 , \1495 );
and \U$1464 ( \1589 , \1033 , \1580 );
and \U$1465 ( \1590 , \1588 , \1589 );
xor \U$1466 ( \1591 , \1588 , \1589 );
xor \U$1467 ( \1592 , \1412 , \1493 );
and \U$1468 ( \1593 , \1041 , \1580 );
and \U$1469 ( \1594 , \1592 , \1593 );
xor \U$1470 ( \1595 , \1592 , \1593 );
xor \U$1471 ( \1596 , \1416 , \1491 );
and \U$1472 ( \1597 , \1049 , \1580 );
and \U$1473 ( \1598 , \1596 , \1597 );
xor \U$1474 ( \1599 , \1596 , \1597 );
xor \U$1475 ( \1600 , \1420 , \1489 );
and \U$1476 ( \1601 , \1057 , \1580 );
and \U$1477 ( \1602 , \1600 , \1601 );
xor \U$1478 ( \1603 , \1600 , \1601 );
xor \U$1479 ( \1604 , \1424 , \1487 );
and \U$1480 ( \1605 , \1065 , \1580 );
and \U$1481 ( \1606 , \1604 , \1605 );
xor \U$1482 ( \1607 , \1604 , \1605 );
xor \U$1483 ( \1608 , \1428 , \1485 );
and \U$1484 ( \1609 , \1073 , \1580 );
and \U$1485 ( \1610 , \1608 , \1609 );
xor \U$1486 ( \1611 , \1608 , \1609 );
xor \U$1487 ( \1612 , \1432 , \1483 );
and \U$1488 ( \1613 , \1081 , \1580 );
and \U$1489 ( \1614 , \1612 , \1613 );
xor \U$1490 ( \1615 , \1612 , \1613 );
xor \U$1491 ( \1616 , \1436 , \1481 );
and \U$1492 ( \1617 , \1089 , \1580 );
and \U$1493 ( \1618 , \1616 , \1617 );
xor \U$1494 ( \1619 , \1616 , \1617 );
xor \U$1495 ( \1620 , \1440 , \1479 );
and \U$1496 ( \1621 , \1097 , \1580 );
and \U$1497 ( \1622 , \1620 , \1621 );
xor \U$1498 ( \1623 , \1620 , \1621 );
xor \U$1499 ( \1624 , \1444 , \1477 );
and \U$1500 ( \1625 , \1105 , \1580 );
and \U$1501 ( \1626 , \1624 , \1625 );
xor \U$1502 ( \1627 , \1624 , \1625 );
xor \U$1503 ( \1628 , \1448 , \1475 );
and \U$1504 ( \1629 , \1113 , \1580 );
and \U$1505 ( \1630 , \1628 , \1629 );
xor \U$1506 ( \1631 , \1628 , \1629 );
xor \U$1507 ( \1632 , \1452 , \1473 );
and \U$1508 ( \1633 , \1121 , \1580 );
and \U$1509 ( \1634 , \1632 , \1633 );
xor \U$1510 ( \1635 , \1632 , \1633 );
xor \U$1511 ( \1636 , \1456 , \1471 );
and \U$1512 ( \1637 , \1129 , \1580 );
and \U$1513 ( \1638 , \1636 , \1637 );
xor \U$1514 ( \1639 , \1636 , \1637 );
xor \U$1515 ( \1640 , \1460 , \1469 );
and \U$1516 ( \1641 , \1137 , \1580 );
and \U$1517 ( \1642 , \1640 , \1641 );
xor \U$1518 ( \1643 , \1640 , \1641 );
xor \U$1519 ( \1644 , \1464 , \1467 );
and \U$1520 ( \1645 , \1144 , \1580 );
and \U$1521 ( \1646 , \1644 , \1645 );
and \U$1522 ( \1647 , \1643 , \1646 );
or \U$1523 ( \1648 , \1642 , \1647 );
and \U$1524 ( \1649 , \1639 , \1648 );
or \U$1525 ( \1650 , \1638 , \1649 );
and \U$1526 ( \1651 , \1635 , \1650 );
or \U$1527 ( \1652 , \1634 , \1651 );
and \U$1528 ( \1653 , \1631 , \1652 );
or \U$1529 ( \1654 , \1630 , \1653 );
and \U$1530 ( \1655 , \1627 , \1654 );
or \U$1531 ( \1656 , \1626 , \1655 );
and \U$1532 ( \1657 , \1623 , \1656 );
or \U$1533 ( \1658 , \1622 , \1657 );
and \U$1534 ( \1659 , \1619 , \1658 );
or \U$1535 ( \1660 , \1618 , \1659 );
and \U$1536 ( \1661 , \1615 , \1660 );
or \U$1537 ( \1662 , \1614 , \1661 );
and \U$1538 ( \1663 , \1611 , \1662 );
or \U$1539 ( \1664 , \1610 , \1663 );
and \U$1540 ( \1665 , \1607 , \1664 );
or \U$1541 ( \1666 , \1606 , \1665 );
and \U$1542 ( \1667 , \1603 , \1666 );
or \U$1543 ( \1668 , \1602 , \1667 );
and \U$1544 ( \1669 , \1599 , \1668 );
or \U$1545 ( \1670 , \1598 , \1669 );
and \U$1546 ( \1671 , \1595 , \1670 );
or \U$1547 ( \1672 , \1594 , \1671 );
and \U$1548 ( \1673 , \1591 , \1672 );
or \U$1549 ( \1674 , \1590 , \1673 );
and \U$1550 ( \1675 , \1587 , \1674 );
or \U$1551 ( \1676 , \1586 , \1675 );
and \U$1552 ( \1677 , \1583 , \1676 );
or \U$1553 ( \1678 , \1582 , \1677 );
_DC g683 ( \1679_nG683 , 1'b0 , \941 );
or \U$1555 ( \1680 , RI8928bf0_11, RI892a270_59);
and \U$1556 ( \1681 , \1680 , \940 );
and \U$1557 ( \1682 , RI8929370_27, RI8929af0_43);
and \U$1558 ( \1683 , \1682 , \938 );
or \U$1559 ( \1684 , RI8928bf0_11, RI8929370_27);
and \U$1560 ( \1685 , \1684 , \936 );
xor \U$1561 ( \1686 , RI8929af0_43, RI892a270_59);
and \U$1562 ( \1687 , \1686 , \934 );
buf \U$1563 ( \1688 , RI8929370_27);
and \U$1564 ( \1689 , \1688 , \952 );
and \U$1565 ( \1690 , \1509 , \955 );
xor \U$1566 ( \1691 , \1689 , \1690 );
and \U$1567 ( \1692 , \1510 , \1511 );
and \U$1568 ( \1693 , \1512 , \1515 );
or \U$1569 ( \1694 , \1692 , \1693 );
xor \U$1570 ( \1695 , \1691 , \1694 );
and \U$1571 ( \1696 , \1342 , \1193 );
xor \U$1572 ( \1697 , \1695 , \1696 );
and \U$1573 ( \1698 , \1516 , \1517 );
and \U$1574 ( \1699 , \1518 , \1521 );
or \U$1575 ( \1700 , \1698 , \1699 );
xor \U$1576 ( \1701 , \1697 , \1700 );
and \U$1577 ( \1702 , \1187 , \1354 );
xor \U$1578 ( \1703 , \1701 , \1702 );
and \U$1579 ( \1704 , \1522 , \1523 );
and \U$1580 ( \1705 , \1524 , \1525 );
or \U$1581 ( \1706 , \1704 , \1705 );
xor \U$1582 ( \1707 , \1703 , \1706 );
and \U$1583 ( \1708 , \951 , \1527 );
xor \U$1584 ( \1709 , \1707 , \1708 );
and \U$1585 ( \1710 , \1526 , \1528 );
xor \U$1586 ( \1711 , \1709 , \1710 );
buf \U$1587 ( \1712 , RI8929af0_43);
and \U$1588 ( \1713 , \954 , \1712 );
xor \U$1589 ( \1714 , \1711 , \1713 );
buf \U$1590 ( \1715 , \1714 );
and \U$1591 ( \1716 , \1715 , \932 );
buf \U$1592 ( \1717 , RI8928bf0_11);
and \U$1593 ( \1718 , \1717 , \961 );
and \U$1594 ( \1719 , \1532 , \964 );
xor \U$1595 ( \1720 , \1718 , \1719 );
and \U$1596 ( \1721 , \1533 , \1534 );
and \U$1597 ( \1722 , \1535 , \1538 );
or \U$1598 ( \1723 , \1721 , \1722 );
xor \U$1599 ( \1724 , \1720 , \1723 );
and \U$1600 ( \1725 , \1359 , \1204 );
xor \U$1601 ( \1726 , \1724 , \1725 );
and \U$1602 ( \1727 , \1539 , \1540 );
and \U$1603 ( \1728 , \1541 , \1544 );
or \U$1604 ( \1729 , \1727 , \1728 );
xor \U$1605 ( \1730 , \1726 , \1729 );
and \U$1606 ( \1731 , \1198 , \1371 );
xor \U$1607 ( \1732 , \1730 , \1731 );
and \U$1608 ( \1733 , \1545 , \1546 );
and \U$1609 ( \1734 , \1547 , \1548 );
or \U$1610 ( \1735 , \1733 , \1734 );
xor \U$1611 ( \1736 , \1732 , \1735 );
and \U$1612 ( \1737 , \960 , \1550 );
xor \U$1613 ( \1738 , \1736 , \1737 );
and \U$1614 ( \1739 , \1549 , \1551 );
xor \U$1615 ( \1740 , \1738 , \1739 );
buf \U$1616 ( \1741 , RI892a270_59);
and \U$1617 ( \1742 , \963 , \1741 );
xor \U$1618 ( \1743 , \1740 , \1742 );
buf \U$1619 ( \1744 , \1743 );
and \U$1620 ( \1745 , \1744 , \930 );
buf \U$1621 ( \1746 , RI8929370_27);
buf \U$1622 ( \1747 , RI892a270_59);
xor \U$1623 ( \1748 , \1746 , \1747 );
and \U$1624 ( \1749 , \1555 , \1556 );
and \U$1625 ( \1750 , \1556 , \1561 );
and \U$1626 ( \1751 , \1555 , \1561 );
or \U$1627 ( \1752 , \1749 , \1750 , \1751 );
xor \U$1628 ( \1753 , \1748 , \1752 );
buf \U$1629 ( \1754 , \1753 );
and \U$1630 ( \1755 , \1754 , \928 );
buf \U$1631 ( \1756 , RI8928bf0_11);
buf \U$1632 ( \1757 , RI8929af0_43);
xor \U$1633 ( \1758 , \1756 , \1757 );
and \U$1634 ( \1759 , \1565 , \1566 );
and \U$1635 ( \1760 , \1566 , \1571 );
and \U$1636 ( \1761 , \1565 , \1571 );
or \U$1637 ( \1762 , \1759 , \1760 , \1761 );
xor \U$1638 ( \1763 , \1758 , \1762 );
buf \U$1639 ( \1764 , \1763 );
and \U$1640 ( \1765 , \1764 , \926 );
and \U$1641 ( \1766 , RI892a270_59, \924 );
and \U$1642 ( \1767 , RI8929af0_43, \922 );
and \U$1643 ( \1768 , RI8929370_27, \920 );
and \U$1644 ( \1769 , RI8928bf0_11, \918 );
or \U$1645 ( \1770 , \1679_nG683 , \1681 , \1683 , \1685 , \1687 , \1716 , \1745 , \1755 , \1765 , \1766 , \1767 , \1768 , \1769 );
buf \U$1646 ( \1771 , \1770 );
and \U$1647 ( \1772 , \220 , \1771 );
and \U$1648 ( \1773 , \1678 , \1772 );
xor \U$1649 ( \1774 , \1678 , \1772 );
xor \U$1650 ( \1775 , \1583 , \1676 );
and \U$1651 ( \1776 , \1025 , \1771 );
and \U$1652 ( \1777 , \1775 , \1776 );
xor \U$1653 ( \1778 , \1775 , \1776 );
xor \U$1654 ( \1779 , \1587 , \1674 );
and \U$1655 ( \1780 , \1033 , \1771 );
and \U$1656 ( \1781 , \1779 , \1780 );
xor \U$1657 ( \1782 , \1779 , \1780 );
xor \U$1658 ( \1783 , \1591 , \1672 );
and \U$1659 ( \1784 , \1041 , \1771 );
and \U$1660 ( \1785 , \1783 , \1784 );
xor \U$1661 ( \1786 , \1783 , \1784 );
xor \U$1662 ( \1787 , \1595 , \1670 );
and \U$1663 ( \1788 , \1049 , \1771 );
and \U$1664 ( \1789 , \1787 , \1788 );
xor \U$1665 ( \1790 , \1787 , \1788 );
xor \U$1666 ( \1791 , \1599 , \1668 );
and \U$1667 ( \1792 , \1057 , \1771 );
and \U$1668 ( \1793 , \1791 , \1792 );
xor \U$1669 ( \1794 , \1791 , \1792 );
xor \U$1670 ( \1795 , \1603 , \1666 );
and \U$1671 ( \1796 , \1065 , \1771 );
and \U$1672 ( \1797 , \1795 , \1796 );
xor \U$1673 ( \1798 , \1795 , \1796 );
xor \U$1674 ( \1799 , \1607 , \1664 );
and \U$1675 ( \1800 , \1073 , \1771 );
and \U$1676 ( \1801 , \1799 , \1800 );
xor \U$1677 ( \1802 , \1799 , \1800 );
xor \U$1678 ( \1803 , \1611 , \1662 );
and \U$1679 ( \1804 , \1081 , \1771 );
and \U$1680 ( \1805 , \1803 , \1804 );
xor \U$1681 ( \1806 , \1803 , \1804 );
xor \U$1682 ( \1807 , \1615 , \1660 );
and \U$1683 ( \1808 , \1089 , \1771 );
and \U$1684 ( \1809 , \1807 , \1808 );
xor \U$1685 ( \1810 , \1807 , \1808 );
xor \U$1686 ( \1811 , \1619 , \1658 );
and \U$1687 ( \1812 , \1097 , \1771 );
and \U$1688 ( \1813 , \1811 , \1812 );
xor \U$1689 ( \1814 , \1811 , \1812 );
xor \U$1690 ( \1815 , \1623 , \1656 );
and \U$1691 ( \1816 , \1105 , \1771 );
and \U$1692 ( \1817 , \1815 , \1816 );
xor \U$1693 ( \1818 , \1815 , \1816 );
xor \U$1694 ( \1819 , \1627 , \1654 );
and \U$1695 ( \1820 , \1113 , \1771 );
and \U$1696 ( \1821 , \1819 , \1820 );
xor \U$1697 ( \1822 , \1819 , \1820 );
xor \U$1698 ( \1823 , \1631 , \1652 );
and \U$1699 ( \1824 , \1121 , \1771 );
and \U$1700 ( \1825 , \1823 , \1824 );
xor \U$1701 ( \1826 , \1823 , \1824 );
xor \U$1702 ( \1827 , \1635 , \1650 );
and \U$1703 ( \1828 , \1129 , \1771 );
and \U$1704 ( \1829 , \1827 , \1828 );
xor \U$1705 ( \1830 , \1827 , \1828 );
xor \U$1706 ( \1831 , \1639 , \1648 );
and \U$1707 ( \1832 , \1137 , \1771 );
and \U$1708 ( \1833 , \1831 , \1832 );
xor \U$1709 ( \1834 , \1831 , \1832 );
xor \U$1710 ( \1835 , \1643 , \1646 );
and \U$1711 ( \1836 , \1144 , \1771 );
and \U$1712 ( \1837 , \1835 , \1836 );
and \U$1713 ( \1838 , \1834 , \1837 );
or \U$1714 ( \1839 , \1833 , \1838 );
and \U$1715 ( \1840 , \1830 , \1839 );
or \U$1716 ( \1841 , \1829 , \1840 );
and \U$1717 ( \1842 , \1826 , \1841 );
or \U$1718 ( \1843 , \1825 , \1842 );
and \U$1719 ( \1844 , \1822 , \1843 );
or \U$1720 ( \1845 , \1821 , \1844 );
and \U$1721 ( \1846 , \1818 , \1845 );
or \U$1722 ( \1847 , \1817 , \1846 );
and \U$1723 ( \1848 , \1814 , \1847 );
or \U$1724 ( \1849 , \1813 , \1848 );
and \U$1725 ( \1850 , \1810 , \1849 );
or \U$1726 ( \1851 , \1809 , \1850 );
and \U$1727 ( \1852 , \1806 , \1851 );
or \U$1728 ( \1853 , \1805 , \1852 );
and \U$1729 ( \1854 , \1802 , \1853 );
or \U$1730 ( \1855 , \1801 , \1854 );
and \U$1731 ( \1856 , \1798 , \1855 );
or \U$1732 ( \1857 , \1797 , \1856 );
and \U$1733 ( \1858 , \1794 , \1857 );
or \U$1734 ( \1859 , \1793 , \1858 );
and \U$1735 ( \1860 , \1790 , \1859 );
or \U$1736 ( \1861 , \1789 , \1860 );
and \U$1737 ( \1862 , \1786 , \1861 );
or \U$1738 ( \1863 , \1785 , \1862 );
and \U$1739 ( \1864 , \1782 , \1863 );
or \U$1740 ( \1865 , \1781 , \1864 );
and \U$1741 ( \1866 , \1778 , \1865 );
or \U$1742 ( \1867 , \1777 , \1866 );
and \U$1743 ( \1868 , \1774 , \1867 );
or \U$1744 ( \1869 , \1773 , \1868 );
_DC g742 ( \1870_nG742 , 1'b0 , \941 );
or \U$1746 ( \1871 , RI8928b78_10, RI892a1f8_58);
and \U$1747 ( \1872 , \1871 , \940 );
and \U$1748 ( \1873 , RI89292f8_26, RI8929a78_42);
and \U$1749 ( \1874 , \1873 , \938 );
or \U$1750 ( \1875 , RI8928b78_10, RI89292f8_26);
and \U$1751 ( \1876 , \1875 , \936 );
xor \U$1752 ( \1877 , RI8929a78_42, RI892a1f8_58);
and \U$1753 ( \1878 , \1877 , \934 );
buf \U$1754 ( \1879 , RI89292f8_26);
and \U$1755 ( \1880 , \1879 , \952 );
and \U$1756 ( \1881 , \1688 , \955 );
xor \U$1757 ( \1882 , \1880 , \1881 );
and \U$1758 ( \1883 , \1689 , \1690 );
and \U$1759 ( \1884 , \1691 , \1694 );
or \U$1760 ( \1885 , \1883 , \1884 );
xor \U$1761 ( \1886 , \1882 , \1885 );
and \U$1762 ( \1887 , \1509 , \1193 );
xor \U$1763 ( \1888 , \1886 , \1887 );
and \U$1764 ( \1889 , \1695 , \1696 );
and \U$1765 ( \1890 , \1697 , \1700 );
or \U$1766 ( \1891 , \1889 , \1890 );
xor \U$1767 ( \1892 , \1888 , \1891 );
and \U$1768 ( \1893 , \1342 , \1354 );
xor \U$1769 ( \1894 , \1892 , \1893 );
and \U$1770 ( \1895 , \1701 , \1702 );
and \U$1771 ( \1896 , \1703 , \1706 );
or \U$1772 ( \1897 , \1895 , \1896 );
xor \U$1773 ( \1898 , \1894 , \1897 );
and \U$1774 ( \1899 , \1187 , \1527 );
xor \U$1775 ( \1900 , \1898 , \1899 );
and \U$1776 ( \1901 , \1707 , \1708 );
and \U$1777 ( \1902 , \1709 , \1710 );
or \U$1778 ( \1903 , \1901 , \1902 );
xor \U$1779 ( \1904 , \1900 , \1903 );
and \U$1780 ( \1905 , \951 , \1712 );
xor \U$1781 ( \1906 , \1904 , \1905 );
and \U$1782 ( \1907 , \1711 , \1713 );
xor \U$1783 ( \1908 , \1906 , \1907 );
buf \U$1784 ( \1909 , RI8929a78_42);
and \U$1785 ( \1910 , \954 , \1909 );
xor \U$1786 ( \1911 , \1908 , \1910 );
buf \U$1787 ( \1912 , \1911 );
and \U$1788 ( \1913 , \1912 , \932 );
buf \U$1789 ( \1914 , RI8928b78_10);
and \U$1790 ( \1915 , \1914 , \961 );
and \U$1791 ( \1916 , \1717 , \964 );
xor \U$1792 ( \1917 , \1915 , \1916 );
and \U$1793 ( \1918 , \1718 , \1719 );
and \U$1794 ( \1919 , \1720 , \1723 );
or \U$1795 ( \1920 , \1918 , \1919 );
xor \U$1796 ( \1921 , \1917 , \1920 );
and \U$1797 ( \1922 , \1532 , \1204 );
xor \U$1798 ( \1923 , \1921 , \1922 );
and \U$1799 ( \1924 , \1724 , \1725 );
and \U$1800 ( \1925 , \1726 , \1729 );
or \U$1801 ( \1926 , \1924 , \1925 );
xor \U$1802 ( \1927 , \1923 , \1926 );
and \U$1803 ( \1928 , \1359 , \1371 );
xor \U$1804 ( \1929 , \1927 , \1928 );
and \U$1805 ( \1930 , \1730 , \1731 );
and \U$1806 ( \1931 , \1732 , \1735 );
or \U$1807 ( \1932 , \1930 , \1931 );
xor \U$1808 ( \1933 , \1929 , \1932 );
and \U$1809 ( \1934 , \1198 , \1550 );
xor \U$1810 ( \1935 , \1933 , \1934 );
and \U$1811 ( \1936 , \1736 , \1737 );
and \U$1812 ( \1937 , \1738 , \1739 );
or \U$1813 ( \1938 , \1936 , \1937 );
xor \U$1814 ( \1939 , \1935 , \1938 );
and \U$1815 ( \1940 , \960 , \1741 );
xor \U$1816 ( \1941 , \1939 , \1940 );
and \U$1817 ( \1942 , \1740 , \1742 );
xor \U$1818 ( \1943 , \1941 , \1942 );
buf \U$1819 ( \1944 , RI892a1f8_58);
and \U$1820 ( \1945 , \963 , \1944 );
xor \U$1821 ( \1946 , \1943 , \1945 );
buf \U$1822 ( \1947 , \1946 );
and \U$1823 ( \1948 , \1947 , \930 );
buf \U$1824 ( \1949 , RI89292f8_26);
buf \U$1825 ( \1950 , RI892a1f8_58);
xor \U$1826 ( \1951 , \1949 , \1950 );
and \U$1827 ( \1952 , \1746 , \1747 );
and \U$1828 ( \1953 , \1747 , \1752 );
and \U$1829 ( \1954 , \1746 , \1752 );
or \U$1830 ( \1955 , \1952 , \1953 , \1954 );
xor \U$1831 ( \1956 , \1951 , \1955 );
buf \U$1832 ( \1957 , \1956 );
and \U$1833 ( \1958 , \1957 , \928 );
buf \U$1834 ( \1959 , RI8928b78_10);
buf \U$1835 ( \1960 , RI8929a78_42);
xor \U$1836 ( \1961 , \1959 , \1960 );
and \U$1837 ( \1962 , \1756 , \1757 );
and \U$1838 ( \1963 , \1757 , \1762 );
and \U$1839 ( \1964 , \1756 , \1762 );
or \U$1840 ( \1965 , \1962 , \1963 , \1964 );
xor \U$1841 ( \1966 , \1961 , \1965 );
buf \U$1842 ( \1967 , \1966 );
and \U$1843 ( \1968 , \1967 , \926 );
and \U$1844 ( \1969 , RI892a1f8_58, \924 );
and \U$1845 ( \1970 , RI8929a78_42, \922 );
and \U$1846 ( \1971 , RI89292f8_26, \920 );
and \U$1847 ( \1972 , RI8928b78_10, \918 );
or \U$1848 ( \1973 , \1870_nG742 , \1872 , \1874 , \1876 , \1878 , \1913 , \1948 , \1958 , \1968 , \1969 , \1970 , \1971 , \1972 );
buf \U$1849 ( \1974 , \1973 );
and \U$1850 ( \1975 , \220 , \1974 );
and \U$1851 ( \1976 , \1869 , \1975 );
xor \U$1852 ( \1977 , \1869 , \1975 );
xor \U$1853 ( \1978 , \1774 , \1867 );
and \U$1854 ( \1979 , \1025 , \1974 );
and \U$1855 ( \1980 , \1978 , \1979 );
xor \U$1856 ( \1981 , \1978 , \1979 );
xor \U$1857 ( \1982 , \1778 , \1865 );
and \U$1858 ( \1983 , \1033 , \1974 );
and \U$1859 ( \1984 , \1982 , \1983 );
xor \U$1860 ( \1985 , \1982 , \1983 );
xor \U$1861 ( \1986 , \1782 , \1863 );
and \U$1862 ( \1987 , \1041 , \1974 );
and \U$1863 ( \1988 , \1986 , \1987 );
xor \U$1864 ( \1989 , \1986 , \1987 );
xor \U$1865 ( \1990 , \1786 , \1861 );
and \U$1866 ( \1991 , \1049 , \1974 );
and \U$1867 ( \1992 , \1990 , \1991 );
xor \U$1868 ( \1993 , \1990 , \1991 );
xor \U$1869 ( \1994 , \1790 , \1859 );
and \U$1870 ( \1995 , \1057 , \1974 );
and \U$1871 ( \1996 , \1994 , \1995 );
xor \U$1872 ( \1997 , \1994 , \1995 );
xor \U$1873 ( \1998 , \1794 , \1857 );
and \U$1874 ( \1999 , \1065 , \1974 );
and \U$1875 ( \2000 , \1998 , \1999 );
xor \U$1876 ( \2001 , \1998 , \1999 );
xor \U$1877 ( \2002 , \1798 , \1855 );
and \U$1878 ( \2003 , \1073 , \1974 );
and \U$1879 ( \2004 , \2002 , \2003 );
xor \U$1880 ( \2005 , \2002 , \2003 );
xor \U$1881 ( \2006 , \1802 , \1853 );
and \U$1882 ( \2007 , \1081 , \1974 );
and \U$1883 ( \2008 , \2006 , \2007 );
xor \U$1884 ( \2009 , \2006 , \2007 );
xor \U$1885 ( \2010 , \1806 , \1851 );
and \U$1886 ( \2011 , \1089 , \1974 );
and \U$1887 ( \2012 , \2010 , \2011 );
xor \U$1888 ( \2013 , \2010 , \2011 );
xor \U$1889 ( \2014 , \1810 , \1849 );
and \U$1890 ( \2015 , \1097 , \1974 );
and \U$1891 ( \2016 , \2014 , \2015 );
xor \U$1892 ( \2017 , \2014 , \2015 );
xor \U$1893 ( \2018 , \1814 , \1847 );
and \U$1894 ( \2019 , \1105 , \1974 );
and \U$1895 ( \2020 , \2018 , \2019 );
xor \U$1896 ( \2021 , \2018 , \2019 );
xor \U$1897 ( \2022 , \1818 , \1845 );
and \U$1898 ( \2023 , \1113 , \1974 );
and \U$1899 ( \2024 , \2022 , \2023 );
xor \U$1900 ( \2025 , \2022 , \2023 );
xor \U$1901 ( \2026 , \1822 , \1843 );
and \U$1902 ( \2027 , \1121 , \1974 );
and \U$1903 ( \2028 , \2026 , \2027 );
xor \U$1904 ( \2029 , \2026 , \2027 );
xor \U$1905 ( \2030 , \1826 , \1841 );
and \U$1906 ( \2031 , \1129 , \1974 );
and \U$1907 ( \2032 , \2030 , \2031 );
xor \U$1908 ( \2033 , \2030 , \2031 );
xor \U$1909 ( \2034 , \1830 , \1839 );
and \U$1910 ( \2035 , \1137 , \1974 );
and \U$1911 ( \2036 , \2034 , \2035 );
xor \U$1912 ( \2037 , \2034 , \2035 );
xor \U$1913 ( \2038 , \1834 , \1837 );
and \U$1914 ( \2039 , \1144 , \1974 );
and \U$1915 ( \2040 , \2038 , \2039 );
and \U$1916 ( \2041 , \2037 , \2040 );
or \U$1917 ( \2042 , \2036 , \2041 );
and \U$1918 ( \2043 , \2033 , \2042 );
or \U$1919 ( \2044 , \2032 , \2043 );
and \U$1920 ( \2045 , \2029 , \2044 );
or \U$1921 ( \2046 , \2028 , \2045 );
and \U$1922 ( \2047 , \2025 , \2046 );
or \U$1923 ( \2048 , \2024 , \2047 );
and \U$1924 ( \2049 , \2021 , \2048 );
or \U$1925 ( \2050 , \2020 , \2049 );
and \U$1926 ( \2051 , \2017 , \2050 );
or \U$1927 ( \2052 , \2016 , \2051 );
and \U$1928 ( \2053 , \2013 , \2052 );
or \U$1929 ( \2054 , \2012 , \2053 );
and \U$1930 ( \2055 , \2009 , \2054 );
or \U$1931 ( \2056 , \2008 , \2055 );
and \U$1932 ( \2057 , \2005 , \2056 );
or \U$1933 ( \2058 , \2004 , \2057 );
and \U$1934 ( \2059 , \2001 , \2058 );
or \U$1935 ( \2060 , \2000 , \2059 );
and \U$1936 ( \2061 , \1997 , \2060 );
or \U$1937 ( \2062 , \1996 , \2061 );
and \U$1938 ( \2063 , \1993 , \2062 );
or \U$1939 ( \2064 , \1992 , \2063 );
and \U$1940 ( \2065 , \1989 , \2064 );
or \U$1941 ( \2066 , \1988 , \2065 );
and \U$1942 ( \2067 , \1985 , \2066 );
or \U$1943 ( \2068 , \1984 , \2067 );
and \U$1944 ( \2069 , \1981 , \2068 );
or \U$1945 ( \2070 , \1980 , \2069 );
and \U$1946 ( \2071 , \1977 , \2070 );
or \U$1947 ( \2072 , \1976 , \2071 );
_DC g80d ( \2073_nG80d , 1'b0 , \941 );
or \U$1949 ( \2074 , RI8928b00_9, RI892a180_57);
and \U$1950 ( \2075 , \2074 , \940 );
and \U$1951 ( \2076 , RI8929280_25, RI8929a00_41);
and \U$1952 ( \2077 , \2076 , \938 );
or \U$1953 ( \2078 , RI8928b00_9, RI8929280_25);
and \U$1954 ( \2079 , \2078 , \936 );
xor \U$1955 ( \2080 , RI8929a00_41, RI892a180_57);
and \U$1956 ( \2081 , \2080 , \934 );
buf \U$1957 ( \2082 , RI8929280_25);
and \U$1958 ( \2083 , \2082 , \952 );
and \U$1959 ( \2084 , \1879 , \955 );
xor \U$1960 ( \2085 , \2083 , \2084 );
and \U$1961 ( \2086 , \1880 , \1881 );
and \U$1962 ( \2087 , \1882 , \1885 );
or \U$1963 ( \2088 , \2086 , \2087 );
xor \U$1964 ( \2089 , \2085 , \2088 );
and \U$1965 ( \2090 , \1688 , \1193 );
xor \U$1966 ( \2091 , \2089 , \2090 );
and \U$1967 ( \2092 , \1886 , \1887 );
and \U$1968 ( \2093 , \1888 , \1891 );
or \U$1969 ( \2094 , \2092 , \2093 );
xor \U$1970 ( \2095 , \2091 , \2094 );
and \U$1971 ( \2096 , \1509 , \1354 );
xor \U$1972 ( \2097 , \2095 , \2096 );
and \U$1973 ( \2098 , \1892 , \1893 );
and \U$1974 ( \2099 , \1894 , \1897 );
or \U$1975 ( \2100 , \2098 , \2099 );
xor \U$1976 ( \2101 , \2097 , \2100 );
and \U$1977 ( \2102 , \1342 , \1527 );
xor \U$1978 ( \2103 , \2101 , \2102 );
and \U$1979 ( \2104 , \1898 , \1899 );
and \U$1980 ( \2105 , \1900 , \1903 );
or \U$1981 ( \2106 , \2104 , \2105 );
xor \U$1982 ( \2107 , \2103 , \2106 );
and \U$1983 ( \2108 , \1187 , \1712 );
xor \U$1984 ( \2109 , \2107 , \2108 );
and \U$1985 ( \2110 , \1904 , \1905 );
and \U$1986 ( \2111 , \1906 , \1907 );
or \U$1987 ( \2112 , \2110 , \2111 );
xor \U$1988 ( \2113 , \2109 , \2112 );
and \U$1989 ( \2114 , \951 , \1909 );
xor \U$1990 ( \2115 , \2113 , \2114 );
and \U$1991 ( \2116 , \1908 , \1910 );
xor \U$1992 ( \2117 , \2115 , \2116 );
buf \U$1993 ( \2118 , RI8929a00_41);
and \U$1994 ( \2119 , \954 , \2118 );
xor \U$1995 ( \2120 , \2117 , \2119 );
buf \U$1996 ( \2121 , \2120 );
and \U$1997 ( \2122 , \2121 , \932 );
buf \U$1998 ( \2123 , RI8928b00_9);
and \U$1999 ( \2124 , \2123 , \961 );
and \U$2000 ( \2125 , \1914 , \964 );
xor \U$2001 ( \2126 , \2124 , \2125 );
and \U$2002 ( \2127 , \1915 , \1916 );
and \U$2003 ( \2128 , \1917 , \1920 );
or \U$2004 ( \2129 , \2127 , \2128 );
xor \U$2005 ( \2130 , \2126 , \2129 );
and \U$2006 ( \2131 , \1717 , \1204 );
xor \U$2007 ( \2132 , \2130 , \2131 );
and \U$2008 ( \2133 , \1921 , \1922 );
and \U$2009 ( \2134 , \1923 , \1926 );
or \U$2010 ( \2135 , \2133 , \2134 );
xor \U$2011 ( \2136 , \2132 , \2135 );
and \U$2012 ( \2137 , \1532 , \1371 );
xor \U$2013 ( \2138 , \2136 , \2137 );
and \U$2014 ( \2139 , \1927 , \1928 );
and \U$2015 ( \2140 , \1929 , \1932 );
or \U$2016 ( \2141 , \2139 , \2140 );
xor \U$2017 ( \2142 , \2138 , \2141 );
and \U$2018 ( \2143 , \1359 , \1550 );
xor \U$2019 ( \2144 , \2142 , \2143 );
and \U$2020 ( \2145 , \1933 , \1934 );
and \U$2021 ( \2146 , \1935 , \1938 );
or \U$2022 ( \2147 , \2145 , \2146 );
xor \U$2023 ( \2148 , \2144 , \2147 );
and \U$2024 ( \2149 , \1198 , \1741 );
xor \U$2025 ( \2150 , \2148 , \2149 );
and \U$2026 ( \2151 , \1939 , \1940 );
and \U$2027 ( \2152 , \1941 , \1942 );
or \U$2028 ( \2153 , \2151 , \2152 );
xor \U$2029 ( \2154 , \2150 , \2153 );
and \U$2030 ( \2155 , \960 , \1944 );
xor \U$2031 ( \2156 , \2154 , \2155 );
and \U$2032 ( \2157 , \1943 , \1945 );
xor \U$2033 ( \2158 , \2156 , \2157 );
buf \U$2034 ( \2159 , RI892a180_57);
and \U$2035 ( \2160 , \963 , \2159 );
xor \U$2036 ( \2161 , \2158 , \2160 );
buf \U$2037 ( \2162 , \2161 );
and \U$2038 ( \2163 , \2162 , \930 );
buf \U$2039 ( \2164 , RI8929280_25);
buf \U$2040 ( \2165 , RI892a180_57);
xor \U$2041 ( \2166 , \2164 , \2165 );
and \U$2042 ( \2167 , \1949 , \1950 );
and \U$2043 ( \2168 , \1950 , \1955 );
and \U$2044 ( \2169 , \1949 , \1955 );
or \U$2045 ( \2170 , \2167 , \2168 , \2169 );
xor \U$2046 ( \2171 , \2166 , \2170 );
buf \U$2047 ( \2172 , \2171 );
and \U$2048 ( \2173 , \2172 , \928 );
buf \U$2049 ( \2174 , RI8928b00_9);
buf \U$2050 ( \2175 , RI8929a00_41);
xor \U$2051 ( \2176 , \2174 , \2175 );
and \U$2052 ( \2177 , \1959 , \1960 );
and \U$2053 ( \2178 , \1960 , \1965 );
and \U$2054 ( \2179 , \1959 , \1965 );
or \U$2055 ( \2180 , \2177 , \2178 , \2179 );
xor \U$2056 ( \2181 , \2176 , \2180 );
buf \U$2057 ( \2182 , \2181 );
and \U$2058 ( \2183 , \2182 , \926 );
and \U$2059 ( \2184 , RI892a180_57, \924 );
and \U$2060 ( \2185 , RI8929a00_41, \922 );
and \U$2061 ( \2186 , RI8929280_25, \920 );
and \U$2062 ( \2187 , RI8928b00_9, \918 );
or \U$2063 ( \2188 , \2073_nG80d , \2075 , \2077 , \2079 , \2081 , \2122 , \2163 , \2173 , \2183 , \2184 , \2185 , \2186 , \2187 );
buf \U$2064 ( \2189 , \2188 );
and \U$2065 ( \2190 , \220 , \2189 );
and \U$2066 ( \2191 , \2072 , \2190 );
xor \U$2067 ( \2192 , \2072 , \2190 );
xor \U$2068 ( \2193 , \1977 , \2070 );
and \U$2069 ( \2194 , \1025 , \2189 );
and \U$2070 ( \2195 , \2193 , \2194 );
xor \U$2071 ( \2196 , \2193 , \2194 );
xor \U$2072 ( \2197 , \1981 , \2068 );
and \U$2073 ( \2198 , \1033 , \2189 );
and \U$2074 ( \2199 , \2197 , \2198 );
xor \U$2075 ( \2200 , \2197 , \2198 );
xor \U$2076 ( \2201 , \1985 , \2066 );
and \U$2077 ( \2202 , \1041 , \2189 );
and \U$2078 ( \2203 , \2201 , \2202 );
xor \U$2079 ( \2204 , \2201 , \2202 );
xor \U$2080 ( \2205 , \1989 , \2064 );
and \U$2081 ( \2206 , \1049 , \2189 );
and \U$2082 ( \2207 , \2205 , \2206 );
xor \U$2083 ( \2208 , \2205 , \2206 );
xor \U$2084 ( \2209 , \1993 , \2062 );
and \U$2085 ( \2210 , \1057 , \2189 );
and \U$2086 ( \2211 , \2209 , \2210 );
xor \U$2087 ( \2212 , \2209 , \2210 );
xor \U$2088 ( \2213 , \1997 , \2060 );
and \U$2089 ( \2214 , \1065 , \2189 );
and \U$2090 ( \2215 , \2213 , \2214 );
xor \U$2091 ( \2216 , \2213 , \2214 );
xor \U$2092 ( \2217 , \2001 , \2058 );
and \U$2093 ( \2218 , \1073 , \2189 );
and \U$2094 ( \2219 , \2217 , \2218 );
xor \U$2095 ( \2220 , \2217 , \2218 );
xor \U$2096 ( \2221 , \2005 , \2056 );
and \U$2097 ( \2222 , \1081 , \2189 );
and \U$2098 ( \2223 , \2221 , \2222 );
xor \U$2099 ( \2224 , \2221 , \2222 );
xor \U$2100 ( \2225 , \2009 , \2054 );
and \U$2101 ( \2226 , \1089 , \2189 );
and \U$2102 ( \2227 , \2225 , \2226 );
xor \U$2103 ( \2228 , \2225 , \2226 );
xor \U$2104 ( \2229 , \2013 , \2052 );
and \U$2105 ( \2230 , \1097 , \2189 );
and \U$2106 ( \2231 , \2229 , \2230 );
xor \U$2107 ( \2232 , \2229 , \2230 );
xor \U$2108 ( \2233 , \2017 , \2050 );
and \U$2109 ( \2234 , \1105 , \2189 );
and \U$2110 ( \2235 , \2233 , \2234 );
xor \U$2111 ( \2236 , \2233 , \2234 );
xor \U$2112 ( \2237 , \2021 , \2048 );
and \U$2113 ( \2238 , \1113 , \2189 );
and \U$2114 ( \2239 , \2237 , \2238 );
xor \U$2115 ( \2240 , \2237 , \2238 );
xor \U$2116 ( \2241 , \2025 , \2046 );
and \U$2117 ( \2242 , \1121 , \2189 );
and \U$2118 ( \2243 , \2241 , \2242 );
xor \U$2119 ( \2244 , \2241 , \2242 );
xor \U$2120 ( \2245 , \2029 , \2044 );
and \U$2121 ( \2246 , \1129 , \2189 );
and \U$2122 ( \2247 , \2245 , \2246 );
xor \U$2123 ( \2248 , \2245 , \2246 );
xor \U$2124 ( \2249 , \2033 , \2042 );
and \U$2125 ( \2250 , \1137 , \2189 );
and \U$2126 ( \2251 , \2249 , \2250 );
xor \U$2127 ( \2252 , \2249 , \2250 );
xor \U$2128 ( \2253 , \2037 , \2040 );
and \U$2129 ( \2254 , \1144 , \2189 );
and \U$2130 ( \2255 , \2253 , \2254 );
and \U$2131 ( \2256 , \2252 , \2255 );
or \U$2132 ( \2257 , \2251 , \2256 );
and \U$2133 ( \2258 , \2248 , \2257 );
or \U$2134 ( \2259 , \2247 , \2258 );
and \U$2135 ( \2260 , \2244 , \2259 );
or \U$2136 ( \2261 , \2243 , \2260 );
and \U$2137 ( \2262 , \2240 , \2261 );
or \U$2138 ( \2263 , \2239 , \2262 );
and \U$2139 ( \2264 , \2236 , \2263 );
or \U$2140 ( \2265 , \2235 , \2264 );
and \U$2141 ( \2266 , \2232 , \2265 );
or \U$2142 ( \2267 , \2231 , \2266 );
and \U$2143 ( \2268 , \2228 , \2267 );
or \U$2144 ( \2269 , \2227 , \2268 );
and \U$2145 ( \2270 , \2224 , \2269 );
or \U$2146 ( \2271 , \2223 , \2270 );
and \U$2147 ( \2272 , \2220 , \2271 );
or \U$2148 ( \2273 , \2219 , \2272 );
and \U$2149 ( \2274 , \2216 , \2273 );
or \U$2150 ( \2275 , \2215 , \2274 );
and \U$2151 ( \2276 , \2212 , \2275 );
or \U$2152 ( \2277 , \2211 , \2276 );
and \U$2153 ( \2278 , \2208 , \2277 );
or \U$2154 ( \2279 , \2207 , \2278 );
and \U$2155 ( \2280 , \2204 , \2279 );
or \U$2156 ( \2281 , \2203 , \2280 );
and \U$2157 ( \2282 , \2200 , \2281 );
or \U$2158 ( \2283 , \2199 , \2282 );
and \U$2159 ( \2284 , \2196 , \2283 );
or \U$2160 ( \2285 , \2195 , \2284 );
and \U$2161 ( \2286 , \2192 , \2285 );
or \U$2162 ( \2287 , \2191 , \2286 );
_DC g8e4 ( \2288_nG8e4 , 1'b0 , \941 );
or \U$2164 ( \2289 , RI8928a88_8, RI892a108_56);
and \U$2165 ( \2290 , \2289 , \940 );
and \U$2166 ( \2291 , RI8929208_24, RI8929988_40);
and \U$2167 ( \2292 , \2291 , \938 );
or \U$2168 ( \2293 , RI8928a88_8, RI8929208_24);
and \U$2169 ( \2294 , \2293 , \936 );
xor \U$2170 ( \2295 , RI8929988_40, RI892a108_56);
and \U$2171 ( \2296 , \2295 , \934 );
buf \U$2172 ( \2297 , RI8929208_24);
and \U$2173 ( \2298 , \2297 , \952 );
and \U$2174 ( \2299 , \2082 , \955 );
xor \U$2175 ( \2300 , \2298 , \2299 );
and \U$2176 ( \2301 , \2083 , \2084 );
and \U$2177 ( \2302 , \2085 , \2088 );
or \U$2178 ( \2303 , \2301 , \2302 );
xor \U$2179 ( \2304 , \2300 , \2303 );
and \U$2180 ( \2305 , \1879 , \1193 );
xor \U$2181 ( \2306 , \2304 , \2305 );
and \U$2182 ( \2307 , \2089 , \2090 );
and \U$2183 ( \2308 , \2091 , \2094 );
or \U$2184 ( \2309 , \2307 , \2308 );
xor \U$2185 ( \2310 , \2306 , \2309 );
and \U$2186 ( \2311 , \1688 , \1354 );
xor \U$2187 ( \2312 , \2310 , \2311 );
and \U$2188 ( \2313 , \2095 , \2096 );
and \U$2189 ( \2314 , \2097 , \2100 );
or \U$2190 ( \2315 , \2313 , \2314 );
xor \U$2191 ( \2316 , \2312 , \2315 );
and \U$2192 ( \2317 , \1509 , \1527 );
xor \U$2193 ( \2318 , \2316 , \2317 );
and \U$2194 ( \2319 , \2101 , \2102 );
and \U$2195 ( \2320 , \2103 , \2106 );
or \U$2196 ( \2321 , \2319 , \2320 );
xor \U$2197 ( \2322 , \2318 , \2321 );
and \U$2198 ( \2323 , \1342 , \1712 );
xor \U$2199 ( \2324 , \2322 , \2323 );
and \U$2200 ( \2325 , \2107 , \2108 );
and \U$2201 ( \2326 , \2109 , \2112 );
or \U$2202 ( \2327 , \2325 , \2326 );
xor \U$2203 ( \2328 , \2324 , \2327 );
and \U$2204 ( \2329 , \1187 , \1909 );
xor \U$2205 ( \2330 , \2328 , \2329 );
and \U$2206 ( \2331 , \2113 , \2114 );
and \U$2207 ( \2332 , \2115 , \2116 );
or \U$2208 ( \2333 , \2331 , \2332 );
xor \U$2209 ( \2334 , \2330 , \2333 );
and \U$2210 ( \2335 , \951 , \2118 );
xor \U$2211 ( \2336 , \2334 , \2335 );
and \U$2212 ( \2337 , \2117 , \2119 );
xor \U$2213 ( \2338 , \2336 , \2337 );
buf \U$2214 ( \2339 , RI8929988_40);
and \U$2215 ( \2340 , \954 , \2339 );
xor \U$2216 ( \2341 , \2338 , \2340 );
buf \U$2217 ( \2342 , \2341 );
and \U$2218 ( \2343 , \2342 , \932 );
buf \U$2219 ( \2344 , RI8928a88_8);
and \U$2220 ( \2345 , \2344 , \961 );
and \U$2221 ( \2346 , \2123 , \964 );
xor \U$2222 ( \2347 , \2345 , \2346 );
and \U$2223 ( \2348 , \2124 , \2125 );
and \U$2224 ( \2349 , \2126 , \2129 );
or \U$2225 ( \2350 , \2348 , \2349 );
xor \U$2226 ( \2351 , \2347 , \2350 );
and \U$2227 ( \2352 , \1914 , \1204 );
xor \U$2228 ( \2353 , \2351 , \2352 );
and \U$2229 ( \2354 , \2130 , \2131 );
and \U$2230 ( \2355 , \2132 , \2135 );
or \U$2231 ( \2356 , \2354 , \2355 );
xor \U$2232 ( \2357 , \2353 , \2356 );
and \U$2233 ( \2358 , \1717 , \1371 );
xor \U$2234 ( \2359 , \2357 , \2358 );
and \U$2235 ( \2360 , \2136 , \2137 );
and \U$2236 ( \2361 , \2138 , \2141 );
or \U$2237 ( \2362 , \2360 , \2361 );
xor \U$2238 ( \2363 , \2359 , \2362 );
and \U$2239 ( \2364 , \1532 , \1550 );
xor \U$2240 ( \2365 , \2363 , \2364 );
and \U$2241 ( \2366 , \2142 , \2143 );
and \U$2242 ( \2367 , \2144 , \2147 );
or \U$2243 ( \2368 , \2366 , \2367 );
xor \U$2244 ( \2369 , \2365 , \2368 );
and \U$2245 ( \2370 , \1359 , \1741 );
xor \U$2246 ( \2371 , \2369 , \2370 );
and \U$2247 ( \2372 , \2148 , \2149 );
and \U$2248 ( \2373 , \2150 , \2153 );
or \U$2249 ( \2374 , \2372 , \2373 );
xor \U$2250 ( \2375 , \2371 , \2374 );
and \U$2251 ( \2376 , \1198 , \1944 );
xor \U$2252 ( \2377 , \2375 , \2376 );
and \U$2253 ( \2378 , \2154 , \2155 );
and \U$2254 ( \2379 , \2156 , \2157 );
or \U$2255 ( \2380 , \2378 , \2379 );
xor \U$2256 ( \2381 , \2377 , \2380 );
and \U$2257 ( \2382 , \960 , \2159 );
xor \U$2258 ( \2383 , \2381 , \2382 );
and \U$2259 ( \2384 , \2158 , \2160 );
xor \U$2260 ( \2385 , \2383 , \2384 );
buf \U$2261 ( \2386 , RI892a108_56);
and \U$2262 ( \2387 , \963 , \2386 );
xor \U$2263 ( \2388 , \2385 , \2387 );
buf \U$2264 ( \2389 , \2388 );
and \U$2265 ( \2390 , \2389 , \930 );
buf \U$2266 ( \2391 , RI8929208_24);
buf \U$2267 ( \2392 , RI892a108_56);
xor \U$2268 ( \2393 , \2391 , \2392 );
and \U$2269 ( \2394 , \2164 , \2165 );
and \U$2270 ( \2395 , \2165 , \2170 );
and \U$2271 ( \2396 , \2164 , \2170 );
or \U$2272 ( \2397 , \2394 , \2395 , \2396 );
xor \U$2273 ( \2398 , \2393 , \2397 );
buf \U$2274 ( \2399 , \2398 );
and \U$2275 ( \2400 , \2399 , \928 );
buf \U$2276 ( \2401 , RI8928a88_8);
buf \U$2277 ( \2402 , RI8929988_40);
xor \U$2278 ( \2403 , \2401 , \2402 );
and \U$2279 ( \2404 , \2174 , \2175 );
and \U$2280 ( \2405 , \2175 , \2180 );
and \U$2281 ( \2406 , \2174 , \2180 );
or \U$2282 ( \2407 , \2404 , \2405 , \2406 );
xor \U$2283 ( \2408 , \2403 , \2407 );
buf \U$2284 ( \2409 , \2408 );
and \U$2285 ( \2410 , \2409 , \926 );
and \U$2286 ( \2411 , RI892a108_56, \924 );
and \U$2287 ( \2412 , RI8929988_40, \922 );
and \U$2288 ( \2413 , RI8929208_24, \920 );
and \U$2289 ( \2414 , RI8928a88_8, \918 );
or \U$2290 ( \2415 , \2288_nG8e4 , \2290 , \2292 , \2294 , \2296 , \2343 , \2390 , \2400 , \2410 , \2411 , \2412 , \2413 , \2414 );
buf \U$2291 ( \2416 , \2415 );
and \U$2292 ( \2417 , \220 , \2416 );
and \U$2293 ( \2418 , \2287 , \2417 );
xor \U$2294 ( \2419 , \2287 , \2417 );
xor \U$2295 ( \2420 , \2192 , \2285 );
and \U$2296 ( \2421 , \1025 , \2416 );
and \U$2297 ( \2422 , \2420 , \2421 );
xor \U$2298 ( \2423 , \2420 , \2421 );
xor \U$2299 ( \2424 , \2196 , \2283 );
and \U$2300 ( \2425 , \1033 , \2416 );
and \U$2301 ( \2426 , \2424 , \2425 );
xor \U$2302 ( \2427 , \2424 , \2425 );
xor \U$2303 ( \2428 , \2200 , \2281 );
and \U$2304 ( \2429 , \1041 , \2416 );
and \U$2305 ( \2430 , \2428 , \2429 );
xor \U$2306 ( \2431 , \2428 , \2429 );
xor \U$2307 ( \2432 , \2204 , \2279 );
and \U$2308 ( \2433 , \1049 , \2416 );
and \U$2309 ( \2434 , \2432 , \2433 );
xor \U$2310 ( \2435 , \2432 , \2433 );
xor \U$2311 ( \2436 , \2208 , \2277 );
and \U$2312 ( \2437 , \1057 , \2416 );
and \U$2313 ( \2438 , \2436 , \2437 );
xor \U$2314 ( \2439 , \2436 , \2437 );
xor \U$2315 ( \2440 , \2212 , \2275 );
and \U$2316 ( \2441 , \1065 , \2416 );
and \U$2317 ( \2442 , \2440 , \2441 );
xor \U$2318 ( \2443 , \2440 , \2441 );
xor \U$2319 ( \2444 , \2216 , \2273 );
and \U$2320 ( \2445 , \1073 , \2416 );
and \U$2321 ( \2446 , \2444 , \2445 );
xor \U$2322 ( \2447 , \2444 , \2445 );
xor \U$2323 ( \2448 , \2220 , \2271 );
and \U$2324 ( \2449 , \1081 , \2416 );
and \U$2325 ( \2450 , \2448 , \2449 );
xor \U$2326 ( \2451 , \2448 , \2449 );
xor \U$2327 ( \2452 , \2224 , \2269 );
and \U$2328 ( \2453 , \1089 , \2416 );
and \U$2329 ( \2454 , \2452 , \2453 );
xor \U$2330 ( \2455 , \2452 , \2453 );
xor \U$2331 ( \2456 , \2228 , \2267 );
and \U$2332 ( \2457 , \1097 , \2416 );
and \U$2333 ( \2458 , \2456 , \2457 );
xor \U$2334 ( \2459 , \2456 , \2457 );
xor \U$2335 ( \2460 , \2232 , \2265 );
and \U$2336 ( \2461 , \1105 , \2416 );
and \U$2337 ( \2462 , \2460 , \2461 );
xor \U$2338 ( \2463 , \2460 , \2461 );
xor \U$2339 ( \2464 , \2236 , \2263 );
and \U$2340 ( \2465 , \1113 , \2416 );
and \U$2341 ( \2466 , \2464 , \2465 );
xor \U$2342 ( \2467 , \2464 , \2465 );
xor \U$2343 ( \2468 , \2240 , \2261 );
and \U$2344 ( \2469 , \1121 , \2416 );
and \U$2345 ( \2470 , \2468 , \2469 );
xor \U$2346 ( \2471 , \2468 , \2469 );
xor \U$2347 ( \2472 , \2244 , \2259 );
and \U$2348 ( \2473 , \1129 , \2416 );
and \U$2349 ( \2474 , \2472 , \2473 );
xor \U$2350 ( \2475 , \2472 , \2473 );
xor \U$2351 ( \2476 , \2248 , \2257 );
and \U$2352 ( \2477 , \1137 , \2416 );
and \U$2353 ( \2478 , \2476 , \2477 );
xor \U$2354 ( \2479 , \2476 , \2477 );
xor \U$2355 ( \2480 , \2252 , \2255 );
and \U$2356 ( \2481 , \1144 , \2416 );
and \U$2357 ( \2482 , \2480 , \2481 );
and \U$2358 ( \2483 , \2479 , \2482 );
or \U$2359 ( \2484 , \2478 , \2483 );
and \U$2360 ( \2485 , \2475 , \2484 );
or \U$2361 ( \2486 , \2474 , \2485 );
and \U$2362 ( \2487 , \2471 , \2486 );
or \U$2363 ( \2488 , \2470 , \2487 );
and \U$2364 ( \2489 , \2467 , \2488 );
or \U$2365 ( \2490 , \2466 , \2489 );
and \U$2366 ( \2491 , \2463 , \2490 );
or \U$2367 ( \2492 , \2462 , \2491 );
and \U$2368 ( \2493 , \2459 , \2492 );
or \U$2369 ( \2494 , \2458 , \2493 );
and \U$2370 ( \2495 , \2455 , \2494 );
or \U$2371 ( \2496 , \2454 , \2495 );
and \U$2372 ( \2497 , \2451 , \2496 );
or \U$2373 ( \2498 , \2450 , \2497 );
and \U$2374 ( \2499 , \2447 , \2498 );
or \U$2375 ( \2500 , \2446 , \2499 );
and \U$2376 ( \2501 , \2443 , \2500 );
or \U$2377 ( \2502 , \2442 , \2501 );
and \U$2378 ( \2503 , \2439 , \2502 );
or \U$2379 ( \2504 , \2438 , \2503 );
and \U$2380 ( \2505 , \2435 , \2504 );
or \U$2381 ( \2506 , \2434 , \2505 );
and \U$2382 ( \2507 , \2431 , \2506 );
or \U$2383 ( \2508 , \2430 , \2507 );
and \U$2384 ( \2509 , \2427 , \2508 );
or \U$2385 ( \2510 , \2426 , \2509 );
and \U$2386 ( \2511 , \2423 , \2510 );
or \U$2387 ( \2512 , \2422 , \2511 );
and \U$2388 ( \2513 , \2419 , \2512 );
or \U$2389 ( \2514 , \2418 , \2513 );
_DC g9c7 ( \2515_nG9c7 , 1'b0 , \941 );
or \U$2391 ( \2516 , RI8928a10_7, RI892a090_55);
and \U$2392 ( \2517 , \2516 , \940 );
and \U$2393 ( \2518 , RI8929190_23, RI8929910_39);
and \U$2394 ( \2519 , \2518 , \938 );
or \U$2395 ( \2520 , RI8928a10_7, RI8929190_23);
and \U$2396 ( \2521 , \2520 , \936 );
xor \U$2397 ( \2522 , RI8929910_39, RI892a090_55);
and \U$2398 ( \2523 , \2522 , \934 );
buf \U$2399 ( \2524 , RI8929190_23);
and \U$2400 ( \2525 , \2524 , \952 );
and \U$2401 ( \2526 , \2297 , \955 );
xor \U$2402 ( \2527 , \2525 , \2526 );
and \U$2403 ( \2528 , \2298 , \2299 );
and \U$2404 ( \2529 , \2300 , \2303 );
or \U$2405 ( \2530 , \2528 , \2529 );
xor \U$2406 ( \2531 , \2527 , \2530 );
and \U$2407 ( \2532 , \2082 , \1193 );
xor \U$2408 ( \2533 , \2531 , \2532 );
and \U$2409 ( \2534 , \2304 , \2305 );
and \U$2410 ( \2535 , \2306 , \2309 );
or \U$2411 ( \2536 , \2534 , \2535 );
xor \U$2412 ( \2537 , \2533 , \2536 );
and \U$2413 ( \2538 , \1879 , \1354 );
xor \U$2414 ( \2539 , \2537 , \2538 );
and \U$2415 ( \2540 , \2310 , \2311 );
and \U$2416 ( \2541 , \2312 , \2315 );
or \U$2417 ( \2542 , \2540 , \2541 );
xor \U$2418 ( \2543 , \2539 , \2542 );
and \U$2419 ( \2544 , \1688 , \1527 );
xor \U$2420 ( \2545 , \2543 , \2544 );
and \U$2421 ( \2546 , \2316 , \2317 );
and \U$2422 ( \2547 , \2318 , \2321 );
or \U$2423 ( \2548 , \2546 , \2547 );
xor \U$2424 ( \2549 , \2545 , \2548 );
and \U$2425 ( \2550 , \1509 , \1712 );
xor \U$2426 ( \2551 , \2549 , \2550 );
and \U$2427 ( \2552 , \2322 , \2323 );
and \U$2428 ( \2553 , \2324 , \2327 );
or \U$2429 ( \2554 , \2552 , \2553 );
xor \U$2430 ( \2555 , \2551 , \2554 );
and \U$2431 ( \2556 , \1342 , \1909 );
xor \U$2432 ( \2557 , \2555 , \2556 );
and \U$2433 ( \2558 , \2328 , \2329 );
and \U$2434 ( \2559 , \2330 , \2333 );
or \U$2435 ( \2560 , \2558 , \2559 );
xor \U$2436 ( \2561 , \2557 , \2560 );
and \U$2437 ( \2562 , \1187 , \2118 );
xor \U$2438 ( \2563 , \2561 , \2562 );
and \U$2439 ( \2564 , \2334 , \2335 );
and \U$2440 ( \2565 , \2336 , \2337 );
or \U$2441 ( \2566 , \2564 , \2565 );
xor \U$2442 ( \2567 , \2563 , \2566 );
and \U$2443 ( \2568 , \951 , \2339 );
xor \U$2444 ( \2569 , \2567 , \2568 );
and \U$2445 ( \2570 , \2338 , \2340 );
xor \U$2446 ( \2571 , \2569 , \2570 );
buf \U$2447 ( \2572 , RI8929910_39);
and \U$2448 ( \2573 , \954 , \2572 );
xor \U$2449 ( \2574 , \2571 , \2573 );
buf \U$2450 ( \2575 , \2574 );
and \U$2451 ( \2576 , \2575 , \932 );
buf \U$2452 ( \2577 , RI8928a10_7);
and \U$2453 ( \2578 , \2577 , \961 );
and \U$2454 ( \2579 , \2344 , \964 );
xor \U$2455 ( \2580 , \2578 , \2579 );
and \U$2456 ( \2581 , \2345 , \2346 );
and \U$2457 ( \2582 , \2347 , \2350 );
or \U$2458 ( \2583 , \2581 , \2582 );
xor \U$2459 ( \2584 , \2580 , \2583 );
and \U$2460 ( \2585 , \2123 , \1204 );
xor \U$2461 ( \2586 , \2584 , \2585 );
and \U$2462 ( \2587 , \2351 , \2352 );
and \U$2463 ( \2588 , \2353 , \2356 );
or \U$2464 ( \2589 , \2587 , \2588 );
xor \U$2465 ( \2590 , \2586 , \2589 );
and \U$2466 ( \2591 , \1914 , \1371 );
xor \U$2467 ( \2592 , \2590 , \2591 );
and \U$2468 ( \2593 , \2357 , \2358 );
and \U$2469 ( \2594 , \2359 , \2362 );
or \U$2470 ( \2595 , \2593 , \2594 );
xor \U$2471 ( \2596 , \2592 , \2595 );
and \U$2472 ( \2597 , \1717 , \1550 );
xor \U$2473 ( \2598 , \2596 , \2597 );
and \U$2474 ( \2599 , \2363 , \2364 );
and \U$2475 ( \2600 , \2365 , \2368 );
or \U$2476 ( \2601 , \2599 , \2600 );
xor \U$2477 ( \2602 , \2598 , \2601 );
and \U$2478 ( \2603 , \1532 , \1741 );
xor \U$2479 ( \2604 , \2602 , \2603 );
and \U$2480 ( \2605 , \2369 , \2370 );
and \U$2481 ( \2606 , \2371 , \2374 );
or \U$2482 ( \2607 , \2605 , \2606 );
xor \U$2483 ( \2608 , \2604 , \2607 );
and \U$2484 ( \2609 , \1359 , \1944 );
xor \U$2485 ( \2610 , \2608 , \2609 );
and \U$2486 ( \2611 , \2375 , \2376 );
and \U$2487 ( \2612 , \2377 , \2380 );
or \U$2488 ( \2613 , \2611 , \2612 );
xor \U$2489 ( \2614 , \2610 , \2613 );
and \U$2490 ( \2615 , \1198 , \2159 );
xor \U$2491 ( \2616 , \2614 , \2615 );
and \U$2492 ( \2617 , \2381 , \2382 );
and \U$2493 ( \2618 , \2383 , \2384 );
or \U$2494 ( \2619 , \2617 , \2618 );
xor \U$2495 ( \2620 , \2616 , \2619 );
and \U$2496 ( \2621 , \960 , \2386 );
xor \U$2497 ( \2622 , \2620 , \2621 );
and \U$2498 ( \2623 , \2385 , \2387 );
xor \U$2499 ( \2624 , \2622 , \2623 );
buf \U$2500 ( \2625 , RI892a090_55);
and \U$2501 ( \2626 , \963 , \2625 );
xor \U$2502 ( \2627 , \2624 , \2626 );
buf \U$2503 ( \2628 , \2627 );
and \U$2504 ( \2629 , \2628 , \930 );
buf \U$2505 ( \2630 , RI8929190_23);
buf \U$2506 ( \2631 , RI892a090_55);
xor \U$2507 ( \2632 , \2630 , \2631 );
and \U$2508 ( \2633 , \2391 , \2392 );
and \U$2509 ( \2634 , \2392 , \2397 );
and \U$2510 ( \2635 , \2391 , \2397 );
or \U$2511 ( \2636 , \2633 , \2634 , \2635 );
xor \U$2512 ( \2637 , \2632 , \2636 );
buf \U$2513 ( \2638 , \2637 );
and \U$2514 ( \2639 , \2638 , \928 );
buf \U$2515 ( \2640 , RI8928a10_7);
buf \U$2516 ( \2641 , RI8929910_39);
xor \U$2517 ( \2642 , \2640 , \2641 );
and \U$2518 ( \2643 , \2401 , \2402 );
and \U$2519 ( \2644 , \2402 , \2407 );
and \U$2520 ( \2645 , \2401 , \2407 );
or \U$2521 ( \2646 , \2643 , \2644 , \2645 );
xor \U$2522 ( \2647 , \2642 , \2646 );
buf \U$2523 ( \2648 , \2647 );
and \U$2524 ( \2649 , \2648 , \926 );
and \U$2525 ( \2650 , RI892a090_55, \924 );
and \U$2526 ( \2651 , RI8929910_39, \922 );
and \U$2527 ( \2652 , RI8929190_23, \920 );
and \U$2528 ( \2653 , RI8928a10_7, \918 );
or \U$2529 ( \2654 , \2515_nG9c7 , \2517 , \2519 , \2521 , \2523 , \2576 , \2629 , \2639 , \2649 , \2650 , \2651 , \2652 , \2653 );
buf \U$2530 ( \2655 , \2654 );
and \U$2531 ( \2656 , \220 , \2655 );
and \U$2532 ( \2657 , \2514 , \2656 );
xor \U$2533 ( \2658 , \2514 , \2656 );
xor \U$2534 ( \2659 , \2419 , \2512 );
and \U$2535 ( \2660 , \1025 , \2655 );
and \U$2536 ( \2661 , \2659 , \2660 );
xor \U$2537 ( \2662 , \2659 , \2660 );
xor \U$2538 ( \2663 , \2423 , \2510 );
and \U$2539 ( \2664 , \1033 , \2655 );
and \U$2540 ( \2665 , \2663 , \2664 );
xor \U$2541 ( \2666 , \2663 , \2664 );
xor \U$2542 ( \2667 , \2427 , \2508 );
and \U$2543 ( \2668 , \1041 , \2655 );
and \U$2544 ( \2669 , \2667 , \2668 );
xor \U$2545 ( \2670 , \2667 , \2668 );
xor \U$2546 ( \2671 , \2431 , \2506 );
and \U$2547 ( \2672 , \1049 , \2655 );
and \U$2548 ( \2673 , \2671 , \2672 );
xor \U$2549 ( \2674 , \2671 , \2672 );
xor \U$2550 ( \2675 , \2435 , \2504 );
and \U$2551 ( \2676 , \1057 , \2655 );
and \U$2552 ( \2677 , \2675 , \2676 );
xor \U$2553 ( \2678 , \2675 , \2676 );
xor \U$2554 ( \2679 , \2439 , \2502 );
and \U$2555 ( \2680 , \1065 , \2655 );
and \U$2556 ( \2681 , \2679 , \2680 );
xor \U$2557 ( \2682 , \2679 , \2680 );
xor \U$2558 ( \2683 , \2443 , \2500 );
and \U$2559 ( \2684 , \1073 , \2655 );
and \U$2560 ( \2685 , \2683 , \2684 );
xor \U$2561 ( \2686 , \2683 , \2684 );
xor \U$2562 ( \2687 , \2447 , \2498 );
and \U$2563 ( \2688 , \1081 , \2655 );
and \U$2564 ( \2689 , \2687 , \2688 );
xor \U$2565 ( \2690 , \2687 , \2688 );
xor \U$2566 ( \2691 , \2451 , \2496 );
and \U$2567 ( \2692 , \1089 , \2655 );
and \U$2568 ( \2693 , \2691 , \2692 );
xor \U$2569 ( \2694 , \2691 , \2692 );
xor \U$2570 ( \2695 , \2455 , \2494 );
and \U$2571 ( \2696 , \1097 , \2655 );
and \U$2572 ( \2697 , \2695 , \2696 );
xor \U$2573 ( \2698 , \2695 , \2696 );
xor \U$2574 ( \2699 , \2459 , \2492 );
and \U$2575 ( \2700 , \1105 , \2655 );
and \U$2576 ( \2701 , \2699 , \2700 );
xor \U$2577 ( \2702 , \2699 , \2700 );
xor \U$2578 ( \2703 , \2463 , \2490 );
and \U$2579 ( \2704 , \1113 , \2655 );
and \U$2580 ( \2705 , \2703 , \2704 );
xor \U$2581 ( \2706 , \2703 , \2704 );
xor \U$2582 ( \2707 , \2467 , \2488 );
and \U$2583 ( \2708 , \1121 , \2655 );
and \U$2584 ( \2709 , \2707 , \2708 );
xor \U$2585 ( \2710 , \2707 , \2708 );
xor \U$2586 ( \2711 , \2471 , \2486 );
and \U$2587 ( \2712 , \1129 , \2655 );
and \U$2588 ( \2713 , \2711 , \2712 );
xor \U$2589 ( \2714 , \2711 , \2712 );
xor \U$2590 ( \2715 , \2475 , \2484 );
and \U$2591 ( \2716 , \1137 , \2655 );
and \U$2592 ( \2717 , \2715 , \2716 );
xor \U$2593 ( \2718 , \2715 , \2716 );
xor \U$2594 ( \2719 , \2479 , \2482 );
and \U$2595 ( \2720 , \1144 , \2655 );
and \U$2596 ( \2721 , \2719 , \2720 );
and \U$2597 ( \2722 , \2718 , \2721 );
or \U$2598 ( \2723 , \2717 , \2722 );
and \U$2599 ( \2724 , \2714 , \2723 );
or \U$2600 ( \2725 , \2713 , \2724 );
and \U$2601 ( \2726 , \2710 , \2725 );
or \U$2602 ( \2727 , \2709 , \2726 );
and \U$2603 ( \2728 , \2706 , \2727 );
or \U$2604 ( \2729 , \2705 , \2728 );
and \U$2605 ( \2730 , \2702 , \2729 );
or \U$2606 ( \2731 , \2701 , \2730 );
and \U$2607 ( \2732 , \2698 , \2731 );
or \U$2608 ( \2733 , \2697 , \2732 );
and \U$2609 ( \2734 , \2694 , \2733 );
or \U$2610 ( \2735 , \2693 , \2734 );
and \U$2611 ( \2736 , \2690 , \2735 );
or \U$2612 ( \2737 , \2689 , \2736 );
and \U$2613 ( \2738 , \2686 , \2737 );
or \U$2614 ( \2739 , \2685 , \2738 );
and \U$2615 ( \2740 , \2682 , \2739 );
or \U$2616 ( \2741 , \2681 , \2740 );
and \U$2617 ( \2742 , \2678 , \2741 );
or \U$2618 ( \2743 , \2677 , \2742 );
and \U$2619 ( \2744 , \2674 , \2743 );
or \U$2620 ( \2745 , \2673 , \2744 );
and \U$2621 ( \2746 , \2670 , \2745 );
or \U$2622 ( \2747 , \2669 , \2746 );
and \U$2623 ( \2748 , \2666 , \2747 );
or \U$2624 ( \2749 , \2665 , \2748 );
and \U$2625 ( \2750 , \2662 , \2749 );
or \U$2626 ( \2751 , \2661 , \2750 );
and \U$2627 ( \2752 , \2658 , \2751 );
or \U$2628 ( \2753 , \2657 , \2752 );
_DC gab6 ( \2754_nGab6 , 1'b0 , \941 );
or \U$2630 ( \2755 , RI8928998_6, RI892a018_54);
and \U$2631 ( \2756 , \2755 , \940 );
and \U$2632 ( \2757 , RI8929118_22, RI8929898_38);
and \U$2633 ( \2758 , \2757 , \938 );
or \U$2634 ( \2759 , RI8928998_6, RI8929118_22);
and \U$2635 ( \2760 , \2759 , \936 );
xor \U$2636 ( \2761 , RI8929898_38, RI892a018_54);
and \U$2637 ( \2762 , \2761 , \934 );
buf \U$2638 ( \2763 , RI8929118_22);
and \U$2639 ( \2764 , \2763 , \952 );
and \U$2640 ( \2765 , \2524 , \955 );
xor \U$2641 ( \2766 , \2764 , \2765 );
and \U$2642 ( \2767 , \2525 , \2526 );
and \U$2643 ( \2768 , \2527 , \2530 );
or \U$2644 ( \2769 , \2767 , \2768 );
xor \U$2645 ( \2770 , \2766 , \2769 );
and \U$2646 ( \2771 , \2297 , \1193 );
xor \U$2647 ( \2772 , \2770 , \2771 );
and \U$2648 ( \2773 , \2531 , \2532 );
and \U$2649 ( \2774 , \2533 , \2536 );
or \U$2650 ( \2775 , \2773 , \2774 );
xor \U$2651 ( \2776 , \2772 , \2775 );
and \U$2652 ( \2777 , \2082 , \1354 );
xor \U$2653 ( \2778 , \2776 , \2777 );
and \U$2654 ( \2779 , \2537 , \2538 );
and \U$2655 ( \2780 , \2539 , \2542 );
or \U$2656 ( \2781 , \2779 , \2780 );
xor \U$2657 ( \2782 , \2778 , \2781 );
and \U$2658 ( \2783 , \1879 , \1527 );
xor \U$2659 ( \2784 , \2782 , \2783 );
and \U$2660 ( \2785 , \2543 , \2544 );
and \U$2661 ( \2786 , \2545 , \2548 );
or \U$2662 ( \2787 , \2785 , \2786 );
xor \U$2663 ( \2788 , \2784 , \2787 );
and \U$2664 ( \2789 , \1688 , \1712 );
xor \U$2665 ( \2790 , \2788 , \2789 );
and \U$2666 ( \2791 , \2549 , \2550 );
and \U$2667 ( \2792 , \2551 , \2554 );
or \U$2668 ( \2793 , \2791 , \2792 );
xor \U$2669 ( \2794 , \2790 , \2793 );
and \U$2670 ( \2795 , \1509 , \1909 );
xor \U$2671 ( \2796 , \2794 , \2795 );
and \U$2672 ( \2797 , \2555 , \2556 );
and \U$2673 ( \2798 , \2557 , \2560 );
or \U$2674 ( \2799 , \2797 , \2798 );
xor \U$2675 ( \2800 , \2796 , \2799 );
and \U$2676 ( \2801 , \1342 , \2118 );
xor \U$2677 ( \2802 , \2800 , \2801 );
and \U$2678 ( \2803 , \2561 , \2562 );
and \U$2679 ( \2804 , \2563 , \2566 );
or \U$2680 ( \2805 , \2803 , \2804 );
xor \U$2681 ( \2806 , \2802 , \2805 );
and \U$2682 ( \2807 , \1187 , \2339 );
xor \U$2683 ( \2808 , \2806 , \2807 );
and \U$2684 ( \2809 , \2567 , \2568 );
and \U$2685 ( \2810 , \2569 , \2570 );
or \U$2686 ( \2811 , \2809 , \2810 );
xor \U$2687 ( \2812 , \2808 , \2811 );
and \U$2688 ( \2813 , \951 , \2572 );
xor \U$2689 ( \2814 , \2812 , \2813 );
and \U$2690 ( \2815 , \2571 , \2573 );
xor \U$2691 ( \2816 , \2814 , \2815 );
buf \U$2692 ( \2817 , RI8929898_38);
and \U$2693 ( \2818 , \954 , \2817 );
xor \U$2694 ( \2819 , \2816 , \2818 );
buf \U$2695 ( \2820 , \2819 );
and \U$2696 ( \2821 , \2820 , \932 );
buf \U$2697 ( \2822 , RI8928998_6);
and \U$2698 ( \2823 , \2822 , \961 );
and \U$2699 ( \2824 , \2577 , \964 );
xor \U$2700 ( \2825 , \2823 , \2824 );
and \U$2701 ( \2826 , \2578 , \2579 );
and \U$2702 ( \2827 , \2580 , \2583 );
or \U$2703 ( \2828 , \2826 , \2827 );
xor \U$2704 ( \2829 , \2825 , \2828 );
and \U$2705 ( \2830 , \2344 , \1204 );
xor \U$2706 ( \2831 , \2829 , \2830 );
and \U$2707 ( \2832 , \2584 , \2585 );
and \U$2708 ( \2833 , \2586 , \2589 );
or \U$2709 ( \2834 , \2832 , \2833 );
xor \U$2710 ( \2835 , \2831 , \2834 );
and \U$2711 ( \2836 , \2123 , \1371 );
xor \U$2712 ( \2837 , \2835 , \2836 );
and \U$2713 ( \2838 , \2590 , \2591 );
and \U$2714 ( \2839 , \2592 , \2595 );
or \U$2715 ( \2840 , \2838 , \2839 );
xor \U$2716 ( \2841 , \2837 , \2840 );
and \U$2717 ( \2842 , \1914 , \1550 );
xor \U$2718 ( \2843 , \2841 , \2842 );
and \U$2719 ( \2844 , \2596 , \2597 );
and \U$2720 ( \2845 , \2598 , \2601 );
or \U$2721 ( \2846 , \2844 , \2845 );
xor \U$2722 ( \2847 , \2843 , \2846 );
and \U$2723 ( \2848 , \1717 , \1741 );
xor \U$2724 ( \2849 , \2847 , \2848 );
and \U$2725 ( \2850 , \2602 , \2603 );
and \U$2726 ( \2851 , \2604 , \2607 );
or \U$2727 ( \2852 , \2850 , \2851 );
xor \U$2728 ( \2853 , \2849 , \2852 );
and \U$2729 ( \2854 , \1532 , \1944 );
xor \U$2730 ( \2855 , \2853 , \2854 );
and \U$2731 ( \2856 , \2608 , \2609 );
and \U$2732 ( \2857 , \2610 , \2613 );
or \U$2733 ( \2858 , \2856 , \2857 );
xor \U$2734 ( \2859 , \2855 , \2858 );
and \U$2735 ( \2860 , \1359 , \2159 );
xor \U$2736 ( \2861 , \2859 , \2860 );
and \U$2737 ( \2862 , \2614 , \2615 );
and \U$2738 ( \2863 , \2616 , \2619 );
or \U$2739 ( \2864 , \2862 , \2863 );
xor \U$2740 ( \2865 , \2861 , \2864 );
and \U$2741 ( \2866 , \1198 , \2386 );
xor \U$2742 ( \2867 , \2865 , \2866 );
and \U$2743 ( \2868 , \2620 , \2621 );
and \U$2744 ( \2869 , \2622 , \2623 );
or \U$2745 ( \2870 , \2868 , \2869 );
xor \U$2746 ( \2871 , \2867 , \2870 );
and \U$2747 ( \2872 , \960 , \2625 );
xor \U$2748 ( \2873 , \2871 , \2872 );
and \U$2749 ( \2874 , \2624 , \2626 );
xor \U$2750 ( \2875 , \2873 , \2874 );
buf \U$2751 ( \2876 , RI892a018_54);
and \U$2752 ( \2877 , \963 , \2876 );
xor \U$2753 ( \2878 , \2875 , \2877 );
buf \U$2754 ( \2879 , \2878 );
and \U$2755 ( \2880 , \2879 , \930 );
buf \U$2756 ( \2881 , RI8929118_22);
buf \U$2757 ( \2882 , RI892a018_54);
xor \U$2758 ( \2883 , \2881 , \2882 );
and \U$2759 ( \2884 , \2630 , \2631 );
and \U$2760 ( \2885 , \2631 , \2636 );
and \U$2761 ( \2886 , \2630 , \2636 );
or \U$2762 ( \2887 , \2884 , \2885 , \2886 );
xor \U$2763 ( \2888 , \2883 , \2887 );
buf \U$2764 ( \2889 , \2888 );
and \U$2765 ( \2890 , \2889 , \928 );
buf \U$2766 ( \2891 , RI8928998_6);
buf \U$2767 ( \2892 , RI8929898_38);
xor \U$2768 ( \2893 , \2891 , \2892 );
and \U$2769 ( \2894 , \2640 , \2641 );
and \U$2770 ( \2895 , \2641 , \2646 );
and \U$2771 ( \2896 , \2640 , \2646 );
or \U$2772 ( \2897 , \2894 , \2895 , \2896 );
xor \U$2773 ( \2898 , \2893 , \2897 );
buf \U$2774 ( \2899 , \2898 );
and \U$2775 ( \2900 , \2899 , \926 );
and \U$2776 ( \2901 , RI892a018_54, \924 );
and \U$2777 ( \2902 , RI8929898_38, \922 );
and \U$2778 ( \2903 , RI8929118_22, \920 );
and \U$2779 ( \2904 , RI8928998_6, \918 );
or \U$2780 ( \2905 , \2754_nGab6 , \2756 , \2758 , \2760 , \2762 , \2821 , \2880 , \2890 , \2900 , \2901 , \2902 , \2903 , \2904 );
buf \U$2781 ( \2906 , \2905 );
and \U$2782 ( \2907 , \220 , \2906 );
and \U$2783 ( \2908 , \2753 , \2907 );
xor \U$2784 ( \2909 , \2753 , \2907 );
xor \U$2785 ( \2910 , \2658 , \2751 );
and \U$2786 ( \2911 , \1025 , \2906 );
and \U$2787 ( \2912 , \2910 , \2911 );
xor \U$2788 ( \2913 , \2910 , \2911 );
xor \U$2789 ( \2914 , \2662 , \2749 );
and \U$2790 ( \2915 , \1033 , \2906 );
and \U$2791 ( \2916 , \2914 , \2915 );
xor \U$2792 ( \2917 , \2914 , \2915 );
xor \U$2793 ( \2918 , \2666 , \2747 );
and \U$2794 ( \2919 , \1041 , \2906 );
and \U$2795 ( \2920 , \2918 , \2919 );
xor \U$2796 ( \2921 , \2918 , \2919 );
xor \U$2797 ( \2922 , \2670 , \2745 );
and \U$2798 ( \2923 , \1049 , \2906 );
and \U$2799 ( \2924 , \2922 , \2923 );
xor \U$2800 ( \2925 , \2922 , \2923 );
xor \U$2801 ( \2926 , \2674 , \2743 );
and \U$2802 ( \2927 , \1057 , \2906 );
and \U$2803 ( \2928 , \2926 , \2927 );
xor \U$2804 ( \2929 , \2926 , \2927 );
xor \U$2805 ( \2930 , \2678 , \2741 );
and \U$2806 ( \2931 , \1065 , \2906 );
and \U$2807 ( \2932 , \2930 , \2931 );
xor \U$2808 ( \2933 , \2930 , \2931 );
xor \U$2809 ( \2934 , \2682 , \2739 );
and \U$2810 ( \2935 , \1073 , \2906 );
and \U$2811 ( \2936 , \2934 , \2935 );
xor \U$2812 ( \2937 , \2934 , \2935 );
xor \U$2813 ( \2938 , \2686 , \2737 );
and \U$2814 ( \2939 , \1081 , \2906 );
and \U$2815 ( \2940 , \2938 , \2939 );
xor \U$2816 ( \2941 , \2938 , \2939 );
xor \U$2817 ( \2942 , \2690 , \2735 );
and \U$2818 ( \2943 , \1089 , \2906 );
and \U$2819 ( \2944 , \2942 , \2943 );
xor \U$2820 ( \2945 , \2942 , \2943 );
xor \U$2821 ( \2946 , \2694 , \2733 );
and \U$2822 ( \2947 , \1097 , \2906 );
and \U$2823 ( \2948 , \2946 , \2947 );
xor \U$2824 ( \2949 , \2946 , \2947 );
xor \U$2825 ( \2950 , \2698 , \2731 );
and \U$2826 ( \2951 , \1105 , \2906 );
and \U$2827 ( \2952 , \2950 , \2951 );
xor \U$2828 ( \2953 , \2950 , \2951 );
xor \U$2829 ( \2954 , \2702 , \2729 );
and \U$2830 ( \2955 , \1113 , \2906 );
and \U$2831 ( \2956 , \2954 , \2955 );
xor \U$2832 ( \2957 , \2954 , \2955 );
xor \U$2833 ( \2958 , \2706 , \2727 );
and \U$2834 ( \2959 , \1121 , \2906 );
and \U$2835 ( \2960 , \2958 , \2959 );
xor \U$2836 ( \2961 , \2958 , \2959 );
xor \U$2837 ( \2962 , \2710 , \2725 );
and \U$2838 ( \2963 , \1129 , \2906 );
and \U$2839 ( \2964 , \2962 , \2963 );
xor \U$2840 ( \2965 , \2962 , \2963 );
xor \U$2841 ( \2966 , \2714 , \2723 );
and \U$2842 ( \2967 , \1137 , \2906 );
and \U$2843 ( \2968 , \2966 , \2967 );
xor \U$2844 ( \2969 , \2966 , \2967 );
xor \U$2845 ( \2970 , \2718 , \2721 );
and \U$2846 ( \2971 , \1144 , \2906 );
and \U$2847 ( \2972 , \2970 , \2971 );
and \U$2848 ( \2973 , \2969 , \2972 );
or \U$2849 ( \2974 , \2968 , \2973 );
and \U$2850 ( \2975 , \2965 , \2974 );
or \U$2851 ( \2976 , \2964 , \2975 );
and \U$2852 ( \2977 , \2961 , \2976 );
or \U$2853 ( \2978 , \2960 , \2977 );
and \U$2854 ( \2979 , \2957 , \2978 );
or \U$2855 ( \2980 , \2956 , \2979 );
and \U$2856 ( \2981 , \2953 , \2980 );
or \U$2857 ( \2982 , \2952 , \2981 );
and \U$2858 ( \2983 , \2949 , \2982 );
or \U$2859 ( \2984 , \2948 , \2983 );
and \U$2860 ( \2985 , \2945 , \2984 );
or \U$2861 ( \2986 , \2944 , \2985 );
and \U$2862 ( \2987 , \2941 , \2986 );
or \U$2863 ( \2988 , \2940 , \2987 );
and \U$2864 ( \2989 , \2937 , \2988 );
or \U$2865 ( \2990 , \2936 , \2989 );
and \U$2866 ( \2991 , \2933 , \2990 );
or \U$2867 ( \2992 , \2932 , \2991 );
and \U$2868 ( \2993 , \2929 , \2992 );
or \U$2869 ( \2994 , \2928 , \2993 );
and \U$2870 ( \2995 , \2925 , \2994 );
or \U$2871 ( \2996 , \2924 , \2995 );
and \U$2872 ( \2997 , \2921 , \2996 );
or \U$2873 ( \2998 , \2920 , \2997 );
and \U$2874 ( \2999 , \2917 , \2998 );
or \U$2875 ( \3000 , \2916 , \2999 );
and \U$2876 ( \3001 , \2913 , \3000 );
or \U$2877 ( \3002 , \2912 , \3001 );
and \U$2878 ( \3003 , \2909 , \3002 );
or \U$2879 ( \3004 , \2908 , \3003 );
_DC gbb1 ( \3005_nGbb1 , 1'b0 , \941 );
or \U$2881 ( \3006 , RI8928920_5, RI8929fa0_53);
and \U$2882 ( \3007 , \3006 , \940 );
and \U$2883 ( \3008 , RI89290a0_21, RI8929820_37);
and \U$2884 ( \3009 , \3008 , \938 );
or \U$2885 ( \3010 , RI8928920_5, RI89290a0_21);
and \U$2886 ( \3011 , \3010 , \936 );
xor \U$2887 ( \3012 , RI8929820_37, RI8929fa0_53);
and \U$2888 ( \3013 , \3012 , \934 );
buf \U$2889 ( \3014 , RI89290a0_21);
and \U$2890 ( \3015 , \3014 , \952 );
and \U$2891 ( \3016 , \2763 , \955 );
xor \U$2892 ( \3017 , \3015 , \3016 );
and \U$2893 ( \3018 , \2764 , \2765 );
and \U$2894 ( \3019 , \2766 , \2769 );
or \U$2895 ( \3020 , \3018 , \3019 );
xor \U$2896 ( \3021 , \3017 , \3020 );
and \U$2897 ( \3022 , \2524 , \1193 );
xor \U$2898 ( \3023 , \3021 , \3022 );
and \U$2899 ( \3024 , \2770 , \2771 );
and \U$2900 ( \3025 , \2772 , \2775 );
or \U$2901 ( \3026 , \3024 , \3025 );
xor \U$2902 ( \3027 , \3023 , \3026 );
and \U$2903 ( \3028 , \2297 , \1354 );
xor \U$2904 ( \3029 , \3027 , \3028 );
and \U$2905 ( \3030 , \2776 , \2777 );
and \U$2906 ( \3031 , \2778 , \2781 );
or \U$2907 ( \3032 , \3030 , \3031 );
xor \U$2908 ( \3033 , \3029 , \3032 );
and \U$2909 ( \3034 , \2082 , \1527 );
xor \U$2910 ( \3035 , \3033 , \3034 );
and \U$2911 ( \3036 , \2782 , \2783 );
and \U$2912 ( \3037 , \2784 , \2787 );
or \U$2913 ( \3038 , \3036 , \3037 );
xor \U$2914 ( \3039 , \3035 , \3038 );
and \U$2915 ( \3040 , \1879 , \1712 );
xor \U$2916 ( \3041 , \3039 , \3040 );
and \U$2917 ( \3042 , \2788 , \2789 );
and \U$2918 ( \3043 , \2790 , \2793 );
or \U$2919 ( \3044 , \3042 , \3043 );
xor \U$2920 ( \3045 , \3041 , \3044 );
and \U$2921 ( \3046 , \1688 , \1909 );
xor \U$2922 ( \3047 , \3045 , \3046 );
and \U$2923 ( \3048 , \2794 , \2795 );
and \U$2924 ( \3049 , \2796 , \2799 );
or \U$2925 ( \3050 , \3048 , \3049 );
xor \U$2926 ( \3051 , \3047 , \3050 );
and \U$2927 ( \3052 , \1509 , \2118 );
xor \U$2928 ( \3053 , \3051 , \3052 );
and \U$2929 ( \3054 , \2800 , \2801 );
and \U$2930 ( \3055 , \2802 , \2805 );
or \U$2931 ( \3056 , \3054 , \3055 );
xor \U$2932 ( \3057 , \3053 , \3056 );
and \U$2933 ( \3058 , \1342 , \2339 );
xor \U$2934 ( \3059 , \3057 , \3058 );
and \U$2935 ( \3060 , \2806 , \2807 );
and \U$2936 ( \3061 , \2808 , \2811 );
or \U$2937 ( \3062 , \3060 , \3061 );
xor \U$2938 ( \3063 , \3059 , \3062 );
and \U$2939 ( \3064 , \1187 , \2572 );
xor \U$2940 ( \3065 , \3063 , \3064 );
and \U$2941 ( \3066 , \2812 , \2813 );
and \U$2942 ( \3067 , \2814 , \2815 );
or \U$2943 ( \3068 , \3066 , \3067 );
xor \U$2944 ( \3069 , \3065 , \3068 );
and \U$2945 ( \3070 , \951 , \2817 );
xor \U$2946 ( \3071 , \3069 , \3070 );
and \U$2947 ( \3072 , \2816 , \2818 );
xor \U$2948 ( \3073 , \3071 , \3072 );
buf \U$2949 ( \3074 , RI8929820_37);
and \U$2950 ( \3075 , \954 , \3074 );
xor \U$2951 ( \3076 , \3073 , \3075 );
buf \U$2952 ( \3077 , \3076 );
and \U$2953 ( \3078 , \3077 , \932 );
buf \U$2954 ( \3079 , RI8928920_5);
and \U$2955 ( \3080 , \3079 , \961 );
and \U$2956 ( \3081 , \2822 , \964 );
xor \U$2957 ( \3082 , \3080 , \3081 );
and \U$2958 ( \3083 , \2823 , \2824 );
and \U$2959 ( \3084 , \2825 , \2828 );
or \U$2960 ( \3085 , \3083 , \3084 );
xor \U$2961 ( \3086 , \3082 , \3085 );
and \U$2962 ( \3087 , \2577 , \1204 );
xor \U$2963 ( \3088 , \3086 , \3087 );
and \U$2964 ( \3089 , \2829 , \2830 );
and \U$2965 ( \3090 , \2831 , \2834 );
or \U$2966 ( \3091 , \3089 , \3090 );
xor \U$2967 ( \3092 , \3088 , \3091 );
and \U$2968 ( \3093 , \2344 , \1371 );
xor \U$2969 ( \3094 , \3092 , \3093 );
and \U$2970 ( \3095 , \2835 , \2836 );
and \U$2971 ( \3096 , \2837 , \2840 );
or \U$2972 ( \3097 , \3095 , \3096 );
xor \U$2973 ( \3098 , \3094 , \3097 );
and \U$2974 ( \3099 , \2123 , \1550 );
xor \U$2975 ( \3100 , \3098 , \3099 );
and \U$2976 ( \3101 , \2841 , \2842 );
and \U$2977 ( \3102 , \2843 , \2846 );
or \U$2978 ( \3103 , \3101 , \3102 );
xor \U$2979 ( \3104 , \3100 , \3103 );
and \U$2980 ( \3105 , \1914 , \1741 );
xor \U$2981 ( \3106 , \3104 , \3105 );
and \U$2982 ( \3107 , \2847 , \2848 );
and \U$2983 ( \3108 , \2849 , \2852 );
or \U$2984 ( \3109 , \3107 , \3108 );
xor \U$2985 ( \3110 , \3106 , \3109 );
and \U$2986 ( \3111 , \1717 , \1944 );
xor \U$2987 ( \3112 , \3110 , \3111 );
and \U$2988 ( \3113 , \2853 , \2854 );
and \U$2989 ( \3114 , \2855 , \2858 );
or \U$2990 ( \3115 , \3113 , \3114 );
xor \U$2991 ( \3116 , \3112 , \3115 );
and \U$2992 ( \3117 , \1532 , \2159 );
xor \U$2993 ( \3118 , \3116 , \3117 );
and \U$2994 ( \3119 , \2859 , \2860 );
and \U$2995 ( \3120 , \2861 , \2864 );
or \U$2996 ( \3121 , \3119 , \3120 );
xor \U$2997 ( \3122 , \3118 , \3121 );
and \U$2998 ( \3123 , \1359 , \2386 );
xor \U$2999 ( \3124 , \3122 , \3123 );
and \U$3000 ( \3125 , \2865 , \2866 );
and \U$3001 ( \3126 , \2867 , \2870 );
or \U$3002 ( \3127 , \3125 , \3126 );
xor \U$3003 ( \3128 , \3124 , \3127 );
and \U$3004 ( \3129 , \1198 , \2625 );
xor \U$3005 ( \3130 , \3128 , \3129 );
and \U$3006 ( \3131 , \2871 , \2872 );
and \U$3007 ( \3132 , \2873 , \2874 );
or \U$3008 ( \3133 , \3131 , \3132 );
xor \U$3009 ( \3134 , \3130 , \3133 );
and \U$3010 ( \3135 , \960 , \2876 );
xor \U$3011 ( \3136 , \3134 , \3135 );
and \U$3012 ( \3137 , \2875 , \2877 );
xor \U$3013 ( \3138 , \3136 , \3137 );
buf \U$3014 ( \3139 , RI8929fa0_53);
and \U$3015 ( \3140 , \963 , \3139 );
xor \U$3016 ( \3141 , \3138 , \3140 );
buf \U$3017 ( \3142 , \3141 );
and \U$3018 ( \3143 , \3142 , \930 );
buf \U$3019 ( \3144 , RI89290a0_21);
buf \U$3020 ( \3145 , RI8929fa0_53);
xor \U$3021 ( \3146 , \3144 , \3145 );
and \U$3022 ( \3147 , \2881 , \2882 );
and \U$3023 ( \3148 , \2882 , \2887 );
and \U$3024 ( \3149 , \2881 , \2887 );
or \U$3025 ( \3150 , \3147 , \3148 , \3149 );
xor \U$3026 ( \3151 , \3146 , \3150 );
buf \U$3027 ( \3152 , \3151 );
and \U$3028 ( \3153 , \3152 , \928 );
buf \U$3029 ( \3154 , RI8928920_5);
buf \U$3030 ( \3155 , RI8929820_37);
xor \U$3031 ( \3156 , \3154 , \3155 );
and \U$3032 ( \3157 , \2891 , \2892 );
and \U$3033 ( \3158 , \2892 , \2897 );
and \U$3034 ( \3159 , \2891 , \2897 );
or \U$3035 ( \3160 , \3157 , \3158 , \3159 );
xor \U$3036 ( \3161 , \3156 , \3160 );
buf \U$3037 ( \3162 , \3161 );
and \U$3038 ( \3163 , \3162 , \926 );
and \U$3039 ( \3164 , RI8929fa0_53, \924 );
and \U$3040 ( \3165 , RI8929820_37, \922 );
and \U$3041 ( \3166 , RI89290a0_21, \920 );
and \U$3042 ( \3167 , RI8928920_5, \918 );
or \U$3043 ( \3168 , \3005_nGbb1 , \3007 , \3009 , \3011 , \3013 , \3078 , \3143 , \3153 , \3163 , \3164 , \3165 , \3166 , \3167 );
buf \U$3044 ( \3169 , \3168 );
and \U$3045 ( \3170 , \220 , \3169 );
and \U$3046 ( \3171 , \3004 , \3170 );
xor \U$3047 ( \3172 , \3004 , \3170 );
xor \U$3048 ( \3173 , \2909 , \3002 );
and \U$3049 ( \3174 , \1025 , \3169 );
and \U$3050 ( \3175 , \3173 , \3174 );
xor \U$3051 ( \3176 , \3173 , \3174 );
xor \U$3052 ( \3177 , \2913 , \3000 );
and \U$3053 ( \3178 , \1033 , \3169 );
and \U$3054 ( \3179 , \3177 , \3178 );
xor \U$3055 ( \3180 , \3177 , \3178 );
xor \U$3056 ( \3181 , \2917 , \2998 );
and \U$3057 ( \3182 , \1041 , \3169 );
and \U$3058 ( \3183 , \3181 , \3182 );
xor \U$3059 ( \3184 , \3181 , \3182 );
xor \U$3060 ( \3185 , \2921 , \2996 );
and \U$3061 ( \3186 , \1049 , \3169 );
and \U$3062 ( \3187 , \3185 , \3186 );
xor \U$3063 ( \3188 , \3185 , \3186 );
xor \U$3064 ( \3189 , \2925 , \2994 );
and \U$3065 ( \3190 , \1057 , \3169 );
and \U$3066 ( \3191 , \3189 , \3190 );
xor \U$3067 ( \3192 , \3189 , \3190 );
xor \U$3068 ( \3193 , \2929 , \2992 );
and \U$3069 ( \3194 , \1065 , \3169 );
and \U$3070 ( \3195 , \3193 , \3194 );
xor \U$3071 ( \3196 , \3193 , \3194 );
xor \U$3072 ( \3197 , \2933 , \2990 );
and \U$3073 ( \3198 , \1073 , \3169 );
and \U$3074 ( \3199 , \3197 , \3198 );
xor \U$3075 ( \3200 , \3197 , \3198 );
xor \U$3076 ( \3201 , \2937 , \2988 );
and \U$3077 ( \3202 , \1081 , \3169 );
and \U$3078 ( \3203 , \3201 , \3202 );
xor \U$3079 ( \3204 , \3201 , \3202 );
xor \U$3080 ( \3205 , \2941 , \2986 );
and \U$3081 ( \3206 , \1089 , \3169 );
and \U$3082 ( \3207 , \3205 , \3206 );
xor \U$3083 ( \3208 , \3205 , \3206 );
xor \U$3084 ( \3209 , \2945 , \2984 );
and \U$3085 ( \3210 , \1097 , \3169 );
and \U$3086 ( \3211 , \3209 , \3210 );
xor \U$3087 ( \3212 , \3209 , \3210 );
xor \U$3088 ( \3213 , \2949 , \2982 );
and \U$3089 ( \3214 , \1105 , \3169 );
and \U$3090 ( \3215 , \3213 , \3214 );
xor \U$3091 ( \3216 , \3213 , \3214 );
xor \U$3092 ( \3217 , \2953 , \2980 );
and \U$3093 ( \3218 , \1113 , \3169 );
and \U$3094 ( \3219 , \3217 , \3218 );
xor \U$3095 ( \3220 , \3217 , \3218 );
xor \U$3096 ( \3221 , \2957 , \2978 );
and \U$3097 ( \3222 , \1121 , \3169 );
and \U$3098 ( \3223 , \3221 , \3222 );
xor \U$3099 ( \3224 , \3221 , \3222 );
xor \U$3100 ( \3225 , \2961 , \2976 );
and \U$3101 ( \3226 , \1129 , \3169 );
and \U$3102 ( \3227 , \3225 , \3226 );
xor \U$3103 ( \3228 , \3225 , \3226 );
xor \U$3104 ( \3229 , \2965 , \2974 );
and \U$3105 ( \3230 , \1137 , \3169 );
and \U$3106 ( \3231 , \3229 , \3230 );
xor \U$3107 ( \3232 , \3229 , \3230 );
xor \U$3108 ( \3233 , \2969 , \2972 );
and \U$3109 ( \3234 , \1144 , \3169 );
and \U$3110 ( \3235 , \3233 , \3234 );
and \U$3111 ( \3236 , \3232 , \3235 );
or \U$3112 ( \3237 , \3231 , \3236 );
and \U$3113 ( \3238 , \3228 , \3237 );
or \U$3114 ( \3239 , \3227 , \3238 );
and \U$3115 ( \3240 , \3224 , \3239 );
or \U$3116 ( \3241 , \3223 , \3240 );
and \U$3117 ( \3242 , \3220 , \3241 );
or \U$3118 ( \3243 , \3219 , \3242 );
and \U$3119 ( \3244 , \3216 , \3243 );
or \U$3120 ( \3245 , \3215 , \3244 );
and \U$3121 ( \3246 , \3212 , \3245 );
or \U$3122 ( \3247 , \3211 , \3246 );
and \U$3123 ( \3248 , \3208 , \3247 );
or \U$3124 ( \3249 , \3207 , \3248 );
and \U$3125 ( \3250 , \3204 , \3249 );
or \U$3126 ( \3251 , \3203 , \3250 );
and \U$3127 ( \3252 , \3200 , \3251 );
or \U$3128 ( \3253 , \3199 , \3252 );
and \U$3129 ( \3254 , \3196 , \3253 );
or \U$3130 ( \3255 , \3195 , \3254 );
and \U$3131 ( \3256 , \3192 , \3255 );
or \U$3132 ( \3257 , \3191 , \3256 );
and \U$3133 ( \3258 , \3188 , \3257 );
or \U$3134 ( \3259 , \3187 , \3258 );
and \U$3135 ( \3260 , \3184 , \3259 );
or \U$3136 ( \3261 , \3183 , \3260 );
and \U$3137 ( \3262 , \3180 , \3261 );
or \U$3138 ( \3263 , \3179 , \3262 );
and \U$3139 ( \3264 , \3176 , \3263 );
or \U$3140 ( \3265 , \3175 , \3264 );
and \U$3141 ( \3266 , \3172 , \3265 );
or \U$3142 ( \3267 , \3171 , \3266 );
_DC gcb8 ( \3268_nGcb8 , 1'b0 , \941 );
or \U$3144 ( \3269 , RI89288a8_4, RI8929f28_52);
and \U$3145 ( \3270 , \3269 , \940 );
and \U$3146 ( \3271 , RI8929028_20, RI89297a8_36);
and \U$3147 ( \3272 , \3271 , \938 );
or \U$3148 ( \3273 , RI89288a8_4, RI8929028_20);
and \U$3149 ( \3274 , \3273 , \936 );
xor \U$3150 ( \3275 , RI89297a8_36, RI8929f28_52);
and \U$3151 ( \3276 , \3275 , \934 );
buf \U$3152 ( \3277 , RI8929028_20);
and \U$3153 ( \3278 , \3277 , \952 );
and \U$3154 ( \3279 , \3014 , \955 );
xor \U$3155 ( \3280 , \3278 , \3279 );
and \U$3156 ( \3281 , \3015 , \3016 );
and \U$3157 ( \3282 , \3017 , \3020 );
or \U$3158 ( \3283 , \3281 , \3282 );
xor \U$3159 ( \3284 , \3280 , \3283 );
and \U$3160 ( \3285 , \2763 , \1193 );
xor \U$3161 ( \3286 , \3284 , \3285 );
and \U$3162 ( \3287 , \3021 , \3022 );
and \U$3163 ( \3288 , \3023 , \3026 );
or \U$3164 ( \3289 , \3287 , \3288 );
xor \U$3165 ( \3290 , \3286 , \3289 );
and \U$3166 ( \3291 , \2524 , \1354 );
xor \U$3167 ( \3292 , \3290 , \3291 );
and \U$3168 ( \3293 , \3027 , \3028 );
and \U$3169 ( \3294 , \3029 , \3032 );
or \U$3170 ( \3295 , \3293 , \3294 );
xor \U$3171 ( \3296 , \3292 , \3295 );
and \U$3172 ( \3297 , \2297 , \1527 );
xor \U$3173 ( \3298 , \3296 , \3297 );
and \U$3174 ( \3299 , \3033 , \3034 );
and \U$3175 ( \3300 , \3035 , \3038 );
or \U$3176 ( \3301 , \3299 , \3300 );
xor \U$3177 ( \3302 , \3298 , \3301 );
and \U$3178 ( \3303 , \2082 , \1712 );
xor \U$3179 ( \3304 , \3302 , \3303 );
and \U$3180 ( \3305 , \3039 , \3040 );
and \U$3181 ( \3306 , \3041 , \3044 );
or \U$3182 ( \3307 , \3305 , \3306 );
xor \U$3183 ( \3308 , \3304 , \3307 );
and \U$3184 ( \3309 , \1879 , \1909 );
xor \U$3185 ( \3310 , \3308 , \3309 );
and \U$3186 ( \3311 , \3045 , \3046 );
and \U$3187 ( \3312 , \3047 , \3050 );
or \U$3188 ( \3313 , \3311 , \3312 );
xor \U$3189 ( \3314 , \3310 , \3313 );
and \U$3190 ( \3315 , \1688 , \2118 );
xor \U$3191 ( \3316 , \3314 , \3315 );
and \U$3192 ( \3317 , \3051 , \3052 );
and \U$3193 ( \3318 , \3053 , \3056 );
or \U$3194 ( \3319 , \3317 , \3318 );
xor \U$3195 ( \3320 , \3316 , \3319 );
and \U$3196 ( \3321 , \1509 , \2339 );
xor \U$3197 ( \3322 , \3320 , \3321 );
and \U$3198 ( \3323 , \3057 , \3058 );
and \U$3199 ( \3324 , \3059 , \3062 );
or \U$3200 ( \3325 , \3323 , \3324 );
xor \U$3201 ( \3326 , \3322 , \3325 );
and \U$3202 ( \3327 , \1342 , \2572 );
xor \U$3203 ( \3328 , \3326 , \3327 );
and \U$3204 ( \3329 , \3063 , \3064 );
and \U$3205 ( \3330 , \3065 , \3068 );
or \U$3206 ( \3331 , \3329 , \3330 );
xor \U$3207 ( \3332 , \3328 , \3331 );
and \U$3208 ( \3333 , \1187 , \2817 );
xor \U$3209 ( \3334 , \3332 , \3333 );
and \U$3210 ( \3335 , \3069 , \3070 );
and \U$3211 ( \3336 , \3071 , \3072 );
or \U$3212 ( \3337 , \3335 , \3336 );
xor \U$3213 ( \3338 , \3334 , \3337 );
and \U$3214 ( \3339 , \951 , \3074 );
xor \U$3215 ( \3340 , \3338 , \3339 );
and \U$3216 ( \3341 , \3073 , \3075 );
xor \U$3217 ( \3342 , \3340 , \3341 );
buf \U$3218 ( \3343 , RI89297a8_36);
and \U$3219 ( \3344 , \954 , \3343 );
xor \U$3220 ( \3345 , \3342 , \3344 );
buf \U$3221 ( \3346 , \3345 );
and \U$3222 ( \3347 , \3346 , \932 );
buf \U$3223 ( \3348 , RI89288a8_4);
and \U$3224 ( \3349 , \3348 , \961 );
and \U$3225 ( \3350 , \3079 , \964 );
xor \U$3226 ( \3351 , \3349 , \3350 );
and \U$3227 ( \3352 , \3080 , \3081 );
and \U$3228 ( \3353 , \3082 , \3085 );
or \U$3229 ( \3354 , \3352 , \3353 );
xor \U$3230 ( \3355 , \3351 , \3354 );
and \U$3231 ( \3356 , \2822 , \1204 );
xor \U$3232 ( \3357 , \3355 , \3356 );
and \U$3233 ( \3358 , \3086 , \3087 );
and \U$3234 ( \3359 , \3088 , \3091 );
or \U$3235 ( \3360 , \3358 , \3359 );
xor \U$3236 ( \3361 , \3357 , \3360 );
and \U$3237 ( \3362 , \2577 , \1371 );
xor \U$3238 ( \3363 , \3361 , \3362 );
and \U$3239 ( \3364 , \3092 , \3093 );
and \U$3240 ( \3365 , \3094 , \3097 );
or \U$3241 ( \3366 , \3364 , \3365 );
xor \U$3242 ( \3367 , \3363 , \3366 );
and \U$3243 ( \3368 , \2344 , \1550 );
xor \U$3244 ( \3369 , \3367 , \3368 );
and \U$3245 ( \3370 , \3098 , \3099 );
and \U$3246 ( \3371 , \3100 , \3103 );
or \U$3247 ( \3372 , \3370 , \3371 );
xor \U$3248 ( \3373 , \3369 , \3372 );
and \U$3249 ( \3374 , \2123 , \1741 );
xor \U$3250 ( \3375 , \3373 , \3374 );
and \U$3251 ( \3376 , \3104 , \3105 );
and \U$3252 ( \3377 , \3106 , \3109 );
or \U$3253 ( \3378 , \3376 , \3377 );
xor \U$3254 ( \3379 , \3375 , \3378 );
and \U$3255 ( \3380 , \1914 , \1944 );
xor \U$3256 ( \3381 , \3379 , \3380 );
and \U$3257 ( \3382 , \3110 , \3111 );
and \U$3258 ( \3383 , \3112 , \3115 );
or \U$3259 ( \3384 , \3382 , \3383 );
xor \U$3260 ( \3385 , \3381 , \3384 );
and \U$3261 ( \3386 , \1717 , \2159 );
xor \U$3262 ( \3387 , \3385 , \3386 );
and \U$3263 ( \3388 , \3116 , \3117 );
and \U$3264 ( \3389 , \3118 , \3121 );
or \U$3265 ( \3390 , \3388 , \3389 );
xor \U$3266 ( \3391 , \3387 , \3390 );
and \U$3267 ( \3392 , \1532 , \2386 );
xor \U$3268 ( \3393 , \3391 , \3392 );
and \U$3269 ( \3394 , \3122 , \3123 );
and \U$3270 ( \3395 , \3124 , \3127 );
or \U$3271 ( \3396 , \3394 , \3395 );
xor \U$3272 ( \3397 , \3393 , \3396 );
and \U$3273 ( \3398 , \1359 , \2625 );
xor \U$3274 ( \3399 , \3397 , \3398 );
and \U$3275 ( \3400 , \3128 , \3129 );
and \U$3276 ( \3401 , \3130 , \3133 );
or \U$3277 ( \3402 , \3400 , \3401 );
xor \U$3278 ( \3403 , \3399 , \3402 );
and \U$3279 ( \3404 , \1198 , \2876 );
xor \U$3280 ( \3405 , \3403 , \3404 );
and \U$3281 ( \3406 , \3134 , \3135 );
and \U$3282 ( \3407 , \3136 , \3137 );
or \U$3283 ( \3408 , \3406 , \3407 );
xor \U$3284 ( \3409 , \3405 , \3408 );
and \U$3285 ( \3410 , \960 , \3139 );
xor \U$3286 ( \3411 , \3409 , \3410 );
and \U$3287 ( \3412 , \3138 , \3140 );
xor \U$3288 ( \3413 , \3411 , \3412 );
buf \U$3289 ( \3414 , RI8929f28_52);
and \U$3290 ( \3415 , \963 , \3414 );
xor \U$3291 ( \3416 , \3413 , \3415 );
buf \U$3292 ( \3417 , \3416 );
and \U$3293 ( \3418 , \3417 , \930 );
buf \U$3294 ( \3419 , RI8929028_20);
buf \U$3295 ( \3420 , RI8929f28_52);
xor \U$3296 ( \3421 , \3419 , \3420 );
and \U$3297 ( \3422 , \3144 , \3145 );
and \U$3298 ( \3423 , \3145 , \3150 );
and \U$3299 ( \3424 , \3144 , \3150 );
or \U$3300 ( \3425 , \3422 , \3423 , \3424 );
xor \U$3301 ( \3426 , \3421 , \3425 );
buf \U$3302 ( \3427 , \3426 );
and \U$3303 ( \3428 , \3427 , \928 );
buf \U$3304 ( \3429 , RI89288a8_4);
buf \U$3305 ( \3430 , RI89297a8_36);
xor \U$3306 ( \3431 , \3429 , \3430 );
and \U$3307 ( \3432 , \3154 , \3155 );
and \U$3308 ( \3433 , \3155 , \3160 );
and \U$3309 ( \3434 , \3154 , \3160 );
or \U$3310 ( \3435 , \3432 , \3433 , \3434 );
xor \U$3311 ( \3436 , \3431 , \3435 );
buf \U$3312 ( \3437 , \3436 );
and \U$3313 ( \3438 , \3437 , \926 );
and \U$3314 ( \3439 , RI8929f28_52, \924 );
and \U$3315 ( \3440 , RI89297a8_36, \922 );
and \U$3316 ( \3441 , RI8929028_20, \920 );
and \U$3317 ( \3442 , RI89288a8_4, \918 );
or \U$3318 ( \3443 , \3268_nGcb8 , \3270 , \3272 , \3274 , \3276 , \3347 , \3418 , \3428 , \3438 , \3439 , \3440 , \3441 , \3442 );
buf \U$3319 ( \3444 , \3443 );
and \U$3320 ( \3445 , \220 , \3444 );
and \U$3321 ( \3446 , \3267 , \3445 );
xor \U$3322 ( \3447 , \3267 , \3445 );
xor \U$3323 ( \3448 , \3172 , \3265 );
and \U$3324 ( \3449 , \1025 , \3444 );
and \U$3325 ( \3450 , \3448 , \3449 );
xor \U$3326 ( \3451 , \3448 , \3449 );
xor \U$3327 ( \3452 , \3176 , \3263 );
and \U$3328 ( \3453 , \1033 , \3444 );
and \U$3329 ( \3454 , \3452 , \3453 );
xor \U$3330 ( \3455 , \3452 , \3453 );
xor \U$3331 ( \3456 , \3180 , \3261 );
and \U$3332 ( \3457 , \1041 , \3444 );
and \U$3333 ( \3458 , \3456 , \3457 );
xor \U$3334 ( \3459 , \3456 , \3457 );
xor \U$3335 ( \3460 , \3184 , \3259 );
and \U$3336 ( \3461 , \1049 , \3444 );
and \U$3337 ( \3462 , \3460 , \3461 );
xor \U$3338 ( \3463 , \3460 , \3461 );
xor \U$3339 ( \3464 , \3188 , \3257 );
and \U$3340 ( \3465 , \1057 , \3444 );
and \U$3341 ( \3466 , \3464 , \3465 );
xor \U$3342 ( \3467 , \3464 , \3465 );
xor \U$3343 ( \3468 , \3192 , \3255 );
and \U$3344 ( \3469 , \1065 , \3444 );
and \U$3345 ( \3470 , \3468 , \3469 );
xor \U$3346 ( \3471 , \3468 , \3469 );
xor \U$3347 ( \3472 , \3196 , \3253 );
and \U$3348 ( \3473 , \1073 , \3444 );
and \U$3349 ( \3474 , \3472 , \3473 );
xor \U$3350 ( \3475 , \3472 , \3473 );
xor \U$3351 ( \3476 , \3200 , \3251 );
and \U$3352 ( \3477 , \1081 , \3444 );
and \U$3353 ( \3478 , \3476 , \3477 );
xor \U$3354 ( \3479 , \3476 , \3477 );
xor \U$3355 ( \3480 , \3204 , \3249 );
and \U$3356 ( \3481 , \1089 , \3444 );
and \U$3357 ( \3482 , \3480 , \3481 );
xor \U$3358 ( \3483 , \3480 , \3481 );
xor \U$3359 ( \3484 , \3208 , \3247 );
and \U$3360 ( \3485 , \1097 , \3444 );
and \U$3361 ( \3486 , \3484 , \3485 );
xor \U$3362 ( \3487 , \3484 , \3485 );
xor \U$3363 ( \3488 , \3212 , \3245 );
and \U$3364 ( \3489 , \1105 , \3444 );
and \U$3365 ( \3490 , \3488 , \3489 );
xor \U$3366 ( \3491 , \3488 , \3489 );
xor \U$3367 ( \3492 , \3216 , \3243 );
and \U$3368 ( \3493 , \1113 , \3444 );
and \U$3369 ( \3494 , \3492 , \3493 );
xor \U$3370 ( \3495 , \3492 , \3493 );
xor \U$3371 ( \3496 , \3220 , \3241 );
and \U$3372 ( \3497 , \1121 , \3444 );
and \U$3373 ( \3498 , \3496 , \3497 );
xor \U$3374 ( \3499 , \3496 , \3497 );
xor \U$3375 ( \3500 , \3224 , \3239 );
and \U$3376 ( \3501 , \1129 , \3444 );
and \U$3377 ( \3502 , \3500 , \3501 );
xor \U$3378 ( \3503 , \3500 , \3501 );
xor \U$3379 ( \3504 , \3228 , \3237 );
and \U$3380 ( \3505 , \1137 , \3444 );
and \U$3381 ( \3506 , \3504 , \3505 );
xor \U$3382 ( \3507 , \3504 , \3505 );
xor \U$3383 ( \3508 , \3232 , \3235 );
and \U$3384 ( \3509 , \1144 , \3444 );
and \U$3385 ( \3510 , \3508 , \3509 );
and \U$3386 ( \3511 , \3507 , \3510 );
or \U$3387 ( \3512 , \3506 , \3511 );
and \U$3388 ( \3513 , \3503 , \3512 );
or \U$3389 ( \3514 , \3502 , \3513 );
and \U$3390 ( \3515 , \3499 , \3514 );
or \U$3391 ( \3516 , \3498 , \3515 );
and \U$3392 ( \3517 , \3495 , \3516 );
or \U$3393 ( \3518 , \3494 , \3517 );
and \U$3394 ( \3519 , \3491 , \3518 );
or \U$3395 ( \3520 , \3490 , \3519 );
and \U$3396 ( \3521 , \3487 , \3520 );
or \U$3397 ( \3522 , \3486 , \3521 );
and \U$3398 ( \3523 , \3483 , \3522 );
or \U$3399 ( \3524 , \3482 , \3523 );
and \U$3400 ( \3525 , \3479 , \3524 );
or \U$3401 ( \3526 , \3478 , \3525 );
and \U$3402 ( \3527 , \3475 , \3526 );
or \U$3403 ( \3528 , \3474 , \3527 );
and \U$3404 ( \3529 , \3471 , \3528 );
or \U$3405 ( \3530 , \3470 , \3529 );
and \U$3406 ( \3531 , \3467 , \3530 );
or \U$3407 ( \3532 , \3466 , \3531 );
and \U$3408 ( \3533 , \3463 , \3532 );
or \U$3409 ( \3534 , \3462 , \3533 );
and \U$3410 ( \3535 , \3459 , \3534 );
or \U$3411 ( \3536 , \3458 , \3535 );
and \U$3412 ( \3537 , \3455 , \3536 );
or \U$3413 ( \3538 , \3454 , \3537 );
and \U$3414 ( \3539 , \3451 , \3538 );
or \U$3415 ( \3540 , \3450 , \3539 );
and \U$3416 ( \3541 , \3447 , \3540 );
or \U$3417 ( \3542 , \3446 , \3541 );
_DC gdcb ( \3543_nGdcb , 1'b0 , \941 );
or \U$3419 ( \3544 , RI8928830_3, RI8929eb0_51);
and \U$3420 ( \3545 , \3544 , \940 );
and \U$3421 ( \3546 , RI8928fb0_19, RI8929730_35);
and \U$3422 ( \3547 , \3546 , \938 );
or \U$3423 ( \3548 , RI8928830_3, RI8928fb0_19);
and \U$3424 ( \3549 , \3548 , \936 );
xor \U$3425 ( \3550 , RI8929730_35, RI8929eb0_51);
and \U$3426 ( \3551 , \3550 , \934 );
buf \U$3427 ( \3552 , RI8928fb0_19);
and \U$3428 ( \3553 , \3552 , \952 );
and \U$3429 ( \3554 , \3277 , \955 );
xor \U$3430 ( \3555 , \3553 , \3554 );
and \U$3431 ( \3556 , \3278 , \3279 );
and \U$3432 ( \3557 , \3280 , \3283 );
or \U$3433 ( \3558 , \3556 , \3557 );
xor \U$3434 ( \3559 , \3555 , \3558 );
and \U$3435 ( \3560 , \3014 , \1193 );
xor \U$3436 ( \3561 , \3559 , \3560 );
and \U$3437 ( \3562 , \3284 , \3285 );
and \U$3438 ( \3563 , \3286 , \3289 );
or \U$3439 ( \3564 , \3562 , \3563 );
xor \U$3440 ( \3565 , \3561 , \3564 );
and \U$3441 ( \3566 , \2763 , \1354 );
xor \U$3442 ( \3567 , \3565 , \3566 );
and \U$3443 ( \3568 , \3290 , \3291 );
and \U$3444 ( \3569 , \3292 , \3295 );
or \U$3445 ( \3570 , \3568 , \3569 );
xor \U$3446 ( \3571 , \3567 , \3570 );
and \U$3447 ( \3572 , \2524 , \1527 );
xor \U$3448 ( \3573 , \3571 , \3572 );
and \U$3449 ( \3574 , \3296 , \3297 );
and \U$3450 ( \3575 , \3298 , \3301 );
or \U$3451 ( \3576 , \3574 , \3575 );
xor \U$3452 ( \3577 , \3573 , \3576 );
and \U$3453 ( \3578 , \2297 , \1712 );
xor \U$3454 ( \3579 , \3577 , \3578 );
and \U$3455 ( \3580 , \3302 , \3303 );
and \U$3456 ( \3581 , \3304 , \3307 );
or \U$3457 ( \3582 , \3580 , \3581 );
xor \U$3458 ( \3583 , \3579 , \3582 );
and \U$3459 ( \3584 , \2082 , \1909 );
xor \U$3460 ( \3585 , \3583 , \3584 );
and \U$3461 ( \3586 , \3308 , \3309 );
and \U$3462 ( \3587 , \3310 , \3313 );
or \U$3463 ( \3588 , \3586 , \3587 );
xor \U$3464 ( \3589 , \3585 , \3588 );
and \U$3465 ( \3590 , \1879 , \2118 );
xor \U$3466 ( \3591 , \3589 , \3590 );
and \U$3467 ( \3592 , \3314 , \3315 );
and \U$3468 ( \3593 , \3316 , \3319 );
or \U$3469 ( \3594 , \3592 , \3593 );
xor \U$3470 ( \3595 , \3591 , \3594 );
and \U$3471 ( \3596 , \1688 , \2339 );
xor \U$3472 ( \3597 , \3595 , \3596 );
and \U$3473 ( \3598 , \3320 , \3321 );
and \U$3474 ( \3599 , \3322 , \3325 );
or \U$3475 ( \3600 , \3598 , \3599 );
xor \U$3476 ( \3601 , \3597 , \3600 );
and \U$3477 ( \3602 , \1509 , \2572 );
xor \U$3478 ( \3603 , \3601 , \3602 );
and \U$3479 ( \3604 , \3326 , \3327 );
and \U$3480 ( \3605 , \3328 , \3331 );
or \U$3481 ( \3606 , \3604 , \3605 );
xor \U$3482 ( \3607 , \3603 , \3606 );
and \U$3483 ( \3608 , \1342 , \2817 );
xor \U$3484 ( \3609 , \3607 , \3608 );
and \U$3485 ( \3610 , \3332 , \3333 );
and \U$3486 ( \3611 , \3334 , \3337 );
or \U$3487 ( \3612 , \3610 , \3611 );
xor \U$3488 ( \3613 , \3609 , \3612 );
and \U$3489 ( \3614 , \1187 , \3074 );
xor \U$3490 ( \3615 , \3613 , \3614 );
and \U$3491 ( \3616 , \3338 , \3339 );
and \U$3492 ( \3617 , \3340 , \3341 );
or \U$3493 ( \3618 , \3616 , \3617 );
xor \U$3494 ( \3619 , \3615 , \3618 );
and \U$3495 ( \3620 , \951 , \3343 );
xor \U$3496 ( \3621 , \3619 , \3620 );
and \U$3497 ( \3622 , \3342 , \3344 );
xor \U$3498 ( \3623 , \3621 , \3622 );
buf \U$3499 ( \3624 , RI8929730_35);
and \U$3500 ( \3625 , \954 , \3624 );
xor \U$3501 ( \3626 , \3623 , \3625 );
buf \U$3502 ( \3627 , \3626 );
and \U$3503 ( \3628 , \3627 , \932 );
buf \U$3504 ( \3629 , RI8928830_3);
and \U$3505 ( \3630 , \3629 , \961 );
and \U$3506 ( \3631 , \3348 , \964 );
xor \U$3507 ( \3632 , \3630 , \3631 );
and \U$3508 ( \3633 , \3349 , \3350 );
and \U$3509 ( \3634 , \3351 , \3354 );
or \U$3510 ( \3635 , \3633 , \3634 );
xor \U$3511 ( \3636 , \3632 , \3635 );
and \U$3512 ( \3637 , \3079 , \1204 );
xor \U$3513 ( \3638 , \3636 , \3637 );
and \U$3514 ( \3639 , \3355 , \3356 );
and \U$3515 ( \3640 , \3357 , \3360 );
or \U$3516 ( \3641 , \3639 , \3640 );
xor \U$3517 ( \3642 , \3638 , \3641 );
and \U$3518 ( \3643 , \2822 , \1371 );
xor \U$3519 ( \3644 , \3642 , \3643 );
and \U$3520 ( \3645 , \3361 , \3362 );
and \U$3521 ( \3646 , \3363 , \3366 );
or \U$3522 ( \3647 , \3645 , \3646 );
xor \U$3523 ( \3648 , \3644 , \3647 );
and \U$3524 ( \3649 , \2577 , \1550 );
xor \U$3525 ( \3650 , \3648 , \3649 );
and \U$3526 ( \3651 , \3367 , \3368 );
and \U$3527 ( \3652 , \3369 , \3372 );
or \U$3528 ( \3653 , \3651 , \3652 );
xor \U$3529 ( \3654 , \3650 , \3653 );
and \U$3530 ( \3655 , \2344 , \1741 );
xor \U$3531 ( \3656 , \3654 , \3655 );
and \U$3532 ( \3657 , \3373 , \3374 );
and \U$3533 ( \3658 , \3375 , \3378 );
or \U$3534 ( \3659 , \3657 , \3658 );
xor \U$3535 ( \3660 , \3656 , \3659 );
and \U$3536 ( \3661 , \2123 , \1944 );
xor \U$3537 ( \3662 , \3660 , \3661 );
and \U$3538 ( \3663 , \3379 , \3380 );
and \U$3539 ( \3664 , \3381 , \3384 );
or \U$3540 ( \3665 , \3663 , \3664 );
xor \U$3541 ( \3666 , \3662 , \3665 );
and \U$3542 ( \3667 , \1914 , \2159 );
xor \U$3543 ( \3668 , \3666 , \3667 );
and \U$3544 ( \3669 , \3385 , \3386 );
and \U$3545 ( \3670 , \3387 , \3390 );
or \U$3546 ( \3671 , \3669 , \3670 );
xor \U$3547 ( \3672 , \3668 , \3671 );
and \U$3548 ( \3673 , \1717 , \2386 );
xor \U$3549 ( \3674 , \3672 , \3673 );
and \U$3550 ( \3675 , \3391 , \3392 );
and \U$3551 ( \3676 , \3393 , \3396 );
or \U$3552 ( \3677 , \3675 , \3676 );
xor \U$3553 ( \3678 , \3674 , \3677 );
and \U$3554 ( \3679 , \1532 , \2625 );
xor \U$3555 ( \3680 , \3678 , \3679 );
and \U$3556 ( \3681 , \3397 , \3398 );
and \U$3557 ( \3682 , \3399 , \3402 );
or \U$3558 ( \3683 , \3681 , \3682 );
xor \U$3559 ( \3684 , \3680 , \3683 );
and \U$3560 ( \3685 , \1359 , \2876 );
xor \U$3561 ( \3686 , \3684 , \3685 );
and \U$3562 ( \3687 , \3403 , \3404 );
and \U$3563 ( \3688 , \3405 , \3408 );
or \U$3564 ( \3689 , \3687 , \3688 );
xor \U$3565 ( \3690 , \3686 , \3689 );
and \U$3566 ( \3691 , \1198 , \3139 );
xor \U$3567 ( \3692 , \3690 , \3691 );
and \U$3568 ( \3693 , \3409 , \3410 );
and \U$3569 ( \3694 , \3411 , \3412 );
or \U$3570 ( \3695 , \3693 , \3694 );
xor \U$3571 ( \3696 , \3692 , \3695 );
and \U$3572 ( \3697 , \960 , \3414 );
xor \U$3573 ( \3698 , \3696 , \3697 );
and \U$3574 ( \3699 , \3413 , \3415 );
xor \U$3575 ( \3700 , \3698 , \3699 );
buf \U$3576 ( \3701 , RI8929eb0_51);
and \U$3577 ( \3702 , \963 , \3701 );
xor \U$3578 ( \3703 , \3700 , \3702 );
buf \U$3579 ( \3704 , \3703 );
and \U$3580 ( \3705 , \3704 , \930 );
buf \U$3581 ( \3706 , RI8928fb0_19);
buf \U$3582 ( \3707 , RI8929eb0_51);
xor \U$3583 ( \3708 , \3706 , \3707 );
and \U$3584 ( \3709 , \3419 , \3420 );
and \U$3585 ( \3710 , \3420 , \3425 );
and \U$3586 ( \3711 , \3419 , \3425 );
or \U$3587 ( \3712 , \3709 , \3710 , \3711 );
xor \U$3588 ( \3713 , \3708 , \3712 );
buf \U$3589 ( \3714 , \3713 );
and \U$3590 ( \3715 , \3714 , \928 );
buf \U$3591 ( \3716 , RI8928830_3);
buf \U$3592 ( \3717 , RI8929730_35);
xor \U$3593 ( \3718 , \3716 , \3717 );
and \U$3594 ( \3719 , \3429 , \3430 );
and \U$3595 ( \3720 , \3430 , \3435 );
and \U$3596 ( \3721 , \3429 , \3435 );
or \U$3597 ( \3722 , \3719 , \3720 , \3721 );
xor \U$3598 ( \3723 , \3718 , \3722 );
buf \U$3599 ( \3724 , \3723 );
and \U$3600 ( \3725 , \3724 , \926 );
and \U$3601 ( \3726 , RI8929eb0_51, \924 );
and \U$3602 ( \3727 , RI8929730_35, \922 );
and \U$3603 ( \3728 , RI8928fb0_19, \920 );
and \U$3604 ( \3729 , RI8928830_3, \918 );
or \U$3605 ( \3730 , \3543_nGdcb , \3545 , \3547 , \3549 , \3551 , \3628 , \3705 , \3715 , \3725 , \3726 , \3727 , \3728 , \3729 );
buf \U$3606 ( \3731 , \3730 );
and \U$3607 ( \3732 , \220 , \3731 );
and \U$3608 ( \3733 , \3542 , \3732 );
xor \U$3609 ( \3734 , \3542 , \3732 );
xor \U$3610 ( \3735 , \3447 , \3540 );
and \U$3611 ( \3736 , \1025 , \3731 );
and \U$3612 ( \3737 , \3735 , \3736 );
xor \U$3613 ( \3738 , \3735 , \3736 );
xor \U$3614 ( \3739 , \3451 , \3538 );
and \U$3615 ( \3740 , \1033 , \3731 );
and \U$3616 ( \3741 , \3739 , \3740 );
xor \U$3617 ( \3742 , \3739 , \3740 );
xor \U$3618 ( \3743 , \3455 , \3536 );
and \U$3619 ( \3744 , \1041 , \3731 );
and \U$3620 ( \3745 , \3743 , \3744 );
xor \U$3621 ( \3746 , \3743 , \3744 );
xor \U$3622 ( \3747 , \3459 , \3534 );
and \U$3623 ( \3748 , \1049 , \3731 );
and \U$3624 ( \3749 , \3747 , \3748 );
xor \U$3625 ( \3750 , \3747 , \3748 );
xor \U$3626 ( \3751 , \3463 , \3532 );
and \U$3627 ( \3752 , \1057 , \3731 );
and \U$3628 ( \3753 , \3751 , \3752 );
xor \U$3629 ( \3754 , \3751 , \3752 );
xor \U$3630 ( \3755 , \3467 , \3530 );
and \U$3631 ( \3756 , \1065 , \3731 );
and \U$3632 ( \3757 , \3755 , \3756 );
xor \U$3633 ( \3758 , \3755 , \3756 );
xor \U$3634 ( \3759 , \3471 , \3528 );
and \U$3635 ( \3760 , \1073 , \3731 );
and \U$3636 ( \3761 , \3759 , \3760 );
xor \U$3637 ( \3762 , \3759 , \3760 );
xor \U$3638 ( \3763 , \3475 , \3526 );
and \U$3639 ( \3764 , \1081 , \3731 );
and \U$3640 ( \3765 , \3763 , \3764 );
xor \U$3641 ( \3766 , \3763 , \3764 );
xor \U$3642 ( \3767 , \3479 , \3524 );
and \U$3643 ( \3768 , \1089 , \3731 );
and \U$3644 ( \3769 , \3767 , \3768 );
xor \U$3645 ( \3770 , \3767 , \3768 );
xor \U$3646 ( \3771 , \3483 , \3522 );
and \U$3647 ( \3772 , \1097 , \3731 );
and \U$3648 ( \3773 , \3771 , \3772 );
xor \U$3649 ( \3774 , \3771 , \3772 );
xor \U$3650 ( \3775 , \3487 , \3520 );
and \U$3651 ( \3776 , \1105 , \3731 );
and \U$3652 ( \3777 , \3775 , \3776 );
xor \U$3653 ( \3778 , \3775 , \3776 );
xor \U$3654 ( \3779 , \3491 , \3518 );
and \U$3655 ( \3780 , \1113 , \3731 );
and \U$3656 ( \3781 , \3779 , \3780 );
xor \U$3657 ( \3782 , \3779 , \3780 );
xor \U$3658 ( \3783 , \3495 , \3516 );
and \U$3659 ( \3784 , \1121 , \3731 );
and \U$3660 ( \3785 , \3783 , \3784 );
xor \U$3661 ( \3786 , \3783 , \3784 );
xor \U$3662 ( \3787 , \3499 , \3514 );
and \U$3663 ( \3788 , \1129 , \3731 );
and \U$3664 ( \3789 , \3787 , \3788 );
xor \U$3665 ( \3790 , \3787 , \3788 );
xor \U$3666 ( \3791 , \3503 , \3512 );
and \U$3667 ( \3792 , \1137 , \3731 );
and \U$3668 ( \3793 , \3791 , \3792 );
xor \U$3669 ( \3794 , \3791 , \3792 );
xor \U$3670 ( \3795 , \3507 , \3510 );
and \U$3671 ( \3796 , \1144 , \3731 );
and \U$3672 ( \3797 , \3795 , \3796 );
and \U$3673 ( \3798 , \3794 , \3797 );
or \U$3674 ( \3799 , \3793 , \3798 );
and \U$3675 ( \3800 , \3790 , \3799 );
or \U$3676 ( \3801 , \3789 , \3800 );
and \U$3677 ( \3802 , \3786 , \3801 );
or \U$3678 ( \3803 , \3785 , \3802 );
and \U$3679 ( \3804 , \3782 , \3803 );
or \U$3680 ( \3805 , \3781 , \3804 );
and \U$3681 ( \3806 , \3778 , \3805 );
or \U$3682 ( \3807 , \3777 , \3806 );
and \U$3683 ( \3808 , \3774 , \3807 );
or \U$3684 ( \3809 , \3773 , \3808 );
and \U$3685 ( \3810 , \3770 , \3809 );
or \U$3686 ( \3811 , \3769 , \3810 );
and \U$3687 ( \3812 , \3766 , \3811 );
or \U$3688 ( \3813 , \3765 , \3812 );
and \U$3689 ( \3814 , \3762 , \3813 );
or \U$3690 ( \3815 , \3761 , \3814 );
and \U$3691 ( \3816 , \3758 , \3815 );
or \U$3692 ( \3817 , \3757 , \3816 );
and \U$3693 ( \3818 , \3754 , \3817 );
or \U$3694 ( \3819 , \3753 , \3818 );
and \U$3695 ( \3820 , \3750 , \3819 );
or \U$3696 ( \3821 , \3749 , \3820 );
and \U$3697 ( \3822 , \3746 , \3821 );
or \U$3698 ( \3823 , \3745 , \3822 );
and \U$3699 ( \3824 , \3742 , \3823 );
or \U$3700 ( \3825 , \3741 , \3824 );
and \U$3701 ( \3826 , \3738 , \3825 );
or \U$3702 ( \3827 , \3737 , \3826 );
and \U$3703 ( \3828 , \3734 , \3827 );
or \U$3704 ( \3829 , \3733 , \3828 );
_DC geea ( \3830_nGeea , 1'b0 , \941 );
or \U$3706 ( \3831 , RI89287b8_2, RI8929e38_50);
and \U$3707 ( \3832 , \3831 , \940 );
and \U$3708 ( \3833 , RI8928f38_18, RI89296b8_34);
and \U$3709 ( \3834 , \3833 , \938 );
or \U$3710 ( \3835 , RI89287b8_2, RI8928f38_18);
and \U$3711 ( \3836 , \3835 , \936 );
xor \U$3712 ( \3837 , RI89296b8_34, RI8929e38_50);
and \U$3713 ( \3838 , \3837 , \934 );
buf \U$3714 ( \3839 , RI8928f38_18);
and \U$3715 ( \3840 , \3839 , \952 );
and \U$3716 ( \3841 , \3552 , \955 );
xor \U$3717 ( \3842 , \3840 , \3841 );
and \U$3718 ( \3843 , \3553 , \3554 );
and \U$3719 ( \3844 , \3555 , \3558 );
or \U$3720 ( \3845 , \3843 , \3844 );
xor \U$3721 ( \3846 , \3842 , \3845 );
and \U$3722 ( \3847 , \3277 , \1193 );
xor \U$3723 ( \3848 , \3846 , \3847 );
and \U$3724 ( \3849 , \3559 , \3560 );
and \U$3725 ( \3850 , \3561 , \3564 );
or \U$3726 ( \3851 , \3849 , \3850 );
xor \U$3727 ( \3852 , \3848 , \3851 );
and \U$3728 ( \3853 , \3014 , \1354 );
xor \U$3729 ( \3854 , \3852 , \3853 );
and \U$3730 ( \3855 , \3565 , \3566 );
and \U$3731 ( \3856 , \3567 , \3570 );
or \U$3732 ( \3857 , \3855 , \3856 );
xor \U$3733 ( \3858 , \3854 , \3857 );
and \U$3734 ( \3859 , \2763 , \1527 );
xor \U$3735 ( \3860 , \3858 , \3859 );
and \U$3736 ( \3861 , \3571 , \3572 );
and \U$3737 ( \3862 , \3573 , \3576 );
or \U$3738 ( \3863 , \3861 , \3862 );
xor \U$3739 ( \3864 , \3860 , \3863 );
and \U$3740 ( \3865 , \2524 , \1712 );
xor \U$3741 ( \3866 , \3864 , \3865 );
and \U$3742 ( \3867 , \3577 , \3578 );
and \U$3743 ( \3868 , \3579 , \3582 );
or \U$3744 ( \3869 , \3867 , \3868 );
xor \U$3745 ( \3870 , \3866 , \3869 );
and \U$3746 ( \3871 , \2297 , \1909 );
xor \U$3747 ( \3872 , \3870 , \3871 );
and \U$3748 ( \3873 , \3583 , \3584 );
and \U$3749 ( \3874 , \3585 , \3588 );
or \U$3750 ( \3875 , \3873 , \3874 );
xor \U$3751 ( \3876 , \3872 , \3875 );
and \U$3752 ( \3877 , \2082 , \2118 );
xor \U$3753 ( \3878 , \3876 , \3877 );
and \U$3754 ( \3879 , \3589 , \3590 );
and \U$3755 ( \3880 , \3591 , \3594 );
or \U$3756 ( \3881 , \3879 , \3880 );
xor \U$3757 ( \3882 , \3878 , \3881 );
and \U$3758 ( \3883 , \1879 , \2339 );
xor \U$3759 ( \3884 , \3882 , \3883 );
and \U$3760 ( \3885 , \3595 , \3596 );
and \U$3761 ( \3886 , \3597 , \3600 );
or \U$3762 ( \3887 , \3885 , \3886 );
xor \U$3763 ( \3888 , \3884 , \3887 );
and \U$3764 ( \3889 , \1688 , \2572 );
xor \U$3765 ( \3890 , \3888 , \3889 );
and \U$3766 ( \3891 , \3601 , \3602 );
and \U$3767 ( \3892 , \3603 , \3606 );
or \U$3768 ( \3893 , \3891 , \3892 );
xor \U$3769 ( \3894 , \3890 , \3893 );
and \U$3770 ( \3895 , \1509 , \2817 );
xor \U$3771 ( \3896 , \3894 , \3895 );
and \U$3772 ( \3897 , \3607 , \3608 );
and \U$3773 ( \3898 , \3609 , \3612 );
or \U$3774 ( \3899 , \3897 , \3898 );
xor \U$3775 ( \3900 , \3896 , \3899 );
and \U$3776 ( \3901 , \1342 , \3074 );
xor \U$3777 ( \3902 , \3900 , \3901 );
and \U$3778 ( \3903 , \3613 , \3614 );
and \U$3779 ( \3904 , \3615 , \3618 );
or \U$3780 ( \3905 , \3903 , \3904 );
xor \U$3781 ( \3906 , \3902 , \3905 );
and \U$3782 ( \3907 , \1187 , \3343 );
xor \U$3783 ( \3908 , \3906 , \3907 );
and \U$3784 ( \3909 , \3619 , \3620 );
and \U$3785 ( \3910 , \3621 , \3622 );
or \U$3786 ( \3911 , \3909 , \3910 );
xor \U$3787 ( \3912 , \3908 , \3911 );
and \U$3788 ( \3913 , \951 , \3624 );
xor \U$3789 ( \3914 , \3912 , \3913 );
and \U$3790 ( \3915 , \3623 , \3625 );
xor \U$3791 ( \3916 , \3914 , \3915 );
buf \U$3792 ( \3917 , RI89296b8_34);
and \U$3793 ( \3918 , \954 , \3917 );
xor \U$3794 ( \3919 , \3916 , \3918 );
buf \U$3795 ( \3920 , \3919 );
and \U$3796 ( \3921 , \3920 , \932 );
buf \U$3797 ( \3922 , RI89287b8_2);
and \U$3798 ( \3923 , \3922 , \961 );
and \U$3799 ( \3924 , \3629 , \964 );
xor \U$3800 ( \3925 , \3923 , \3924 );
and \U$3801 ( \3926 , \3630 , \3631 );
and \U$3802 ( \3927 , \3632 , \3635 );
or \U$3803 ( \3928 , \3926 , \3927 );
xor \U$3804 ( \3929 , \3925 , \3928 );
and \U$3805 ( \3930 , \3348 , \1204 );
xor \U$3806 ( \3931 , \3929 , \3930 );
and \U$3807 ( \3932 , \3636 , \3637 );
and \U$3808 ( \3933 , \3638 , \3641 );
or \U$3809 ( \3934 , \3932 , \3933 );
xor \U$3810 ( \3935 , \3931 , \3934 );
and \U$3811 ( \3936 , \3079 , \1371 );
xor \U$3812 ( \3937 , \3935 , \3936 );
and \U$3813 ( \3938 , \3642 , \3643 );
and \U$3814 ( \3939 , \3644 , \3647 );
or \U$3815 ( \3940 , \3938 , \3939 );
xor \U$3816 ( \3941 , \3937 , \3940 );
and \U$3817 ( \3942 , \2822 , \1550 );
xor \U$3818 ( \3943 , \3941 , \3942 );
and \U$3819 ( \3944 , \3648 , \3649 );
and \U$3820 ( \3945 , \3650 , \3653 );
or \U$3821 ( \3946 , \3944 , \3945 );
xor \U$3822 ( \3947 , \3943 , \3946 );
and \U$3823 ( \3948 , \2577 , \1741 );
xor \U$3824 ( \3949 , \3947 , \3948 );
and \U$3825 ( \3950 , \3654 , \3655 );
and \U$3826 ( \3951 , \3656 , \3659 );
or \U$3827 ( \3952 , \3950 , \3951 );
xor \U$3828 ( \3953 , \3949 , \3952 );
and \U$3829 ( \3954 , \2344 , \1944 );
xor \U$3830 ( \3955 , \3953 , \3954 );
and \U$3831 ( \3956 , \3660 , \3661 );
and \U$3832 ( \3957 , \3662 , \3665 );
or \U$3833 ( \3958 , \3956 , \3957 );
xor \U$3834 ( \3959 , \3955 , \3958 );
and \U$3835 ( \3960 , \2123 , \2159 );
xor \U$3836 ( \3961 , \3959 , \3960 );
and \U$3837 ( \3962 , \3666 , \3667 );
and \U$3838 ( \3963 , \3668 , \3671 );
or \U$3839 ( \3964 , \3962 , \3963 );
xor \U$3840 ( \3965 , \3961 , \3964 );
and \U$3841 ( \3966 , \1914 , \2386 );
xor \U$3842 ( \3967 , \3965 , \3966 );
and \U$3843 ( \3968 , \3672 , \3673 );
and \U$3844 ( \3969 , \3674 , \3677 );
or \U$3845 ( \3970 , \3968 , \3969 );
xor \U$3846 ( \3971 , \3967 , \3970 );
and \U$3847 ( \3972 , \1717 , \2625 );
xor \U$3848 ( \3973 , \3971 , \3972 );
and \U$3849 ( \3974 , \3678 , \3679 );
and \U$3850 ( \3975 , \3680 , \3683 );
or \U$3851 ( \3976 , \3974 , \3975 );
xor \U$3852 ( \3977 , \3973 , \3976 );
and \U$3853 ( \3978 , \1532 , \2876 );
xor \U$3854 ( \3979 , \3977 , \3978 );
and \U$3855 ( \3980 , \3684 , \3685 );
and \U$3856 ( \3981 , \3686 , \3689 );
or \U$3857 ( \3982 , \3980 , \3981 );
xor \U$3858 ( \3983 , \3979 , \3982 );
and \U$3859 ( \3984 , \1359 , \3139 );
xor \U$3860 ( \3985 , \3983 , \3984 );
and \U$3861 ( \3986 , \3690 , \3691 );
and \U$3862 ( \3987 , \3692 , \3695 );
or \U$3863 ( \3988 , \3986 , \3987 );
xor \U$3864 ( \3989 , \3985 , \3988 );
and \U$3865 ( \3990 , \1198 , \3414 );
xor \U$3866 ( \3991 , \3989 , \3990 );
and \U$3867 ( \3992 , \3696 , \3697 );
and \U$3868 ( \3993 , \3698 , \3699 );
or \U$3869 ( \3994 , \3992 , \3993 );
xor \U$3870 ( \3995 , \3991 , \3994 );
and \U$3871 ( \3996 , \960 , \3701 );
xor \U$3872 ( \3997 , \3995 , \3996 );
and \U$3873 ( \3998 , \3700 , \3702 );
xor \U$3874 ( \3999 , \3997 , \3998 );
buf \U$3875 ( \4000 , RI8929e38_50);
and \U$3876 ( \4001 , \963 , \4000 );
xor \U$3877 ( \4002 , \3999 , \4001 );
buf \U$3878 ( \4003 , \4002 );
and \U$3879 ( \4004 , \4003 , \930 );
buf \U$3880 ( \4005 , RI8928f38_18);
buf \U$3881 ( \4006 , RI8929e38_50);
xor \U$3882 ( \4007 , \4005 , \4006 );
and \U$3883 ( \4008 , \3706 , \3707 );
and \U$3884 ( \4009 , \3707 , \3712 );
and \U$3885 ( \4010 , \3706 , \3712 );
or \U$3886 ( \4011 , \4008 , \4009 , \4010 );
xor \U$3887 ( \4012 , \4007 , \4011 );
buf \U$3888 ( \4013 , \4012 );
and \U$3889 ( \4014 , \4013 , \928 );
buf \U$3890 ( \4015 , RI89287b8_2);
buf \U$3891 ( \4016 , RI89296b8_34);
xor \U$3892 ( \4017 , \4015 , \4016 );
and \U$3893 ( \4018 , \3716 , \3717 );
and \U$3894 ( \4019 , \3717 , \3722 );
and \U$3895 ( \4020 , \3716 , \3722 );
or \U$3896 ( \4021 , \4018 , \4019 , \4020 );
xor \U$3897 ( \4022 , \4017 , \4021 );
buf \U$3898 ( \4023 , \4022 );
and \U$3899 ( \4024 , \4023 , \926 );
and \U$3900 ( \4025 , RI8929e38_50, \924 );
and \U$3901 ( \4026 , RI89296b8_34, \922 );
and \U$3902 ( \4027 , RI8928f38_18, \920 );
and \U$3903 ( \4028 , RI89287b8_2, \918 );
or \U$3904 ( \4029 , \3830_nGeea , \3832 , \3834 , \3836 , \3838 , \3921 , \4004 , \4014 , \4024 , \4025 , \4026 , \4027 , \4028 );
buf \U$3905 ( \4030 , \4029 );
and \U$3906 ( \4031 , \220 , \4030 );
and \U$3907 ( \4032 , \3829 , \4031 );
xor \U$3908 ( \4033 , \3829 , \4031 );
xor \U$3909 ( \4034 , \3734 , \3827 );
and \U$3910 ( \4035 , \1025 , \4030 );
and \U$3911 ( \4036 , \4034 , \4035 );
xor \U$3912 ( \4037 , \4034 , \4035 );
xor \U$3913 ( \4038 , \3738 , \3825 );
and \U$3914 ( \4039 , \1033 , \4030 );
and \U$3915 ( \4040 , \4038 , \4039 );
xor \U$3916 ( \4041 , \4038 , \4039 );
xor \U$3917 ( \4042 , \3742 , \3823 );
and \U$3918 ( \4043 , \1041 , \4030 );
and \U$3919 ( \4044 , \4042 , \4043 );
xor \U$3920 ( \4045 , \4042 , \4043 );
xor \U$3921 ( \4046 , \3746 , \3821 );
and \U$3922 ( \4047 , \1049 , \4030 );
and \U$3923 ( \4048 , \4046 , \4047 );
xor \U$3924 ( \4049 , \4046 , \4047 );
xor \U$3925 ( \4050 , \3750 , \3819 );
and \U$3926 ( \4051 , \1057 , \4030 );
and \U$3927 ( \4052 , \4050 , \4051 );
xor \U$3928 ( \4053 , \4050 , \4051 );
xor \U$3929 ( \4054 , \3754 , \3817 );
and \U$3930 ( \4055 , \1065 , \4030 );
and \U$3931 ( \4056 , \4054 , \4055 );
xor \U$3932 ( \4057 , \4054 , \4055 );
xor \U$3933 ( \4058 , \3758 , \3815 );
and \U$3934 ( \4059 , \1073 , \4030 );
and \U$3935 ( \4060 , \4058 , \4059 );
xor \U$3936 ( \4061 , \4058 , \4059 );
xor \U$3937 ( \4062 , \3762 , \3813 );
and \U$3938 ( \4063 , \1081 , \4030 );
and \U$3939 ( \4064 , \4062 , \4063 );
xor \U$3940 ( \4065 , \4062 , \4063 );
xor \U$3941 ( \4066 , \3766 , \3811 );
and \U$3942 ( \4067 , \1089 , \4030 );
and \U$3943 ( \4068 , \4066 , \4067 );
xor \U$3944 ( \4069 , \4066 , \4067 );
xor \U$3945 ( \4070 , \3770 , \3809 );
and \U$3946 ( \4071 , \1097 , \4030 );
and \U$3947 ( \4072 , \4070 , \4071 );
xor \U$3948 ( \4073 , \4070 , \4071 );
xor \U$3949 ( \4074 , \3774 , \3807 );
and \U$3950 ( \4075 , \1105 , \4030 );
and \U$3951 ( \4076 , \4074 , \4075 );
xor \U$3952 ( \4077 , \4074 , \4075 );
xor \U$3953 ( \4078 , \3778 , \3805 );
and \U$3954 ( \4079 , \1113 , \4030 );
and \U$3955 ( \4080 , \4078 , \4079 );
xor \U$3956 ( \4081 , \4078 , \4079 );
xor \U$3957 ( \4082 , \3782 , \3803 );
and \U$3958 ( \4083 , \1121 , \4030 );
and \U$3959 ( \4084 , \4082 , \4083 );
xor \U$3960 ( \4085 , \4082 , \4083 );
xor \U$3961 ( \4086 , \3786 , \3801 );
and \U$3962 ( \4087 , \1129 , \4030 );
and \U$3963 ( \4088 , \4086 , \4087 );
xor \U$3964 ( \4089 , \4086 , \4087 );
xor \U$3965 ( \4090 , \3790 , \3799 );
and \U$3966 ( \4091 , \1137 , \4030 );
and \U$3967 ( \4092 , \4090 , \4091 );
xor \U$3968 ( \4093 , \4090 , \4091 );
xor \U$3969 ( \4094 , \3794 , \3797 );
and \U$3970 ( \4095 , \1144 , \4030 );
and \U$3971 ( \4096 , \4094 , \4095 );
and \U$3972 ( \4097 , \4093 , \4096 );
or \U$3973 ( \4098 , \4092 , \4097 );
and \U$3974 ( \4099 , \4089 , \4098 );
or \U$3975 ( \4100 , \4088 , \4099 );
and \U$3976 ( \4101 , \4085 , \4100 );
or \U$3977 ( \4102 , \4084 , \4101 );
and \U$3978 ( \4103 , \4081 , \4102 );
or \U$3979 ( \4104 , \4080 , \4103 );
and \U$3980 ( \4105 , \4077 , \4104 );
or \U$3981 ( \4106 , \4076 , \4105 );
and \U$3982 ( \4107 , \4073 , \4106 );
or \U$3983 ( \4108 , \4072 , \4107 );
and \U$3984 ( \4109 , \4069 , \4108 );
or \U$3985 ( \4110 , \4068 , \4109 );
and \U$3986 ( \4111 , \4065 , \4110 );
or \U$3987 ( \4112 , \4064 , \4111 );
and \U$3988 ( \4113 , \4061 , \4112 );
or \U$3989 ( \4114 , \4060 , \4113 );
and \U$3990 ( \4115 , \4057 , \4114 );
or \U$3991 ( \4116 , \4056 , \4115 );
and \U$3992 ( \4117 , \4053 , \4116 );
or \U$3993 ( \4118 , \4052 , \4117 );
and \U$3994 ( \4119 , \4049 , \4118 );
or \U$3995 ( \4120 , \4048 , \4119 );
and \U$3996 ( \4121 , \4045 , \4120 );
or \U$3997 ( \4122 , \4044 , \4121 );
and \U$3998 ( \4123 , \4041 , \4122 );
or \U$3999 ( \4124 , \4040 , \4123 );
and \U$4000 ( \4125 , \4037 , \4124 );
or \U$4001 ( \4126 , \4036 , \4125 );
and \U$4002 ( \4127 , \4033 , \4126 );
or \U$4003 ( \4128 , \4032 , \4127 );
_DC g1015 ( \4129_nG1015 , 1'b0 , \941 );
or \U$4005 ( \4130 , RI8928740_1, RI8929dc0_49);
and \U$4006 ( \4131 , \4130 , \940 );
and \U$4007 ( \4132 , RI8928ec0_17, RI8929640_33);
and \U$4008 ( \4133 , \4132 , \938 );
or \U$4009 ( \4134 , RI8928740_1, RI8928ec0_17);
and \U$4010 ( \4135 , \4134 , \936 );
xor \U$4011 ( \4136 , RI8929640_33, RI8929dc0_49);
and \U$4012 ( \4137 , \4136 , \934 );
buf \U$4013 ( \4138 , RI8928ec0_17);
and \U$4014 ( \4139 , \4138 , \952 );
and \U$4015 ( \4140 , \3839 , \955 );
xor \U$4016 ( \4141 , \4139 , \4140 );
and \U$4017 ( \4142 , \3840 , \3841 );
and \U$4018 ( \4143 , \3842 , \3845 );
or \U$4019 ( \4144 , \4142 , \4143 );
xor \U$4020 ( \4145 , \4141 , \4144 );
and \U$4021 ( \4146 , \3552 , \1193 );
xor \U$4022 ( \4147 , \4145 , \4146 );
and \U$4023 ( \4148 , \3846 , \3847 );
and \U$4024 ( \4149 , \3848 , \3851 );
or \U$4025 ( \4150 , \4148 , \4149 );
xor \U$4026 ( \4151 , \4147 , \4150 );
and \U$4027 ( \4152 , \3277 , \1354 );
xor \U$4028 ( \4153 , \4151 , \4152 );
and \U$4029 ( \4154 , \3852 , \3853 );
and \U$4030 ( \4155 , \3854 , \3857 );
or \U$4031 ( \4156 , \4154 , \4155 );
xor \U$4032 ( \4157 , \4153 , \4156 );
and \U$4033 ( \4158 , \3014 , \1527 );
xor \U$4034 ( \4159 , \4157 , \4158 );
and \U$4035 ( \4160 , \3858 , \3859 );
and \U$4036 ( \4161 , \3860 , \3863 );
or \U$4037 ( \4162 , \4160 , \4161 );
xor \U$4038 ( \4163 , \4159 , \4162 );
and \U$4039 ( \4164 , \2763 , \1712 );
xor \U$4040 ( \4165 , \4163 , \4164 );
and \U$4041 ( \4166 , \3864 , \3865 );
and \U$4042 ( \4167 , \3866 , \3869 );
or \U$4043 ( \4168 , \4166 , \4167 );
xor \U$4044 ( \4169 , \4165 , \4168 );
and \U$4045 ( \4170 , \2524 , \1909 );
xor \U$4046 ( \4171 , \4169 , \4170 );
and \U$4047 ( \4172 , \3870 , \3871 );
and \U$4048 ( \4173 , \3872 , \3875 );
or \U$4049 ( \4174 , \4172 , \4173 );
xor \U$4050 ( \4175 , \4171 , \4174 );
and \U$4051 ( \4176 , \2297 , \2118 );
xor \U$4052 ( \4177 , \4175 , \4176 );
and \U$4053 ( \4178 , \3876 , \3877 );
and \U$4054 ( \4179 , \3878 , \3881 );
or \U$4055 ( \4180 , \4178 , \4179 );
xor \U$4056 ( \4181 , \4177 , \4180 );
and \U$4057 ( \4182 , \2082 , \2339 );
xor \U$4058 ( \4183 , \4181 , \4182 );
and \U$4059 ( \4184 , \3882 , \3883 );
and \U$4060 ( \4185 , \3884 , \3887 );
or \U$4061 ( \4186 , \4184 , \4185 );
xor \U$4062 ( \4187 , \4183 , \4186 );
and \U$4063 ( \4188 , \1879 , \2572 );
xor \U$4064 ( \4189 , \4187 , \4188 );
and \U$4065 ( \4190 , \3888 , \3889 );
and \U$4066 ( \4191 , \3890 , \3893 );
or \U$4067 ( \4192 , \4190 , \4191 );
xor \U$4068 ( \4193 , \4189 , \4192 );
and \U$4069 ( \4194 , \1688 , \2817 );
xor \U$4070 ( \4195 , \4193 , \4194 );
and \U$4071 ( \4196 , \3894 , \3895 );
and \U$4072 ( \4197 , \3896 , \3899 );
or \U$4073 ( \4198 , \4196 , \4197 );
xor \U$4074 ( \4199 , \4195 , \4198 );
and \U$4075 ( \4200 , \1509 , \3074 );
xor \U$4076 ( \4201 , \4199 , \4200 );
and \U$4077 ( \4202 , \3900 , \3901 );
and \U$4078 ( \4203 , \3902 , \3905 );
or \U$4079 ( \4204 , \4202 , \4203 );
xor \U$4080 ( \4205 , \4201 , \4204 );
and \U$4081 ( \4206 , \1342 , \3343 );
xor \U$4082 ( \4207 , \4205 , \4206 );
and \U$4083 ( \4208 , \3906 , \3907 );
and \U$4084 ( \4209 , \3908 , \3911 );
or \U$4085 ( \4210 , \4208 , \4209 );
xor \U$4086 ( \4211 , \4207 , \4210 );
and \U$4087 ( \4212 , \1187 , \3624 );
xor \U$4088 ( \4213 , \4211 , \4212 );
and \U$4089 ( \4214 , \3912 , \3913 );
and \U$4090 ( \4215 , \3914 , \3915 );
or \U$4091 ( \4216 , \4214 , \4215 );
xor \U$4092 ( \4217 , \4213 , \4216 );
and \U$4093 ( \4218 , \951 , \3917 );
xor \U$4094 ( \4219 , \4217 , \4218 );
and \U$4095 ( \4220 , \3916 , \3918 );
xor \U$4096 ( \4221 , \4219 , \4220 );
buf \U$4097 ( \4222 , RI8929640_33);
and \U$4098 ( \4223 , \954 , \4222 );
xor \U$4099 ( \4224 , \4221 , \4223 );
buf \U$4100 ( \4225 , \4224 );
and \U$4101 ( \4226 , \4225 , \932 );
buf \U$4102 ( \4227 , RI8928740_1);
and \U$4103 ( \4228 , \4227 , \961 );
and \U$4104 ( \4229 , \3922 , \964 );
xor \U$4105 ( \4230 , \4228 , \4229 );
and \U$4106 ( \4231 , \3923 , \3924 );
and \U$4107 ( \4232 , \3925 , \3928 );
or \U$4108 ( \4233 , \4231 , \4232 );
xor \U$4109 ( \4234 , \4230 , \4233 );
and \U$4110 ( \4235 , \3629 , \1204 );
xor \U$4111 ( \4236 , \4234 , \4235 );
and \U$4112 ( \4237 , \3929 , \3930 );
and \U$4113 ( \4238 , \3931 , \3934 );
or \U$4114 ( \4239 , \4237 , \4238 );
xor \U$4115 ( \4240 , \4236 , \4239 );
and \U$4116 ( \4241 , \3348 , \1371 );
xor \U$4117 ( \4242 , \4240 , \4241 );
and \U$4118 ( \4243 , \3935 , \3936 );
and \U$4119 ( \4244 , \3937 , \3940 );
or \U$4120 ( \4245 , \4243 , \4244 );
xor \U$4121 ( \4246 , \4242 , \4245 );
and \U$4122 ( \4247 , \3079 , \1550 );
xor \U$4123 ( \4248 , \4246 , \4247 );
and \U$4124 ( \4249 , \3941 , \3942 );
and \U$4125 ( \4250 , \3943 , \3946 );
or \U$4126 ( \4251 , \4249 , \4250 );
xor \U$4127 ( \4252 , \4248 , \4251 );
and \U$4128 ( \4253 , \2822 , \1741 );
xor \U$4129 ( \4254 , \4252 , \4253 );
and \U$4130 ( \4255 , \3947 , \3948 );
and \U$4131 ( \4256 , \3949 , \3952 );
or \U$4132 ( \4257 , \4255 , \4256 );
xor \U$4133 ( \4258 , \4254 , \4257 );
and \U$4134 ( \4259 , \2577 , \1944 );
xor \U$4135 ( \4260 , \4258 , \4259 );
and \U$4136 ( \4261 , \3953 , \3954 );
and \U$4137 ( \4262 , \3955 , \3958 );
or \U$4138 ( \4263 , \4261 , \4262 );
xor \U$4139 ( \4264 , \4260 , \4263 );
and \U$4140 ( \4265 , \2344 , \2159 );
xor \U$4141 ( \4266 , \4264 , \4265 );
and \U$4142 ( \4267 , \3959 , \3960 );
and \U$4143 ( \4268 , \3961 , \3964 );
or \U$4144 ( \4269 , \4267 , \4268 );
xor \U$4145 ( \4270 , \4266 , \4269 );
and \U$4146 ( \4271 , \2123 , \2386 );
xor \U$4147 ( \4272 , \4270 , \4271 );
and \U$4148 ( \4273 , \3965 , \3966 );
and \U$4149 ( \4274 , \3967 , \3970 );
or \U$4150 ( \4275 , \4273 , \4274 );
xor \U$4151 ( \4276 , \4272 , \4275 );
and \U$4152 ( \4277 , \1914 , \2625 );
xor \U$4153 ( \4278 , \4276 , \4277 );
and \U$4154 ( \4279 , \3971 , \3972 );
and \U$4155 ( \4280 , \3973 , \3976 );
or \U$4156 ( \4281 , \4279 , \4280 );
xor \U$4157 ( \4282 , \4278 , \4281 );
and \U$4158 ( \4283 , \1717 , \2876 );
xor \U$4159 ( \4284 , \4282 , \4283 );
and \U$4160 ( \4285 , \3977 , \3978 );
and \U$4161 ( \4286 , \3979 , \3982 );
or \U$4162 ( \4287 , \4285 , \4286 );
xor \U$4163 ( \4288 , \4284 , \4287 );
and \U$4164 ( \4289 , \1532 , \3139 );
xor \U$4165 ( \4290 , \4288 , \4289 );
and \U$4166 ( \4291 , \3983 , \3984 );
and \U$4167 ( \4292 , \3985 , \3988 );
or \U$4168 ( \4293 , \4291 , \4292 );
xor \U$4169 ( \4294 , \4290 , \4293 );
and \U$4170 ( \4295 , \1359 , \3414 );
xor \U$4171 ( \4296 , \4294 , \4295 );
and \U$4172 ( \4297 , \3989 , \3990 );
and \U$4173 ( \4298 , \3991 , \3994 );
or \U$4174 ( \4299 , \4297 , \4298 );
xor \U$4175 ( \4300 , \4296 , \4299 );
and \U$4176 ( \4301 , \1198 , \3701 );
xor \U$4177 ( \4302 , \4300 , \4301 );
and \U$4178 ( \4303 , \3995 , \3996 );
and \U$4179 ( \4304 , \3997 , \3998 );
or \U$4180 ( \4305 , \4303 , \4304 );
xor \U$4181 ( \4306 , \4302 , \4305 );
and \U$4182 ( \4307 , \960 , \4000 );
xor \U$4183 ( \4308 , \4306 , \4307 );
and \U$4184 ( \4309 , \3999 , \4001 );
xor \U$4185 ( \4310 , \4308 , \4309 );
buf \U$4186 ( \4311 , RI8929dc0_49);
and \U$4187 ( \4312 , \963 , \4311 );
xor \U$4188 ( \4313 , \4310 , \4312 );
buf \U$4189 ( \4314 , \4313 );
and \U$4190 ( \4315 , \4314 , \930 );
buf \U$4191 ( \4316 , RI8928ec0_17);
buf \U$4192 ( \4317 , RI8929dc0_49);
xor \U$4193 ( \4318 , \4316 , \4317 );
and \U$4194 ( \4319 , \4005 , \4006 );
and \U$4195 ( \4320 , \4006 , \4011 );
and \U$4196 ( \4321 , \4005 , \4011 );
or \U$4197 ( \4322 , \4319 , \4320 , \4321 );
xor \U$4198 ( \4323 , \4318 , \4322 );
buf \U$4199 ( \4324 , \4323 );
and \U$4200 ( \4325 , \4324 , \928 );
buf \U$4201 ( \4326 , RI8928740_1);
buf \U$4202 ( \4327 , RI8929640_33);
xor \U$4203 ( \4328 , \4326 , \4327 );
and \U$4204 ( \4329 , \4015 , \4016 );
and \U$4205 ( \4330 , \4016 , \4021 );
and \U$4206 ( \4331 , \4015 , \4021 );
or \U$4207 ( \4332 , \4329 , \4330 , \4331 );
xor \U$4208 ( \4333 , \4328 , \4332 );
buf \U$4209 ( \4334 , \4333 );
and \U$4210 ( \4335 , \4334 , \926 );
and \U$4211 ( \4336 , RI8929dc0_49, \924 );
and \U$4212 ( \4337 , RI8929640_33, \922 );
and \U$4213 ( \4338 , RI8928ec0_17, \920 );
and \U$4214 ( \4339 , RI8928740_1, \918 );
or \U$4215 ( \4340 , \4129_nG1015 , \4131 , \4133 , \4135 , \4137 , \4226 , \4315 , \4325 , \4335 , \4336 , \4337 , \4338 , \4339 );
buf \U$4216 ( \4341 , \4340 );
and \U$4217 ( \4342 , \220 , \4341 );
xor \U$4218 ( \4343 , \4128 , \4342 );
xor \U$4219 ( \4344 , \4033 , \4126 );
and \U$4220 ( \4345 , \1025 , \4341 );
and \U$4221 ( \4346 , \4344 , \4345 );
xor \U$4222 ( \4347 , \4344 , \4345 );
xor \U$4223 ( \4348 , \4037 , \4124 );
and \U$4224 ( \4349 , \1033 , \4341 );
and \U$4225 ( \4350 , \4348 , \4349 );
xor \U$4226 ( \4351 , \4348 , \4349 );
xor \U$4227 ( \4352 , \4041 , \4122 );
and \U$4228 ( \4353 , \1041 , \4341 );
and \U$4229 ( \4354 , \4352 , \4353 );
xor \U$4230 ( \4355 , \4352 , \4353 );
xor \U$4231 ( \4356 , \4045 , \4120 );
and \U$4232 ( \4357 , \1049 , \4341 );
and \U$4233 ( \4358 , \4356 , \4357 );
xor \U$4234 ( \4359 , \4356 , \4357 );
xor \U$4235 ( \4360 , \4049 , \4118 );
and \U$4236 ( \4361 , \1057 , \4341 );
and \U$4237 ( \4362 , \4360 , \4361 );
xor \U$4238 ( \4363 , \4360 , \4361 );
xor \U$4239 ( \4364 , \4053 , \4116 );
and \U$4240 ( \4365 , \1065 , \4341 );
and \U$4241 ( \4366 , \4364 , \4365 );
xor \U$4242 ( \4367 , \4364 , \4365 );
xor \U$4243 ( \4368 , \4057 , \4114 );
and \U$4244 ( \4369 , \1073 , \4341 );
and \U$4245 ( \4370 , \4368 , \4369 );
xor \U$4246 ( \4371 , \4368 , \4369 );
xor \U$4247 ( \4372 , \4061 , \4112 );
and \U$4248 ( \4373 , \1081 , \4341 );
and \U$4249 ( \4374 , \4372 , \4373 );
xor \U$4250 ( \4375 , \4372 , \4373 );
xor \U$4251 ( \4376 , \4065 , \4110 );
and \U$4252 ( \4377 , \1089 , \4341 );
and \U$4253 ( \4378 , \4376 , \4377 );
xor \U$4254 ( \4379 , \4376 , \4377 );
xor \U$4255 ( \4380 , \4069 , \4108 );
and \U$4256 ( \4381 , \1097 , \4341 );
and \U$4257 ( \4382 , \4380 , \4381 );
xor \U$4258 ( \4383 , \4380 , \4381 );
xor \U$4259 ( \4384 , \4073 , \4106 );
and \U$4260 ( \4385 , \1105 , \4341 );
and \U$4261 ( \4386 , \4384 , \4385 );
xor \U$4262 ( \4387 , \4384 , \4385 );
xor \U$4263 ( \4388 , \4077 , \4104 );
and \U$4264 ( \4389 , \1113 , \4341 );
and \U$4265 ( \4390 , \4388 , \4389 );
xor \U$4266 ( \4391 , \4388 , \4389 );
xor \U$4267 ( \4392 , \4081 , \4102 );
and \U$4268 ( \4393 , \1121 , \4341 );
and \U$4269 ( \4394 , \4392 , \4393 );
xor \U$4270 ( \4395 , \4392 , \4393 );
xor \U$4271 ( \4396 , \4085 , \4100 );
and \U$4272 ( \4397 , \1129 , \4341 );
and \U$4273 ( \4398 , \4396 , \4397 );
xor \U$4274 ( \4399 , \4396 , \4397 );
xor \U$4275 ( \4400 , \4089 , \4098 );
and \U$4276 ( \4401 , \1137 , \4341 );
and \U$4277 ( \4402 , \4400 , \4401 );
xor \U$4278 ( \4403 , \4400 , \4401 );
xor \U$4279 ( \4404 , \4093 , \4096 );
and \U$4280 ( \4405 , \1144 , \4341 );
and \U$4281 ( \4406 , \4404 , \4405 );
and \U$4282 ( \4407 , \4403 , \4406 );
or \U$4283 ( \4408 , \4402 , \4407 );
and \U$4284 ( \4409 , \4399 , \4408 );
or \U$4285 ( \4410 , \4398 , \4409 );
and \U$4286 ( \4411 , \4395 , \4410 );
or \U$4287 ( \4412 , \4394 , \4411 );
and \U$4288 ( \4413 , \4391 , \4412 );
or \U$4289 ( \4414 , \4390 , \4413 );
and \U$4290 ( \4415 , \4387 , \4414 );
or \U$4291 ( \4416 , \4386 , \4415 );
and \U$4292 ( \4417 , \4383 , \4416 );
or \U$4293 ( \4418 , \4382 , \4417 );
and \U$4294 ( \4419 , \4379 , \4418 );
or \U$4295 ( \4420 , \4378 , \4419 );
and \U$4296 ( \4421 , \4375 , \4420 );
or \U$4297 ( \4422 , \4374 , \4421 );
and \U$4298 ( \4423 , \4371 , \4422 );
or \U$4299 ( \4424 , \4370 , \4423 );
and \U$4300 ( \4425 , \4367 , \4424 );
or \U$4301 ( \4426 , \4366 , \4425 );
and \U$4302 ( \4427 , \4363 , \4426 );
or \U$4303 ( \4428 , \4362 , \4427 );
and \U$4304 ( \4429 , \4359 , \4428 );
or \U$4305 ( \4430 , \4358 , \4429 );
and \U$4306 ( \4431 , \4355 , \4430 );
or \U$4307 ( \4432 , \4354 , \4431 );
and \U$4308 ( \4433 , \4351 , \4432 );
or \U$4309 ( \4434 , \4350 , \4433 );
and \U$4310 ( \4435 , \4347 , \4434 );
or \U$4311 ( \4436 , \4346 , \4435 );
xor \U$4312 ( \4437 , \4343 , \4436 );
buf \U$4313 ( \4438 , \4437 );
buf \U$4315 ( \4439 , \4438 );
xor \U$4316 ( \4440 , \4347 , \4434 );
buf \U$4317 ( \4441 , \4440 );
buf \U$4319 ( \4442 , \4441 );
xor \U$4320 ( \4443 , \4351 , \4432 );
buf \U$4321 ( \4444 , \4443 );
buf \U$4323 ( \4445 , \4444 );
xor \U$4324 ( \4446 , \4355 , \4430 );
buf \U$4325 ( \4447 , \4446 );
buf \U$4327 ( \4448 , \4447 );
xor \U$4328 ( \4449 , \4359 , \4428 );
buf \U$4329 ( \4450 , \4449 );
buf \U$4331 ( \4451 , \4450 );
xor \U$4332 ( \4452 , \4363 , \4426 );
buf \U$4333 ( \4453 , \4452 );
buf \U$4335 ( \4454 , \4453 );
xor \U$4336 ( \4455 , \4367 , \4424 );
buf \U$4337 ( \4456 , \4455 );
buf \U$4339 ( \4457 , \4456 );
xor \U$4340 ( \4458 , \4371 , \4422 );
buf \U$4341 ( \4459 , \4458 );
buf \U$4343 ( \4460 , \4459 );
xor \U$4344 ( \4461 , \4375 , \4420 );
buf \U$4345 ( \4462 , \4461 );
buf \U$4347 ( \4463 , \4462 );
xor \U$4348 ( \4464 , \4379 , \4418 );
buf \U$4349 ( \4465 , \4464 );
buf \U$4351 ( \4466 , \4465 );
xor \U$4352 ( \4467 , \4383 , \4416 );
buf \U$4353 ( \4468 , \4467 );
buf \U$4355 ( \4469 , \4468 );
xor \U$4356 ( \4470 , \4387 , \4414 );
buf \U$4357 ( \4471 , \4470 );
buf \U$4359 ( \4472 , \4471 );
xor \U$4360 ( \4473 , \4391 , \4412 );
buf \U$4361 ( \4474 , \4473 );
buf \U$4363 ( \4475 , \4474 );
xor \U$4364 ( \4476 , \4395 , \4410 );
buf \U$4365 ( \4477 , \4476 );
buf \U$4367 ( \4478 , \4477 );
xor \U$4368 ( \4479 , \4399 , \4408 );
buf \U$4369 ( \4480 , \4479 );
buf \U$4371 ( \4481 , \4480 );
xor \U$4372 ( \4482 , \4403 , \4406 );
buf \U$4373 ( \4483 , \4482 );
buf \U$4375 ( \4484 , \4483 );
xor \U$4376 ( \4485 , \4404 , \4405 );
buf \U$4377 ( \4486 , \4485 );
buf \U$4379 ( \4487 , \4486 );
xor \U$4380 ( \4488 , \4094 , \4095 );
buf \U$4381 ( \4489 , \4488 );
buf \U$4383 ( \4490 , \4489 );
xor \U$4384 ( \4491 , \3795 , \3796 );
buf \U$4385 ( \4492 , \4491 );
buf \U$4387 ( \4493 , \4492 );
xor \U$4388 ( \4494 , \3508 , \3509 );
buf \U$4389 ( \4495 , \4494 );
buf \U$4391 ( \4496 , \4495 );
xor \U$4392 ( \4497 , \3233 , \3234 );
buf \U$4393 ( \4498 , \4497 );
buf \U$4395 ( \4499 , \4498 );
xor \U$4396 ( \4500 , \2970 , \2971 );
buf \U$4397 ( \4501 , \4500 );
buf \U$4399 ( \4502 , \4501 );
xor \U$4400 ( \4503 , \2719 , \2720 );
buf \U$4401 ( \4504 , \4503 );
buf \U$4403 ( \4505 , \4504 );
xor \U$4404 ( \4506 , \2480 , \2481 );
buf \U$4405 ( \4507 , \4506 );
buf \U$4407 ( \4508 , \4507 );
xor \U$4408 ( \4509 , \2253 , \2254 );
buf \U$4409 ( \4510 , \4509 );
buf \U$4411 ( \4511 , \4510 );
xor \U$4412 ( \4512 , \2038 , \2039 );
buf \U$4413 ( \4513 , \4512 );
buf \U$4415 ( \4514 , \4513 );
xor \U$4416 ( \4515 , \1835 , \1836 );
buf \U$4417 ( \4516 , \4515 );
buf \U$4419 ( \4517 , \4516 );
endmodule

