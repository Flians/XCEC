//
// Conformal-LEC Version 20.10-d207 (02-Sep-2020)
//
module top(RIdec64b8_720,RIbc62af0_23,RIbc62a78_22,RIbc62a00_21,RIbc62988_20,RIbc62910_19,RIbc62898_18,RIbc62820_17,RIbc627a8_16,
        RIbc62730_15,RIbc626b8_14,RIbc62640_13,RIdec37b8_688,RIfc8daa0_6634,RIdec0ab8_656,RIfc56348_6003,RIdebddb8_624,RIdebb0b8_592,RIdeb83b8_560,
        RIfc98798_6757,RIdeb29b8_496,RIfcbd098_7173,RIdeafcb8_464,RIfc8dc08_6635,RIdeacb80_432,RIdea6280_400,RIde9f980_368,RIfcd6868_7463,RIfc8ded8_6637,
        RIfc7dd80_6454,RIfc56618_6005,RIde92e10_306,RIde8f300_288,RIde8b160_268,RIde86fc0_248,RIde82ad8_227,RIfc8e040_6638,RIfcd96d0_7496,RIfca1e10_6864,
        RIfcbd200_7174,RIe16c5c0_2610,RIe16a298_2585,RIe168ab0_2568,RIe1664b8_2541,RIe1637b8_2509,RIee37f00_5095,RIe160ab8_2477,RIfc8ea18_6645,RIe15ddb8_2445,
        RIe1583b8_2381,RIe1556b8_2349,RIfe9f828_8159,RIe1529b8_2317,RIfe9f990_8160,RIe14fcb8_2285,RIfcbd368_7175,RIe14cfb8_2253,RIe14a2b8_2221,RIe1475b8_2189,
        RIfc8ee50_6648,RIfc45278_5809,RIfc98360_6754,RIfca2248_6867,RIe141d20_2126,RIe13f9f8_2101,RIdf3d900_2077,RIdf3b470_2051,RIfcd6ca0_7466,RIee2ff08_5004,
        RIfc8ece8_6647,RIee2dd48_4980,RIdf36718_1996,RIdf34120_1969,RIdf31f60_1945,RIfe9f6c0_8158,RIfcb4560_7074,RIfc45db8_5817,RIfc8e1a8_6639,RIfc7d678_6449,
        RIdf2aee0_1865,RIdf28ff0_1843,RIdf26e30_1819,RIdf25378_1800,RIfcb43f8_7073,RIfc8e748_6643,RIdf23488_1778,RIfcc2c00_7238,RIdf21e08_1762,RIdf20788_1746,
        RIdf1b760_1689,RIdf1a248_1674,RIdf18088_1650,RIdf15388_1618,RIdf12688_1586,RIdf0f988_1554,RIdf0cc88_1522,RIdf09f88_1490,RIdf07288_1458,RIdf04588_1426,
        RIdefeb88_1362,RIdefbe88_1330,RIdef9188_1298,RIdef6488_1266,RIdef3788_1234,RIdef0a88_1202,RIdeedd88_1170,RIdeeb088_1138,RIfc8efb8_6649,RIfc44e40_5806,
        RIfc57860_6018,RIfca23b0_6868,RIfe9faf8_8161,RIdee3900_1053,RIdee1740_1029,RIdedf6e8_1006,RIfcbd4d0_7176,RIee22678_4850,RIfc98090_6752,RIee21598_4838,
        RIfe9fc60_8162,RIded80c8_922,RIfe9fdc8_8163,RIded3be0_873,RIded18b8_848,RIdecebb8_816,RIdecbeb8_784,RIdec91b8_752,RIdeb56b8_528,RIde99080_336,
        RIe16f2c0_2642,RIe15b0b8_2413,RIe1448b8_2157,RIdf392b0_2027,RIdf2d910_1895,RIdf1e190_1719,RIdf01888_1394,RIdee8388_1106,RIdedd0f0_979,RIde7efc8_209,
        RIe19e750_3180,RIbc625c8_12,RIbc62550_11,RIbc624d8_10,RIbc62460_9,RIbc623e8_8,RIbc62370_7,RIbc622f8_6,RIbc62280_5,RIbc62208_4,
        RIbc62190_3,RIbc62118_2,RIe19ba50_3148,RIfc479d8_5837,RIe198d50_3116,RIfe9f558_8157,RIe196050_3084,RIe193350_3052,RIe190650_3020,RIe18ac50_2956,
        RIe187f50_2924,RIfc47870_5836,RIe185250_2892,RIf142ef8_5221,RIe182550_2860,RIe17f850_2828,RIe17cb50_2796,RIfcb5208_7083,RIfcbc6c0_7166,RIe177588_2735,
        RIe176610_2724,RIf13fdc0_5186,RIfe9f3f0_8156,RIfce40f8_7617,RIfc47708_5835,RIfc47438_5833,RIfca15a0_6858,RIfc99170_6764,RIe1745b8_2701,RIfc8cc90_6624,
        RIfc556a0_5994,RIfc7ee60_6466,RIfce8e50_7672,RIfe9f288_8155,RIe224aa8_4707,RIfc55808_5995,RIe221da8_4675,RIfcb50a0_7082,RIe21f0a8_4643,RIe2196a8_4579,
        RIe2169a8_4547,RIfcbc828_7167,RIe213ca8_4515,RIfc47000_5830,RIe210fa8_4483,RIfcbc990_7168,RIe20e2a8_4451,RIe20b5a8_4419,RIe2088a8_4387,RIfc46bc8_5827,
        RIfcd6598_7461,RIe2032e0_4326,RIe2016c0_4306,RIfc98ea0_6762,RIfc7eb90_6464,RIfce0318_7573,RIfcbcaf8_7169,RIfc8cf60_6626,RIfcb4dd0_7080,RIe1fd340_4258,
        RIe1fc260_4246,RIf15cf38_5517,RIfe9f120_8154,RIfc7ea28_6463,RIfc8d0c8_6627,RIfcbcc60_7170,RIfc98bd0_6760,RIfce2d48_7603,RIe1fb018_4233,RIfc55f10_6000,
        RIfc7e8c0_6462,RIfc8d230_6628,RIe1f6590_4180,RIfce58e0_7634,RIfc468f8_5825,RIfcc2ed0_7240,RIe1f4100_4154,RIfceedf0_7740,RIfc8d398_6629,RIfc8d500_6630,
        RIe1eef70_4096,RIe1ec810_4068,RIe1e9b10_4036,RIe1e6e10_4004,RIe1e4110_3972,RIe1e1410_3940,RIe1de710_3908,RIe1dba10_3876,RIe1d8d10_3844,RIe1d3310_3780,
        RIe1d0610_3748,RIe1cd910_3716,RIe1cac10_3684,RIe1c7f10_3652,RIe1c5210_3620,RIe1c2510_3588,RIe1bf810_3556,RIf14d0b0_5336,RIfe9efb8_8153,RIe1ba248_3495,
        RIe1b8088_3471,RIfec4dd0_8360,RIfec50a0_8362,RIe1b5ec8_3447,RIe1b46e0_3430,RIfcb4998_7077,RIfcb4c68_7079,RIfec5370_8364,RIfe9ee50_8152,RIfcbcdc8_7171,
        RIfc46358_5821,RIfec5208_8363,RIfec4f38_8361,RIe1a9b50_3308,RIe1a6e50_3276,RIe1a4150_3244,RIe1a1450_3212,RIe18d950_2988,RIe179e50_2764,RIe2277a8_4739,
        RIe21c3a8_4611,RIe205ba8_4355,RIe1ffc08_4287,RIe1f8fc0_4210,RIe1f1b08_4127,RIe1d6010_3812,RIe1bcb10_3524,RIe1af988_3375,RIe171fc0_2674,RIdec6080_717,
        RIdec3380_685,RIee204b8_4826,RIdec0680_653,RIfcd70d8_7469,RIdebd980_621,RIdebac80_589,RIdeb7f80_557,RIfcbe448_7187,RIdeb2580_493,RIfcb3480_7062,
        RIdeaf880_461,RIfc43928_5791,RIdeac1a8_429,RIdea58a8_397,RIde9efa8_365,RIfcd88c0_7486,RIee1c408_4780,RIfcc77f0_7292,RIfea04d0_8168,RIde92438_303,
        RIde8ec70_286,RIde8aad0_266,RIde86930_246,RIfca31c0_6878,RIfc59a20_6042,RIfcd1de0_7410,RIfc91448_6675,RIfc97280_6742,RIe16c188_2607,RIfc97118_6741,
        RIe168948_2567,RIe166080_2538,RIe163380_2506,RIee37ac8_5092,RIe160680_2474,RIfcd1c78_7409,RIe15d980_2442,RIe157f80_2378,RIe155280_2346,RIfc3f530_5746,
        RIe152580_2314,RIee35368_5064,RIe14f880_2282,RIfc7a3d8_6413,RIe14cb80_2250,RIe149e80_2218,RIe147180_2186,RIfc42b18_5781,RIfc7a270_6412,RIfc5a560_6050,
        RIfc96b78_6737,RIfea6fb0_8216,RIe13f5c0_2098,RIdf3d4c8_2074,RIdf3b038_2048,RIfce5bb0_7636,RIee2fc38_5002,RIfc91cb8_6681,RIee2d910_4977,RIdf362e0_1993,
        RIdf33e50_1967,RIdf31c90_1943,RIdf2fda0_1921,RIfc43658_5789,RIfc59e58_6045,RIfc96fb0_6740,RIfc7ac48_6419,RIfea0368_8167,RIdf28bb8_1840,RIdf26cc8_1818,
        RIdf25210_1799,RIfc91718_6677,RIfcb3318_7061,RIfc919e8_6679,RIfc91880_6678,RIfc430b8_5785,RIdf20350_1743,RIfc7a978_6417,RIdf19e10_1671,RIdf17c50_1647,
        RIdf14f50_1615,RIdf12250_1583,RIdf0f550_1551,RIdf0c850_1519,RIdf09b50_1487,RIdf06e50_1455,RIdf04150_1423,RIdefe750_1359,RIdefba50_1327,RIdef8d50_1295,
        RIdef6050_1263,RIdef3350_1231,RIdef0650_1199,RIdeed950_1167,RIdeeac50_1135,RIfcd1b10_7408,RIfc968a8_6735,RIfc91f88_6683,RIfcdfc10_7568,RIfea99e0_8246,
        RIdee3630_1051,RIdee1308_1026,RIdedf2b0_1003,RIfcc7d90_7296,RIfcd85f0_7484,RIfce3888_7611,RIfc5a830_6052,RIdeda3f0_947,RIfea9878_8245,RIded5f08_898,
        RIded37a8_870,RIded1480_845,RIdece780_813,RIdecba80_781,RIdec8d80_749,RIdeb5280_525,RIde986a8_333,RIe16ee88_2639,RIe15ac80_2410,RIe144480_2154,
        RIdf38e78_2024,RIdf2d4d8_1892,RIdf1dd58_1716,RIdf01450_1391,RIdee7f50_1103,RIdedccb8_976,RIde7e5f0_206,RIe19e318_3177,RIe19b618_3145,RIfc8f3f0_6652,
        RIe198918_3113,RIf144b18_5241,RIe195c18_3081,RIe192f18_3049,RIe190218_3017,RIe18a818_2953,RIe187b18_2921,RIf143d08_5231,RIe184e18_2889,RIfcb3cf0_7068,
        RIe182118_2857,RIe17f418_2825,RIe17c718_2793,RIfc448a0_5802,RIf141170_5200,RIfc7c9d0_6440,RIfea0098_8165,RIfc57e00_6022,RIf13f550_5180,RIfcd6e08_7467,
        RIee3d900_5159,RIfc8f6c0_6654,RIfce0048_7571,RIfca27e8_6871,RIe1742e8_2699,RIfc7c700_6438,RIfc8f990_6656,RIfce9828_7679,RIfc583a0_6026,RIf16cdc0_5698,
        RIe224670_4704,RIf16c118_5689,RIe221970_4672,RIfc58508_6027,RIe21ec70_4640,RIe219270_4576,RIe216570_4544,RIfc3ff08_5753,RIe213870_4512,RIf1696e8_5659,
        RIe210b70_4480,RIfc58940_6030,RIe20de70_4448,RIe20b170_4416,RIe208470_4384,RIfc8fc60_6658,RIfc97820_6746,RIe202ea8_4323,RIe201288_4303,RIfcc27c8_7235,
        RIfcdfee0_7570,RIfc44198_5797,RIfc58670_6028,RIf1608e0_5558,RIf15e9f0_5536,RIfe9ff30_8164,RIe1fc0f8_4245,RIfc7be90_6432,RIf15bb88_5503,RIfcd8cf8_7489,
        RIfcd8e60_7490,RIfca2d88_6875,RIfcbdea8_7183,RIfcb3a20_7066,RIe1fabe0_4230,RIfc90098_6661,RIfc90200_6662,RIfcd20b0_7412,RIe1f6158_4177,RIfc904d0_6664,
        RIfca2ef0_6876,RIfc97550_6744,RIe1f3e30_4152,RIfc59048_6035,RIfc907a0_6666,RIfc90638_6665,RIe1eeb38_4093,RIe1ec3d8_4065,RIe1e96d8_4033,RIe1e69d8_4001,
        RIe1e3cd8_3969,RIe1e0fd8_3937,RIe1de2d8_3905,RIe1db5d8_3873,RIe1d88d8_3841,RIe1d2ed8_3777,RIe1d01d8_3745,RIe1cd4d8_3713,RIe1ca7d8_3681,RIe1c7ad8_3649,
        RIe1c4dd8_3617,RIe1c20d8_3585,RIe1bf3d8_3553,RIfcc73b8_7289,RIfce3cc0_7614,RIe1b9e10_3492,RIe1b7c50_3468,RIfcd6f70_7468,RIf149e10_5300,RIe1b5a90_3444,
        RIfea0200_8166,RIfc90bd8_6669,RIfcdfd78_7569,RIe1b2ef8_3413,RIe1b15a8_3395,RIfc973e8_6743,RIfcc7520_7290,RIe1acdf0_3344,RIe1ab608_3327,RIe1a9718_3305,
        RIe1a6a18_3273,RIe1a3d18_3241,RIe1a1018_3209,RIe18d518_2985,RIe179a18_2761,RIe227370_4736,RIe21bf70_4608,RIe205770_4352,RIe1ff7d0_4284,RIe1f8b88_4207,
        RIe1f16d0_4124,RIe1d5bd8_3809,RIe1bc6d8_3521,RIe1af550_3372,RIe171b88_2671,RIdec5108_706,RIdec2408_674,RIfc93608_6699,RIdebf708_642,RIfc934a0_6698,
        RIdebca08_610,RIdeb9d08_578,RIdeb7008_546,RIfcdf7d8_7565,RIdeb1608_482,RIfc78218_6389,RIdeae908_450,RIfcc8498_7301,RIdea9d90_418,RIdea3490_386,
        RIde9cb90_354,RIee1cc78_4786,RIee1bb98_4774,RIee1b328_4768,RIee1aab8_4762,RIde909f8_295,RIde8d578_279,RIfea8ea0_8238,RIde85238_239,RIde813e0_220,
        RIfc938d8_6701,RIfce5e80_7638,RIfcbfd98_7205,RIfce8ce8_7671,RIe16b4e0_2598,RIfea8d38_8237,RIfea9f80_8250,RIe165108_2527,RIe162408_2495,RIfc779a8_6383,
        RIe15f708_2463,RIfe9dc08_8139,RIe15ca08_2431,RIe157008_2367,RIe154308_2335,RIfea7550_8220,RIe151608_2303,RIfcd6160_7458,RIe14e908_2271,RIfcd1408_7403,
        RIe14bc08_2239,RIe148f08_2207,RIe146208_2175,RIfceb718_7701,RIfcb19c8_7043,RIfc93e78_6705,RIfce7938_7657,RIe140da8_2115,RIdf3ecb0_2091,RIdf3c988_2066,
        RIfe9daa0_8138,RIfce8478_7665,RIfcdbf98_7525,RIfc776d8_6381,RIfc93fe0_6706,RIdf354d0_1983,RIdf33040_1957,RIdf30fe8_1934,RIdf2ee28_1910,RIee2ba20_4955,
        RIfc93ba8_6703,RIfc77de0_6386,RIee27ad8_4910,RIfe9d668_8135,RIfea8bd0_8236,RIdf26458_1812,RIfe9d7d0_8136,RIfcb1c98_7045,RIee26cc8_4900,RIdf22ab0_1771,
        RIfcc0068_7207,RIdf21598_1756,RIdf1f6a8_1734,RIdf1aef0_1683,RIfe9d938_8137,RIdf16cd8_1636,RIdf13fd8_1604,RIdf112d8_1572,RIdf0e5d8_1540,RIdf0b8d8_1508,
        RIdf08bd8_1476,RIdf05ed8_1444,RIdf031d8_1412,RIdefd7d8_1348,RIdefaad8_1316,RIdef7dd8_1284,RIdef50d8_1252,RIdef23d8_1220,RIdeef6d8_1188,RIdeec9d8_1156,
        RIdee9cd8_1124,RIfc942b0_6708,RIfcde6f8_7553,RIfcd1138_7401,RIfcde860_7554,RIdee4878_1064,RIdee2af0_1043,RIdee0a98_1020,RIdede8d8_996,RIfc5c9f0_6076,
        RIee22240_4847,RIfcc8768_7303,RIee21160_4835,RIded95e0_937,RIded7150_911,RIded5260_889,RIfea76b8_8221,RIded0508_834,RIdecd808_802,RIdecab08_770,
        RIdec7e08_738,RIdeb4308_514,RIde96290_322,RIe16df10_2628,RIe159d08_2399,RIe143508_2143,RIdf37f00_2013,RIdf2c560_1881,RIdf1cde0_1705,RIdf004d8_1380,
        RIdee6fd8_1092,RIdedbd40_965,RIde7c1d8_195,RIe19d3a0_3166,RIe19a6a0_3134,RIfcb2c10_7056,RIe1979a0_3102,RIfc923c0_6686,RIe194ca0_3070,RIe191fa0_3038,
        RIe18f2a0_3006,RIe1898a0_2942,RIe186ba0_2910,RIfc422a8_5775,RIe183ea0_2878,RIfcbecb8_7193,RIe1811a0_2846,RIe17e4a0_2814,RIe17b7a0_2782,RIf142250_5212,
        RIf140bd0_5196,RIfec43f8_8353,RIe175968_2715,RIfc79b68_6407,RIf13efb0_5176,RIfc92528_6687,RIfcb2aa8_7055,RIfcd8320_7482,RIfcea200_7686,RIfc79898_6405,
        RIe1734d8_2689,RIfcd7948_7475,RIfcd7678_7473,RIf16e170_5712,RIfc927f8_6689,RIfc92960_6690,RIe2236f8_4693,RIfc795c8_6403,RIe2209f8_4661,RIf16ad68_5675,
        RIe21dcf8_4629,RIe2182f8_4565,RIe2155f8_4533,RIfe9d398_8133,RIe2128f8_4501,RIfcdb9f8_7521,RIe20fbf8_4469,RIfc41d08_5771,RIe20cef8_4437,RIe20a1f8_4405,
        RIe2074f8_4373,RIfcd7510_7472,RIf166010_5620,RIfe9d230_8132,RIe2008b0_4296,RIf165098_5609,RIfc41ba0_5770,RIfc41a38_5769,RIfc92c30_6692,RIfc418d0_5768,
        RIfc79190_6400,RIe1fcad0_4252,RIfec4560_8354,RIfc79028_6399,RIfcbf258_7197,RIfcc1df0_7228,RIfcd81b8_7481,RIfc92d98_6693,RIfc5b4d8_6061,RIfcd77e0_7474,
        RIe1fa0a0_4222,RIf156188_5439,RIfe9d500_8134,RIf1546d0_5420,RIe1f5348_4167,RIfec4830_8356,RIfec46c8_8355,RIf1508f0_5376,RIe1f3020_4142,RIfce3180_7606,
        RIfce8fb8_7673,RIfcbf690_7200,RIe1edd28_4083,RIe1eb460_4054,RIe1e8760_4022,RIe1e5a60_3990,RIe1e2d60_3958,RIe1e0060_3926,RIe1dd360_3894,RIe1da660_3862,
        RIe1d7960_3830,RIe1d1f60_3766,RIe1cf260_3734,RIe1cc560_3702,RIe1c9860_3670,RIe1c6b60_3638,RIe1c3e60_3606,RIe1c1160_3574,RIe1be460_3542,RIfe9d0c8_8131,
        RIfe9cc90_8128,RIe1b9168_3483,RIe1b7110_3460,RIf14a3b0_5304,RIfe9cb28_8127,RIfe9cf60_8130,RIfe9c9c0_8126,RIfce2208_7595,RIfce9558_7677,RIfe9c858_8125,
        RIfe9cdf8_8129,RIf147110_5268,RIf146468_5259,RIe1ac2b0_3336,RIe1aaac8_3319,RIe1a87a0_3294,RIe1a5aa0_3262,RIe1a2da0_3230,RIe1a00a0_3198,RIe18c5a0_2974,
        RIe178aa0_2750,RIe2263f8_4725,RIe21aff8_4597,RIe2047f8_4341,RIe1fe858_4273,RIe1f7c10_4196,RIe1f0758_4113,RIe1d4c60_3798,RIe1bb760_3510,RIe1ae5d8_3361,
        RIe170c10_2660,RIdec4190_695,RIdec1490_663,RIfceaa70_7692,RIdebe790_631,RIfc954f8_6721,RIdebba90_599,RIdeb8d90_567,RIdeb6090_535,RIfcebb50_7704,
        RIdeb0690_471,RIee1e190_4801,RIdead990_439,RIfcdf0d0_7560,RIdea7978_407,RIdea1078_375,RIde9a778_343,RIee1c840_4783,RIfc957c8_6723,RIfcc8e70_7308,
        RIfc5e610_6096,RIfe9e8b0_8148,RIde8c1c8_273,RIde88028_253,RIde83b40_232,RIfcb0bb8_7033,RIfca4b10_6896,RIfc75d88_6363,RIfca4c78_6897,RIfc95390_6720,
        RIe16a9a0_2590,RIfcc8fd8_7309,RIe166e90_2548,RIe164190_2516,RIe161490_2484,RIfe9e748_8147,RIe15e790_2452,RIfc74f78_6353,RIe15ba90_2420,RIe156090_2356,
        RIe153390_2324,RIfc3ecc0_5740,RIe150690_2292,RIfce8b80_7670,RIe14d990_2260,RIfca6730_6916,RIe14ac90_2228,RIe147f90_2196,RIe145290_2164,RIfcee2b0_7732,
        RIfc5f2b8_6105,RIfc753b0_6356,RIfc74b40_6350,RIe140268_2107,RIdf3e170_2083,RIdf3be48_2058,RIdf39c88_2034,RIfcc1c88_7227,RIfcc1850_7224,RIfc965d8_6733,
        RIfc96038_6729,RIdf34828_1974,RIdf327d0_1951,RIdf301d8_1924,RIdf2e2e8_1902,RIfc5e778_6097,RIfcd0328_7391,RIfc757e8_6359,RIfcee6e8_7735,RIdf296f8_1848,
        RIdf273d0_1823,RIdf257b0_1803,RIdf23b90_1783,RIfc95d68_6727,RIfceda40_7726,RIfe9eb80_8150,RIfc75518_6357,RIfcd01c0_7390,RIdf1eb68_1726,RIfe9ece8_8151,
        RIfe9ea18_8149,RIdf15d60_1625,RIdf13060_1593,RIdf10360_1561,RIdf0d660_1529,RIdf0a960_1497,RIdf07c60_1465,RIdf04f60_1433,RIdf02260_1401,RIdefc860_1337,
        RIdef9b60_1305,RIdef6e60_1273,RIdef4160_1241,RIdef1460_1209,RIdeee760_1177,RIdeeba60_1145,RIdee8d60_1113,RIfc961a0_6730,RIfc96308_6731,RIfc5ee80_6102,
        RIfce6150_7640,RIdee42d8_1060,RIdee1e48_1034,RIdee00c0_1013,RIdeddac8_986,RIfc96470_6732,RIfc75248_6355,RIfc74ca8_6351,RIfcb0618_7029,RIded8938_928,
        RIded6610_903,RIded4450_879,RIded2290_855,RIdecf590_823,RIdecc890_791,RIdec9b90_759,RIdec6e90_727,RIdeb3390_503,RIde93e78_311,RIe16cf98_2617,
        RIe158d90_2388,RIe142590_2132,RIdf36f88_2002,RIdf2b5e8_1870,RIdf1be68_1694,RIdeff560_1369,RIdee6060_1081,RIdedadc8_954,RIde79dc0_184,RIe19c428_3155,
        RIe199728_3123,RIfe9e310_8144,RIe196a28_3091,RIfcc04a0_7210,RIe193d28_3059,RIe191028_3027,RIe18e328_2995,RIe188928_2931,RIe185c28_2899,RIfce1830_7588,
        RIe182f28_2867,RIfe9e478_8145,RIe180228_2835,RIe17d528_2803,RIe17a828_2771,RIf141878_5205,RIfcb12c0_7038,RIfc94418_6709,RIe174f90_2708,RIfc77408_6379,
        RIf13ea10_5172,RIfcdc100_7526,RIfc94580_6710,RIfc946e8_6711,RIfced338_7721,RIfce5fe8_7639,RIe172998_2681,RIfcdc268_7527,RIfcddff0_7548,RIfcc0608_7211,
        RIfce7230_7652,RIfc40340_5756,RIe222780_4682,RIfcdd618_7541,RIe21fa80_4650,RIfcd0b98_7397,RIe21cd80_4618,RIe217380_4554,RIe214680_4522,RIfec4998_8357,
        RIe211980_4490,RIf168608_5647,RIe20ec80_4458,RIfcc0770_7212,RIe20bf80_4426,RIe209280_4394,RIe206580_4362,RIfce2370_7596,RIfcee580_7734,RIfec4c68_8359,
        RIfec4b00_8358,RIfc949b8_6713,RIfcebcb8_7705,RIf162938_5581,RIf1612b8_5565,RIfccd088_7355,RIfcc08d8_7213,RIfe9e040_8142,RIfe9e1a8_8143,RIfcead40_7694,
        RIf15ad78_5493,RIfc94c88_6715,RIfccc3e0_7346,RIfc765f8_6369,RIfc94df0_6716,RIfcc0a40_7214,RIe1f9998_4217,RIfcc8d08_7307,RIfce8748_7667,RIfceb2e0_7698,
        RIe1f4970_4160,RIf152510_5396,RIf1512c8_5383,RIfcb0ff0_7036,RIe1f24e0_4134,RIfc761c0_6366,RIfc950c0_6718,RIfcc0e78_7217,RIe1ed1e8_4075,RIe1ea4e8_4043,
        RIe1e77e8_4011,RIe1e4ae8_3979,RIe1e1de8_3947,RIe1df0e8_3915,RIe1dc3e8_3883,RIe1d96e8_3851,RIe1d69e8_3819,RIe1d0fe8_3755,RIe1ce2e8_3723,RIe1cb5e8_3691,
        RIe1c88e8_3659,RIe1c5be8_3627,RIe1c2ee8_3595,RIe1c01e8_3563,RIe1bd4e8_3531,RIf14bfd0_5324,RIf14ac20_5310,RIfe9ded8_8141,RIe1b65d0_3452,RIfcecd98_7717,
        RIfc76490_6368,RIe1b4c80_3434,RIe1b38d0_3420,RIfcc0fe0_7218,RIfceaea8_7695,RIe1b1f80_3402,RIe1b0360_3382,RIfcd0760_7394,RIf145ec8_5255,RIfe9e5e0_8146,
        RIfe9dd70_8140,RIe1a7828_3283,RIe1a4b28_3251,RIe1a1e28_3219,RIe19f128_3187,RIe18b628_2963,RIe177b28_2739,RIe225480_4714,RIe21a080_4586,RIe203880_4330,
        RIe1fd8e0_4262,RIe1f6c98_4185,RIe1ef7e0_4102,RIe1d3ce8_3787,RIe1ba7e8_3499,RIe1ad660_3350,RIe16fc98_2649,RIdec6788_722,RIdec3a88_690,RIee20788_4828,
        RIdec0d88_658,RIee1f810_4817,RIdebe088_626,RIdebb388_594,RIdeb8688_562,RIfc9b1c8_6787,RIdeb2c88_498,RIfce1f38_7593,RIdeaff88_466,RIfc892e8_6583,
        RIdead210_434,RIdea6910_402,RIdea0010_370,RIee1d650_4793,RIee1c570_4781,RIee1b5f8_4770,RIee1aef0_4765,RIfe99888_8091,RIfe99450_8088,RIfe99720_8090,
        RIfe995b8_8089,RIde83168_229,RIfcc43e8_7255,RIfcd5a58_7453,RIfc89450_6584,RIfcc5798_7269,RIe16c890_2612,RIe16a568_2587,RIe168d80_2570,RIe166788_2543,
        RIe163a88_2511,RIfc83618_6517,RIe160d88_2479,RIee36718_5078,RIe15e088_2447,RIe158688_2383,RIe155988_2351,RIfc3f800_5748,RIe152c88_2319,RIfc895b8_6585,
        RIe14ff88_2287,RIfc51cf8_5953,RIe14d288_2255,RIe14a588_2223,RIe147888_2191,RIee34990_5057,RIee338b0_5045,RIfc831e0_6514,RIfcd3b68_7431,RIe141ff0_2128,
        RIe13fcc8_2103,RIdf3dbd0_2079,RIdf3b740_2053,RIfcb6f90_7104,RIee301d8_5006,RIfcba938_7145,RIee2e018_4982,RIdf369e8_1998,RIdf343f0_1971,RIdf32230_1947,
        RIfe99e28_8095,RIfc83078_6513,RIfcb6e28_7103,RIfc9ad90_6784,RIfcbad70_7148,RIdf2b1b0_1867,RIdf292c0_1845,RIfe99b58_8093,RIfe999f0_8092,RIfc9ac28_6783,
        RIfc4a9a8_5871,RIdf23758_1780,RIfc82da8_6511,RIdf220d8_1764,RIdf20a58_1748,RIdf1ba30_1691,RIfe99cc0_8094,RIdf18358_1652,RIdf15658_1620,RIdf12958_1588,
        RIdf0fc58_1556,RIdf0cf58_1524,RIdf0a258_1492,RIdf07558_1460,RIdf04858_1428,RIdefee58_1364,RIdefc158_1332,RIdef9458_1300,RIdef6758_1268,RIdef3a58_1236,
        RIdef0d58_1204,RIdeee058_1172,RIdeeb358_1140,RIee25918_4886,RIee24b08_4876,RIfc52568_5959,RIfc826a0_6506,RIdee5958_1076,RIdee3bd0_1055,RIfe99f90_8096,
        RIdedf9b8_1008,RIfce4800_7622,RIfc89b58_6589,RIfc9f3e0_6834,RIfc82538_6505,RIdeda828_950,RIded8398_924,RIfeabe70_8272,RIded3eb0_875,RIded1b88_850,
        RIdecee88_818,RIdecc188_786,RIdec9488_754,RIdeb5988_530,RIde99710_338,RIe16f590_2644,RIe15b388_2415,RIe144b88_2159,RIdf39580_2029,RIdf2dbe0_1897,
        RIdf1e460_1721,RIdf01b58_1396,RIdee8658_1108,RIdedd3c0_981,RIde7f658_211,RIe19ea20_3182,RIe19bd20_3150,RIf145928_5251,RIe199020_3118,RIfe98910_8080,
        RIe196320_3086,RIe193620_3054,RIe190920_3022,RIe18af20_2958,RIe188220_2926,RIf143e70_5232,RIe185520_2894,RIfc95c00_6726,RIe182820_2862,RIe17fb20_2830,
        RIe17ce20_2798,RIf142520_5214,RIf141440_5202,RIe1776f0_2736,RIfeab8d0_8268,RIfcc5bd0_7272,RIfc62dc8_6147,RIee3e710_5169,RIfc9cb18_6805,RIee3c820_5147,
        RIee3b470_5133,RIee3a390_5121,RIe174888_2703,RIf170498_5737,RIfc68660_6210,RIf16e878_5717,RIfc6ea38_6281,RIfe98d48_8083,RIe224d78_4709,RIf16c280_5690,
        RIe222078_4677,RIf16b308_5679,RIe21f378_4645,RIe219978_4581,RIe216c78_4549,RIf16a390_5668,RIe213f78_4517,RIf169b20_5662,RIe211278_4485,RIf1681d0_5644,
        RIe20e578_4453,RIe20b878_4421,RIe208b78_4389,RIfcd4ae0_7442,RIfc61478_6129,RIfeab060_8262,RIe201990_4308,RIfc70ec8_6307,RIfc70928_6303,RIfcec528_7711,
        RIfcbe880_7190,RIf160d18_5561,RIf15ee28_5539,RIfe98be0_8082,RIfe98eb0_8084,RIf15d0a0_5518,RIf15bcf0_5504,RIfcd4540_7438,RIf159e00_5482,RIf1592c0_5474,
        RIf158078_5461,RIfca3a30_6884,RIfea7988_8223,RIf156728_5443,RIf155be8_5435,RIf154b08_5423,RIfe98a78_8081,RIf1538c0_5410,RIf1520d8_5393,RIf150e90_5380,
        RIe1f43d0_4156,RIf14fdb0_5368,RIfcd2380_7414,RIf14e2f8_5349,RIe1ef240_4098,RIe1ecae0_4070,RIe1e9de0_4038,RIe1e70e0_4006,RIe1e43e0_3974,RIe1e16e0_3942,
        RIe1de9e0_3910,RIe1dbce0_3878,RIe1d8fe0_3846,RIe1d35e0_3782,RIe1d08e0_3750,RIe1cdbe0_3718,RIe1caee0_3686,RIe1c81e0_3654,RIe1c54e0_3622,RIe1c27e0_3590,
        RIe1bfae0_3558,RIfc44b70_5804,RIf14bd00_5322,RIfe992e8_8087,RIfe987a8_8079,RIf14a950_5308,RIf149f78_5301,RIfe99180_8086,RIfe98640_8078,RIf149438_5293,
        RIfcec7f8_7713,RIfe984d8_8077,RIe1b1b48_3399,RIfc4b650_5880,RIfcda918_7509,RIfe98370_8076,RIfe99018_8085,RIe1a9e20_3310,RIe1a7120_3278,RIe1a4420_3246,
        RIe1a1720_3214,RIe18dc20_2990,RIe17a120_2766,RIe227a78_4741,RIe21c678_4613,RIe205e78_4357,RIe1ffed8_4289,RIe1f9290_4212,RIe1f1dd8_4129,RIe1d62e0_3814,
        RIe1bcde0_3526,RIe1afc58_3377,RIe172290_2676,RIdec6620_721,RIdec3920_689,RIfc49328_5855,RIdec0c20_657,RIfc80eb8_6489,RIdebdf20_625,RIdebb220_593,
        RIdeb8520_561,RIfc80648_6483,RIdeb2b20_497,RIfc8b340_6606,RIdeafe20_465,RIfc491c0_5854,RIdeacec8_433,RIdea65c8_401,RIde9fcc8_369,RIfcd9c70_7500,
        RIfe98208_8075,RIfce4698_7621,RIfe980a0_8074,RIde93158_307,RIde8f648_289,RIde8b4a8_269,RIde87308_249,RIde82e20_228,RIfcbba18_7157,RIfc48d88_5851,
        RIfc99f80_6774,RIfc8b4a8_6607,RIe16c728_2611,RIe16a400_2586,RIe168c18_2569,RIe166620_2542,RIe163920_2510,RIee38068_5096,RIe160c20_2478,RIfc48248_5843,
        RIe15df20_2446,RIe158520_2382,RIe155820_2350,RIfcbbe50_7160,RIe152b20_2318,RIfc47e10_5840,RIe14fe20_2286,RIfca0e98_6853,RIe14d120_2254,RIe14a420_2222,
        RIe147720_2190,RIfc8be80_6614,RIfc7fb08_6475,RIfc480e0_5842,RIfc99878_6769,RIe141e88_2127,RIe13fb60_2102,RIdf3da68_2078,RIdf3b5d8_2052,RIfe97f38_8073,
        RIee30070_5005,RIee2eb58_4990,RIee2deb0_4981,RIdf36880_1997,RIdf34288_1970,RIdf320c8_1946,RIfe97dd0_8072,RIfcc3740_7246,RIfc48ab8_5849,RIfce05e8_7575,
        RIfc80210_6480,RIdf2b048_1866,RIdf29158_1844,RIdf26f98_1820,RIdf254e0_1801,RIfc8bbb0_6612,RIfc48950_5848,RIdf235f0_1779,RIfc8bd18_6613,RIdf21f70_1763,
        RIdf208f0_1747,RIdf1b8c8_1690,RIdf1a3b0_1675,RIdf181f0_1651,RIdf154f0_1619,RIdf127f0_1587,RIdf0faf0_1555,RIdf0cdf0_1523,RIdf0a0f0_1491,RIdf073f0_1459,
        RIdf046f0_1427,RIdefecf0_1363,RIdefbff0_1331,RIdef92f0_1299,RIdef65f0_1267,RIdef38f0_1235,RIdef0bf0_1203,RIdeedef0_1171,RIdeeb1f0_1139,RIfcbc120_7162,
        RIfcd9838_7497,RIfc99710_6768,RIfca1168_6855,RIdee57f0_1075,RIdee3a68_1054,RIdee18a8_1030,RIdedf850_1007,RIfc549f8_5985,RIfcb5370_7084,RIfce43c8_7619,
        RIfce0480_7574,RIdeda6c0_949,RIded8230_923,RIded6070_899,RIded3d48_874,RIded1a20_849,RIdeced20_817,RIdecc020_785,RIdec9320_753,RIdeb5820_529,
        RIde993c8_337,RIe16f428_2643,RIe15b220_2414,RIe144a20_2158,RIdf39418_2028,RIdf2da78_1896,RIdf1e2f8_1720,RIdf019f0_1395,RIdee84f0_1107,RIdedd258_980,
        RIde7f310_210,RIe19e8b8_3181,RIe19bbb8_3149,RIfe976c8_8067,RIe198eb8_3117,RIf144c80_5242,RIe1961b8_3085,RIe1934b8_3053,RIe1907b8_3021,RIe18adb8_2957,
        RIe1880b8_2925,RIfe97560_8066,RIe1853b8_2893,RIfcc3fb0_7252,RIe1826b8_2861,RIe17f9b8_2829,RIe17ccb8_2797,RIfcd3730_7428,RIf1412d8_5201,RIfcc4118_7253,
        RIfe97830_8068,RIfc4a6d8_5869,RIf13f6b8_5181,RIfc9f980_6838,RIfc9fae8_6839,RIfcc3e48_7251,RIfc89e28_6591,RIfc89cc0_6590,RIe174720_2702,RIfc4a408_5867,
        RIfce27a8_7599,RIfc530a8_5967,RIfcd5d28_7455,RIf16cf28_5699,RIe224c10_4708,RIfc53210_5968,RIe221f10_4676,RIf16b1a0_5678,RIe21f210_4644,RIe219810_4580,
        RIe216b10_4548,RIfc401d8_5755,RIe213e10_4516,RIf1699b8_5661,RIe211110_4484,RIfc81cc8_6499,RIe20e410_4452,RIe20b710_4420,RIe208a10_4388,RIfc8a0f8_6593,
        RIfcb6720_7098,RIe203448_4327,RIe201828_4307,RIfc53378_5969,RIfc8a3c8_6595,RIfcb65b8_7097,RIfc49fd0_5864,RIf160bb0_5560,RIf15ecc0_5538,RIe1fd4a8_4259,
        RIfe97b00_8070,RIfc8a530_6596,RIfe97c68_8071,RIfc8a800_6598,RIfc8a698_6597,RIfc9a7f0_6780,RIfc81890_6496,RIfcd5e90_7456,RIe1fb180_4234,RIfc49e68_5863,
        RIfc81728_6495,RIfcbb1a8_7151,RIe1f66f8_4181,RIfcd3460_7426,RIfcb62e8_7095,RIfc9a520_6778,RIe1f4268_4155,RIfc49d00_5862,RIfcd9dd8_7501,RIfcbb310_7152,
        RIe1ef0d8_4097,RIe1ec978_4069,RIe1e9c78_4037,RIe1e6f78_4005,RIe1e4278_3973,RIe1e1578_3941,RIe1de878_3909,RIe1dbb78_3877,RIe1d8e78_3845,RIe1d3478_3781,
        RIe1d0778_3749,RIe1cda78_3717,RIe1cad78_3685,RIe1c8078_3653,RIe1c5378_3621,RIe1c2678_3589,RIe1bf978_3557,RIfc49a30_5860,RIfcb6018_7093,RIe1ba3b0_3496,
        RIe1b81f0_3472,RIfce0a20_7578,RIfcbb5e0_7154,RIe1b6030_3448,RIfe97998_8069,RIfce5610_7632,RIfcc3a10_7248,RIe1b3330_3416,RIe1b19e0_3398,RIfc495f8_5857,
        RIfc81188_6491,RIe1ad228_3347,RIe1aba40_3330,RIe1a9cb8_3309,RIe1a6fb8_3277,RIe1a42b8_3245,RIe1a15b8_3213,RIe18dab8_2989,RIe179fb8_2765,RIe227910_4740,
        RIe21c510_4612,RIe205d10_4356,RIe1ffd70_4288,RIe1f9128_4211,RIe1f1c70_4128,RIe1d6178_3813,RIe1bcc78_3525,RIe1afaf0_3376,RIe172128_2675,RIdec6a58_724,
        RIdec3d58_692,RIfc723e0_6322,RIdec1058_660,RIfc59fc0_6046,RIdebe358_628,RIdebb658_596,RIdeb8958_564,RIfcb96f0_7132,RIdeb2f58_500,RIfce1c68_7591,
        RIdeb0258_468,RIfc9b498_6789,RIdead558_436,RIdea6fa0_404,RIdea06a0_372,RIfc81458_6493,RIfc83780_6518,RIfc4e620_5914,RIfcd3e38_7433,RIde937e8_309,
        RIde8f990_290,RIde8bb38_271,RIde87650_250,RIde834b0_230,RIfc42c80_5782,RIfc65960_6178,RIfc6c710_6256,RIee392b0_5109,RIe16cb60_2614,RIe16a6d0_2588,
        RIe169050_2572,RIe166a58_2545,RIe163d58_2513,RIfec3cf0_8348,RIe161058_2481,RIfcd54b8_7449,RIe15e358_2449,RIe158958_2385,RIe155c58_2353,RIfe9ba48_8115,
        RIe152f58_2321,RIfec4128_8351,RIe150258_2289,RIfcb9b28_7135,RIe14d558_2257,RIe14a858_2225,RIe147b58_2193,RIfcdb2f0_7516,RIfc553d0_5992,RIfc9a0e8_6775,
        RIfcbd908_7179,RIe1422c0_2130,RIe13ff98_2105,RIdf3dea0_2081,RIdf3ba10_2055,RIfc87128_6559,RIee304a8_5008,RIfcc51f8_7265,RIee2e2e8_4984,RIdf36cb8_2000,
        RIfec3fc0_8350,RIdf32500_1949,RIfec3e58_8349,RIee2c830_4965,RIee2ad78_4946,RIee296f8_4930,RIee284b0_4917,RIfe9b8e0_8114,RIfe9b610_8112,RIfe9b778_8113,
        RIfe9b4a8_8111,RIfcb7c38_7113,RIfc86b88_6555,RIdf238c0_1781,RIfc75ab8_6361,RIdf22240_1765,RIfeaa3b8_8253,RIdf1bb98_1692,RIdf1a680_1677,RIdf18628_1654,
        RIdf15928_1622,RIdf12c28_1590,RIdf0ff28_1558,RIdf0d228_1526,RIdf0a528_1494,RIdf07828_1462,RIdf04b28_1430,RIdeff128_1366,RIdefc428_1334,RIdef9728_1302,
        RIdef6a28_1270,RIdef3d28_1238,RIdef1028_1206,RIdeee328_1174,RIdeeb628_1142,RIee25a80_4887,RIee24c70_4877,RIfcddd20_7546,RIfccc110_7344,RIdee5c28_1078,
        RIdee3ea0_1057,RIdee1b78_1032,RIdedfc88_1010,RIfc6a6b8_6233,RIee227e0_4851,RIfc88be0_6578,RIee21868_4840,RIdedaaf8_952,RIded8668_926,RIded6340_901,
        RIded4180_877,RIded1e58_852,RIdecf158_820,RIdecc458_788,RIdec9758_756,RIdeb5c58_532,RIde99da0_340,RIe16f860_2646,RIe15b658_2417,RIe144e58_2161,
        RIdf39850_2031,RIdf2deb0_1899,RIdf1e730_1723,RIdf01e28_1398,RIdee8928_1110,RIdedd690_983,RIde7fce8_213,RIe19ecf0_3184,RIe19bff0_3152,RIf145a90_5252,
        RIe1992f0_3120,RIf144de8_5243,RIe1965f0_3088,RIe1938f0_3056,RIe190bf0_3024,RIe18b1f0_2960,RIe1884f0_2928,RIfc72980_6326,RIe1857f0_2896,RIf143060_5222,
        RIe182af0_2864,RIe17fdf0_2832,RIe17d0f0_2800,RIf142688_5215,RIf141710_5204,RIe177858_2737,RIe176778_2725,RIfcea638_7689,RIfca54e8_6903,RIee3e878_5170,
        RIee3dbd0_5161,RIee3c988_5148,RIee3b5d8_5134,RIee3a4f8_5122,RIe174b58_2705,RIf170600_5738,RIfc76fd0_6376,RIf16e9e0_5718,RIfced608_7723,RIf16d090_5700,
        RIe225048_4711,RIf16c550_5692,RIe222348_4679,RIf16b470_5680,RIe21f648_4647,RIe219c48_4583,RIe216f48_4551,RIf16a4f8_5669,RIe214248_4519,RIf169df0_5664,
        RIe211548_4487,RIf1684a0_5646,RIe20e848_4455,RIe20bb48_4423,RIe208e48_4391,RIf1673c0_5634,RIf166448_5623,RIfe9c6f0_8124,RIfe9c150_8120,RIf1654d0_5612,
        RIfcc4550_7256,RIf1635e0_5590,RIf162500_5578,RIf160fe8_5563,RIf15f0f8_5541,RIfe9bfe8_8119,RIfe9c588_8123,RIf15d208_5519,RIf15bfc0_5506,RIfc4d540_5902,
        RIfc9c848_6803,RIfec4290_8352,RIfe9c2b8_8121,RIfcc01d0_7208,RIe1fb2e8_4235,RIfe9c420_8122,RIfca3e68_6887,RIf154c70_5424,RIe1f69c8_4183,RIf153a28_5411,
        RIf152240_5394,RIf150ff8_5381,RIe1f46a0_4158,RIfca6028_6911,RIfc43bf8_5793,RIf14e460_5350,RIe1ef3a8_4099,RIe1ecdb0_4072,RIe1ea0b0_4040,RIe1e73b0_4008,
        RIe1e46b0_3976,RIe1e19b0_3944,RIe1decb0_3912,RIe1dbfb0_3880,RIe1d92b0_3848,RIe1d38b0_3784,RIe1d0bb0_3752,RIe1cdeb0_3720,RIe1cb1b0_3688,RIe1c84b0_3656,
        RIe1c57b0_3624,RIe1c2ab0_3592,RIe1bfdb0_3560,RIfc4d6a8_5903,RIf14be68_5323,RIe1ba680_3498,RIfe9be80_8118,RIfc86e58_6557,RIfcd46a8_7439,RIe1b6300_3450,
        RIfe9bd18_8117,RIf1495a0_5294,RIf1481f0_5280,RIe1b3600_3418,RIe1b1e18_3401,RIfc69470_6220,RIfcbfac8_7203,RIfe9bbb0_8116,RIe1abd10_3332,RIe1aa0f0_3312,
        RIe1a73f0_3280,RIe1a46f0_3248,RIe1a19f0_3216,RIe18def0_2992,RIe17a3f0_2768,RIe227d48_4743,RIe21c948_4615,RIe206148_4359,RIe2001a8_4291,RIe1f9560_4214,
        RIe1f20a8_4131,RIe1d65b0_3816,RIe1bd0b0_3528,RIe1aff28_3379,RIe172560_2678,RIdec68f0_723,RIdec3bf0_691,RIee208f0_4829,RIdec0ef0_659,RIfc7ce08_6443,
        RIdebe1f0_627,RIdebb4f0_595,RIdeb87f0_563,RIfc9b8d0_6792,RIdeb2df0_499,RIfcc6710_7280,RIdeb00f0_467,RIfc5ff60_6114,RIdead3f0_435,RIdea6c58_403,
        RIdea0358_371,RIfce5070_7628,RIee1c6d8_4782,RIfce70c8_7651,RIee1b058_4766,RIde934a0_308,RIfe9b1d8_8109,RIde8b7f0_270,RIfe9b340_8110,RIfc6b798_6245,
        RIfcb2238_7049,RIfcd3a00_7430,RIfcdb020_7514,RIfc511b8_5945,RIe16c9f8_2613,RIfcb27d8_7053,RIe168ee8_2571,RIe1668f0_2544,RIe163bf0_2512,RIee381d0_5097,
        RIe160ef0_2480,RIfcdfaa8_7567,RIe15e1f0_2448,RIe1587f0_2384,RIe155af0_2352,RIfc3f968_5749,RIe152df0_2320,RIfcd5080_7446,RIe1500f0_2288,RIfc84b30_6532,
        RIe14d3f0_2256,RIe14a6f0_2224,RIe1479f0_2192,RIfcea098_7685,RIfc92f00_6694,RIfc54890_5984,RIfcdcc40_7534,RIe142158_2129,RIe13fe30_2104,RIdf3dd38_2080,
        RIdf3b8a8_2054,RIfc57590_6016,RIee30340_5007,RIfcd0490_7392,RIee2e180_4983,RIdf36b50_1999,RIdf34558_1972,RIdf32398_1948,RIfe9b070_8108,RIfcb1860_7042,
        RIfca1b40_6862,RIfc5c018_6069,RIfe9ada0_8106,RIdf2b318_1868,RIdf29428_1846,RIdf27100_1821,RIfe9af08_8107,RIfc5e1d8_6093,RIfcdcda8_7535,RIfcac400_6982,
        RIfc691a0_6218,RIfcaad80_6966,RIdf20bc0_1749,RIfc61b80_6134,RIdf1a518_1676,RIdf184c0_1653,RIdf157c0_1621,RIdf12ac0_1589,RIdf0fdc0_1557,RIdf0d0c0_1525,
        RIdf0a3c0_1493,RIdf076c0_1461,RIdf049c0_1429,RIdefefc0_1365,RIdefc2c0_1333,RIdef95c0_1301,RIdef68c0_1269,RIdef3bc0_1237,RIdef0ec0_1205,RIdeee1c0_1173,
        RIdeeb4c0_1141,RIfc69b78_6225,RIfc6b900_6246,RIfc4d270_5900,RIfced770_7724,RIdee5ac0_1077,RIdee3d38_1056,RIdee1a10_1031,RIdedfb20_1009,RIfc7ff40_6478,
        RIfca4408_6891,RIfcb5640_7086,RIee21700_4839,RIdeda990_951,RIded8500_925,RIded61d8_900,RIded4018_876,RIded1cf0_851,RIdeceff0_819,RIdecc2f0_787,
        RIdec95f0_755,RIdeb5af0_531,RIde99a58_339,RIe16f6f8_2645,RIe15b4f0_2416,RIe144cf0_2160,RIdf396e8_2030,RIdf2dd48_1898,RIdf1e5c8_1722,RIdf01cc0_1397,
        RIdee87c0_1109,RIdedd528_982,RIde7f9a0_212,RIe19eb88_3183,RIe19be88_3151,RIfe9a698_8101,RIe199188_3119,RIfe9a530_8100,RIe196488_3087,RIe193788_3055,
        RIe190a88_3023,RIe18b088_2959,RIe188388_2927,RIfe9a800_8102,RIe185688_2895,RIfc8d938_6633,RIe182988_2863,RIe17fc88_2831,RIe17cf88_2799,RIfe9a3c8_8099,
        RIf1415a8_5203,RIfe9a260_8098,RIfe9a0f8_8097,RIfcb9150_7128,RIf13f820_5182,RIfc9fc50_6840,RIfce5340_7630,RIfc5cb58_6077,RIfc576f8_6017,RIfc780b0_6388,
        RIe1749f0_2704,RIfc7adb0_6420,RIfc7c2c8_6435,RIfcb2d78_7057,RIfc7e758_6461,RIfe9aad0_8104,RIe224ee0_4710,RIf16c3e8_5691,RIe2221e0_4678,RIfcd3898_7429,
        RIe21f4e0_4646,RIe219ae0_4582,RIe216de0_4550,RIfc880a0_6570,RIe2140e0_4518,RIf169c88_5663,RIe2113e0_4486,RIf168338_5645,RIe20e6e0_4454,RIe20b9e0_4422,
        RIe208ce0_4390,RIfce4c38_7625,RIfc9c6e0_6802,RIe2035b0_4328,RIe201af8_4309,RIfc500d8_5933,RIfc85c10_6544,RIfce81a8_7663,RIfce9c60_7682,RIf160e80_5562,
        RIf15ef90_5540,RIfe9a968_8103,RIfe9ac38_8105,RIfca8d28_6943,RIf15be58_5505,RIfcedba8_7727,RIfc6a988_6235,RIfc71cd8_6317,RIfccb198_7333,RIfcaa3a8_6959,
        RIfec3b88_8347,RIfc4c730_5892,RIfc6d688_6267,RIfca8e90_6944,RIe1f6860_4182,RIfc64e20_6170,RIfcaee30_7012,RIfccee10_7376,RIe1f4538_4157,RIfc63ea8_6159,
        RIfcaecc8_7011,RIfcae458_7005,RIfeab1c8_8263,RIe1ecc48_4071,RIe1e9f48_4039,RIe1e7248_4007,RIe1e4548_3975,RIe1e1848_3943,RIe1deb48_3911,RIe1dbe48_3879,
        RIe1d9148_3847,RIe1d3748_3783,RIe1d0a48_3751,RIe1cdd48_3719,RIe1cb048_3687,RIe1c8348_3655,RIe1c5648_3623,RIe1c2948_3591,RIe1bfc48_3559,RIfcc70e8_7287,
        RIfca7ae0_6930,RIe1ba518_3497,RIe1b8358_3473,RIfc598b8_6041,RIfcc2228_7231,RIe1b6198_3449,RIe1b4848_3431,RIfc82f10_6512,RIfc55970_5996,RIe1b3498_3417,
        RIe1b1cb0_3400,RIfcb7698_7109,RIfc4b4e8_5879,RIe1ad390_3348,RIe1abba8_3331,RIe1a9f88_3311,RIe1a7288_3279,RIe1a4588_3247,RIe1a1888_3215,RIe18dd88_2991,
        RIe17a288_2767,RIe227be0_4742,RIe21c7e0_4614,RIe205fe0_4358,RIe200040_4290,RIe1f93f8_4213,RIe1f1f40_4130,RIe1d6448_3815,RIe1bcf48_3527,RIe1afdc0_3378,
        RIe1723f8_2677,RIdec6d28_726,RIdec4028_694,RIee20bc0_4831,RIdec1328_662,RIfcbaed8_7149,RIdebe628_630,RIdebb928_598,RIdeb8c28_566,RIfc412b8_5767,
        RIdeb3228_502,RIfc9ea08_6827,RIdeb0528_470,RIee1e028_4800,RIdead828_438,RIdea7630_406,RIdea0d30_374,RIfcbac08_7147,RIfc55538_5993,RIfcba668_7143,
        RIfc4af48_5875,RIfe912f0_7996,RIfe91458_7997,RIde8be80_272,RIde87ce0_252,RIfc85238_6537,RIfc88640_6574,RIfcda210_7504,RIfcd5788_7451,RIee39418_5110,
        RIe16ce30_2616,RIfc884d8_6573,RIe169320_2574,RIe166d28_2547,RIe164028_2515,RIfe90918_7989,RIe161328_2483,RIee36880_5079,RIe15e628_2451,RIe158c28_2387,
        RIe155f28_2355,RIfe91188_7995,RIe153228_2323,RIfe91020_7994,RIe150528_2291,RIfcda378_7505,RIe14d828_2259,RIe14ab28_2227,RIe147e28_2195,RIfe90eb8_7993,
        RIfe90d50_7992,RIfcb99c0_7134,RIfc9c2a8_6799,RIfe90be8_7991,RIfe90a80_7990,RIdf3e008_2082,RIdf3bce0_2057,RIfcec690_7712,RIee30778_5010,RIfc87dd0_6568,
        RIee2e5b8_4986,RIdf36e20_2001,RIdf346c0_1973,RIdf32668_1950,RIdf30070_1923,RIee2c998_4966,RIee2aee0_4947,RIee299c8_4932,RIee28618_4918,RIfe90378_7985,
        RIfe907b0_7988,RIfe904e0_7986,RIfe90648_7987,RIfc9d928_6815,RIfc86048_6547,RIfcb92b8_7129,RIfc4ee90_5920,RIfc86a20_6554,RIdf20e90_1751,RIfcb8fe8_7127,
        RIdf1a950_1679,RIdf188f8_1656,RIdf15bf8_1624,RIdf12ef8_1592,RIdf101f8_1560,RIdf0d4f8_1528,RIdf0a7f8_1496,RIdf07af8_1464,RIdf04df8_1432,RIdeff3f8_1368,
        RIdefc6f8_1336,RIdef99f8_1304,RIdef6cf8_1272,RIdef3ff8_1240,RIdef12f8_1208,RIdeee5f8_1176,RIdeeb8f8_1144,RIfc857d8_6541,RIee24dd8_4878,RIfc4ff70_5932,
        RIfc50240_5934,RIdee5ef8_1080,RIdee4170_1059,RIfe915c0_7998,RIdedff58_1012,RIfcd4810_7440,RIee22948_4852,RIfce1560_7586,RIee219d0_4841,RIdedac60_953,
        RIfe91728_7999,RIded64a8_902,RIfe91890_8000,RIded2128_854,RIdecf428_822,RIdecc728_790,RIdec9a28_758,RIdeb5f28_534,RIde9a430_342,RIe16fb30_2648,
        RIe15b928_2419,RIe145128_2163,RIdf39b20_2033,RIdf2e180_1901,RIdf1ea00_1725,RIdf020f8_1400,RIdee8bf8_1112,RIdedd960_985,RIde80378_215,RIe19efc0_3186,
        RIe19c2c0_3154,RIf145d60_5254,RIe1995c0_3122,RIfc637a0_6154,RIe1968c0_3090,RIe193bc0_3058,RIe190ec0_3026,RIe18b4c0_2962,RIe1887c0_2930,RIfc62af8_6145,
        RIe185ac0_2898,RIfe8fc70_7980,RIe182dc0_2866,RIe1800c0_2834,RIe17d3c0_2802,RIfe90210_7984,RIfe8ff40_7982,RIfc72f20_6330,RIe176a48_2727,RIfcaf6a0_7018,
        RIfc61040_6126,RIf13e8a8_5171,RIfe900a8_7983,RIee3caf0_5149,RIee3b740_5135,RIee3a660_5123,RIe174e28_2707,RIf170768_5739,RIfc5fdf8_6113,RIf16eb48_5719,
        RIfcaaab0_6964,RIf16d1f8_5701,RIe225318_4713,RIf16c6b8_5693,RIe222618_4681,RIf16b5d8_5681,RIe21f918_4649,RIe219f18_4585,RIe217218_4553,RIfca62f8_6913,
        RIe214518_4521,RIfcc9578_7313,RIe211818_4489,RIfca5a88_6907,RIe20eb18_4457,RIe20be18_4425,RIe209118_4393,RIf167690_5636,RIf166718_5625,RIfe8f9a0_7978,
        RIfe8f838_7977,RIf165638_5613,RIf164990_5604,RIf1638b0_5592,RIf1627d0_5580,RIf161150_5564,RIf15f260_5542,RIe1fd778_4261,RIe1fc530_4248,RIf15d4d8_5521,
        RIf15c290_5508,RIfca20e0_6866,RIf159f68_5483,RIf159428_5475,RIf1581e0_5462,RIfc5ebb0_6100,RIfe8fdd8_7981,RIfc69e48_6227,RIfc5e8e0_6098,RIf154f40_5426,
        RIe1f6b30_4184,RIf153b90_5412,RIf1523a8_5395,RIfce88b0_7668,RIfe8fb08_7979,RIfcebe20_7706,RIfcb1158_7037,RIf14e730_5352,RIe1ef678_4101,RIe1ed080_4074,
        RIe1ea380_4042,RIe1e7680_4010,RIe1e4980_3978,RIe1e1c80_3946,RIe1def80_3914,RIe1dc280_3882,RIe1d9580_3850,RIe1d3b80_3786,RIe1d0e80_3754,RIe1ce180_3722,
        RIe1cb480_3690,RIe1c8780_3658,RIe1c5a80_3626,RIe1c2d80_3594,RIe1c0080_3562,RIfcc8ba0_7306,RIfc5d698_6085,RIfec35e8_8343,RIfeabd08_8271,RIfc5cf90_6080,
        RIfc5ce28_6079,RIfec31b0_8340,RIe1b4b18_3433,RIf149708_5295,RIf148358_5281,RIe1b3768_3419,RIfec3480_8342,RIfc483b0_5844,RIfc80be8_6487,RIe1ad4f8_3349,
        RIfec3318_8341,RIe1aa3c0_3314,RIe1a76c0_3282,RIe1a49c0_3250,RIe1a1cc0_3218,RIe18e1c0_2994,RIe17a6c0_2770,RIe228018_4745,RIe21cc18_4617,RIe206418_4361,
        RIe200478_4293,RIe1f9830_4216,RIe1f2378_4133,RIe1d6880_3818,RIe1bd380_3530,RIe1b01f8_3381,RIe172830_2680,RIdec6bc0_725,RIdec3ec0_693,RIee20a58_4830,
        RIdec11c0_661,RIee1f978_4818,RIdebe4c0_629,RIdebb7c0_597,RIdeb8ac0_565,RIee1efa0_4811,RIdeb30c0_501,RIfcb04b0_7028,RIdeb03c0_469,RIfc5e4a8_6095,
        RIdead6c0_437,RIdea72e8_405,RIdea09e8_373,RIfcb2508_7051,RIfcd16d8_7405,RIfc5d800_6086,RIfc63d40_6158,RIde93b30_310,RIfea7820_8222,RIfea73e8_8219,
        RIde87998_251,RIde837f8_231,RIfc7bd28_6431,RIfcc7ef8_7297,RIfc7a108_6411,RIfc7a6a8_6415,RIe16ccc8_2615,RIe16a838_2589,RIe1691b8_2573,RIe166bc0_2546,
        RIe163ec0_2514,RIee38338_5098,RIe1611c0_2482,RIfc54b60_5986,RIe15e4c0_2450,RIe158ac0_2386,RIe155dc0_2354,RIee35a70_5069,RIe1530c0_2322,RIee357a0_5067,
        RIe1503c0_2290,RIfc9fdb8_6841,RIe14d6c0_2258,RIe14a9c0_2226,RIe147cc0_2194,RIee34af8_5058,RIee33a18_5046,RIee327d0_5033,RIfcbcf30_7172,RIe142428_2131,
        RIe140100_2106,RIfea7280_8218,RIdf3bb78_2056,RIfc731f0_6332,RIee30610_5009,RIfcbe010_7184,RIee2e450_4985,RIfec2ee0_8338,RIfec3048_8339,RIfec2c10_8336,
        RIfec2d78_8337,RIfcb46c8_7075,RIfcb4830_7076,RIee29860_4931,RIfcb88e0_7122,RIdf2b480_1869,RIdf29590_1847,RIdf27268_1822,RIdf25648_1802,RIfcc9de8_7319,
        RIfc53648_5971,RIdf23a28_1782,RIfc823d0_6504,RIdf223a8_1766,RIdf20d28_1750,RIdf1bd00_1693,RIdf1a7e8_1678,RIdf18790_1655,RIdf15a90_1623,RIdf12d90_1591,
        RIdf10090_1559,RIdf0d390_1527,RIdf0a690_1495,RIdf07990_1463,RIdf04c90_1431,RIdeff290_1367,RIdefc590_1335,RIdef9890_1303,RIdef6b90_1271,RIdef3e90_1239,
        RIdef1190_1207,RIdeee490_1175,RIdeeb790_1143,RIee25be8_4888,RIfc6af28_6239,RIee23fc8_4868,RIfccf680_7382,RIdee5d90_1079,RIdee4008_1058,RIdee1ce0_1033,
        RIdedfdf0_1011,RIfc6b090_6240,RIfc534e0_5970,RIfca5920_6906,RIfc66770_6188,RIfe8f6d0_7976,RIded87d0_927,RIfe8f568_7975,RIded42e8_878,RIded1fc0_853,
        RIdecf2c0_821,RIdecc5c0_789,RIdec98c0_757,RIdeb5dc0_533,RIde9a0e8_341,RIe16f9c8_2647,RIe15b7c0_2418,RIe144fc0_2162,RIdf399b8_2032,RIdf2e018_1900,
        RIdf1e898_1724,RIdf01f90_1399,RIdee8a90_1111,RIdedd7f8_984,RIde80030_214,RIe19ee58_3185,RIe19c158_3153,RIf145bf8_5253,RIe199458_3121,RIfe8f298_7973,
        RIe196758_3089,RIe193a58_3057,RIe190d58_3025,RIe18b358_2961,RIe188658_2929,RIfe8f130_7972,RIe185958_2897,RIfc9f278_6833,RIe182c58_2865,RIe17ff58_2833,
        RIe17d258_2801,RIf1427f0_5216,RIfe8efc8_7971,RIe1779c0_2738,RIe1768e0_2726,RIfc81e30_6500,RIfc9ff20_6842,RIfca0088_6843,RIfc81b60_6498,RIfce5778_7633,
        RIfce08b8_7577,RIfc815c0_6494,RIe174cc0_2706,RIfca04c0_6846,RIfc53eb8_5977,RIfcc65a8_7279,RIfc80d50_6488,RIfc804e0_6482,RIe2251b0_4712,RIfc80378_6481,
        RIe2224b0_4680,RIfcb5910_7088,RIe21f7b0_4648,RIe219db0_4584,RIe2170b0_4552,RIfca01f0_6844,RIe2143b0_4520,RIfc82c40_6510,RIe2116b0_4488,RIfc7f6d0_6472,
        RIe20e9b0_4456,RIe20bcb0_4424,RIe208fb0_4392,RIf167528_5635,RIf1665b0_5624,RIe203718_4329,RIe201c60_4310,RIfc9da90_6816,RIfcc5360_7266,RIf163748_5591,
        RIf162668_5579,RIfc7e320_6458,RIfc87998_6565,RIe1fd610_4260,RIe1fc3c8_4247,RIf15d370_5520,RIf15c128_5507,RIfcc5d38_7273,RIfce7d70_7660,RIfc4bd58_5885,
        RIfc55c40_5998,RIfca2ab8_6873,RIe1fb450_4236,RIf156890_5444,RIfcd5ff8_7457,RIf154dd8_5425,RIfec2aa8_8335,RIfcb4b00_7078,RIfcd9400_7494,RIf151160_5382,
        RIe1f4808_4159,RIfc44738_5801,RIfc90908_6667,RIf14e5c8_5351,RIe1ef510_4100,RIe1ecf18_4073,RIe1ea218_4041,RIe1e7518_4009,RIe1e4818_3977,RIe1e1b18_3945,
        RIe1dee18_3913,RIe1dc118_3881,RIe1d9418_3849,RIe1d3a18_3785,RIe1d0d18_3753,RIe1ce018_3721,RIe1cb318_3689,RIe1c8618_3657,RIe1c5918_3625,RIe1c2c18_3593,
        RIe1bff18_3561,RIf14d218_5337,RIfe8ee60_7970,RIfea8090_8228,RIe1b84c0_3474,RIf14aab8_5309,RIfc6c170_6252,RIe1b6468_3451,RIe1b49b0_3432,RIfcafad8_7021,
        RIfcaa948_6963,RIfe8ecf8_7969,RIfe8f400_7974,RIfc67f58_6205,RIfca8ff8_6945,RIfe8eb90_7968,RIe1abe78_3333,RIe1aa258_3313,RIe1a7558_3281,RIe1a4858_3249,
        RIe1a1b58_3217,RIe18e058_2993,RIe17a558_2769,RIe227eb0_4744,RIe21cab0_4616,RIe2062b0_4360,RIe200310_4292,RIe1f96c8_4215,RIe1f2210_4132,RIe1d6718_3817,
        RIe1bd218_3529,RIe1b0090_3380,RIe1726c8_2679,RIdec4460_697,RIdec1760_665,RIee1fae0_4819,RIdebea60_633,RIee1f108_4812,RIdebbd60_601,RIdeb9060_569,
        RIdeb6360_537,RIee1eb68_4808,RIdeb0960_473,RIee1e460_4803,RIdeadc60_441,RIee1d7b8_4794,RIdea8008_409,RIdea1708_377,RIde9ae08_345,RIfe957d8_8045,
        RIfe95508_8043,RIfe95670_8044,RIee1a7e8_4760,RIfe95aa8_8047,RIfe95238_8041,RIfe95940_8046,RIfe953a0_8042,RIee1a0e0_4755,RIee19ca8_4752,RIee19870_4749,
        RIee19438_4746,RIee38ba8_5104,RIfe95c10_8048,RIee384a0_5099,RIfea9440_8242,RIe164460_2518,RIe161760_2486,RIfe942c0_8030,RIe15ea60_2454,RIfe94158_8029,
        RIe15bd60_2422,RIe156360_2358,RIe153660_2326,RIfe94428_8031,RIe150960_2294,RIfe94590_8032,RIe14dc60_2262,RIfc5c2e8_6071,RIe14af60_2230,RIe148260_2198,
        RIe145560_2166,RIee33ce8_5048,RIee32aa0_5035,RIee31858_5022,RIfc5d530_6084,RIe140538_2109,RIdf3e2d8_2084,RIdf3c118_2060,RIdf39df0_2035,RIfcdd780_7542,
        RIee2ee28_4992,RIfcc88d0_7304,RIee2cc68_4968,RIdf34990_1975,RIdf32aa0_1953,RIdf304a8_1926,RIdf2e5b8_1904,RIee2b1b0_4949,RIfe946f8_8033,RIfcb2940_7054,
        RIee273d0_4905,RIfe949c8_8035,RIdf27538_1824,RIfe94b30_8036,RIfe94860_8034,RIee26f98_4902,RIee269f8_4898,RIee26728_4896,RIee26458_4894,RIee26188_4892,
        RIfe94c98_8037,RIee25d50_4889,RIfea9170_8240,RIdf16030_1627,RIdf13330_1595,RIdf10630_1563,RIdf0d930_1531,RIdf0ac30_1499,RIdf07f30_1467,RIdf05230_1435,
        RIdf02530_1403,RIdefcb30_1339,RIdef9e30_1307,RIdef7130_1275,RIdef4430_1243,RIdef1730_1211,RIdeeea30_1179,RIdeebd30_1147,RIdee9030_1115,RIee250a8_4880,
        RIee24298_4870,RIee23758_4862,RIee22d80_4855,RIfe950d0_8040,RIfe94f68_8039,RIfe94e00_8038,RIdeddd98_988,RIee22ab0_4853,RIee21e08_4844,RIfca46d8_6893,
        RIfc5dad0_6088,RIfeaa250_8252,RIfe96048_8051,RIfe95d78_8049,RIfe95ee0_8050,RIdecf860_825,RIdeccb60_793,RIdec9e60_761,RIdec7160_729,RIdeb3660_505,
        RIde94508_313,RIe16d268_2619,RIe159060_2390,RIe142860_2134,RIdf37258_2004,RIdf2b8b8_1872,RIdf1c138_1696,RIdeff830_1371,RIdee6330_1083,RIdedb098_956,
        RIde7a450_186,RIe19c6f8_3157,RIe1999f8_3125,RIf1450b8_5245,RIe196cf8_3093,RIf143fd8_5233,RIe193ff8_3061,RIe1912f8_3029,RIe18e5f8_2997,RIe188bf8_2933,
        RIe185ef8_2901,RIfe973f8_8065,RIe1831f8_2869,RIf142958_5217,RIe1804f8_2837,RIe17d7f8_2805,RIe17aaf8_2773,RIf141b48_5207,RIfc542f0_5980,RIfc800a8_6479,
        RIe175260_2710,RIfca0bc8_6851,RIfc48680_5846,RIee3dea0_5163,RIfcc6878_7281,RIee3ba10_5137,RIee3a930_5125,RIfe97290_8064,RIe172b00_2682,RIf16f958_5729,
        RIf16ee18_5721,RIf16da68_5707,RIf16d360_5702,RIfe96e58_8061,RIe222a50_4684,RIfe96cf0_8060,RIe21fd50_4652,RIf16a660_5670,RIe21d050_4620,RIe217650_4556,
        RIe214950_4524,RIf169f58_5665,RIe211c50_4492,RIf168770_5648,RIe20ef50_4460,RIf1677f8_5637,RIe20c250_4428,RIe209550_4396,RIe206850_4364,RIf166880_5626,
        RIf1657a0_5614,RIe201dc8_4311,RIe2005e0_4294,RIfe96b88_8059,RIf163b80_5594,RIf162c08_5583,RIf161420_5566,RIf15f530_5544,RIf15d7a8_5523,RIfe968b8_8057,
        RIfe96a20_8058,RIfcb3fc0_7070,RIfc7cf70_6444,RIfc579c8_6019,RIf159590_5476,RIf1584b0_5464,RIf157268_5451,RIf1569f8_5445,RIfe965e8_8055,RIf155d50_5436,
        RIf155210_5428,RIf153e60_5414,RIfe96750_8056,RIf1527e0_5398,RIf151430_5384,RIfcd2650_7416,RIe1f2648_4135,RIf14f108_5359,RIfc7f298_6469,RIf14d4e8_5339,
        RIe1ed350_4076,RIe1ea7b8_4045,RIe1e7ab8_4013,RIe1e4db8_3981,RIe1e20b8_3949,RIe1df3b8_3917,RIe1dc6b8_3885,RIe1d99b8_3853,RIe1d6cb8_3821,RIe1d12b8_3757,
        RIe1ce5b8_3725,RIe1cb8b8_3693,RIe1c8bb8_3661,RIe1c5eb8_3629,RIe1c31b8_3597,RIe1c04b8_3565,RIe1bd7b8_3533,RIf14c138_5325,RIf14ad88_5311,RIe1b8790_3476,
        RIfe96480_8054,RIf14a0e0_5302,RIf149870_5296,RIfe97128_8063,RIfe96318_8053,RIf148628_5283,RIfc58d78_6033,RIe1b20e8_3403,RIe1b04c8_3383,RIf146cd8_5265,
        RIfc591b0_6036,RIfe961b0_8052,RIfe96fc0_8062,RIe1a7af8_3285,RIe1a4df8_3253,RIe1a20f8_3221,RIe19f3f8_3189,RIe18b8f8_2965,RIe177df8_2741,RIe225750_4716,
        RIe21a350_4588,RIe203b50_4332,RIe1fdbb0_4264,RIe1f6f68_4187,RIe1efab0_4104,RIe1d3fb8_3789,RIe1baab8_3501,RIe1ad930_3352,RIe16ff68_2651,RIdec42f8_696,
        RIdec15f8_664,RIfcc6cb0_7284,RIdebe8f8_632,RIfe93780_8022,RIdebbbf8_600,RIdeb8ef8_568,RIdeb61f8_536,RIee1ea00_4807,RIdeb07f8_472,RIee1e2f8_4802,
        RIdeadaf8_440,RIfc5d3c8_6083,RIdea7cc0_408,RIdea13c0_376,RIde9aac0_344,RIfc58238_6025,RIfcc3b78_7249,RIfc7d0d8_6445,RIfc59750_6040,RIfe93a50_8024,
        RIfe938e8_8023,RIde88370_254,RIde83e88_233,RIfc5f420_6106,RIfc976b8_6745,RIfc90a70_6668,RIfc60500_6118,RIee38a40_5103,RIe16ab08_2591,RIe169488_2575,
        RIe166ff8_2549,RIe1642f8_2517,RIe1615f8_2485,RIee369e8_5080,RIe15e8f8_2453,RIee35bd8_5070,RIe15bbf8_2421,RIe1561f8_2357,RIe1534f8_2325,RIfc3ee28_5741,
        RIe1507f8_2293,RIfce6c90_7648,RIe14daf8_2261,RIfcca7c0_7326,RIe14adf8_2229,RIe1480f8_2197,RIe1453f8_2165,RIee33b80_5047,RIee32938_5034,RIee316f0_5021,
        RIee30bb0_5013,RIe1403d0_2108,RIfe93618_8021,RIdf3bfb0_2059,RIfe934b0_8020,RIfcd0d00_7398,RIee2ecc0_4991,RIee2e720_4987,RIee2cb00_4967,RIfe93bb8_8025,
        RIdf32938_1952,RIdf30340_1925,RIdf2e450_1903,RIee2b048_4948,RIee29b30_4933,RIfc67148_6195,RIfc6fb18_6293,RIdf29860_1849,RIfe931e0_8018,RIfe93348_8019,
        RIfe93078_8017,RIfc672b0_6196,RIfca8788_6939,RIdf22510_1767,RIfcea7a0_7690,RIdf20ff8_1752,RIdf1ecd0_1727,RIdf1aab8_1680,RIfea7c58_8225,RIdf15ec8_1626,
        RIdf131c8_1594,RIdf104c8_1562,RIdf0d7c8_1530,RIdf0aac8_1498,RIdf07dc8_1466,RIdf050c8_1434,RIdf023c8_1402,RIdefc9c8_1338,RIdef9cc8_1306,RIdef6fc8_1274,
        RIdef42c8_1242,RIdef15c8_1210,RIdeee8c8_1178,RIdeebbc8_1146,RIdee8ec8_1114,RIee24f40_4879,RIee24130_4869,RIee235f0_4861,RIee22c18_4854,RIfe93d20_8026,
        RIdee1fb0_1035,RIdee0228_1014,RIdeddc30_987,RIfc684f8_6209,RIee21ca0_4843,RIfc68390_6208,RIee20d28_4832,RIded8aa0_929,RIfe93ff0_8028,RIded45b8_880,
        RIfe93e88_8027,RIdecf6f8_824,RIdecc9f8_792,RIdec9cf8_760,RIdec6ff8_728,RIdeb34f8_504,RIde941c0_312,RIe16d100_2618,RIe158ef8_2389,RIe1426f8_2133,
        RIdf370f0_2003,RIdf2b750_1871,RIdf1bfd0_1695,RIdeff6c8_1370,RIdee61c8_1082,RIdedaf30_955,RIde7a108_185,RIe19c590_3156,RIe199890_3124,RIf144f50_5244,
        RIe196b90_3092,RIfc76058_6365,RIe193e90_3060,RIe191190_3028,RIe18e490_2996,RIe188a90_2932,RIe185d90_2900,RIfccd8f8_7361,RIe183090_2868,RIfc76e68_6375,
        RIe180390_2836,RIe17d690_2804,RIe17a990_2772,RIf1419e0_5206,RIf140630_5192,RIe176bb0_2728,RIe1750f8_2709,RIfcd1840_7406,RIfc5f6f0_6108,RIee3dd38_5162,
        RIee3cc58_5150,RIee3b8a8_5136,RIee3a7c8_5124,RIee39580_5111,RIfea9008_8239,RIf16f7f0_5728,RIf16ecb0_5720,RIf16d900_5706,RIfc78ec0_6398,RIfcc8060_7298,
        RIe2228e8_4683,RIfc5a3f8_6049,RIe21fbe8_4651,RIfc74000_6342,RIe21cee8_4619,RIe2174e8_4555,RIe2147e8_4523,RIfca2c20_6874,RIe211ae8_4491,RIfca2950_6872,
        RIe20ede8_4459,RIfcc24f8_7233,RIe20c0e8_4427,RIe2093e8_4395,RIe2066e8_4363,RIfc45110_5808,RIfcc6f80_7286,RIfe92f10_8016,RIfe92970_8012,RIf164af8_5605,
        RIf163a18_5593,RIf162aa0_5582,RIfe92ad8_8013,RIf15f3c8_5543,RIf15d640_5522,RIfe92808_8011,RIfe92c40_8014,RIfe926a0_8010,RIfe92da8_8015,RIfe92538_8009,
        RIfcb5a78_7089,RIf158348_5463,RIf157100_5450,RIfc53be8_5975,RIfec38b8_8345,RIfcc5ea0_7274,RIf1550a8_5427,RIf153cf8_5413,RIfec3a20_8346,RIf152678_5397,
        RIfec3750_8344,RIf14ff18_5369,RIfe923d0_8008,RIf14efa0_5358,RIf14e898_5353,RIf14d380_5338,RIfe92268_8007,RIe1ea650_4044,RIe1e7950_4012,RIe1e4c50_3980,
        RIe1e1f50_3948,RIe1df250_3916,RIe1dc550_3884,RIe1d9850_3852,RIe1d6b50_3820,RIe1d1150_3756,RIe1ce450_3724,RIe1cb750_3692,RIe1c8a50_3660,RIe1c5d50_3628,
        RIe1c3050_3596,RIe1c0350_3564,RIe1bd650_3532,RIfcda4e0_7506,RIfc9d220_6810,RIe1b8628_3475,RIe1b6738_3453,RIfc4f2c8_5923,RIfce16c8_7587,RIfe91cc8_8003,
        RIfe91e30_8004,RIf1484c0_5282,RIf147548_5271,RIfe91f98_8005,RIfe91b60_8002,RIf146b70_5264,RIfc9f548_6835,RIfe92100_8006,RIfe919f8_8001,RIe1a7990_3284,
        RIe1a4c90_3252,RIe1a1f90_3220,RIe19f290_3188,RIe18b790_2964,RIe177c90_2740,RIe2255e8_4715,RIe21a1e8_4587,RIe2039e8_4331,RIe1fda48_4263,RIe1f6e00_4186,
        RIe1ef948_4103,RIe1d3e50_3788,RIe1ba950_3500,RIe1ad7c8_3351,RIe16fe00_2650,RIdec4730_699,RIdec1a30_667,RIfce3f90_7616,RIdebed30_635,RIfcc3308_7243,
        RIdebc030_603,RIdeb9330_571,RIdeb6630_539,RIfc8c588_6619,RIdeb0c30_475,RIfc5a998_6053,RIdeadf30_443,RIfc99b48_6771,RIdea8698_411,RIdea1d98_379,
        RIde9b498_347,RIfc78bf0_6396,RIfcbc558_7165,RIfca12d0_6856,RIfca3fd0_6888,RIfec2670_8332,RIfec2508_8331,RIde88a00_256,RIde84518_235,RIfcc35d8_7245,
        RIfcb57a8_7087,RIfc5a290_6048,RIfca3058_6877,RIee38e78_5106,RIfec27d8_8333,RIfca3328_6879,RIe1672c8_2551,RIe164730_2520,RIe161a30_2488,RIee36cb8_5082,
        RIe15ed30_2456,RIfcc7250_7288,RIe15c030_2424,RIe156630_2360,RIe153930_2328,RIfcc7688_7291,RIe150c30_2296,RIfc8af08_6603,RIe14df30_2264,RIfc9a250_6776,
        RIe14b230_2232,RIe148530_2200,RIe145830_2168,RIfc9aac0_6782,RIfc56bb8_6009,RIfca1ca8_6863,RIfcec960_7714,RIe1406a0_2110,RIdf3e440_2085,RIdf3c280_2061,
        RIdf39f58_2036,RIfc9a958_6781,RIee2f0f8_4994,RIfcdb458_7517,RIee2cf38_4970,RIdf34c60_1977,RIfec2940_8334,RIdf30778_1928,RIdf2e888_1906,RIee2b480_4951,
        RIfec23a0_8330,RIee288e8_4920,RIfec2238_8329,RIdf29b30_1851,RIdf27808_1826,RIdf25a80_1805,RIdf23e60_1785,RIfc55100_5990,RIfcd9f40_7502,RIfc54f98_5989,
        RIfc54cc8_5987,RIfc4b218_5877,RIdf1efa0_1729,RIfcc69e0_7282,RIdf18bc8_1658,RIdf16300_1629,RIdf13600_1597,RIdf10900_1565,RIdf0dc00_1533,RIdf0af00_1501,
        RIdf08200_1469,RIdf05500_1437,RIdf02800_1405,RIdefce00_1341,RIdefa100_1309,RIdef7400_1277,RIdef4700_1245,RIdef1a00_1213,RIdeeed00_1181,RIdeec000_1149,
        RIdee9300_1117,RIfce4ad0_7624,RIfc9e8a0_6826,RIfcc46b8_7257,RIfcd4108_7435,RIdee4440_1061,RIdee2280_1037,RIdee0390_1015,RIdede068_990,RIfcda0a8_7503,
        RIfce54a8_7631,RIfca0790_6848,RIfc50ee8_5943,RIded8d70_931,RIded68e0_905,RIded4888_882,RIded2560_857,RIdecfb30_827,RIdecce30_795,RIdeca130_763,
        RIdec7430_731,RIdeb3930_507,RIde94b98_315,RIe16d538_2621,RIe159330_2392,RIe142b30_2136,RIdf37528_2006,RIdf2bb88_1874,RIdf1c408_1698,RIdeffb00_1373,
        RIdee6600_1085,RIdedb368_958,RIde7aae0_188,RIe19c9c8_3159,RIe199cc8_3127,RIfe8ea28_7967,RIe196fc8_3095,RIfec20d0_8328,RIe1942c8_3063,RIe1915c8_3031,
        RIe18e8c8_2999,RIe188ec8_2935,RIe1861c8_2903,RIfc68228_6207,RIe1834c8_2871,RIfccb5d0_7336,RIe1807c8_2839,RIe17dac8_2807,RIe17adc8_2775,RIf141e18_5209,
        RIf140900_5194,RIf140090_5188,RIe1753c8_2711,RIf13f988_5183,RIf13ece0_5174,RIee3e170_5165,RIee3cf28_5152,RIee3bce0_5139,RIee3ac00_5127,RIee39850_5113,
        RIe172dd0_2684,RIf16fc28_5731,RIf16f0e8_5723,RIf16dd38_5709,RIfce9120_7674,RIfc404a8_5757,RIe222d20_4686,RIf16b8a8_5683,RIe220020_4654,RIf16a930_5672,
        RIe21d320_4622,RIe217920_4558,RIe214c20_4526,RIfc5b910_6064,RIe211f20_4494,RIfe8e8c0_7966,RIe20f220_4462,RIfe8e758_7965,RIe20c520_4430,RIe209820_4398,
        RIe206b20_4366,RIf166b50_5628,RIf165a70_5616,RIfe8dd80_7958,RIfe8dab0_7956,RIf164c60_5606,RIf163e50_5596,RIf162ed8_5585,RIf1616f0_5568,RIf15f800_5546,
        RIf15da78_5525,RIfe8d948_7955,RIfe8dc18_7957,RIf15c560_5510,RIf15b048_5495,RIfc62828_6143,RIf159860_5478,RIf158780_5466,RIf157538_5453,RIfca6e38_6921,
        RIe1f9b00_4218,RIfc61e50_6136,RIfc61748_6131,RIf154130_5416,RIe1f4ad8_4161,RIf152ab0_5400,RIf151700_5386,RIf1501e8_5371,RIe1f27b0_4136,RIfc60ed8_6125,
        RIfc7b620_6426,RIf14d7b8_5341,RIe1ed4b8_4077,RIe1eaa88_4047,RIe1e7d88_4015,RIe1e5088_3983,RIe1e2388_3951,RIe1df688_3919,RIe1dc988_3887,RIe1d9c88_3855,
        RIe1d6f88_3823,RIe1d1588_3759,RIe1ce888_3727,RIe1cbb88_3695,RIe1c8e88_3663,RIe1c6188_3631,RIe1c3488_3599,RIe1c0788_3567,RIe1bda88_3535,RIfca4de0_6898,
        RIfc5ea48_6099,RIe1b8a60_3478,RIe1b6a08_3455,RIfcbd638_7177,RIfc44fa8_5807,RIfe8e5f0_7964,RIfe8e1b8_7961,RIf1488f8_5285,RIf147818_5273,RIfe8e050_7960,
        RIfe8e488_7963,RIf146e40_5266,RIf146030_5256,RIfe8dee8_7959,RIfe8e320_7962,RIe1a7dc8_3287,RIe1a50c8_3255,RIe1a23c8_3223,RIe19f6c8_3191,RIe18bbc8_2967,
        RIe1780c8_2743,RIe225a20_4718,RIe21a620_4590,RIe203e20_4334,RIe1fde80_4266,RIe1f7238_4189,RIe1efd80_4106,RIe1d4288_3791,RIe1bad88_3503,RIe1adc00_3354,
        RIe170238_2653,RIdec45c8_698,RIdec18c8_666,RIfce85e0_7666,RIdebebc8_634,RIfcb8bb0_7124,RIdebbec8_602,RIdeb91c8_570,RIdeb64c8_538,RIfc85d78_6545,
        RIdeb0ac8_474,RIfc85aa8_6543,RIdeaddc8_442,RIfc4d3d8_5901,RIdea8350_410,RIdea1a50_378,RIde9b150_346,RIfc85ee0_6546,RIfc9c9b0_6804,RIfce13f8_7585,
        RIfcb8778_7121,RIfe8d510_7952,RIfe8d3a8_7951,RIde886b8_255,RIde841d0_234,RIde806c0_216,RIfcb8070_7116,RIfce1128_7583,RIfc9c140_6798,RIee38d10_5105,
        RIe16ac70_2592,RIfc850d0_6536,RIe167160_2550,RIe1645c8_2519,RIe1618c8_2487,RIee36b50_5081,RIe15ebc8_2455,RIee35d40_5071,RIe15bec8_2423,RIe1564c8_2359,
        RIe1537c8_2327,RIfc3ef90_5742,RIe150ac8_2295,RIfe8d7e0_7954,RIe14ddc8_2263,RIfce0fc0_7582,RIe14b0c8_2231,RIe1483c8_2199,RIe1456c8_2167,RIee33e50_5049,
        RIee32c08_5036,RIee319c0_5023,RIee30d18_5014,RIfe8cf70_7948,RIfe8ce08_7947,RIfe8d240_7950,RIfe8d0d8_7949,RIfce9dc8_7683,RIee2ef90_4993,RIfce51d8_7629,
        RIee2cdd0_4969,RIdf34af8_1976,RIfe8d678_7953,RIdf30610_1927,RIdf2e720_1905,RIee2b318_4950,RIee29c98_4934,RIee28780_4919,RIee27538_4906,RIdf299c8_1850,
        RIdf276a0_1825,RIdf25918_1804,RIdf23cf8_1784,RIfc83ff0_6524,RIfcb73c8_7107,RIfc51320_5946,RIfcdaa80_7510,RIfc83d20_6522,RIdf1ee38_1728,RIfc51b90_5952,
        RIdf18a60_1657,RIdf16198_1628,RIdf13498_1596,RIdf10798_1564,RIdf0da98_1532,RIdf0ad98_1500,RIdf08098_1468,RIdf05398_1436,RIdf02698_1404,RIdefcc98_1340,
        RIdef9f98_1308,RIdef7298_1276,RIdef4598_1244,RIdef1898_1212,RIdeeeb98_1180,RIdeebe98_1148,RIdee9198_1116,RIee25210_4881,RIee24400_4871,RIee238c0_4863,
        RIee22ee8_4856,RIfe8cca0_7946,RIdee2118_1036,RIfe8cb38_7945,RIdeddf00_989,RIfcc5a68_7271,RIee21f70_4845,RIfcb6cc0_7102,RIee20e90_4833,RIded8c08_930,
        RIded6778_904,RIded4720_881,RIded23f8_856,RIdecf9c8_826,RIdecccc8_794,RIdec9fc8_762,RIdec72c8_730,RIdeb37c8_506,RIde94850_314,RIe16d3d0_2620,
        RIe1591c8_2391,RIe1429c8_2135,RIdf373c0_2005,RIdf2ba20_1873,RIdf1c2a0_1697,RIdeff998_1372,RIdee6498_1084,RIdedb200_957,RIde7a798_187,RIe19c860_3158,
        RIe199b60_3126,RIf145220_5246,RIe196e60_3094,RIf144140_5234,RIe194160_3062,RIe191460_3030,RIe18e760_2998,RIe188d60_2934,RIe186060_2902,RIf1431c8_5223,
        RIe183360_2870,RIf142ac0_5218,RIe180660_2838,RIe17d960_2806,RIe17ac60_2774,RIf141cb0_5208,RIf140798_5193,RIf13ff28_5187,RIfe8be90_7936,RIfceb880_7702,
        RIf13eb78_5173,RIee3e008_5164,RIee3cdc0_5151,RIee3bb78_5138,RIee3aa98_5126,RIee396e8_5112,RIe172c68_2683,RIf16fac0_5730,RIf16ef80_5722,RIf16dbd0_5708,
        RIfcc4af0_7260,RIf16c820_5694,RIe222bb8_4685,RIf16b740_5682,RIe21feb8_4653,RIf16a7c8_5671,RIe21d1b8_4621,RIe2177b8_4557,RIe214ab8_4525,RIfe8c430_7940,
        RIe211db8_4493,RIf1688d8_5649,RIe20f0b8_4461,RIf167960_5638,RIe20c3b8_4429,RIe2096b8_4397,RIe2069b8_4365,RIf1669e8_5627,RIf165908_5615,RIfe8c9d0_7944,
        RIfe8c700_7942,RIfc9c578_6801,RIf163ce8_5595,RIf162d70_5584,RIf161588_5567,RIf15f698_5545,RIf15d910_5524,RIfe8c598_7941,RIfe8c868_7943,RIf15c3f8_5509,
        RIf15aee0_5494,RIf15a0d0_5484,RIf1596f8_5477,RIf158618_5465,RIf1573d0_5452,RIf156b60_5446,RIfec1f68_8327,RIf155eb8_5437,RIf155378_5429,RIf153fc8_5415,
        RIfe8bff8_7937,RIf152948_5399,RIf151598_5385,RIf150080_5370,RIfe8c2c8_7939,RIf14f270_5360,RIfc503a8_5935,RIf14d650_5340,RIfe8c160_7938,RIe1ea920_4046,
        RIe1e7c20_4014,RIe1e4f20_3982,RIe1e2220_3950,RIe1df520_3918,RIe1dc820_3886,RIe1d9b20_3854,RIe1d6e20_3822,RIe1d1420_3758,RIe1ce720_3726,RIe1cba20_3694,
        RIe1c8d20_3662,RIe1c6020_3630,RIe1c3320_3598,RIe1c0620_3566,RIe1bd920_3534,RIf14c2a0_5326,RIf14aef0_5312,RIe1b88f8_3477,RIe1b68a0_3454,RIfcd4db0_7444,
        RIfc4ebc0_5918,RIfec1e00_8326,RIfe8bd28_7935,RIf148790_5284,RIf1476b0_5272,RIfe8ba58_7933,RIfec1b30_8324,RIfc4e788_5915,RIfcb8e80_7126,RIfe8bbc0_7934,
        RIfec1c98_8325,RIe1a7c60_3286,RIe1a4f60_3254,RIe1a2260_3222,RIe19f560_3190,RIe18ba60_2966,RIe177f60_2742,RIe2258b8_4717,RIe21a4b8_4589,RIe203cb8_4333,
        RIe1fdd18_4265,RIe1f70d0_4188,RIe1efc18_4105,RIe1d4120_3790,RIe1bac20_3502,RIe1ada98_3353,RIe1700d0_2652,RIdec4a00_701,RIdec1d00_669,RIfcad7b0_6996,
        RIdebf000_637,RIfc64cb8_6169,RIdebc300_605,RIdeb9600_573,RIdeb6900_541,RIfc6f9b0_6292,RIdeb0f00_477,RIfc657f8_6177,RIdeae200_445,RIfce69c0_7646,
        RIdea8d28_413,RIdea2428_381,RIde9bb28_349,RIfc6fc80_6294,RIee1b760_4771,RIfca8080_6934,RIfe8b8f0_7932,RIde90020_292,RIde8c510_274,RIde89090_258,
        RIde84ba8_237,RIfc65ac8_6179,RIfcad210_6992,RIfcce168_7367,RIfcce2d0_7368,RIfc51488_5947,RIe16af40_2594,RIfc65c30_6180,RIe167598_2553,RIe164a00_2522,
        RIe161d00_2490,RIfc66e78_6193,RIe15f000_2458,RIfc6e498_6277,RIe15c300_2426,RIe156900_2362,RIe153c00_2330,RIfc6e330_6276,RIe150f00_2298,RIfccda60_7362,
        RIe14e200_2266,RIfc6e1c8_6275,RIe14b500_2234,RIe148800_2202,RIe145b00_2170,RIee33fb8_5050,RIee32d70_5037,RIee31c90_5025,RIee30fe8_5016,RIfea8630_8232,
        RIdf3e5a8_2086,RIdf3c550_2063,RIfea8798_8233,RIfc6e060_6274,RIfcac6d0_6984,RIfc56078_6001,RIfc6e600_6278,RIdf34dc8_1978,RIdf32d70_1955,RIfea84c8_8231,
        RIdf2eb58_1908,RIee2b750_4953,RIfc6ee70_6284,RIfc6efd8_6285,RIee27808_4908,RIfe8b788_7931,RIdf27ad8_1828,RIdf25d50_1807,RIdf24130_1787,RIfc66608_6187,
        RIfccde98_7365,RIfc66a40_6190,RIfc668d8_6189,RIfcacf40_6990,RIfeaaef8_8261,RIfc6e8d0_6280,RIdf18d30_1659,RIdf165d0_1631,RIdf138d0_1599,RIdf10bd0_1567,
        RIdf0ded0_1535,RIdf0b1d0_1503,RIdf084d0_1471,RIdf057d0_1439,RIdf02ad0_1407,RIdefd0d0_1343,RIdefa3d0_1311,RIdef76d0_1279,RIdef49d0_1247,RIdef1cd0_1215,
        RIdeeefd0_1183,RIdeec2d0_1151,RIdee95d0_1119,RIfc6dc28_6271,RIfc67c88_6203,RIfccb300_7334,RIfccd4c0_7358,RIfea81f8_8229,RIfea8360_8230,RIdee04f8_1016,
        RIdede338_992,RIfc6def8_6273,RIfcac130_6980,RIfc67b20_6202,RIfc67df0_6204,RIded9040_933,RIded6a48_906,RIded4b58_884,RIded26c8_858,RIdecfe00_829,
        RIdecd100_797,RIdeca400_765,RIdec7700_733,RIdeb3c00_509,RIde95228_317,RIe16d808_2623,RIe159600_2394,RIe142e00_2138,RIdf377f8_2008,RIdf2be58_1876,
        RIdf1c6d8_1700,RIdeffdd0_1375,RIdee68d0_1087,RIdedb638_960,RIde7b170_190,RIe19cc98_3161,RIe199f98_3129,RIfc73088_6331,RIe197298_3097,RIf1442a8_5235,
        RIe194598_3065,RIe191898_3033,RIe18eb98_3001,RIe189198_2937,RIe186498_2905,RIfc72278_6321,RIe183798_2873,RIfc61ce8_6135,RIe180a98_2841,RIe17dd98_2809,
        RIe17b098_2777,RIfcaf268_7015,RIfca6a00_6918,RIfcc9b18_7317,RIe175530_2712,RIfc72818_6325,RIfc726b0_6324,RIfccf7e8_7383,RIfc72548_6323,RIee3be48_5140,
        RIee3ad68_5128,RIfc71fa8_6319,RIe1730a0_2686,RIfcaef98_7013,RIfccf518_7381,RIfc71e40_6318,RIfc62120_6138,RIfe8b350_7928,RIe222ff0_4688,RIfcc9f50_7320,
        RIe2202f0_4656,RIfc4a570_5868,RIe21d5f0_4624,RIe217bf0_4560,RIe214ef0_4528,RIfccf3b0_7380,RIe2121f0_4496,RIf168ba8_5651,RIe20f4f0_4464,RIfc71300_6310,
        RIe20c7f0_4432,RIe209af0_4400,RIe206df0_4368,RIfc718a0_6314,RIfc71a08_6315,RIe202098_4313,RIfe8b1e8_7927,RIfc715d0_6312,RIfce6588_7643,RIfc62c60_6146,
        RIf161858_5569,RIf15fad0_5548,RIf15dbe0_5526,RIe1fc698_4249,RIfe8b4b8_7929,RIfcae5c0_7006,RIfc63098_6149,RIfc63200_6150,RIfc71198_6309,RIf158a50_5468,
        RIf1576a0_5454,RIfcdc808_7531,RIfe8b620_7930,RIfc634d0_6152,RIfcceb40_7374,RIf154400_5418,RIe1f4da8_4163,RIf152c18_5401,RIf151868_5387,RIfc4d108_5899,
        RIe1f2a80_4138,RIfc70a90_6304,RIfc63bd8_6157,RIfca7810_6928,RIe1ed788_4079,RIe1ead58_4049,RIe1e8058_4017,RIe1e5358_3985,RIe1e2658_3953,RIe1df958_3921,
        RIe1dcc58_3889,RIe1d9f58_3857,RIe1d7258_3825,RIe1d1858_3761,RIe1ceb58_3729,RIe1cbe58_3697,RIe1c9158_3665,RIe1c6458_3633,RIe1c3758_3601,RIe1c0a58_3569,
        RIe1bdd58_3537,RIf14c408_5327,RIf14b1c0_5314,RIe1b8d30_3480,RIe1b6cd8_3457,RIfc707c0_6302,RIfca7c48_6931,RIe1b4de8_3435,RIe1b3a38_3421,RIfc70220_6298,
        RIfcce870_7372,RIe1b23b8_3405,RIe1b0630_3384,RIfc645b0_6164,RIfc700b8_6297,RIfeaac28_8259,RIe1aa690_3316,RIe1a8098_3289,RIe1a5398_3257,RIe1a2698_3225,
        RIe19f998_3193,RIe18be98_2969,RIe178398_2745,RIe225cf0_4720,RIe21a8f0_4592,RIe2040f0_4336,RIe1fe150_4268,RIe1f7508_4191,RIe1f0050_4108,RIe1d4558_3793,
        RIe1bb058_3505,RIe1aded0_3356,RIe170508_2655,RIdec4898_700,RIdec1b98_668,RIfc661d0_6184,RIdebee98_636,RIfce6b28_7647,RIdebc198_604,RIdeb9498_572,
        RIdeb6798_540,RIfc40d18_5763,RIdeb0d98_476,RIfcad648_6995,RIdeae098_444,RIfcaa510_6960,RIdea89e0_412,RIdea20e0_380,RIde9b7e0_348,RIfcab320_6970,
        RIfca8350_6936,RIfc6f6e0_6290,RIfcaa240_6958,RIde8fcd8_291,RIfe8aae0_7922,RIde88d48_257,RIde84860_236,RIde80a08_217,RIfc64718_6165,RIfcae020_7002,
        RIfcadeb8_7001,RIee38fe0_5107,RIe16add8_2593,RIe1695f0_2576,RIe167430_2552,RIe164898_2521,RIe161b98_2489,RIfe8a3d8_7917,RIe15ee98_2457,RIfe8a270_7916,
        RIe15c198_2425,RIe156798_2361,RIe153a98_2329,RIfc3f0f8_5743,RIe150d98_2297,RIfcab050_6968,RIe14e098_2265,RIfcca658_7325,RIe14b398_2233,RIe148698_2201,
        RIe145998_2169,RIfe8a810_7920,RIfe8a6a8_7919,RIee31b28_5024,RIee30e80_5015,RIe140808_2111,RIfe8a540_7918,RIdf3c3e8_2062,RIdf3a0c0_2037,RIfc6b1f8_6241,
        RIee2f260_4995,RIfc70d60_6306,RIee2d0a0_4971,RIfe8a978_7921,RIdf32c08_1954,RIdf308e0_1929,RIdf2e9f0_1907,RIee2b5e8_4952,RIee29e00_4935,RIee28a50_4921,
        RIee276a0_4907,RIdf29c98_1852,RIdf27970_1827,RIdf25be8_1806,RIdf23fc8_1786,RIfc6aaf0_6236,RIfc6ac58_6237,RIdf22678_1768,RIfcdd4b0_7540,RIdf21160_1753,
        RIdf1f108_1730,RIdf1ac20_1681,RIfeaa7f0_8256,RIdf16468_1630,RIdf13768_1598,RIdf10a68_1566,RIdf0dd68_1534,RIdf0b068_1502,RIdf08368_1470,RIdf05668_1438,
        RIdf02968_1406,RIdefcf68_1342,RIdefa268_1310,RIdef7568_1278,RIdef4868_1246,RIdef1b68_1214,RIdeeee68_1182,RIdeec168_1150,RIdee9468_1118,RIee25378_4882,
        RIee24568_4872,RIee23a28_4864,RIee23050_4857,RIfe8adb0_7924,RIdee23e8_1038,RIfe8ac48_7923,RIdede1d0_991,RIfca5650_6904,RIee220d8_4846,RIfceeb20_7738,
        RIee20ff8_4834,RIded8ed8_932,RIfe8af18_7925,RIded49f0_883,RIfe8b080_7926,RIdecfc98_828,RIdeccf98_796,RIdeca298_764,RIdec7598_732,RIdeb3a98_508,
        RIde94ee0_316,RIe16d6a0_2622,RIe159498_2393,RIe142c98_2137,RIdf37690_2007,RIdf2bcf0_1875,RIdf1c570_1699,RIdeffc68_1374,RIdee6768_1086,RIdedb4d0_959,
        RIde7ae28_189,RIe19cb30_3160,RIe199e30_3128,RIf145388_5247,RIe197130_3096,RIfe8a108_7915,RIe194430_3064,RIe191730_3032,RIe18ea30_3000,RIe189030_2936,
        RIe186330_2904,RIfc6c878_6257,RIe183630_2872,RIfcabcf8_6977,RIe180930_2840,RIe17dc30_2808,RIe17af30_2776,RIfcccc50_7352,RIfcccdb8_7353,RIe176d18_2729,
        RIfea7af0_8224,RIfe89fa0_7914,RIfe89e38_7913,RIfcdd078_7537,RIfccb738_7337,RIfca9868_6951,RIfcabb90_6976,RIfca99d0_6952,RIe172f38_2685,RIf16fd90_5732,
        RIf16f250_5724,RIfc6c440_6254,RIfcaba28_6975,RIfc40610_5758,RIe222e88_4687,RIfc5d260_6082,RIe220188_4655,RIfcab758_6973,RIe21d488_4623,RIe217a88_4559,
        RIe214d88_4527,RIfe892f8_7905,RIe212088_4495,RIf168a40_5650,RIe20f388_4463,RIf167ac8_5639,RIe20c688_4431,RIe209988_4399,RIe206c88_4367,RIfc6c2d8_6253,
        RIfceec88_7739,RIe201f30_4312,RIe200748_4295,RIf164dc8_5607,RIf163fb8_5597,RIf163040_5586,RIfe895c8_7907,RIf15f968_5547,RIfe89898_7909,RIfe89460_7906,
        RIe1fb5b8_4237,RIf15c6c8_5511,RIfe89730_7908,RIf15a238_5485,RIf1599c8_5479,RIf1588e8_5467,RIfe89cd0_7912,RIfc5ba78_6065,RIe1f9c68_4219,RIfc5bd48_6067,
        RIf1554e0_5430,RIf154298_5417,RIe1f4c40_4162,RIfe89b68_7911,RIfe89a00_7910,RIf150350_5372,RIe1f2918_4137,RIf14f3d8_5361,RIfccc818_7349,RIf14d920_5342,
        RIe1ed620_4078,RIe1eabf0_4048,RIe1e7ef0_4016,RIe1e51f0_3984,RIe1e24f0_3952,RIe1df7f0_3920,RIe1dcaf0_3888,RIe1d9df0_3856,RIe1d70f0_3824,RIe1d16f0_3760,
        RIe1ce9f0_3728,RIe1cbcf0_3696,RIe1c8ff0_3664,RIe1c62f0_3632,RIe1c35f0_3600,RIe1c08f0_3568,RIe1bdbf0_3536,RIfc680c0_6206,RIf14b058_5313,RIe1b8bc8_3479,
        RIe1b6b70_3456,RIfcac298_6981,RIf1499d8_5297,RIfe89190_7904,RIfec19c8_8323,RIf148a60_5286,RIfccdd30_7364,RIe1b2250_3404,RIfec1860_8322,RIfc6e768_6279,
        RIfc54728_5983,RIe1abfe0_3334,RIe1aa528_3315,RIe1a7f30_3288,RIe1a5230_3256,RIe1a2530_3224,RIe19f830_3192,RIe18bd30_2968,RIe178230_2744,RIe225b88_4719,
        RIe21a788_4591,RIe203f88_4335,RIe1fdfe8_4267,RIe1f73a0_4190,RIe1efee8_4107,RIe1d43f0_3792,RIe1baef0_3504,RIe1add68_3355,RIe1703a0_2654,RIdec4cd0_703,
        RIdec1fd0_671,RIfc7b4b8_6425,RIdebf2d0_639,RIfc7b1e8_6423,RIdebc5d0_607,RIdeb98d0_575,RIdeb6bd0_543,RIfe83358_7837,RIdeb11d0_479,RIee1e5c8_4804,
        RIdeae4d0_447,RIfc437c0_5790,RIdea93b8_415,RIdea2ab8_383,RIde9c1b8_351,RIfc90ea8_6671,RIfc7af18_6421,RIfe83088_7835,RIee1a950_4761,RIde906b0_294,
        RIde8cba0_276,RIfe82f20_7834,RIfe82db8_7833,RIee1a248_4756,RIfe831f0_7836,RIfcc2390_7232,RIee195a0_4747,RIfcbe718_7189,RIfea9e18_8249,RIfc43220_5786,
        RIe167868_2555,RIe164cd0_2524,RIe161fd0_2492,RIee36f88_5084,RIe15f2d0_2460,RIee35ea8_5072,RIe15c5d0_2428,RIe156bd0_2364,RIe153ed0_2332,RIfe83628_7839,
        RIe1511d0_2300,RIfebfda8_8303,RIe14e4d0_2268,RIfebfc40_8302,RIe14b7d0_2236,RIe148ad0_2204,RIe145dd0_2172,RIee34120_5051,RIee32ed8_5038,RIee31df8_5026,
        RIfcc1f58_7229,RIe140ad8_2113,RIdf3e878_2088,RIfe834c0_7838,RIdf3a390_2039,RIfc5a6c8_6051,RIfc91e20_6682,RIee2e888_4988,RIfc96a10_6736,RIdf35098_1980,
        RIfeab600_8266,RIdf30bb0_1931,RIfeab768_8267,RIfcbe9e8_7191,RIfc79fa0_6410,RIfc96740_6734,RIfc92258_6685,RIfea7118_8217,RIfea95a8_8243,RIdf26020_1809,
        RIdf24400_1789,RIfc79a00_6406,RIfc5add0_6056,RIfce5d18_7637,RIfc92690_6688,RIfce3018_7605,RIdf1f270_1731,RIfc79730_6404,RIdf19000_1661,RIdf168a0_1633,
        RIdf13ba0_1601,RIdf10ea0_1569,RIdf0e1a0_1537,RIdf0b4a0_1505,RIdf087a0_1473,RIdf05aa0_1441,RIdf02da0_1409,RIdefd3a0_1345,RIdefa6a0_1313,RIdef79a0_1281,
        RIdef4ca0_1249,RIdef1fa0_1217,RIdeef2a0_1185,RIdeec5a0_1153,RIdee98a0_1121,RIfc5b7a8_6063,RIfc5b640_6062,RIfc931d0_6696,RIfcecac8_7715,RIdee4710_1063,
        RIdee26b8_1040,RIdee07c8_1018,RIdede4a0_993,RIfcbf0f0_7196,RIfcbf528_7199,RIfc792f8_6401,RIfc93068_6695,RIded91a8_934,RIded6d18_908,RIded4e28_886,
        RIded2998_860,RIded00d0_831,RIdecd3d0_799,RIdeca6d0_767,RIdec79d0_735,RIdeb3ed0_511,RIde958b8_319,RIe16dad8_2625,RIe1598d0_2396,RIe1430d0_2140,
        RIdf37ac8_2010,RIdf2c128_1878,RIdf1c9a8_1702,RIdf000a0_1377,RIdee6ba0_1089,RIdedb908_962,RIde7b800_192,RIe19cf68_3163,RIe19a268_3131,RIfc8d7d0_6632,
        RIe197568_3099,RIfc561e0_6002,RIe194868_3067,RIe191b68_3035,RIe18ee68_3003,RIe189468_2939,RIe186768_2907,RIf143330_5224,RIe183a68_2875,RIfc7d948_6451,
        RIe180d68_2843,RIe17e068_2811,RIe17b368_2779,RIfc564b0_6004,RIfcd6700_7462,RIfc461f0_5820,RIe175698_2713,RIfc46088_5819,RIfc45f20_5818,RIfc7dc18_6453,
        RIfcd69d0_7464,RIfc98630_6756,RIfcc2a98_7237,RIfc7d510_6448,RIe173208_2687,RIfc8e478_6641,RIfc45ae8_5815,RIfc8e8b0_6644,RIfc45980_5814,RIfe82ae8_7831,
        RIe2232c0_4690,RIf16ba10_5684,RIe2205c0_4658,RIfcd24e8_7415,RIe21d8c0_4626,RIe217ec0_4562,RIe2151c0_4530,RIfebf268_8295,RIe2124c0_4498,RIf168d10_5652,
        RIe20f7c0_4466,RIfc7d240_6446,RIe20cac0_4434,RIe209dc0_4402,RIe2070c0_4370,RIf166e20_5630,RIfebf6a0_8298,RIfebf808_8299,RIfebf538_8297,RIfc8eb80_6646,
        RIf164120_5598,RIfc453e0_5810,RIf161b28_5571,RIf15fc38_5549,RIf15dd48_5527,RIe1fc968_4251,RIe1fb888_4239,RIfebf3d0_8296,RIf15b318_5497,RIfca2518_6869,
        RIfc8f120_6650,RIfebfad8_8301,RIfebf970_8300,RIfc7cca0_6442,RIe1f9dd0_4220,RIfe82c50_7832,RIf155648_5431,RIfc8f288_6651,RIe1f4f10_4164,RIf152d80_5402,
        RIfc8f828_6655,RIfcb3b88_7067,RIe1f2d50_4140,RIfc445d0_5800,RIfc8faf8_6657,RIf14da88_5343,RIe1eda58_4081,RIe1eb028_4051,RIe1e8328_4019,RIe1e5628_3987,
        RIe1e2928_3955,RIe1dfc28_3923,RIe1dcf28_3891,RIe1da228_3859,RIe1d7528_3827,RIe1d1b28_3763,RIe1cee28_3731,RIe1cc128_3699,RIe1c9428_3667,RIe1c6728_3635,
        RIe1c3a28_3603,RIe1c0d28_3571,RIe1be028_3539,RIfc7bff8_6433,RIfc44030_5796,RIe1b9000_3482,RIe1b6fa8_3459,RIfcbdd40_7182,RIfc8ff30_6660,RIe1b50b8_3437,
        RIe1b3d08_3423,RIfcbe178_7185,RIfc43d60_5794,RIe1b2520_3406,RIe1b0798_3385,RIfcdb5c0_7518,RIfc7ba58_6429,RIe1ac148_3335,RIe1aa960_3318,RIe1a8368_3291,
        RIe1a5668_3259,RIe1a2968_3227,RIe19fc68_3195,RIe18c168_2971,RIe178668_2747,RIe225fc0_4722,RIe21abc0_4594,RIe2043c0_4338,RIe1fe420_4270,RIe1f77d8_4193,
        RIe1f0320_4110,RIe1d4828_3795,RIe1bb328_3507,RIe1ae1a0_3358,RIe1707d8_2657,RIdec4b68_702,RIdec1e68_670,RIfc5df08_6091,RIdebf168_638,RIfce6df8_7649,
        RIdebc468_606,RIdeb9768_574,RIdeb6a68_542,RIfc75ef0_6364,RIdeb1068_478,RIfcc12b0_7220,RIdeae368_446,RIfc5e340_6094,RIdea9070_414,RIdea2770_382,
        RIde9be70_350,RIfced4a0_7722,RIfcc1418_7221,RIfc95930_6724,RIfcec0f0_7708,RIde90368_293,RIde8c858_275,RIde893d8_259,RIde84ef0_238,RIde80d50_218,
        RIfc95a98_6725,RIfced068_7719,RIfced1d0_7720,RIfcedfe0_7730,RIe16b0a8_2595,RIe169758_2577,RIe167700_2554,RIe164b68_2523,RIe161e68_2491,RIee36e20_5083,
        RIe15f168_2459,RIfc426e0_5778,RIe15c468_2427,RIe156a68_2363,RIe153d68_2331,RIfe82818_7829,RIe151068_2299,RIee34c60_5059,RIe14e368_2267,RIfc5f9c0_6110,
        RIe14b668_2235,RIe148968_2203,RIe145c68_2171,RIfccfef0_7388,RIfca57b8_6905,RIfc600c8_6115,RIfcafda8_7023,RIe140970_2112,RIdf3e710_2087,RIdf3c6b8_2064,
        RIdf3a228_2038,RIfc5fc90_6112,RIee2f3c8_4996,RIfc742d0_6344,RIee2d208_4972,RIdf34f30_1979,RIfebf100_8294,RIdf30a48_1930,RIdf2ecc0_1909,RIfcb08e8_7031,
        RIfcee418_7733,RIfc95ed0_6728,RIfcdef68_7559,RIdf29e00_1853,RIdf27c40_1829,RIdf25eb8_1808,RIdf24298_1788,RIfc5ed18_6101,RIfcee850_7736,RIdf227e0_1769,
        RIfc5efe8_6103,RIdf212c8_1754,RIfeaa520_8254,RIdf1ad88_1682,RIdf18e98_1660,RIdf16738_1632,RIdf13a38_1600,RIdf10d38_1568,RIdf0e038_1536,RIdf0b338_1504,
        RIdf08638_1472,RIdf05938_1440,RIdf02c38_1408,RIdefd238_1344,RIdefa538_1312,RIdef7838_1280,RIdef4b38_1248,RIdef1e38_1216,RIdeef138_1184,RIdeec438_1152,
        RIdee9738_1120,RIfcc96e0_7314,RIfccfd88_7387,RIfc60aa0_6122,RIfca5ec0_6910,RIdee45a8_1062,RIdee2550_1039,RIdee0660_1017,RIfe826b0_7828,RIfcdeb30_7556,
        RIfc73bc8_6339,RIfca5bf0_6908,RIfc73a60_6338,RIfe82980_7830,RIded6bb0_907,RIded4cc0_885,RIded2830_859,RIdecff68_830,RIdecd268_798,RIdeca568_766,
        RIdec7868_734,RIdeb3d68_510,RIde95570_318,RIe16d970_2624,RIe159768_2395,RIe142f68_2139,RIdf37960_2009,RIdf2bfc0_1877,RIdf1c840_1701,RIdefff38_1376,
        RIdee6a38_1088,RIdedb7a0_961,RIde7b4b8_191,RIe19ce00_3162,RIe19a100_3130,RIfce96c0_7678,RIe197400_3098,RIf144410_5236,RIe194700_3066,RIe191a00_3034,
        RIe18ed00_3002,RIe189300_2938,RIe186600_2906,RIfebee30_8292,RIe183900_2874,RIfcdbcc8_7523,RIe180c00_2842,RIe17df00_2810,RIe17b200_2778,RIf141f80_5210,
        RIfce7398_7653,RIfcb1e00_7046,RIfe82548_7827,RIfca42a0_6890,RIfcbff00_7206,RIfcaaee8_6967,RIee3d090_5153,RIfc5c180_6070,RIfce35b8_7609,RIee399b8_5114,
        RIfea8a68_8235,RIf16fef8_5733,RIfebecc8_8291,RIfc5c450_6072,RIfce9288_7675,RIfc40778_5759,RIe223158_4689,RIfce77d0_7656,RIe220458_4657,RIfce24d8_7597,
        RIe21d758_4625,RIe217d58_4561,RIe215058_4529,RIfce8a18_7669,RIe212358_4497,RIfce1998_7589,RIe20f658_4465,RIfc77840_6382,RIe20c958_4433,RIe209c58_4401,
        RIe206f58_4369,RIf166cb8_5629,RIf165bd8_5617,RIfe81fa8_7823,RIfe81e40_7822,RIfc5c888_6075,RIfceb178_7697,RIf1631a8_5587,RIf1619c0_5570,RIfccf248_7379,
        RIfc77570_6380,RIe1fc800_4250,RIe1fb720_4238,RIf15c830_5512,RIf15b1b0_5496,RIfcd0fd0_7400,RIfccc6b0_7348,RIf158bb8_5469,RIf157808_5455,RIfc5d0f8_6081,
        RIfebef98_8293,RIfcc8a38_7305,RIfcd7ab0_7476,RIfcb1428_7039,RIfeaa0e8_8251,RIfccc548_7347,RIfce3450_7608,RIf1504b8_5373,RIe1f2be8_4139,RIf14f540_5362,
        RIfc772a0_6378,RIfcec258_7709,RIe1ed8f0_4080,RIe1eaec0_4050,RIe1e81c0_4018,RIe1e54c0_3986,RIe1e27c0_3954,RIe1dfac0_3922,RIe1dcdc0_3890,RIe1da0c0_3858,
        RIe1d73c0_3826,RIe1d19c0_3762,RIe1cecc0_3730,RIe1cbfc0_3698,RIe1c92c0_3666,RIe1c65c0_3634,RIe1c38c0_3602,RIe1c0bc0_3570,RIe1bdec0_3538,RIf14c570_5328,
        RIf14b328_5315,RIe1b8e98_3481,RIe1b6e40_3458,RIfc76760_6370,RIfc94b20_6714,RIe1b4f50_3436,RIe1b3ba0_3422,RIfcec3c0_7710,RIfceb010_7696,RIfe823e0_7826,
        RIfe82110_7824,RIfcdd8e8_7543,RIfcc0ba8_7215,RIfe82278_7825,RIe1aa7f8_3317,RIe1a8200_3290,RIe1a5500_3258,RIe1a2800_3226,RIe19fb00_3194,RIe18c000_2970,
        RIe178500_2746,RIe225e58_4721,RIe21aa58_4593,RIe204258_4337,RIe1fe2b8_4269,RIe1f7670_4192,RIe1f01b8_4109,RIe1d46c0_3794,RIe1bb1c0_3506,RIe1ae038_3357,
        RIe170670_2656,RIdec4fa0_705,RIdec22a0_673,RIee1fdb0_4821,RIdebf5a0_641,RIee1f270_4813,RIdebc8a0_609,RIdeb9ba0_577,RIdeb6ea0_545,RIee1ecd0_4809,
        RIdeb14a0_481,RIee1e730_4805,RIdeae7a0_449,RIee1d920_4795,RIdea9a48_417,RIdea3148_385,RIde9c848_353,RIee1cb10_4785,RIee1ba30_4773,RIee1b1c0_4767,
        RIfec04b0_8308,RIfe850e0_7858,RIde8d230_278,RIfea9cb0_8248,RIfe84f78_7857,RIee1a3b0_4757,RIfe853b0_7860,RIee199d8_4750,RIfe85248_7859,RIee39148_5108,
        RIe16b378_2597,RIee38608_5100,RIe167b38_2557,RIe164fa0_2526,RIe1622a0_2494,RIfe85950_7864,RIe15f5a0_2462,RIee36010_5073,RIe15c8a0_2430,RIe156ea0_2366,
        RIe1541a0_2334,RIfe85c20_7866,RIe1514a0_2302,RIee34dc8_5060,RIe14e7a0_2270,RIfc861b0_6548,RIe14baa0_2238,RIe148da0_2206,RIe1460a0_2174,RIee343f0_5053,
        RIfe85518_7861,RIfe857e8_7863,RIfe85680_7862,RIe140c40_2114,RIdf3eb48_2090,RIdf3c820_2065,RIdf3a660_2041,RIfc9d4f0_6812,RIee2f698_4998,RIfc52298_5957,
        RIee2d4d8_4974,RIdf35368_1982,RIdf32ed8_1956,RIdf30e80_1933,RIfe85ab8_7865,RIee2b8b8_4954,RIee29f68_4936,RIee28bb8_4922,RIee27970_4909,RIdf2a0d0_1855,
        RIfe84e10_7856,RIdf262f0_1811,RIfe84ca8_7855,RIee27100_4903,RIee26b60_4899,RIfcd32f8_7425,RIee265c0_4895,RIfc9e300_6822,RIdf1f540_1733,RIee25eb8_4890,
        RIfe84b40_7854,RIdf16b70_1635,RIdf13e70_1603,RIdf11170_1571,RIdf0e470_1539,RIdf0b770_1507,RIdf08a70_1475,RIdf05d70_1443,RIdf03070_1411,RIdefd670_1347,
        RIdefa970_1315,RIdef7c70_1283,RIdef4f70_1251,RIdef2270_1219,RIdeef570_1187,RIdeec870_1155,RIdee9b70_1123,RIfec0348_8307,RIfcb54d8_7085,RIee23cf8_4866,
        RIfc54e30_5988,RIfec0078_8305,RIdee2988_1042,RIfec01e0_8306,RIdede770_995,RIfcd7ee8_7479,RIfcd43d8_7437,RIfc88eb0_6580,RIfc9e5d0_6824,RIded9478_936,
        RIded6fe8_910,RIded50f8_888,RIfeab330_8264,RIded03a0_833,RIdecd6a0_801,RIdeca9a0_769,RIdec7ca0_737,RIdeb41a0_513,RIde95f48_321,RIe16dda8_2627,
        RIe159ba0_2398,RIe1433a0_2142,RIdf37d98_2012,RIdf2c3f8_1880,RIdf1cc78_1704,RIdf00370_1379,RIdee6e70_1091,RIdedbbd8_964,RIde7be90_194,RIe19d238_3165,
        RIe19a538_3133,RIf145658_5249,RIe197838_3101,RIf1446e0_5238,RIe194b38_3069,RIe191e38_3037,RIe18f138_3005,RIe189738_2941,RIe186a38_2909,RIf143600_5226,
        RIe183d38_2877,RIf142c28_5219,RIe181038_2845,RIe17e338_2813,RIe17b638_2781,RIf1420e8_5211,RIf140a68_5195,RIf1401f8_5189,RIfebff10_8304,RIf13faf0_5184,
        RIf13ee48_5175,RIee3e2d8_5166,RIee3d1f8_5154,RIee3c118_5142,RIee3b038_5130,RIee39c88_5116,RIfe838f8_7841,RIf1701c8_5735,RIfc5ab00_6054,RIf16e008_5711,
        RIfcb0e88_7035,RIf16caf0_5696,RIe223590_4692,RIf16bce0_5686,RIe220890_4660,RIf16ac00_5674,RIe21db90_4628,RIe218190_4564,RIe215490_4532,RIf16a228_5667,
        RIe212790_4500,RIf168fe0_5654,RIe20fa90_4468,RIf167d98_5641,RIe20cd90_4436,RIe20a090_4404,RIe207390_4372,RIf1670f0_5632,RIf165ea8_5619,RIe202200_4314,
        RIfe83e98_7845,RIf164f30_5608,RIf1643f0_5600,RIfce8310_7664,RIf161df8_5573,RIf15ff08_5551,RIf15e018_5529,RIfe83d30_7844,RIfe84000_7846,RIf15cb00_5514,
        RIf15b5e8_5499,RIf15a508_5487,RIfc887a8_6575,RIf158d20_5470,RIf157970_5456,RIf156cc8_5447,RIfe84438_7849,RIf156020_5438,RIfc51fc8_5955,RIf154568_5419,
        RIe1f51e0_4166,RIf153050_5404,RIf1519d0_5388,RIf150788_5375,RIfe842d0_7848,RIf14f810_5364,RIf14eb68_5355,RIf14dd58_5345,RIfe84168_7847,RIe1eb2f8_4053,
        RIe1e85f8_4021,RIe1e58f8_3989,RIe1e2bf8_3957,RIe1dfef8_3925,RIe1dd1f8_3893,RIe1da4f8_3861,RIe1d77f8_3829,RIe1d1df8_3765,RIe1cf0f8_3733,RIe1cc3f8_3701,
        RIe1c96f8_3669,RIe1c69f8_3637,RIe1c3cf8_3605,RIe1c0ff8_3573,RIe1be2f8_3541,RIf14c840_5330,RIf14b5f8_5317,RIfe83a60_7842,RIfe849d8_7853,RIfc74168_6343,
        RIf149b40_5298,RIfe83bc8_7843,RIfe84708_7851,RIf148d30_5288,RIf147ae8_5275,RIfe84870_7852,RIe1b0900_3386,RIf146fa8_5267,RIf146300_5258,RIfe845a0_7850,
        RIfe83790_7840,RIe1a8638_3293,RIe1a5938_3261,RIe1a2c38_3229,RIe19ff38_3197,RIe18c438_2973,RIe178938_2749,RIe226290_4724,RIe21ae90_4596,RIe204690_4340,
        RIe1fe6f0_4272,RIe1f7aa8_4195,RIe1f05f0_4112,RIe1d4af8_3797,RIe1bb5f8_3509,RIe1ae470_3360,RIe170aa8_2659,RIdec4e38_704,RIdec2138_672,RIee1fc48_4820,
        RIdebf438_640,RIfc49490_5856,RIdebc738_608,RIdeb9a38_576,RIdeb6d38_544,RIfc48ef0_5852,RIdeb1338_480,RIfcd9b08_7499,RIdeae638_448,RIfc8b610_6608,
        RIdea9700_416,RIdea2e00_384,RIde9c500_352,RIee1c9a8_4784,RIee1b8c8_4772,RIfc80918_6485,RIfcdad50_7512,RIfe86e68_7879,RIde8cee8_277,RIfe86d00_7878,
        RIfec0d20_8314,RIde81098_219,RIfc8b8e0_6610,RIfcd2d58_7421,RIfce4530_7620,RIfc8ba48_6611,RIe16b210_2596,RIe1698c0_2578,RIe1679d0_2556,RIe164e38_2525,
        RIe162138_2493,RIee370f0_5085,RIe15f438_2461,RIfc999e0_6770,RIe15c738_2429,RIe156d38_2365,RIe154038_2333,RIfc3f260_5744,RIe151338_2301,RIfc48518_5845,
        RIe14e638_2269,RIfc99e18_6773,RIe14b938_2237,RIe148c38_2205,RIe145f38_2173,RIee34288_5052,RIee33040_5039,RIee31f60_5027,RIfcd99a0_7498,RIfe86b98_7877,
        RIdf3e9e0_2089,RIfe86a30_7876,RIdf3a4f8_2040,RIfcc3470_7244,RIee2f530_4997,RIfc7fdd8_6477,RIee2d370_4973,RIdf35200_1981,RIfec0ff0_8316,RIdf30d18_1932,
        RIfec0e88_8315,RIfcd2a88_7419,RIfc8c858_6621,RIfc47ca8_5839,RIfcd6430_7460,RIdf29f68_1854,RIdf27da8_1830,RIdf26188_1810,RIdf24568_1790,RIfc8cb28_6623,
        RIfcdb188_7515,RIdf22948_1770,RIfc475a0_5834,RIdf21430_1755,RIdf1f3d8_1732,RIfec0bb8_8313,RIfe868c8_7875,RIdf16a08_1634,RIdf13d08_1602,RIdf11008_1570,
        RIdf0e308_1538,RIdf0b608_1506,RIdf08908_1474,RIdf05c08_1442,RIdf02f08_1410,RIdefd508_1346,RIdefa808_1314,RIdef7b08_1282,RIdef4e08_1250,RIdef2108_1218,
        RIdeef408_1186,RIdeec708_1154,RIdee9a08_1122,RIee254e0_4883,RIee246d0_4873,RIee23b90_4865,RIee231b8_4858,RIfe86fd0_7880,RIdee2820_1041,RIdee0930_1019,
        RIdede608_994,RIfc55da8_5999,RIfc98a68_6759,RIfcc3038_7241,RIfc464c0_5822,RIded9310_935,RIded6e80_909,RIded4f90_887,RIded2b00_861,RIded0238_832,
        RIdecd538_800,RIdeca838_768,RIdec7b38_736,RIdeb4038_512,RIde95c00_320,RIe16dc40_2626,RIe159a38_2397,RIe143238_2141,RIdf37c30_2011,RIdf2c290_1879,
        RIdf1cb10_1703,RIdf00208_1378,RIdee6d08_1090,RIdedba70_963,RIde7bb48_193,RIe19d0d0_3164,RIe19a3d0_3132,RIf1454f0_5248,RIe1976d0_3100,RIf144578_5237,
        RIe1949d0_3068,RIe191cd0_3036,RIe18efd0_3004,RIe1895d0_2940,RIe1868d0_2908,RIf143498_5225,RIe183bd0_2876,RIfc51758_5949,RIe180ed0_2844,RIe17e1d0_2812,
        RIe17b4d0_2780,RIfc9b060_6786,RIfc9ee40_6830,RIe176e80_2730,RIe175800_2714,RIfcb70f8_7105,RIfce0cf0_7580,RIfcc4280_7254,RIfcba7d0_7144,RIee3bfb0_5141,
        RIee3aed0_5129,RIee39b20_5115,RIe173370_2688,RIf170060_5734,RIf16f3b8_5725,RIf16dea0_5710,RIf16d4c8_5703,RIf16c988_5695,RIe223428_4691,RIf16bb78_5685,
        RIe220728_4659,RIf16aa98_5673,RIe21da28_4627,RIe218028_4563,RIe215328_4531,RIf16a0c0_5666,RIe212628_4499,RIf168e78_5653,RIe20f928_4467,RIf167c30_5640,
        RIe20cc28_4435,RIe209f28_4403,RIe207228_4371,RIf166f88_5631,RIf165d40_5618,RIfec0618_8309,RIfe86760_7874,RIfc52b08_5963,RIf164288_5599,RIf163310_5588,
        RIf161c90_5572,RIf15fda0_5550,RIf15deb0_5528,RIfe865f8_7873,RIfe85d88_7867,RIf15c998_5513,RIf15b480_5498,RIf15a3a0_5486,RIf159b30_5480,RIfc83348_6515,
        RIfc4ade0_5874,RIfc89720_6586,RIe1f9f38_4221,RIfc4ac78_5873,RIfc9f110_6832,RIfc4ab10_5872,RIe1f5078_4165,RIf152ee8_5403,RIfc899f0_6588,RIf150620_5374,
        RIe1f2eb8_4141,RIf14f6a8_5363,RIf14ea00_5354,RIf14dbf0_5344,RIe1edbc0_4082,RIe1eb190_4052,RIe1e8490_4020,RIe1e5790_3988,RIe1e2a90_3956,RIe1dfd90_3924,
        RIe1dd090_3892,RIe1da390_3860,RIe1d7690_3828,RIe1d1c90_3764,RIe1cef90_3732,RIe1cc290_3700,RIe1c9590_3668,RIe1c6890_3636,RIe1c3b90_3604,RIe1c0e90_3572,
        RIe1be190_3540,RIf14c6d8_5329,RIf14b490_5316,RIfe85ef0_7868,RIfe86490_7872,RIf14a248_5303,RIfc819f8_6497,RIfec0a50_8312,RIfe861c0_7870,RIf148bc8_5287,
        RIf147980_5274,RIfe86328_7871,RIfec0780_8310,RIfcbb478_7153,RIf146198_5257,RIfe86058_7869,RIfec08e8_8311,RIe1a84d0_3292,RIe1a57d0_3260,RIe1a2ad0_3228,
        RIe19fdd0_3196,RIe18c2d0_2972,RIe1787d0_2748,RIe226128_4723,RIe21ad28_4595,RIe204528_4339,RIe1fe588_4271,RIe1f7940_4194,RIe1f0488_4111,RIe1d4990_3796,
        RIe1bb490_3508,RIe1ae308_3359,RIe170940_2658,RIdec53d8_708,RIdec26d8_676,RIee20080_4823,RIdebf9d8_644,RIee1f3d8_4814,RIdebccd8_612,RIdeb9fd8_580,
        RIdeb72d8_548,RIee1ee38_4810,RIdeb18d8_484,RIee1e898_4806,RIdeaebd8_452,RIee1da88_4796,RIdeaa420_420,RIdea3b20_388,RIde9d220_356,RIee1cde0_4787,
        RIee1bd00_4775,RIee1b490_4769,RIfcd8a28_7487,RIde91088_297,RIde8d8c0_280,RIfe7dac0_7774,RIfe7d958_7773,RIee1a518_4758,RIee19e10_4753,RIee19b40_4751,
        RIfc768c8_6371,RIfcd05f8_7393,RIfe7dd90_7776,RIee38770_5101,RIfe7dc28_7775,RIe1653d8_2529,RIe1626d8_2497,RIee373c0_5087,RIe15f9d8_2465,RIee362e0_5075,
        RIe15ccd8_2433,RIe1572d8_2369,RIe1545d8_2337,RIfe7def8_7777,RIe1518d8_2305,RIfebdeb8_8281,RIe14ebd8_2273,RIfc649e8_6167,RIe14bed8_2241,RIe1491d8_2209,
        RIe1464d8_2177,RIfe7d7f0_7772,RIfe7d688_7771,RIee32230_5029,RIfceb9e8_7703,RIfebdd50_8280,RIfe7d520_7770,RIfebdbe8_8279,RIfe7d3b8_7769,RIfc734c0_6334,
        RIee2f968_5000,RIfccfab8_7385,RIee2d7a8_4976,RIdf357a0_1985,RIdf33310_1959,RIdf312b8_1936,RIdf2f0f8_1912,RIee2bcf0_4957,RIee2a238_4938,RIee28e88_4924,
        RIee27c40_4911,RIfe7ce18_7765,RIfe7ccb0_7764,RIfe7cf80_7766,RIfe7cb48_7763,RIee27268_4904,RIee26e30_4901,RIee26890_4897,RIfcaa0d8_6957,RIee262f0_4893,
        RIfe7d250_7768,RIee26020_4891,RIfe7d0e8_7767,RIdf16fa8_1638,RIdf142a8_1606,RIdf115a8_1574,RIdf0e8a8_1542,RIdf0bba8_1510,RIdf08ea8_1478,RIdf061a8_1446,
        RIdf034a8_1414,RIdefdaa8_1350,RIdefada8_1318,RIdef80a8_1286,RIdef53a8_1254,RIdef26a8_1222,RIdeef9a8_1190,RIdeecca8_1158,RIdee9fa8_1126,RIee25648_4884,
        RIee249a0_4875,RIfebe020_8282,RIee23488_4860,RIfebe2f0_8284,RIfebe188_8283,RIfe7e1c8_7779,RIfe7e060_7778,RIfcbf7f8_7201,RIfc7aae0_6418,RIfc787b8_6393,
        RIfc618b0_6132,RIded98b0_939,RIded72b8_912,RIded5530_891,RIded2dd0_863,RIded07d8_836,RIdecdad8_804,RIdecadd8_772,RIdec80d8_740,RIdeb45d8_516,
        RIde96920_324,RIe16e1e0_2630,RIe159fd8_2401,RIe1437d8_2145,RIdf381d0_2015,RIdf2c830_1883,RIdf1d0b0_1707,RIdf007a8_1382,RIdee72a8_1094,RIdedc010_967,
        RIde7c868_197,RIe19d670_3168,RIe19a970_3136,RIfe7b630_7748,RIe197c70_3104,RIfe7b4c8_7747,RIe194f70_3072,RIe192270_3040,RIe18f570_3008,RIe189b70_2944,
        RIe186e70_2912,RIfe7b360_7746,RIe184170_2880,RIfe7b1f8_7745,RIe181470_2848,RIe17e770_2816,RIe17ba70_2784,RIf1423b8_5213,RIf140ea0_5198,RIf140360_5190,
        RIfe7b798_7749,RIf13fc58_5185,RIf13f280_5178,RIfc79460_6402,RIee3d4c8_5156,RIfe7b090_7744,RIfe7af28_7743,RIee39df0_5117,RIe1737a8_2691,RIfe7adc0_7742,
        RIfe7ac58_7741,RIf16e440_5714,RIfcb20d0_7048,RIfe7bd38_7753,RIe2239c8_4695,RIf16be48_5687,RIe220cc8_4663,RIf16aed0_5676,RIe21dfc8_4631,RIe2185c8_4567,
        RIe2158c8_4535,RIfebd7b0_8276,RIe212bc8_4503,RIfebd648_8275,RIe20fec8_4471,RIfe7b900_7750,RIe20d1c8_4439,RIe20a4c8_4407,RIe2077c8_4375,RIf167258_5633,
        RIf166178_5621,RIe2024d0_4316,RIfe7bbd0_7752,RIf165368_5611,RIf1646c0_5602,RIfcd0a30_7396,RIf1620c8_5575,RIf1601d8_5553,RIf15e2e8_5531,RIfe7ba68_7751,
        RIfe7bea0_7754,RIf15cdd0_5516,RIf15b8b8_5501,RIf15a7d8_5489,RIfca4840_6894,RIf158ff0_5472,RIf157c40_5458,RIf156f98_5449,RIfe7c170_7756,RIf156458_5441,
        RIf155918_5433,RIf1549a0_5422,RIe1f54b0_4168,RIfe7c008_7755,RIf151b38_5389,RIf150bc0_5378,RIe1f32f0_4144,RIf14fae0_5366,RIf14ee38_5357,RIf14e028_5347,
        RIe1edff8_4085,RIe1eb730_4056,RIe1e8a30_4024,RIe1e5d30_3992,RIe1e3030_3960,RIe1e0330_3928,RIe1dd630_3896,RIe1da930_3864,RIe1d7c30_3832,RIe1d2230_3768,
        RIe1cf530_3736,RIe1cc830_3704,RIe1c9b30_3672,RIe1c6e30_3640,RIe1c4130_3608,RIe1c1430_3576,RIe1be730_3544,RIf14cb10_5332,RIf14b8c8_5319,RIfebda80_8278,
        RIfe7c878_7761,RIf14a680_5306,RIfe7c2d8_7757,RIfe7c9e0_7762,RIfe7c440_7758,RIf149000_5290,RIf147db8_5277,RIe1b2688_3407,RIfebd918_8277,RIfe7c5a8_7759,
        RIf146738_5261,RIfe7c710_7760,RIe1aad98_3321,RIe1a8a70_3296,RIe1a5d70_3264,RIe1a3070_3232,RIe1a0370_3200,RIe18c870_2976,RIe178d70_2752,RIe2266c8_4727,
        RIe21b2c8_4599,RIe204ac8_4343,RIe1feb28_4275,RIe1f7ee0_4198,RIe1f0a28_4115,RIe1d4f30_3800,RIe1bba30_3512,RIe1ae8a8_3363,RIe170ee0_2662,RIdec5270_707,
        RIdec2570_675,RIee1ff18_4822,RIdebf870_643,RIfe7f848_7795,RIdebcb70_611,RIdeb9e70_579,RIdeb7170_547,RIfe7fc80_7798,RIdeb1770_483,RIfca5d58_6909,
        RIdeaea70_451,RIfcaf808_7019,RIdeaa0d8_419,RIdea37d8_387,RIde9ced8_355,RIfcdc3d0_7528,RIfcce438_7369,RIfcb0a50_7032,RIfc75680_6358,RIde90d40_296,
        RIfe7f9b0_7796,RIde89720_260,RIde85580_240,RIde81728_221,RIfc52f40_5966,RIfc82100_6502,RIfca7108_6923,RIfe7fb18_7797,RIe16b648_2599,RIe169a28_2579,
        RIe167ca0_2558,RIe165270_2528,RIe162570_2496,RIee37258_5086,RIe15f870_2464,RIee36178_5074,RIe15cb70_2432,RIe157170_2368,RIe154470_2336,RIfc86fc0_6558,
        RIe151770_2304,RIfc4eff8_5921,RIe14ea70_2272,RIfce1290_7584,RIe14bd70_2240,RIe149070_2208,RIe146370_2176,RIee34558_5054,RIee331a8_5040,RIee320c8_5028,
        RIee31150_5017,RIfe800b8_7801,RIfe7ff50_7800,RIdf3caf0_2067,RIfe7fde8_7799,RIfcc8330_7300,RIee2f800_4999,RIfca0d30_6852,RIee2d640_4975,RIdf35638_1984,
        RIdf331a8_1958,RIdf31150_1935,RIdf2ef90_1911,RIee2bb88_4956,RIee2a0d0_4937,RIee28d20_4923,RIfe7f578_7793,RIdf2a238_1856,RIdf27f10_1831,RIfe7f6e0_7794,
        RIdf246d0_1791,RIfcce9d8_7373,RIfc63638_6153,RIdf22c18_1772,RIfc62990_6144,RIdf21700_1757,RIdf1f810_1735,RIfeaa958_8257,RIdf19168_1662,RIdf16e40_1637,
        RIdf14140_1605,RIdf11440_1573,RIdf0e740_1541,RIdf0ba40_1509,RIdf08d40_1477,RIdf06040_1445,RIdf03340_1413,RIdefd940_1349,RIdefac40_1317,RIdef7f40_1285,
        RIdef5240_1253,RIdef2540_1221,RIdeef840_1189,RIdeecb40_1157,RIdee9e40_1125,RIfcb7800_7110,RIee24838_4874,RIfc4cb68_5895,RIee23320_4859,RIfe80388_7803,
        RIdee2c58_1044,RIfe80220_7802,RIdedea40_997,RIfc98900_6758,RIee223a8_4848,RIfcc8600_7302,RIee212c8_4836,RIded9748_938,RIfe804f0_7804,RIded53c8_890,
        RIded2c68_862,RIded0670_835,RIdecd970_803,RIdecac70_771,RIdec7f70_739,RIdeb4470_515,RIde965d8_323,RIe16e078_2629,RIe159e70_2400,RIe143670_2144,
        RIdf38068_2014,RIdf2c6c8_1882,RIdf1cf48_1706,RIdf00640_1381,RIdee7140_1093,RIdedbea8_966,RIde7c520_196,RIe19d508_3167,RIe19a808_3135,RIfe7ee70_7788,
        RIe197b08_3103,RIfe7efd8_7789,RIe194e08_3071,RIe192108_3039,RIe18f408_3007,RIe189a08_2943,RIe186d08_2911,RIf143768_5227,RIe184008_2879,RIfc4bbf0_5884,
        RIe181308_2847,RIe17e608_2815,RIe17b908_2783,RIfe7f410_7792,RIf140d38_5197,RIe176fe8_2731,RIe175ad0_2716,RIfe7f2a8_7791,RIf13f118_5177,RIee3e440_5167,
        RIee3d360_5155,RIee3c280_5143,RIee3b1a0_5131,RIfe7f140_7790,RIe173640_2690,RIf170330_5736,RIf16f520_5726,RIf16e2d8_5713,RIf16d630_5704,RIfe7ea38_7785,
        RIe223860_4694,RIfc9c410_6800,RIe220b60_4662,RIfcb8340_7118,RIe21de60_4630,RIe218460_4566,RIe215760_4534,RIfc9cc80_6806,RIe212a60_4502,RIfc4ddb0_5908,
        RIe20fd60_4470,RIfc873f8_6561,RIe20d060_4438,RIe20a360_4406,RIe207660_4374,RIfc86750_6552,RIfc4e4b8_5913,RIe202368_4315,RIe200a18_4297,RIf165200_5610,
        RIf164558_5601,RIf163478_5589,RIf161f60_5574,RIf160070_5552,RIf15e180_5530,RIe1fcc38_4253,RIe1fb9f0_4240,RIf15cc68_5515,RIf15b750_5500,RIf15a670_5488,
        RIf159c98_5481,RIf158e88_5471,RIf157ad8_5457,RIf156e30_5448,RIfe7e768_7783,RIf1562f0_5440,RIf1557b0_5432,RIf154838_5421,RIfe7e8d0_7784,RIf1531b8_5405,
        RIfc52400_5958,RIf150a58_5377,RIe1f3188_4143,RIf14f978_5365,RIf14ecd0_5356,RIf14dec0_5346,RIe1ede90_4084,RIe1eb5c8_4055,RIe1e88c8_4023,RIe1e5bc8_3991,
        RIe1e2ec8_3959,RIe1e01c8_3927,RIe1dd4c8_3895,RIe1da7c8_3863,RIe1d7ac8_3831,RIe1d20c8_3767,RIe1cf3c8_3735,RIe1cc6c8_3703,RIe1c99c8_3671,RIe1c6cc8_3639,
        RIe1c3fc8_3607,RIe1c12c8_3575,RIe1be5c8_3543,RIf14c9a8_5331,RIf14b760_5318,RIfe7ed08_7787,RIfe7e600_7782,RIf14a518_5305,RIfca1f78_6865,RIfe7eba0_7786,
        RIfe7e498_7781,RIf148e98_5289,RIf147c50_5276,RIfe7e330_7780,RIe1b0a68_3387,RIf147278_5269,RIf1465d0_5260,RIe1ac418_3337,RIe1aac30_3320,RIe1a8908_3295,
        RIe1a5c08_3263,RIe1a2f08_3231,RIe1a0208_3199,RIe18c708_2975,RIe178c08_2751,RIe226560_4726,RIe21b160_4598,RIe204960_4342,RIe1fe9c0_4274,RIe1f7d78_4197,
        RIe1f08c0_4114,RIe1d4dc8_3799,RIe1bb8c8_3511,RIe1ae740_3362,RIe170d78_2661,RIdec56a8_710,RIdec29a8_678,RIfc54020_5978,RIdebfca8_646,RIee1f540_4815,
        RIdebcfa8_614,RIdeba2a8_582,RIdeb75a8_550,RIfc4fe08_5931,RIdeb1ba8_486,RIfc6b630_6244,RIdeaeea8_454,RIfc6a118_6229,RIdeaaab0_422,RIdea41b0_390,
        RIde9d8b0_358,RIfc69ce0_6226,RIee1be68_4776,RIfc653c0_6174,RIee1ac20_4763,RIde91718_299,RIde8df50_282,RIde89db0_262,RIde85c10_242,RIde81db8_223,
        RIfca76a8_6927,RIfcca4f0_7324,RIfc4ce38_5897,RIfc6b360_6242,RIe16b918_2601,RIe169cf8_2581,RIe167f70_2560,RIe1656a8_2531,RIe1629a8_2499,RIee37690_5089,
        RIe15fca8_2467,RIfce93f0_7676,RIe15cfa8_2435,RIe1575a8_2371,RIe1548a8_2339,RIee35908_5068,RIe151ba8_2307,RIee34f30_5061,RIe14eea8_2275,RIfce32e8_7607,
        RIe14c1a8_2243,RIe1494a8_2211,RIe1467a8_2179,RIfcde2c0_7550,RIfc687c8_6211,RIfca9160_6946,RIfcb1590_7040,RIe141078_2117,RIdf3ef80_2093,RIdf3cdc0_2069,
        RIfebeb60_8290,RIfc64448_6163,RIee2fad0_5001,RIfca7978_6929,RIfc676e8_6199,RIdf35a70_1987,RIdf335e0_1961,RIdf31420_1937,RIdf2f3c8_1914,RIfccef78_7377,
        RIfca6fa0_6922,RIfc62558_6141,RIfc61fb8_6137,RIfe81b70_7820,RIdf281e0_1833,RIfe81cd8_7821,RIdf249a0_1793,RIfc44300_5798,RIfcafc40_7022,RIdf22ee8_1774,
        RIfcaac18_6965,RIdf219d0_1759,RIdf1fae0_1737,RIdf1b1c0_1685,RIdf19438_1664,RIdf17278_1640,RIdf14578_1608,RIdf11878_1576,RIdf0eb78_1544,RIdf0be78_1512,
        RIdf09178_1480,RIdf06478_1448,RIdf03778_1416,RIdefdd78_1352,RIdefb078_1320,RIdef8378_1288,RIdef5678_1256,RIdef2978_1224,RIdeefc78_1192,RIdeecf78_1160,
        RIdeea278_1128,RIfc611a8_6127,RIfc61a18_6133,RIfca65c8_6915,RIfca6b68_6919,RIdee4b48_1066,RIdee2dc0_1045,RIdee0c00_1021,RIdedeba8_998,RIfc626c0_6142,
        RIfc738f8_6337,RIfcb31b0_7060,RIee21430_4837,RIded9a18_940,RIded7588_914,RIded5698_892,RIded30a0_865,RIded0aa8_838,RIdecdda8_806,RIdecb0a8_774,
        RIdec83a8_742,RIdeb48a8_518,RIde96fb0_326,RIe16e4b0_2632,RIe15a2a8_2403,RIe143aa8_2147,RIdf384a0_2017,RIdf2cb00_1885,RIdf1d380_1709,RIdf00a78_1384,
        RIdee7578_1096,RIdedc2e0_969,RIde7cef8_199,RIe19d940_3170,RIe19ac40_3138,RIfc64880_6166,RIe197f40_3106,RIf144848_5239,RIe195240_3074,RIe192540_3042,
        RIe18f840_3010,RIe189e40_2946,RIe187140_2914,RIf143a38_5229,RIe184440_2882,RIfc6f140_6286,RIe181740_2850,RIe17ea40_2818,RIe17bd40_2786,RIfc64f88_6171,
        RIf141008_5199,RIe177150_2732,RIfe81738_7817,RIfccabf8_7329,RIf13f3e8_5179,RIfca81e8_6935,RIee3d630_5157,RIfc66068_6183,RIfc6ed08_6283,RIfcdde88_7547,
        RIe173a78_2693,RIfc66338_6185,RIfc6eba0_6282,RIfc664a0_6186,RIfcacdd8_6989,RIfe81468_7815,RIe223c98_4697,RIfc66d10_6192,RIe220f98_4665,RIf16b038_5677,
        RIe21e298_4633,RIe218898_4569,RIe215b98_4537,RIfc3fc38_5751,RIe212e98_4505,RIfc67850_6200,RIe210198_4473,RIf167f00_5642,RIe20d498_4441,RIe20a798_4409,
        RIe207a98_4377,RIfcacb08_6987,RIfcac9a0_6986,RIfea8900_8234,RIfe818a0_7818,RIfca8a58_6941,RIfccad60_7330,RIfcac838_6985,RIfc67418_6197,RIf160340_5554,
        RIf15e450_5532,RIfe81a08_7819,RIfe81300_7814,RIfc6dac0_6270,RIf15ba20_5502,RIfc6d958_6269,RIfc6d7f0_6268,RIfc587d8_6029,RIfc6cf80_6262,RIfc6d3b8_6265,
        RIfe815d0_7816,RIfc6d520_6266,RIfcabe60_6978,RIfc6d0e8_6263,RIe1f5780_4170,RIfc6c5a8_6255,RIfc68d68_6215,RIfc68c00_6214,RIe1f3458_4145,RIfc68a98_6213,
        RIfccb8a0_7338,RIfca9b38_6953,RIe1ee160_4086,RIe1eba00_4058,RIe1e8d00_4026,RIe1e6000_3994,RIe1e3300_3962,RIe1e0600_3930,RIe1dd900_3898,RIe1dac00_3866,
        RIe1d7f00_3834,RIe1d2500_3770,RIe1cf800_3738,RIe1ccb00_3706,RIe1c9e00_3674,RIe1c7100_3642,RIe1c4400_3610,RIe1c1700_3578,RIe1bea00_3546,RIfc6bbd0_6248,
        RIfcdd348_7539,RIe1b9438_3485,RIe1b73e0_3462,RIfcab5f0_6972,RIfccbb70_7340,RIe1b5220_3438,RIe1b3e70_3424,RIfc6c9e0_6258,RIfcab488_6971,RIfea7dc0_8226,
        RIe1b0bd0_3388,RIfc6ce18_6261,RIfcabfc8_6979,RIe1ac580_3338,RIe1aaf00_3322,RIe1a8d40_3298,RIe1a6040_3266,RIe1a3340_3234,RIe1a0640_3202,RIe18cb40_2978,
        RIe179040_2754,RIe226998_4729,RIe21b598_4601,RIe204d98_4345,RIe1fedf8_4277,RIe1f81b0_4200,RIe1f0cf8_4117,RIe1d5200_3802,RIe1bbd00_3514,RIe1aeb78_3365,
        RIe1711b0_2664,RIdec5540_709,RIdec2840_677,RIfcc4dc0_7262,RIdebfb40_645,RIfc9d7c0_6814,RIdebce40_613,RIdeba140_581,RIdeb7440_549,RIfc4d978_5905,
        RIdeb1a40_485,RIfc9dbf8_6817,RIdeaed40_453,RIfcb8610_7120,RIdeaa768_421,RIdea3e68_389,RIde9d568_357,RIfc50678_5937,RIfc507e0_5938,RIfc9dec8_6819,
        RIfc853a0_6538,RIde913d0_298,RIde8dc08_281,RIde89a68_261,RIde858c8_241,RIde81a70_222,RIfc84860_6530,RIfc50948_5939,RIfc84c98_6533,RIfcb7da0_7114,
        RIe16b7b0_2600,RIe169b90_2580,RIe167e08_2559,RIe165540_2530,RIe162840_2498,RIee37528_5088,RIe15fb40_2466,RIfcb5be0_7090,RIe15ce40_2434,RIe157440_2370,
        RIe154740_2338,RIfcd35c8_7427,RIe151a40_2306,RIfc53a80_5974,RIe14ed40_2274,RIfcc6170_7276,RIe14c040_2242,RIe149340_2210,RIe146640_2178,RIfc7f130_6468,
        RIee33310_5041,RIfcb4f38_7081,RIfc47f78_5841,RIe140f10_2116,RIdf3ee18_2092,RIdf3cc58_2068,RIdf3a7c8_2042,RIfc7fc70_6476,RIfcd27b8_7417,RIfca1000_6854,
        RIfcc6b48_7283,RIdf35908_1986,RIdf33478_1960,RIfebe9f8_8289,RIdf2f260_1913,RIfcb7968_7111,RIee2a3a0_4939,RIfc51050_5944,RIfcd3fa0_7434,RIdf2a3a0_1857,
        RIdf28078_1832,RIfe81198_7813,RIdf24838_1792,RIfc84428_6527,RIfce7ed8_7661,RIdf22d80_1773,RIfc515f0_5948,RIdf21868_1758,RIdf1f978_1736,RIdf1b058_1684,
        RIdf192d0_1663,RIdf17110_1639,RIdf14410_1607,RIdf11710_1575,RIdf0ea10_1543,RIdf0bd10_1511,RIdf09010_1479,RIdf06310_1447,RIdf03610_1415,RIdefdc10_1351,
        RIdefaf10_1319,RIdef8210_1287,RIdef5510_1255,RIdef2810_1223,RIdeefb10_1191,RIdeece10_1159,RIdeea110_1127,RIfc7e1b8_6457,RIfca19d8_6861,RIfc7dab0_6452,
        RIfc7e488_6459,RIdee49e0_1065,RIfe80d60_7810,RIfeabba0_8270,RIfe80bf8_7809,RIfcb3750_7064,RIfce9f30_7684,RIfc7e5f0_6460,RIfc56a50_6008,RIfe81030_7812,
        RIded7420_913,RIfe80ec8_7811,RIded2f38_864,RIded0940_837,RIdecdc40_805,RIdecaf40_773,RIdec8240_741,RIdeb4740_517,RIde96c68_325,RIe16e348_2631,
        RIe15a140_2402,RIe143940_2146,RIdf38338_2016,RIdf2c998_1884,RIdf1d218_1708,RIdf00910_1383,RIdee7410_1095,RIdedc178_968,RIde7cbb0_198,RIe19d7d8_3169,
        RIe19aad8_3137,RIfcc2d68_7239,RIe197dd8_3105,RIfc5c5b8_6073,RIe1950d8_3073,RIe1923d8_3041,RIe18f6d8_3009,RIe189cd8_2945,RIe186fd8_2913,RIf1438d0_5228,
        RIe1842d8_2881,RIfc5b370_6060,RIe1815d8_2849,RIe17e8d8_2817,RIe17bbd8_2785,RIfcbb748_7155,RIfc59480_6038,RIfcbbce8_7159,RIe175c38_2717,RIfcdb890_7520,
        RIfc59b88_6043,RIfc8ada0_6602,RIfcb5eb0_7092,RIfc57c98_6021,RIfc57158_6013,RIfc58aa8_6031,RIe173910_2692,RIfcc62d8_7277,RIfc8a968_6599,RIfc57428_6015,
        RIfc56d20_6010,RIfc408e0_5760,RIe223b30_4696,RIfc82970_6508,RIe220e30_4664,RIfcecc30_7716,RIe21e130_4632,RIe218730_4568,RIe215a30_4536,RIfc3fad0_5750,
        RIe212d30_4504,RIf169148_5655,RIe210030_4472,RIfc545c0_5982,RIe20d330_4440,RIe20a630_4408,RIe207930_4376,RIfc88d48_6579,RIfc4bec0_5886,RIe202638_4317,
        RIe200b80_4298,RIfc88910_6576,RIfc4c190_5888,RIfc4c2f8_5889,RIfcba398_7141,RIfcd4270_7436,RIfcba0c8_7139,RIe1fcda0_4254,RIe1fbb58_4241,RIfc53d50_5976,
        RIfc9b768_6791,RIfc537b0_5972,RIfc4c5c8_5891,RIfc9e468_6823,RIf157da8_5459,RIfcb9f60_7138,RIe1fa208_4223,RIfc849c8_6531,RIfc529a0_5962,RIfc9f6b0_6836,
        RIe1f5618_4169,RIf153320_5406,RIfcc4988_7259,RIf150d28_5379,RIfebe458_8285,RIfc87f38_6569,RIfcb7f08_7115,RIf14e190_5348,RIfe80658_7805,RIe1eb898_4057,
        RIe1e8b98_4025,RIe1e5e98_3993,RIe1e3198_3961,RIe1e0498_3929,RIe1dd798_3897,RIe1daa98_3865,RIe1d7d98_3833,RIe1d2398_3769,RIe1cf698_3737,RIe1cc998_3705,
        RIe1c9c98_3673,RIe1c6f98_3641,RIe1c4298_3609,RIe1c1598_3577,RIe1be898_3545,RIf14cc78_5333,RIf14ba30_5320,RIe1b92d0_3484,RIe1b7278_3461,RIf14a7e8_5307,
        RIf149ca8_5299,RIfebe5c0_8286,RIfe807c0_7806,RIfc50510_5936,RIfce4f08_7627,RIfe80a90_7808,RIfebe890_8288,RIfc9cde8_6807,RIfc87560_6562,RIfe80928_7807,
        RIfebe728_8287,RIe1a8bd8_3297,RIe1a5ed8_3265,RIe1a31d8_3233,RIe1a04d8_3201,RIe18c9d8_2977,RIe178ed8_2753,RIe226830_4728,RIe21b430_4600,RIe204c30_4344,
        RIe1fec90_4276,RIe1f8048_4199,RIe1f0b90_4116,RIe1d5098_3801,RIe1bbb98_3513,RIe1aea10_3364,RIe171048_2663,RIdec5978_712,RIdec2c78_680,RIfc8aad0_6600,
        RIdebff78_648,RIfc8ac38_6601,RIdebd278_616,RIdeba578_584,RIdeb7878_552,RIfc40e80_5764,RIdeb1e78_488,RIfcdaeb8_7513,RIdeaf178_456,RIee1dbf0_4797,
        RIdeab140_424,RIdea4840_392,RIde9df40_360,RIfc8b070_6604,RIfcc38a8_7247,RIfc807b0_6484,RIfcbb8b0_7156,RIde91a60_300,RIde8e298_283,RIde8a440_264,
        RIde862a0_244,RIde82100_224,RIfcbbb80_7158,RIfc8c150_6616,RIfcbbfb8_7161,RIfc54458_5981,RIe16bbe8_2603,RIfc8c2b8_6617,RIe168240_2562,RIe165978_2533,
        RIe162c78_2501,RIee37960_5091,RIe15ff78_2469,RIfcd6b38_7465,RIe15d278_2437,RIe157878_2373,RIe154b78_2341,RIfc8e5e0_6642,RIe151e78_2309,RIfcb4290_7072,
        RIe14f178_2277,RIfc56ff0_6012,RIe14c478_2245,RIe149778_2213,RIe146a78_2181,RIee346c0_5055,RIee335e0_5043,RIee32398_5030,RIee31420_5019,RIe141348_2119,
        RIe13f020_2094,RIfec16f8_8321,RIdf3a930_2043,RIfce3e28_7615,RIfc56780_6006,RIfcb4128_7071,RIfce2eb0_7604,RIdf35d40_1989,RIfe88218_7893,RIdf316f0_1939,
        RIdf2f698_1916,RIfc7f9a0_6474,RIfce4260_7618,RIfcd62c8_7459,RIfce9990_7680,RIdf2a670_1859,RIdf284b0_1835,RIdf26728_1814,RIdf24c70_1795,RIfc7ecf8_6465,
        RIfcc31a0_7242,RIfc99008_6763,RIfc46e98_5829,RIfce2a78_7601,RIdf1fdb0_1739,RIfcc6e18_7285,RIdf19708_1666,RIdf17548_1642,RIdf14848_1610,RIdf11b48_1578,
        RIdf0ee48_1546,RIdf0c148_1514,RIdf09448_1482,RIdf06748_1450,RIdf03a48_1418,RIdefe048_1354,RIdefb348_1322,RIdef8648_1290,RIdef5948_1258,RIdef2c48_1226,
        RIdeeff48_1194,RIdeed248_1162,RIdeea548_1130,RIfcd9130_7492,RIfc7cb38_6441,RIfc97af0_6748,RIfcb3e58_7069,RIdee4e18_1068,RIdee3090_1047,RIdee0ed0_1023,
        RIfe88380_7894,RIfc97dc0_6750,RIfcc2930_7236,RIfcd9298_7493,RIfc7c868_6439,RIded9ce8_942,RIded76f0_915,RIded5968_894,RIded3370_867,RIded0d78_840,
        RIdece078_808,RIdecb378_776,RIdec8678_744,RIdeb4b78_520,RIde97640_328,RIe16e780_2634,RIe15a578_2405,RIe143d78_2149,RIdf38770_2019,RIdf2cdd0_1887,
        RIdf1d650_1711,RIdf00d48_1386,RIdee7848_1098,RIdedc5b0_971,RIde7d588_201,RIe19dc10_3172,RIe19af10_3140,RIfec1590_8320,RIe198210_3108,RIfec1428_8319,
        RIe195510_3076,RIe192810_3044,RIe18fb10_3012,RIe18a110_2948,RIe187410_2916,RIfec12c0_8318,RIe184710_2884,RIfc88370_6572,RIe181a10_2852,RIe17ed10_2820,
        RIe17c010_2788,RIfc6ccb0_6260,RIfc5f858_6109,RIfca88f0_6940,RIe175f08_2719,RIfc81020_6490,RIfcc6008_7275,RIfc4ea58_5917,RIfc42140_5774,RIfca3b98_6885,
        RIfc5ac68_6055,RIfc984c8_6755,RIe173d48_2695,RIfc9b330_6788,RIf16f688_5727,RIfc42410_5776,RIfc5f588_6107,RIfe880b0_7892,RIe223f68_4699,RIf16bfb0_5688,
        RIe221268_4667,RIfc86cf0_6556,RIe21e568_4635,RIe218b68_4571,RIe215e68_4539,RIfe87de0_7890,RIe213168_4507,RIf1692b0_5656,RIe210468_4475,RIfcdf670_7564,
        RIe20d768_4443,RIe20aa68_4411,RIe207d68_4379,RIfca6460_6914,RIf1662e0_5622,RIe202908_4319,RIfe87b10_7888,RIfc58c10_6032,RIfc50ab0_5940,RIfccd790_7360,
        RIfccd1f0_7356,RIf160610_5556,RIf15e720_5534,RIfe87c78_7889,RIfe87f48_7891,RIfce7668_7655,RIfc86480_6550,RIfcd2218_7413,RIfcb01e0_7026,RIfc47b40_5838,
        RIfc84158_6525,RIfc4b920_5882,RIe1fa4d8_4225,RIfc4ba88_5883,RIfcb7530_7108,RIfcd58f0_7452,RIe1f5a50_4172,RIf153488_5407,RIf151ca0_5390,RIfc51e60_5954,
        RIe1f3728_4147,RIfc9aef8_6785,RIfcbaaa0_7146,RIfc52130_5956,RIe1ee430_4088,RIe1ebcd0_4060,RIe1e8fd0_4028,RIe1e62d0_3996,RIe1e35d0_3964,RIe1e08d0_3932,
        RIe1ddbd0_3900,RIe1daed0_3868,RIe1d81d0_3836,RIe1d27d0_3772,RIe1cfad0_3740,RIe1ccdd0_3708,RIe1ca0d0_3676,RIe1c73d0_3644,RIe1c46d0_3612,RIe1c19d0_3580,
        RIe1becd0_3548,RIfce0b88_7579,RIfc82808_6507,RIe1b9708_3487,RIe1b76b0_3464,RIfcd5bc0_7454,RIfcb69f0_7100,RIe1b54f0_3440,RIe1b4140_3426,RIfc89f90_6592,
        RIfce9af8_7681,RIe1b2958_3409,RIe1b0ea0_3390,RIfc4a138_5865,RIfc8a260_6594,RIe1ac850_3340,RIe1ab1d0_3324,RIe1a9010_3300,RIe1a6310_3268,RIe1a3610_3236,
        RIe1a0910_3204,RIe18ce10_2980,RIe179310_2756,RIe226c68_4731,RIe21b868_4603,RIe205068_4347,RIe1ff0c8_4279,RIe1f8480_4202,RIe1f0fc8_4119,RIe1d54d0_3804,
        RIe1bbfd0_3516,RIe1aee48_3367,RIe171480_2666,RIdec5810_711,RIdec2b10_679,RIfce6f60_7650,RIdebfe10_647,RIfc95228_6719,RIdebd110_615,RIdeba410_583,
        RIdeb7710_551,RIfe879a8_7887,RIdeb1d10_487,RIfcc16e8_7223,RIdeaf010_455,RIfca4f48_6899,RIdeaadf8_423,RIdea44f8_391,RIde9dbf8_359,RIee1cf48_4788,
        RIee1bfd0_4777,RIfc95660_6722,RIfcee148_7731,RIfe87840_7886,RIfe876d8_7885,RIde8a0f8_263,RIde85f58_243,RIfcb0780_7030,RIfcee9b8_7737,RIfc5f150_6104,
        RIfcdee00_7558,RIfcd8050_7480,RIe16ba80_2602,RIfca5380_6902,RIe1680d8_2561,RIe165810_2532,RIe162b10_2500,RIee377f8_5090,RIe15fe10_2468,RIee36448_5076,
        RIe15d110_2436,RIe157710_2372,RIe154a10_2340,RIfc3f3c8_5745,RIe151d10_2308,RIfcde9c8_7555,RIe14f010_2276,RIfc4a2a0_5866,RIe14c310_2244,RIe149610_2212,
        RIe146910_2180,RIfc62288_6139,RIee33478_5042,RIfc71b70_6316,RIee312b8_5018,RIe1411e0_2118,RIfe87570_7884,RIdf3cf28_2070,RIfe87408_7883,RIfcc99b0_7316,
        RIfccf0e0_7378,RIfcaeb60_7010,RIfcca220_7322,RIdf35bd8_1988,RIdf33748_1962,RIdf31588_1938,RIdf2f530_1915,RIee2be58_4958,RIee2a508_4940,RIee28ff0_4925,
        RIee27da8_4912,RIdf2a508_1858,RIdf28348_1834,RIdf265c0_1813,RIdf24b08_1794,RIfc74708_6347,RIfc42578_5777,RIfc43388_5787,RIfc745a0_6346,RIfcb0078_7025,
        RIdf1fc48_1738,RIfcaff10_7024,RIdf195a0_1665,RIdf173e0_1641,RIdf146e0_1609,RIdf119e0_1577,RIdf0ece0_1545,RIdf0bfe0_1513,RIdf092e0_1481,RIdf065e0_1449,
        RIdf038e0_1417,RIdefdee0_1353,RIdefb1e0_1321,RIdef84e0_1289,RIdef57e0_1257,RIdef2ae0_1225,RIdeefde0_1193,RIdeed0e0_1161,RIdeea3e0_1129,RIee257b0_4885,
        RIfca73d8_6925,RIee23e60_4867,RIfce66f0_7644,RIdee4cb0_1067,RIdee2f28_1046,RIdee0d68_1022,RIdeded10_999,RIfcca388_7323,RIfce6858_7645,RIfcceca8_7375,
        RIfcdc970_7532,RIded9b80_941,RIfeaaac0_8258,RIded5800_893,RIded3208_866,RIded0c10_839,RIdecdf10_807,RIdecb210_775,RIdec8510_743,RIdeb4a10_519,
        RIde972f8_327,RIe16e618_2633,RIe15a410_2404,RIe143c10_2148,RIdf38608_2018,RIdf2cc68_1886,RIdf1d4e8_1710,RIdf00be0_1385,RIdee76e0_1097,RIdedc448_970,
        RIde7d240_200,RIe19daa8_3171,RIe19ada8_3139,RIf1457c0_5250,RIe1980a8_3107,RIf1449b0_5240,RIe1953a8_3075,RIe1926a8_3043,RIe18f9a8_3011,RIe189fa8_2947,
        RIe1872a8_2915,RIf143ba0_5230,RIe1845a8_2883,RIfc912e0_6674,RIe1818a8_2851,RIe17eba8_2819,RIe17bea8_2787,RIfc915b0_6676,RIfcbe5b0_7188,RIfce3b58_7613,
        RIe175da0_2718,RIfceb448_7699,RIfcc7958_7293,RIfc42de8_5783,RIfc96e48_6739,RIfc7a810_6416,RIfc96ce0_6738,RIfcc7ac0_7294,RIe173be0_2694,RIfce39f0_7612,
        RIfc7a540_6414,RIfc91b50_6680,RIfc429b0_5780,RIfea9710_8244,RIe223e00_4698,RIfcd8488_7483,RIe221100_4666,RIfc920f0_6684,RIe21e400_4634,RIe218a00_4570,
        RIe215d00_4538,RIfc79e38_6409,RIe213000_4506,RIfcbee20_7194,RIe210300_4474,RIf168068_5643,RIe20d600_4442,RIe20a900_4410,RIe207c00_4378,RIfc5af38_6057,
        RIfcd73a8_7471,RIe2027a0_4318,RIe200ce8_4299,RIfcb2670_7052,RIfcdf940_7566,RIfc5b208_6059,RIfcbf3c0_7198,RIf1604a8_5555,RIf15e5b8_5533,RIfe872a0_7882,
        RIfe87138_7881,RIfc78920_6394,RIfec1158_8317,RIfc93338_6697,RIfcea368_7687,RIfcb23a0_7050,RIfc5bbe0_6066,RIfcede78_7729,RIe1fa370_4224,RIfcd4c48_7443,
        RIfce1dd0_7592,RIfcbf960_7202,RIe1f58e8_4171,RIfcbfc30_7204,RIfc78380_6390,RIfc93770_6700,RIe1f35c0_4146,RIfcb1f68_7047,RIfce1b00_7590,RIfc93a40_6702,
        RIe1ee2c8_4087,RIe1ebb68_4059,RIe1e8e68_4027,RIe1e6168_3995,RIe1e3468_3963,RIe1e0768_3931,RIe1dda68_3899,RIe1dad68_3867,RIe1d8068_3835,RIe1d2668_3771,
        RIe1cf968_3739,RIe1ccc68_3707,RIe1c9f68_3675,RIe1c7268_3643,RIe1c4568_3611,RIe1c1868_3579,RIe1beb68_3547,RIfcdec98_7557,RIfc94148_6707,RIe1b95a0_3486,
        RIe1b7548_3463,RIfcd12a0_7402,RIfceabd8_7693,RIe1b5388_3439,RIe1b3fd8_3425,RIfc94850_6712,RIfcd7c18_7477,RIe1b27f0_3408,RIe1b0d38_3389,RIfc76a30_6372,
        RIfce2640_7598,RIe1ac6e8_3339,RIe1ab068_3323,RIe1a8ea8_3299,RIe1a61a8_3267,RIe1a34a8_3235,RIe1a07a8_3203,RIe18cca8_2979,RIe1791a8_2755,RIe226b00_4730,
        RIe21b700_4602,RIe204f00_4346,RIe1fef60_4278,RIe1f8318_4201,RIe1f0e60_4118,RIe1d5368_3803,RIe1bbe68_3515,RIe1aece0_3366,RIe171318_2665,RIdec5c48_714,
        RIdec2f48_682,RIfc7c160_6434,RIdec0248_650,RIfcb38b8_7065,RIdebd548_618,RIdeba848_586,RIdeb7b48_554,RIfce7c08_7659,RIdeb2148_490,RIfce7aa0_7658,
        RIdeaf448_458,RIfca38c8_6883,RIdeab7d0_426,RIdea4ed0_394,RIde9e5d0_362,RIfc41e70_5772,RIfc5b0a0_6058,RIfcdbb60_7522,RIfc78650_6392,RIfea92d8_8241,
        RIde8e5e0_284,RIfea0d40_8174,RIfea0bd8_8173,RIfcdf508_7563,RIfcb1b30_7044,RIfc5ccc0_6078,RIfcb16f8_7041,RIfc77b10_6384,RIe16beb8_2605,RIe169e60_2582,
        RIe168510_2564,RIe165c48_2535,RIe162f48_2503,RIfc4f9d0_5928,RIe160248_2471,RIfc4e8f0_5916,RIe15d548_2439,RIe157b48_2375,RIe154e48_2343,RIfc4e1e8_5911,
        RIe152148_2311,RIfc868b8_6553,RIe14f448_2279,RIfc865e8_6551,RIe14c748_2247,RIe149a48_2215,RIe146d48_2183,RIfc9eb70_6828,RIfc9ecd8_6829,RIfcc5630_7268,
        RIfc83bb8_6521,RIe141618_2121,RIfea0ea8_8175,RIdf3d1f8_2072,RIdf3ac00_2045,RIee308e0_5011,RIfcd3cd0_7432,RIfc84e00_6534,RIfc834b0_6516,RIdf36010_1991,
        RIdf33a18_1964,RIdf31858_1940,RIdf2f968_1918,RIee2c128_4960,RIee2a7d8_4942,RIee292c0_4927,RIee28078_4914,RIdf2a940_1861,RIdf28780_1837,RIfea0a70_8172,
        RIfea0908_8171,RIfcd4f18_7445,RIfca0628_6847,RIdf23050_1775,RIfcd3190_7424,RIdf21b38_1760,RIdf20080_1741,RIdf1b328_1686,RIdf199d8_1668,RIdf17818_1644,
        RIdf14b18_1612,RIdf11e18_1580,RIdf0f118_1548,RIdf0c418_1516,RIdf09718_1484,RIdf06a18_1452,RIdf03d18_1420,RIdefe318_1356,RIdefb618_1324,RIdef8918_1292,
        RIdef5c18_1260,RIdef2f18_1228,RIdef0218_1196,RIdeed518_1164,RIdeea818_1132,RIfcdf3a0_7562,RIfca5218_6901,RIfcdc538_7529,RIfcdc6a0_7530,RIdee50e8_1070,
        RIdee3360_1049,RIfea07a0_8170,RIdedefe0_1001,RIfcb0d20_7034,RIfcd4978_7441,RIfca49a8_6895,RIfca1708_6859,RIded9fb8_944,RIded79c0_917,RIded5ad0_895,
        RIfeab498_8265,RIded1048_842,RIdece348_810,RIdecb648_778,RIdec8948_746,RIdeb4e48_522,RIde97cd0_330,RIe16ea50_2636,RIe15a848_2407,RIe144048_2151,
        RIdf38a40_2021,RIdf2d0a0_1889,RIdf1d920_1713,RIdf01018_1388,RIdee7b18_1100,RIdedc880_973,RIde7dc18_203,RIe19dee0_3174,RIe19b1e0_3142,RIfc67580_6198,
        RIe1984e0_3110,RIfccb030_7332,RIe1957e0_3078,RIe192ae0_3046,RIe18fde0_3014,RIe18a3e0_2950,RIe1876e0_2918,RIfc6a550_6232,RIe1849e0_2886,RIfcaa7e0_6962,
        RIe181ce0_2854,RIe17efe0_2822,RIe17c2e0_2790,RIfc65d98_6181,RIfc65690_6176,RIe1772b8_2733,RIfea0638_8169,RIfcca928_7327,RIfc607d0_6120,RIfc65258_6173,
        RIee3d798_5158,RIee3c3e8_5144,RIfca9430_6948,RIee39f58_5118,RIe174018_2697,RIfcecf00_7718,RIfc650f0_6172,RIf16e5a8_5715,RIfc43a90_5792,RIfc65528_6175,
        RIe224238_4701,RIfca9f70_6956,RIe221538_4669,RIfc6b4c8_6243,RIe21e838_4637,RIe218e38_4573,RIe216138_4541,RIfc3fda0_5752,RIe213438_4509,RIfc61310_6128,
        RIe210738_4477,RIfc60c08_6123,RIe20da38_4445,RIe20ad38_4413,RIe208038_4381,RIfc66ba8_6191,RIfccbcd8_7341,RIe202bd8_4321,RIe200fb8_4301,RIfcadbe8_6999,
        RIfccbe40_7342,RIfca7540_6926,RIfc6a3e8_6231,RIfca6898_6917,RIfc73358_6333,RIe1fd070_4256,RIe1fbe28_4243,RIfcc2660_7234,RIfc44468_5799,RIf15a940_5490,
        RIfca7270_6924,RIfc5e070_6092,RIfc5dda0_6090,RIfc7e050_6456,RIe1fa7a8_4227,RIfc5d968_6087,RIfcd9568_7495,RIfc8d668_6631,RIe1f5d20_4174,RIfca4138_6889,
        RIfc8cdf8_6625,RIfcc7c28_7295,RIe1f39f8_4149,RIfc99440_6766,RIfcbc3f0_7164,RIfc5a128_6047,RIe1ee700_4090,RIe1ebfa0_4062,RIe1e92a0_4030,RIe1e65a0_3998,
        RIe1e38a0_3966,RIe1e0ba0_3934,RIe1ddea0_3902,RIe1db1a0_3870,RIe1d84a0_3838,RIe1d2aa0_3774,RIe1cfda0_3742,RIe1cd0a0_3710,RIe1ca3a0_3678,RIe1c76a0_3646,
        RIe1c49a0_3614,RIe1c1ca0_3582,RIe1befa0_3550,RIf14cde0_5334,RIf14bb98_5321,RIe1b99d8_3489,RIe1b7980_3466,RIfc4c460_5890,RIfc9e738_6825,RIe1b5658_3441,
        RIfec54d8_8365,RIf149168_5291,RIf147f20_5278,RIe1b2ac0_3410,RIe1b1170_3392,RIf1473e0_5270,RIf1468a0_5262,RIe1acb20_3342,RIe1ab338_3325,RIe1a92e0_3302,
        RIe1a65e0_3270,RIe1a38e0_3238,RIe1a0be0_3206,RIe18d0e0_2982,RIe1795e0_2758,RIe226f38_4733,RIe21bb38_4605,RIe205338_4349,RIe1ff398_4281,RIe1f8750_4204,
        RIe1f1298_4121,RIe1d57a0_3806,RIe1bc2a0_3518,RIe1af118_3369,RIe171750_2668,RIdec5ae0_713,RIdec2de0_681,RIfc82268_6503,RIdec00e0_649,RIfcb8d18_7125,
        RIdebd3e0_617,RIdeba6e0_585,RIdeb79e0_553,RIfcb9858_7133,RIdeb1fe0_489,RIfc9efa8_6831,RIdeaf2e0_457,RIfce0750_7576,RIdeab488_425,RIdea4b88_393,
        RIde9e288_361,RIee1d0b0_4789,RIee1c138_4778,RIfcd0e68_7399,RIfc76d00_6374,RIfe89028_7903,RIfe88d58_7901,RIfe88ec0_7902,RIfe88bf0_7900,RIfcda7b0_7508,
        RIfc4d810_5904,RIfc52dd8_5965,RIfcde590_7552,RIfc4f868_5927,RIe16bd50_2604,RIfc68930_6212,RIe1683a8_2563,RIe165ae0_2534,RIe162de0_2502,RIfe88a88_7899,
        RIe1600e0_2470,RIfcc9140_7310,RIe15d3e0_2438,RIe1579e0_2374,RIe154ce0_2342,RIfc698a8_6223,RIe151fe0_2310,RIee35098_5062,RIe14f2e0_2278,RIfcc0338_7209,
        RIe14c5e0_2246,RIe1498e0_2214,RIe146be0_2182,RIfc88208_6571,RIfc85670_6540,RIfc81f98_6501,RIfcc4f28_7263,RIe1414b0_2120,RIe13f188_2095,RIdf3d090_2071,
        RIdf3aa98_2044,RIfcd2920_7418,RIfc7d7e0_6450,RIfc49760_5858,RIfce5a48_7635,RIdf35ea8_1990,RIdf338b0_1963,RIfe88920_7898,RIdf2f800_1917,RIee2bfc0_4959,
        RIee2a670_4941,RIee29158_4926,RIee27f10_4913,RIdf2a7d8_1860,RIdf28618_1836,RIdf26890_1815,RIdf24dd8_1796,RIfcad918_6997,RIfc69fb0_6228,RIfc63368_6151,
        RIfc623f0_6140,RIfc60938_6121,RIdf1ff18_1740,RIfcba500_7142,RIdf19870_1667,RIdf176b0_1643,RIdf149b0_1611,RIdf11cb0_1579,RIdf0efb0_1547,RIdf0c2b0_1515,
        RIdf095b0_1483,RIdf068b0_1451,RIdf03bb0_1419,RIdefe1b0_1355,RIdefb4b0_1323,RIdef87b0_1291,RIdef5ab0_1259,RIdef2db0_1227,RIdef00b0_1195,RIdeed3b0_1163,
        RIdeea6b0_1131,RIfcc9848_7315,RIfc69a10_6224,RIfcacc70_6988,RIfccbfa8_7343,RIdee4f80_1069,RIdee31f8_1048,RIdee1038_1024,RIdedee78_1000,RIfc84590_6528,
        RIfc9bba0_6794,RIee21b38_4842,RIfc47168_5831,RIded9e50_943,RIded7858_916,RIfe887b8_7897,RIded34d8_868,RIded0ee0_841,RIdece1e0_809,RIdecb4e0_777,
        RIdec87e0_745,RIdeb4ce0_521,RIde97988_329,RIe16e8e8_2635,RIe15a6e0_2406,RIe143ee0_2150,RIdf388d8_2020,RIdf2cf38_1888,RIdf1d7b8_1712,RIdf00eb0_1387,
        RIdee79b0_1099,RIdedc718_972,RIde7d8d0_202,RIe19dd78_3173,RIe19b078_3141,RIfca1438_6857,RIe198378_3109,RIfca35f8_6881,RIe195678_3077,RIe192978_3045,
        RIe18fc78_3013,RIe18a278_2949,RIe187578_2917,RIfcba230_7140,RIe184878_2885,RIf142d90_5220,RIe181b78_2853,RIe17ee78_2821,RIe17c178_2789,RIfc9be70_6796,
        RIfc9bd08_6795,RIfc4ccd0_5896,RIe176070_2720,RIfc87c68_6567,RIfc87b00_6566,RIfcc4c58_7261,RIfc4fca0_5930,RIfc4f598_5925,RIfc876c8_6563,RIfc4dae0_5906,
        RIe173eb0_2696,RIfcb9420_7130,RIfc4e080_5910,RIfc4e350_5912,RIfc9d388_6811,RIfc40a48_5761,RIe2240d0_4700,RIfc85508_6539,RIe2213d0_4668,RIfc9ba38_6793,
        RIe21e6d0_4636,RIe218cd0_4572,RIe215fd0_4540,RIfc52c70_5964,RIe2132d0_4508,RIfca3760_6882,RIe2105d0_4476,RIfc97988_6747,RIe20d8d0_4444,RIe20abd0_4412,
        RIe207ed0_4380,RIfceb5b0_7700,RIfcddbb8_7545,RIe202a70_4320,RIe200e50_4300,RIfc73d30_6340,RIfcaf100_7014,RIfc71468_6311,RIfcdcad8_7533,RIfcdda50_7544,
        RIfca8620_6938,RIe1fcf08_4255,RIe1fbcc0_4242,RIfc6c008_6251,RIfcdd1e0_7538,RIfca9700_6950,RIfca92c8_6947,RIfcce5a0_7370,RIfc6ba68_6247,RIfc6f410_6288,
        RIe1fa640_4226,RIfcce000_7366,RIfc53918_5973,RIfcce708_7371,RIe1f5bb8_4173,RIf1535f0_5408,RIf151e08_5391,RIfc72db8_6329,RIe1f3890_4148,RIf14fc48_5367,
        RIfc72c50_6328,RIfc73e98_6341,RIe1ee598_4089,RIe1ebe38_4061,RIe1e9138_4029,RIe1e6438_3997,RIe1e3738_3965,RIe1e0a38_3933,RIe1ddd38_3901,RIe1db038_3869,
        RIe1d8338_3837,RIe1d2938_3773,RIe1cfc38_3741,RIe1ccf38_3709,RIe1ca238_3677,RIe1c7538_3645,RIe1c4838_3613,RIe1c1b38_3581,RIe1bee38_3549,RIfcb8a48_7123,
        RIfcb84a8_7119,RIe1b9870_3488,RIe1b7818_3465,RIfc85940_6542,RIfc9e198_6821,RIfeac140_8274,RIe1b42a8_3427,RIfc518c0_5950,RIfc838e8_6519,RIfe884e8_7895,
        RIe1b1008_3391,RIfcc5900_7270,RIfc82ad8_6509,RIe1ac9b8_3341,RIfe88650_7896,RIe1a9178_3301,RIe1a6478_3269,RIe1a3778_3237,RIe1a0a78_3205,RIe18cf78_2981,
        RIe179478_2757,RIe226dd0_4732,RIe21b9d0_4604,RIe2051d0_4348,RIe1ff230_4280,RIe1f85e8_4203,RIe1f1130_4120,RIe1d5638_3805,RIe1bc138_3517,RIe1aefb0_3368,
        RIe1715e8_2667,RIdec5f18_716,RIdec3218_684,RIee20350_4825,RIdec0518_652,RIee1f6a8_4816,RIdebd818_620,RIdebab18_588,RIdeb7e18_556,RIfce4da0_7626,
        RIdeb2418_492,RIfcea908_7691,RIdeaf718_460,RIfce20a0_7594,RIdeabe60_428,RIdea5560_396,RIde9ec60_364,RIfce6420_7642,RIee1c2a0_4779,RIfc75950_6360,
        RIee1ad88_4764,RIde920f0_302,RIfea4148_8211,RIfeaa688_8255,RIfea3fe0_8210,RIde82790_226,RIfc6f848_6291,RIfc5dc38_6089,RIfc76b98_6373,RIfcae2f0_7004,
        RIe16c020_2606,RIe16a130_2584,RIe1687e0_2566,RIe165f18_2537,RIe163218_2505,RIfcadd50_7000,RIe160518_2473,RIfc55268_5991,RIe15d818_2441,RIe157e18_2377,
        RIe155118_2345,RIfc45548_5811,RIe152418_2313,RIfc498c8_5859,RIe14f718_2281,RIfcbda70_7180,RIe14ca18_2249,RIe149d18_2217,RIe147018_2185,RIee34828_5056,
        RIee33748_5044,RIee32668_5032,RIee31588_5020,RIe1418e8_2123,RIe13f458_2097,RIdf3d360_2073,RIdf3aed0_2047,RIfc526d0_5960,RIfc42848_5779,RIfcae9f8_7009,
        RIfcb7260_7106,RIfea42b0_8212,RIdf33ce8_1966,RIdf31b28_1942,RIdf2fc38_1920,RIee2c3f8_4962,RIfc4cfa0_5898,RIfc572c0_6014,RIfc4f430_5924,RIfea3e78_8209,
        RIdf28a50_1839,RIdf26b60_1817,RIdf250a8_1798,RIfc9b600_6790,RIfcb9df8_7137,RIdf23320_1777,RIfc86318_6549,RIfeabfd8_8273,RIdf201e8_1742,RIdf1b5f8_1688,
        RIdf19ca8_1670,RIdf17ae8_1646,RIdf14de8_1614,RIdf120e8_1582,RIdf0f3e8_1550,RIdf0c6e8_1518,RIdf099e8_1486,RIdf06ce8_1454,RIdf03fe8_1422,RIdefe5e8_1358,
        RIdefb8e8_1326,RIdef8be8_1294,RIdef5ee8_1262,RIdef31e8_1230,RIdef04e8_1198,RIdeed7e8_1166,RIdeeaae8_1134,RIfc89018_6581,RIfcc54c8_7267,RIfc89180_6582,
        RIfc4b380_5878,RIdee53b8_1072,RIdee34c8_1050,RIfea3d10_8208,RIdedf148_1002,RIfcae188_7003,RIfc4b0b0_5876,RIfc74870_6348,RIfce4968_7623,RIdeda288_946,
        RIded7c90_919,RIded5da0_897,RIded3640_869,RIded1318_844,RIdece618_812,RIdecb918_780,RIdec8c18_748,RIdeb5118_524,RIde98360_332,RIe16ed20_2638,
        RIe15ab18_2409,RIe144318_2153,RIdf38d10_2023,RIdf2d370_1891,RIdf1dbf0_1715,RIdf012e8_1390,RIdee7de8_1102,RIdedcb50_975,RIde7e2a8_205,RIe19e1b0_3176,
        RIe19b4b0_3144,RIfc9cf50_6808,RIe1987b0_3112,RIfc87290_6560,RIe195ab0_3080,RIe192db0_3048,RIe1900b0_3016,RIe18a6b0_2952,RIe1879b0_2920,RIfc842c0_6526,
        RIe184cb0_2888,RIfc83a50_6520,RIe181fb0_2856,RIe17f2b0_2824,RIe17c5b0_2792,RIfc9d0b8_6809,RIfc9e030_6820,RIe177420_2734,RIe176340_2722,RIfc4f700_5926,
        RIfcc4820_7258,RIfc4fb38_5929,RIfce8040_7662,RIee3c6b8_5146,RIee3b308_5132,RIfc812f0_6492,RIe174180_2698,RIfcd3028_7423,RIfc7f400_6470,RIfc46a60_5826,
        RIfc472d0_5832,RIf16cc58_5697,RIe224508_4703,RIfc7d3a8_6447,RIe221808_4671,RIfc97c58_6749,RIe21eb08_4639,RIe219108_4575,RIe216408_4543,RIfcdbe30_7524,
        RIe213708_4511,RIf169580_5658,RIe210a08_4479,RIfca4570_6892,RIe20dd08_4447,RIe20b008_4415,RIe208308_4383,RIfc7b080_6422,RIfc59cf0_6044,RIfea9b48_8247,
        RIfea4418_8213,RIfc79cd0_6408,RIfcd19a8_7407,RIfcc81c8_7299,RIf162230_5576,RIf160778_5557,RIf15e888_5535,RIfea4580_8214,RIfea46e8_8215,RIfc77f48_6387,
        RIfc41fd8_5773,RIf15aaa8_5491,RIfc7c430_6436,RIf159158_5473,RIf157f10_5460,RIfcae890_7008,RIe1faa78_4229,RIfc4a840_5870,RIfc4ed28_5919,RIfce0e58_7581,
        RIe1f5ff0_4176,RIf153758_5409,RIf151f70_5392,RIfccb468_7335,RIe1f3cc8_4151,RIfc68ed0_6216,RIfc6d250_6264,RIfca9ca0_6954,RIe1ee9d0_4092,RIe1ec270_4064,
        RIe1e9570_4032,RIe1e6870_4000,RIe1e3b70_3968,RIe1e0e70_3936,RIe1de170_3904,RIe1db470_3872,RIe1d8770_3840,RIe1d2d70_3776,RIe1d0070_3744,RIe1cd370_3712,
        RIe1ca670_3680,RIe1c7970_3648,RIe1c4c70_3616,RIe1c1f70_3584,RIe1bf270_3552,RIfc784e8_6391,RIfcbef88_7195,RIe1b9ca8_3491,RIe1b7ae8_3467,RIfcc20c0_7230,
        RIfca6190_6912,RIe1b5928_3443,RIe1b4410_3428,RIfcb81d8_7117,RIfcc5090_7264,RIe1b2d90_3412,RIe1b1440_3394,RIfcd5350_7448,RIfcb9588_7131,RIe1acc88_3343,
        RIe1ab4a0_3326,RIe1a95b0_3304,RIe1a68b0_3272,RIe1a3bb0_3240,RIe1a0eb0_3208,RIe18d3b0_2984,RIe1798b0_2760,RIe227208_4735,RIe21be08_4607,RIe205608_4351,
        RIe1ff668_4283,RIe1f8a20_4206,RIe1f1568_4123,RIe1d5a70_3808,RIe1bc570_3520,RIe1af3e8_3371,RIe171a20_2670,RIdec5db0_715,RIdec30b0_683,RIee201e8_4824,
        RIdec03b0_651,RIfcaf538_7017,RIdebd6b0_619,RIdeba9b0_587,RIdeb7cb0_555,RIfc40fe8_5765,RIdeb22b0_491,RIfcd08c8_7395,RIdeaf5b0_459,RIee1dd58_4798,
        RIdeabb18_427,RIdea5218_395,RIde9e918_363,RIee1d218_4790,RIfcedd10_7728,RIfce62b8_7641,RIfcc92a8_7311,RIde91da8_301,RIde8e928_285,RIde8a788_265,
        RIde865e8_245,RIde82448_225,RIfea1448_8179,RIfc750e0_6354,RIfcc19b8_7225,RIfced8d8_7725,RIfec5eb0_8372,RIe169fc8_2583,RIe168678_2565,RIe165db0_2536,
        RIe1630b0_2504,RIfccfc20_7386,RIe1603b0_2472,RIee365b0_5077,RIe15d6b0_2440,RIe157cb0_2376,RIe154fb0_2344,RIfea1718_8181,RIe1522b0_2312,RIee35200_5063,
        RIe14f5b0_2280,RIfcb0348_7027,RIe14c8b0_2248,RIe149bb0_2216,RIe146eb0_2184,RIfc73790_6336,RIfcdf238_7561,RIee32500_5031,RIfc94f58_6717,RIe141780_2122,
        RIe13f2f0_2096,RIfec5be0_8370,RIdf3ad68_2046,RIfea15b0_8180,RIfc5fb28_6111,RIfcae728_7007,RIfc74438_6345,RIdf36178_1992,RIdf33b80_1965,RIdf319c0_1941,
        RIdf2fad0_1919,RIee2c290_4961,RIee2a940_4943,RIfc70658_6301,RIfc704f0_6300,RIdf2aaa8_1862,RIdf288e8_1838,RIdf269f8_1816,RIdf24f40_1797,RIfc64b50_6168,
        RIfccaa90_7328,RIdf231b8_1776,RIfcad4e0_6994,RIdf21ca0_1761,RIfeaad90_8260,RIdf1b490_1687,RIdf19b40_1669,RIdf17980_1645,RIdf14c80_1613,RIdf11f80_1581,
        RIdf0f280_1549,RIdf0c580_1517,RIdf09880_1485,RIdf06b80_1453,RIdf03e80_1421,RIdefe480_1357,RIdefb780_1325,RIdef8a80_1293,RIdef5d80_1261,RIdef3080_1229,
        RIdef0380_1197,RIdeed680_1165,RIdeea980_1133,RIfc595e8_6039,RIfcac568_6983,RIfcccf20_7354,RIfccd358_7357,RIdee5250_1071,RIfea7f28_8227,RIdee11a0_1025,
        RIfea12e0_8178,RIfc679b8_6201,RIee22510_4849,RIfc6dd90_6272,RIfc6cb48_6259,RIdeda120_945,RIded7b28_918,RIded5c38_896,RIfec5d48_8371,RIded11b0_843,
        RIdece4b0_811,RIdecb7b0_779,RIdec8ab0_747,RIdeb4fb0_523,RIde98018_331,RIe16ebb8_2637,RIe15a9b0_2408,RIe1441b0_2152,RIdf38ba8_2022,RIdf2d208_1890,
        RIdf1da88_1714,RIdf01180_1389,RIdee7c80_1101,RIdedc9e8_974,RIde7df60_204,RIe19e048_3175,RIe19b348_3143,RIfcc3ce0_7250,RIe198648_3111,RIfc7efc8_6467,
        RIe195948_3079,RIe192c48_3047,RIe18ff48_3015,RIe18a548_2951,RIe187848_2919,RIfc46790_5824,RIe184b48_2887,RIfc98d38_6761,RIe181e48_2855,RIe17f148_2823,
        RIe17c448_2791,RIfcb5d48_7091,RIfc995a8_6767,RIfc9a3b8_6777,RIe1761d8_2721,RIfc54188_5979,RIfcd2bf0_7420,RIfc8b778_6609,RIfc7dee8_6455,RIee3c550_5145,
        RIfc8c420_6618,RIee3a0c0_5119,RIfeaba38_8269,RIfc46628_5823,RIfcbc288_7163,RIf16e710_5716,RIfc8fdc8_6659,RIfc48c20_5850,RIe2243a0_4702,RIfca0358_6845,
        RIe2216a0_4670,RIfc9a688_6779,RIe21e9a0_4638,RIe218fa0_4574,RIe2162a0_4542,RIfc456b0_5812,RIe2135a0_4510,RIf169418_5657,RIe2108a0_4478,RIfc8bfe8_6615,
        RIe20dba0_4446,RIe20aea0_4414,RIe2081a0_4382,RIfc8c9c0_6622,RIfc7f568_6471,RIe202d40_4322,RIe201120_4302,RIfce2910_7600,RIfc487e8_5847,RIfc46d30_5828,
        RIfc992d8_6765,RIfca2680_6870,RIfc44a08_5803,RIe1fd1d8_4257,RIe1fbf90_4244,RIfc580d0_6024,RIfcbdbd8_7181,RIfc8dd70_6636,RIfce01b0_7572,RIfc7bbc0_6430,
        RIfc90368_6663,RIfc7b8f0_6428,RIe1fa910_4228,RIfcd8b90_7488,RIfc43ec8_5795,RIfc7b788_6427,RIe1f5e88_4175,RIfc7b350_6424,RIfc90d40_6670,RIfca3490_6880,
        RIe1f3b60_4150,RIfc91010_6672,RIfcdb728_7519,RIfcd8758_7485,RIe1ee868_4091,RIe1ec108_4063,RIe1e9408_4031,RIe1e6708_3999,RIe1e3a08_3967,RIe1e0d08_3935,
        RIe1de008_3903,RIe1db308_3871,RIe1d8608_3839,RIe1d2c08_3775,RIe1cff08_3743,RIe1cd208_3711,RIe1ca508_3679,RIe1c7808_3647,RIe1c4b08_3615,RIe1c1e08_3583,
        RIe1bf108_3551,RIf14cf48_5335,RIfc78d58_6397,RIe1b9b40_3490,RIfec5910_8368,RIfc78a88_6395,RIfcd51e8_7447,RIe1b57c0_3442,RIfea1010_8176,RIf1492d0_5292,
        RIfec5a78_8369,RIe1b2c28_3411,RIe1b12d8_3393,RIfec5640_8366,RIf146a08_5263,RIfec57a8_8367,RIfea1178_8177,RIe1a9448_3303,RIe1a6748_3271,RIe1a3a48_3239,
        RIe1a0d48_3207,RIe18d248_2983,RIe179748_2759,RIe2270a0_4734,RIe21bca0_4606,RIe2054a0_4350,RIe1ff500_4282,RIe1f88b8_4205,RIe1f1400_4122,RIe1d5908_3807,
        RIe1bc408_3519,RIe1af280_3370,RIe1718b8_2669,RIdec6350_719,RIdec3650_687,RIfcaf3d0_7016,RIdec0950_655,RIfc6a280_6230,RIdebdc50_623,RIdebaf50_591,
        RIdeb8250_559,RIfc42f50_5784,RIdeb2850_495,RIfc981f8_6753,RIdeafb50_463,RIfc8c6f0_6620,RIdeac838_431,RIdea5f38_399,RIde9f638_367,RIee1d4e8_4792,
        RIfcda648_7507,RIfcc6440_7278,RIfcd5620_7450,RIde92ac8_305,RIfea34a0_8202,RIfea31d0_8200,RIfea3338_8201,RIfcb6b58_7101,RIfcb6888_7099,RIfc9dd60_6818,
        RIee19708_4748,RIfc50c18_5941,RIe16c458_2609,RIfc80a80_6486,RIfec62e8_8375,RIe166350_2540,RIe163650_2508,RIee37d98_5094,RIe160950_2476,RIfcaa678_6961,
        RIe15dc50_2444,RIe158250_2380,RIe155550_2348,RIfea3ba8_8207,RIe152850_2316,RIee35638_5066,RIe14fb50_2284,RIfc62f30_6148,RIe14ce50_2252,RIe14a150_2220,
        RIe147450_2188,RIfc97f28_6751,RIfc89888_6587,RIfc8f558_6653,RIfc52838_5961,RIe141bb8_2125,RIe13f890_2100,RIdf3d798_2076,RIdf3b308_2050,RIee30a48_5012,
        RIfc568e8_6007,RIee2e9f0_4989,RIee2dbe0_4979,RIdf365b0_1995,RIfea38d8_8205,RIfea3a40_8206,RIdf2ff08_1922,RIee2c6c8_4964,RIee2ac10_4945,RIee29590_4929,
        RIee28348_4916,RIdf2ad78_1864,RIdf28e88_1842,RIfea3608_8203,RIfea3770_8204,RIfcc0d10_7216,RIfc75c20_6362,RIfca50b0_6900,RIfc74e10_6352,RIfcc9410_7312,
        RIdf20620_1745,RIfc73628_6335,RIdf1a0e0_1673,RIdf17f20_1649,RIdf15220_1617,RIdf12520_1585,RIdf0f820_1553,RIdf0cb20_1521,RIdf09e20_1489,RIdf07120_1457,
        RIdf04420_1425,RIdefea20_1361,RIdefbd20_1329,RIdef9020_1297,RIdef6320_1265,RIdef3620_1233,RIdef0920_1201,RIdeedc20_1169,RIdeeaf20_1137,RIfcab8c0_6974,
        RIfc7c598_6437,RIfc5beb0_6068,RIfc58ee0_6034,RIdee5688_1074,RIdee3798_1052,RIdee15d8_1028,RIdedf580_1005,RIfcb3048_7059,RIfc72ae8_6327,RIfca3d00_6886,
        RIfcb6450_7096,RIdeda558_948,RIded7f60_921,RIfea3068_8199,RIded3a78_872,RIded1750_847,RIdecea50_815,RIdecbd50_783,RIdec9050_751,RIdeb5550_527,
        RIde98d38_335,RIe16f158_2641,RIe15af50_2412,RIe144750_2156,RIdf39148_2026,RIdf2d7a8_1894,RIdf1e028_1718,RIdf01720_1393,RIdee8220_1105,RIdedcf88_978,
        RIde7ec80_208,RIe19e5e8_3179,RIe19b8e8_3147,RIfca84b8_6937,RIe198be8_3115,RIfc846f8_6529,RIe195ee8_3083,RIe1931e8_3051,RIe1904e8_3019,RIe18aae8_2955,
        RIe187de8_2923,RIfce2be0_7602,RIe1850e8_2891,RIfc8e310_6640,RIe1823e8_2859,RIe17f6e8_2827,RIe17c9e8_2795,RIfcd1570_7404,RIfccc278_7345,RIf1404c8_5191,
        RIfea2d98_8197,RIfcc1b20_7226,RIfc60398_6117,RIee3e5a8_5168,RIee3da68_5160,RIfc642e0_6162,RIfca7f18_6933,RIee3a228_5120,RIfec6180_8374,RIfca9598_6949,
        RIfc5c720_6074,RIfc6bea0_6250,RIfccaec8_7331,RIfc44cd8_5805,RIe224940_4706,RIfcb6180_7094,RIe221c40_4674,RIfc55ad8_5997,RIe21ef40_4642,RIe219540_4578,
        RIe216840_4546,RIfc4dc48_5907,RIe213b40_4514,RIfcdcf10_7536,RIe210e40_4482,RIfcab1b8_6969,RIe20e140_4450,RIe20b440_4418,RIe208740_4386,RIfce3720_7610,
        RIfc64178_6161,RIe203178_4325,RIe201558_4305,RIfcd2ec0_7422,RIf164828_5603,RIfc7f838_6473,RIf162398_5577,RIfcc9c80_7318,RIfca8bc0_6942,RIfea2ac8_8195,
        RIfea2c30_8196,RIfc59318_6037,RIfc4f160_5922,RIf15ac10_5492,RIfcebf88_7707,RIfcbb040_7150,RIfca1870_6860,RIfc93d10_6704,RIe1faeb0_4232,RIf1565c0_5442,
        RIf155a80_5434,RIfc45c50_5816,RIe1f6428_4179,RIfccdbc8_7363,RIfcccae8_7351,RIfca6cd0_6920,RIfec6018_8373,RIfc64010_6160,RIfc434f0_5788,RIfc4c028_5887,
        RIe1eee08_4095,RIe1ec6a8_4067,RIe1e99a8_4035,RIe1e6ca8_4003,RIe1e3fa8_3971,RIe1e12a8_3939,RIe1de5a8_3907,RIe1db8a8_3875,RIe1d8ba8_3843,RIe1d31a8_3779,
        RIe1d04a8_3747,RIe1cd7a8_3715,RIe1caaa8_3683,RIe1c7da8_3651,RIe1c50a8_3619,RIe1c23a8_3587,RIe1bf6a8_3555,RIfc63908_6155,RIfc6bd38_6249,RIe1ba0e0_3494,
        RIe1b7f20_3470,RIfc66fe0_6194,RIfc92ac8_6691,RIe1b5d60_3446,RIfea2f00_8198,RIfc9bfd8_6797,RIfc50d80_5942,RIe1b31c8_3415,RIe1b1878_3397,RIfc4df18_5909,
        RIfc9d658_6813,RIe1ad0c0_3346,RIe1ab8d8_3329,RIe1a99e8_3307,RIe1a6ce8_3275,RIe1a3fe8_3243,RIe1a12e8_3211,RIe18d7e8_2987,RIe179ce8_2763,RIe227640_4738,
        RIe21c240_4610,RIe205a40_4354,RIe1ffaa0_4286,RIe1f8e58_4209,RIe1f19a0_4126,RIe1d5ea8_3811,RIe1bc9a8_3523,RIe1af820_3374,RIe171e58_2673,RIdec61e8_718,
        RIdec34e8_686,RIee20620_4827,RIdec07e8_654,RIfc4b7b8_5881,RIdebdae8_622,RIdebade8_590,RIdeb80e8_558,RIfc41150_5766,RIdeb26e8_494,RIfc87830_6564,
        RIdeaf9e8_462,RIee1dec0_4799,RIdeac4f0_430,RIdea5bf0_398,RIde9f2f0_366,RIee1d380_4791,RIfc77c78_6385,RIfc84f68_6535,RIfc6ff50_6296,RIde92780_304,
        RIde8efb8_287,RIde8ae18_267,RIde86c78_247,RIee1a680_4759,RIee19f78_4754,RIfcd7240_7470,RIfcbeb50_7192,RIfc76328_6367,RIe16c2f0_2608,RIee388d8_5102,
        RIfea20f0_8188,RIe1661e8_2539,RIe1634e8_2507,RIee37c30_5093,RIe1607e8_2475,RIfce7500_7654,RIe15dae8_2443,RIe1580e8_2379,RIe1553e8_2347,RIfc3f698_5747,
        RIe1526e8_2315,RIee354d0_5065,RIe14f9e8_2283,RIfc83e88_6523,RIe14cce8_2251,RIe149fe8_2219,RIe1472e8_2187,RIfcea4d0_7688,RIfcb7ad0_7112,RIfc695d8_6221,
        RIfc51a28_5951,RIe141a50_2124,RIe13f728_2099,RIdf3d630_2075,RIdf3b1a0_2049,RIfca9e08_6955,RIee2fda0_5003,RIfc88a78_6577,RIee2da78_4978,RIdf36448_1994,
        RIdf33fb8_1968,RIdf31df8_1944,RIfea2258_8189,RIee2c560_4963,RIee2aaa8_4944,RIee29428_4928,RIee281e0_4915,RIdf2ac10_1863,RIdf28d20_1841,RIfea27f8_8193,
        RIfea2960_8194,RIfcdabe8_7511,RIfca08f8_6849,RIfc8b1d8_6605,RIfc49058_5853,RIfca0a60_6850,RIdf204b8_1744,RIfc99cb0_6772,RIdf19f78_1672,RIdf17db8_1648,
        RIdf150b8_1616,RIdf123b8_1584,RIdf0f6b8_1552,RIdf0c9b8_1520,RIdf09cb8_1488,RIdf06fb8_1456,RIdf042b8_1424,RIdefe8b8_1360,RIdefbbb8_1328,RIdef8eb8_1296,
        RIdef61b8_1264,RIdef34b8_1232,RIdef07b8_1200,RIdeedab8_1168,RIdeeadb8_1136,RIfcd1f48_7411,RIfc57f68_6023,RIfcbe2e0_7186,RIfcd8fc8_7491,RIdee5520_1073,
        RIfea2690_8192,RIdee1470_1027,RIdedf418_1004,RIfc57b30_6020,RIfcb35e8_7063,RIfcbd7a0_7178,RIfc91178_6673,RIfea2528_8191,RIded7df8_920,RIfea23c0_8190,
        RIded3910_871,RIded15e8_846,RIdece8e8_814,RIdecbbe8_782,RIdec8ee8_750,RIdeb53e8_526,RIde989f0_334,RIe16eff0_2640,RIe15ade8_2411,RIe1445e8_2155,
        RIdf38fe0_2025,RIdf2d640_1893,RIdf1dec0_1717,RIdf015b8_1392,RIdee80b8_1104,RIdedce20_977,RIde7e938_207,RIe19e480_3178,RIe19b780_3146,RIfccc980_7350,
        RIe198a80_3114,RIfcc1148_7219,RIe195d80_3082,RIe193080_3050,RIe190380_3018,RIe18a980_2954,RIe187c80_2922,RIfcb2ee0_7058,RIe184f80_2890,RIfc615e0_6130,
        RIe182280_2858,RIe17f580_2826,RIe17c880_2794,RIfc69038_6217,RIfc4c898_5893,RIfc6f2a8_6287,RIe1764a8_2723,RIfcad0a8_6991,RIfc6adc0_6238,RIfc70388_6299,
        RIfea1b50_8184,RIfea1f88_8187,RIfc56e88_6011,RIfea1cb8_8185,RIe174450_2700,RIfc60d70_6124,RIfc6a820_6234,RIfea1e20_8186,RIf16d798_5705,RIfc40bb0_5762,
        RIe2247d8_4705,RIfc77138_6377,RIe221ad8_4673,RIfcd7d80_7478,RIe21edd8_4641,RIe2193d8_4577,RIe2166d8_4545,RIfc40070_5754,RIe2139d8_4513,RIf169850_5660,
        RIe210cd8_4481,RIfcc1580_7222,RIe20dfd8_4449,RIe20b2d8_4417,RIe2085d8_4385,RIfcd0058_7389,RIfc749d8_6349,RIe203010_4324,RIe2013f0_4304,RIfc60230_6116,
        RIfc60668_6119,RIfcaf970_7020,RIfc45818_5813,RIf160a48_5559,RIf15eb58_5537,RIfea1880_8182,RIfea19e8_8183,RIfc72110_6320,RIfc49b98_5861,RIfcca0b8_7321,
        RIfc71738_6313,RIfc4ca00_5894,RIfc71030_6308,RIfcde428_7551,RIe1fad48_4231,RIfc70bf8_6305,RIfc63a70_6156,RIfca7db0_6932,RIe1f62c0_4178,RIfcada80_6998,
        RIfc6fde8_6295,RIfc6f578_6289,RIe1f3f98_4153,RIfcde158_7549,RIfcad378_6993,RIfc65f00_6182,RIe1eeca0_4094,RIe1ec540_4066,RIe1e9840_4034,RIe1e6b40_4002,
        RIe1e3e40_3970,RIe1e1140_3938,RIe1de440_3906,RIe1db740_3874,RIe1d8a40_3842,RIe1d3040_3778,RIe1d0340_3746,RIe1cd640_3714,RIe1ca940_3682,RIe1c7c40_3650,
        RIe1c4f40_3618,RIe1c2240_3586,RIe1bf540_3554,RIfc69308_6219,RIfccba08_7339,RIe1b9f78_3493,RIe1b7db8_3469,RIfccd628_7359,RIfc69740_6222,RIe1b5bf8_3445,
        RIe1b4578_3429,RIfccf950_7384,RIf148088_5279,RIe1b3060_3414,RIe1b1710_3396,RIfc9f818_6837,RIfcb9c90_7136,RIe1acf58_3345,RIe1ab770_3328,RIe1a9880_3306,
        RIe1a6b80_3274,RIe1a3e80_3242,RIe1a1180_3210,RIe18d680_2986,RIe179b80_2762,RIe2274d8_4737,RIe21c0d8_4609,RIe2058d8_4353,RIe1ff938_4285,RIe1f8cf0_4208,
        RIe1f1838_4125,RIe1d5d40_3810,RIe1bc840_3522,RIe1af6b8_3373,RIe171cf0_2672,R_58_102f1b78,R_59_be1fc68,R_5a_10279198,R_5b_102299e8,R_5c_101d0448,
        R_5d_f7f82f0,R_5e_be21600,R_5f_f7fa5b8,R_60_1027d530,R_61_10205ae8,R_62_10283510,R_63_f82b578,R_64_ace4e68,R_65_f8204e0,R_66_1027a0b0,
        R_67_1022dc30,R_68_102478a8,R_69_10286f78,R_6a_f7edd80,R_6b_101c3628,R_6c_f7fbe00,R_6d_f7ce9f8,R_6e_f7c8830,R_6f_101ffc68,R_70_f7d4000,
        R_71_acee958,R_72_94046c0,R_73_101ee420,R_74_102eb268,R_75_b320c50,R_76_ad80a90,R_77_1027fd48,R_78_f7ce4b8,R_79_ad77048,R_7a_102a6ae0,
        R_7b_f7e4c78,R_7c_e2a6ce0,R_7d_101e86e0,R_7e_e2a9cc8,R_7f_10292be0,R_80_b33cde8,R_81_101e2908,R_82_102e9780,R_83_f8157a0,R_84_f819358,
        R_85_ace8b70,R_86_be142b0,R_87_f81b770,R_88_b330278,R_89_f7fe9f8,R_8a_101cf488,R_8b_f8225c0,R_8c_101d4738,R_8d_101c4000,R_8e_101fe960,
        R_8f_102a0330,R_90_f7f4bd0,R_91_1023e5a8,R_92_10248da8,R_93_be2c938,R_94_f7f5458,R_95_f7c6808,R_96_be316a8,R_97_e2a0328,R_98_be2d850,
        R_99_10217db0,R_9a_f7ec340,R_9b_be23ec0,R_9c_101d4540,R_9d_f800828,R_9e_102970c8,R_9f_10221de0,R_a0_ad8d568,R_a1_be4eb58,R_a2_f7c5500,
        R_a3_ad88f30,R_a4_f82f088,R_a5_f7dcbc8,R_a6_10292940,R_a7_be138d8,R_a8_acee418,R_a9_ad84450,R_aa_be10838,R_ab_be31fd8,R_ac_acdaef0,
        R_ad_acea908,R_ae_101f8830,R_af_f7dec98,R_b0_101e2c50,R_b1_f801b30,R_b2_be16e00,R_b3_102e3cf0,R_b4_10291788);
input RIdec64b8_720,RIbc62af0_23,RIbc62a78_22,RIbc62a00_21,RIbc62988_20,RIbc62910_19,RIbc62898_18,RIbc62820_17,RIbc627a8_16,
        RIbc62730_15,RIbc626b8_14,RIbc62640_13,RIdec37b8_688,RIfc8daa0_6634,RIdec0ab8_656,RIfc56348_6003,RIdebddb8_624,RIdebb0b8_592,RIdeb83b8_560,
        RIfc98798_6757,RIdeb29b8_496,RIfcbd098_7173,RIdeafcb8_464,RIfc8dc08_6635,RIdeacb80_432,RIdea6280_400,RIde9f980_368,RIfcd6868_7463,RIfc8ded8_6637,
        RIfc7dd80_6454,RIfc56618_6005,RIde92e10_306,RIde8f300_288,RIde8b160_268,RIde86fc0_248,RIde82ad8_227,RIfc8e040_6638,RIfcd96d0_7496,RIfca1e10_6864,
        RIfcbd200_7174,RIe16c5c0_2610,RIe16a298_2585,RIe168ab0_2568,RIe1664b8_2541,RIe1637b8_2509,RIee37f00_5095,RIe160ab8_2477,RIfc8ea18_6645,RIe15ddb8_2445,
        RIe1583b8_2381,RIe1556b8_2349,RIfe9f828_8159,RIe1529b8_2317,RIfe9f990_8160,RIe14fcb8_2285,RIfcbd368_7175,RIe14cfb8_2253,RIe14a2b8_2221,RIe1475b8_2189,
        RIfc8ee50_6648,RIfc45278_5809,RIfc98360_6754,RIfca2248_6867,RIe141d20_2126,RIe13f9f8_2101,RIdf3d900_2077,RIdf3b470_2051,RIfcd6ca0_7466,RIee2ff08_5004,
        RIfc8ece8_6647,RIee2dd48_4980,RIdf36718_1996,RIdf34120_1969,RIdf31f60_1945,RIfe9f6c0_8158,RIfcb4560_7074,RIfc45db8_5817,RIfc8e1a8_6639,RIfc7d678_6449,
        RIdf2aee0_1865,RIdf28ff0_1843,RIdf26e30_1819,RIdf25378_1800,RIfcb43f8_7073,RIfc8e748_6643,RIdf23488_1778,RIfcc2c00_7238,RIdf21e08_1762,RIdf20788_1746,
        RIdf1b760_1689,RIdf1a248_1674,RIdf18088_1650,RIdf15388_1618,RIdf12688_1586,RIdf0f988_1554,RIdf0cc88_1522,RIdf09f88_1490,RIdf07288_1458,RIdf04588_1426,
        RIdefeb88_1362,RIdefbe88_1330,RIdef9188_1298,RIdef6488_1266,RIdef3788_1234,RIdef0a88_1202,RIdeedd88_1170,RIdeeb088_1138,RIfc8efb8_6649,RIfc44e40_5806,
        RIfc57860_6018,RIfca23b0_6868,RIfe9faf8_8161,RIdee3900_1053,RIdee1740_1029,RIdedf6e8_1006,RIfcbd4d0_7176,RIee22678_4850,RIfc98090_6752,RIee21598_4838,
        RIfe9fc60_8162,RIded80c8_922,RIfe9fdc8_8163,RIded3be0_873,RIded18b8_848,RIdecebb8_816,RIdecbeb8_784,RIdec91b8_752,RIdeb56b8_528,RIde99080_336,
        RIe16f2c0_2642,RIe15b0b8_2413,RIe1448b8_2157,RIdf392b0_2027,RIdf2d910_1895,RIdf1e190_1719,RIdf01888_1394,RIdee8388_1106,RIdedd0f0_979,RIde7efc8_209,
        RIe19e750_3180,RIbc625c8_12,RIbc62550_11,RIbc624d8_10,RIbc62460_9,RIbc623e8_8,RIbc62370_7,RIbc622f8_6,RIbc62280_5,RIbc62208_4,
        RIbc62190_3,RIbc62118_2,RIe19ba50_3148,RIfc479d8_5837,RIe198d50_3116,RIfe9f558_8157,RIe196050_3084,RIe193350_3052,RIe190650_3020,RIe18ac50_2956,
        RIe187f50_2924,RIfc47870_5836,RIe185250_2892,RIf142ef8_5221,RIe182550_2860,RIe17f850_2828,RIe17cb50_2796,RIfcb5208_7083,RIfcbc6c0_7166,RIe177588_2735,
        RIe176610_2724,RIf13fdc0_5186,RIfe9f3f0_8156,RIfce40f8_7617,RIfc47708_5835,RIfc47438_5833,RIfca15a0_6858,RIfc99170_6764,RIe1745b8_2701,RIfc8cc90_6624,
        RIfc556a0_5994,RIfc7ee60_6466,RIfce8e50_7672,RIfe9f288_8155,RIe224aa8_4707,RIfc55808_5995,RIe221da8_4675,RIfcb50a0_7082,RIe21f0a8_4643,RIe2196a8_4579,
        RIe2169a8_4547,RIfcbc828_7167,RIe213ca8_4515,RIfc47000_5830,RIe210fa8_4483,RIfcbc990_7168,RIe20e2a8_4451,RIe20b5a8_4419,RIe2088a8_4387,RIfc46bc8_5827,
        RIfcd6598_7461,RIe2032e0_4326,RIe2016c0_4306,RIfc98ea0_6762,RIfc7eb90_6464,RIfce0318_7573,RIfcbcaf8_7169,RIfc8cf60_6626,RIfcb4dd0_7080,RIe1fd340_4258,
        RIe1fc260_4246,RIf15cf38_5517,RIfe9f120_8154,RIfc7ea28_6463,RIfc8d0c8_6627,RIfcbcc60_7170,RIfc98bd0_6760,RIfce2d48_7603,RIe1fb018_4233,RIfc55f10_6000,
        RIfc7e8c0_6462,RIfc8d230_6628,RIe1f6590_4180,RIfce58e0_7634,RIfc468f8_5825,RIfcc2ed0_7240,RIe1f4100_4154,RIfceedf0_7740,RIfc8d398_6629,RIfc8d500_6630,
        RIe1eef70_4096,RIe1ec810_4068,RIe1e9b10_4036,RIe1e6e10_4004,RIe1e4110_3972,RIe1e1410_3940,RIe1de710_3908,RIe1dba10_3876,RIe1d8d10_3844,RIe1d3310_3780,
        RIe1d0610_3748,RIe1cd910_3716,RIe1cac10_3684,RIe1c7f10_3652,RIe1c5210_3620,RIe1c2510_3588,RIe1bf810_3556,RIf14d0b0_5336,RIfe9efb8_8153,RIe1ba248_3495,
        RIe1b8088_3471,RIfec4dd0_8360,RIfec50a0_8362,RIe1b5ec8_3447,RIe1b46e0_3430,RIfcb4998_7077,RIfcb4c68_7079,RIfec5370_8364,RIfe9ee50_8152,RIfcbcdc8_7171,
        RIfc46358_5821,RIfec5208_8363,RIfec4f38_8361,RIe1a9b50_3308,RIe1a6e50_3276,RIe1a4150_3244,RIe1a1450_3212,RIe18d950_2988,RIe179e50_2764,RIe2277a8_4739,
        RIe21c3a8_4611,RIe205ba8_4355,RIe1ffc08_4287,RIe1f8fc0_4210,RIe1f1b08_4127,RIe1d6010_3812,RIe1bcb10_3524,RIe1af988_3375,RIe171fc0_2674,RIdec6080_717,
        RIdec3380_685,RIee204b8_4826,RIdec0680_653,RIfcd70d8_7469,RIdebd980_621,RIdebac80_589,RIdeb7f80_557,RIfcbe448_7187,RIdeb2580_493,RIfcb3480_7062,
        RIdeaf880_461,RIfc43928_5791,RIdeac1a8_429,RIdea58a8_397,RIde9efa8_365,RIfcd88c0_7486,RIee1c408_4780,RIfcc77f0_7292,RIfea04d0_8168,RIde92438_303,
        RIde8ec70_286,RIde8aad0_266,RIde86930_246,RIfca31c0_6878,RIfc59a20_6042,RIfcd1de0_7410,RIfc91448_6675,RIfc97280_6742,RIe16c188_2607,RIfc97118_6741,
        RIe168948_2567,RIe166080_2538,RIe163380_2506,RIee37ac8_5092,RIe160680_2474,RIfcd1c78_7409,RIe15d980_2442,RIe157f80_2378,RIe155280_2346,RIfc3f530_5746,
        RIe152580_2314,RIee35368_5064,RIe14f880_2282,RIfc7a3d8_6413,RIe14cb80_2250,RIe149e80_2218,RIe147180_2186,RIfc42b18_5781,RIfc7a270_6412,RIfc5a560_6050,
        RIfc96b78_6737,RIfea6fb0_8216,RIe13f5c0_2098,RIdf3d4c8_2074,RIdf3b038_2048,RIfce5bb0_7636,RIee2fc38_5002,RIfc91cb8_6681,RIee2d910_4977,RIdf362e0_1993,
        RIdf33e50_1967,RIdf31c90_1943,RIdf2fda0_1921,RIfc43658_5789,RIfc59e58_6045,RIfc96fb0_6740,RIfc7ac48_6419,RIfea0368_8167,RIdf28bb8_1840,RIdf26cc8_1818,
        RIdf25210_1799,RIfc91718_6677,RIfcb3318_7061,RIfc919e8_6679,RIfc91880_6678,RIfc430b8_5785,RIdf20350_1743,RIfc7a978_6417,RIdf19e10_1671,RIdf17c50_1647,
        RIdf14f50_1615,RIdf12250_1583,RIdf0f550_1551,RIdf0c850_1519,RIdf09b50_1487,RIdf06e50_1455,RIdf04150_1423,RIdefe750_1359,RIdefba50_1327,RIdef8d50_1295,
        RIdef6050_1263,RIdef3350_1231,RIdef0650_1199,RIdeed950_1167,RIdeeac50_1135,RIfcd1b10_7408,RIfc968a8_6735,RIfc91f88_6683,RIfcdfc10_7568,RIfea99e0_8246,
        RIdee3630_1051,RIdee1308_1026,RIdedf2b0_1003,RIfcc7d90_7296,RIfcd85f0_7484,RIfce3888_7611,RIfc5a830_6052,RIdeda3f0_947,RIfea9878_8245,RIded5f08_898,
        RIded37a8_870,RIded1480_845,RIdece780_813,RIdecba80_781,RIdec8d80_749,RIdeb5280_525,RIde986a8_333,RIe16ee88_2639,RIe15ac80_2410,RIe144480_2154,
        RIdf38e78_2024,RIdf2d4d8_1892,RIdf1dd58_1716,RIdf01450_1391,RIdee7f50_1103,RIdedccb8_976,RIde7e5f0_206,RIe19e318_3177,RIe19b618_3145,RIfc8f3f0_6652,
        RIe198918_3113,RIf144b18_5241,RIe195c18_3081,RIe192f18_3049,RIe190218_3017,RIe18a818_2953,RIe187b18_2921,RIf143d08_5231,RIe184e18_2889,RIfcb3cf0_7068,
        RIe182118_2857,RIe17f418_2825,RIe17c718_2793,RIfc448a0_5802,RIf141170_5200,RIfc7c9d0_6440,RIfea0098_8165,RIfc57e00_6022,RIf13f550_5180,RIfcd6e08_7467,
        RIee3d900_5159,RIfc8f6c0_6654,RIfce0048_7571,RIfca27e8_6871,RIe1742e8_2699,RIfc7c700_6438,RIfc8f990_6656,RIfce9828_7679,RIfc583a0_6026,RIf16cdc0_5698,
        RIe224670_4704,RIf16c118_5689,RIe221970_4672,RIfc58508_6027,RIe21ec70_4640,RIe219270_4576,RIe216570_4544,RIfc3ff08_5753,RIe213870_4512,RIf1696e8_5659,
        RIe210b70_4480,RIfc58940_6030,RIe20de70_4448,RIe20b170_4416,RIe208470_4384,RIfc8fc60_6658,RIfc97820_6746,RIe202ea8_4323,RIe201288_4303,RIfcc27c8_7235,
        RIfcdfee0_7570,RIfc44198_5797,RIfc58670_6028,RIf1608e0_5558,RIf15e9f0_5536,RIfe9ff30_8164,RIe1fc0f8_4245,RIfc7be90_6432,RIf15bb88_5503,RIfcd8cf8_7489,
        RIfcd8e60_7490,RIfca2d88_6875,RIfcbdea8_7183,RIfcb3a20_7066,RIe1fabe0_4230,RIfc90098_6661,RIfc90200_6662,RIfcd20b0_7412,RIe1f6158_4177,RIfc904d0_6664,
        RIfca2ef0_6876,RIfc97550_6744,RIe1f3e30_4152,RIfc59048_6035,RIfc907a0_6666,RIfc90638_6665,RIe1eeb38_4093,RIe1ec3d8_4065,RIe1e96d8_4033,RIe1e69d8_4001,
        RIe1e3cd8_3969,RIe1e0fd8_3937,RIe1de2d8_3905,RIe1db5d8_3873,RIe1d88d8_3841,RIe1d2ed8_3777,RIe1d01d8_3745,RIe1cd4d8_3713,RIe1ca7d8_3681,RIe1c7ad8_3649,
        RIe1c4dd8_3617,RIe1c20d8_3585,RIe1bf3d8_3553,RIfcc73b8_7289,RIfce3cc0_7614,RIe1b9e10_3492,RIe1b7c50_3468,RIfcd6f70_7468,RIf149e10_5300,RIe1b5a90_3444,
        RIfea0200_8166,RIfc90bd8_6669,RIfcdfd78_7569,RIe1b2ef8_3413,RIe1b15a8_3395,RIfc973e8_6743,RIfcc7520_7290,RIe1acdf0_3344,RIe1ab608_3327,RIe1a9718_3305,
        RIe1a6a18_3273,RIe1a3d18_3241,RIe1a1018_3209,RIe18d518_2985,RIe179a18_2761,RIe227370_4736,RIe21bf70_4608,RIe205770_4352,RIe1ff7d0_4284,RIe1f8b88_4207,
        RIe1f16d0_4124,RIe1d5bd8_3809,RIe1bc6d8_3521,RIe1af550_3372,RIe171b88_2671,RIdec5108_706,RIdec2408_674,RIfc93608_6699,RIdebf708_642,RIfc934a0_6698,
        RIdebca08_610,RIdeb9d08_578,RIdeb7008_546,RIfcdf7d8_7565,RIdeb1608_482,RIfc78218_6389,RIdeae908_450,RIfcc8498_7301,RIdea9d90_418,RIdea3490_386,
        RIde9cb90_354,RIee1cc78_4786,RIee1bb98_4774,RIee1b328_4768,RIee1aab8_4762,RIde909f8_295,RIde8d578_279,RIfea8ea0_8238,RIde85238_239,RIde813e0_220,
        RIfc938d8_6701,RIfce5e80_7638,RIfcbfd98_7205,RIfce8ce8_7671,RIe16b4e0_2598,RIfea8d38_8237,RIfea9f80_8250,RIe165108_2527,RIe162408_2495,RIfc779a8_6383,
        RIe15f708_2463,RIfe9dc08_8139,RIe15ca08_2431,RIe157008_2367,RIe154308_2335,RIfea7550_8220,RIe151608_2303,RIfcd6160_7458,RIe14e908_2271,RIfcd1408_7403,
        RIe14bc08_2239,RIe148f08_2207,RIe146208_2175,RIfceb718_7701,RIfcb19c8_7043,RIfc93e78_6705,RIfce7938_7657,RIe140da8_2115,RIdf3ecb0_2091,RIdf3c988_2066,
        RIfe9daa0_8138,RIfce8478_7665,RIfcdbf98_7525,RIfc776d8_6381,RIfc93fe0_6706,RIdf354d0_1983,RIdf33040_1957,RIdf30fe8_1934,RIdf2ee28_1910,RIee2ba20_4955,
        RIfc93ba8_6703,RIfc77de0_6386,RIee27ad8_4910,RIfe9d668_8135,RIfea8bd0_8236,RIdf26458_1812,RIfe9d7d0_8136,RIfcb1c98_7045,RIee26cc8_4900,RIdf22ab0_1771,
        RIfcc0068_7207,RIdf21598_1756,RIdf1f6a8_1734,RIdf1aef0_1683,RIfe9d938_8137,RIdf16cd8_1636,RIdf13fd8_1604,RIdf112d8_1572,RIdf0e5d8_1540,RIdf0b8d8_1508,
        RIdf08bd8_1476,RIdf05ed8_1444,RIdf031d8_1412,RIdefd7d8_1348,RIdefaad8_1316,RIdef7dd8_1284,RIdef50d8_1252,RIdef23d8_1220,RIdeef6d8_1188,RIdeec9d8_1156,
        RIdee9cd8_1124,RIfc942b0_6708,RIfcde6f8_7553,RIfcd1138_7401,RIfcde860_7554,RIdee4878_1064,RIdee2af0_1043,RIdee0a98_1020,RIdede8d8_996,RIfc5c9f0_6076,
        RIee22240_4847,RIfcc8768_7303,RIee21160_4835,RIded95e0_937,RIded7150_911,RIded5260_889,RIfea76b8_8221,RIded0508_834,RIdecd808_802,RIdecab08_770,
        RIdec7e08_738,RIdeb4308_514,RIde96290_322,RIe16df10_2628,RIe159d08_2399,RIe143508_2143,RIdf37f00_2013,RIdf2c560_1881,RIdf1cde0_1705,RIdf004d8_1380,
        RIdee6fd8_1092,RIdedbd40_965,RIde7c1d8_195,RIe19d3a0_3166,RIe19a6a0_3134,RIfcb2c10_7056,RIe1979a0_3102,RIfc923c0_6686,RIe194ca0_3070,RIe191fa0_3038,
        RIe18f2a0_3006,RIe1898a0_2942,RIe186ba0_2910,RIfc422a8_5775,RIe183ea0_2878,RIfcbecb8_7193,RIe1811a0_2846,RIe17e4a0_2814,RIe17b7a0_2782,RIf142250_5212,
        RIf140bd0_5196,RIfec43f8_8353,RIe175968_2715,RIfc79b68_6407,RIf13efb0_5176,RIfc92528_6687,RIfcb2aa8_7055,RIfcd8320_7482,RIfcea200_7686,RIfc79898_6405,
        RIe1734d8_2689,RIfcd7948_7475,RIfcd7678_7473,RIf16e170_5712,RIfc927f8_6689,RIfc92960_6690,RIe2236f8_4693,RIfc795c8_6403,RIe2209f8_4661,RIf16ad68_5675,
        RIe21dcf8_4629,RIe2182f8_4565,RIe2155f8_4533,RIfe9d398_8133,RIe2128f8_4501,RIfcdb9f8_7521,RIe20fbf8_4469,RIfc41d08_5771,RIe20cef8_4437,RIe20a1f8_4405,
        RIe2074f8_4373,RIfcd7510_7472,RIf166010_5620,RIfe9d230_8132,RIe2008b0_4296,RIf165098_5609,RIfc41ba0_5770,RIfc41a38_5769,RIfc92c30_6692,RIfc418d0_5768,
        RIfc79190_6400,RIe1fcad0_4252,RIfec4560_8354,RIfc79028_6399,RIfcbf258_7197,RIfcc1df0_7228,RIfcd81b8_7481,RIfc92d98_6693,RIfc5b4d8_6061,RIfcd77e0_7474,
        RIe1fa0a0_4222,RIf156188_5439,RIfe9d500_8134,RIf1546d0_5420,RIe1f5348_4167,RIfec4830_8356,RIfec46c8_8355,RIf1508f0_5376,RIe1f3020_4142,RIfce3180_7606,
        RIfce8fb8_7673,RIfcbf690_7200,RIe1edd28_4083,RIe1eb460_4054,RIe1e8760_4022,RIe1e5a60_3990,RIe1e2d60_3958,RIe1e0060_3926,RIe1dd360_3894,RIe1da660_3862,
        RIe1d7960_3830,RIe1d1f60_3766,RIe1cf260_3734,RIe1cc560_3702,RIe1c9860_3670,RIe1c6b60_3638,RIe1c3e60_3606,RIe1c1160_3574,RIe1be460_3542,RIfe9d0c8_8131,
        RIfe9cc90_8128,RIe1b9168_3483,RIe1b7110_3460,RIf14a3b0_5304,RIfe9cb28_8127,RIfe9cf60_8130,RIfe9c9c0_8126,RIfce2208_7595,RIfce9558_7677,RIfe9c858_8125,
        RIfe9cdf8_8129,RIf147110_5268,RIf146468_5259,RIe1ac2b0_3336,RIe1aaac8_3319,RIe1a87a0_3294,RIe1a5aa0_3262,RIe1a2da0_3230,RIe1a00a0_3198,RIe18c5a0_2974,
        RIe178aa0_2750,RIe2263f8_4725,RIe21aff8_4597,RIe2047f8_4341,RIe1fe858_4273,RIe1f7c10_4196,RIe1f0758_4113,RIe1d4c60_3798,RIe1bb760_3510,RIe1ae5d8_3361,
        RIe170c10_2660,RIdec4190_695,RIdec1490_663,RIfceaa70_7692,RIdebe790_631,RIfc954f8_6721,RIdebba90_599,RIdeb8d90_567,RIdeb6090_535,RIfcebb50_7704,
        RIdeb0690_471,RIee1e190_4801,RIdead990_439,RIfcdf0d0_7560,RIdea7978_407,RIdea1078_375,RIde9a778_343,RIee1c840_4783,RIfc957c8_6723,RIfcc8e70_7308,
        RIfc5e610_6096,RIfe9e8b0_8148,RIde8c1c8_273,RIde88028_253,RIde83b40_232,RIfcb0bb8_7033,RIfca4b10_6896,RIfc75d88_6363,RIfca4c78_6897,RIfc95390_6720,
        RIe16a9a0_2590,RIfcc8fd8_7309,RIe166e90_2548,RIe164190_2516,RIe161490_2484,RIfe9e748_8147,RIe15e790_2452,RIfc74f78_6353,RIe15ba90_2420,RIe156090_2356,
        RIe153390_2324,RIfc3ecc0_5740,RIe150690_2292,RIfce8b80_7670,RIe14d990_2260,RIfca6730_6916,RIe14ac90_2228,RIe147f90_2196,RIe145290_2164,RIfcee2b0_7732,
        RIfc5f2b8_6105,RIfc753b0_6356,RIfc74b40_6350,RIe140268_2107,RIdf3e170_2083,RIdf3be48_2058,RIdf39c88_2034,RIfcc1c88_7227,RIfcc1850_7224,RIfc965d8_6733,
        RIfc96038_6729,RIdf34828_1974,RIdf327d0_1951,RIdf301d8_1924,RIdf2e2e8_1902,RIfc5e778_6097,RIfcd0328_7391,RIfc757e8_6359,RIfcee6e8_7735,RIdf296f8_1848,
        RIdf273d0_1823,RIdf257b0_1803,RIdf23b90_1783,RIfc95d68_6727,RIfceda40_7726,RIfe9eb80_8150,RIfc75518_6357,RIfcd01c0_7390,RIdf1eb68_1726,RIfe9ece8_8151,
        RIfe9ea18_8149,RIdf15d60_1625,RIdf13060_1593,RIdf10360_1561,RIdf0d660_1529,RIdf0a960_1497,RIdf07c60_1465,RIdf04f60_1433,RIdf02260_1401,RIdefc860_1337,
        RIdef9b60_1305,RIdef6e60_1273,RIdef4160_1241,RIdef1460_1209,RIdeee760_1177,RIdeeba60_1145,RIdee8d60_1113,RIfc961a0_6730,RIfc96308_6731,RIfc5ee80_6102,
        RIfce6150_7640,RIdee42d8_1060,RIdee1e48_1034,RIdee00c0_1013,RIdeddac8_986,RIfc96470_6732,RIfc75248_6355,RIfc74ca8_6351,RIfcb0618_7029,RIded8938_928,
        RIded6610_903,RIded4450_879,RIded2290_855,RIdecf590_823,RIdecc890_791,RIdec9b90_759,RIdec6e90_727,RIdeb3390_503,RIde93e78_311,RIe16cf98_2617,
        RIe158d90_2388,RIe142590_2132,RIdf36f88_2002,RIdf2b5e8_1870,RIdf1be68_1694,RIdeff560_1369,RIdee6060_1081,RIdedadc8_954,RIde79dc0_184,RIe19c428_3155,
        RIe199728_3123,RIfe9e310_8144,RIe196a28_3091,RIfcc04a0_7210,RIe193d28_3059,RIe191028_3027,RIe18e328_2995,RIe188928_2931,RIe185c28_2899,RIfce1830_7588,
        RIe182f28_2867,RIfe9e478_8145,RIe180228_2835,RIe17d528_2803,RIe17a828_2771,RIf141878_5205,RIfcb12c0_7038,RIfc94418_6709,RIe174f90_2708,RIfc77408_6379,
        RIf13ea10_5172,RIfcdc100_7526,RIfc94580_6710,RIfc946e8_6711,RIfced338_7721,RIfce5fe8_7639,RIe172998_2681,RIfcdc268_7527,RIfcddff0_7548,RIfcc0608_7211,
        RIfce7230_7652,RIfc40340_5756,RIe222780_4682,RIfcdd618_7541,RIe21fa80_4650,RIfcd0b98_7397,RIe21cd80_4618,RIe217380_4554,RIe214680_4522,RIfec4998_8357,
        RIe211980_4490,RIf168608_5647,RIe20ec80_4458,RIfcc0770_7212,RIe20bf80_4426,RIe209280_4394,RIe206580_4362,RIfce2370_7596,RIfcee580_7734,RIfec4c68_8359,
        RIfec4b00_8358,RIfc949b8_6713,RIfcebcb8_7705,RIf162938_5581,RIf1612b8_5565,RIfccd088_7355,RIfcc08d8_7213,RIfe9e040_8142,RIfe9e1a8_8143,RIfcead40_7694,
        RIf15ad78_5493,RIfc94c88_6715,RIfccc3e0_7346,RIfc765f8_6369,RIfc94df0_6716,RIfcc0a40_7214,RIe1f9998_4217,RIfcc8d08_7307,RIfce8748_7667,RIfceb2e0_7698,
        RIe1f4970_4160,RIf152510_5396,RIf1512c8_5383,RIfcb0ff0_7036,RIe1f24e0_4134,RIfc761c0_6366,RIfc950c0_6718,RIfcc0e78_7217,RIe1ed1e8_4075,RIe1ea4e8_4043,
        RIe1e77e8_4011,RIe1e4ae8_3979,RIe1e1de8_3947,RIe1df0e8_3915,RIe1dc3e8_3883,RIe1d96e8_3851,RIe1d69e8_3819,RIe1d0fe8_3755,RIe1ce2e8_3723,RIe1cb5e8_3691,
        RIe1c88e8_3659,RIe1c5be8_3627,RIe1c2ee8_3595,RIe1c01e8_3563,RIe1bd4e8_3531,RIf14bfd0_5324,RIf14ac20_5310,RIfe9ded8_8141,RIe1b65d0_3452,RIfcecd98_7717,
        RIfc76490_6368,RIe1b4c80_3434,RIe1b38d0_3420,RIfcc0fe0_7218,RIfceaea8_7695,RIe1b1f80_3402,RIe1b0360_3382,RIfcd0760_7394,RIf145ec8_5255,RIfe9e5e0_8146,
        RIfe9dd70_8140,RIe1a7828_3283,RIe1a4b28_3251,RIe1a1e28_3219,RIe19f128_3187,RIe18b628_2963,RIe177b28_2739,RIe225480_4714,RIe21a080_4586,RIe203880_4330,
        RIe1fd8e0_4262,RIe1f6c98_4185,RIe1ef7e0_4102,RIe1d3ce8_3787,RIe1ba7e8_3499,RIe1ad660_3350,RIe16fc98_2649,RIdec6788_722,RIdec3a88_690,RIee20788_4828,
        RIdec0d88_658,RIee1f810_4817,RIdebe088_626,RIdebb388_594,RIdeb8688_562,RIfc9b1c8_6787,RIdeb2c88_498,RIfce1f38_7593,RIdeaff88_466,RIfc892e8_6583,
        RIdead210_434,RIdea6910_402,RIdea0010_370,RIee1d650_4793,RIee1c570_4781,RIee1b5f8_4770,RIee1aef0_4765,RIfe99888_8091,RIfe99450_8088,RIfe99720_8090,
        RIfe995b8_8089,RIde83168_229,RIfcc43e8_7255,RIfcd5a58_7453,RIfc89450_6584,RIfcc5798_7269,RIe16c890_2612,RIe16a568_2587,RIe168d80_2570,RIe166788_2543,
        RIe163a88_2511,RIfc83618_6517,RIe160d88_2479,RIee36718_5078,RIe15e088_2447,RIe158688_2383,RIe155988_2351,RIfc3f800_5748,RIe152c88_2319,RIfc895b8_6585,
        RIe14ff88_2287,RIfc51cf8_5953,RIe14d288_2255,RIe14a588_2223,RIe147888_2191,RIee34990_5057,RIee338b0_5045,RIfc831e0_6514,RIfcd3b68_7431,RIe141ff0_2128,
        RIe13fcc8_2103,RIdf3dbd0_2079,RIdf3b740_2053,RIfcb6f90_7104,RIee301d8_5006,RIfcba938_7145,RIee2e018_4982,RIdf369e8_1998,RIdf343f0_1971,RIdf32230_1947,
        RIfe99e28_8095,RIfc83078_6513,RIfcb6e28_7103,RIfc9ad90_6784,RIfcbad70_7148,RIdf2b1b0_1867,RIdf292c0_1845,RIfe99b58_8093,RIfe999f0_8092,RIfc9ac28_6783,
        RIfc4a9a8_5871,RIdf23758_1780,RIfc82da8_6511,RIdf220d8_1764,RIdf20a58_1748,RIdf1ba30_1691,RIfe99cc0_8094,RIdf18358_1652,RIdf15658_1620,RIdf12958_1588,
        RIdf0fc58_1556,RIdf0cf58_1524,RIdf0a258_1492,RIdf07558_1460,RIdf04858_1428,RIdefee58_1364,RIdefc158_1332,RIdef9458_1300,RIdef6758_1268,RIdef3a58_1236,
        RIdef0d58_1204,RIdeee058_1172,RIdeeb358_1140,RIee25918_4886,RIee24b08_4876,RIfc52568_5959,RIfc826a0_6506,RIdee5958_1076,RIdee3bd0_1055,RIfe99f90_8096,
        RIdedf9b8_1008,RIfce4800_7622,RIfc89b58_6589,RIfc9f3e0_6834,RIfc82538_6505,RIdeda828_950,RIded8398_924,RIfeabe70_8272,RIded3eb0_875,RIded1b88_850,
        RIdecee88_818,RIdecc188_786,RIdec9488_754,RIdeb5988_530,RIde99710_338,RIe16f590_2644,RIe15b388_2415,RIe144b88_2159,RIdf39580_2029,RIdf2dbe0_1897,
        RIdf1e460_1721,RIdf01b58_1396,RIdee8658_1108,RIdedd3c0_981,RIde7f658_211,RIe19ea20_3182,RIe19bd20_3150,RIf145928_5251,RIe199020_3118,RIfe98910_8080,
        RIe196320_3086,RIe193620_3054,RIe190920_3022,RIe18af20_2958,RIe188220_2926,RIf143e70_5232,RIe185520_2894,RIfc95c00_6726,RIe182820_2862,RIe17fb20_2830,
        RIe17ce20_2798,RIf142520_5214,RIf141440_5202,RIe1776f0_2736,RIfeab8d0_8268,RIfcc5bd0_7272,RIfc62dc8_6147,RIee3e710_5169,RIfc9cb18_6805,RIee3c820_5147,
        RIee3b470_5133,RIee3a390_5121,RIe174888_2703,RIf170498_5737,RIfc68660_6210,RIf16e878_5717,RIfc6ea38_6281,RIfe98d48_8083,RIe224d78_4709,RIf16c280_5690,
        RIe222078_4677,RIf16b308_5679,RIe21f378_4645,RIe219978_4581,RIe216c78_4549,RIf16a390_5668,RIe213f78_4517,RIf169b20_5662,RIe211278_4485,RIf1681d0_5644,
        RIe20e578_4453,RIe20b878_4421,RIe208b78_4389,RIfcd4ae0_7442,RIfc61478_6129,RIfeab060_8262,RIe201990_4308,RIfc70ec8_6307,RIfc70928_6303,RIfcec528_7711,
        RIfcbe880_7190,RIf160d18_5561,RIf15ee28_5539,RIfe98be0_8082,RIfe98eb0_8084,RIf15d0a0_5518,RIf15bcf0_5504,RIfcd4540_7438,RIf159e00_5482,RIf1592c0_5474,
        RIf158078_5461,RIfca3a30_6884,RIfea7988_8223,RIf156728_5443,RIf155be8_5435,RIf154b08_5423,RIfe98a78_8081,RIf1538c0_5410,RIf1520d8_5393,RIf150e90_5380,
        RIe1f43d0_4156,RIf14fdb0_5368,RIfcd2380_7414,RIf14e2f8_5349,RIe1ef240_4098,RIe1ecae0_4070,RIe1e9de0_4038,RIe1e70e0_4006,RIe1e43e0_3974,RIe1e16e0_3942,
        RIe1de9e0_3910,RIe1dbce0_3878,RIe1d8fe0_3846,RIe1d35e0_3782,RIe1d08e0_3750,RIe1cdbe0_3718,RIe1caee0_3686,RIe1c81e0_3654,RIe1c54e0_3622,RIe1c27e0_3590,
        RIe1bfae0_3558,RIfc44b70_5804,RIf14bd00_5322,RIfe992e8_8087,RIfe987a8_8079,RIf14a950_5308,RIf149f78_5301,RIfe99180_8086,RIfe98640_8078,RIf149438_5293,
        RIfcec7f8_7713,RIfe984d8_8077,RIe1b1b48_3399,RIfc4b650_5880,RIfcda918_7509,RIfe98370_8076,RIfe99018_8085,RIe1a9e20_3310,RIe1a7120_3278,RIe1a4420_3246,
        RIe1a1720_3214,RIe18dc20_2990,RIe17a120_2766,RIe227a78_4741,RIe21c678_4613,RIe205e78_4357,RIe1ffed8_4289,RIe1f9290_4212,RIe1f1dd8_4129,RIe1d62e0_3814,
        RIe1bcde0_3526,RIe1afc58_3377,RIe172290_2676,RIdec6620_721,RIdec3920_689,RIfc49328_5855,RIdec0c20_657,RIfc80eb8_6489,RIdebdf20_625,RIdebb220_593,
        RIdeb8520_561,RIfc80648_6483,RIdeb2b20_497,RIfc8b340_6606,RIdeafe20_465,RIfc491c0_5854,RIdeacec8_433,RIdea65c8_401,RIde9fcc8_369,RIfcd9c70_7500,
        RIfe98208_8075,RIfce4698_7621,RIfe980a0_8074,RIde93158_307,RIde8f648_289,RIde8b4a8_269,RIde87308_249,RIde82e20_228,RIfcbba18_7157,RIfc48d88_5851,
        RIfc99f80_6774,RIfc8b4a8_6607,RIe16c728_2611,RIe16a400_2586,RIe168c18_2569,RIe166620_2542,RIe163920_2510,RIee38068_5096,RIe160c20_2478,RIfc48248_5843,
        RIe15df20_2446,RIe158520_2382,RIe155820_2350,RIfcbbe50_7160,RIe152b20_2318,RIfc47e10_5840,RIe14fe20_2286,RIfca0e98_6853,RIe14d120_2254,RIe14a420_2222,
        RIe147720_2190,RIfc8be80_6614,RIfc7fb08_6475,RIfc480e0_5842,RIfc99878_6769,RIe141e88_2127,RIe13fb60_2102,RIdf3da68_2078,RIdf3b5d8_2052,RIfe97f38_8073,
        RIee30070_5005,RIee2eb58_4990,RIee2deb0_4981,RIdf36880_1997,RIdf34288_1970,RIdf320c8_1946,RIfe97dd0_8072,RIfcc3740_7246,RIfc48ab8_5849,RIfce05e8_7575,
        RIfc80210_6480,RIdf2b048_1866,RIdf29158_1844,RIdf26f98_1820,RIdf254e0_1801,RIfc8bbb0_6612,RIfc48950_5848,RIdf235f0_1779,RIfc8bd18_6613,RIdf21f70_1763,
        RIdf208f0_1747,RIdf1b8c8_1690,RIdf1a3b0_1675,RIdf181f0_1651,RIdf154f0_1619,RIdf127f0_1587,RIdf0faf0_1555,RIdf0cdf0_1523,RIdf0a0f0_1491,RIdf073f0_1459,
        RIdf046f0_1427,RIdefecf0_1363,RIdefbff0_1331,RIdef92f0_1299,RIdef65f0_1267,RIdef38f0_1235,RIdef0bf0_1203,RIdeedef0_1171,RIdeeb1f0_1139,RIfcbc120_7162,
        RIfcd9838_7497,RIfc99710_6768,RIfca1168_6855,RIdee57f0_1075,RIdee3a68_1054,RIdee18a8_1030,RIdedf850_1007,RIfc549f8_5985,RIfcb5370_7084,RIfce43c8_7619,
        RIfce0480_7574,RIdeda6c0_949,RIded8230_923,RIded6070_899,RIded3d48_874,RIded1a20_849,RIdeced20_817,RIdecc020_785,RIdec9320_753,RIdeb5820_529,
        RIde993c8_337,RIe16f428_2643,RIe15b220_2414,RIe144a20_2158,RIdf39418_2028,RIdf2da78_1896,RIdf1e2f8_1720,RIdf019f0_1395,RIdee84f0_1107,RIdedd258_980,
        RIde7f310_210,RIe19e8b8_3181,RIe19bbb8_3149,RIfe976c8_8067,RIe198eb8_3117,RIf144c80_5242,RIe1961b8_3085,RIe1934b8_3053,RIe1907b8_3021,RIe18adb8_2957,
        RIe1880b8_2925,RIfe97560_8066,RIe1853b8_2893,RIfcc3fb0_7252,RIe1826b8_2861,RIe17f9b8_2829,RIe17ccb8_2797,RIfcd3730_7428,RIf1412d8_5201,RIfcc4118_7253,
        RIfe97830_8068,RIfc4a6d8_5869,RIf13f6b8_5181,RIfc9f980_6838,RIfc9fae8_6839,RIfcc3e48_7251,RIfc89e28_6591,RIfc89cc0_6590,RIe174720_2702,RIfc4a408_5867,
        RIfce27a8_7599,RIfc530a8_5967,RIfcd5d28_7455,RIf16cf28_5699,RIe224c10_4708,RIfc53210_5968,RIe221f10_4676,RIf16b1a0_5678,RIe21f210_4644,RIe219810_4580,
        RIe216b10_4548,RIfc401d8_5755,RIe213e10_4516,RIf1699b8_5661,RIe211110_4484,RIfc81cc8_6499,RIe20e410_4452,RIe20b710_4420,RIe208a10_4388,RIfc8a0f8_6593,
        RIfcb6720_7098,RIe203448_4327,RIe201828_4307,RIfc53378_5969,RIfc8a3c8_6595,RIfcb65b8_7097,RIfc49fd0_5864,RIf160bb0_5560,RIf15ecc0_5538,RIe1fd4a8_4259,
        RIfe97b00_8070,RIfc8a530_6596,RIfe97c68_8071,RIfc8a800_6598,RIfc8a698_6597,RIfc9a7f0_6780,RIfc81890_6496,RIfcd5e90_7456,RIe1fb180_4234,RIfc49e68_5863,
        RIfc81728_6495,RIfcbb1a8_7151,RIe1f66f8_4181,RIfcd3460_7426,RIfcb62e8_7095,RIfc9a520_6778,RIe1f4268_4155,RIfc49d00_5862,RIfcd9dd8_7501,RIfcbb310_7152,
        RIe1ef0d8_4097,RIe1ec978_4069,RIe1e9c78_4037,RIe1e6f78_4005,RIe1e4278_3973,RIe1e1578_3941,RIe1de878_3909,RIe1dbb78_3877,RIe1d8e78_3845,RIe1d3478_3781,
        RIe1d0778_3749,RIe1cda78_3717,RIe1cad78_3685,RIe1c8078_3653,RIe1c5378_3621,RIe1c2678_3589,RIe1bf978_3557,RIfc49a30_5860,RIfcb6018_7093,RIe1ba3b0_3496,
        RIe1b81f0_3472,RIfce0a20_7578,RIfcbb5e0_7154,RIe1b6030_3448,RIfe97998_8069,RIfce5610_7632,RIfcc3a10_7248,RIe1b3330_3416,RIe1b19e0_3398,RIfc495f8_5857,
        RIfc81188_6491,RIe1ad228_3347,RIe1aba40_3330,RIe1a9cb8_3309,RIe1a6fb8_3277,RIe1a42b8_3245,RIe1a15b8_3213,RIe18dab8_2989,RIe179fb8_2765,RIe227910_4740,
        RIe21c510_4612,RIe205d10_4356,RIe1ffd70_4288,RIe1f9128_4211,RIe1f1c70_4128,RIe1d6178_3813,RIe1bcc78_3525,RIe1afaf0_3376,RIe172128_2675,RIdec6a58_724,
        RIdec3d58_692,RIfc723e0_6322,RIdec1058_660,RIfc59fc0_6046,RIdebe358_628,RIdebb658_596,RIdeb8958_564,RIfcb96f0_7132,RIdeb2f58_500,RIfce1c68_7591,
        RIdeb0258_468,RIfc9b498_6789,RIdead558_436,RIdea6fa0_404,RIdea06a0_372,RIfc81458_6493,RIfc83780_6518,RIfc4e620_5914,RIfcd3e38_7433,RIde937e8_309,
        RIde8f990_290,RIde8bb38_271,RIde87650_250,RIde834b0_230,RIfc42c80_5782,RIfc65960_6178,RIfc6c710_6256,RIee392b0_5109,RIe16cb60_2614,RIe16a6d0_2588,
        RIe169050_2572,RIe166a58_2545,RIe163d58_2513,RIfec3cf0_8348,RIe161058_2481,RIfcd54b8_7449,RIe15e358_2449,RIe158958_2385,RIe155c58_2353,RIfe9ba48_8115,
        RIe152f58_2321,RIfec4128_8351,RIe150258_2289,RIfcb9b28_7135,RIe14d558_2257,RIe14a858_2225,RIe147b58_2193,RIfcdb2f0_7516,RIfc553d0_5992,RIfc9a0e8_6775,
        RIfcbd908_7179,RIe1422c0_2130,RIe13ff98_2105,RIdf3dea0_2081,RIdf3ba10_2055,RIfc87128_6559,RIee304a8_5008,RIfcc51f8_7265,RIee2e2e8_4984,RIdf36cb8_2000,
        RIfec3fc0_8350,RIdf32500_1949,RIfec3e58_8349,RIee2c830_4965,RIee2ad78_4946,RIee296f8_4930,RIee284b0_4917,RIfe9b8e0_8114,RIfe9b610_8112,RIfe9b778_8113,
        RIfe9b4a8_8111,RIfcb7c38_7113,RIfc86b88_6555,RIdf238c0_1781,RIfc75ab8_6361,RIdf22240_1765,RIfeaa3b8_8253,RIdf1bb98_1692,RIdf1a680_1677,RIdf18628_1654,
        RIdf15928_1622,RIdf12c28_1590,RIdf0ff28_1558,RIdf0d228_1526,RIdf0a528_1494,RIdf07828_1462,RIdf04b28_1430,RIdeff128_1366,RIdefc428_1334,RIdef9728_1302,
        RIdef6a28_1270,RIdef3d28_1238,RIdef1028_1206,RIdeee328_1174,RIdeeb628_1142,RIee25a80_4887,RIee24c70_4877,RIfcddd20_7546,RIfccc110_7344,RIdee5c28_1078,
        RIdee3ea0_1057,RIdee1b78_1032,RIdedfc88_1010,RIfc6a6b8_6233,RIee227e0_4851,RIfc88be0_6578,RIee21868_4840,RIdedaaf8_952,RIded8668_926,RIded6340_901,
        RIded4180_877,RIded1e58_852,RIdecf158_820,RIdecc458_788,RIdec9758_756,RIdeb5c58_532,RIde99da0_340,RIe16f860_2646,RIe15b658_2417,RIe144e58_2161,
        RIdf39850_2031,RIdf2deb0_1899,RIdf1e730_1723,RIdf01e28_1398,RIdee8928_1110,RIdedd690_983,RIde7fce8_213,RIe19ecf0_3184,RIe19bff0_3152,RIf145a90_5252,
        RIe1992f0_3120,RIf144de8_5243,RIe1965f0_3088,RIe1938f0_3056,RIe190bf0_3024,RIe18b1f0_2960,RIe1884f0_2928,RIfc72980_6326,RIe1857f0_2896,RIf143060_5222,
        RIe182af0_2864,RIe17fdf0_2832,RIe17d0f0_2800,RIf142688_5215,RIf141710_5204,RIe177858_2737,RIe176778_2725,RIfcea638_7689,RIfca54e8_6903,RIee3e878_5170,
        RIee3dbd0_5161,RIee3c988_5148,RIee3b5d8_5134,RIee3a4f8_5122,RIe174b58_2705,RIf170600_5738,RIfc76fd0_6376,RIf16e9e0_5718,RIfced608_7723,RIf16d090_5700,
        RIe225048_4711,RIf16c550_5692,RIe222348_4679,RIf16b470_5680,RIe21f648_4647,RIe219c48_4583,RIe216f48_4551,RIf16a4f8_5669,RIe214248_4519,RIf169df0_5664,
        RIe211548_4487,RIf1684a0_5646,RIe20e848_4455,RIe20bb48_4423,RIe208e48_4391,RIf1673c0_5634,RIf166448_5623,RIfe9c6f0_8124,RIfe9c150_8120,RIf1654d0_5612,
        RIfcc4550_7256,RIf1635e0_5590,RIf162500_5578,RIf160fe8_5563,RIf15f0f8_5541,RIfe9bfe8_8119,RIfe9c588_8123,RIf15d208_5519,RIf15bfc0_5506,RIfc4d540_5902,
        RIfc9c848_6803,RIfec4290_8352,RIfe9c2b8_8121,RIfcc01d0_7208,RIe1fb2e8_4235,RIfe9c420_8122,RIfca3e68_6887,RIf154c70_5424,RIe1f69c8_4183,RIf153a28_5411,
        RIf152240_5394,RIf150ff8_5381,RIe1f46a0_4158,RIfca6028_6911,RIfc43bf8_5793,RIf14e460_5350,RIe1ef3a8_4099,RIe1ecdb0_4072,RIe1ea0b0_4040,RIe1e73b0_4008,
        RIe1e46b0_3976,RIe1e19b0_3944,RIe1decb0_3912,RIe1dbfb0_3880,RIe1d92b0_3848,RIe1d38b0_3784,RIe1d0bb0_3752,RIe1cdeb0_3720,RIe1cb1b0_3688,RIe1c84b0_3656,
        RIe1c57b0_3624,RIe1c2ab0_3592,RIe1bfdb0_3560,RIfc4d6a8_5903,RIf14be68_5323,RIe1ba680_3498,RIfe9be80_8118,RIfc86e58_6557,RIfcd46a8_7439,RIe1b6300_3450,
        RIfe9bd18_8117,RIf1495a0_5294,RIf1481f0_5280,RIe1b3600_3418,RIe1b1e18_3401,RIfc69470_6220,RIfcbfac8_7203,RIfe9bbb0_8116,RIe1abd10_3332,RIe1aa0f0_3312,
        RIe1a73f0_3280,RIe1a46f0_3248,RIe1a19f0_3216,RIe18def0_2992,RIe17a3f0_2768,RIe227d48_4743,RIe21c948_4615,RIe206148_4359,RIe2001a8_4291,RIe1f9560_4214,
        RIe1f20a8_4131,RIe1d65b0_3816,RIe1bd0b0_3528,RIe1aff28_3379,RIe172560_2678,RIdec68f0_723,RIdec3bf0_691,RIee208f0_4829,RIdec0ef0_659,RIfc7ce08_6443,
        RIdebe1f0_627,RIdebb4f0_595,RIdeb87f0_563,RIfc9b8d0_6792,RIdeb2df0_499,RIfcc6710_7280,RIdeb00f0_467,RIfc5ff60_6114,RIdead3f0_435,RIdea6c58_403,
        RIdea0358_371,RIfce5070_7628,RIee1c6d8_4782,RIfce70c8_7651,RIee1b058_4766,RIde934a0_308,RIfe9b1d8_8109,RIde8b7f0_270,RIfe9b340_8110,RIfc6b798_6245,
        RIfcb2238_7049,RIfcd3a00_7430,RIfcdb020_7514,RIfc511b8_5945,RIe16c9f8_2613,RIfcb27d8_7053,RIe168ee8_2571,RIe1668f0_2544,RIe163bf0_2512,RIee381d0_5097,
        RIe160ef0_2480,RIfcdfaa8_7567,RIe15e1f0_2448,RIe1587f0_2384,RIe155af0_2352,RIfc3f968_5749,RIe152df0_2320,RIfcd5080_7446,RIe1500f0_2288,RIfc84b30_6532,
        RIe14d3f0_2256,RIe14a6f0_2224,RIe1479f0_2192,RIfcea098_7685,RIfc92f00_6694,RIfc54890_5984,RIfcdcc40_7534,RIe142158_2129,RIe13fe30_2104,RIdf3dd38_2080,
        RIdf3b8a8_2054,RIfc57590_6016,RIee30340_5007,RIfcd0490_7392,RIee2e180_4983,RIdf36b50_1999,RIdf34558_1972,RIdf32398_1948,RIfe9b070_8108,RIfcb1860_7042,
        RIfca1b40_6862,RIfc5c018_6069,RIfe9ada0_8106,RIdf2b318_1868,RIdf29428_1846,RIdf27100_1821,RIfe9af08_8107,RIfc5e1d8_6093,RIfcdcda8_7535,RIfcac400_6982,
        RIfc691a0_6218,RIfcaad80_6966,RIdf20bc0_1749,RIfc61b80_6134,RIdf1a518_1676,RIdf184c0_1653,RIdf157c0_1621,RIdf12ac0_1589,RIdf0fdc0_1557,RIdf0d0c0_1525,
        RIdf0a3c0_1493,RIdf076c0_1461,RIdf049c0_1429,RIdefefc0_1365,RIdefc2c0_1333,RIdef95c0_1301,RIdef68c0_1269,RIdef3bc0_1237,RIdef0ec0_1205,RIdeee1c0_1173,
        RIdeeb4c0_1141,RIfc69b78_6225,RIfc6b900_6246,RIfc4d270_5900,RIfced770_7724,RIdee5ac0_1077,RIdee3d38_1056,RIdee1a10_1031,RIdedfb20_1009,RIfc7ff40_6478,
        RIfca4408_6891,RIfcb5640_7086,RIee21700_4839,RIdeda990_951,RIded8500_925,RIded61d8_900,RIded4018_876,RIded1cf0_851,RIdeceff0_819,RIdecc2f0_787,
        RIdec95f0_755,RIdeb5af0_531,RIde99a58_339,RIe16f6f8_2645,RIe15b4f0_2416,RIe144cf0_2160,RIdf396e8_2030,RIdf2dd48_1898,RIdf1e5c8_1722,RIdf01cc0_1397,
        RIdee87c0_1109,RIdedd528_982,RIde7f9a0_212,RIe19eb88_3183,RIe19be88_3151,RIfe9a698_8101,RIe199188_3119,RIfe9a530_8100,RIe196488_3087,RIe193788_3055,
        RIe190a88_3023,RIe18b088_2959,RIe188388_2927,RIfe9a800_8102,RIe185688_2895,RIfc8d938_6633,RIe182988_2863,RIe17fc88_2831,RIe17cf88_2799,RIfe9a3c8_8099,
        RIf1415a8_5203,RIfe9a260_8098,RIfe9a0f8_8097,RIfcb9150_7128,RIf13f820_5182,RIfc9fc50_6840,RIfce5340_7630,RIfc5cb58_6077,RIfc576f8_6017,RIfc780b0_6388,
        RIe1749f0_2704,RIfc7adb0_6420,RIfc7c2c8_6435,RIfcb2d78_7057,RIfc7e758_6461,RIfe9aad0_8104,RIe224ee0_4710,RIf16c3e8_5691,RIe2221e0_4678,RIfcd3898_7429,
        RIe21f4e0_4646,RIe219ae0_4582,RIe216de0_4550,RIfc880a0_6570,RIe2140e0_4518,RIf169c88_5663,RIe2113e0_4486,RIf168338_5645,RIe20e6e0_4454,RIe20b9e0_4422,
        RIe208ce0_4390,RIfce4c38_7625,RIfc9c6e0_6802,RIe2035b0_4328,RIe201af8_4309,RIfc500d8_5933,RIfc85c10_6544,RIfce81a8_7663,RIfce9c60_7682,RIf160e80_5562,
        RIf15ef90_5540,RIfe9a968_8103,RIfe9ac38_8105,RIfca8d28_6943,RIf15be58_5505,RIfcedba8_7727,RIfc6a988_6235,RIfc71cd8_6317,RIfccb198_7333,RIfcaa3a8_6959,
        RIfec3b88_8347,RIfc4c730_5892,RIfc6d688_6267,RIfca8e90_6944,RIe1f6860_4182,RIfc64e20_6170,RIfcaee30_7012,RIfccee10_7376,RIe1f4538_4157,RIfc63ea8_6159,
        RIfcaecc8_7011,RIfcae458_7005,RIfeab1c8_8263,RIe1ecc48_4071,RIe1e9f48_4039,RIe1e7248_4007,RIe1e4548_3975,RIe1e1848_3943,RIe1deb48_3911,RIe1dbe48_3879,
        RIe1d9148_3847,RIe1d3748_3783,RIe1d0a48_3751,RIe1cdd48_3719,RIe1cb048_3687,RIe1c8348_3655,RIe1c5648_3623,RIe1c2948_3591,RIe1bfc48_3559,RIfcc70e8_7287,
        RIfca7ae0_6930,RIe1ba518_3497,RIe1b8358_3473,RIfc598b8_6041,RIfcc2228_7231,RIe1b6198_3449,RIe1b4848_3431,RIfc82f10_6512,RIfc55970_5996,RIe1b3498_3417,
        RIe1b1cb0_3400,RIfcb7698_7109,RIfc4b4e8_5879,RIe1ad390_3348,RIe1abba8_3331,RIe1a9f88_3311,RIe1a7288_3279,RIe1a4588_3247,RIe1a1888_3215,RIe18dd88_2991,
        RIe17a288_2767,RIe227be0_4742,RIe21c7e0_4614,RIe205fe0_4358,RIe200040_4290,RIe1f93f8_4213,RIe1f1f40_4130,RIe1d6448_3815,RIe1bcf48_3527,RIe1afdc0_3378,
        RIe1723f8_2677,RIdec6d28_726,RIdec4028_694,RIee20bc0_4831,RIdec1328_662,RIfcbaed8_7149,RIdebe628_630,RIdebb928_598,RIdeb8c28_566,RIfc412b8_5767,
        RIdeb3228_502,RIfc9ea08_6827,RIdeb0528_470,RIee1e028_4800,RIdead828_438,RIdea7630_406,RIdea0d30_374,RIfcbac08_7147,RIfc55538_5993,RIfcba668_7143,
        RIfc4af48_5875,RIfe912f0_7996,RIfe91458_7997,RIde8be80_272,RIde87ce0_252,RIfc85238_6537,RIfc88640_6574,RIfcda210_7504,RIfcd5788_7451,RIee39418_5110,
        RIe16ce30_2616,RIfc884d8_6573,RIe169320_2574,RIe166d28_2547,RIe164028_2515,RIfe90918_7989,RIe161328_2483,RIee36880_5079,RIe15e628_2451,RIe158c28_2387,
        RIe155f28_2355,RIfe91188_7995,RIe153228_2323,RIfe91020_7994,RIe150528_2291,RIfcda378_7505,RIe14d828_2259,RIe14ab28_2227,RIe147e28_2195,RIfe90eb8_7993,
        RIfe90d50_7992,RIfcb99c0_7134,RIfc9c2a8_6799,RIfe90be8_7991,RIfe90a80_7990,RIdf3e008_2082,RIdf3bce0_2057,RIfcec690_7712,RIee30778_5010,RIfc87dd0_6568,
        RIee2e5b8_4986,RIdf36e20_2001,RIdf346c0_1973,RIdf32668_1950,RIdf30070_1923,RIee2c998_4966,RIee2aee0_4947,RIee299c8_4932,RIee28618_4918,RIfe90378_7985,
        RIfe907b0_7988,RIfe904e0_7986,RIfe90648_7987,RIfc9d928_6815,RIfc86048_6547,RIfcb92b8_7129,RIfc4ee90_5920,RIfc86a20_6554,RIdf20e90_1751,RIfcb8fe8_7127,
        RIdf1a950_1679,RIdf188f8_1656,RIdf15bf8_1624,RIdf12ef8_1592,RIdf101f8_1560,RIdf0d4f8_1528,RIdf0a7f8_1496,RIdf07af8_1464,RIdf04df8_1432,RIdeff3f8_1368,
        RIdefc6f8_1336,RIdef99f8_1304,RIdef6cf8_1272,RIdef3ff8_1240,RIdef12f8_1208,RIdeee5f8_1176,RIdeeb8f8_1144,RIfc857d8_6541,RIee24dd8_4878,RIfc4ff70_5932,
        RIfc50240_5934,RIdee5ef8_1080,RIdee4170_1059,RIfe915c0_7998,RIdedff58_1012,RIfcd4810_7440,RIee22948_4852,RIfce1560_7586,RIee219d0_4841,RIdedac60_953,
        RIfe91728_7999,RIded64a8_902,RIfe91890_8000,RIded2128_854,RIdecf428_822,RIdecc728_790,RIdec9a28_758,RIdeb5f28_534,RIde9a430_342,RIe16fb30_2648,
        RIe15b928_2419,RIe145128_2163,RIdf39b20_2033,RIdf2e180_1901,RIdf1ea00_1725,RIdf020f8_1400,RIdee8bf8_1112,RIdedd960_985,RIde80378_215,RIe19efc0_3186,
        RIe19c2c0_3154,RIf145d60_5254,RIe1995c0_3122,RIfc637a0_6154,RIe1968c0_3090,RIe193bc0_3058,RIe190ec0_3026,RIe18b4c0_2962,RIe1887c0_2930,RIfc62af8_6145,
        RIe185ac0_2898,RIfe8fc70_7980,RIe182dc0_2866,RIe1800c0_2834,RIe17d3c0_2802,RIfe90210_7984,RIfe8ff40_7982,RIfc72f20_6330,RIe176a48_2727,RIfcaf6a0_7018,
        RIfc61040_6126,RIf13e8a8_5171,RIfe900a8_7983,RIee3caf0_5149,RIee3b740_5135,RIee3a660_5123,RIe174e28_2707,RIf170768_5739,RIfc5fdf8_6113,RIf16eb48_5719,
        RIfcaaab0_6964,RIf16d1f8_5701,RIe225318_4713,RIf16c6b8_5693,RIe222618_4681,RIf16b5d8_5681,RIe21f918_4649,RIe219f18_4585,RIe217218_4553,RIfca62f8_6913,
        RIe214518_4521,RIfcc9578_7313,RIe211818_4489,RIfca5a88_6907,RIe20eb18_4457,RIe20be18_4425,RIe209118_4393,RIf167690_5636,RIf166718_5625,RIfe8f9a0_7978,
        RIfe8f838_7977,RIf165638_5613,RIf164990_5604,RIf1638b0_5592,RIf1627d0_5580,RIf161150_5564,RIf15f260_5542,RIe1fd778_4261,RIe1fc530_4248,RIf15d4d8_5521,
        RIf15c290_5508,RIfca20e0_6866,RIf159f68_5483,RIf159428_5475,RIf1581e0_5462,RIfc5ebb0_6100,RIfe8fdd8_7981,RIfc69e48_6227,RIfc5e8e0_6098,RIf154f40_5426,
        RIe1f6b30_4184,RIf153b90_5412,RIf1523a8_5395,RIfce88b0_7668,RIfe8fb08_7979,RIfcebe20_7706,RIfcb1158_7037,RIf14e730_5352,RIe1ef678_4101,RIe1ed080_4074,
        RIe1ea380_4042,RIe1e7680_4010,RIe1e4980_3978,RIe1e1c80_3946,RIe1def80_3914,RIe1dc280_3882,RIe1d9580_3850,RIe1d3b80_3786,RIe1d0e80_3754,RIe1ce180_3722,
        RIe1cb480_3690,RIe1c8780_3658,RIe1c5a80_3626,RIe1c2d80_3594,RIe1c0080_3562,RIfcc8ba0_7306,RIfc5d698_6085,RIfec35e8_8343,RIfeabd08_8271,RIfc5cf90_6080,
        RIfc5ce28_6079,RIfec31b0_8340,RIe1b4b18_3433,RIf149708_5295,RIf148358_5281,RIe1b3768_3419,RIfec3480_8342,RIfc483b0_5844,RIfc80be8_6487,RIe1ad4f8_3349,
        RIfec3318_8341,RIe1aa3c0_3314,RIe1a76c0_3282,RIe1a49c0_3250,RIe1a1cc0_3218,RIe18e1c0_2994,RIe17a6c0_2770,RIe228018_4745,RIe21cc18_4617,RIe206418_4361,
        RIe200478_4293,RIe1f9830_4216,RIe1f2378_4133,RIe1d6880_3818,RIe1bd380_3530,RIe1b01f8_3381,RIe172830_2680,RIdec6bc0_725,RIdec3ec0_693,RIee20a58_4830,
        RIdec11c0_661,RIee1f978_4818,RIdebe4c0_629,RIdebb7c0_597,RIdeb8ac0_565,RIee1efa0_4811,RIdeb30c0_501,RIfcb04b0_7028,RIdeb03c0_469,RIfc5e4a8_6095,
        RIdead6c0_437,RIdea72e8_405,RIdea09e8_373,RIfcb2508_7051,RIfcd16d8_7405,RIfc5d800_6086,RIfc63d40_6158,RIde93b30_310,RIfea7820_8222,RIfea73e8_8219,
        RIde87998_251,RIde837f8_231,RIfc7bd28_6431,RIfcc7ef8_7297,RIfc7a108_6411,RIfc7a6a8_6415,RIe16ccc8_2615,RIe16a838_2589,RIe1691b8_2573,RIe166bc0_2546,
        RIe163ec0_2514,RIee38338_5098,RIe1611c0_2482,RIfc54b60_5986,RIe15e4c0_2450,RIe158ac0_2386,RIe155dc0_2354,RIee35a70_5069,RIe1530c0_2322,RIee357a0_5067,
        RIe1503c0_2290,RIfc9fdb8_6841,RIe14d6c0_2258,RIe14a9c0_2226,RIe147cc0_2194,RIee34af8_5058,RIee33a18_5046,RIee327d0_5033,RIfcbcf30_7172,RIe142428_2131,
        RIe140100_2106,RIfea7280_8218,RIdf3bb78_2056,RIfc731f0_6332,RIee30610_5009,RIfcbe010_7184,RIee2e450_4985,RIfec2ee0_8338,RIfec3048_8339,RIfec2c10_8336,
        RIfec2d78_8337,RIfcb46c8_7075,RIfcb4830_7076,RIee29860_4931,RIfcb88e0_7122,RIdf2b480_1869,RIdf29590_1847,RIdf27268_1822,RIdf25648_1802,RIfcc9de8_7319,
        RIfc53648_5971,RIdf23a28_1782,RIfc823d0_6504,RIdf223a8_1766,RIdf20d28_1750,RIdf1bd00_1693,RIdf1a7e8_1678,RIdf18790_1655,RIdf15a90_1623,RIdf12d90_1591,
        RIdf10090_1559,RIdf0d390_1527,RIdf0a690_1495,RIdf07990_1463,RIdf04c90_1431,RIdeff290_1367,RIdefc590_1335,RIdef9890_1303,RIdef6b90_1271,RIdef3e90_1239,
        RIdef1190_1207,RIdeee490_1175,RIdeeb790_1143,RIee25be8_4888,RIfc6af28_6239,RIee23fc8_4868,RIfccf680_7382,RIdee5d90_1079,RIdee4008_1058,RIdee1ce0_1033,
        RIdedfdf0_1011,RIfc6b090_6240,RIfc534e0_5970,RIfca5920_6906,RIfc66770_6188,RIfe8f6d0_7976,RIded87d0_927,RIfe8f568_7975,RIded42e8_878,RIded1fc0_853,
        RIdecf2c0_821,RIdecc5c0_789,RIdec98c0_757,RIdeb5dc0_533,RIde9a0e8_341,RIe16f9c8_2647,RIe15b7c0_2418,RIe144fc0_2162,RIdf399b8_2032,RIdf2e018_1900,
        RIdf1e898_1724,RIdf01f90_1399,RIdee8a90_1111,RIdedd7f8_984,RIde80030_214,RIe19ee58_3185,RIe19c158_3153,RIf145bf8_5253,RIe199458_3121,RIfe8f298_7973,
        RIe196758_3089,RIe193a58_3057,RIe190d58_3025,RIe18b358_2961,RIe188658_2929,RIfe8f130_7972,RIe185958_2897,RIfc9f278_6833,RIe182c58_2865,RIe17ff58_2833,
        RIe17d258_2801,RIf1427f0_5216,RIfe8efc8_7971,RIe1779c0_2738,RIe1768e0_2726,RIfc81e30_6500,RIfc9ff20_6842,RIfca0088_6843,RIfc81b60_6498,RIfce5778_7633,
        RIfce08b8_7577,RIfc815c0_6494,RIe174cc0_2706,RIfca04c0_6846,RIfc53eb8_5977,RIfcc65a8_7279,RIfc80d50_6488,RIfc804e0_6482,RIe2251b0_4712,RIfc80378_6481,
        RIe2224b0_4680,RIfcb5910_7088,RIe21f7b0_4648,RIe219db0_4584,RIe2170b0_4552,RIfca01f0_6844,RIe2143b0_4520,RIfc82c40_6510,RIe2116b0_4488,RIfc7f6d0_6472,
        RIe20e9b0_4456,RIe20bcb0_4424,RIe208fb0_4392,RIf167528_5635,RIf1665b0_5624,RIe203718_4329,RIe201c60_4310,RIfc9da90_6816,RIfcc5360_7266,RIf163748_5591,
        RIf162668_5579,RIfc7e320_6458,RIfc87998_6565,RIe1fd610_4260,RIe1fc3c8_4247,RIf15d370_5520,RIf15c128_5507,RIfcc5d38_7273,RIfce7d70_7660,RIfc4bd58_5885,
        RIfc55c40_5998,RIfca2ab8_6873,RIe1fb450_4236,RIf156890_5444,RIfcd5ff8_7457,RIf154dd8_5425,RIfec2aa8_8335,RIfcb4b00_7078,RIfcd9400_7494,RIf151160_5382,
        RIe1f4808_4159,RIfc44738_5801,RIfc90908_6667,RIf14e5c8_5351,RIe1ef510_4100,RIe1ecf18_4073,RIe1ea218_4041,RIe1e7518_4009,RIe1e4818_3977,RIe1e1b18_3945,
        RIe1dee18_3913,RIe1dc118_3881,RIe1d9418_3849,RIe1d3a18_3785,RIe1d0d18_3753,RIe1ce018_3721,RIe1cb318_3689,RIe1c8618_3657,RIe1c5918_3625,RIe1c2c18_3593,
        RIe1bff18_3561,RIf14d218_5337,RIfe8ee60_7970,RIfea8090_8228,RIe1b84c0_3474,RIf14aab8_5309,RIfc6c170_6252,RIe1b6468_3451,RIe1b49b0_3432,RIfcafad8_7021,
        RIfcaa948_6963,RIfe8ecf8_7969,RIfe8f400_7974,RIfc67f58_6205,RIfca8ff8_6945,RIfe8eb90_7968,RIe1abe78_3333,RIe1aa258_3313,RIe1a7558_3281,RIe1a4858_3249,
        RIe1a1b58_3217,RIe18e058_2993,RIe17a558_2769,RIe227eb0_4744,RIe21cab0_4616,RIe2062b0_4360,RIe200310_4292,RIe1f96c8_4215,RIe1f2210_4132,RIe1d6718_3817,
        RIe1bd218_3529,RIe1b0090_3380,RIe1726c8_2679,RIdec4460_697,RIdec1760_665,RIee1fae0_4819,RIdebea60_633,RIee1f108_4812,RIdebbd60_601,RIdeb9060_569,
        RIdeb6360_537,RIee1eb68_4808,RIdeb0960_473,RIee1e460_4803,RIdeadc60_441,RIee1d7b8_4794,RIdea8008_409,RIdea1708_377,RIde9ae08_345,RIfe957d8_8045,
        RIfe95508_8043,RIfe95670_8044,RIee1a7e8_4760,RIfe95aa8_8047,RIfe95238_8041,RIfe95940_8046,RIfe953a0_8042,RIee1a0e0_4755,RIee19ca8_4752,RIee19870_4749,
        RIee19438_4746,RIee38ba8_5104,RIfe95c10_8048,RIee384a0_5099,RIfea9440_8242,RIe164460_2518,RIe161760_2486,RIfe942c0_8030,RIe15ea60_2454,RIfe94158_8029,
        RIe15bd60_2422,RIe156360_2358,RIe153660_2326,RIfe94428_8031,RIe150960_2294,RIfe94590_8032,RIe14dc60_2262,RIfc5c2e8_6071,RIe14af60_2230,RIe148260_2198,
        RIe145560_2166,RIee33ce8_5048,RIee32aa0_5035,RIee31858_5022,RIfc5d530_6084,RIe140538_2109,RIdf3e2d8_2084,RIdf3c118_2060,RIdf39df0_2035,RIfcdd780_7542,
        RIee2ee28_4992,RIfcc88d0_7304,RIee2cc68_4968,RIdf34990_1975,RIdf32aa0_1953,RIdf304a8_1926,RIdf2e5b8_1904,RIee2b1b0_4949,RIfe946f8_8033,RIfcb2940_7054,
        RIee273d0_4905,RIfe949c8_8035,RIdf27538_1824,RIfe94b30_8036,RIfe94860_8034,RIee26f98_4902,RIee269f8_4898,RIee26728_4896,RIee26458_4894,RIee26188_4892,
        RIfe94c98_8037,RIee25d50_4889,RIfea9170_8240,RIdf16030_1627,RIdf13330_1595,RIdf10630_1563,RIdf0d930_1531,RIdf0ac30_1499,RIdf07f30_1467,RIdf05230_1435,
        RIdf02530_1403,RIdefcb30_1339,RIdef9e30_1307,RIdef7130_1275,RIdef4430_1243,RIdef1730_1211,RIdeeea30_1179,RIdeebd30_1147,RIdee9030_1115,RIee250a8_4880,
        RIee24298_4870,RIee23758_4862,RIee22d80_4855,RIfe950d0_8040,RIfe94f68_8039,RIfe94e00_8038,RIdeddd98_988,RIee22ab0_4853,RIee21e08_4844,RIfca46d8_6893,
        RIfc5dad0_6088,RIfeaa250_8252,RIfe96048_8051,RIfe95d78_8049,RIfe95ee0_8050,RIdecf860_825,RIdeccb60_793,RIdec9e60_761,RIdec7160_729,RIdeb3660_505,
        RIde94508_313,RIe16d268_2619,RIe159060_2390,RIe142860_2134,RIdf37258_2004,RIdf2b8b8_1872,RIdf1c138_1696,RIdeff830_1371,RIdee6330_1083,RIdedb098_956,
        RIde7a450_186,RIe19c6f8_3157,RIe1999f8_3125,RIf1450b8_5245,RIe196cf8_3093,RIf143fd8_5233,RIe193ff8_3061,RIe1912f8_3029,RIe18e5f8_2997,RIe188bf8_2933,
        RIe185ef8_2901,RIfe973f8_8065,RIe1831f8_2869,RIf142958_5217,RIe1804f8_2837,RIe17d7f8_2805,RIe17aaf8_2773,RIf141b48_5207,RIfc542f0_5980,RIfc800a8_6479,
        RIe175260_2710,RIfca0bc8_6851,RIfc48680_5846,RIee3dea0_5163,RIfcc6878_7281,RIee3ba10_5137,RIee3a930_5125,RIfe97290_8064,RIe172b00_2682,RIf16f958_5729,
        RIf16ee18_5721,RIf16da68_5707,RIf16d360_5702,RIfe96e58_8061,RIe222a50_4684,RIfe96cf0_8060,RIe21fd50_4652,RIf16a660_5670,RIe21d050_4620,RIe217650_4556,
        RIe214950_4524,RIf169f58_5665,RIe211c50_4492,RIf168770_5648,RIe20ef50_4460,RIf1677f8_5637,RIe20c250_4428,RIe209550_4396,RIe206850_4364,RIf166880_5626,
        RIf1657a0_5614,RIe201dc8_4311,RIe2005e0_4294,RIfe96b88_8059,RIf163b80_5594,RIf162c08_5583,RIf161420_5566,RIf15f530_5544,RIf15d7a8_5523,RIfe968b8_8057,
        RIfe96a20_8058,RIfcb3fc0_7070,RIfc7cf70_6444,RIfc579c8_6019,RIf159590_5476,RIf1584b0_5464,RIf157268_5451,RIf1569f8_5445,RIfe965e8_8055,RIf155d50_5436,
        RIf155210_5428,RIf153e60_5414,RIfe96750_8056,RIf1527e0_5398,RIf151430_5384,RIfcd2650_7416,RIe1f2648_4135,RIf14f108_5359,RIfc7f298_6469,RIf14d4e8_5339,
        RIe1ed350_4076,RIe1ea7b8_4045,RIe1e7ab8_4013,RIe1e4db8_3981,RIe1e20b8_3949,RIe1df3b8_3917,RIe1dc6b8_3885,RIe1d99b8_3853,RIe1d6cb8_3821,RIe1d12b8_3757,
        RIe1ce5b8_3725,RIe1cb8b8_3693,RIe1c8bb8_3661,RIe1c5eb8_3629,RIe1c31b8_3597,RIe1c04b8_3565,RIe1bd7b8_3533,RIf14c138_5325,RIf14ad88_5311,RIe1b8790_3476,
        RIfe96480_8054,RIf14a0e0_5302,RIf149870_5296,RIfe97128_8063,RIfe96318_8053,RIf148628_5283,RIfc58d78_6033,RIe1b20e8_3403,RIe1b04c8_3383,RIf146cd8_5265,
        RIfc591b0_6036,RIfe961b0_8052,RIfe96fc0_8062,RIe1a7af8_3285,RIe1a4df8_3253,RIe1a20f8_3221,RIe19f3f8_3189,RIe18b8f8_2965,RIe177df8_2741,RIe225750_4716,
        RIe21a350_4588,RIe203b50_4332,RIe1fdbb0_4264,RIe1f6f68_4187,RIe1efab0_4104,RIe1d3fb8_3789,RIe1baab8_3501,RIe1ad930_3352,RIe16ff68_2651,RIdec42f8_696,
        RIdec15f8_664,RIfcc6cb0_7284,RIdebe8f8_632,RIfe93780_8022,RIdebbbf8_600,RIdeb8ef8_568,RIdeb61f8_536,RIee1ea00_4807,RIdeb07f8_472,RIee1e2f8_4802,
        RIdeadaf8_440,RIfc5d3c8_6083,RIdea7cc0_408,RIdea13c0_376,RIde9aac0_344,RIfc58238_6025,RIfcc3b78_7249,RIfc7d0d8_6445,RIfc59750_6040,RIfe93a50_8024,
        RIfe938e8_8023,RIde88370_254,RIde83e88_233,RIfc5f420_6106,RIfc976b8_6745,RIfc90a70_6668,RIfc60500_6118,RIee38a40_5103,RIe16ab08_2591,RIe169488_2575,
        RIe166ff8_2549,RIe1642f8_2517,RIe1615f8_2485,RIee369e8_5080,RIe15e8f8_2453,RIee35bd8_5070,RIe15bbf8_2421,RIe1561f8_2357,RIe1534f8_2325,RIfc3ee28_5741,
        RIe1507f8_2293,RIfce6c90_7648,RIe14daf8_2261,RIfcca7c0_7326,RIe14adf8_2229,RIe1480f8_2197,RIe1453f8_2165,RIee33b80_5047,RIee32938_5034,RIee316f0_5021,
        RIee30bb0_5013,RIe1403d0_2108,RIfe93618_8021,RIdf3bfb0_2059,RIfe934b0_8020,RIfcd0d00_7398,RIee2ecc0_4991,RIee2e720_4987,RIee2cb00_4967,RIfe93bb8_8025,
        RIdf32938_1952,RIdf30340_1925,RIdf2e450_1903,RIee2b048_4948,RIee29b30_4933,RIfc67148_6195,RIfc6fb18_6293,RIdf29860_1849,RIfe931e0_8018,RIfe93348_8019,
        RIfe93078_8017,RIfc672b0_6196,RIfca8788_6939,RIdf22510_1767,RIfcea7a0_7690,RIdf20ff8_1752,RIdf1ecd0_1727,RIdf1aab8_1680,RIfea7c58_8225,RIdf15ec8_1626,
        RIdf131c8_1594,RIdf104c8_1562,RIdf0d7c8_1530,RIdf0aac8_1498,RIdf07dc8_1466,RIdf050c8_1434,RIdf023c8_1402,RIdefc9c8_1338,RIdef9cc8_1306,RIdef6fc8_1274,
        RIdef42c8_1242,RIdef15c8_1210,RIdeee8c8_1178,RIdeebbc8_1146,RIdee8ec8_1114,RIee24f40_4879,RIee24130_4869,RIee235f0_4861,RIee22c18_4854,RIfe93d20_8026,
        RIdee1fb0_1035,RIdee0228_1014,RIdeddc30_987,RIfc684f8_6209,RIee21ca0_4843,RIfc68390_6208,RIee20d28_4832,RIded8aa0_929,RIfe93ff0_8028,RIded45b8_880,
        RIfe93e88_8027,RIdecf6f8_824,RIdecc9f8_792,RIdec9cf8_760,RIdec6ff8_728,RIdeb34f8_504,RIde941c0_312,RIe16d100_2618,RIe158ef8_2389,RIe1426f8_2133,
        RIdf370f0_2003,RIdf2b750_1871,RIdf1bfd0_1695,RIdeff6c8_1370,RIdee61c8_1082,RIdedaf30_955,RIde7a108_185,RIe19c590_3156,RIe199890_3124,RIf144f50_5244,
        RIe196b90_3092,RIfc76058_6365,RIe193e90_3060,RIe191190_3028,RIe18e490_2996,RIe188a90_2932,RIe185d90_2900,RIfccd8f8_7361,RIe183090_2868,RIfc76e68_6375,
        RIe180390_2836,RIe17d690_2804,RIe17a990_2772,RIf1419e0_5206,RIf140630_5192,RIe176bb0_2728,RIe1750f8_2709,RIfcd1840_7406,RIfc5f6f0_6108,RIee3dd38_5162,
        RIee3cc58_5150,RIee3b8a8_5136,RIee3a7c8_5124,RIee39580_5111,RIfea9008_8239,RIf16f7f0_5728,RIf16ecb0_5720,RIf16d900_5706,RIfc78ec0_6398,RIfcc8060_7298,
        RIe2228e8_4683,RIfc5a3f8_6049,RIe21fbe8_4651,RIfc74000_6342,RIe21cee8_4619,RIe2174e8_4555,RIe2147e8_4523,RIfca2c20_6874,RIe211ae8_4491,RIfca2950_6872,
        RIe20ede8_4459,RIfcc24f8_7233,RIe20c0e8_4427,RIe2093e8_4395,RIe2066e8_4363,RIfc45110_5808,RIfcc6f80_7286,RIfe92f10_8016,RIfe92970_8012,RIf164af8_5605,
        RIf163a18_5593,RIf162aa0_5582,RIfe92ad8_8013,RIf15f3c8_5543,RIf15d640_5522,RIfe92808_8011,RIfe92c40_8014,RIfe926a0_8010,RIfe92da8_8015,RIfe92538_8009,
        RIfcb5a78_7089,RIf158348_5463,RIf157100_5450,RIfc53be8_5975,RIfec38b8_8345,RIfcc5ea0_7274,RIf1550a8_5427,RIf153cf8_5413,RIfec3a20_8346,RIf152678_5397,
        RIfec3750_8344,RIf14ff18_5369,RIfe923d0_8008,RIf14efa0_5358,RIf14e898_5353,RIf14d380_5338,RIfe92268_8007,RIe1ea650_4044,RIe1e7950_4012,RIe1e4c50_3980,
        RIe1e1f50_3948,RIe1df250_3916,RIe1dc550_3884,RIe1d9850_3852,RIe1d6b50_3820,RIe1d1150_3756,RIe1ce450_3724,RIe1cb750_3692,RIe1c8a50_3660,RIe1c5d50_3628,
        RIe1c3050_3596,RIe1c0350_3564,RIe1bd650_3532,RIfcda4e0_7506,RIfc9d220_6810,RIe1b8628_3475,RIe1b6738_3453,RIfc4f2c8_5923,RIfce16c8_7587,RIfe91cc8_8003,
        RIfe91e30_8004,RIf1484c0_5282,RIf147548_5271,RIfe91f98_8005,RIfe91b60_8002,RIf146b70_5264,RIfc9f548_6835,RIfe92100_8006,RIfe919f8_8001,RIe1a7990_3284,
        RIe1a4c90_3252,RIe1a1f90_3220,RIe19f290_3188,RIe18b790_2964,RIe177c90_2740,RIe2255e8_4715,RIe21a1e8_4587,RIe2039e8_4331,RIe1fda48_4263,RIe1f6e00_4186,
        RIe1ef948_4103,RIe1d3e50_3788,RIe1ba950_3500,RIe1ad7c8_3351,RIe16fe00_2650,RIdec4730_699,RIdec1a30_667,RIfce3f90_7616,RIdebed30_635,RIfcc3308_7243,
        RIdebc030_603,RIdeb9330_571,RIdeb6630_539,RIfc8c588_6619,RIdeb0c30_475,RIfc5a998_6053,RIdeadf30_443,RIfc99b48_6771,RIdea8698_411,RIdea1d98_379,
        RIde9b498_347,RIfc78bf0_6396,RIfcbc558_7165,RIfca12d0_6856,RIfca3fd0_6888,RIfec2670_8332,RIfec2508_8331,RIde88a00_256,RIde84518_235,RIfcc35d8_7245,
        RIfcb57a8_7087,RIfc5a290_6048,RIfca3058_6877,RIee38e78_5106,RIfec27d8_8333,RIfca3328_6879,RIe1672c8_2551,RIe164730_2520,RIe161a30_2488,RIee36cb8_5082,
        RIe15ed30_2456,RIfcc7250_7288,RIe15c030_2424,RIe156630_2360,RIe153930_2328,RIfcc7688_7291,RIe150c30_2296,RIfc8af08_6603,RIe14df30_2264,RIfc9a250_6776,
        RIe14b230_2232,RIe148530_2200,RIe145830_2168,RIfc9aac0_6782,RIfc56bb8_6009,RIfca1ca8_6863,RIfcec960_7714,RIe1406a0_2110,RIdf3e440_2085,RIdf3c280_2061,
        RIdf39f58_2036,RIfc9a958_6781,RIee2f0f8_4994,RIfcdb458_7517,RIee2cf38_4970,RIdf34c60_1977,RIfec2940_8334,RIdf30778_1928,RIdf2e888_1906,RIee2b480_4951,
        RIfec23a0_8330,RIee288e8_4920,RIfec2238_8329,RIdf29b30_1851,RIdf27808_1826,RIdf25a80_1805,RIdf23e60_1785,RIfc55100_5990,RIfcd9f40_7502,RIfc54f98_5989,
        RIfc54cc8_5987,RIfc4b218_5877,RIdf1efa0_1729,RIfcc69e0_7282,RIdf18bc8_1658,RIdf16300_1629,RIdf13600_1597,RIdf10900_1565,RIdf0dc00_1533,RIdf0af00_1501,
        RIdf08200_1469,RIdf05500_1437,RIdf02800_1405,RIdefce00_1341,RIdefa100_1309,RIdef7400_1277,RIdef4700_1245,RIdef1a00_1213,RIdeeed00_1181,RIdeec000_1149,
        RIdee9300_1117,RIfce4ad0_7624,RIfc9e8a0_6826,RIfcc46b8_7257,RIfcd4108_7435,RIdee4440_1061,RIdee2280_1037,RIdee0390_1015,RIdede068_990,RIfcda0a8_7503,
        RIfce54a8_7631,RIfca0790_6848,RIfc50ee8_5943,RIded8d70_931,RIded68e0_905,RIded4888_882,RIded2560_857,RIdecfb30_827,RIdecce30_795,RIdeca130_763,
        RIdec7430_731,RIdeb3930_507,RIde94b98_315,RIe16d538_2621,RIe159330_2392,RIe142b30_2136,RIdf37528_2006,RIdf2bb88_1874,RIdf1c408_1698,RIdeffb00_1373,
        RIdee6600_1085,RIdedb368_958,RIde7aae0_188,RIe19c9c8_3159,RIe199cc8_3127,RIfe8ea28_7967,RIe196fc8_3095,RIfec20d0_8328,RIe1942c8_3063,RIe1915c8_3031,
        RIe18e8c8_2999,RIe188ec8_2935,RIe1861c8_2903,RIfc68228_6207,RIe1834c8_2871,RIfccb5d0_7336,RIe1807c8_2839,RIe17dac8_2807,RIe17adc8_2775,RIf141e18_5209,
        RIf140900_5194,RIf140090_5188,RIe1753c8_2711,RIf13f988_5183,RIf13ece0_5174,RIee3e170_5165,RIee3cf28_5152,RIee3bce0_5139,RIee3ac00_5127,RIee39850_5113,
        RIe172dd0_2684,RIf16fc28_5731,RIf16f0e8_5723,RIf16dd38_5709,RIfce9120_7674,RIfc404a8_5757,RIe222d20_4686,RIf16b8a8_5683,RIe220020_4654,RIf16a930_5672,
        RIe21d320_4622,RIe217920_4558,RIe214c20_4526,RIfc5b910_6064,RIe211f20_4494,RIfe8e8c0_7966,RIe20f220_4462,RIfe8e758_7965,RIe20c520_4430,RIe209820_4398,
        RIe206b20_4366,RIf166b50_5628,RIf165a70_5616,RIfe8dd80_7958,RIfe8dab0_7956,RIf164c60_5606,RIf163e50_5596,RIf162ed8_5585,RIf1616f0_5568,RIf15f800_5546,
        RIf15da78_5525,RIfe8d948_7955,RIfe8dc18_7957,RIf15c560_5510,RIf15b048_5495,RIfc62828_6143,RIf159860_5478,RIf158780_5466,RIf157538_5453,RIfca6e38_6921,
        RIe1f9b00_4218,RIfc61e50_6136,RIfc61748_6131,RIf154130_5416,RIe1f4ad8_4161,RIf152ab0_5400,RIf151700_5386,RIf1501e8_5371,RIe1f27b0_4136,RIfc60ed8_6125,
        RIfc7b620_6426,RIf14d7b8_5341,RIe1ed4b8_4077,RIe1eaa88_4047,RIe1e7d88_4015,RIe1e5088_3983,RIe1e2388_3951,RIe1df688_3919,RIe1dc988_3887,RIe1d9c88_3855,
        RIe1d6f88_3823,RIe1d1588_3759,RIe1ce888_3727,RIe1cbb88_3695,RIe1c8e88_3663,RIe1c6188_3631,RIe1c3488_3599,RIe1c0788_3567,RIe1bda88_3535,RIfca4de0_6898,
        RIfc5ea48_6099,RIe1b8a60_3478,RIe1b6a08_3455,RIfcbd638_7177,RIfc44fa8_5807,RIfe8e5f0_7964,RIfe8e1b8_7961,RIf1488f8_5285,RIf147818_5273,RIfe8e050_7960,
        RIfe8e488_7963,RIf146e40_5266,RIf146030_5256,RIfe8dee8_7959,RIfe8e320_7962,RIe1a7dc8_3287,RIe1a50c8_3255,RIe1a23c8_3223,RIe19f6c8_3191,RIe18bbc8_2967,
        RIe1780c8_2743,RIe225a20_4718,RIe21a620_4590,RIe203e20_4334,RIe1fde80_4266,RIe1f7238_4189,RIe1efd80_4106,RIe1d4288_3791,RIe1bad88_3503,RIe1adc00_3354,
        RIe170238_2653,RIdec45c8_698,RIdec18c8_666,RIfce85e0_7666,RIdebebc8_634,RIfcb8bb0_7124,RIdebbec8_602,RIdeb91c8_570,RIdeb64c8_538,RIfc85d78_6545,
        RIdeb0ac8_474,RIfc85aa8_6543,RIdeaddc8_442,RIfc4d3d8_5901,RIdea8350_410,RIdea1a50_378,RIde9b150_346,RIfc85ee0_6546,RIfc9c9b0_6804,RIfce13f8_7585,
        RIfcb8778_7121,RIfe8d510_7952,RIfe8d3a8_7951,RIde886b8_255,RIde841d0_234,RIde806c0_216,RIfcb8070_7116,RIfce1128_7583,RIfc9c140_6798,RIee38d10_5105,
        RIe16ac70_2592,RIfc850d0_6536,RIe167160_2550,RIe1645c8_2519,RIe1618c8_2487,RIee36b50_5081,RIe15ebc8_2455,RIee35d40_5071,RIe15bec8_2423,RIe1564c8_2359,
        RIe1537c8_2327,RIfc3ef90_5742,RIe150ac8_2295,RIfe8d7e0_7954,RIe14ddc8_2263,RIfce0fc0_7582,RIe14b0c8_2231,RIe1483c8_2199,RIe1456c8_2167,RIee33e50_5049,
        RIee32c08_5036,RIee319c0_5023,RIee30d18_5014,RIfe8cf70_7948,RIfe8ce08_7947,RIfe8d240_7950,RIfe8d0d8_7949,RIfce9dc8_7683,RIee2ef90_4993,RIfce51d8_7629,
        RIee2cdd0_4969,RIdf34af8_1976,RIfe8d678_7953,RIdf30610_1927,RIdf2e720_1905,RIee2b318_4950,RIee29c98_4934,RIee28780_4919,RIee27538_4906,RIdf299c8_1850,
        RIdf276a0_1825,RIdf25918_1804,RIdf23cf8_1784,RIfc83ff0_6524,RIfcb73c8_7107,RIfc51320_5946,RIfcdaa80_7510,RIfc83d20_6522,RIdf1ee38_1728,RIfc51b90_5952,
        RIdf18a60_1657,RIdf16198_1628,RIdf13498_1596,RIdf10798_1564,RIdf0da98_1532,RIdf0ad98_1500,RIdf08098_1468,RIdf05398_1436,RIdf02698_1404,RIdefcc98_1340,
        RIdef9f98_1308,RIdef7298_1276,RIdef4598_1244,RIdef1898_1212,RIdeeeb98_1180,RIdeebe98_1148,RIdee9198_1116,RIee25210_4881,RIee24400_4871,RIee238c0_4863,
        RIee22ee8_4856,RIfe8cca0_7946,RIdee2118_1036,RIfe8cb38_7945,RIdeddf00_989,RIfcc5a68_7271,RIee21f70_4845,RIfcb6cc0_7102,RIee20e90_4833,RIded8c08_930,
        RIded6778_904,RIded4720_881,RIded23f8_856,RIdecf9c8_826,RIdecccc8_794,RIdec9fc8_762,RIdec72c8_730,RIdeb37c8_506,RIde94850_314,RIe16d3d0_2620,
        RIe1591c8_2391,RIe1429c8_2135,RIdf373c0_2005,RIdf2ba20_1873,RIdf1c2a0_1697,RIdeff998_1372,RIdee6498_1084,RIdedb200_957,RIde7a798_187,RIe19c860_3158,
        RIe199b60_3126,RIf145220_5246,RIe196e60_3094,RIf144140_5234,RIe194160_3062,RIe191460_3030,RIe18e760_2998,RIe188d60_2934,RIe186060_2902,RIf1431c8_5223,
        RIe183360_2870,RIf142ac0_5218,RIe180660_2838,RIe17d960_2806,RIe17ac60_2774,RIf141cb0_5208,RIf140798_5193,RIf13ff28_5187,RIfe8be90_7936,RIfceb880_7702,
        RIf13eb78_5173,RIee3e008_5164,RIee3cdc0_5151,RIee3bb78_5138,RIee3aa98_5126,RIee396e8_5112,RIe172c68_2683,RIf16fac0_5730,RIf16ef80_5722,RIf16dbd0_5708,
        RIfcc4af0_7260,RIf16c820_5694,RIe222bb8_4685,RIf16b740_5682,RIe21feb8_4653,RIf16a7c8_5671,RIe21d1b8_4621,RIe2177b8_4557,RIe214ab8_4525,RIfe8c430_7940,
        RIe211db8_4493,RIf1688d8_5649,RIe20f0b8_4461,RIf167960_5638,RIe20c3b8_4429,RIe2096b8_4397,RIe2069b8_4365,RIf1669e8_5627,RIf165908_5615,RIfe8c9d0_7944,
        RIfe8c700_7942,RIfc9c578_6801,RIf163ce8_5595,RIf162d70_5584,RIf161588_5567,RIf15f698_5545,RIf15d910_5524,RIfe8c598_7941,RIfe8c868_7943,RIf15c3f8_5509,
        RIf15aee0_5494,RIf15a0d0_5484,RIf1596f8_5477,RIf158618_5465,RIf1573d0_5452,RIf156b60_5446,RIfec1f68_8327,RIf155eb8_5437,RIf155378_5429,RIf153fc8_5415,
        RIfe8bff8_7937,RIf152948_5399,RIf151598_5385,RIf150080_5370,RIfe8c2c8_7939,RIf14f270_5360,RIfc503a8_5935,RIf14d650_5340,RIfe8c160_7938,RIe1ea920_4046,
        RIe1e7c20_4014,RIe1e4f20_3982,RIe1e2220_3950,RIe1df520_3918,RIe1dc820_3886,RIe1d9b20_3854,RIe1d6e20_3822,RIe1d1420_3758,RIe1ce720_3726,RIe1cba20_3694,
        RIe1c8d20_3662,RIe1c6020_3630,RIe1c3320_3598,RIe1c0620_3566,RIe1bd920_3534,RIf14c2a0_5326,RIf14aef0_5312,RIe1b88f8_3477,RIe1b68a0_3454,RIfcd4db0_7444,
        RIfc4ebc0_5918,RIfec1e00_8326,RIfe8bd28_7935,RIf148790_5284,RIf1476b0_5272,RIfe8ba58_7933,RIfec1b30_8324,RIfc4e788_5915,RIfcb8e80_7126,RIfe8bbc0_7934,
        RIfec1c98_8325,RIe1a7c60_3286,RIe1a4f60_3254,RIe1a2260_3222,RIe19f560_3190,RIe18ba60_2966,RIe177f60_2742,RIe2258b8_4717,RIe21a4b8_4589,RIe203cb8_4333,
        RIe1fdd18_4265,RIe1f70d0_4188,RIe1efc18_4105,RIe1d4120_3790,RIe1bac20_3502,RIe1ada98_3353,RIe1700d0_2652,RIdec4a00_701,RIdec1d00_669,RIfcad7b0_6996,
        RIdebf000_637,RIfc64cb8_6169,RIdebc300_605,RIdeb9600_573,RIdeb6900_541,RIfc6f9b0_6292,RIdeb0f00_477,RIfc657f8_6177,RIdeae200_445,RIfce69c0_7646,
        RIdea8d28_413,RIdea2428_381,RIde9bb28_349,RIfc6fc80_6294,RIee1b760_4771,RIfca8080_6934,RIfe8b8f0_7932,RIde90020_292,RIde8c510_274,RIde89090_258,
        RIde84ba8_237,RIfc65ac8_6179,RIfcad210_6992,RIfcce168_7367,RIfcce2d0_7368,RIfc51488_5947,RIe16af40_2594,RIfc65c30_6180,RIe167598_2553,RIe164a00_2522,
        RIe161d00_2490,RIfc66e78_6193,RIe15f000_2458,RIfc6e498_6277,RIe15c300_2426,RIe156900_2362,RIe153c00_2330,RIfc6e330_6276,RIe150f00_2298,RIfccda60_7362,
        RIe14e200_2266,RIfc6e1c8_6275,RIe14b500_2234,RIe148800_2202,RIe145b00_2170,RIee33fb8_5050,RIee32d70_5037,RIee31c90_5025,RIee30fe8_5016,RIfea8630_8232,
        RIdf3e5a8_2086,RIdf3c550_2063,RIfea8798_8233,RIfc6e060_6274,RIfcac6d0_6984,RIfc56078_6001,RIfc6e600_6278,RIdf34dc8_1978,RIdf32d70_1955,RIfea84c8_8231,
        RIdf2eb58_1908,RIee2b750_4953,RIfc6ee70_6284,RIfc6efd8_6285,RIee27808_4908,RIfe8b788_7931,RIdf27ad8_1828,RIdf25d50_1807,RIdf24130_1787,RIfc66608_6187,
        RIfccde98_7365,RIfc66a40_6190,RIfc668d8_6189,RIfcacf40_6990,RIfeaaef8_8261,RIfc6e8d0_6280,RIdf18d30_1659,RIdf165d0_1631,RIdf138d0_1599,RIdf10bd0_1567,
        RIdf0ded0_1535,RIdf0b1d0_1503,RIdf084d0_1471,RIdf057d0_1439,RIdf02ad0_1407,RIdefd0d0_1343,RIdefa3d0_1311,RIdef76d0_1279,RIdef49d0_1247,RIdef1cd0_1215,
        RIdeeefd0_1183,RIdeec2d0_1151,RIdee95d0_1119,RIfc6dc28_6271,RIfc67c88_6203,RIfccb300_7334,RIfccd4c0_7358,RIfea81f8_8229,RIfea8360_8230,RIdee04f8_1016,
        RIdede338_992,RIfc6def8_6273,RIfcac130_6980,RIfc67b20_6202,RIfc67df0_6204,RIded9040_933,RIded6a48_906,RIded4b58_884,RIded26c8_858,RIdecfe00_829,
        RIdecd100_797,RIdeca400_765,RIdec7700_733,RIdeb3c00_509,RIde95228_317,RIe16d808_2623,RIe159600_2394,RIe142e00_2138,RIdf377f8_2008,RIdf2be58_1876,
        RIdf1c6d8_1700,RIdeffdd0_1375,RIdee68d0_1087,RIdedb638_960,RIde7b170_190,RIe19cc98_3161,RIe199f98_3129,RIfc73088_6331,RIe197298_3097,RIf1442a8_5235,
        RIe194598_3065,RIe191898_3033,RIe18eb98_3001,RIe189198_2937,RIe186498_2905,RIfc72278_6321,RIe183798_2873,RIfc61ce8_6135,RIe180a98_2841,RIe17dd98_2809,
        RIe17b098_2777,RIfcaf268_7015,RIfca6a00_6918,RIfcc9b18_7317,RIe175530_2712,RIfc72818_6325,RIfc726b0_6324,RIfccf7e8_7383,RIfc72548_6323,RIee3be48_5140,
        RIee3ad68_5128,RIfc71fa8_6319,RIe1730a0_2686,RIfcaef98_7013,RIfccf518_7381,RIfc71e40_6318,RIfc62120_6138,RIfe8b350_7928,RIe222ff0_4688,RIfcc9f50_7320,
        RIe2202f0_4656,RIfc4a570_5868,RIe21d5f0_4624,RIe217bf0_4560,RIe214ef0_4528,RIfccf3b0_7380,RIe2121f0_4496,RIf168ba8_5651,RIe20f4f0_4464,RIfc71300_6310,
        RIe20c7f0_4432,RIe209af0_4400,RIe206df0_4368,RIfc718a0_6314,RIfc71a08_6315,RIe202098_4313,RIfe8b1e8_7927,RIfc715d0_6312,RIfce6588_7643,RIfc62c60_6146,
        RIf161858_5569,RIf15fad0_5548,RIf15dbe0_5526,RIe1fc698_4249,RIfe8b4b8_7929,RIfcae5c0_7006,RIfc63098_6149,RIfc63200_6150,RIfc71198_6309,RIf158a50_5468,
        RIf1576a0_5454,RIfcdc808_7531,RIfe8b620_7930,RIfc634d0_6152,RIfcceb40_7374,RIf154400_5418,RIe1f4da8_4163,RIf152c18_5401,RIf151868_5387,RIfc4d108_5899,
        RIe1f2a80_4138,RIfc70a90_6304,RIfc63bd8_6157,RIfca7810_6928,RIe1ed788_4079,RIe1ead58_4049,RIe1e8058_4017,RIe1e5358_3985,RIe1e2658_3953,RIe1df958_3921,
        RIe1dcc58_3889,RIe1d9f58_3857,RIe1d7258_3825,RIe1d1858_3761,RIe1ceb58_3729,RIe1cbe58_3697,RIe1c9158_3665,RIe1c6458_3633,RIe1c3758_3601,RIe1c0a58_3569,
        RIe1bdd58_3537,RIf14c408_5327,RIf14b1c0_5314,RIe1b8d30_3480,RIe1b6cd8_3457,RIfc707c0_6302,RIfca7c48_6931,RIe1b4de8_3435,RIe1b3a38_3421,RIfc70220_6298,
        RIfcce870_7372,RIe1b23b8_3405,RIe1b0630_3384,RIfc645b0_6164,RIfc700b8_6297,RIfeaac28_8259,RIe1aa690_3316,RIe1a8098_3289,RIe1a5398_3257,RIe1a2698_3225,
        RIe19f998_3193,RIe18be98_2969,RIe178398_2745,RIe225cf0_4720,RIe21a8f0_4592,RIe2040f0_4336,RIe1fe150_4268,RIe1f7508_4191,RIe1f0050_4108,RIe1d4558_3793,
        RIe1bb058_3505,RIe1aded0_3356,RIe170508_2655,RIdec4898_700,RIdec1b98_668,RIfc661d0_6184,RIdebee98_636,RIfce6b28_7647,RIdebc198_604,RIdeb9498_572,
        RIdeb6798_540,RIfc40d18_5763,RIdeb0d98_476,RIfcad648_6995,RIdeae098_444,RIfcaa510_6960,RIdea89e0_412,RIdea20e0_380,RIde9b7e0_348,RIfcab320_6970,
        RIfca8350_6936,RIfc6f6e0_6290,RIfcaa240_6958,RIde8fcd8_291,RIfe8aae0_7922,RIde88d48_257,RIde84860_236,RIde80a08_217,RIfc64718_6165,RIfcae020_7002,
        RIfcadeb8_7001,RIee38fe0_5107,RIe16add8_2593,RIe1695f0_2576,RIe167430_2552,RIe164898_2521,RIe161b98_2489,RIfe8a3d8_7917,RIe15ee98_2457,RIfe8a270_7916,
        RIe15c198_2425,RIe156798_2361,RIe153a98_2329,RIfc3f0f8_5743,RIe150d98_2297,RIfcab050_6968,RIe14e098_2265,RIfcca658_7325,RIe14b398_2233,RIe148698_2201,
        RIe145998_2169,RIfe8a810_7920,RIfe8a6a8_7919,RIee31b28_5024,RIee30e80_5015,RIe140808_2111,RIfe8a540_7918,RIdf3c3e8_2062,RIdf3a0c0_2037,RIfc6b1f8_6241,
        RIee2f260_4995,RIfc70d60_6306,RIee2d0a0_4971,RIfe8a978_7921,RIdf32c08_1954,RIdf308e0_1929,RIdf2e9f0_1907,RIee2b5e8_4952,RIee29e00_4935,RIee28a50_4921,
        RIee276a0_4907,RIdf29c98_1852,RIdf27970_1827,RIdf25be8_1806,RIdf23fc8_1786,RIfc6aaf0_6236,RIfc6ac58_6237,RIdf22678_1768,RIfcdd4b0_7540,RIdf21160_1753,
        RIdf1f108_1730,RIdf1ac20_1681,RIfeaa7f0_8256,RIdf16468_1630,RIdf13768_1598,RIdf10a68_1566,RIdf0dd68_1534,RIdf0b068_1502,RIdf08368_1470,RIdf05668_1438,
        RIdf02968_1406,RIdefcf68_1342,RIdefa268_1310,RIdef7568_1278,RIdef4868_1246,RIdef1b68_1214,RIdeeee68_1182,RIdeec168_1150,RIdee9468_1118,RIee25378_4882,
        RIee24568_4872,RIee23a28_4864,RIee23050_4857,RIfe8adb0_7924,RIdee23e8_1038,RIfe8ac48_7923,RIdede1d0_991,RIfca5650_6904,RIee220d8_4846,RIfceeb20_7738,
        RIee20ff8_4834,RIded8ed8_932,RIfe8af18_7925,RIded49f0_883,RIfe8b080_7926,RIdecfc98_828,RIdeccf98_796,RIdeca298_764,RIdec7598_732,RIdeb3a98_508,
        RIde94ee0_316,RIe16d6a0_2622,RIe159498_2393,RIe142c98_2137,RIdf37690_2007,RIdf2bcf0_1875,RIdf1c570_1699,RIdeffc68_1374,RIdee6768_1086,RIdedb4d0_959,
        RIde7ae28_189,RIe19cb30_3160,RIe199e30_3128,RIf145388_5247,RIe197130_3096,RIfe8a108_7915,RIe194430_3064,RIe191730_3032,RIe18ea30_3000,RIe189030_2936,
        RIe186330_2904,RIfc6c878_6257,RIe183630_2872,RIfcabcf8_6977,RIe180930_2840,RIe17dc30_2808,RIe17af30_2776,RIfcccc50_7352,RIfcccdb8_7353,RIe176d18_2729,
        RIfea7af0_8224,RIfe89fa0_7914,RIfe89e38_7913,RIfcdd078_7537,RIfccb738_7337,RIfca9868_6951,RIfcabb90_6976,RIfca99d0_6952,RIe172f38_2685,RIf16fd90_5732,
        RIf16f250_5724,RIfc6c440_6254,RIfcaba28_6975,RIfc40610_5758,RIe222e88_4687,RIfc5d260_6082,RIe220188_4655,RIfcab758_6973,RIe21d488_4623,RIe217a88_4559,
        RIe214d88_4527,RIfe892f8_7905,RIe212088_4495,RIf168a40_5650,RIe20f388_4463,RIf167ac8_5639,RIe20c688_4431,RIe209988_4399,RIe206c88_4367,RIfc6c2d8_6253,
        RIfceec88_7739,RIe201f30_4312,RIe200748_4295,RIf164dc8_5607,RIf163fb8_5597,RIf163040_5586,RIfe895c8_7907,RIf15f968_5547,RIfe89898_7909,RIfe89460_7906,
        RIe1fb5b8_4237,RIf15c6c8_5511,RIfe89730_7908,RIf15a238_5485,RIf1599c8_5479,RIf1588e8_5467,RIfe89cd0_7912,RIfc5ba78_6065,RIe1f9c68_4219,RIfc5bd48_6067,
        RIf1554e0_5430,RIf154298_5417,RIe1f4c40_4162,RIfe89b68_7911,RIfe89a00_7910,RIf150350_5372,RIe1f2918_4137,RIf14f3d8_5361,RIfccc818_7349,RIf14d920_5342,
        RIe1ed620_4078,RIe1eabf0_4048,RIe1e7ef0_4016,RIe1e51f0_3984,RIe1e24f0_3952,RIe1df7f0_3920,RIe1dcaf0_3888,RIe1d9df0_3856,RIe1d70f0_3824,RIe1d16f0_3760,
        RIe1ce9f0_3728,RIe1cbcf0_3696,RIe1c8ff0_3664,RIe1c62f0_3632,RIe1c35f0_3600,RIe1c08f0_3568,RIe1bdbf0_3536,RIfc680c0_6206,RIf14b058_5313,RIe1b8bc8_3479,
        RIe1b6b70_3456,RIfcac298_6981,RIf1499d8_5297,RIfe89190_7904,RIfec19c8_8323,RIf148a60_5286,RIfccdd30_7364,RIe1b2250_3404,RIfec1860_8322,RIfc6e768_6279,
        RIfc54728_5983,RIe1abfe0_3334,RIe1aa528_3315,RIe1a7f30_3288,RIe1a5230_3256,RIe1a2530_3224,RIe19f830_3192,RIe18bd30_2968,RIe178230_2744,RIe225b88_4719,
        RIe21a788_4591,RIe203f88_4335,RIe1fdfe8_4267,RIe1f73a0_4190,RIe1efee8_4107,RIe1d43f0_3792,RIe1baef0_3504,RIe1add68_3355,RIe1703a0_2654,RIdec4cd0_703,
        RIdec1fd0_671,RIfc7b4b8_6425,RIdebf2d0_639,RIfc7b1e8_6423,RIdebc5d0_607,RIdeb98d0_575,RIdeb6bd0_543,RIfe83358_7837,RIdeb11d0_479,RIee1e5c8_4804,
        RIdeae4d0_447,RIfc437c0_5790,RIdea93b8_415,RIdea2ab8_383,RIde9c1b8_351,RIfc90ea8_6671,RIfc7af18_6421,RIfe83088_7835,RIee1a950_4761,RIde906b0_294,
        RIde8cba0_276,RIfe82f20_7834,RIfe82db8_7833,RIee1a248_4756,RIfe831f0_7836,RIfcc2390_7232,RIee195a0_4747,RIfcbe718_7189,RIfea9e18_8249,RIfc43220_5786,
        RIe167868_2555,RIe164cd0_2524,RIe161fd0_2492,RIee36f88_5084,RIe15f2d0_2460,RIee35ea8_5072,RIe15c5d0_2428,RIe156bd0_2364,RIe153ed0_2332,RIfe83628_7839,
        RIe1511d0_2300,RIfebfda8_8303,RIe14e4d0_2268,RIfebfc40_8302,RIe14b7d0_2236,RIe148ad0_2204,RIe145dd0_2172,RIee34120_5051,RIee32ed8_5038,RIee31df8_5026,
        RIfcc1f58_7229,RIe140ad8_2113,RIdf3e878_2088,RIfe834c0_7838,RIdf3a390_2039,RIfc5a6c8_6051,RIfc91e20_6682,RIee2e888_4988,RIfc96a10_6736,RIdf35098_1980,
        RIfeab600_8266,RIdf30bb0_1931,RIfeab768_8267,RIfcbe9e8_7191,RIfc79fa0_6410,RIfc96740_6734,RIfc92258_6685,RIfea7118_8217,RIfea95a8_8243,RIdf26020_1809,
        RIdf24400_1789,RIfc79a00_6406,RIfc5add0_6056,RIfce5d18_7637,RIfc92690_6688,RIfce3018_7605,RIdf1f270_1731,RIfc79730_6404,RIdf19000_1661,RIdf168a0_1633,
        RIdf13ba0_1601,RIdf10ea0_1569,RIdf0e1a0_1537,RIdf0b4a0_1505,RIdf087a0_1473,RIdf05aa0_1441,RIdf02da0_1409,RIdefd3a0_1345,RIdefa6a0_1313,RIdef79a0_1281,
        RIdef4ca0_1249,RIdef1fa0_1217,RIdeef2a0_1185,RIdeec5a0_1153,RIdee98a0_1121,RIfc5b7a8_6063,RIfc5b640_6062,RIfc931d0_6696,RIfcecac8_7715,RIdee4710_1063,
        RIdee26b8_1040,RIdee07c8_1018,RIdede4a0_993,RIfcbf0f0_7196,RIfcbf528_7199,RIfc792f8_6401,RIfc93068_6695,RIded91a8_934,RIded6d18_908,RIded4e28_886,
        RIded2998_860,RIded00d0_831,RIdecd3d0_799,RIdeca6d0_767,RIdec79d0_735,RIdeb3ed0_511,RIde958b8_319,RIe16dad8_2625,RIe1598d0_2396,RIe1430d0_2140,
        RIdf37ac8_2010,RIdf2c128_1878,RIdf1c9a8_1702,RIdf000a0_1377,RIdee6ba0_1089,RIdedb908_962,RIde7b800_192,RIe19cf68_3163,RIe19a268_3131,RIfc8d7d0_6632,
        RIe197568_3099,RIfc561e0_6002,RIe194868_3067,RIe191b68_3035,RIe18ee68_3003,RIe189468_2939,RIe186768_2907,RIf143330_5224,RIe183a68_2875,RIfc7d948_6451,
        RIe180d68_2843,RIe17e068_2811,RIe17b368_2779,RIfc564b0_6004,RIfcd6700_7462,RIfc461f0_5820,RIe175698_2713,RIfc46088_5819,RIfc45f20_5818,RIfc7dc18_6453,
        RIfcd69d0_7464,RIfc98630_6756,RIfcc2a98_7237,RIfc7d510_6448,RIe173208_2687,RIfc8e478_6641,RIfc45ae8_5815,RIfc8e8b0_6644,RIfc45980_5814,RIfe82ae8_7831,
        RIe2232c0_4690,RIf16ba10_5684,RIe2205c0_4658,RIfcd24e8_7415,RIe21d8c0_4626,RIe217ec0_4562,RIe2151c0_4530,RIfebf268_8295,RIe2124c0_4498,RIf168d10_5652,
        RIe20f7c0_4466,RIfc7d240_6446,RIe20cac0_4434,RIe209dc0_4402,RIe2070c0_4370,RIf166e20_5630,RIfebf6a0_8298,RIfebf808_8299,RIfebf538_8297,RIfc8eb80_6646,
        RIf164120_5598,RIfc453e0_5810,RIf161b28_5571,RIf15fc38_5549,RIf15dd48_5527,RIe1fc968_4251,RIe1fb888_4239,RIfebf3d0_8296,RIf15b318_5497,RIfca2518_6869,
        RIfc8f120_6650,RIfebfad8_8301,RIfebf970_8300,RIfc7cca0_6442,RIe1f9dd0_4220,RIfe82c50_7832,RIf155648_5431,RIfc8f288_6651,RIe1f4f10_4164,RIf152d80_5402,
        RIfc8f828_6655,RIfcb3b88_7067,RIe1f2d50_4140,RIfc445d0_5800,RIfc8faf8_6657,RIf14da88_5343,RIe1eda58_4081,RIe1eb028_4051,RIe1e8328_4019,RIe1e5628_3987,
        RIe1e2928_3955,RIe1dfc28_3923,RIe1dcf28_3891,RIe1da228_3859,RIe1d7528_3827,RIe1d1b28_3763,RIe1cee28_3731,RIe1cc128_3699,RIe1c9428_3667,RIe1c6728_3635,
        RIe1c3a28_3603,RIe1c0d28_3571,RIe1be028_3539,RIfc7bff8_6433,RIfc44030_5796,RIe1b9000_3482,RIe1b6fa8_3459,RIfcbdd40_7182,RIfc8ff30_6660,RIe1b50b8_3437,
        RIe1b3d08_3423,RIfcbe178_7185,RIfc43d60_5794,RIe1b2520_3406,RIe1b0798_3385,RIfcdb5c0_7518,RIfc7ba58_6429,RIe1ac148_3335,RIe1aa960_3318,RIe1a8368_3291,
        RIe1a5668_3259,RIe1a2968_3227,RIe19fc68_3195,RIe18c168_2971,RIe178668_2747,RIe225fc0_4722,RIe21abc0_4594,RIe2043c0_4338,RIe1fe420_4270,RIe1f77d8_4193,
        RIe1f0320_4110,RIe1d4828_3795,RIe1bb328_3507,RIe1ae1a0_3358,RIe1707d8_2657,RIdec4b68_702,RIdec1e68_670,RIfc5df08_6091,RIdebf168_638,RIfce6df8_7649,
        RIdebc468_606,RIdeb9768_574,RIdeb6a68_542,RIfc75ef0_6364,RIdeb1068_478,RIfcc12b0_7220,RIdeae368_446,RIfc5e340_6094,RIdea9070_414,RIdea2770_382,
        RIde9be70_350,RIfced4a0_7722,RIfcc1418_7221,RIfc95930_6724,RIfcec0f0_7708,RIde90368_293,RIde8c858_275,RIde893d8_259,RIde84ef0_238,RIde80d50_218,
        RIfc95a98_6725,RIfced068_7719,RIfced1d0_7720,RIfcedfe0_7730,RIe16b0a8_2595,RIe169758_2577,RIe167700_2554,RIe164b68_2523,RIe161e68_2491,RIee36e20_5083,
        RIe15f168_2459,RIfc426e0_5778,RIe15c468_2427,RIe156a68_2363,RIe153d68_2331,RIfe82818_7829,RIe151068_2299,RIee34c60_5059,RIe14e368_2267,RIfc5f9c0_6110,
        RIe14b668_2235,RIe148968_2203,RIe145c68_2171,RIfccfef0_7388,RIfca57b8_6905,RIfc600c8_6115,RIfcafda8_7023,RIe140970_2112,RIdf3e710_2087,RIdf3c6b8_2064,
        RIdf3a228_2038,RIfc5fc90_6112,RIee2f3c8_4996,RIfc742d0_6344,RIee2d208_4972,RIdf34f30_1979,RIfebf100_8294,RIdf30a48_1930,RIdf2ecc0_1909,RIfcb08e8_7031,
        RIfcee418_7733,RIfc95ed0_6728,RIfcdef68_7559,RIdf29e00_1853,RIdf27c40_1829,RIdf25eb8_1808,RIdf24298_1788,RIfc5ed18_6101,RIfcee850_7736,RIdf227e0_1769,
        RIfc5efe8_6103,RIdf212c8_1754,RIfeaa520_8254,RIdf1ad88_1682,RIdf18e98_1660,RIdf16738_1632,RIdf13a38_1600,RIdf10d38_1568,RIdf0e038_1536,RIdf0b338_1504,
        RIdf08638_1472,RIdf05938_1440,RIdf02c38_1408,RIdefd238_1344,RIdefa538_1312,RIdef7838_1280,RIdef4b38_1248,RIdef1e38_1216,RIdeef138_1184,RIdeec438_1152,
        RIdee9738_1120,RIfcc96e0_7314,RIfccfd88_7387,RIfc60aa0_6122,RIfca5ec0_6910,RIdee45a8_1062,RIdee2550_1039,RIdee0660_1017,RIfe826b0_7828,RIfcdeb30_7556,
        RIfc73bc8_6339,RIfca5bf0_6908,RIfc73a60_6338,RIfe82980_7830,RIded6bb0_907,RIded4cc0_885,RIded2830_859,RIdecff68_830,RIdecd268_798,RIdeca568_766,
        RIdec7868_734,RIdeb3d68_510,RIde95570_318,RIe16d970_2624,RIe159768_2395,RIe142f68_2139,RIdf37960_2009,RIdf2bfc0_1877,RIdf1c840_1701,RIdefff38_1376,
        RIdee6a38_1088,RIdedb7a0_961,RIde7b4b8_191,RIe19ce00_3162,RIe19a100_3130,RIfce96c0_7678,RIe197400_3098,RIf144410_5236,RIe194700_3066,RIe191a00_3034,
        RIe18ed00_3002,RIe189300_2938,RIe186600_2906,RIfebee30_8292,RIe183900_2874,RIfcdbcc8_7523,RIe180c00_2842,RIe17df00_2810,RIe17b200_2778,RIf141f80_5210,
        RIfce7398_7653,RIfcb1e00_7046,RIfe82548_7827,RIfca42a0_6890,RIfcbff00_7206,RIfcaaee8_6967,RIee3d090_5153,RIfc5c180_6070,RIfce35b8_7609,RIee399b8_5114,
        RIfea8a68_8235,RIf16fef8_5733,RIfebecc8_8291,RIfc5c450_6072,RIfce9288_7675,RIfc40778_5759,RIe223158_4689,RIfce77d0_7656,RIe220458_4657,RIfce24d8_7597,
        RIe21d758_4625,RIe217d58_4561,RIe215058_4529,RIfce8a18_7669,RIe212358_4497,RIfce1998_7589,RIe20f658_4465,RIfc77840_6382,RIe20c958_4433,RIe209c58_4401,
        RIe206f58_4369,RIf166cb8_5629,RIf165bd8_5617,RIfe81fa8_7823,RIfe81e40_7822,RIfc5c888_6075,RIfceb178_7697,RIf1631a8_5587,RIf1619c0_5570,RIfccf248_7379,
        RIfc77570_6380,RIe1fc800_4250,RIe1fb720_4238,RIf15c830_5512,RIf15b1b0_5496,RIfcd0fd0_7400,RIfccc6b0_7348,RIf158bb8_5469,RIf157808_5455,RIfc5d0f8_6081,
        RIfebef98_8293,RIfcc8a38_7305,RIfcd7ab0_7476,RIfcb1428_7039,RIfeaa0e8_8251,RIfccc548_7347,RIfce3450_7608,RIf1504b8_5373,RIe1f2be8_4139,RIf14f540_5362,
        RIfc772a0_6378,RIfcec258_7709,RIe1ed8f0_4080,RIe1eaec0_4050,RIe1e81c0_4018,RIe1e54c0_3986,RIe1e27c0_3954,RIe1dfac0_3922,RIe1dcdc0_3890,RIe1da0c0_3858,
        RIe1d73c0_3826,RIe1d19c0_3762,RIe1cecc0_3730,RIe1cbfc0_3698,RIe1c92c0_3666,RIe1c65c0_3634,RIe1c38c0_3602,RIe1c0bc0_3570,RIe1bdec0_3538,RIf14c570_5328,
        RIf14b328_5315,RIe1b8e98_3481,RIe1b6e40_3458,RIfc76760_6370,RIfc94b20_6714,RIe1b4f50_3436,RIe1b3ba0_3422,RIfcec3c0_7710,RIfceb010_7696,RIfe823e0_7826,
        RIfe82110_7824,RIfcdd8e8_7543,RIfcc0ba8_7215,RIfe82278_7825,RIe1aa7f8_3317,RIe1a8200_3290,RIe1a5500_3258,RIe1a2800_3226,RIe19fb00_3194,RIe18c000_2970,
        RIe178500_2746,RIe225e58_4721,RIe21aa58_4593,RIe204258_4337,RIe1fe2b8_4269,RIe1f7670_4192,RIe1f01b8_4109,RIe1d46c0_3794,RIe1bb1c0_3506,RIe1ae038_3357,
        RIe170670_2656,RIdec4fa0_705,RIdec22a0_673,RIee1fdb0_4821,RIdebf5a0_641,RIee1f270_4813,RIdebc8a0_609,RIdeb9ba0_577,RIdeb6ea0_545,RIee1ecd0_4809,
        RIdeb14a0_481,RIee1e730_4805,RIdeae7a0_449,RIee1d920_4795,RIdea9a48_417,RIdea3148_385,RIde9c848_353,RIee1cb10_4785,RIee1ba30_4773,RIee1b1c0_4767,
        RIfec04b0_8308,RIfe850e0_7858,RIde8d230_278,RIfea9cb0_8248,RIfe84f78_7857,RIee1a3b0_4757,RIfe853b0_7860,RIee199d8_4750,RIfe85248_7859,RIee39148_5108,
        RIe16b378_2597,RIee38608_5100,RIe167b38_2557,RIe164fa0_2526,RIe1622a0_2494,RIfe85950_7864,RIe15f5a0_2462,RIee36010_5073,RIe15c8a0_2430,RIe156ea0_2366,
        RIe1541a0_2334,RIfe85c20_7866,RIe1514a0_2302,RIee34dc8_5060,RIe14e7a0_2270,RIfc861b0_6548,RIe14baa0_2238,RIe148da0_2206,RIe1460a0_2174,RIee343f0_5053,
        RIfe85518_7861,RIfe857e8_7863,RIfe85680_7862,RIe140c40_2114,RIdf3eb48_2090,RIdf3c820_2065,RIdf3a660_2041,RIfc9d4f0_6812,RIee2f698_4998,RIfc52298_5957,
        RIee2d4d8_4974,RIdf35368_1982,RIdf32ed8_1956,RIdf30e80_1933,RIfe85ab8_7865,RIee2b8b8_4954,RIee29f68_4936,RIee28bb8_4922,RIee27970_4909,RIdf2a0d0_1855,
        RIfe84e10_7856,RIdf262f0_1811,RIfe84ca8_7855,RIee27100_4903,RIee26b60_4899,RIfcd32f8_7425,RIee265c0_4895,RIfc9e300_6822,RIdf1f540_1733,RIee25eb8_4890,
        RIfe84b40_7854,RIdf16b70_1635,RIdf13e70_1603,RIdf11170_1571,RIdf0e470_1539,RIdf0b770_1507,RIdf08a70_1475,RIdf05d70_1443,RIdf03070_1411,RIdefd670_1347,
        RIdefa970_1315,RIdef7c70_1283,RIdef4f70_1251,RIdef2270_1219,RIdeef570_1187,RIdeec870_1155,RIdee9b70_1123,RIfec0348_8307,RIfcb54d8_7085,RIee23cf8_4866,
        RIfc54e30_5988,RIfec0078_8305,RIdee2988_1042,RIfec01e0_8306,RIdede770_995,RIfcd7ee8_7479,RIfcd43d8_7437,RIfc88eb0_6580,RIfc9e5d0_6824,RIded9478_936,
        RIded6fe8_910,RIded50f8_888,RIfeab330_8264,RIded03a0_833,RIdecd6a0_801,RIdeca9a0_769,RIdec7ca0_737,RIdeb41a0_513,RIde95f48_321,RIe16dda8_2627,
        RIe159ba0_2398,RIe1433a0_2142,RIdf37d98_2012,RIdf2c3f8_1880,RIdf1cc78_1704,RIdf00370_1379,RIdee6e70_1091,RIdedbbd8_964,RIde7be90_194,RIe19d238_3165,
        RIe19a538_3133,RIf145658_5249,RIe197838_3101,RIf1446e0_5238,RIe194b38_3069,RIe191e38_3037,RIe18f138_3005,RIe189738_2941,RIe186a38_2909,RIf143600_5226,
        RIe183d38_2877,RIf142c28_5219,RIe181038_2845,RIe17e338_2813,RIe17b638_2781,RIf1420e8_5211,RIf140a68_5195,RIf1401f8_5189,RIfebff10_8304,RIf13faf0_5184,
        RIf13ee48_5175,RIee3e2d8_5166,RIee3d1f8_5154,RIee3c118_5142,RIee3b038_5130,RIee39c88_5116,RIfe838f8_7841,RIf1701c8_5735,RIfc5ab00_6054,RIf16e008_5711,
        RIfcb0e88_7035,RIf16caf0_5696,RIe223590_4692,RIf16bce0_5686,RIe220890_4660,RIf16ac00_5674,RIe21db90_4628,RIe218190_4564,RIe215490_4532,RIf16a228_5667,
        RIe212790_4500,RIf168fe0_5654,RIe20fa90_4468,RIf167d98_5641,RIe20cd90_4436,RIe20a090_4404,RIe207390_4372,RIf1670f0_5632,RIf165ea8_5619,RIe202200_4314,
        RIfe83e98_7845,RIf164f30_5608,RIf1643f0_5600,RIfce8310_7664,RIf161df8_5573,RIf15ff08_5551,RIf15e018_5529,RIfe83d30_7844,RIfe84000_7846,RIf15cb00_5514,
        RIf15b5e8_5499,RIf15a508_5487,RIfc887a8_6575,RIf158d20_5470,RIf157970_5456,RIf156cc8_5447,RIfe84438_7849,RIf156020_5438,RIfc51fc8_5955,RIf154568_5419,
        RIe1f51e0_4166,RIf153050_5404,RIf1519d0_5388,RIf150788_5375,RIfe842d0_7848,RIf14f810_5364,RIf14eb68_5355,RIf14dd58_5345,RIfe84168_7847,RIe1eb2f8_4053,
        RIe1e85f8_4021,RIe1e58f8_3989,RIe1e2bf8_3957,RIe1dfef8_3925,RIe1dd1f8_3893,RIe1da4f8_3861,RIe1d77f8_3829,RIe1d1df8_3765,RIe1cf0f8_3733,RIe1cc3f8_3701,
        RIe1c96f8_3669,RIe1c69f8_3637,RIe1c3cf8_3605,RIe1c0ff8_3573,RIe1be2f8_3541,RIf14c840_5330,RIf14b5f8_5317,RIfe83a60_7842,RIfe849d8_7853,RIfc74168_6343,
        RIf149b40_5298,RIfe83bc8_7843,RIfe84708_7851,RIf148d30_5288,RIf147ae8_5275,RIfe84870_7852,RIe1b0900_3386,RIf146fa8_5267,RIf146300_5258,RIfe845a0_7850,
        RIfe83790_7840,RIe1a8638_3293,RIe1a5938_3261,RIe1a2c38_3229,RIe19ff38_3197,RIe18c438_2973,RIe178938_2749,RIe226290_4724,RIe21ae90_4596,RIe204690_4340,
        RIe1fe6f0_4272,RIe1f7aa8_4195,RIe1f05f0_4112,RIe1d4af8_3797,RIe1bb5f8_3509,RIe1ae470_3360,RIe170aa8_2659,RIdec4e38_704,RIdec2138_672,RIee1fc48_4820,
        RIdebf438_640,RIfc49490_5856,RIdebc738_608,RIdeb9a38_576,RIdeb6d38_544,RIfc48ef0_5852,RIdeb1338_480,RIfcd9b08_7499,RIdeae638_448,RIfc8b610_6608,
        RIdea9700_416,RIdea2e00_384,RIde9c500_352,RIee1c9a8_4784,RIee1b8c8_4772,RIfc80918_6485,RIfcdad50_7512,RIfe86e68_7879,RIde8cee8_277,RIfe86d00_7878,
        RIfec0d20_8314,RIde81098_219,RIfc8b8e0_6610,RIfcd2d58_7421,RIfce4530_7620,RIfc8ba48_6611,RIe16b210_2596,RIe1698c0_2578,RIe1679d0_2556,RIe164e38_2525,
        RIe162138_2493,RIee370f0_5085,RIe15f438_2461,RIfc999e0_6770,RIe15c738_2429,RIe156d38_2365,RIe154038_2333,RIfc3f260_5744,RIe151338_2301,RIfc48518_5845,
        RIe14e638_2269,RIfc99e18_6773,RIe14b938_2237,RIe148c38_2205,RIe145f38_2173,RIee34288_5052,RIee33040_5039,RIee31f60_5027,RIfcd99a0_7498,RIfe86b98_7877,
        RIdf3e9e0_2089,RIfe86a30_7876,RIdf3a4f8_2040,RIfcc3470_7244,RIee2f530_4997,RIfc7fdd8_6477,RIee2d370_4973,RIdf35200_1981,RIfec0ff0_8316,RIdf30d18_1932,
        RIfec0e88_8315,RIfcd2a88_7419,RIfc8c858_6621,RIfc47ca8_5839,RIfcd6430_7460,RIdf29f68_1854,RIdf27da8_1830,RIdf26188_1810,RIdf24568_1790,RIfc8cb28_6623,
        RIfcdb188_7515,RIdf22948_1770,RIfc475a0_5834,RIdf21430_1755,RIdf1f3d8_1732,RIfec0bb8_8313,RIfe868c8_7875,RIdf16a08_1634,RIdf13d08_1602,RIdf11008_1570,
        RIdf0e308_1538,RIdf0b608_1506,RIdf08908_1474,RIdf05c08_1442,RIdf02f08_1410,RIdefd508_1346,RIdefa808_1314,RIdef7b08_1282,RIdef4e08_1250,RIdef2108_1218,
        RIdeef408_1186,RIdeec708_1154,RIdee9a08_1122,RIee254e0_4883,RIee246d0_4873,RIee23b90_4865,RIee231b8_4858,RIfe86fd0_7880,RIdee2820_1041,RIdee0930_1019,
        RIdede608_994,RIfc55da8_5999,RIfc98a68_6759,RIfcc3038_7241,RIfc464c0_5822,RIded9310_935,RIded6e80_909,RIded4f90_887,RIded2b00_861,RIded0238_832,
        RIdecd538_800,RIdeca838_768,RIdec7b38_736,RIdeb4038_512,RIde95c00_320,RIe16dc40_2626,RIe159a38_2397,RIe143238_2141,RIdf37c30_2011,RIdf2c290_1879,
        RIdf1cb10_1703,RIdf00208_1378,RIdee6d08_1090,RIdedba70_963,RIde7bb48_193,RIe19d0d0_3164,RIe19a3d0_3132,RIf1454f0_5248,RIe1976d0_3100,RIf144578_5237,
        RIe1949d0_3068,RIe191cd0_3036,RIe18efd0_3004,RIe1895d0_2940,RIe1868d0_2908,RIf143498_5225,RIe183bd0_2876,RIfc51758_5949,RIe180ed0_2844,RIe17e1d0_2812,
        RIe17b4d0_2780,RIfc9b060_6786,RIfc9ee40_6830,RIe176e80_2730,RIe175800_2714,RIfcb70f8_7105,RIfce0cf0_7580,RIfcc4280_7254,RIfcba7d0_7144,RIee3bfb0_5141,
        RIee3aed0_5129,RIee39b20_5115,RIe173370_2688,RIf170060_5734,RIf16f3b8_5725,RIf16dea0_5710,RIf16d4c8_5703,RIf16c988_5695,RIe223428_4691,RIf16bb78_5685,
        RIe220728_4659,RIf16aa98_5673,RIe21da28_4627,RIe218028_4563,RIe215328_4531,RIf16a0c0_5666,RIe212628_4499,RIf168e78_5653,RIe20f928_4467,RIf167c30_5640,
        RIe20cc28_4435,RIe209f28_4403,RIe207228_4371,RIf166f88_5631,RIf165d40_5618,RIfec0618_8309,RIfe86760_7874,RIfc52b08_5963,RIf164288_5599,RIf163310_5588,
        RIf161c90_5572,RIf15fda0_5550,RIf15deb0_5528,RIfe865f8_7873,RIfe85d88_7867,RIf15c998_5513,RIf15b480_5498,RIf15a3a0_5486,RIf159b30_5480,RIfc83348_6515,
        RIfc4ade0_5874,RIfc89720_6586,RIe1f9f38_4221,RIfc4ac78_5873,RIfc9f110_6832,RIfc4ab10_5872,RIe1f5078_4165,RIf152ee8_5403,RIfc899f0_6588,RIf150620_5374,
        RIe1f2eb8_4141,RIf14f6a8_5363,RIf14ea00_5354,RIf14dbf0_5344,RIe1edbc0_4082,RIe1eb190_4052,RIe1e8490_4020,RIe1e5790_3988,RIe1e2a90_3956,RIe1dfd90_3924,
        RIe1dd090_3892,RIe1da390_3860,RIe1d7690_3828,RIe1d1c90_3764,RIe1cef90_3732,RIe1cc290_3700,RIe1c9590_3668,RIe1c6890_3636,RIe1c3b90_3604,RIe1c0e90_3572,
        RIe1be190_3540,RIf14c6d8_5329,RIf14b490_5316,RIfe85ef0_7868,RIfe86490_7872,RIf14a248_5303,RIfc819f8_6497,RIfec0a50_8312,RIfe861c0_7870,RIf148bc8_5287,
        RIf147980_5274,RIfe86328_7871,RIfec0780_8310,RIfcbb478_7153,RIf146198_5257,RIfe86058_7869,RIfec08e8_8311,RIe1a84d0_3292,RIe1a57d0_3260,RIe1a2ad0_3228,
        RIe19fdd0_3196,RIe18c2d0_2972,RIe1787d0_2748,RIe226128_4723,RIe21ad28_4595,RIe204528_4339,RIe1fe588_4271,RIe1f7940_4194,RIe1f0488_4111,RIe1d4990_3796,
        RIe1bb490_3508,RIe1ae308_3359,RIe170940_2658,RIdec53d8_708,RIdec26d8_676,RIee20080_4823,RIdebf9d8_644,RIee1f3d8_4814,RIdebccd8_612,RIdeb9fd8_580,
        RIdeb72d8_548,RIee1ee38_4810,RIdeb18d8_484,RIee1e898_4806,RIdeaebd8_452,RIee1da88_4796,RIdeaa420_420,RIdea3b20_388,RIde9d220_356,RIee1cde0_4787,
        RIee1bd00_4775,RIee1b490_4769,RIfcd8a28_7487,RIde91088_297,RIde8d8c0_280,RIfe7dac0_7774,RIfe7d958_7773,RIee1a518_4758,RIee19e10_4753,RIee19b40_4751,
        RIfc768c8_6371,RIfcd05f8_7393,RIfe7dd90_7776,RIee38770_5101,RIfe7dc28_7775,RIe1653d8_2529,RIe1626d8_2497,RIee373c0_5087,RIe15f9d8_2465,RIee362e0_5075,
        RIe15ccd8_2433,RIe1572d8_2369,RIe1545d8_2337,RIfe7def8_7777,RIe1518d8_2305,RIfebdeb8_8281,RIe14ebd8_2273,RIfc649e8_6167,RIe14bed8_2241,RIe1491d8_2209,
        RIe1464d8_2177,RIfe7d7f0_7772,RIfe7d688_7771,RIee32230_5029,RIfceb9e8_7703,RIfebdd50_8280,RIfe7d520_7770,RIfebdbe8_8279,RIfe7d3b8_7769,RIfc734c0_6334,
        RIee2f968_5000,RIfccfab8_7385,RIee2d7a8_4976,RIdf357a0_1985,RIdf33310_1959,RIdf312b8_1936,RIdf2f0f8_1912,RIee2bcf0_4957,RIee2a238_4938,RIee28e88_4924,
        RIee27c40_4911,RIfe7ce18_7765,RIfe7ccb0_7764,RIfe7cf80_7766,RIfe7cb48_7763,RIee27268_4904,RIee26e30_4901,RIee26890_4897,RIfcaa0d8_6957,RIee262f0_4893,
        RIfe7d250_7768,RIee26020_4891,RIfe7d0e8_7767,RIdf16fa8_1638,RIdf142a8_1606,RIdf115a8_1574,RIdf0e8a8_1542,RIdf0bba8_1510,RIdf08ea8_1478,RIdf061a8_1446,
        RIdf034a8_1414,RIdefdaa8_1350,RIdefada8_1318,RIdef80a8_1286,RIdef53a8_1254,RIdef26a8_1222,RIdeef9a8_1190,RIdeecca8_1158,RIdee9fa8_1126,RIee25648_4884,
        RIee249a0_4875,RIfebe020_8282,RIee23488_4860,RIfebe2f0_8284,RIfebe188_8283,RIfe7e1c8_7779,RIfe7e060_7778,RIfcbf7f8_7201,RIfc7aae0_6418,RIfc787b8_6393,
        RIfc618b0_6132,RIded98b0_939,RIded72b8_912,RIded5530_891,RIded2dd0_863,RIded07d8_836,RIdecdad8_804,RIdecadd8_772,RIdec80d8_740,RIdeb45d8_516,
        RIde96920_324,RIe16e1e0_2630,RIe159fd8_2401,RIe1437d8_2145,RIdf381d0_2015,RIdf2c830_1883,RIdf1d0b0_1707,RIdf007a8_1382,RIdee72a8_1094,RIdedc010_967,
        RIde7c868_197,RIe19d670_3168,RIe19a970_3136,RIfe7b630_7748,RIe197c70_3104,RIfe7b4c8_7747,RIe194f70_3072,RIe192270_3040,RIe18f570_3008,RIe189b70_2944,
        RIe186e70_2912,RIfe7b360_7746,RIe184170_2880,RIfe7b1f8_7745,RIe181470_2848,RIe17e770_2816,RIe17ba70_2784,RIf1423b8_5213,RIf140ea0_5198,RIf140360_5190,
        RIfe7b798_7749,RIf13fc58_5185,RIf13f280_5178,RIfc79460_6402,RIee3d4c8_5156,RIfe7b090_7744,RIfe7af28_7743,RIee39df0_5117,RIe1737a8_2691,RIfe7adc0_7742,
        RIfe7ac58_7741,RIf16e440_5714,RIfcb20d0_7048,RIfe7bd38_7753,RIe2239c8_4695,RIf16be48_5687,RIe220cc8_4663,RIf16aed0_5676,RIe21dfc8_4631,RIe2185c8_4567,
        RIe2158c8_4535,RIfebd7b0_8276,RIe212bc8_4503,RIfebd648_8275,RIe20fec8_4471,RIfe7b900_7750,RIe20d1c8_4439,RIe20a4c8_4407,RIe2077c8_4375,RIf167258_5633,
        RIf166178_5621,RIe2024d0_4316,RIfe7bbd0_7752,RIf165368_5611,RIf1646c0_5602,RIfcd0a30_7396,RIf1620c8_5575,RIf1601d8_5553,RIf15e2e8_5531,RIfe7ba68_7751,
        RIfe7bea0_7754,RIf15cdd0_5516,RIf15b8b8_5501,RIf15a7d8_5489,RIfca4840_6894,RIf158ff0_5472,RIf157c40_5458,RIf156f98_5449,RIfe7c170_7756,RIf156458_5441,
        RIf155918_5433,RIf1549a0_5422,RIe1f54b0_4168,RIfe7c008_7755,RIf151b38_5389,RIf150bc0_5378,RIe1f32f0_4144,RIf14fae0_5366,RIf14ee38_5357,RIf14e028_5347,
        RIe1edff8_4085,RIe1eb730_4056,RIe1e8a30_4024,RIe1e5d30_3992,RIe1e3030_3960,RIe1e0330_3928,RIe1dd630_3896,RIe1da930_3864,RIe1d7c30_3832,RIe1d2230_3768,
        RIe1cf530_3736,RIe1cc830_3704,RIe1c9b30_3672,RIe1c6e30_3640,RIe1c4130_3608,RIe1c1430_3576,RIe1be730_3544,RIf14cb10_5332,RIf14b8c8_5319,RIfebda80_8278,
        RIfe7c878_7761,RIf14a680_5306,RIfe7c2d8_7757,RIfe7c9e0_7762,RIfe7c440_7758,RIf149000_5290,RIf147db8_5277,RIe1b2688_3407,RIfebd918_8277,RIfe7c5a8_7759,
        RIf146738_5261,RIfe7c710_7760,RIe1aad98_3321,RIe1a8a70_3296,RIe1a5d70_3264,RIe1a3070_3232,RIe1a0370_3200,RIe18c870_2976,RIe178d70_2752,RIe2266c8_4727,
        RIe21b2c8_4599,RIe204ac8_4343,RIe1feb28_4275,RIe1f7ee0_4198,RIe1f0a28_4115,RIe1d4f30_3800,RIe1bba30_3512,RIe1ae8a8_3363,RIe170ee0_2662,RIdec5270_707,
        RIdec2570_675,RIee1ff18_4822,RIdebf870_643,RIfe7f848_7795,RIdebcb70_611,RIdeb9e70_579,RIdeb7170_547,RIfe7fc80_7798,RIdeb1770_483,RIfca5d58_6909,
        RIdeaea70_451,RIfcaf808_7019,RIdeaa0d8_419,RIdea37d8_387,RIde9ced8_355,RIfcdc3d0_7528,RIfcce438_7369,RIfcb0a50_7032,RIfc75680_6358,RIde90d40_296,
        RIfe7f9b0_7796,RIde89720_260,RIde85580_240,RIde81728_221,RIfc52f40_5966,RIfc82100_6502,RIfca7108_6923,RIfe7fb18_7797,RIe16b648_2599,RIe169a28_2579,
        RIe167ca0_2558,RIe165270_2528,RIe162570_2496,RIee37258_5086,RIe15f870_2464,RIee36178_5074,RIe15cb70_2432,RIe157170_2368,RIe154470_2336,RIfc86fc0_6558,
        RIe151770_2304,RIfc4eff8_5921,RIe14ea70_2272,RIfce1290_7584,RIe14bd70_2240,RIe149070_2208,RIe146370_2176,RIee34558_5054,RIee331a8_5040,RIee320c8_5028,
        RIee31150_5017,RIfe800b8_7801,RIfe7ff50_7800,RIdf3caf0_2067,RIfe7fde8_7799,RIfcc8330_7300,RIee2f800_4999,RIfca0d30_6852,RIee2d640_4975,RIdf35638_1984,
        RIdf331a8_1958,RIdf31150_1935,RIdf2ef90_1911,RIee2bb88_4956,RIee2a0d0_4937,RIee28d20_4923,RIfe7f578_7793,RIdf2a238_1856,RIdf27f10_1831,RIfe7f6e0_7794,
        RIdf246d0_1791,RIfcce9d8_7373,RIfc63638_6153,RIdf22c18_1772,RIfc62990_6144,RIdf21700_1757,RIdf1f810_1735,RIfeaa958_8257,RIdf19168_1662,RIdf16e40_1637,
        RIdf14140_1605,RIdf11440_1573,RIdf0e740_1541,RIdf0ba40_1509,RIdf08d40_1477,RIdf06040_1445,RIdf03340_1413,RIdefd940_1349,RIdefac40_1317,RIdef7f40_1285,
        RIdef5240_1253,RIdef2540_1221,RIdeef840_1189,RIdeecb40_1157,RIdee9e40_1125,RIfcb7800_7110,RIee24838_4874,RIfc4cb68_5895,RIee23320_4859,RIfe80388_7803,
        RIdee2c58_1044,RIfe80220_7802,RIdedea40_997,RIfc98900_6758,RIee223a8_4848,RIfcc8600_7302,RIee212c8_4836,RIded9748_938,RIfe804f0_7804,RIded53c8_890,
        RIded2c68_862,RIded0670_835,RIdecd970_803,RIdecac70_771,RIdec7f70_739,RIdeb4470_515,RIde965d8_323,RIe16e078_2629,RIe159e70_2400,RIe143670_2144,
        RIdf38068_2014,RIdf2c6c8_1882,RIdf1cf48_1706,RIdf00640_1381,RIdee7140_1093,RIdedbea8_966,RIde7c520_196,RIe19d508_3167,RIe19a808_3135,RIfe7ee70_7788,
        RIe197b08_3103,RIfe7efd8_7789,RIe194e08_3071,RIe192108_3039,RIe18f408_3007,RIe189a08_2943,RIe186d08_2911,RIf143768_5227,RIe184008_2879,RIfc4bbf0_5884,
        RIe181308_2847,RIe17e608_2815,RIe17b908_2783,RIfe7f410_7792,RIf140d38_5197,RIe176fe8_2731,RIe175ad0_2716,RIfe7f2a8_7791,RIf13f118_5177,RIee3e440_5167,
        RIee3d360_5155,RIee3c280_5143,RIee3b1a0_5131,RIfe7f140_7790,RIe173640_2690,RIf170330_5736,RIf16f520_5726,RIf16e2d8_5713,RIf16d630_5704,RIfe7ea38_7785,
        RIe223860_4694,RIfc9c410_6800,RIe220b60_4662,RIfcb8340_7118,RIe21de60_4630,RIe218460_4566,RIe215760_4534,RIfc9cc80_6806,RIe212a60_4502,RIfc4ddb0_5908,
        RIe20fd60_4470,RIfc873f8_6561,RIe20d060_4438,RIe20a360_4406,RIe207660_4374,RIfc86750_6552,RIfc4e4b8_5913,RIe202368_4315,RIe200a18_4297,RIf165200_5610,
        RIf164558_5601,RIf163478_5589,RIf161f60_5574,RIf160070_5552,RIf15e180_5530,RIe1fcc38_4253,RIe1fb9f0_4240,RIf15cc68_5515,RIf15b750_5500,RIf15a670_5488,
        RIf159c98_5481,RIf158e88_5471,RIf157ad8_5457,RIf156e30_5448,RIfe7e768_7783,RIf1562f0_5440,RIf1557b0_5432,RIf154838_5421,RIfe7e8d0_7784,RIf1531b8_5405,
        RIfc52400_5958,RIf150a58_5377,RIe1f3188_4143,RIf14f978_5365,RIf14ecd0_5356,RIf14dec0_5346,RIe1ede90_4084,RIe1eb5c8_4055,RIe1e88c8_4023,RIe1e5bc8_3991,
        RIe1e2ec8_3959,RIe1e01c8_3927,RIe1dd4c8_3895,RIe1da7c8_3863,RIe1d7ac8_3831,RIe1d20c8_3767,RIe1cf3c8_3735,RIe1cc6c8_3703,RIe1c99c8_3671,RIe1c6cc8_3639,
        RIe1c3fc8_3607,RIe1c12c8_3575,RIe1be5c8_3543,RIf14c9a8_5331,RIf14b760_5318,RIfe7ed08_7787,RIfe7e600_7782,RIf14a518_5305,RIfca1f78_6865,RIfe7eba0_7786,
        RIfe7e498_7781,RIf148e98_5289,RIf147c50_5276,RIfe7e330_7780,RIe1b0a68_3387,RIf147278_5269,RIf1465d0_5260,RIe1ac418_3337,RIe1aac30_3320,RIe1a8908_3295,
        RIe1a5c08_3263,RIe1a2f08_3231,RIe1a0208_3199,RIe18c708_2975,RIe178c08_2751,RIe226560_4726,RIe21b160_4598,RIe204960_4342,RIe1fe9c0_4274,RIe1f7d78_4197,
        RIe1f08c0_4114,RIe1d4dc8_3799,RIe1bb8c8_3511,RIe1ae740_3362,RIe170d78_2661,RIdec56a8_710,RIdec29a8_678,RIfc54020_5978,RIdebfca8_646,RIee1f540_4815,
        RIdebcfa8_614,RIdeba2a8_582,RIdeb75a8_550,RIfc4fe08_5931,RIdeb1ba8_486,RIfc6b630_6244,RIdeaeea8_454,RIfc6a118_6229,RIdeaaab0_422,RIdea41b0_390,
        RIde9d8b0_358,RIfc69ce0_6226,RIee1be68_4776,RIfc653c0_6174,RIee1ac20_4763,RIde91718_299,RIde8df50_282,RIde89db0_262,RIde85c10_242,RIde81db8_223,
        RIfca76a8_6927,RIfcca4f0_7324,RIfc4ce38_5897,RIfc6b360_6242,RIe16b918_2601,RIe169cf8_2581,RIe167f70_2560,RIe1656a8_2531,RIe1629a8_2499,RIee37690_5089,
        RIe15fca8_2467,RIfce93f0_7676,RIe15cfa8_2435,RIe1575a8_2371,RIe1548a8_2339,RIee35908_5068,RIe151ba8_2307,RIee34f30_5061,RIe14eea8_2275,RIfce32e8_7607,
        RIe14c1a8_2243,RIe1494a8_2211,RIe1467a8_2179,RIfcde2c0_7550,RIfc687c8_6211,RIfca9160_6946,RIfcb1590_7040,RIe141078_2117,RIdf3ef80_2093,RIdf3cdc0_2069,
        RIfebeb60_8290,RIfc64448_6163,RIee2fad0_5001,RIfca7978_6929,RIfc676e8_6199,RIdf35a70_1987,RIdf335e0_1961,RIdf31420_1937,RIdf2f3c8_1914,RIfccef78_7377,
        RIfca6fa0_6922,RIfc62558_6141,RIfc61fb8_6137,RIfe81b70_7820,RIdf281e0_1833,RIfe81cd8_7821,RIdf249a0_1793,RIfc44300_5798,RIfcafc40_7022,RIdf22ee8_1774,
        RIfcaac18_6965,RIdf219d0_1759,RIdf1fae0_1737,RIdf1b1c0_1685,RIdf19438_1664,RIdf17278_1640,RIdf14578_1608,RIdf11878_1576,RIdf0eb78_1544,RIdf0be78_1512,
        RIdf09178_1480,RIdf06478_1448,RIdf03778_1416,RIdefdd78_1352,RIdefb078_1320,RIdef8378_1288,RIdef5678_1256,RIdef2978_1224,RIdeefc78_1192,RIdeecf78_1160,
        RIdeea278_1128,RIfc611a8_6127,RIfc61a18_6133,RIfca65c8_6915,RIfca6b68_6919,RIdee4b48_1066,RIdee2dc0_1045,RIdee0c00_1021,RIdedeba8_998,RIfc626c0_6142,
        RIfc738f8_6337,RIfcb31b0_7060,RIee21430_4837,RIded9a18_940,RIded7588_914,RIded5698_892,RIded30a0_865,RIded0aa8_838,RIdecdda8_806,RIdecb0a8_774,
        RIdec83a8_742,RIdeb48a8_518,RIde96fb0_326,RIe16e4b0_2632,RIe15a2a8_2403,RIe143aa8_2147,RIdf384a0_2017,RIdf2cb00_1885,RIdf1d380_1709,RIdf00a78_1384,
        RIdee7578_1096,RIdedc2e0_969,RIde7cef8_199,RIe19d940_3170,RIe19ac40_3138,RIfc64880_6166,RIe197f40_3106,RIf144848_5239,RIe195240_3074,RIe192540_3042,
        RIe18f840_3010,RIe189e40_2946,RIe187140_2914,RIf143a38_5229,RIe184440_2882,RIfc6f140_6286,RIe181740_2850,RIe17ea40_2818,RIe17bd40_2786,RIfc64f88_6171,
        RIf141008_5199,RIe177150_2732,RIfe81738_7817,RIfccabf8_7329,RIf13f3e8_5179,RIfca81e8_6935,RIee3d630_5157,RIfc66068_6183,RIfc6ed08_6283,RIfcdde88_7547,
        RIe173a78_2693,RIfc66338_6185,RIfc6eba0_6282,RIfc664a0_6186,RIfcacdd8_6989,RIfe81468_7815,RIe223c98_4697,RIfc66d10_6192,RIe220f98_4665,RIf16b038_5677,
        RIe21e298_4633,RIe218898_4569,RIe215b98_4537,RIfc3fc38_5751,RIe212e98_4505,RIfc67850_6200,RIe210198_4473,RIf167f00_5642,RIe20d498_4441,RIe20a798_4409,
        RIe207a98_4377,RIfcacb08_6987,RIfcac9a0_6986,RIfea8900_8234,RIfe818a0_7818,RIfca8a58_6941,RIfccad60_7330,RIfcac838_6985,RIfc67418_6197,RIf160340_5554,
        RIf15e450_5532,RIfe81a08_7819,RIfe81300_7814,RIfc6dac0_6270,RIf15ba20_5502,RIfc6d958_6269,RIfc6d7f0_6268,RIfc587d8_6029,RIfc6cf80_6262,RIfc6d3b8_6265,
        RIfe815d0_7816,RIfc6d520_6266,RIfcabe60_6978,RIfc6d0e8_6263,RIe1f5780_4170,RIfc6c5a8_6255,RIfc68d68_6215,RIfc68c00_6214,RIe1f3458_4145,RIfc68a98_6213,
        RIfccb8a0_7338,RIfca9b38_6953,RIe1ee160_4086,RIe1eba00_4058,RIe1e8d00_4026,RIe1e6000_3994,RIe1e3300_3962,RIe1e0600_3930,RIe1dd900_3898,RIe1dac00_3866,
        RIe1d7f00_3834,RIe1d2500_3770,RIe1cf800_3738,RIe1ccb00_3706,RIe1c9e00_3674,RIe1c7100_3642,RIe1c4400_3610,RIe1c1700_3578,RIe1bea00_3546,RIfc6bbd0_6248,
        RIfcdd348_7539,RIe1b9438_3485,RIe1b73e0_3462,RIfcab5f0_6972,RIfccbb70_7340,RIe1b5220_3438,RIe1b3e70_3424,RIfc6c9e0_6258,RIfcab488_6971,RIfea7dc0_8226,
        RIe1b0bd0_3388,RIfc6ce18_6261,RIfcabfc8_6979,RIe1ac580_3338,RIe1aaf00_3322,RIe1a8d40_3298,RIe1a6040_3266,RIe1a3340_3234,RIe1a0640_3202,RIe18cb40_2978,
        RIe179040_2754,RIe226998_4729,RIe21b598_4601,RIe204d98_4345,RIe1fedf8_4277,RIe1f81b0_4200,RIe1f0cf8_4117,RIe1d5200_3802,RIe1bbd00_3514,RIe1aeb78_3365,
        RIe1711b0_2664,RIdec5540_709,RIdec2840_677,RIfcc4dc0_7262,RIdebfb40_645,RIfc9d7c0_6814,RIdebce40_613,RIdeba140_581,RIdeb7440_549,RIfc4d978_5905,
        RIdeb1a40_485,RIfc9dbf8_6817,RIdeaed40_453,RIfcb8610_7120,RIdeaa768_421,RIdea3e68_389,RIde9d568_357,RIfc50678_5937,RIfc507e0_5938,RIfc9dec8_6819,
        RIfc853a0_6538,RIde913d0_298,RIde8dc08_281,RIde89a68_261,RIde858c8_241,RIde81a70_222,RIfc84860_6530,RIfc50948_5939,RIfc84c98_6533,RIfcb7da0_7114,
        RIe16b7b0_2600,RIe169b90_2580,RIe167e08_2559,RIe165540_2530,RIe162840_2498,RIee37528_5088,RIe15fb40_2466,RIfcb5be0_7090,RIe15ce40_2434,RIe157440_2370,
        RIe154740_2338,RIfcd35c8_7427,RIe151a40_2306,RIfc53a80_5974,RIe14ed40_2274,RIfcc6170_7276,RIe14c040_2242,RIe149340_2210,RIe146640_2178,RIfc7f130_6468,
        RIee33310_5041,RIfcb4f38_7081,RIfc47f78_5841,RIe140f10_2116,RIdf3ee18_2092,RIdf3cc58_2068,RIdf3a7c8_2042,RIfc7fc70_6476,RIfcd27b8_7417,RIfca1000_6854,
        RIfcc6b48_7283,RIdf35908_1986,RIdf33478_1960,RIfebe9f8_8289,RIdf2f260_1913,RIfcb7968_7111,RIee2a3a0_4939,RIfc51050_5944,RIfcd3fa0_7434,RIdf2a3a0_1857,
        RIdf28078_1832,RIfe81198_7813,RIdf24838_1792,RIfc84428_6527,RIfce7ed8_7661,RIdf22d80_1773,RIfc515f0_5948,RIdf21868_1758,RIdf1f978_1736,RIdf1b058_1684,
        RIdf192d0_1663,RIdf17110_1639,RIdf14410_1607,RIdf11710_1575,RIdf0ea10_1543,RIdf0bd10_1511,RIdf09010_1479,RIdf06310_1447,RIdf03610_1415,RIdefdc10_1351,
        RIdefaf10_1319,RIdef8210_1287,RIdef5510_1255,RIdef2810_1223,RIdeefb10_1191,RIdeece10_1159,RIdeea110_1127,RIfc7e1b8_6457,RIfca19d8_6861,RIfc7dab0_6452,
        RIfc7e488_6459,RIdee49e0_1065,RIfe80d60_7810,RIfeabba0_8270,RIfe80bf8_7809,RIfcb3750_7064,RIfce9f30_7684,RIfc7e5f0_6460,RIfc56a50_6008,RIfe81030_7812,
        RIded7420_913,RIfe80ec8_7811,RIded2f38_864,RIded0940_837,RIdecdc40_805,RIdecaf40_773,RIdec8240_741,RIdeb4740_517,RIde96c68_325,RIe16e348_2631,
        RIe15a140_2402,RIe143940_2146,RIdf38338_2016,RIdf2c998_1884,RIdf1d218_1708,RIdf00910_1383,RIdee7410_1095,RIdedc178_968,RIde7cbb0_198,RIe19d7d8_3169,
        RIe19aad8_3137,RIfcc2d68_7239,RIe197dd8_3105,RIfc5c5b8_6073,RIe1950d8_3073,RIe1923d8_3041,RIe18f6d8_3009,RIe189cd8_2945,RIe186fd8_2913,RIf1438d0_5228,
        RIe1842d8_2881,RIfc5b370_6060,RIe1815d8_2849,RIe17e8d8_2817,RIe17bbd8_2785,RIfcbb748_7155,RIfc59480_6038,RIfcbbce8_7159,RIe175c38_2717,RIfcdb890_7520,
        RIfc59b88_6043,RIfc8ada0_6602,RIfcb5eb0_7092,RIfc57c98_6021,RIfc57158_6013,RIfc58aa8_6031,RIe173910_2692,RIfcc62d8_7277,RIfc8a968_6599,RIfc57428_6015,
        RIfc56d20_6010,RIfc408e0_5760,RIe223b30_4696,RIfc82970_6508,RIe220e30_4664,RIfcecc30_7716,RIe21e130_4632,RIe218730_4568,RIe215a30_4536,RIfc3fad0_5750,
        RIe212d30_4504,RIf169148_5655,RIe210030_4472,RIfc545c0_5982,RIe20d330_4440,RIe20a630_4408,RIe207930_4376,RIfc88d48_6579,RIfc4bec0_5886,RIe202638_4317,
        RIe200b80_4298,RIfc88910_6576,RIfc4c190_5888,RIfc4c2f8_5889,RIfcba398_7141,RIfcd4270_7436,RIfcba0c8_7139,RIe1fcda0_4254,RIe1fbb58_4241,RIfc53d50_5976,
        RIfc9b768_6791,RIfc537b0_5972,RIfc4c5c8_5891,RIfc9e468_6823,RIf157da8_5459,RIfcb9f60_7138,RIe1fa208_4223,RIfc849c8_6531,RIfc529a0_5962,RIfc9f6b0_6836,
        RIe1f5618_4169,RIf153320_5406,RIfcc4988_7259,RIf150d28_5379,RIfebe458_8285,RIfc87f38_6569,RIfcb7f08_7115,RIf14e190_5348,RIfe80658_7805,RIe1eb898_4057,
        RIe1e8b98_4025,RIe1e5e98_3993,RIe1e3198_3961,RIe1e0498_3929,RIe1dd798_3897,RIe1daa98_3865,RIe1d7d98_3833,RIe1d2398_3769,RIe1cf698_3737,RIe1cc998_3705,
        RIe1c9c98_3673,RIe1c6f98_3641,RIe1c4298_3609,RIe1c1598_3577,RIe1be898_3545,RIf14cc78_5333,RIf14ba30_5320,RIe1b92d0_3484,RIe1b7278_3461,RIf14a7e8_5307,
        RIf149ca8_5299,RIfebe5c0_8286,RIfe807c0_7806,RIfc50510_5936,RIfce4f08_7627,RIfe80a90_7808,RIfebe890_8288,RIfc9cde8_6807,RIfc87560_6562,RIfe80928_7807,
        RIfebe728_8287,RIe1a8bd8_3297,RIe1a5ed8_3265,RIe1a31d8_3233,RIe1a04d8_3201,RIe18c9d8_2977,RIe178ed8_2753,RIe226830_4728,RIe21b430_4600,RIe204c30_4344,
        RIe1fec90_4276,RIe1f8048_4199,RIe1f0b90_4116,RIe1d5098_3801,RIe1bbb98_3513,RIe1aea10_3364,RIe171048_2663,RIdec5978_712,RIdec2c78_680,RIfc8aad0_6600,
        RIdebff78_648,RIfc8ac38_6601,RIdebd278_616,RIdeba578_584,RIdeb7878_552,RIfc40e80_5764,RIdeb1e78_488,RIfcdaeb8_7513,RIdeaf178_456,RIee1dbf0_4797,
        RIdeab140_424,RIdea4840_392,RIde9df40_360,RIfc8b070_6604,RIfcc38a8_7247,RIfc807b0_6484,RIfcbb8b0_7156,RIde91a60_300,RIde8e298_283,RIde8a440_264,
        RIde862a0_244,RIde82100_224,RIfcbbb80_7158,RIfc8c150_6616,RIfcbbfb8_7161,RIfc54458_5981,RIe16bbe8_2603,RIfc8c2b8_6617,RIe168240_2562,RIe165978_2533,
        RIe162c78_2501,RIee37960_5091,RIe15ff78_2469,RIfcd6b38_7465,RIe15d278_2437,RIe157878_2373,RIe154b78_2341,RIfc8e5e0_6642,RIe151e78_2309,RIfcb4290_7072,
        RIe14f178_2277,RIfc56ff0_6012,RIe14c478_2245,RIe149778_2213,RIe146a78_2181,RIee346c0_5055,RIee335e0_5043,RIee32398_5030,RIee31420_5019,RIe141348_2119,
        RIe13f020_2094,RIfec16f8_8321,RIdf3a930_2043,RIfce3e28_7615,RIfc56780_6006,RIfcb4128_7071,RIfce2eb0_7604,RIdf35d40_1989,RIfe88218_7893,RIdf316f0_1939,
        RIdf2f698_1916,RIfc7f9a0_6474,RIfce4260_7618,RIfcd62c8_7459,RIfce9990_7680,RIdf2a670_1859,RIdf284b0_1835,RIdf26728_1814,RIdf24c70_1795,RIfc7ecf8_6465,
        RIfcc31a0_7242,RIfc99008_6763,RIfc46e98_5829,RIfce2a78_7601,RIdf1fdb0_1739,RIfcc6e18_7285,RIdf19708_1666,RIdf17548_1642,RIdf14848_1610,RIdf11b48_1578,
        RIdf0ee48_1546,RIdf0c148_1514,RIdf09448_1482,RIdf06748_1450,RIdf03a48_1418,RIdefe048_1354,RIdefb348_1322,RIdef8648_1290,RIdef5948_1258,RIdef2c48_1226,
        RIdeeff48_1194,RIdeed248_1162,RIdeea548_1130,RIfcd9130_7492,RIfc7cb38_6441,RIfc97af0_6748,RIfcb3e58_7069,RIdee4e18_1068,RIdee3090_1047,RIdee0ed0_1023,
        RIfe88380_7894,RIfc97dc0_6750,RIfcc2930_7236,RIfcd9298_7493,RIfc7c868_6439,RIded9ce8_942,RIded76f0_915,RIded5968_894,RIded3370_867,RIded0d78_840,
        RIdece078_808,RIdecb378_776,RIdec8678_744,RIdeb4b78_520,RIde97640_328,RIe16e780_2634,RIe15a578_2405,RIe143d78_2149,RIdf38770_2019,RIdf2cdd0_1887,
        RIdf1d650_1711,RIdf00d48_1386,RIdee7848_1098,RIdedc5b0_971,RIde7d588_201,RIe19dc10_3172,RIe19af10_3140,RIfec1590_8320,RIe198210_3108,RIfec1428_8319,
        RIe195510_3076,RIe192810_3044,RIe18fb10_3012,RIe18a110_2948,RIe187410_2916,RIfec12c0_8318,RIe184710_2884,RIfc88370_6572,RIe181a10_2852,RIe17ed10_2820,
        RIe17c010_2788,RIfc6ccb0_6260,RIfc5f858_6109,RIfca88f0_6940,RIe175f08_2719,RIfc81020_6490,RIfcc6008_7275,RIfc4ea58_5917,RIfc42140_5774,RIfca3b98_6885,
        RIfc5ac68_6055,RIfc984c8_6755,RIe173d48_2695,RIfc9b330_6788,RIf16f688_5727,RIfc42410_5776,RIfc5f588_6107,RIfe880b0_7892,RIe223f68_4699,RIf16bfb0_5688,
        RIe221268_4667,RIfc86cf0_6556,RIe21e568_4635,RIe218b68_4571,RIe215e68_4539,RIfe87de0_7890,RIe213168_4507,RIf1692b0_5656,RIe210468_4475,RIfcdf670_7564,
        RIe20d768_4443,RIe20aa68_4411,RIe207d68_4379,RIfca6460_6914,RIf1662e0_5622,RIe202908_4319,RIfe87b10_7888,RIfc58c10_6032,RIfc50ab0_5940,RIfccd790_7360,
        RIfccd1f0_7356,RIf160610_5556,RIf15e720_5534,RIfe87c78_7889,RIfe87f48_7891,RIfce7668_7655,RIfc86480_6550,RIfcd2218_7413,RIfcb01e0_7026,RIfc47b40_5838,
        RIfc84158_6525,RIfc4b920_5882,RIe1fa4d8_4225,RIfc4ba88_5883,RIfcb7530_7108,RIfcd58f0_7452,RIe1f5a50_4172,RIf153488_5407,RIf151ca0_5390,RIfc51e60_5954,
        RIe1f3728_4147,RIfc9aef8_6785,RIfcbaaa0_7146,RIfc52130_5956,RIe1ee430_4088,RIe1ebcd0_4060,RIe1e8fd0_4028,RIe1e62d0_3996,RIe1e35d0_3964,RIe1e08d0_3932,
        RIe1ddbd0_3900,RIe1daed0_3868,RIe1d81d0_3836,RIe1d27d0_3772,RIe1cfad0_3740,RIe1ccdd0_3708,RIe1ca0d0_3676,RIe1c73d0_3644,RIe1c46d0_3612,RIe1c19d0_3580,
        RIe1becd0_3548,RIfce0b88_7579,RIfc82808_6507,RIe1b9708_3487,RIe1b76b0_3464,RIfcd5bc0_7454,RIfcb69f0_7100,RIe1b54f0_3440,RIe1b4140_3426,RIfc89f90_6592,
        RIfce9af8_7681,RIe1b2958_3409,RIe1b0ea0_3390,RIfc4a138_5865,RIfc8a260_6594,RIe1ac850_3340,RIe1ab1d0_3324,RIe1a9010_3300,RIe1a6310_3268,RIe1a3610_3236,
        RIe1a0910_3204,RIe18ce10_2980,RIe179310_2756,RIe226c68_4731,RIe21b868_4603,RIe205068_4347,RIe1ff0c8_4279,RIe1f8480_4202,RIe1f0fc8_4119,RIe1d54d0_3804,
        RIe1bbfd0_3516,RIe1aee48_3367,RIe171480_2666,RIdec5810_711,RIdec2b10_679,RIfce6f60_7650,RIdebfe10_647,RIfc95228_6719,RIdebd110_615,RIdeba410_583,
        RIdeb7710_551,RIfe879a8_7887,RIdeb1d10_487,RIfcc16e8_7223,RIdeaf010_455,RIfca4f48_6899,RIdeaadf8_423,RIdea44f8_391,RIde9dbf8_359,RIee1cf48_4788,
        RIee1bfd0_4777,RIfc95660_6722,RIfcee148_7731,RIfe87840_7886,RIfe876d8_7885,RIde8a0f8_263,RIde85f58_243,RIfcb0780_7030,RIfcee9b8_7737,RIfc5f150_6104,
        RIfcdee00_7558,RIfcd8050_7480,RIe16ba80_2602,RIfca5380_6902,RIe1680d8_2561,RIe165810_2532,RIe162b10_2500,RIee377f8_5090,RIe15fe10_2468,RIee36448_5076,
        RIe15d110_2436,RIe157710_2372,RIe154a10_2340,RIfc3f3c8_5745,RIe151d10_2308,RIfcde9c8_7555,RIe14f010_2276,RIfc4a2a0_5866,RIe14c310_2244,RIe149610_2212,
        RIe146910_2180,RIfc62288_6139,RIee33478_5042,RIfc71b70_6316,RIee312b8_5018,RIe1411e0_2118,RIfe87570_7884,RIdf3cf28_2070,RIfe87408_7883,RIfcc99b0_7316,
        RIfccf0e0_7378,RIfcaeb60_7010,RIfcca220_7322,RIdf35bd8_1988,RIdf33748_1962,RIdf31588_1938,RIdf2f530_1915,RIee2be58_4958,RIee2a508_4940,RIee28ff0_4925,
        RIee27da8_4912,RIdf2a508_1858,RIdf28348_1834,RIdf265c0_1813,RIdf24b08_1794,RIfc74708_6347,RIfc42578_5777,RIfc43388_5787,RIfc745a0_6346,RIfcb0078_7025,
        RIdf1fc48_1738,RIfcaff10_7024,RIdf195a0_1665,RIdf173e0_1641,RIdf146e0_1609,RIdf119e0_1577,RIdf0ece0_1545,RIdf0bfe0_1513,RIdf092e0_1481,RIdf065e0_1449,
        RIdf038e0_1417,RIdefdee0_1353,RIdefb1e0_1321,RIdef84e0_1289,RIdef57e0_1257,RIdef2ae0_1225,RIdeefde0_1193,RIdeed0e0_1161,RIdeea3e0_1129,RIee257b0_4885,
        RIfca73d8_6925,RIee23e60_4867,RIfce66f0_7644,RIdee4cb0_1067,RIdee2f28_1046,RIdee0d68_1022,RIdeded10_999,RIfcca388_7323,RIfce6858_7645,RIfcceca8_7375,
        RIfcdc970_7532,RIded9b80_941,RIfeaaac0_8258,RIded5800_893,RIded3208_866,RIded0c10_839,RIdecdf10_807,RIdecb210_775,RIdec8510_743,RIdeb4a10_519,
        RIde972f8_327,RIe16e618_2633,RIe15a410_2404,RIe143c10_2148,RIdf38608_2018,RIdf2cc68_1886,RIdf1d4e8_1710,RIdf00be0_1385,RIdee76e0_1097,RIdedc448_970,
        RIde7d240_200,RIe19daa8_3171,RIe19ada8_3139,RIf1457c0_5250,RIe1980a8_3107,RIf1449b0_5240,RIe1953a8_3075,RIe1926a8_3043,RIe18f9a8_3011,RIe189fa8_2947,
        RIe1872a8_2915,RIf143ba0_5230,RIe1845a8_2883,RIfc912e0_6674,RIe1818a8_2851,RIe17eba8_2819,RIe17bea8_2787,RIfc915b0_6676,RIfcbe5b0_7188,RIfce3b58_7613,
        RIe175da0_2718,RIfceb448_7699,RIfcc7958_7293,RIfc42de8_5783,RIfc96e48_6739,RIfc7a810_6416,RIfc96ce0_6738,RIfcc7ac0_7294,RIe173be0_2694,RIfce39f0_7612,
        RIfc7a540_6414,RIfc91b50_6680,RIfc429b0_5780,RIfea9710_8244,RIe223e00_4698,RIfcd8488_7483,RIe221100_4666,RIfc920f0_6684,RIe21e400_4634,RIe218a00_4570,
        RIe215d00_4538,RIfc79e38_6409,RIe213000_4506,RIfcbee20_7194,RIe210300_4474,RIf168068_5643,RIe20d600_4442,RIe20a900_4410,RIe207c00_4378,RIfc5af38_6057,
        RIfcd73a8_7471,RIe2027a0_4318,RIe200ce8_4299,RIfcb2670_7052,RIfcdf940_7566,RIfc5b208_6059,RIfcbf3c0_7198,RIf1604a8_5555,RIf15e5b8_5533,RIfe872a0_7882,
        RIfe87138_7881,RIfc78920_6394,RIfec1158_8317,RIfc93338_6697,RIfcea368_7687,RIfcb23a0_7050,RIfc5bbe0_6066,RIfcede78_7729,RIe1fa370_4224,RIfcd4c48_7443,
        RIfce1dd0_7592,RIfcbf960_7202,RIe1f58e8_4171,RIfcbfc30_7204,RIfc78380_6390,RIfc93770_6700,RIe1f35c0_4146,RIfcb1f68_7047,RIfce1b00_7590,RIfc93a40_6702,
        RIe1ee2c8_4087,RIe1ebb68_4059,RIe1e8e68_4027,RIe1e6168_3995,RIe1e3468_3963,RIe1e0768_3931,RIe1dda68_3899,RIe1dad68_3867,RIe1d8068_3835,RIe1d2668_3771,
        RIe1cf968_3739,RIe1ccc68_3707,RIe1c9f68_3675,RIe1c7268_3643,RIe1c4568_3611,RIe1c1868_3579,RIe1beb68_3547,RIfcdec98_7557,RIfc94148_6707,RIe1b95a0_3486,
        RIe1b7548_3463,RIfcd12a0_7402,RIfceabd8_7693,RIe1b5388_3439,RIe1b3fd8_3425,RIfc94850_6712,RIfcd7c18_7477,RIe1b27f0_3408,RIe1b0d38_3389,RIfc76a30_6372,
        RIfce2640_7598,RIe1ac6e8_3339,RIe1ab068_3323,RIe1a8ea8_3299,RIe1a61a8_3267,RIe1a34a8_3235,RIe1a07a8_3203,RIe18cca8_2979,RIe1791a8_2755,RIe226b00_4730,
        RIe21b700_4602,RIe204f00_4346,RIe1fef60_4278,RIe1f8318_4201,RIe1f0e60_4118,RIe1d5368_3803,RIe1bbe68_3515,RIe1aece0_3366,RIe171318_2665,RIdec5c48_714,
        RIdec2f48_682,RIfc7c160_6434,RIdec0248_650,RIfcb38b8_7065,RIdebd548_618,RIdeba848_586,RIdeb7b48_554,RIfce7c08_7659,RIdeb2148_490,RIfce7aa0_7658,
        RIdeaf448_458,RIfca38c8_6883,RIdeab7d0_426,RIdea4ed0_394,RIde9e5d0_362,RIfc41e70_5772,RIfc5b0a0_6058,RIfcdbb60_7522,RIfc78650_6392,RIfea92d8_8241,
        RIde8e5e0_284,RIfea0d40_8174,RIfea0bd8_8173,RIfcdf508_7563,RIfcb1b30_7044,RIfc5ccc0_6078,RIfcb16f8_7041,RIfc77b10_6384,RIe16beb8_2605,RIe169e60_2582,
        RIe168510_2564,RIe165c48_2535,RIe162f48_2503,RIfc4f9d0_5928,RIe160248_2471,RIfc4e8f0_5916,RIe15d548_2439,RIe157b48_2375,RIe154e48_2343,RIfc4e1e8_5911,
        RIe152148_2311,RIfc868b8_6553,RIe14f448_2279,RIfc865e8_6551,RIe14c748_2247,RIe149a48_2215,RIe146d48_2183,RIfc9eb70_6828,RIfc9ecd8_6829,RIfcc5630_7268,
        RIfc83bb8_6521,RIe141618_2121,RIfea0ea8_8175,RIdf3d1f8_2072,RIdf3ac00_2045,RIee308e0_5011,RIfcd3cd0_7432,RIfc84e00_6534,RIfc834b0_6516,RIdf36010_1991,
        RIdf33a18_1964,RIdf31858_1940,RIdf2f968_1918,RIee2c128_4960,RIee2a7d8_4942,RIee292c0_4927,RIee28078_4914,RIdf2a940_1861,RIdf28780_1837,RIfea0a70_8172,
        RIfea0908_8171,RIfcd4f18_7445,RIfca0628_6847,RIdf23050_1775,RIfcd3190_7424,RIdf21b38_1760,RIdf20080_1741,RIdf1b328_1686,RIdf199d8_1668,RIdf17818_1644,
        RIdf14b18_1612,RIdf11e18_1580,RIdf0f118_1548,RIdf0c418_1516,RIdf09718_1484,RIdf06a18_1452,RIdf03d18_1420,RIdefe318_1356,RIdefb618_1324,RIdef8918_1292,
        RIdef5c18_1260,RIdef2f18_1228,RIdef0218_1196,RIdeed518_1164,RIdeea818_1132,RIfcdf3a0_7562,RIfca5218_6901,RIfcdc538_7529,RIfcdc6a0_7530,RIdee50e8_1070,
        RIdee3360_1049,RIfea07a0_8170,RIdedefe0_1001,RIfcb0d20_7034,RIfcd4978_7441,RIfca49a8_6895,RIfca1708_6859,RIded9fb8_944,RIded79c0_917,RIded5ad0_895,
        RIfeab498_8265,RIded1048_842,RIdece348_810,RIdecb648_778,RIdec8948_746,RIdeb4e48_522,RIde97cd0_330,RIe16ea50_2636,RIe15a848_2407,RIe144048_2151,
        RIdf38a40_2021,RIdf2d0a0_1889,RIdf1d920_1713,RIdf01018_1388,RIdee7b18_1100,RIdedc880_973,RIde7dc18_203,RIe19dee0_3174,RIe19b1e0_3142,RIfc67580_6198,
        RIe1984e0_3110,RIfccb030_7332,RIe1957e0_3078,RIe192ae0_3046,RIe18fde0_3014,RIe18a3e0_2950,RIe1876e0_2918,RIfc6a550_6232,RIe1849e0_2886,RIfcaa7e0_6962,
        RIe181ce0_2854,RIe17efe0_2822,RIe17c2e0_2790,RIfc65d98_6181,RIfc65690_6176,RIe1772b8_2733,RIfea0638_8169,RIfcca928_7327,RIfc607d0_6120,RIfc65258_6173,
        RIee3d798_5158,RIee3c3e8_5144,RIfca9430_6948,RIee39f58_5118,RIe174018_2697,RIfcecf00_7718,RIfc650f0_6172,RIf16e5a8_5715,RIfc43a90_5792,RIfc65528_6175,
        RIe224238_4701,RIfca9f70_6956,RIe221538_4669,RIfc6b4c8_6243,RIe21e838_4637,RIe218e38_4573,RIe216138_4541,RIfc3fda0_5752,RIe213438_4509,RIfc61310_6128,
        RIe210738_4477,RIfc60c08_6123,RIe20da38_4445,RIe20ad38_4413,RIe208038_4381,RIfc66ba8_6191,RIfccbcd8_7341,RIe202bd8_4321,RIe200fb8_4301,RIfcadbe8_6999,
        RIfccbe40_7342,RIfca7540_6926,RIfc6a3e8_6231,RIfca6898_6917,RIfc73358_6333,RIe1fd070_4256,RIe1fbe28_4243,RIfcc2660_7234,RIfc44468_5799,RIf15a940_5490,
        RIfca7270_6924,RIfc5e070_6092,RIfc5dda0_6090,RIfc7e050_6456,RIe1fa7a8_4227,RIfc5d968_6087,RIfcd9568_7495,RIfc8d668_6631,RIe1f5d20_4174,RIfca4138_6889,
        RIfc8cdf8_6625,RIfcc7c28_7295,RIe1f39f8_4149,RIfc99440_6766,RIfcbc3f0_7164,RIfc5a128_6047,RIe1ee700_4090,RIe1ebfa0_4062,RIe1e92a0_4030,RIe1e65a0_3998,
        RIe1e38a0_3966,RIe1e0ba0_3934,RIe1ddea0_3902,RIe1db1a0_3870,RIe1d84a0_3838,RIe1d2aa0_3774,RIe1cfda0_3742,RIe1cd0a0_3710,RIe1ca3a0_3678,RIe1c76a0_3646,
        RIe1c49a0_3614,RIe1c1ca0_3582,RIe1befa0_3550,RIf14cde0_5334,RIf14bb98_5321,RIe1b99d8_3489,RIe1b7980_3466,RIfc4c460_5890,RIfc9e738_6825,RIe1b5658_3441,
        RIfec54d8_8365,RIf149168_5291,RIf147f20_5278,RIe1b2ac0_3410,RIe1b1170_3392,RIf1473e0_5270,RIf1468a0_5262,RIe1acb20_3342,RIe1ab338_3325,RIe1a92e0_3302,
        RIe1a65e0_3270,RIe1a38e0_3238,RIe1a0be0_3206,RIe18d0e0_2982,RIe1795e0_2758,RIe226f38_4733,RIe21bb38_4605,RIe205338_4349,RIe1ff398_4281,RIe1f8750_4204,
        RIe1f1298_4121,RIe1d57a0_3806,RIe1bc2a0_3518,RIe1af118_3369,RIe171750_2668,RIdec5ae0_713,RIdec2de0_681,RIfc82268_6503,RIdec00e0_649,RIfcb8d18_7125,
        RIdebd3e0_617,RIdeba6e0_585,RIdeb79e0_553,RIfcb9858_7133,RIdeb1fe0_489,RIfc9efa8_6831,RIdeaf2e0_457,RIfce0750_7576,RIdeab488_425,RIdea4b88_393,
        RIde9e288_361,RIee1d0b0_4789,RIee1c138_4778,RIfcd0e68_7399,RIfc76d00_6374,RIfe89028_7903,RIfe88d58_7901,RIfe88ec0_7902,RIfe88bf0_7900,RIfcda7b0_7508,
        RIfc4d810_5904,RIfc52dd8_5965,RIfcde590_7552,RIfc4f868_5927,RIe16bd50_2604,RIfc68930_6212,RIe1683a8_2563,RIe165ae0_2534,RIe162de0_2502,RIfe88a88_7899,
        RIe1600e0_2470,RIfcc9140_7310,RIe15d3e0_2438,RIe1579e0_2374,RIe154ce0_2342,RIfc698a8_6223,RIe151fe0_2310,RIee35098_5062,RIe14f2e0_2278,RIfcc0338_7209,
        RIe14c5e0_2246,RIe1498e0_2214,RIe146be0_2182,RIfc88208_6571,RIfc85670_6540,RIfc81f98_6501,RIfcc4f28_7263,RIe1414b0_2120,RIe13f188_2095,RIdf3d090_2071,
        RIdf3aa98_2044,RIfcd2920_7418,RIfc7d7e0_6450,RIfc49760_5858,RIfce5a48_7635,RIdf35ea8_1990,RIdf338b0_1963,RIfe88920_7898,RIdf2f800_1917,RIee2bfc0_4959,
        RIee2a670_4941,RIee29158_4926,RIee27f10_4913,RIdf2a7d8_1860,RIdf28618_1836,RIdf26890_1815,RIdf24dd8_1796,RIfcad918_6997,RIfc69fb0_6228,RIfc63368_6151,
        RIfc623f0_6140,RIfc60938_6121,RIdf1ff18_1740,RIfcba500_7142,RIdf19870_1667,RIdf176b0_1643,RIdf149b0_1611,RIdf11cb0_1579,RIdf0efb0_1547,RIdf0c2b0_1515,
        RIdf095b0_1483,RIdf068b0_1451,RIdf03bb0_1419,RIdefe1b0_1355,RIdefb4b0_1323,RIdef87b0_1291,RIdef5ab0_1259,RIdef2db0_1227,RIdef00b0_1195,RIdeed3b0_1163,
        RIdeea6b0_1131,RIfcc9848_7315,RIfc69a10_6224,RIfcacc70_6988,RIfccbfa8_7343,RIdee4f80_1069,RIdee31f8_1048,RIdee1038_1024,RIdedee78_1000,RIfc84590_6528,
        RIfc9bba0_6794,RIee21b38_4842,RIfc47168_5831,RIded9e50_943,RIded7858_916,RIfe887b8_7897,RIded34d8_868,RIded0ee0_841,RIdece1e0_809,RIdecb4e0_777,
        RIdec87e0_745,RIdeb4ce0_521,RIde97988_329,RIe16e8e8_2635,RIe15a6e0_2406,RIe143ee0_2150,RIdf388d8_2020,RIdf2cf38_1888,RIdf1d7b8_1712,RIdf00eb0_1387,
        RIdee79b0_1099,RIdedc718_972,RIde7d8d0_202,RIe19dd78_3173,RIe19b078_3141,RIfca1438_6857,RIe198378_3109,RIfca35f8_6881,RIe195678_3077,RIe192978_3045,
        RIe18fc78_3013,RIe18a278_2949,RIe187578_2917,RIfcba230_7140,RIe184878_2885,RIf142d90_5220,RIe181b78_2853,RIe17ee78_2821,RIe17c178_2789,RIfc9be70_6796,
        RIfc9bd08_6795,RIfc4ccd0_5896,RIe176070_2720,RIfc87c68_6567,RIfc87b00_6566,RIfcc4c58_7261,RIfc4fca0_5930,RIfc4f598_5925,RIfc876c8_6563,RIfc4dae0_5906,
        RIe173eb0_2696,RIfcb9420_7130,RIfc4e080_5910,RIfc4e350_5912,RIfc9d388_6811,RIfc40a48_5761,RIe2240d0_4700,RIfc85508_6539,RIe2213d0_4668,RIfc9ba38_6793,
        RIe21e6d0_4636,RIe218cd0_4572,RIe215fd0_4540,RIfc52c70_5964,RIe2132d0_4508,RIfca3760_6882,RIe2105d0_4476,RIfc97988_6747,RIe20d8d0_4444,RIe20abd0_4412,
        RIe207ed0_4380,RIfceb5b0_7700,RIfcddbb8_7545,RIe202a70_4320,RIe200e50_4300,RIfc73d30_6340,RIfcaf100_7014,RIfc71468_6311,RIfcdcad8_7533,RIfcdda50_7544,
        RIfca8620_6938,RIe1fcf08_4255,RIe1fbcc0_4242,RIfc6c008_6251,RIfcdd1e0_7538,RIfca9700_6950,RIfca92c8_6947,RIfcce5a0_7370,RIfc6ba68_6247,RIfc6f410_6288,
        RIe1fa640_4226,RIfcce000_7366,RIfc53918_5973,RIfcce708_7371,RIe1f5bb8_4173,RIf1535f0_5408,RIf151e08_5391,RIfc72db8_6329,RIe1f3890_4148,RIf14fc48_5367,
        RIfc72c50_6328,RIfc73e98_6341,RIe1ee598_4089,RIe1ebe38_4061,RIe1e9138_4029,RIe1e6438_3997,RIe1e3738_3965,RIe1e0a38_3933,RIe1ddd38_3901,RIe1db038_3869,
        RIe1d8338_3837,RIe1d2938_3773,RIe1cfc38_3741,RIe1ccf38_3709,RIe1ca238_3677,RIe1c7538_3645,RIe1c4838_3613,RIe1c1b38_3581,RIe1bee38_3549,RIfcb8a48_7123,
        RIfcb84a8_7119,RIe1b9870_3488,RIe1b7818_3465,RIfc85940_6542,RIfc9e198_6821,RIfeac140_8274,RIe1b42a8_3427,RIfc518c0_5950,RIfc838e8_6519,RIfe884e8_7895,
        RIe1b1008_3391,RIfcc5900_7270,RIfc82ad8_6509,RIe1ac9b8_3341,RIfe88650_7896,RIe1a9178_3301,RIe1a6478_3269,RIe1a3778_3237,RIe1a0a78_3205,RIe18cf78_2981,
        RIe179478_2757,RIe226dd0_4732,RIe21b9d0_4604,RIe2051d0_4348,RIe1ff230_4280,RIe1f85e8_4203,RIe1f1130_4120,RIe1d5638_3805,RIe1bc138_3517,RIe1aefb0_3368,
        RIe1715e8_2667,RIdec5f18_716,RIdec3218_684,RIee20350_4825,RIdec0518_652,RIee1f6a8_4816,RIdebd818_620,RIdebab18_588,RIdeb7e18_556,RIfce4da0_7626,
        RIdeb2418_492,RIfcea908_7691,RIdeaf718_460,RIfce20a0_7594,RIdeabe60_428,RIdea5560_396,RIde9ec60_364,RIfce6420_7642,RIee1c2a0_4779,RIfc75950_6360,
        RIee1ad88_4764,RIde920f0_302,RIfea4148_8211,RIfeaa688_8255,RIfea3fe0_8210,RIde82790_226,RIfc6f848_6291,RIfc5dc38_6089,RIfc76b98_6373,RIfcae2f0_7004,
        RIe16c020_2606,RIe16a130_2584,RIe1687e0_2566,RIe165f18_2537,RIe163218_2505,RIfcadd50_7000,RIe160518_2473,RIfc55268_5991,RIe15d818_2441,RIe157e18_2377,
        RIe155118_2345,RIfc45548_5811,RIe152418_2313,RIfc498c8_5859,RIe14f718_2281,RIfcbda70_7180,RIe14ca18_2249,RIe149d18_2217,RIe147018_2185,RIee34828_5056,
        RIee33748_5044,RIee32668_5032,RIee31588_5020,RIe1418e8_2123,RIe13f458_2097,RIdf3d360_2073,RIdf3aed0_2047,RIfc526d0_5960,RIfc42848_5779,RIfcae9f8_7009,
        RIfcb7260_7106,RIfea42b0_8212,RIdf33ce8_1966,RIdf31b28_1942,RIdf2fc38_1920,RIee2c3f8_4962,RIfc4cfa0_5898,RIfc572c0_6014,RIfc4f430_5924,RIfea3e78_8209,
        RIdf28a50_1839,RIdf26b60_1817,RIdf250a8_1798,RIfc9b600_6790,RIfcb9df8_7137,RIdf23320_1777,RIfc86318_6549,RIfeabfd8_8273,RIdf201e8_1742,RIdf1b5f8_1688,
        RIdf19ca8_1670,RIdf17ae8_1646,RIdf14de8_1614,RIdf120e8_1582,RIdf0f3e8_1550,RIdf0c6e8_1518,RIdf099e8_1486,RIdf06ce8_1454,RIdf03fe8_1422,RIdefe5e8_1358,
        RIdefb8e8_1326,RIdef8be8_1294,RIdef5ee8_1262,RIdef31e8_1230,RIdef04e8_1198,RIdeed7e8_1166,RIdeeaae8_1134,RIfc89018_6581,RIfcc54c8_7267,RIfc89180_6582,
        RIfc4b380_5878,RIdee53b8_1072,RIdee34c8_1050,RIfea3d10_8208,RIdedf148_1002,RIfcae188_7003,RIfc4b0b0_5876,RIfc74870_6348,RIfce4968_7623,RIdeda288_946,
        RIded7c90_919,RIded5da0_897,RIded3640_869,RIded1318_844,RIdece618_812,RIdecb918_780,RIdec8c18_748,RIdeb5118_524,RIde98360_332,RIe16ed20_2638,
        RIe15ab18_2409,RIe144318_2153,RIdf38d10_2023,RIdf2d370_1891,RIdf1dbf0_1715,RIdf012e8_1390,RIdee7de8_1102,RIdedcb50_975,RIde7e2a8_205,RIe19e1b0_3176,
        RIe19b4b0_3144,RIfc9cf50_6808,RIe1987b0_3112,RIfc87290_6560,RIe195ab0_3080,RIe192db0_3048,RIe1900b0_3016,RIe18a6b0_2952,RIe1879b0_2920,RIfc842c0_6526,
        RIe184cb0_2888,RIfc83a50_6520,RIe181fb0_2856,RIe17f2b0_2824,RIe17c5b0_2792,RIfc9d0b8_6809,RIfc9e030_6820,RIe177420_2734,RIe176340_2722,RIfc4f700_5926,
        RIfcc4820_7258,RIfc4fb38_5929,RIfce8040_7662,RIee3c6b8_5146,RIee3b308_5132,RIfc812f0_6492,RIe174180_2698,RIfcd3028_7423,RIfc7f400_6470,RIfc46a60_5826,
        RIfc472d0_5832,RIf16cc58_5697,RIe224508_4703,RIfc7d3a8_6447,RIe221808_4671,RIfc97c58_6749,RIe21eb08_4639,RIe219108_4575,RIe216408_4543,RIfcdbe30_7524,
        RIe213708_4511,RIf169580_5658,RIe210a08_4479,RIfca4570_6892,RIe20dd08_4447,RIe20b008_4415,RIe208308_4383,RIfc7b080_6422,RIfc59cf0_6044,RIfea9b48_8247,
        RIfea4418_8213,RIfc79cd0_6408,RIfcd19a8_7407,RIfcc81c8_7299,RIf162230_5576,RIf160778_5557,RIf15e888_5535,RIfea4580_8214,RIfea46e8_8215,RIfc77f48_6387,
        RIfc41fd8_5773,RIf15aaa8_5491,RIfc7c430_6436,RIf159158_5473,RIf157f10_5460,RIfcae890_7008,RIe1faa78_4229,RIfc4a840_5870,RIfc4ed28_5919,RIfce0e58_7581,
        RIe1f5ff0_4176,RIf153758_5409,RIf151f70_5392,RIfccb468_7335,RIe1f3cc8_4151,RIfc68ed0_6216,RIfc6d250_6264,RIfca9ca0_6954,RIe1ee9d0_4092,RIe1ec270_4064,
        RIe1e9570_4032,RIe1e6870_4000,RIe1e3b70_3968,RIe1e0e70_3936,RIe1de170_3904,RIe1db470_3872,RIe1d8770_3840,RIe1d2d70_3776,RIe1d0070_3744,RIe1cd370_3712,
        RIe1ca670_3680,RIe1c7970_3648,RIe1c4c70_3616,RIe1c1f70_3584,RIe1bf270_3552,RIfc784e8_6391,RIfcbef88_7195,RIe1b9ca8_3491,RIe1b7ae8_3467,RIfcc20c0_7230,
        RIfca6190_6912,RIe1b5928_3443,RIe1b4410_3428,RIfcb81d8_7117,RIfcc5090_7264,RIe1b2d90_3412,RIe1b1440_3394,RIfcd5350_7448,RIfcb9588_7131,RIe1acc88_3343,
        RIe1ab4a0_3326,RIe1a95b0_3304,RIe1a68b0_3272,RIe1a3bb0_3240,RIe1a0eb0_3208,RIe18d3b0_2984,RIe1798b0_2760,RIe227208_4735,RIe21be08_4607,RIe205608_4351,
        RIe1ff668_4283,RIe1f8a20_4206,RIe1f1568_4123,RIe1d5a70_3808,RIe1bc570_3520,RIe1af3e8_3371,RIe171a20_2670,RIdec5db0_715,RIdec30b0_683,RIee201e8_4824,
        RIdec03b0_651,RIfcaf538_7017,RIdebd6b0_619,RIdeba9b0_587,RIdeb7cb0_555,RIfc40fe8_5765,RIdeb22b0_491,RIfcd08c8_7395,RIdeaf5b0_459,RIee1dd58_4798,
        RIdeabb18_427,RIdea5218_395,RIde9e918_363,RIee1d218_4790,RIfcedd10_7728,RIfce62b8_7641,RIfcc92a8_7311,RIde91da8_301,RIde8e928_285,RIde8a788_265,
        RIde865e8_245,RIde82448_225,RIfea1448_8179,RIfc750e0_6354,RIfcc19b8_7225,RIfced8d8_7725,RIfec5eb0_8372,RIe169fc8_2583,RIe168678_2565,RIe165db0_2536,
        RIe1630b0_2504,RIfccfc20_7386,RIe1603b0_2472,RIee365b0_5077,RIe15d6b0_2440,RIe157cb0_2376,RIe154fb0_2344,RIfea1718_8181,RIe1522b0_2312,RIee35200_5063,
        RIe14f5b0_2280,RIfcb0348_7027,RIe14c8b0_2248,RIe149bb0_2216,RIe146eb0_2184,RIfc73790_6336,RIfcdf238_7561,RIee32500_5031,RIfc94f58_6717,RIe141780_2122,
        RIe13f2f0_2096,RIfec5be0_8370,RIdf3ad68_2046,RIfea15b0_8180,RIfc5fb28_6111,RIfcae728_7007,RIfc74438_6345,RIdf36178_1992,RIdf33b80_1965,RIdf319c0_1941,
        RIdf2fad0_1919,RIee2c290_4961,RIee2a940_4943,RIfc70658_6301,RIfc704f0_6300,RIdf2aaa8_1862,RIdf288e8_1838,RIdf269f8_1816,RIdf24f40_1797,RIfc64b50_6168,
        RIfccaa90_7328,RIdf231b8_1776,RIfcad4e0_6994,RIdf21ca0_1761,RIfeaad90_8260,RIdf1b490_1687,RIdf19b40_1669,RIdf17980_1645,RIdf14c80_1613,RIdf11f80_1581,
        RIdf0f280_1549,RIdf0c580_1517,RIdf09880_1485,RIdf06b80_1453,RIdf03e80_1421,RIdefe480_1357,RIdefb780_1325,RIdef8a80_1293,RIdef5d80_1261,RIdef3080_1229,
        RIdef0380_1197,RIdeed680_1165,RIdeea980_1133,RIfc595e8_6039,RIfcac568_6983,RIfcccf20_7354,RIfccd358_7357,RIdee5250_1071,RIfea7f28_8227,RIdee11a0_1025,
        RIfea12e0_8178,RIfc679b8_6201,RIee22510_4849,RIfc6dd90_6272,RIfc6cb48_6259,RIdeda120_945,RIded7b28_918,RIded5c38_896,RIfec5d48_8371,RIded11b0_843,
        RIdece4b0_811,RIdecb7b0_779,RIdec8ab0_747,RIdeb4fb0_523,RIde98018_331,RIe16ebb8_2637,RIe15a9b0_2408,RIe1441b0_2152,RIdf38ba8_2022,RIdf2d208_1890,
        RIdf1da88_1714,RIdf01180_1389,RIdee7c80_1101,RIdedc9e8_974,RIde7df60_204,RIe19e048_3175,RIe19b348_3143,RIfcc3ce0_7250,RIe198648_3111,RIfc7efc8_6467,
        RIe195948_3079,RIe192c48_3047,RIe18ff48_3015,RIe18a548_2951,RIe187848_2919,RIfc46790_5824,RIe184b48_2887,RIfc98d38_6761,RIe181e48_2855,RIe17f148_2823,
        RIe17c448_2791,RIfcb5d48_7091,RIfc995a8_6767,RIfc9a3b8_6777,RIe1761d8_2721,RIfc54188_5979,RIfcd2bf0_7420,RIfc8b778_6609,RIfc7dee8_6455,RIee3c550_5145,
        RIfc8c420_6618,RIee3a0c0_5119,RIfeaba38_8269,RIfc46628_5823,RIfcbc288_7163,RIf16e710_5716,RIfc8fdc8_6659,RIfc48c20_5850,RIe2243a0_4702,RIfca0358_6845,
        RIe2216a0_4670,RIfc9a688_6779,RIe21e9a0_4638,RIe218fa0_4574,RIe2162a0_4542,RIfc456b0_5812,RIe2135a0_4510,RIf169418_5657,RIe2108a0_4478,RIfc8bfe8_6615,
        RIe20dba0_4446,RIe20aea0_4414,RIe2081a0_4382,RIfc8c9c0_6622,RIfc7f568_6471,RIe202d40_4322,RIe201120_4302,RIfce2910_7600,RIfc487e8_5847,RIfc46d30_5828,
        RIfc992d8_6765,RIfca2680_6870,RIfc44a08_5803,RIe1fd1d8_4257,RIe1fbf90_4244,RIfc580d0_6024,RIfcbdbd8_7181,RIfc8dd70_6636,RIfce01b0_7572,RIfc7bbc0_6430,
        RIfc90368_6663,RIfc7b8f0_6428,RIe1fa910_4228,RIfcd8b90_7488,RIfc43ec8_5795,RIfc7b788_6427,RIe1f5e88_4175,RIfc7b350_6424,RIfc90d40_6670,RIfca3490_6880,
        RIe1f3b60_4150,RIfc91010_6672,RIfcdb728_7519,RIfcd8758_7485,RIe1ee868_4091,RIe1ec108_4063,RIe1e9408_4031,RIe1e6708_3999,RIe1e3a08_3967,RIe1e0d08_3935,
        RIe1de008_3903,RIe1db308_3871,RIe1d8608_3839,RIe1d2c08_3775,RIe1cff08_3743,RIe1cd208_3711,RIe1ca508_3679,RIe1c7808_3647,RIe1c4b08_3615,RIe1c1e08_3583,
        RIe1bf108_3551,RIf14cf48_5335,RIfc78d58_6397,RIe1b9b40_3490,RIfec5910_8368,RIfc78a88_6395,RIfcd51e8_7447,RIe1b57c0_3442,RIfea1010_8176,RIf1492d0_5292,
        RIfec5a78_8369,RIe1b2c28_3411,RIe1b12d8_3393,RIfec5640_8366,RIf146a08_5263,RIfec57a8_8367,RIfea1178_8177,RIe1a9448_3303,RIe1a6748_3271,RIe1a3a48_3239,
        RIe1a0d48_3207,RIe18d248_2983,RIe179748_2759,RIe2270a0_4734,RIe21bca0_4606,RIe2054a0_4350,RIe1ff500_4282,RIe1f88b8_4205,RIe1f1400_4122,RIe1d5908_3807,
        RIe1bc408_3519,RIe1af280_3370,RIe1718b8_2669,RIdec6350_719,RIdec3650_687,RIfcaf3d0_7016,RIdec0950_655,RIfc6a280_6230,RIdebdc50_623,RIdebaf50_591,
        RIdeb8250_559,RIfc42f50_5784,RIdeb2850_495,RIfc981f8_6753,RIdeafb50_463,RIfc8c6f0_6620,RIdeac838_431,RIdea5f38_399,RIde9f638_367,RIee1d4e8_4792,
        RIfcda648_7507,RIfcc6440_7278,RIfcd5620_7450,RIde92ac8_305,RIfea34a0_8202,RIfea31d0_8200,RIfea3338_8201,RIfcb6b58_7101,RIfcb6888_7099,RIfc9dd60_6818,
        RIee19708_4748,RIfc50c18_5941,RIe16c458_2609,RIfc80a80_6486,RIfec62e8_8375,RIe166350_2540,RIe163650_2508,RIee37d98_5094,RIe160950_2476,RIfcaa678_6961,
        RIe15dc50_2444,RIe158250_2380,RIe155550_2348,RIfea3ba8_8207,RIe152850_2316,RIee35638_5066,RIe14fb50_2284,RIfc62f30_6148,RIe14ce50_2252,RIe14a150_2220,
        RIe147450_2188,RIfc97f28_6751,RIfc89888_6587,RIfc8f558_6653,RIfc52838_5961,RIe141bb8_2125,RIe13f890_2100,RIdf3d798_2076,RIdf3b308_2050,RIee30a48_5012,
        RIfc568e8_6007,RIee2e9f0_4989,RIee2dbe0_4979,RIdf365b0_1995,RIfea38d8_8205,RIfea3a40_8206,RIdf2ff08_1922,RIee2c6c8_4964,RIee2ac10_4945,RIee29590_4929,
        RIee28348_4916,RIdf2ad78_1864,RIdf28e88_1842,RIfea3608_8203,RIfea3770_8204,RIfcc0d10_7216,RIfc75c20_6362,RIfca50b0_6900,RIfc74e10_6352,RIfcc9410_7312,
        RIdf20620_1745,RIfc73628_6335,RIdf1a0e0_1673,RIdf17f20_1649,RIdf15220_1617,RIdf12520_1585,RIdf0f820_1553,RIdf0cb20_1521,RIdf09e20_1489,RIdf07120_1457,
        RIdf04420_1425,RIdefea20_1361,RIdefbd20_1329,RIdef9020_1297,RIdef6320_1265,RIdef3620_1233,RIdef0920_1201,RIdeedc20_1169,RIdeeaf20_1137,RIfcab8c0_6974,
        RIfc7c598_6437,RIfc5beb0_6068,RIfc58ee0_6034,RIdee5688_1074,RIdee3798_1052,RIdee15d8_1028,RIdedf580_1005,RIfcb3048_7059,RIfc72ae8_6327,RIfca3d00_6886,
        RIfcb6450_7096,RIdeda558_948,RIded7f60_921,RIfea3068_8199,RIded3a78_872,RIded1750_847,RIdecea50_815,RIdecbd50_783,RIdec9050_751,RIdeb5550_527,
        RIde98d38_335,RIe16f158_2641,RIe15af50_2412,RIe144750_2156,RIdf39148_2026,RIdf2d7a8_1894,RIdf1e028_1718,RIdf01720_1393,RIdee8220_1105,RIdedcf88_978,
        RIde7ec80_208,RIe19e5e8_3179,RIe19b8e8_3147,RIfca84b8_6937,RIe198be8_3115,RIfc846f8_6529,RIe195ee8_3083,RIe1931e8_3051,RIe1904e8_3019,RIe18aae8_2955,
        RIe187de8_2923,RIfce2be0_7602,RIe1850e8_2891,RIfc8e310_6640,RIe1823e8_2859,RIe17f6e8_2827,RIe17c9e8_2795,RIfcd1570_7404,RIfccc278_7345,RIf1404c8_5191,
        RIfea2d98_8197,RIfcc1b20_7226,RIfc60398_6117,RIee3e5a8_5168,RIee3da68_5160,RIfc642e0_6162,RIfca7f18_6933,RIee3a228_5120,RIfec6180_8374,RIfca9598_6949,
        RIfc5c720_6074,RIfc6bea0_6250,RIfccaec8_7331,RIfc44cd8_5805,RIe224940_4706,RIfcb6180_7094,RIe221c40_4674,RIfc55ad8_5997,RIe21ef40_4642,RIe219540_4578,
        RIe216840_4546,RIfc4dc48_5907,RIe213b40_4514,RIfcdcf10_7536,RIe210e40_4482,RIfcab1b8_6969,RIe20e140_4450,RIe20b440_4418,RIe208740_4386,RIfce3720_7610,
        RIfc64178_6161,RIe203178_4325,RIe201558_4305,RIfcd2ec0_7422,RIf164828_5603,RIfc7f838_6473,RIf162398_5577,RIfcc9c80_7318,RIfca8bc0_6942,RIfea2ac8_8195,
        RIfea2c30_8196,RIfc59318_6037,RIfc4f160_5922,RIf15ac10_5492,RIfcebf88_7707,RIfcbb040_7150,RIfca1870_6860,RIfc93d10_6704,RIe1faeb0_4232,RIf1565c0_5442,
        RIf155a80_5434,RIfc45c50_5816,RIe1f6428_4179,RIfccdbc8_7363,RIfcccae8_7351,RIfca6cd0_6920,RIfec6018_8373,RIfc64010_6160,RIfc434f0_5788,RIfc4c028_5887,
        RIe1eee08_4095,RIe1ec6a8_4067,RIe1e99a8_4035,RIe1e6ca8_4003,RIe1e3fa8_3971,RIe1e12a8_3939,RIe1de5a8_3907,RIe1db8a8_3875,RIe1d8ba8_3843,RIe1d31a8_3779,
        RIe1d04a8_3747,RIe1cd7a8_3715,RIe1caaa8_3683,RIe1c7da8_3651,RIe1c50a8_3619,RIe1c23a8_3587,RIe1bf6a8_3555,RIfc63908_6155,RIfc6bd38_6249,RIe1ba0e0_3494,
        RIe1b7f20_3470,RIfc66fe0_6194,RIfc92ac8_6691,RIe1b5d60_3446,RIfea2f00_8198,RIfc9bfd8_6797,RIfc50d80_5942,RIe1b31c8_3415,RIe1b1878_3397,RIfc4df18_5909,
        RIfc9d658_6813,RIe1ad0c0_3346,RIe1ab8d8_3329,RIe1a99e8_3307,RIe1a6ce8_3275,RIe1a3fe8_3243,RIe1a12e8_3211,RIe18d7e8_2987,RIe179ce8_2763,RIe227640_4738,
        RIe21c240_4610,RIe205a40_4354,RIe1ffaa0_4286,RIe1f8e58_4209,RIe1f19a0_4126,RIe1d5ea8_3811,RIe1bc9a8_3523,RIe1af820_3374,RIe171e58_2673,RIdec61e8_718,
        RIdec34e8_686,RIee20620_4827,RIdec07e8_654,RIfc4b7b8_5881,RIdebdae8_622,RIdebade8_590,RIdeb80e8_558,RIfc41150_5766,RIdeb26e8_494,RIfc87830_6564,
        RIdeaf9e8_462,RIee1dec0_4799,RIdeac4f0_430,RIdea5bf0_398,RIde9f2f0_366,RIee1d380_4791,RIfc77c78_6385,RIfc84f68_6535,RIfc6ff50_6296,RIde92780_304,
        RIde8efb8_287,RIde8ae18_267,RIde86c78_247,RIee1a680_4759,RIee19f78_4754,RIfcd7240_7470,RIfcbeb50_7192,RIfc76328_6367,RIe16c2f0_2608,RIee388d8_5102,
        RIfea20f0_8188,RIe1661e8_2539,RIe1634e8_2507,RIee37c30_5093,RIe1607e8_2475,RIfce7500_7654,RIe15dae8_2443,RIe1580e8_2379,RIe1553e8_2347,RIfc3f698_5747,
        RIe1526e8_2315,RIee354d0_5065,RIe14f9e8_2283,RIfc83e88_6523,RIe14cce8_2251,RIe149fe8_2219,RIe1472e8_2187,RIfcea4d0_7688,RIfcb7ad0_7112,RIfc695d8_6221,
        RIfc51a28_5951,RIe141a50_2124,RIe13f728_2099,RIdf3d630_2075,RIdf3b1a0_2049,RIfca9e08_6955,RIee2fda0_5003,RIfc88a78_6577,RIee2da78_4978,RIdf36448_1994,
        RIdf33fb8_1968,RIdf31df8_1944,RIfea2258_8189,RIee2c560_4963,RIee2aaa8_4944,RIee29428_4928,RIee281e0_4915,RIdf2ac10_1863,RIdf28d20_1841,RIfea27f8_8193,
        RIfea2960_8194,RIfcdabe8_7511,RIfca08f8_6849,RIfc8b1d8_6605,RIfc49058_5853,RIfca0a60_6850,RIdf204b8_1744,RIfc99cb0_6772,RIdf19f78_1672,RIdf17db8_1648,
        RIdf150b8_1616,RIdf123b8_1584,RIdf0f6b8_1552,RIdf0c9b8_1520,RIdf09cb8_1488,RIdf06fb8_1456,RIdf042b8_1424,RIdefe8b8_1360,RIdefbbb8_1328,RIdef8eb8_1296,
        RIdef61b8_1264,RIdef34b8_1232,RIdef07b8_1200,RIdeedab8_1168,RIdeeadb8_1136,RIfcd1f48_7411,RIfc57f68_6023,RIfcbe2e0_7186,RIfcd8fc8_7491,RIdee5520_1073,
        RIfea2690_8192,RIdee1470_1027,RIdedf418_1004,RIfc57b30_6020,RIfcb35e8_7063,RIfcbd7a0_7178,RIfc91178_6673,RIfea2528_8191,RIded7df8_920,RIfea23c0_8190,
        RIded3910_871,RIded15e8_846,RIdece8e8_814,RIdecbbe8_782,RIdec8ee8_750,RIdeb53e8_526,RIde989f0_334,RIe16eff0_2640,RIe15ade8_2411,RIe1445e8_2155,
        RIdf38fe0_2025,RIdf2d640_1893,RIdf1dec0_1717,RIdf015b8_1392,RIdee80b8_1104,RIdedce20_977,RIde7e938_207,RIe19e480_3178,RIe19b780_3146,RIfccc980_7350,
        RIe198a80_3114,RIfcc1148_7219,RIe195d80_3082,RIe193080_3050,RIe190380_3018,RIe18a980_2954,RIe187c80_2922,RIfcb2ee0_7058,RIe184f80_2890,RIfc615e0_6130,
        RIe182280_2858,RIe17f580_2826,RIe17c880_2794,RIfc69038_6217,RIfc4c898_5893,RIfc6f2a8_6287,RIe1764a8_2723,RIfcad0a8_6991,RIfc6adc0_6238,RIfc70388_6299,
        RIfea1b50_8184,RIfea1f88_8187,RIfc56e88_6011,RIfea1cb8_8185,RIe174450_2700,RIfc60d70_6124,RIfc6a820_6234,RIfea1e20_8186,RIf16d798_5705,RIfc40bb0_5762,
        RIe2247d8_4705,RIfc77138_6377,RIe221ad8_4673,RIfcd7d80_7478,RIe21edd8_4641,RIe2193d8_4577,RIe2166d8_4545,RIfc40070_5754,RIe2139d8_4513,RIf169850_5660,
        RIe210cd8_4481,RIfcc1580_7222,RIe20dfd8_4449,RIe20b2d8_4417,RIe2085d8_4385,RIfcd0058_7389,RIfc749d8_6349,RIe203010_4324,RIe2013f0_4304,RIfc60230_6116,
        RIfc60668_6119,RIfcaf970_7020,RIfc45818_5813,RIf160a48_5559,RIf15eb58_5537,RIfea1880_8182,RIfea19e8_8183,RIfc72110_6320,RIfc49b98_5861,RIfcca0b8_7321,
        RIfc71738_6313,RIfc4ca00_5894,RIfc71030_6308,RIfcde428_7551,RIe1fad48_4231,RIfc70bf8_6305,RIfc63a70_6156,RIfca7db0_6932,RIe1f62c0_4178,RIfcada80_6998,
        RIfc6fde8_6295,RIfc6f578_6289,RIe1f3f98_4153,RIfcde158_7549,RIfcad378_6993,RIfc65f00_6182,RIe1eeca0_4094,RIe1ec540_4066,RIe1e9840_4034,RIe1e6b40_4002,
        RIe1e3e40_3970,RIe1e1140_3938,RIe1de440_3906,RIe1db740_3874,RIe1d8a40_3842,RIe1d3040_3778,RIe1d0340_3746,RIe1cd640_3714,RIe1ca940_3682,RIe1c7c40_3650,
        RIe1c4f40_3618,RIe1c2240_3586,RIe1bf540_3554,RIfc69308_6219,RIfccba08_7339,RIe1b9f78_3493,RIe1b7db8_3469,RIfccd628_7359,RIfc69740_6222,RIe1b5bf8_3445,
        RIe1b4578_3429,RIfccf950_7384,RIf148088_5279,RIe1b3060_3414,RIe1b1710_3396,RIfc9f818_6837,RIfcb9c90_7136,RIe1acf58_3345,RIe1ab770_3328,RIe1a9880_3306,
        RIe1a6b80_3274,RIe1a3e80_3242,RIe1a1180_3210,RIe18d680_2986,RIe179b80_2762,RIe2274d8_4737,RIe21c0d8_4609,RIe2058d8_4353,RIe1ff938_4285,RIe1f8cf0_4208,
        RIe1f1838_4125,RIe1d5d40_3810,RIe1bc840_3522,RIe1af6b8_3373,RIe171cf0_2672;
output R_58_102f1b78,R_59_be1fc68,R_5a_10279198,R_5b_102299e8,R_5c_101d0448,R_5d_f7f82f0,R_5e_be21600,R_5f_f7fa5b8,R_60_1027d530,
        R_61_10205ae8,R_62_10283510,R_63_f82b578,R_64_ace4e68,R_65_f8204e0,R_66_1027a0b0,R_67_1022dc30,R_68_102478a8,R_69_10286f78,R_6a_f7edd80,
        R_6b_101c3628,R_6c_f7fbe00,R_6d_f7ce9f8,R_6e_f7c8830,R_6f_101ffc68,R_70_f7d4000,R_71_acee958,R_72_94046c0,R_73_101ee420,R_74_102eb268,
        R_75_b320c50,R_76_ad80a90,R_77_1027fd48,R_78_f7ce4b8,R_79_ad77048,R_7a_102a6ae0,R_7b_f7e4c78,R_7c_e2a6ce0,R_7d_101e86e0,R_7e_e2a9cc8,
        R_7f_10292be0,R_80_b33cde8,R_81_101e2908,R_82_102e9780,R_83_f8157a0,R_84_f819358,R_85_ace8b70,R_86_be142b0,R_87_f81b770,R_88_b330278,
        R_89_f7fe9f8,R_8a_101cf488,R_8b_f8225c0,R_8c_101d4738,R_8d_101c4000,R_8e_101fe960,R_8f_102a0330,R_90_f7f4bd0,R_91_1023e5a8,R_92_10248da8,
        R_93_be2c938,R_94_f7f5458,R_95_f7c6808,R_96_be316a8,R_97_e2a0328,R_98_be2d850,R_99_10217db0,R_9a_f7ec340,R_9b_be23ec0,R_9c_101d4540,
        R_9d_f800828,R_9e_102970c8,R_9f_10221de0,R_a0_ad8d568,R_a1_be4eb58,R_a2_f7c5500,R_a3_ad88f30,R_a4_f82f088,R_a5_f7dcbc8,R_a6_10292940,
        R_a7_be138d8,R_a8_acee418,R_a9_ad84450,R_aa_be10838,R_ab_be31fd8,R_ac_acdaef0,R_ad_acea908,R_ae_101f8830,R_af_f7dec98,R_b0_101e2c50,
        R_b1_f801b30,R_b2_be16e00,R_b3_102e3cf0,R_b4_10291788;

wire \8308 , \8309_ZERO , \8310_ONE , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 ,
         \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 ,
         \8327 , \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 ,
         \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345 , \8346 ,
         \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 ,
         \8357 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 , \8366 ,
         \8367 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 ,
         \8377 , \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 ,
         \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 ,
         \8397 , \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 ,
         \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 ,
         \8417 , \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 ,
         \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 ,
         \8437 , \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 ,
         \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 , \8455 , \8456 ,
         \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 , \8465 , \8466 ,
         \8467 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 , \8475 , \8476 ,
         \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 ,
         \8487 , \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 ,
         \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 ,
         \8507 , \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 , \8515 , \8516 ,
         \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 ,
         \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 ,
         \8537 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 ,
         \8547 , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556 ,
         \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 , \8565 , \8566 ,
         \8567 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 ,
         \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 ,
         \8587 , \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 ,
         \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 ,
         \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 ,
         \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 ,
         \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 ,
         \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 ,
         \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 ,
         \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 ,
         \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 ,
         \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 ,
         \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 ,
         \8697 , \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 , \8705 , \8706 ,
         \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 ,
         \8717 , \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 ,
         \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 ,
         \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 ,
         \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 ,
         \8757 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 , \8765 , \8766 ,
         \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 ,
         \8777 , \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 , \8786 ,
         \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 ,
         \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 ,
         \8807 , \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 ,
         \8817 , \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 ,
         \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 ,
         \8837 , \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 , \8845 , \8846 ,
         \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 ,
         \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 , \8865 , \8866 ,
         \8867 , \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 ,
         \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 ,
         \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 , \8895 , \8896 ,
         \8897 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 ,
         \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 ,
         \8917 , \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 , \8925 , \8926 ,
         \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 ,
         \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 , \8945 , \8946 ,
         \8947 , \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 , \8955 , \8956 ,
         \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966 ,
         \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 ,
         \8977 , \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 , \8985 , \8986 ,
         \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 ,
         \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 ,
         \9007 , \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 ,
         \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 ,
         \9027 , \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 , \9035 , \9036 ,
         \9037 , \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046 ,
         \9047 , \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 , \9055 , \9056 ,
         \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 , \9065 , \9066 ,
         \9067 , \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 , \9075 , \9076 ,
         \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 , \9085 , \9086 ,
         \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 ,
         \9097 , \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 , \9105 , \9106 ,
         \9107 , \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 , \9115 , \9116 ,
         \9117 , \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 , \9125 , \9126 ,
         \9127 , \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 , \9135 , \9136 ,
         \9137 , \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 , \9145 , \9146 ,
         \9147 , \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 , \9155 , \9156 ,
         \9157 , \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 , \9165 , \9166 ,
         \9167 , \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 , \9175 , \9176 ,
         \9177 , \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 , \9185 , \9186 ,
         \9187 , \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 , \9195 , \9196 ,
         \9197 , \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 , \9205 , \9206 ,
         \9207 , \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 , \9215 , \9216 ,
         \9217 , \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 , \9225 , \9226 ,
         \9227 , \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 , \9235 , \9236 ,
         \9237 , \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 , \9245 , \9246 ,
         \9247 , \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 , \9255 , \9256 ,
         \9257 , \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 , \9265 , \9266 ,
         \9267 , \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 , \9275 , \9276 ,
         \9277 , \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 , \9285 , \9286 ,
         \9287 , \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 , \9295 , \9296 ,
         \9297 , \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 , \9305 , \9306 ,
         \9307 , \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 , \9315 , \9316 ,
         \9317 , \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 , \9325 , \9326 ,
         \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 , \9335 , \9336 ,
         \9337 , \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 , \9345 , \9346 ,
         \9347 , \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 , \9355 , \9356 ,
         \9357 , \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 , \9365 , \9366 ,
         \9367 , \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 , \9375 , \9376 ,
         \9377 , \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 , \9385 , \9386 ,
         \9387 , \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 , \9395 , \9396 ,
         \9397 , \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 , \9405 , \9406 ,
         \9407 , \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 , \9415 , \9416 ,
         \9417 , \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 , \9425 , \9426 ,
         \9427 , \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 , \9435 , \9436 ,
         \9437 , \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 , \9445 , \9446 ,
         \9447 , \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 , \9455 , \9456 ,
         \9457 , \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 , \9465 , \9466 ,
         \9467 , \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 , \9475 , \9476 ,
         \9477 , \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 , \9485 , \9486 ,
         \9487 , \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 , \9495 , \9496 ,
         \9497 , \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 , \9505 , \9506 ,
         \9507 , \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 , \9515 , \9516 ,
         \9517 , \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 , \9525 , \9526 ,
         \9527 , \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 , \9535 , \9536 ,
         \9537 , \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 , \9545 , \9546 ,
         \9547 , \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 , \9555 , \9556 ,
         \9557 , \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 , \9565 , \9566 ,
         \9567 , \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 , \9575 , \9576 ,
         \9577 , \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 , \9585 , \9586 ,
         \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 , \9595 , \9596 ,
         \9597 , \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 ,
         \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 , \9615 , \9616 ,
         \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 ,
         \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 ,
         \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 , \9645 , \9646 ,
         \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 ,
         \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 , \9665 , \9666 ,
         \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 , \9675 , \9676 ,
         \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 ,
         \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 ,
         \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 ,
         \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 ,
         \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 ,
         \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 ,
         \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 ,
         \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 ,
         \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 ,
         \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 ,
         \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 ,
         \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 ,
         \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 ,
         \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 ,
         \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 ,
         \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 ,
         \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 ,
         \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 ,
         \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 ,
         \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 ,
         \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 ,
         \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 ,
         \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 ,
         \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 ,
         \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 ,
         \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 ,
         \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 ,
         \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 ,
         \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 ,
         \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 ,
         \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 ,
         \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 ,
         \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 ,
         \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 ,
         \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 ,
         \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 ,
         \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 ,
         \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 ,
         \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 , \10065 , \10066 ,
         \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 ,
         \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 ,
         \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 ,
         \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 ,
         \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 ,
         \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 ,
         \10127 , \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 ,
         \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 ,
         \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 ,
         \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 ,
         \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 ,
         \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 ,
         \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 ,
         \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 ,
         \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 ,
         \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 ,
         \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 ,
         \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 ,
         \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 ,
         \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 , \10265 , \10266 ,
         \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 ,
         \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 ,
         \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 ,
         \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 ,
         \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 ,
         \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 ,
         \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 ,
         \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 ,
         \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 ,
         \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 ,
         \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 ,
         \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 ,
         \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 ,
         \10397 , \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 ,
         \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 ,
         \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 , \10425 , \10426 ,
         \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 ,
         \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 ,
         \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 ,
         \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 ,
         \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 ,
         \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 ,
         \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 ,
         \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506 ,
         \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 ,
         \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 ,
         \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 ,
         \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 ,
         \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 ,
         \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 ,
         \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 ,
         \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 ,
         \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 ,
         \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 ,
         \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 ,
         \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 ,
         \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 ,
         \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 ,
         \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 , \10656 ,
         \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 ,
         \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 ,
         \10677 , \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 , \10685 , \10686 ,
         \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 ,
         \10697 , \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 , \10705 , \10706 ,
         \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 ,
         \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 ,
         \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 ,
         \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 ,
         \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 ,
         \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 ,
         \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 ,
         \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 ,
         \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 ,
         \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 ,
         \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 ,
         \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 ,
         \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 ,
         \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 ,
         \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 ,
         \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 ,
         \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 ,
         \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 ,
         \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 ,
         \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 ,
         \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 ,
         \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 ,
         \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 ,
         \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 ,
         \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 ,
         \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 ,
         \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 ,
         \10977 , \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 , \10985 , \10986 ,
         \10987 , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 ,
         \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 ,
         \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 ,
         \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 ,
         \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 ,
         \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 ,
         \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 ,
         \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 ,
         \11067 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 ,
         \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 ,
         \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 ,
         \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 ,
         \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 ,
         \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 ,
         \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136 ,
         \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 ,
         \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 ,
         \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 ,
         \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 ,
         \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 ,
         \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 ,
         \11197 , \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 , \11205 , \11206 ,
         \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 ,
         \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 ,
         \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 ,
         \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 ,
         \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 ,
         \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 ,
         \11267 , \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 , \11275 , \11276 ,
         \11277 , \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 , \11285 , \11286 ,
         \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 ,
         \11297 , \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 , \11305 , \11306 ,
         \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 ,
         \11317 , \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 ,
         \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 ,
         \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 ,
         \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 ,
         \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 ,
         \11367 , \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 ,
         \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 ,
         \11387 , \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 ,
         \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 ,
         \11407 , \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 ,
         \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 ,
         \11427 , \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 , \11435 , \11436 ,
         \11437 , \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 ,
         \11447 , \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 ,
         \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 ,
         \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 ,
         \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486 ,
         \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 ,
         \11497 , \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 , \11505 , \11506 ,
         \11507 , \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515 , \11516 ,
         \11517 , \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 ,
         \11527 , \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 ,
         \11537 , \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 , \11545 , \11546 ,
         \11547 , \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 ,
         \11557 , \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 , \11565 , \11566 ,
         \11567 , \11568 , \11569 , \11570 , \11571 , \11572 , \11573 , \11574 , \11575 , \11576 ,
         \11577 , \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 , \11585 , \11586 ,
         \11587 , \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 , \11595 , \11596 ,
         \11597 , \11598 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 , \11605 , \11606 ,
         \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 ,
         \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 ,
         \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 , \11635 , \11636 ,
         \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 ,
         \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 ,
         \11657 , \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 ,
         \11667 , \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 ,
         \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 ,
         \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 ,
         \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 ,
         \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 ,
         \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 ,
         \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 , \11735 , \11736 ,
         \11737 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 ,
         \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 ,
         \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 ,
         \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 ,
         \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 , \11786 ,
         \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 ,
         \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 ,
         \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 ,
         \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 ,
         \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 ,
         \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 ,
         \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 ,
         \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 ,
         \11867 , \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 , \11875 , \11876 ,
         \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 ,
         \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 ,
         \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 ,
         \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 ,
         \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 ,
         \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 ,
         \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 ,
         \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 ,
         \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 ,
         \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 , \11975 , \11976 ,
         \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 ,
         \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 ,
         \11997 , \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 , \12005 , \12006 ,
         \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 ,
         \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 ,
         \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 ,
         \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 ,
         \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 ,
         \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 ,
         \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 ,
         \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 ,
         \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 ,
         \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 ,
         \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 ,
         \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 ,
         \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 ,
         \12137 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 , \12145 , \12146 ,
         \12147 , \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 , \12155 , \12156 ,
         \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 ,
         \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 ,
         \12177 , \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 , \12185 , \12186 ,
         \12187 , \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 ,
         \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 ,
         \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 ,
         \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 ,
         \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 ,
         \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 ,
         \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 ,
         \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 ,
         \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 ,
         \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 ,
         \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 ,
         \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 ,
         \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 , \12315 , \12316 ,
         \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 ,
         \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 ,
         \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 ,
         \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 ,
         \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 ,
         \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 ,
         \12377 , \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 ,
         \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 ,
         \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 ,
         \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 ,
         \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 ,
         \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 ,
         \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446 ,
         \12447 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 ,
         \12457 , \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 ,
         \12467 , \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 ,
         \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 , \12486 ,
         \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 ,
         \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 ,
         \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 ,
         \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 ,
         \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 ,
         \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 ,
         \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 ,
         \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 ,
         \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 ,
         \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 ,
         \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 ,
         \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 ,
         \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 ,
         \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 ,
         \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635 , \12636 ,
         \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 ,
         \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 ,
         \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 ,
         \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 ,
         \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 ,
         \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 ,
         \12697 , \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 ,
         \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 ,
         \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 ,
         \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 ,
         \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 ,
         \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 ,
         \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 ,
         \12767 , \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 , \12775 , \12776 ,
         \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 ,
         \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 ,
         \12797 , \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 , \12805 , \12806 ,
         \12807 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 ,
         \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 ,
         \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 ,
         \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 ,
         \12847 , \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 ,
         \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 ,
         \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 ,
         \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 , \12885 , \12886 ,
         \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 ,
         \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 ,
         \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 ,
         \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 ,
         \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 ,
         \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 ,
         \12947 , \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 , \12955 , \12956 ,
         \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 ,
         \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 ,
         \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 ,
         \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 ,
         \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 ,
         \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 ,
         \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 ,
         \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 ,
         \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 ,
         \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 ,
         \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 ,
         \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 ,
         \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 ,
         \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 ,
         \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 ,
         \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 ,
         \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 ,
         \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 ,
         \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 ,
         \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 ,
         \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 ,
         \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 ,
         \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 ,
         \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 ,
         \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 ,
         \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 ,
         \13217 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 ,
         \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 ,
         \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 ,
         \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 ,
         \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 ,
         \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 ,
         \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 ,
         \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 , \13295 , \13296 ,
         \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 ,
         \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 ,
         \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 , \13326 ,
         \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 ,
         \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 ,
         \13347 , \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 ,
         \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 , \13365 , \13366 ,
         \13367 , \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 , \13375 , \13376 ,
         \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 ,
         \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 ,
         \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 , \13405 , \13406 ,
         \13407 , \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 , \13415 , \13416 ,
         \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 ,
         \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 ,
         \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 ,
         \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 ,
         \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 ,
         \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 ,
         \13477 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 ,
         \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 ,
         \13497 , \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 ,
         \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 ,
         \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 ,
         \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 ,
         \13537 , \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 ,
         \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 ,
         \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 ,
         \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 ,
         \13577 , \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 , \13585 , \13586 ,
         \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 ,
         \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 ,
         \13607 , \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 ,
         \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 ,
         \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 ,
         \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 ,
         \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 ,
         \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 ,
         \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 , \13675 , \13676 ,
         \13677 , \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685 , \13686 ,
         \13687 , \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 ,
         \13697 , \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705 , \13706 ,
         \13707 , \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 ,
         \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726 ,
         \13727 , \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 , \13735 , \13736 ,
         \13737 , \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 ,
         \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 ,
         \13757 , \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 ,
         \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 ,
         \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 ,
         \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 ,
         \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 ,
         \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 ,
         \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826 ,
         \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 ,
         \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 ,
         \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 ,
         \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 ,
         \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 ,
         \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 ,
         \13887 , \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 ,
         \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 ,
         \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 ,
         \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 ,
         \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 ,
         \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 ,
         \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 , \13955 , \13956 ,
         \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 ,
         \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 ,
         \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 ,
         \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 ,
         \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 ,
         \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 ,
         \14017 , \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 , \14025 , \14026 ,
         \14027 , \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 , \14035 , \14036 ,
         \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 ,
         \14047 , \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 , \14055 , \14056 ,
         \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 ,
         \14067 , \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 ,
         \14077 , \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 ,
         \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 ,
         \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 ,
         \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 ,
         \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 ,
         \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 ,
         \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 ,
         \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 ,
         \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 ,
         \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 ,
         \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 ,
         \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 ,
         \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 ,
         \14207 , \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 , \14215 , \14216 ,
         \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 ,
         \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 ,
         \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 ,
         \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 ,
         \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 ,
         \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 ,
         \14277 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 ,
         \14287 , \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 ,
         \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 ,
         \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 ,
         \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 ,
         \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 ,
         \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 , \14345 , \14346 ,
         \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 ,
         \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 ,
         \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 ,
         \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 ,
         \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 ,
         \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 ,
         \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 , \14415 , \14416 ,
         \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 ,
         \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 ,
         \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 ,
         \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 ,
         \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 ,
         \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 ,
         \14477 , \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 ,
         \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 ,
         \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 ,
         \14507 , \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 ,
         \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 ,
         \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 ,
         \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 ,
         \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 ,
         \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 ,
         \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 ,
         \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 ,
         \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 ,
         \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 ,
         \14607 , \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 , \14615 , \14616 ,
         \14617 , \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 , \14625 , \14626 ,
         \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 , \14635 , \14636 ,
         \14637 , \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 , \14645 , \14646 ,
         \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 , \14655 , \14656 ,
         \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 , \14665 , \14666 ,
         \14667 , \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 , \14675 , \14676 ,
         \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 , \14685 , \14686 ,
         \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 , \14695 , \14696 ,
         \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 ,
         \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 ,
         \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 , \14725 , \14726 ,
         \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 ,
         \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 ,
         \14747 , \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 , \14755 , \14756 ,
         \14757 , \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 , \14765 , \14766 ,
         \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 ,
         \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786 ,
         \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 , \14795 , \14796 ,
         \14797 , \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 , \14805 , \14806 ,
         \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816 ,
         \14817 , \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 ,
         \14827 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 ,
         \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 , \14845 , \14846 ,
         \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 , \14855 , \14856 ,
         \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865 , \14866 ,
         \14867 , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875 , \14876 ,
         \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885 , \14886 ,
         \14887 , \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 , \14895 , \14896 ,
         \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 , \14905 , \14906 ,
         \14907 , \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 ,
         \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 ,
         \14927 , \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 , \14935 , \14936 ,
         \14937 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 ,
         \14947 , \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 , \14955 , \14956 ,
         \14957 , \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 , \14965 , \14966 ,
         \14967 , \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 ,
         \14977 , \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 , \14985 , \14986 ,
         \14987 , \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995 , \14996 ,
         \14997 , \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 , \15005 , \15006 ,
         \15007 , \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 , \15015 , \15016 ,
         \15017 , \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 , \15025 , \15026 ,
         \15027 , \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 , \15035 , \15036 ,
         \15037 , \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 , \15045 , \15046 ,
         \15047 , \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 , \15055 , \15056 ,
         \15057 , \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 ,
         \15067 , \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 , \15075 , \15076 ,
         \15077 , \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 , \15085 , \15086 ,
         \15087 , \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 , \15095 , \15096 ,
         \15097 , \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 , \15105 , \15106 ,
         \15107 , \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115 , \15116 ,
         \15117 , \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 , \15125 , \15126 ,
         \15127 , \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 , \15135 , \15136 ,
         \15137 , \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 , \15145 , \15146 ,
         \15147 , \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 , \15155 , \15156 ,
         \15157 , \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 , \15165 , \15166 ,
         \15167 , \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 , \15175 , \15176 ,
         \15177 , \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 , \15185 , \15186 ,
         \15187 , \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 , \15195 , \15196 ,
         \15197 , \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 , \15205 , \15206 ,
         \15207 , \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 , \15215 , \15216 ,
         \15217 , \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 , \15225 , \15226 ,
         \15227 , \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 , \15235 , \15236 ,
         \15237 , \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 , \15245 , \15246 ,
         \15247 , \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 , \15255 , \15256 ,
         \15257 , \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 , \15265 , \15266 ,
         \15267 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 ,
         \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 , \15285 , \15286 ,
         \15287 , \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 , \15295 , \15296 ,
         \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 ,
         \15307 , \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 , \15315 , \15316 ,
         \15317 , \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 , \15325 , \15326 ,
         \15327 , \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 , \15335 , \15336 ,
         \15337 , \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 , \15345 , \15346 ,
         \15347 , \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 , \15355 , \15356 ,
         \15357 , \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 , \15365 , \15366 ,
         \15367 , \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 , \15375 , \15376 ,
         \15377 , \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 , \15385 , \15386 ,
         \15387 , \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 , \15395 , \15396 ,
         \15397 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 , \15405 , \15406 ,
         \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 , \15415 , \15416 ,
         \15417 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 , \15425 , \15426 ,
         \15427 , \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 , \15435 , \15436 ,
         \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 , \15445 , \15446 ,
         \15447 , \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 , \15455 , \15456 ,
         \15457 , \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 , \15465 , \15466 ,
         \15467 , \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 , \15475 , \15476 ,
         \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 , \15485 , \15486 ,
         \15487 , \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 , \15495 , \15496 ,
         \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 , \15505 , \15506 ,
         \15507 , \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 , \15515 , \15516 ,
         \15517 , \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 , \15525 , \15526 ,
         \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 , \15535 , \15536 ,
         \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 ,
         \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 , \15555 , \15556 ,
         \15557 , \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 , \15565 , \15566 ,
         \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 , \15575 , \15576 ,
         \15577 , \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 , \15585 , \15586 ,
         \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 ,
         \15597 , \15598 , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 , \15605 , \15606 ,
         \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 , \15615 , \15616 ,
         \15617 , \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 , \15625 , \15626 ,
         \15627 , \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 , \15635 , \15636 ,
         \15637 , \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 , \15645 , \15646 ,
         \15647 , \15648 , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 , \15655 , \15656 ,
         \15657 , \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 , \15665 , \15666 ,
         \15667 , \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 , \15675 , \15676 ,
         \15677 , \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 , \15685 , \15686 ,
         \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 , \15696 ,
         \15697 , \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 , \15705 , \15706 ,
         \15707 , \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 , \15715 , \15716 ,
         \15717 , \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 , \15725 , \15726 ,
         \15727 , \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , \15736 ,
         \15737 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 , \15745 , \15746 ,
         \15747 , \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 , \15755 , \15756 ,
         \15757 , \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 , \15765 , \15766 ,
         \15767 , \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 , \15775 , \15776 ,
         \15777 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 , \15785 , \15786 ,
         \15787 , \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 , \15795 , \15796 ,
         \15797 , \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 , \15805 , \15806 ,
         \15807 , \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 , \15815 , \15816 ,
         \15817 , \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 , \15825 , \15826 ,
         \15827 , \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 , \15835 , \15836 ,
         \15837 , \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 , \15845 , \15846 ,
         \15847 , \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 , \15855 , \15856 ,
         \15857 , \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 , \15865 , \15866 ,
         \15867 , \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 , \15875 , \15876 ,
         \15877 , \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 , \15885 , \15886 ,
         \15887 , \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 , \15895 , \15896 ,
         \15897 , \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 , \15905 , \15906 ,
         \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 , \15915 , \15916 ,
         \15917 , \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 , \15925 , \15926 ,
         \15927 , \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 , \15935 , \15936 ,
         \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 , \15945 , \15946 ,
         \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 , \15955 , \15956 ,
         \15957 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 , \15965 , \15966 ,
         \15967 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 , \15975 , \15976 ,
         \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 , \15985 , \15986 ,
         \15987 , \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 , \15995 , \15996 ,
         \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 , \16006 ,
         \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 , \16015 , \16016 ,
         \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 ,
         \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 ,
         \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 , \16045 , \16046 ,
         \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 , \16055 , \16056 ,
         \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 , \16066 ,
         \16067 , \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 , \16075 , \16076 ,
         \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 ,
         \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 , \16095 , \16096 ,
         \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 ,
         \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 , \16115 , \16116 ,
         \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 , \16125 , \16126 ,
         \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 , \16135 , \16136 ,
         \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 ,
         \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 , \16155 , \16156 ,
         \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 ,
         \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 , \16176 ,
         \16177 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 ,
         \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 , \16195 , \16196 ,
         \16197 , \16198 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 , \16205 , \16206 ,
         \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 , \16216 ,
         \16217 , \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 , \16225 , \16226 ,
         \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 , \16235 , \16236 ,
         \16237 , \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 , \16245 , \16246 ,
         \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 ,
         \16257 , \16258 , \16259 , \16260 , \16261 , \16262 , \16263 , \16264 , \16265 , \16266 ,
         \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 , \16275 , \16276 ,
         \16277 , \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 , \16285 , \16286 ,
         \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 , \16295 , \16296 ,
         \16297 , \16298 , \16299 , \16300 , \16301 , \16302 , \16303 , \16304 , \16305 , \16306 ,
         \16307 , \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 , \16315 , \16316 ,
         \16317 , \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 , \16325 , \16326 ,
         \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 , \16335 , \16336 ,
         \16337 , \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 , \16345 , \16346 ,
         \16347 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 , \16355 , \16356 ,
         \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 , \16365 , \16366 ,
         \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 , \16375 , \16376 ,
         \16377 , \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 , \16385 , \16386 ,
         \16387 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 , \16395 , \16396 ,
         \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 , \16405 , \16406 ,
         \16407 , \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 , \16415 , \16416 ,
         \16417 , \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 , \16425 , \16426 ,
         \16427 , \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 , \16435 , \16436 ,
         \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 , \16445 , \16446 ,
         \16447 , \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 , \16455 , \16456 ,
         \16457 , \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 , \16465 , \16466 ,
         \16467 , \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 , \16475 , \16476 ,
         \16477 , \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 , \16485 , \16486 ,
         \16487 , \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 , \16495 , \16496 ,
         \16497 , \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 , \16505 , \16506 ,
         \16507 , \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 , \16515 , \16516 ,
         \16517 , \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 , \16525 , \16526 ,
         \16527 , \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 , \16535 , \16536 ,
         \16537 , \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 , \16545 , \16546 ,
         \16547 , \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 , \16555 , \16556 ,
         \16557 , \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 , \16565 , \16566 ,
         \16567 , \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 , \16575 , \16576 ,
         \16577 , \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 , \16585 , \16586 ,
         \16587 , \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 , \16595 , \16596 ,
         \16597 , \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 , \16605 , \16606 ,
         \16607 , \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 , \16615 , \16616 ,
         \16617 , \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 , \16625 , \16626 ,
         \16627 , \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 , \16635 , \16636 ,
         \16637 , \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 , \16645 , \16646 ,
         \16647 , \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 , \16655 , \16656 ,
         \16657 , \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 , \16665 , \16666 ,
         \16667 , \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 , \16675 , \16676 ,
         \16677 , \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684 , \16685 , \16686 ,
         \16687 , \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 , \16695 , \16696 ,
         \16697 , \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 , \16705 , \16706 ,
         \16707 , \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 , \16715 , \16716 ,
         \16717 , \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 , \16725 , \16726 ,
         \16727 , \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 , \16735 , \16736 ,
         \16737 , \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 , \16745 , \16746 ,
         \16747 , \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 , \16755 , \16756 ,
         \16757 , \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 , \16765 , \16766 ,
         \16767 , \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 , \16775 , \16776 ,
         \16777 , \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 , \16785 , \16786 ,
         \16787 , \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 , \16795 , \16796 ,
         \16797 , \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 , \16805 , \16806 ,
         \16807 , \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 , \16815 , \16816 ,
         \16817 , \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 , \16825 , \16826 ,
         \16827 , \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 , \16835 , \16836 ,
         \16837 , \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 , \16845 , \16846 ,
         \16847 , \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 , \16855 , \16856 ,
         \16857 , \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 , \16865 , \16866 ,
         \16867 , \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 , \16875 , \16876 ,
         \16877 , \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 , \16885 , \16886 ,
         \16887 , \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 , \16895 , \16896 ,
         \16897 , \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 , \16905 , \16906 ,
         \16907 , \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 , \16915 , \16916 ,
         \16917 , \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 , \16925 , \16926 ,
         \16927 , \16928 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 , \16935 , \16936 ,
         \16937 , \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 , \16945 , \16946 ,
         \16947 , \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954 , \16955 , \16956 ,
         \16957 , \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 , \16965 , \16966 ,
         \16967 , \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 , \16975 , \16976 ,
         \16977 , \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 , \16985 , \16986 ,
         \16987 , \16988 , \16989 , \16990 , \16991 , \16992 , \16993 , \16994 , \16995 , \16996 ,
         \16997 , \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 , \17005 , \17006 ,
         \17007 , \17008 , \17009 , \17010 , \17011 , \17012 , \17013 , \17014 , \17015 , \17016 ,
         \17017 , \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 , \17025 , \17026 ,
         \17027 , \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 , \17035 , \17036 ,
         \17037 , \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 , \17045 , \17046 ,
         \17047 , \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 , \17055 , \17056 ,
         \17057 , \17058 , \17059 , \17060 , \17061 , \17062 , \17063 , \17064 , \17065 , \17066 ,
         \17067 , \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 , \17075 , \17076 ,
         \17077 , \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084 , \17085 , \17086 ,
         \17087 , \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 , \17095 , \17096 ,
         \17097 , \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 , \17105 , \17106 ,
         \17107 , \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 , \17115 , \17116 ,
         \17117 , \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 , \17125 , \17126 ,
         \17127 , \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 , \17135 , \17136 ,
         \17137 , \17138 , \17139 , \17140 , \17141 , \17142 , \17143 , \17144 , \17145 , \17146 ,
         \17147 , \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 , \17155 , \17156 ,
         \17157 , \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 , \17165 , \17166 ,
         \17167 , \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 , \17175 , \17176 ,
         \17177 , \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 , \17185 , \17186 ,
         \17187 , \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 , \17195 , \17196 ,
         \17197 , \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 , \17205 , \17206 ,
         \17207 , \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 , \17215 , \17216 ,
         \17217 , \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 , \17225 , \17226 ,
         \17227 , \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 , \17235 , \17236 ,
         \17237 , \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 , \17245 , \17246 ,
         \17247 , \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 , \17255 , \17256 ,
         \17257 , \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 , \17265 , \17266 ,
         \17267 , \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 , \17275 , \17276 ,
         \17277 , \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 , \17285 , \17286 ,
         \17287 , \17288 , \17289 , \17290 , \17291 , \17292 , \17293 , \17294 , \17295 , \17296 ,
         \17297 , \17298 , \17299 , \17300 , \17301 , \17302 , \17303 , \17304 , \17305 , \17306 ,
         \17307 , \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 , \17315 , \17316 ,
         \17317 , \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 , \17325 , \17326 ,
         \17327 , \17328 , \17329 , \17330 , \17331 , \17332 , \17333 , \17334 , \17335 , \17336 ,
         \17337 , \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 , \17345 , \17346 ,
         \17347 , \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 , \17355 , \17356 ,
         \17357 , \17358 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 , \17365 , \17366 ,
         \17367 , \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 , \17375 , \17376 ,
         \17377 , \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 , \17385 , \17386 ,
         \17387 , \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 , \17395 , \17396 ,
         \17397 , \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 , \17405 , \17406 ,
         \17407 , \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 , \17415 , \17416 ,
         \17417 , \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 , \17425 , \17426 ,
         \17427 , \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 , \17435 , \17436 ,
         \17437 , \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 , \17445 , \17446 ,
         \17447 , \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 , \17455 , \17456 ,
         \17457 , \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 , \17465 , \17466 ,
         \17467 , \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 , \17475 , \17476 ,
         \17477 , \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 , \17485 , \17486 ,
         \17487 , \17488 , \17489 , \17490 , \17491 , \17492 , \17493 , \17494 , \17495 , \17496 ,
         \17497 , \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 , \17505 , \17506 ,
         \17507 , \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 , \17515 , \17516 ,
         \17517 , \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 , \17525 , \17526 ,
         \17527 , \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 , \17535 , \17536 ,
         \17537 , \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 , \17545 , \17546 ,
         \17547 , \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 , \17555 , \17556 ,
         \17557 , \17558 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 , \17565 , \17566 ,
         \17567 , \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 , \17575 , \17576 ,
         \17577 , \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 , \17585 , \17586 ,
         \17587 , \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 , \17595 , \17596 ,
         \17597 , \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 , \17605 , \17606 ,
         \17607 , \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 , \17615 , \17616 ,
         \17617 , \17618 , \17619 , \17620 , \17621 , \17622 , \17623 , \17624 , \17625 , \17626 ,
         \17627 , \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 , \17635 , \17636 ,
         \17637 , \17638 , \17639 , \17640 , \17641 , \17642 , \17643 , \17644 , \17645 , \17646 ,
         \17647 , \17648 , \17649 , \17650 , \17651 , \17652 , \17653 , \17654 , \17655 , \17656 ,
         \17657 , \17658 , \17659 , \17660 , \17661 , \17662 , \17663 , \17664 , \17665 , \17666 ,
         \17667 , \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 , \17675 , \17676 ,
         \17677 , \17678 , \17679 , \17680 , \17681 , \17682 , \17683 , \17684 , \17685 , \17686 ,
         \17687 , \17688 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 , \17695 , \17696 ,
         \17697 , \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 , \17705 , \17706 ,
         \17707 , \17708 , \17709 , \17710 , \17711 , \17712 , \17713 , \17714 , \17715 , \17716 ,
         \17717 , \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 , \17725 , \17726 ,
         \17727 , \17728 , \17729 , \17730 , \17731 , \17732 , \17733 , \17734 , \17735 , \17736 ,
         \17737 , \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 , \17745 , \17746 ,
         \17747 , \17748 , \17749 , \17750 , \17751 , \17752 , \17753 , \17754 , \17755 , \17756 ,
         \17757 , \17758 , \17759 , \17760 , \17761 , \17762 , \17763 , \17764 , \17765 , \17766 ,
         \17767 , \17768 , \17769 , \17770 , \17771 , \17772 , \17773 , \17774 , \17775 , \17776 ,
         \17777 , \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 , \17785 , \17786 ,
         \17787 , \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 , \17795 , \17796 ,
         \17797 , \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 , \17805 , \17806 ,
         \17807 , \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 , \17815 , \17816 ,
         \17817 , \17818 , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 , \17825 , \17826 ,
         \17827 , \17828 , \17829 , \17830 , \17831 , \17832 , \17833 , \17834 , \17835 , \17836 ,
         \17837 , \17838 , \17839 , \17840 , \17841 , \17842 , \17843 , \17844 , \17845 , \17846 ,
         \17847 , \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854 , \17855 , \17856 ,
         \17857 , \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 , \17865 , \17866 ,
         \17867 , \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 , \17875 , \17876 ,
         \17877 , \17878 , \17879 , \17880 , \17881 , \17882 , \17883 , \17884 , \17885 , \17886 ,
         \17887 , \17888 , \17889 , \17890 , \17891 , \17892 , \17893 , \17894 , \17895 , \17896 ,
         \17897 , \17898 , \17899 , \17900 , \17901 , \17902 , \17903 , \17904 , \17905 , \17906 ,
         \17907 , \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 , \17915 , \17916 ,
         \17917 , \17918 , \17919 , \17920 , \17921 , \17922 , \17923 , \17924 , \17925 , \17926 ,
         \17927 , \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934 , \17935 , \17936 ,
         \17937 , \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 , \17945 , \17946 ,
         \17947 , \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 , \17955 , \17956 ,
         \17957 , \17958 , \17959 , \17960 , \17961 , \17962 , \17963 , \17964 , \17965 , \17966 ,
         \17967 , \17968 , \17969 , \17970 , \17971 , \17972 , \17973 , \17974 , \17975 , \17976 ,
         \17977 , \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 , \17985 , \17986 ,
         \17987 , \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 , \17995 , \17996 ,
         \17997 , \17998 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 , \18005 , \18006 ,
         \18007 , \18008 , \18009 , \18010 , \18011 , \18012 , \18013 , \18014 , \18015 , \18016 ,
         \18017 , \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024 , \18025 , \18026 ,
         \18027 , \18028 , \18029 , \18030 , \18031 , \18032 , \18033 , \18034 , \18035 , \18036 ,
         \18037 , \18038 , \18039 , \18040 , \18041 , \18042 , \18043 , \18044 , \18045 , \18046 ,
         \18047 , \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 , \18055 , \18056 ,
         \18057 , \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 , \18065 , \18066 ,
         \18067 , \18068 , \18069 , \18070 , \18071 , \18072 , \18073 , \18074 , \18075 , \18076 ,
         \18077 , \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 , \18085 , \18086 ,
         \18087 , \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 , \18095 , \18096 ,
         \18097 , \18098 , \18099 , \18100 , \18101 , \18102 , \18103 , \18104 , \18105 , \18106 ,
         \18107 , \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 , \18115 , \18116 ,
         \18117 , \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 , \18125 , \18126 ,
         \18127 , \18128 , \18129 , \18130 , \18131 , \18132 , \18133 , \18134 , \18135 , \18136 ,
         \18137 , \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 , \18145 , \18146 ,
         \18147 , \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 , \18155 , \18156 ,
         \18157 , \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 , \18165 , \18166 ,
         \18167 , \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 , \18175 , \18176 ,
         \18177 , \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 , \18185 , \18186 ,
         \18187 , \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 , \18195 , \18196 ,
         \18197 , \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 , \18205 , \18206 ,
         \18207 , \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 , \18215 , \18216 ,
         \18217 , \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 , \18225 , \18226 ,
         \18227 , \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 , \18235 , \18236 ,
         \18237 , \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 , \18245 , \18246 ,
         \18247 , \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 , \18255 , \18256 ,
         \18257 , \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 , \18265 , \18266 ,
         \18267 , \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 , \18275 , \18276 ,
         \18277 , \18278 , \18279 , \18280 , \18281 , \18282 , \18283 , \18284 , \18285 , \18286 ,
         \18287 , \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 , \18295 , \18296 ,
         \18297 , \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 , \18305 , \18306 ,
         \18307 , \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 , \18315 , \18316 ,
         \18317 , \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 , \18325 , \18326 ,
         \18327 , \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 , \18335 , \18336 ,
         \18337 , \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 , \18345 , \18346 ,
         \18347 , \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 , \18355 , \18356 ,
         \18357 , \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 , \18365 , \18366 ,
         \18367 , \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 , \18375 , \18376 ,
         \18377 , \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 , \18385 , \18386 ,
         \18387 , \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 , \18395 , \18396 ,
         \18397 , \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 , \18405 , \18406 ,
         \18407 , \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 , \18415 , \18416 ,
         \18417 , \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 , \18425 , \18426 ,
         \18427 , \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 , \18435 , \18436 ,
         \18437 , \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 , \18445 , \18446 ,
         \18447 , \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 , \18455 , \18456 ,
         \18457 , \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 , \18465 , \18466 ,
         \18467 , \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 , \18475 , \18476 ,
         \18477 , \18478 , \18479 , \18480 , \18481 , \18482 , \18483 , \18484 , \18485 , \18486 ,
         \18487 , \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 , \18495 , \18496 ,
         \18497 , \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 , \18505 , \18506 ,
         \18507 , \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 , \18515 , \18516 ,
         \18517 , \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 , \18525 , \18526 ,
         \18527 , \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 , \18535 , \18536 ,
         \18537 , \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 , \18545 , \18546 ,
         \18547 , \18548 , \18549 , \18550 , \18551 , \18552 , \18553 , \18554 , \18555 , \18556 ,
         \18557 , \18558 , \18559 , \18560 , \18561 , \18562 , \18563 , \18564 , \18565 , \18566 ,
         \18567 , \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 , \18575 , \18576 ,
         \18577 , \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 , \18585 , \18586 ,
         \18587 , \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 , \18595 , \18596 ,
         \18597 , \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 , \18605 , \18606 ,
         \18607 , \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 , \18615 , \18616 ,
         \18617 , \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 , \18625 , \18626 ,
         \18627 , \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 , \18635 , \18636 ,
         \18637 , \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 , \18645 , \18646 ,
         \18647 , \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 , \18655 , \18656 ,
         \18657 , \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 , \18665 , \18666 ,
         \18667 , \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 , \18675 , \18676 ,
         \18677 , \18678 , \18679 , \18680 , \18681 , \18682 , \18683 , \18684 , \18685 , \18686 ,
         \18687 , \18688 , \18689 , \18690 , \18691 , \18692 , \18693 , \18694 , \18695 , \18696 ,
         \18697 , \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 , \18705 , \18706 ,
         \18707 , \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 , \18715 , \18716 ,
         \18717 , \18718 , \18719 , \18720 , \18721 , \18722 , \18723 , \18724 , \18725 , \18726 ,
         \18727 , \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 , \18735 , \18736 ,
         \18737 , \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 , \18745 , \18746 ,
         \18747 , \18748 , \18749 , \18750 , \18751 , \18752 , \18753 , \18754 , \18755 , \18756 ,
         \18757 , \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 , \18765 , \18766 ,
         \18767 , \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 , \18775 , \18776 ,
         \18777 , \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 , \18785 , \18786 ,
         \18787 , \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 , \18795 , \18796 ,
         \18797 , \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 , \18805 , \18806 ,
         \18807 , \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 , \18815 , \18816 ,
         \18817 , \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 , \18825 , \18826 ,
         \18827 , \18828 , \18829 , \18830 , \18831 , \18832 , \18833 , \18834 , \18835 , \18836 ,
         \18837 , \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 , \18845 , \18846 ,
         \18847 , \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 , \18855 , \18856 ,
         \18857 , \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 , \18865 , \18866 ,
         \18867 , \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 , \18875 , \18876 ,
         \18877 , \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 , \18885 , \18886 ,
         \18887 , \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 , \18895 , \18896 ,
         \18897 , \18898 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 , \18905 , \18906 ,
         \18907 , \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 , \18915 , \18916 ,
         \18917 , \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 , \18925 , \18926 ,
         \18927 , \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 , \18935 , \18936 ,
         \18937 , \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 , \18945 , \18946 ,
         \18947 , \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 , \18955 , \18956 ,
         \18957 , \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 , \18965 , \18966 ,
         \18967 , \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 , \18975 , \18976 ,
         \18977 , \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 , \18985 , \18986 ,
         \18987 , \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 , \18995 , \18996 ,
         \18997 , \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 , \19005 , \19006 ,
         \19007 , \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 , \19015 , \19016 ,
         \19017 , \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 , \19025 , \19026 ,
         \19027 , \19028 , \19029 , \19030 , \19031 , \19032 , \19033 , \19034 , \19035 , \19036 ,
         \19037 , \19038 , \19039 , \19040 , \19041 , \19042 , \19043 , \19044 , \19045 , \19046 ,
         \19047 , \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 , \19055 , \19056 ,
         \19057 , \19058 , \19059 , \19060 , \19061 , \19062 , \19063 , \19064 , \19065 , \19066 ,
         \19067 , \19068 , \19069 , \19070 , \19071 , \19072 , \19073 , \19074 , \19075 , \19076 ,
         \19077 , \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 , \19085 , \19086 ,
         \19087 , \19088 , \19089 , \19090 , \19091 , \19092 , \19093 , \19094 , \19095 , \19096 ,
         \19097 , \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 , \19105 , \19106 ,
         \19107 , \19108 , \19109 , \19110 , \19111 , \19112 , \19113 , \19114 , \19115 , \19116 ,
         \19117 , \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 , \19125 , \19126 ,
         \19127 , \19128 , \19129 , \19130 , \19131 , \19132 , \19133 , \19134 , \19135 , \19136 ,
         \19137 , \19138 , \19139 , \19140 , \19141 , \19142 , \19143 , \19144 , \19145 , \19146 ,
         \19147 , \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 , \19155 , \19156 ,
         \19157 , \19158 , \19159 , \19160 , \19161 , \19162 , \19163 , \19164 , \19165 , \19166 ,
         \19167 , \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 , \19175 , \19176 ,
         \19177 , \19178 , \19179 , \19180 , \19181 , \19182 , \19183 , \19184 , \19185 , \19186 ,
         \19187 , \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 , \19195 , \19196 ,
         \19197 , \19198 , \19199 , \19200 , \19201 , \19202 , \19203 , \19204 , \19205 , \19206 ,
         \19207 , \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 , \19215 , \19216 ,
         \19217 , \19218 , \19219 , \19220 , \19221 , \19222 , \19223 , \19224 , \19225 , \19226 ,
         \19227 , \19228 , \19229 , \19230 , \19231 , \19232 , \19233 , \19234 , \19235 , \19236 ,
         \19237 , \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 , \19245 , \19246 ,
         \19247 , \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 , \19255 , \19256 ,
         \19257 , \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 , \19265 , \19266 ,
         \19267 , \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 , \19275 , \19276 ,
         \19277 , \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 , \19285 , \19286 ,
         \19287 , \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 , \19295 , \19296 ,
         \19297 , \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 , \19305 , \19306 ,
         \19307 , \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 , \19315 , \19316 ,
         \19317 , \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 , \19325 , \19326 ,
         \19327 , \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 , \19335 , \19336 ,
         \19337 , \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 , \19345 , \19346 ,
         \19347 , \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 , \19355 , \19356 ,
         \19357 , \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 , \19365 , \19366 ,
         \19367 , \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 , \19375 , \19376 ,
         \19377 , \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 , \19385 , \19386 ,
         \19387 , \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 , \19395 , \19396 ,
         \19397 , \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 , \19405 , \19406 ,
         \19407 , \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 , \19415 , \19416 ,
         \19417 , \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 , \19425 , \19426 ,
         \19427 , \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 , \19435 , \19436 ,
         \19437 , \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 , \19445 , \19446 ,
         \19447 , \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 , \19455 , \19456 ,
         \19457 , \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 , \19465 , \19466 ,
         \19467 , \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 , \19475 , \19476 ,
         \19477 , \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 , \19485 , \19486 ,
         \19487 , \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 , \19495 , \19496 ,
         \19497 , \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 , \19505 , \19506 ,
         \19507 , \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 , \19515 , \19516 ,
         \19517 , \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 , \19525 , \19526 ,
         \19527 , \19528 , \19529 , \19530 , \19531 , \19532 , \19533 , \19534 , \19535 , \19536 ,
         \19537 , \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 , \19545 , \19546 ,
         \19547 , \19548 , \19549 , \19550 , \19551 , \19552 , \19553 , \19554 , \19555 , \19556 ,
         \19557 , \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 , \19565 , \19566 ,
         \19567 , \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 , \19575 , \19576 ,
         \19577 , \19578 , \19579 , \19580 , \19581 , \19582 , \19583 , \19584 , \19585 , \19586 ,
         \19587 , \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 , \19595 , \19596 ,
         \19597 , \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 , \19605 , \19606 ,
         \19607 , \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 , \19615 , \19616 ,
         \19617 , \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 , \19625 , \19626 ,
         \19627 , \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 , \19635 , \19636 ,
         \19637 , \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 , \19645 , \19646 ,
         \19647 , \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 , \19655 , \19656 ,
         \19657 , \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 , \19665 , \19666 ,
         \19667 , \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 , \19675 , \19676 ,
         \19677 , \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 , \19685 , \19686 ,
         \19687 , \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 , \19695 , \19696 ,
         \19697 , \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 , \19705 , \19706 ,
         \19707 , \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 , \19715 , \19716 ,
         \19717 , \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 , \19725 , \19726 ,
         \19727 , \19728 , \19729 , \19730 , \19731 , \19732 , \19733 , \19734 , \19735 , \19736 ,
         \19737 , \19738 , \19739 , \19740 , \19741 , \19742 , \19743 , \19744 , \19745 , \19746 ,
         \19747 , \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 , \19755 , \19756 ,
         \19757 , \19758 , \19759 , \19760 , \19761 , \19762 , \19763 , \19764 , \19765 , \19766 ,
         \19767 , \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 , \19775 , \19776 ,
         \19777 , \19778 , \19779 , \19780 , \19781 , \19782 , \19783 , \19784 , \19785 , \19786 ,
         \19787 , \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 , \19795 , \19796 ,
         \19797 , \19798 , \19799 , \19800 , \19801 , \19802 , \19803 , \19804 , \19805 , \19806 ,
         \19807 , \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 , \19815 , \19816 ,
         \19817 , \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 , \19825 , \19826 ,
         \19827 , \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 , \19835 , \19836 ,
         \19837 , \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 , \19845 , \19846 ,
         \19847 , \19848 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 , \19855 , \19856 ,
         \19857 , \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 , \19865 , \19866 ,
         \19867 , \19868 , \19869 , \19870 , \19871 , \19872 , \19873 , \19874 , \19875 , \19876 ,
         \19877 , \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 , \19885 , \19886 ,
         \19887 , \19888 , \19889 , \19890 , \19891 , \19892 , \19893 , \19894 , \19895 , \19896 ,
         \19897 , \19898 , \19899 , \19900 , \19901 , \19902 , \19903 , \19904 , \19905 , \19906 ,
         \19907 , \19908 , \19909 , \19910 , \19911 , \19912 , \19913 , \19914 , \19915 , \19916 ,
         \19917 , \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 , \19925 , \19926 ,
         \19927 , \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 , \19935 , \19936 ,
         \19937 , \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 , \19945 , \19946 ,
         \19947 , \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 , \19955 , \19956 ,
         \19957 , \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964 , \19965 , \19966 ,
         \19967 , \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 , \19975 , \19976 ,
         \19977 , \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 , \19985 , \19986 ,
         \19987 , \19988 , \19989 , \19990 , \19991 , \19992 , \19993 , \19994 , \19995 , \19996 ,
         \19997 , \19998 , \19999 , \20000 , \20001 , \20002 , \20003 , \20004 , \20005 , \20006 ,
         \20007 , \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 , \20015 , \20016 ,
         \20017 , \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 , \20025 , \20026 ,
         \20027 , \20028 , \20029 , \20030 , \20031 , \20032 , \20033 , \20034 , \20035 , \20036 ,
         \20037 , \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 , \20045 , \20046 ,
         \20047 , \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 , \20055 , \20056 ,
         \20057 , \20058 , \20059 , \20060 , \20061 , \20062 , \20063 , \20064 , \20065 , \20066 ,
         \20067 , \20068 , \20069 , \20070 , \20071 , \20072 , \20073 , \20074 , \20075 , \20076 ,
         \20077 , \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 , \20085 , \20086 ,
         \20087 , \20088 , \20089 , \20090 , \20091 , \20092 , \20093 , \20094 , \20095 , \20096 ,
         \20097 , \20098 , \20099 , \20100 , \20101 , \20102 , \20103 , \20104 , \20105 , \20106 ,
         \20107 , \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 , \20115 , \20116 ,
         \20117 , \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 , \20125 , \20126 ,
         \20127 , \20128 , \20129 , \20130 , \20131 , \20132 , \20133 , \20134 , \20135 , \20136 ,
         \20137 , \20138 , \20139 , \20140 , \20141 , \20142 , \20143 , \20144 , \20145 , \20146 ,
         \20147 , \20148 , \20149 , \20150 , \20151 , \20152 , \20153 , \20154 , \20155 , \20156 ,
         \20157 , \20158 , \20159 , \20160 , \20161 , \20162 , \20163 , \20164 , \20165 , \20166 ,
         \20167 , \20168 , \20169 , \20170 , \20171 , \20172 , \20173 , \20174 , \20175 , \20176 ,
         \20177 , \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 , \20185 , \20186 ,
         \20187 , \20188 , \20189 , \20190 , \20191 , \20192 , \20193 , \20194 , \20195 , \20196 ,
         \20197 , \20198 , \20199 , \20200 , \20201 , \20202 , \20203 , \20204 , \20205 , \20206 ,
         \20207 , \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 , \20215 , \20216 ,
         \20217 , \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 , \20225 , \20226 ,
         \20227 , \20228 , \20229 , \20230 , \20231 , \20232 , \20233 , \20234 , \20235 , \20236 ,
         \20237 , \20238 , \20239 , \20240 , \20241 , \20242 , \20243 , \20244 , \20245 , \20246 ,
         \20247 , \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 , \20255 , \20256 ,
         \20257 , \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 , \20265 , \20266 ,
         \20267 , \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 , \20275 , \20276 ,
         \20277 , \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 , \20285 , \20286 ,
         \20287 , \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 , \20295 , \20296 ,
         \20297 , \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 , \20305 , \20306 ,
         \20307 , \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 , \20315 , \20316 ,
         \20317 , \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 , \20325 , \20326 ,
         \20327 , \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 , \20335 , \20336 ,
         \20337 , \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 , \20345 , \20346 ,
         \20347 , \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 , \20355 , \20356 ,
         \20357 , \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 , \20365 , \20366 ,
         \20367 , \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 , \20375 , \20376 ,
         \20377 , \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 , \20385 , \20386 ,
         \20387 , \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 , \20395 , \20396 ,
         \20397 , \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 , \20405 , \20406 ,
         \20407 , \20408 , \20409 , \20410 , \20411 , \20412 , \20413 , \20414 , \20415 , \20416 ,
         \20417 , \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 , \20425 , \20426 ,
         \20427 , \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 , \20435 , \20436 ,
         \20437 , \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 , \20445 , \20446 ,
         \20447 , \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 , \20455 , \20456 ,
         \20457 , \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 , \20465 , \20466 ,
         \20467 , \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 , \20475 , \20476 ,
         \20477 , \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 , \20485 , \20486 ,
         \20487 , \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 , \20495 , \20496 ,
         \20497 , \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 , \20505 , \20506 ,
         \20507 , \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 , \20515 , \20516 ,
         \20517 , \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 , \20525 , \20526 ,
         \20527 , \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 , \20535 , \20536 ,
         \20537 , \20538 , \20539 , \20540 , \20541 , \20542 , \20543 , \20544 , \20545 , \20546 ,
         \20547 , \20548 , \20549 , \20550 , \20551 , \20552 , \20553 , \20554 , \20555 , \20556 ,
         \20557 , \20558 , \20559 , \20560 , \20561 , \20562 , \20563 , \20564 , \20565 , \20566 ,
         \20567 , \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 , \20575 , \20576 ,
         \20577 , \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 , \20585 , \20586 ,
         \20587 , \20588 , \20589 , \20590 , \20591 , \20592 , \20593 , \20594 , \20595 , \20596 ,
         \20597 , \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 , \20605 , \20606 ,
         \20607 , \20608 , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 , \20615 , \20616 ,
         \20617 , \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 , \20625 , \20626 ,
         \20627 , \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 , \20635 , \20636 ,
         \20637 , \20638 , \20639 , \20640 , \20641 , \20642 , \20643 , \20644 , \20645 , \20646 ,
         \20647 , \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 , \20655 , \20656 ,
         \20657 , \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 , \20665 , \20666 ,
         \20667 , \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 , \20675 , \20676 ,
         \20677 , \20678 , \20679 , \20680 , \20681 , \20682 , \20683 , \20684 , \20685 , \20686 ,
         \20687 , \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 , \20695 , \20696 ,
         \20697 , \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 , \20705 , \20706 ,
         \20707 , \20708 , \20709 , \20710 , \20711 , \20712 , \20713 , \20714 , \20715 , \20716 ,
         \20717 , \20718 , \20719 , \20720 , \20721 , \20722 , \20723 , \20724 , \20725 , \20726 ,
         \20727 , \20728 , \20729 , \20730 , \20731 , \20732 , \20733 , \20734 , \20735 , \20736 ,
         \20737 , \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 , \20745 , \20746 ,
         \20747 , \20748 , \20749 , \20750 , \20751 , \20752 , \20753 , \20754 , \20755 , \20756 ,
         \20757 , \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 , \20765 , \20766 ,
         \20767 , \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 , \20775 , \20776 ,
         \20777 , \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 , \20785 , \20786 ,
         \20787 , \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 , \20795 , \20796 ,
         \20797 , \20798 , \20799 , \20800 , \20801 , \20802 , \20803 , \20804 , \20805 , \20806 ,
         \20807 , \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 , \20815 , \20816 ,
         \20817 , \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 , \20825 , \20826 ,
         \20827 , \20828 , \20829 , \20830 , \20831 , \20832 , \20833 , \20834 , \20835 , \20836 ,
         \20837 , \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 , \20845 , \20846 ,
         \20847 , \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 , \20855 , \20856 ,
         \20857 , \20858 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 , \20865 , \20866 ,
         \20867 , \20868 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 , \20875 , \20876 ,
         \20877 , \20878 , \20879 , \20880 , \20881 , \20882 , \20883 , \20884 , \20885 , \20886 ,
         \20887 , \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 , \20895 , \20896 ,
         \20897 , \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 , \20905 , \20906 ,
         \20907 , \20908 , \20909 , \20910 , \20911 , \20912 , \20913 , \20914 , \20915 , \20916 ,
         \20917 , \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 , \20925 , \20926 ,
         \20927 , \20928 , \20929 , \20930 , \20931 , \20932 , \20933 , \20934 , \20935 , \20936 ,
         \20937 , \20938 , \20939 , \20940 , \20941 , \20942 , \20943 , \20944 , \20945 , \20946 ,
         \20947 , \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 , \20955 , \20956 ,
         \20957 , \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 , \20965 , \20966 ,
         \20967 , \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 , \20975 , \20976 ,
         \20977 , \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 , \20985 , \20986 ,
         \20987 , \20988 , \20989 , \20990 , \20991 , \20992 , \20993 , \20994 , \20995 , \20996 ,
         \20997 , \20998 , \20999 , \21000 , \21001 , \21002 , \21003 , \21004 , \21005 , \21006 ,
         \21007 , \21008 , \21009 , \21010 , \21011 , \21012 , \21013 , \21014 , \21015 , \21016 ,
         \21017 , \21018 , \21019 , \21020 , \21021 , \21022 , \21023 , \21024 , \21025 , \21026 ,
         \21027 , \21028 , \21029 , \21030 , \21031 , \21032 , \21033 , \21034 , \21035 , \21036 ,
         \21037 , \21038 , \21039 , \21040 , \21041 , \21042 , \21043 , \21044 , \21045 , \21046 ,
         \21047 , \21048 , \21049 , \21050 , \21051 , \21052 , \21053 , \21054 , \21055 , \21056 ,
         \21057 , \21058 , \21059 , \21060 , \21061 , \21062 , \21063 , \21064 , \21065 , \21066 ,
         \21067 , \21068 , \21069 , \21070 , \21071 , \21072 , \21073 , \21074 , \21075 , \21076 ,
         \21077 , \21078 , \21079 , \21080 , \21081 , \21082 , \21083 , \21084 , \21085 , \21086 ,
         \21087 , \21088 , \21089 , \21090 , \21091 , \21092 , \21093 , \21094 , \21095 , \21096 ,
         \21097 , \21098 , \21099 , \21100 , \21101 , \21102 , \21103 , \21104 , \21105 , \21106 ,
         \21107 , \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 , \21115 , \21116 ,
         \21117 , \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 , \21125 , \21126 ,
         \21127 , \21128 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 , \21135 , \21136 ,
         \21137 , \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 , \21145 , \21146 ,
         \21147 , \21148 , \21149 , \21150 , \21151 , \21152 , \21153 , \21154 , \21155 , \21156 ,
         \21157 , \21158 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 , \21165 , \21166 ,
         \21167 , \21168 , \21169 , \21170 , \21171 , \21172 , \21173 , \21174 , \21175 , \21176 ,
         \21177 , \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 , \21185 , \21186 ,
         \21187 , \21188 , \21189 , \21190 , \21191 , \21192 , \21193 , \21194 , \21195 , \21196 ,
         \21197 , \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 , \21205 , \21206 ,
         \21207 , \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 , \21215 , \21216 ,
         \21217 , \21218 , \21219 , \21220 , \21221 , \21222 , \21223 , \21224 , \21225 , \21226 ,
         \21227 , \21228 , \21229 , \21230 , \21231 , \21232 , \21233 , \21234 , \21235 , \21236 ,
         \21237 , \21238 , \21239 , \21240 , \21241 , \21242 , \21243 , \21244 , \21245 , \21246 ,
         \21247 , \21248 , \21249 , \21250 , \21251 , \21252 , \21253 , \21254 , \21255 , \21256 ,
         \21257 , \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 , \21265 , \21266 ,
         \21267 , \21268 , \21269 , \21270 , \21271 , \21272 , \21273 , \21274 , \21275 , \21276 ,
         \21277 , \21278 , \21279 , \21280 , \21281 , \21282 , \21283 , \21284 , \21285 , \21286 ,
         \21287 , \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 , \21295 , \21296 ,
         \21297 , \21298 , \21299 , \21300 , \21301 , \21302 , \21303 , \21304 , \21305 , \21306 ,
         \21307 , \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 , \21315 , \21316 ,
         \21317 , \21318 , \21319 , \21320 , \21321 , \21322 , \21323 , \21324 , \21325 , \21326 ,
         \21327 , \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 , \21335 , \21336 ,
         \21337 , \21338 , \21339 , \21340 , \21341 , \21342 , \21343 , \21344 , \21345 , \21346 ,
         \21347 , \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 , \21355 , \21356 ,
         \21357 , \21358 , \21359 , \21360 , \21361 , \21362 , \21363 , \21364 , \21365 , \21366 ,
         \21367 , \21368 , \21369 , \21370 , \21371 , \21372 , \21373 , \21374 , \21375 , \21376 ,
         \21377 , \21378 , \21379 , \21380 , \21381 , \21382 , \21383 , \21384 , \21385 , \21386 ,
         \21387 , \21388 , \21389 , \21390 , \21391 , \21392 , \21393 , \21394 , \21395 , \21396 ,
         \21397 , \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 , \21405 , \21406 ,
         \21407 , \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 , \21415 , \21416 ,
         \21417 , \21418 , \21419 , \21420 , \21421 , \21422 , \21423 , \21424 , \21425 , \21426 ,
         \21427 , \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 , \21435 , \21436 ,
         \21437 , \21438 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 , \21445 , \21446 ,
         \21447 , \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 , \21455 , \21456 ,
         \21457 , \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 , \21465 , \21466 ,
         \21467 , \21468 , \21469 , \21470 , \21471 , \21472 , \21473 , \21474 , \21475 , \21476 ,
         \21477 , \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 , \21485 , \21486 ,
         \21487 , \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 , \21495 , \21496 ,
         \21497 , \21498 , \21499 , \21500 , \21501 , \21502 , \21503 , \21504 , \21505 , \21506 ,
         \21507 , \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 , \21515 , \21516 ,
         \21517 , \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 , \21525 , \21526 ,
         \21527 , \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 , \21535 , \21536 ,
         \21537 , \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 , \21545 , \21546 ,
         \21547 , \21548 , \21549 , \21550 , \21551 , \21552 , \21553 , \21554 , \21555 , \21556 ,
         \21557 , \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 , \21565 , \21566 ,
         \21567 , \21568 , \21569 , \21570 , \21571 , \21572 , \21573 , \21574 , \21575 , \21576 ,
         \21577 , \21578 , \21579 , \21580 , \21581 , \21582 , \21583 , \21584 , \21585 , \21586 ,
         \21587 , \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 , \21595 , \21596 ,
         \21597 , \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 , \21605 , \21606 ,
         \21607 , \21608 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 , \21615 , \21616 ,
         \21617 , \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 , \21625 , \21626 ,
         \21627 , \21628 , \21629 , \21630 , \21631 , \21632 , \21633 , \21634 , \21635 , \21636 ,
         \21637 , \21638 , \21639 , \21640 , \21641 , \21642 , \21643 , \21644 , \21645 , \21646 ,
         \21647 , \21648 , \21649 , \21650 , \21651 , \21652 , \21653 , \21654 , \21655 , \21656 ,
         \21657 , \21658 , \21659 , \21660 , \21661 , \21662 , \21663 , \21664 , \21665 , \21666 ,
         \21667 , \21668 , \21669 , \21670 , \21671 , \21672 , \21673 , \21674 , \21675 , \21676 ,
         \21677 , \21678 , \21679 , \21680 , \21681 , \21682 , \21683 , \21684 , \21685 , \21686 ,
         \21687 , \21688 , \21689 , \21690 , \21691 , \21692 , \21693 , \21694 , \21695 , \21696 ,
         \21697 , \21698 , \21699 , \21700 , \21701 , \21702 , \21703 , \21704 , \21705 , \21706 ,
         \21707 , \21708 , \21709 , \21710 , \21711 , \21712 , \21713 , \21714 , \21715 , \21716 ,
         \21717 , \21718 , \21719 , \21720 , \21721 , \21722 , \21723 , \21724 , \21725 , \21726 ,
         \21727 , \21728 , \21729 , \21730 , \21731 , \21732 , \21733 , \21734 , \21735 , \21736 ,
         \21737 , \21738 , \21739 , \21740 , \21741 , \21742 , \21743 , \21744 , \21745 , \21746 ,
         \21747 , \21748 , \21749 , \21750 , \21751 , \21752 , \21753 , \21754 , \21755 , \21756 ,
         \21757 , \21758 , \21759 , \21760 , \21761 , \21762 , \21763 , \21764 , \21765 , \21766 ,
         \21767 , \21768 , \21769 , \21770 , \21771 , \21772 , \21773 , \21774 , \21775 , \21776 ,
         \21777 , \21778 , \21779 , \21780 , \21781 , \21782 , \21783 , \21784 , \21785 , \21786 ,
         \21787 , \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 , \21795 , \21796 ,
         \21797 , \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 , \21805 , \21806 ,
         \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 , \21815 , \21816 ,
         \21817 , \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 , \21825 , \21826 ,
         \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 , \21835 , \21836 ,
         \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 , \21845 , \21846 ,
         \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 , \21855 , \21856 ,
         \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 , \21865 , \21866 ,
         \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 , \21875 , \21876 ,
         \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 , \21885 , \21886 ,
         \21887 , \21888 , \21889 , \21890 , \21891 , \21892 , \21893 , \21894 , \21895 , \21896 ,
         \21897 , \21898 , \21899 , \21900 , \21901 , \21902 , \21903 , \21904 , \21905 , \21906 ,
         \21907 , \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 , \21915 , \21916 ,
         \21917 , \21918 , \21919 , \21920 , \21921 , \21922 , \21923 , \21924 , \21925 , \21926 ,
         \21927 , \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 , \21935 , \21936 ,
         \21937 , \21938 , \21939 , \21940 , \21941 , \21942 , \21943 , \21944 , \21945 , \21946 ,
         \21947 , \21948 , \21949 , \21950 , \21951 , \21952 , \21953 , \21954 , \21955 , \21956 ,
         \21957 , \21958 , \21959 , \21960 , \21961 , \21962 , \21963 , \21964 , \21965 , \21966 ,
         \21967 , \21968 , \21969 , \21970 , \21971 , \21972 , \21973 , \21974 , \21975 , \21976 ,
         \21977 , \21978 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 , \21985 , \21986 ,
         \21987 , \21988 , \21989 , \21990 , \21991 , \21992 , \21993 , \21994 , \21995 , \21996 ,
         \21997 , \21998 , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 , \22005 , \22006 ,
         \22007 , \22008 , \22009 , \22010 , \22011 , \22012 , \22013 , \22014 , \22015 , \22016 ,
         \22017 , \22018 , \22019 , \22020 , \22021 , \22022 , \22023 , \22024 , \22025 , \22026 ,
         \22027 , \22028 , \22029 , \22030 , \22031 , \22032 , \22033 , \22034 , \22035 , \22036 ,
         \22037 , \22038 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 , \22045 , \22046 ,
         \22047 , \22048 , \22049 , \22050 , \22051 , \22052 , \22053 , \22054 , \22055 , \22056 ,
         \22057 , \22058 , \22059 , \22060 , \22061 , \22062 , \22063 , \22064 , \22065 , \22066 ,
         \22067 , \22068 , \22069 , \22070 , \22071 , \22072 , \22073 , \22074 , \22075 , \22076 ,
         \22077 , \22078 , \22079 , \22080 , \22081 , \22082 , \22083 , \22084 , \22085 , \22086 ,
         \22087 , \22088 , \22089 , \22090 , \22091 , \22092 , \22093 , \22094 , \22095 , \22096 ,
         \22097 , \22098 , \22099 , \22100 , \22101 , \22102 , \22103 , \22104 , \22105 , \22106 ,
         \22107 , \22108 , \22109 , \22110 , \22111 , \22112 , \22113 , \22114 , \22115 , \22116 ,
         \22117 , \22118 , \22119 , \22120 , \22121 , \22122 , \22123 , \22124 , \22125 , \22126 ,
         \22127 , \22128 , \22129 , \22130 , \22131 , \22132 , \22133 , \22134 , \22135 , \22136 ,
         \22137 , \22138 , \22139 , \22140 , \22141 , \22142 , \22143 , \22144 , \22145 , \22146 ,
         \22147 , \22148 , \22149 , \22150 , \22151 , \22152 , \22153 , \22154 , \22155 , \22156 ,
         \22157 , \22158 , \22159 , \22160 , \22161 , \22162 , \22163 , \22164 , \22165 , \22166 ,
         \22167 , \22168 , \22169 , \22170 , \22171 , \22172 , \22173 , \22174 , \22175 , \22176 ,
         \22177 , \22178 , \22179 , \22180 , \22181 , \22182 , \22183 , \22184 , \22185 , \22186 ,
         \22187 , \22188 , \22189 , \22190 , \22191 , \22192 , \22193 , \22194 , \22195 , \22196 ,
         \22197 , \22198 , \22199 , \22200 , \22201 , \22202 , \22203 , \22204 , \22205 , \22206 ,
         \22207 , \22208 , \22209 , \22210 , \22211 , \22212 , \22213 , \22214 , \22215 , \22216 ,
         \22217 , \22218 , \22219 , \22220 , \22221 , \22222 , \22223 , \22224 , \22225 , \22226 ,
         \22227 , \22228 , \22229 , \22230 , \22231 , \22232 , \22233 , \22234 , \22235 , \22236 ,
         \22237 , \22238 , \22239 , \22240 , \22241 , \22242 , \22243 , \22244 , \22245 , \22246 ,
         \22247 , \22248 , \22249 , \22250 , \22251 , \22252 , \22253 , \22254 , \22255 , \22256 ,
         \22257 , \22258 , \22259 , \22260 , \22261 , \22262 , \22263 , \22264 , \22265 , \22266 ,
         \22267 , \22268 , \22269 , \22270 , \22271 , \22272 , \22273 , \22274 , \22275 , \22276 ,
         \22277 , \22278 , \22279 , \22280 , \22281 , \22282 , \22283 , \22284 , \22285 , \22286 ,
         \22287 , \22288 , \22289 , \22290 , \22291 , \22292 , \22293 , \22294 , \22295 , \22296 ,
         \22297 , \22298 , \22299 , \22300 , \22301 , \22302 , \22303 , \22304 , \22305 , \22306 ,
         \22307 , \22308 , \22309 , \22310 , \22311 , \22312 , \22313 , \22314 , \22315 , \22316 ,
         \22317 , \22318 , \22319 , \22320 , \22321 , \22322 , \22323 , \22324 , \22325 , \22326 ,
         \22327 , \22328 , \22329 , \22330 , \22331 , \22332 , \22333 , \22334 , \22335 , \22336 ,
         \22337 , \22338 , \22339 , \22340 , \22341 , \22342 , \22343 , \22344 , \22345 , \22346 ,
         \22347 , \22348 , \22349 , \22350 , \22351 , \22352 , \22353 , \22354 , \22355 , \22356 ,
         \22357 , \22358 , \22359 , \22360 , \22361 , \22362 , \22363 , \22364 , \22365 , \22366 ,
         \22367 , \22368 , \22369 , \22370 , \22371 , \22372 , \22373 , \22374 , \22375 , \22376 ,
         \22377 , \22378 , \22379 , \22380 , \22381 , \22382 , \22383 , \22384 , \22385 , \22386 ,
         \22387 , \22388 , \22389 , \22390 , \22391 , \22392 , \22393 , \22394 , \22395 , \22396 ,
         \22397 , \22398 , \22399 , \22400 , \22401 , \22402 , \22403 , \22404 , \22405 , \22406 ,
         \22407 , \22408 , \22409 , \22410 , \22411 , \22412 , \22413 , \22414 , \22415 , \22416 ,
         \22417 , \22418 , \22419 , \22420 , \22421 , \22422 , \22423 , \22424 , \22425 , \22426 ,
         \22427 , \22428 , \22429 , \22430 , \22431 , \22432 , \22433 , \22434 , \22435 , \22436 ,
         \22437 , \22438 , \22439 , \22440 , \22441 , \22442 , \22443 , \22444 , \22445 , \22446 ,
         \22447 , \22448 , \22449 , \22450 , \22451 , \22452 , \22453 , \22454 , \22455 , \22456 ,
         \22457 , \22458 , \22459 , \22460 , \22461 , \22462 , \22463 , \22464 , \22465 , \22466 ,
         \22467 , \22468 , \22469 , \22470 , \22471 , \22472 , \22473 , \22474 , \22475 , \22476 ,
         \22477 , \22478 , \22479 , \22480 , \22481 , \22482 , \22483 , \22484 , \22485 , \22486 ,
         \22487 , \22488 , \22489 , \22490 , \22491 , \22492 , \22493 , \22494 , \22495 , \22496 ,
         \22497 , \22498 , \22499 , \22500 , \22501 , \22502 , \22503 , \22504 , \22505 , \22506 ,
         \22507 , \22508 , \22509 , \22510 , \22511 , \22512 , \22513 , \22514 , \22515 , \22516 ,
         \22517 , \22518 , \22519 , \22520 , \22521 , \22522 , \22523 , \22524 , \22525 , \22526 ,
         \22527 , \22528 , \22529 , \22530 , \22531 , \22532 , \22533 , \22534 , \22535 , \22536 ,
         \22537 , \22538 , \22539 , \22540 , \22541 , \22542 , \22543 , \22544 , \22545 , \22546 ,
         \22547 , \22548 , \22549 , \22550 , \22551 , \22552 , \22553 , \22554 , \22555 , \22556 ,
         \22557 , \22558 , \22559 , \22560 , \22561 , \22562 , \22563 , \22564 , \22565 , \22566 ,
         \22567 , \22568 , \22569 , \22570 , \22571 , \22572 , \22573 , \22574 , \22575 , \22576 ,
         \22577 , \22578 , \22579 , \22580 , \22581 , \22582 , \22583 , \22584 , \22585 , \22586 ,
         \22587 , \22588 , \22589 , \22590 , \22591 , \22592 , \22593 , \22594 , \22595 , \22596 ,
         \22597 , \22598 , \22599 , \22600 , \22601 , \22602 , \22603 , \22604 , \22605 , \22606 ,
         \22607 , \22608 , \22609 , \22610 , \22611 , \22612 , \22613 , \22614 , \22615 , \22616 ,
         \22617 , \22618 , \22619 , \22620 , \22621 , \22622 , \22623 , \22624 , \22625 , \22626 ,
         \22627 , \22628 , \22629 , \22630 , \22631 , \22632 , \22633 , \22634 , \22635 , \22636 ,
         \22637 , \22638 , \22639 , \22640 , \22641 , \22642 , \22643 , \22644 , \22645 , \22646 ,
         \22647 , \22648 , \22649 , \22650 , \22651 , \22652 , \22653 , \22654 , \22655 , \22656 ,
         \22657 , \22658 , \22659 , \22660 , \22661 , \22662 , \22663 , \22664 , \22665 , \22666 ,
         \22667 , \22668 , \22669 , \22670 , \22671 , \22672 , \22673 , \22674 , \22675 , \22676 ,
         \22677 , \22678 , \22679 , \22680 , \22681 , \22682 , \22683 , \22684 , \22685 , \22686 ,
         \22687 , \22688 , \22689 , \22690 , \22691 , \22692 , \22693 , \22694 , \22695 , \22696 ,
         \22697 , \22698 , \22699 , \22700 , \22701 , \22702 , \22703 , \22704 , \22705 , \22706 ,
         \22707 , \22708 , \22709 , \22710 , \22711 , \22712 , \22713 , \22714 , \22715 , \22716 ,
         \22717 , \22718 , \22719 , \22720 , \22721 , \22722 , \22723 , \22724 , \22725 , \22726 ,
         \22727 , \22728 , \22729 , \22730 , \22731 , \22732 , \22733 , \22734 , \22735 , \22736 ,
         \22737 , \22738 , \22739 , \22740 , \22741 , \22742 , \22743 , \22744 , \22745 , \22746 ,
         \22747 , \22748 , \22749 , \22750 , \22751 , \22752 , \22753 , \22754 , \22755 , \22756 ,
         \22757 , \22758 , \22759 , \22760 , \22761 , \22762 , \22763 , \22764 , \22765 , \22766 ,
         \22767 , \22768 , \22769 , \22770 , \22771 , \22772 , \22773 , \22774 , \22775 , \22776 ,
         \22777 , \22778 , \22779 , \22780 , \22781 , \22782 , \22783 , \22784 , \22785 , \22786 ,
         \22787 , \22788 , \22789 , \22790 , \22791 , \22792 , \22793 , \22794 , \22795 , \22796 ,
         \22797 , \22798 , \22799 , \22800 , \22801 , \22802 , \22803 , \22804 , \22805 , \22806 ,
         \22807 , \22808 , \22809 , \22810 , \22811 , \22812 , \22813 , \22814 , \22815 , \22816 ,
         \22817 , \22818 , \22819 , \22820 , \22821 , \22822 , \22823 , \22824 , \22825 , \22826 ,
         \22827 , \22828 , \22829 , \22830 , \22831 , \22832 , \22833 , \22834 , \22835 , \22836 ,
         \22837 , \22838 , \22839 , \22840 , \22841 , \22842 , \22843 , \22844 , \22845 , \22846 ,
         \22847 , \22848 , \22849 , \22850 , \22851 , \22852 , \22853 , \22854 , \22855 , \22856 ,
         \22857 , \22858 , \22859 , \22860 , \22861 , \22862 , \22863 , \22864 , \22865 , \22866 ,
         \22867 , \22868 , \22869 , \22870 , \22871 , \22872 , \22873 , \22874 , \22875 , \22876 ,
         \22877 , \22878 , \22879 , \22880 , \22881 , \22882 , \22883 , \22884 , \22885 , \22886 ,
         \22887 , \22888 , \22889 , \22890 , \22891 , \22892 , \22893 , \22894 , \22895 , \22896 ,
         \22897 , \22898 , \22899 , \22900 , \22901 , \22902 , \22903 , \22904 , \22905 , \22906 ,
         \22907 , \22908 , \22909 , \22910 , \22911 , \22912 , \22913 , \22914 , \22915 , \22916 ,
         \22917 , \22918 , \22919 , \22920 , \22921 , \22922 , \22923 , \22924 , \22925 , \22926 ,
         \22927 , \22928 , \22929 , \22930 , \22931 , \22932 , \22933 , \22934 , \22935 , \22936 ,
         \22937 , \22938 , \22939 , \22940 , \22941 , \22942 , \22943 , \22944 , \22945 , \22946 ,
         \22947 , \22948 , \22949 , \22950 , \22951 , \22952 , \22953 , \22954 , \22955 , \22956 ,
         \22957 , \22958 , \22959 , \22960 , \22961 , \22962 , \22963 , \22964 , \22965 , \22966 ,
         \22967 , \22968 , \22969 , \22970 , \22971 , \22972 , \22973 , \22974 , \22975 , \22976 ,
         \22977 , \22978 , \22979 , \22980 , \22981 , \22982 , \22983 , \22984 , \22985 , \22986 ,
         \22987 , \22988 , \22989 , \22990 , \22991 , \22992 , \22993 , \22994 , \22995 , \22996 ,
         \22997 , \22998 , \22999 , \23000 , \23001 , \23002 , \23003 , \23004 , \23005 , \23006 ,
         \23007 , \23008 , \23009 , \23010 , \23011 , \23012 , \23013 , \23014 , \23015 , \23016 ,
         \23017 , \23018 , \23019 , \23020 , \23021 , \23022 , \23023 , \23024 , \23025 , \23026 ,
         \23027 , \23028 , \23029 , \23030 , \23031 , \23032 , \23033 , \23034 , \23035 , \23036 ,
         \23037 , \23038 , \23039 , \23040 , \23041 , \23042 , \23043 , \23044 , \23045 , \23046 ,
         \23047 , \23048 , \23049 , \23050 , \23051 , \23052 , \23053 , \23054 , \23055 , \23056 ,
         \23057 , \23058 , \23059 , \23060 , \23061 , \23062 , \23063 , \23064 , \23065 , \23066 ,
         \23067 , \23068 , \23069 , \23070 , \23071 , \23072 , \23073 , \23074 , \23075 , \23076 ,
         \23077 , \23078 , \23079 , \23080 , \23081 , \23082 , \23083 , \23084 , \23085 , \23086 ,
         \23087 , \23088 , \23089 , \23090 , \23091 , \23092 , \23093 , \23094 , \23095 , \23096 ,
         \23097 , \23098 , \23099 , \23100 , \23101 , \23102 , \23103 , \23104 , \23105 , \23106 ,
         \23107 , \23108 , \23109 , \23110 , \23111 , \23112 , \23113 , \23114 , \23115 , \23116 ,
         \23117 , \23118 , \23119 , \23120 , \23121 , \23122 , \23123 , \23124 , \23125 , \23126 ,
         \23127 , \23128 , \23129 , \23130 , \23131 , \23132 , \23133 , \23134 , \23135 , \23136 ,
         \23137 , \23138 , \23139 , \23140 , \23141 , \23142 , \23143 , \23144 , \23145 , \23146 ,
         \23147 , \23148 , \23149 , \23150 , \23151 , \23152 , \23153 , \23154 , \23155 , \23156 ,
         \23157 , \23158 , \23159 , \23160 , \23161 , \23162 , \23163 , \23164 , \23165 , \23166 ,
         \23167 , \23168 , \23169 , \23170 , \23171 , \23172 , \23173 , \23174 , \23175 , \23176 ,
         \23177 , \23178 , \23179 , \23180 , \23181 , \23182 , \23183 , \23184 , \23185 , \23186 ,
         \23187 , \23188 , \23189 , \23190 , \23191 , \23192 , \23193 , \23194 , \23195 , \23196 ,
         \23197 , \23198 , \23199 , \23200 , \23201 , \23202 , \23203 , \23204 , \23205 , \23206 ,
         \23207 , \23208 , \23209 , \23210 , \23211 , \23212 , \23213 , \23214 , \23215 , \23216 ,
         \23217 , \23218 , \23219 , \23220 , \23221 , \23222 , \23223 , \23224 , \23225 , \23226 ,
         \23227 , \23228 , \23229 , \23230 , \23231 , \23232 , \23233 , \23234 , \23235 , \23236 ,
         \23237 , \23238 , \23239 , \23240 , \23241 , \23242 , \23243 , \23244 , \23245 , \23246 ,
         \23247 , \23248 , \23249 , \23250 , \23251 , \23252 , \23253 , \23254 , \23255 , \23256 ,
         \23257 , \23258 , \23259 , \23260 , \23261 , \23262 , \23263 , \23264 , \23265 , \23266 ,
         \23267 , \23268 , \23269 , \23270 , \23271 , \23272 , \23273 , \23274 , \23275 , \23276 ,
         \23277 , \23278 , \23279 , \23280 , \23281 , \23282 , \23283 , \23284 , \23285 , \23286 ,
         \23287 , \23288 , \23289 , \23290 , \23291 , \23292 , \23293 , \23294 , \23295 , \23296 ,
         \23297 , \23298 , \23299 , \23300 , \23301 , \23302 , \23303 , \23304 , \23305 , \23306 ,
         \23307 , \23308 , \23309 , \23310 , \23311 , \23312 , \23313 , \23314 , \23315 , \23316 ,
         \23317 , \23318 , \23319 , \23320 , \23321 , \23322 , \23323 , \23324 , \23325 , \23326 ,
         \23327 , \23328 , \23329 , \23330 , \23331 , \23332 , \23333 , \23334 , \23335 , \23336 ,
         \23337 , \23338 , \23339 , \23340 , \23341 , \23342 , \23343 , \23344 , \23345 , \23346 ,
         \23347 , \23348 , \23349 , \23350 , \23351 , \23352 , \23353 , \23354 , \23355 , \23356 ,
         \23357 , \23358 , \23359 , \23360 , \23361 , \23362 , \23363 , \23364 , \23365 , \23366 ,
         \23367 , \23368 , \23369 , \23370 , \23371 , \23372 , \23373 , \23374 , \23375 , \23376 ,
         \23377 , \23378 , \23379 , \23380 , \23381 , \23382 , \23383 , \23384 , \23385 , \23386 ,
         \23387 , \23388 , \23389 , \23390 , \23391 , \23392 , \23393 , \23394 , \23395 , \23396 ,
         \23397 , \23398 , \23399 , \23400 , \23401 , \23402 , \23403 , \23404 , \23405 , \23406 ,
         \23407 , \23408 , \23409 , \23410 , \23411 , \23412 , \23413 , \23414 , \23415 , \23416 ,
         \23417 , \23418 , \23419 , \23420 , \23421 , \23422 , \23423 , \23424 , \23425 , \23426 ,
         \23427 , \23428 , \23429 , \23430 , \23431 , \23432 , \23433 , \23434 , \23435 , \23436 ,
         \23437 , \23438 , \23439 , \23440 , \23441 , \23442 , \23443 , \23444 , \23445 , \23446 ,
         \23447 , \23448 , \23449 , \23450 , \23451 , \23452 , \23453 , \23454 , \23455 , \23456 ,
         \23457 , \23458 , \23459 , \23460 , \23461 , \23462 , \23463 , \23464 , \23465 , \23466 ,
         \23467 , \23468 , \23469 , \23470 , \23471 , \23472 , \23473 , \23474 , \23475 , \23476 ,
         \23477 , \23478 , \23479 , \23480 , \23481 , \23482 , \23483 , \23484 , \23485 , \23486 ,
         \23487 , \23488 , \23489 , \23490 , \23491 , \23492 , \23493 , \23494 , \23495 , \23496 ,
         \23497 , \23498 , \23499 , \23500 , \23501 , \23502 , \23503 , \23504 , \23505 , \23506 ,
         \23507 , \23508 , \23509 , \23510 , \23511 , \23512 , \23513 , \23514 , \23515 , \23516 ,
         \23517 , \23518 , \23519 , \23520 , \23521 , \23522 , \23523 , \23524 , \23525 , \23526 ,
         \23527 , \23528 , \23529 , \23530 , \23531 , \23532 , \23533 , \23534 , \23535 , \23536 ,
         \23537 , \23538 , \23539 , \23540 , \23541 , \23542 , \23543 , \23544 , \23545 , \23546 ,
         \23547 , \23548 , \23549 , \23550 , \23551 , \23552 , \23553 , \23554 , \23555 , \23556 ,
         \23557 , \23558 , \23559 , \23560 , \23561 , \23562 , \23563 , \23564 , \23565 , \23566 ,
         \23567 , \23568 , \23569 , \23570 , \23571 , \23572 , \23573 , \23574 , \23575 , \23576 ,
         \23577 , \23578 , \23579 , \23580 , \23581 , \23582 , \23583 , \23584 , \23585 , \23586 ,
         \23587 , \23588 , \23589 , \23590 , \23591 , \23592 , \23593 , \23594 , \23595 , \23596 ,
         \23597 , \23598 , \23599 , \23600 , \23601 , \23602 , \23603 , \23604 , \23605 , \23606 ,
         \23607 , \23608 , \23609 , \23610 , \23611 , \23612 , \23613 , \23614 , \23615 , \23616 ,
         \23617 , \23618 , \23619 , \23620 , \23621 , \23622 , \23623 , \23624 , \23625 , \23626 ,
         \23627 , \23628 , \23629 , \23630 , \23631 , \23632 , \23633 , \23634 , \23635 , \23636 ,
         \23637 , \23638 , \23639 , \23640 , \23641 , \23642 , \23643 , \23644 , \23645 , \23646 ,
         \23647 , \23648 , \23649 , \23650 , \23651 , \23652 , \23653 , \23654 , \23655 , \23656 ,
         \23657 , \23658 , \23659 , \23660 , \23661 , \23662 , \23663 , \23664 , \23665 , \23666 ,
         \23667 , \23668 , \23669 , \23670 , \23671 , \23672 , \23673 , \23674 , \23675 , \23676 ,
         \23677 , \23678 , \23679 , \23680 , \23681 , \23682 , \23683 , \23684 , \23685 , \23686 ,
         \23687 , \23688 , \23689 , \23690 , \23691 , \23692 , \23693 , \23694 , \23695 , \23696 ,
         \23697 , \23698 , \23699 , \23700 , \23701 , \23702 , \23703 , \23704 , \23705 , \23706 ,
         \23707 , \23708 , \23709 , \23710 , \23711 , \23712 , \23713 , \23714 , \23715 , \23716 ,
         \23717 , \23718 , \23719 , \23720 , \23721 , \23722 , \23723 , \23724 , \23725 , \23726 ,
         \23727 , \23728 , \23729 , \23730 , \23731 , \23732 , \23733 , \23734 , \23735 , \23736 ,
         \23737 , \23738 , \23739 , \23740 , \23741 , \23742 , \23743 , \23744 , \23745 , \23746 ,
         \23747 , \23748 , \23749 , \23750 , \23751 , \23752 , \23753 , \23754 , \23755 , \23756 ,
         \23757 , \23758 , \23759 , \23760 , \23761 , \23762 , \23763 , \23764 , \23765 , \23766 ,
         \23767 , \23768 , \23769 , \23770 , \23771 , \23772 , \23773 , \23774 , \23775 , \23776 ,
         \23777 , \23778 , \23779 , \23780 , \23781 , \23782 , \23783 , \23784 , \23785 , \23786 ,
         \23787 , \23788 , \23789 , \23790 , \23791 , \23792 , \23793 , \23794 , \23795 , \23796 ,
         \23797 , \23798 , \23799 , \23800 , \23801 , \23802 , \23803 , \23804 , \23805 , \23806 ,
         \23807 , \23808 , \23809 , \23810 , \23811 , \23812 , \23813 , \23814 , \23815 , \23816 ,
         \23817 , \23818 , \23819 , \23820 , \23821 , \23822 , \23823 , \23824 , \23825 , \23826 ,
         \23827 , \23828 , \23829 , \23830 , \23831 , \23832 , \23833 , \23834 , \23835 , \23836 ,
         \23837 , \23838 , \23839 , \23840 , \23841 , \23842 , \23843 , \23844 , \23845 , \23846 ,
         \23847 , \23848 , \23849 , \23850 , \23851 , \23852 , \23853 , \23854 , \23855 , \23856 ,
         \23857 , \23858 , \23859 , \23860 , \23861 , \23862 , \23863 , \23864 , \23865 , \23866 ,
         \23867 , \23868 , \23869 , \23870 , \23871 , \23872 , \23873 , \23874 , \23875 , \23876 ,
         \23877 , \23878 , \23879 , \23880 , \23881 , \23882 , \23883 , \23884 , \23885 , \23886 ,
         \23887 , \23888 , \23889 , \23890 , \23891 , \23892 , \23893 , \23894 , \23895 , \23896 ,
         \23897 , \23898 , \23899 , \23900 , \23901 , \23902 , \23903 , \23904 , \23905 , \23906 ,
         \23907 , \23908 , \23909 , \23910 , \23911 , \23912 , \23913 , \23914 , \23915 , \23916 ,
         \23917 , \23918 , \23919 , \23920 , \23921 , \23922 , \23923 , \23924 , \23925 , \23926 ,
         \23927 , \23928 , \23929 , \23930 , \23931 , \23932 , \23933 , \23934 , \23935 , \23936 ,
         \23937 , \23938 , \23939 , \23940 , \23941 , \23942 , \23943 , \23944 , \23945 , \23946 ,
         \23947 , \23948 , \23949 , \23950 , \23951 , \23952 , \23953 , \23954 , \23955 , \23956 ,
         \23957 , \23958 , \23959 , \23960 , \23961 , \23962 , \23963 , \23964 , \23965 , \23966 ,
         \23967 , \23968 , \23969 , \23970 , \23971 , \23972 , \23973 , \23974 , \23975 , \23976 ,
         \23977 , \23978 , \23979 , \23980 , \23981 , \23982 , \23983 , \23984 , \23985 , \23986 ,
         \23987 , \23988 , \23989 , \23990 , \23991 , \23992 , \23993 , \23994 , \23995 , \23996 ,
         \23997 , \23998 , \23999 , \24000 , \24001 , \24002 , \24003 , \24004 , \24005 , \24006 ,
         \24007 , \24008 , \24009 , \24010 , \24011 , \24012 , \24013 , \24014 , \24015 , \24016 ,
         \24017 , \24018 , \24019 , \24020 , \24021 , \24022 , \24023 , \24024 , \24025 , \24026 ,
         \24027 , \24028 , \24029 , \24030 , \24031 , \24032 , \24033 , \24034 , \24035 , \24036 ,
         \24037 , \24038 , \24039 , \24040 , \24041 , \24042 , \24043 , \24044 , \24045 , \24046 ,
         \24047 , \24048 , \24049 , \24050 , \24051 , \24052 , \24053 , \24054 , \24055 , \24056 ,
         \24057 , \24058 , \24059 , \24060 , \24061 , \24062 , \24063 , \24064 , \24065 , \24066 ,
         \24067 , \24068 , \24069 , \24070 , \24071 , \24072 , \24073 , \24074 , \24075 , \24076 ,
         \24077 , \24078 , \24079 , \24080 , \24081 , \24082 , \24083 , \24084 , \24085 , \24086 ,
         \24087 , \24088 , \24089 , \24090 , \24091 , \24092 , \24093 , \24094 , \24095 , \24096 ,
         \24097 , \24098 , \24099 , \24100 , \24101 , \24102 , \24103 , \24104 , \24105 , \24106 ,
         \24107 , \24108 , \24109 , \24110 , \24111 , \24112 , \24113 , \24114 , \24115 , \24116 ,
         \24117 , \24118 , \24119 , \24120 , \24121 , \24122 , \24123 , \24124 , \24125 , \24126 ,
         \24127 , \24128 , \24129 , \24130 , \24131 , \24132 , \24133 , \24134 , \24135 , \24136 ,
         \24137 , \24138 , \24139 , \24140 , \24141 , \24142 , \24143 , \24144 , \24145 , \24146 ,
         \24147 , \24148 , \24149 , \24150 , \24151 , \24152 , \24153 , \24154 , \24155 , \24156 ,
         \24157 , \24158 , \24159 , \24160 , \24161 , \24162 , \24163 , \24164 , \24165 , \24166 ,
         \24167 , \24168 , \24169 , \24170 , \24171 , \24172 , \24173 , \24174 , \24175 , \24176 ,
         \24177 , \24178 , \24179 , \24180 , \24181 , \24182 , \24183 , \24184 , \24185 , \24186 ,
         \24187 , \24188 , \24189 , \24190 , \24191 , \24192 , \24193 , \24194 , \24195 , \24196 ,
         \24197 , \24198 , \24199 , \24200 , \24201 , \24202 , \24203 , \24204 , \24205 , \24206 ,
         \24207 , \24208 , \24209 , \24210 , \24211 , \24212 , \24213 , \24214 , \24215 , \24216 ,
         \24217 , \24218 , \24219 , \24220 , \24221 , \24222 , \24223 , \24224 , \24225 , \24226 ,
         \24227 , \24228 , \24229 , \24230 , \24231 , \24232 , \24233 , \24234 , \24235 , \24236 ,
         \24237 , \24238 , \24239 , \24240 , \24241 , \24242 , \24243 , \24244 , \24245 , \24246 ,
         \24247 , \24248 , \24249 , \24250 , \24251 , \24252 , \24253 , \24254 , \24255 , \24256 ,
         \24257 , \24258 , \24259 , \24260 , \24261 , \24262 , \24263 , \24264 , \24265 , \24266 ,
         \24267 , \24268 , \24269 , \24270 , \24271 , \24272 , \24273 , \24274 , \24275 , \24276 ,
         \24277 , \24278 , \24279 , \24280 , \24281 , \24282 , \24283 , \24284 , \24285 , \24286 ,
         \24287 , \24288 , \24289 , \24290 , \24291 , \24292 , \24293 , \24294 , \24295 , \24296 ,
         \24297 , \24298 , \24299 , \24300 , \24301 , \24302 , \24303 , \24304 , \24305 , \24306 ,
         \24307 , \24308 , \24309 , \24310 , \24311 , \24312 , \24313 , \24314 , \24315 , \24316 ,
         \24317 , \24318 , \24319 , \24320 , \24321 , \24322 , \24323 , \24324 , \24325 , \24326 ,
         \24327 , \24328 , \24329 , \24330 , \24331 , \24332 , \24333 , \24334 , \24335 , \24336 ,
         \24337 , \24338 , \24339 , \24340 , \24341 , \24342 , \24343 , \24344 , \24345 , \24346 ,
         \24347 , \24348 , \24349 , \24350 , \24351 , \24352 , \24353 , \24354 , \24355 , \24356 ,
         \24357 , \24358 , \24359 , \24360 , \24361 , \24362 , \24363 , \24364 , \24365 , \24366 ,
         \24367 , \24368 , \24369 , \24370 , \24371 , \24372 , \24373 , \24374 , \24375 , \24376 ,
         \24377 , \24378 , \24379 , \24380 , \24381 , \24382 , \24383 , \24384 , \24385 , \24386 ,
         \24387 , \24388 , \24389 , \24390 , \24391 , \24392 , \24393 , \24394 , \24395 , \24396 ,
         \24397 , \24398 , \24399 , \24400 , \24401 , \24402 , \24403 , \24404 , \24405 , \24406 ,
         \24407 , \24408 , \24409 , \24410 , \24411 , \24412 , \24413 , \24414 , \24415 , \24416 ,
         \24417 , \24418 , \24419 , \24420 , \24421 , \24422 , \24423 , \24424 , \24425 , \24426 ,
         \24427 , \24428 , \24429 , \24430 , \24431 , \24432 , \24433 , \24434 , \24435 , \24436 ,
         \24437 , \24438 , \24439 , \24440 , \24441 , \24442 , \24443 , \24444 , \24445 , \24446 ,
         \24447 , \24448 , \24449 , \24450 , \24451 , \24452 , \24453 , \24454 , \24455 , \24456 ,
         \24457 , \24458 , \24459 , \24460 , \24461 , \24462 , \24463 , \24464 , \24465 , \24466 ,
         \24467 , \24468 , \24469 , \24470 , \24471 , \24472 , \24473 , \24474 , \24475 , \24476 ,
         \24477 , \24478 , \24479 , \24480 , \24481 , \24482 , \24483 , \24484 , \24485 , \24486 ,
         \24487 , \24488 , \24489 , \24490 , \24491 , \24492 , \24493 , \24494 , \24495 , \24496 ,
         \24497 , \24498 , \24499 , \24500 , \24501 , \24502 , \24503 , \24504 , \24505 , \24506 ,
         \24507 , \24508 , \24509 , \24510 , \24511 , \24512 , \24513 , \24514 , \24515 , \24516 ,
         \24517 , \24518 , \24519 , \24520 , \24521 , \24522 , \24523 , \24524 , \24525 , \24526 ,
         \24527 , \24528 , \24529 , \24530 , \24531 , \24532 , \24533 , \24534 , \24535 , \24536 ,
         \24537 , \24538 , \24539 , \24540 , \24541 , \24542 , \24543 , \24544 , \24545 , \24546 ,
         \24547 , \24548 , \24549 , \24550 , \24551 , \24552 , \24553 , \24554 , \24555 , \24556 ,
         \24557 , \24558 , \24559 , \24560 , \24561 , \24562 , \24563 , \24564 , \24565 , \24566 ,
         \24567 , \24568 , \24569 , \24570 , \24571 , \24572 , \24573 , \24574 , \24575 , \24576 ,
         \24577 , \24578 , \24579 , \24580 , \24581 , \24582 , \24583 , \24584 , \24585 , \24586 ,
         \24587 , \24588 , \24589 , \24590 , \24591 , \24592 , \24593 , \24594 , \24595 , \24596 ,
         \24597 , \24598 , \24599 , \24600 , \24601 , \24602 , \24603 , \24604 , \24605 , \24606 ,
         \24607 , \24608 , \24609 , \24610 , \24611 , \24612 , \24613 , \24614 , \24615 , \24616 ,
         \24617 , \24618 , \24619 , \24620 , \24621 , \24622 , \24623 , \24624 , \24625 , \24626 ,
         \24627 , \24628 , \24629 , \24630 , \24631 , \24632 , \24633 , \24634 , \24635 , \24636 ,
         \24637 , \24638 , \24639 , \24640 , \24641 , \24642 , \24643 , \24644 , \24645 , \24646 ,
         \24647 , \24648 , \24649 , \24650 , \24651 , \24652 , \24653 , \24654 , \24655 , \24656 ,
         \24657 , \24658 , \24659 , \24660 , \24661 , \24662 , \24663 , \24664 , \24665 , \24666 ,
         \24667 , \24668 , \24669 , \24670 , \24671 , \24672 , \24673 , \24674 , \24675 , \24676 ,
         \24677 , \24678 , \24679 , \24680 , \24681 , \24682 , \24683 , \24684 , \24685 , \24686 ,
         \24687 , \24688 , \24689 , \24690 , \24691 , \24692 , \24693 , \24694 , \24695 , \24696 ,
         \24697 , \24698 , \24699 , \24700 , \24701 , \24702 , \24703 , \24704 , \24705 , \24706 ,
         \24707 , \24708 , \24709 , \24710 , \24711 , \24712 , \24713 , \24714 , \24715 , \24716 ,
         \24717 , \24718 , \24719 , \24720 , \24721 , \24722 , \24723 , \24724 , \24725 , \24726 ,
         \24727 , \24728 , \24729 , \24730 , \24731 , \24732 , \24733 , \24734 , \24735 , \24736 ,
         \24737 , \24738 , \24739 , \24740 , \24741 , \24742 , \24743 , \24744 , \24745 , \24746 ,
         \24747 , \24748 , \24749 , \24750 , \24751 , \24752 , \24753 , \24754 , \24755 , \24756 ,
         \24757 , \24758 , \24759 , \24760 , \24761 , \24762 , \24763 , \24764 , \24765 , \24766 ,
         \24767 , \24768 , \24769 , \24770 , \24771 , \24772 , \24773 , \24774 , \24775 , \24776 ,
         \24777 , \24778 , \24779 , \24780 , \24781 , \24782 , \24783 , \24784 , \24785 , \24786 ,
         \24787 , \24788 , \24789 , \24790 , \24791 , \24792 , \24793 , \24794 , \24795 , \24796 ,
         \24797 , \24798 , \24799 , \24800 , \24801 , \24802 , \24803 , \24804 , \24805 , \24806 ,
         \24807 , \24808 , \24809 , \24810 , \24811 , \24812 , \24813 , \24814 , \24815 , \24816 ,
         \24817 , \24818 , \24819 , \24820 , \24821 , \24822 , \24823 , \24824 , \24825 , \24826 ,
         \24827 , \24828 , \24829 , \24830 , \24831 , \24832 , \24833 , \24834 , \24835 , \24836 ,
         \24837 , \24838 , \24839 , \24840 , \24841 , \24842 , \24843 , \24844 , \24845 , \24846 ,
         \24847 , \24848 , \24849 , \24850 , \24851 , \24852 , \24853 , \24854 , \24855 , \24856 ,
         \24857 , \24858 , \24859 , \24860 , \24861 , \24862 , \24863 , \24864 , \24865 , \24866 ,
         \24867 , \24868 , \24869 , \24870 , \24871 , \24872 , \24873 , \24874 , \24875 , \24876 ,
         \24877 , \24878 , \24879 , \24880 , \24881 , \24882 , \24883 , \24884 , \24885 , \24886 ,
         \24887 , \24888 , \24889 , \24890 , \24891 , \24892 , \24893 , \24894 , \24895 , \24896 ,
         \24897 , \24898 , \24899 , \24900 , \24901 , \24902 , \24903 , \24904 , \24905 , \24906 ,
         \24907 , \24908 , \24909 , \24910 , \24911 , \24912 , \24913 , \24914 , \24915 , \24916 ,
         \24917 , \24918 , \24919 , \24920 , \24921 , \24922 , \24923 , \24924 , \24925 , \24926 ,
         \24927 , \24928 , \24929 , \24930 , \24931 , \24932 , \24933 , \24934 , \24935 , \24936 ,
         \24937 , \24938 , \24939 , \24940 , \24941 , \24942 , \24943 , \24944 , \24945 , \24946 ,
         \24947 , \24948 , \24949 , \24950 , \24951 , \24952 , \24953 , \24954 , \24955 , \24956 ,
         \24957 , \24958 , \24959 , \24960 , \24961 , \24962 , \24963 , \24964 , \24965 , \24966 ,
         \24967 , \24968 , \24969 , \24970 , \24971 , \24972 , \24973 , \24974 , \24975 , \24976 ,
         \24977 , \24978 , \24979 , \24980 , \24981 , \24982 , \24983 , \24984 , \24985 , \24986 ,
         \24987 , \24988 , \24989 , \24990 , \24991 , \24992 , \24993 , \24994 , \24995 , \24996 ,
         \24997 , \24998 , \24999 , \25000 , \25001 , \25002 , \25003 , \25004 , \25005 , \25006 ,
         \25007 , \25008 , \25009 , \25010 , \25011 , \25012 , \25013 , \25014 , \25015 , \25016 ,
         \25017 , \25018 , \25019 , \25020 , \25021 , \25022 , \25023 , \25024 , \25025 , \25026 ,
         \25027 , \25028 , \25029 , \25030 , \25031 , \25032 , \25033 , \25034 , \25035 , \25036 ,
         \25037 , \25038 , \25039 , \25040 , \25041 , \25042 , \25043 , \25044 , \25045 , \25046 ,
         \25047 , \25048 , \25049 , \25050 , \25051 , \25052 , \25053 , \25054 , \25055 , \25056 ,
         \25057 , \25058 , \25059 , \25060 , \25061 , \25062 , \25063 , \25064 , \25065 , \25066 ,
         \25067 , \25068 , \25069 , \25070 , \25071 , \25072 , \25073 , \25074 , \25075 , \25076 ,
         \25077 , \25078 , \25079 , \25080 , \25081 , \25082 , \25083 , \25084 , \25085 , \25086 ,
         \25087 , \25088 , \25089 , \25090 , \25091 , \25092 , \25093 , \25094 , \25095 , \25096 ,
         \25097 , \25098 , \25099 , \25100 , \25101 , \25102 , \25103 , \25104 , \25105 , \25106 ,
         \25107 , \25108 , \25109 , \25110 , \25111 , \25112 , \25113 , \25114 , \25115 , \25116 ,
         \25117 , \25118 , \25119 , \25120 , \25121 , \25122 , \25123 , \25124 , \25125 , \25126 ,
         \25127 , \25128 , \25129 , \25130 , \25131 , \25132 , \25133 , \25134 , \25135 , \25136 ,
         \25137 , \25138 , \25139 , \25140 , \25141 , \25142 , \25143 , \25144 , \25145 , \25146 ,
         \25147 , \25148 , \25149 , \25150 , \25151 , \25152 , \25153 , \25154 , \25155 , \25156 ,
         \25157 , \25158 , \25159 , \25160 , \25161 , \25162 , \25163 , \25164 , \25165 , \25166 ,
         \25167 , \25168 , \25169 , \25170 , \25171 , \25172 , \25173 , \25174 , \25175 , \25176 ,
         \25177 , \25178 , \25179 , \25180 , \25181 , \25182 , \25183 , \25184 , \25185 , \25186 ,
         \25187 , \25188 , \25189 , \25190 , \25191 , \25192 , \25193 , \25194 , \25195 , \25196 ,
         \25197 , \25198 , \25199 , \25200 , \25201 , \25202 , \25203 , \25204 , \25205 , \25206 ,
         \25207 , \25208 , \25209 , \25210 , \25211 , \25212 , \25213 , \25214 , \25215 , \25216 ,
         \25217 , \25218 , \25219 , \25220 , \25221 , \25222 , \25223 , \25224 , \25225 , \25226 ,
         \25227 , \25228 , \25229 , \25230 , \25231 , \25232 , \25233 , \25234 , \25235 , \25236 ,
         \25237 , \25238 , \25239 , \25240 , \25241 , \25242 , \25243 , \25244 , \25245 , \25246 ,
         \25247 , \25248 , \25249 , \25250 , \25251 , \25252 , \25253 , \25254 , \25255 , \25256 ,
         \25257 , \25258 , \25259 , \25260 , \25261 , \25262 , \25263 , \25264 , \25265 , \25266 ,
         \25267 , \25268 , \25269 , \25270 , \25271 , \25272 , \25273 , \25274 , \25275 , \25276 ,
         \25277 , \25278 , \25279 , \25280 , \25281 , \25282 , \25283 , \25284 , \25285 , \25286 ,
         \25287 , \25288 , \25289 , \25290 , \25291 , \25292 , \25293 , \25294 , \25295 , \25296 ,
         \25297 , \25298 , \25299 , \25300 , \25301 , \25302 , \25303 , \25304 , \25305 , \25306 ,
         \25307 , \25308 , \25309 , \25310 , \25311 , \25312 , \25313 , \25314 , \25315 , \25316 ,
         \25317 , \25318 , \25319 , \25320 , \25321 , \25322 , \25323 , \25324 , \25325 , \25326 ,
         \25327 , \25328 , \25329 , \25330 , \25331 , \25332 , \25333 , \25334 , \25335 , \25336 ,
         \25337 , \25338 , \25339 , \25340 , \25341 , \25342 , \25343 , \25344 , \25345 , \25346 ,
         \25347 , \25348 , \25349 , \25350 , \25351 , \25352 , \25353 , \25354 , \25355 , \25356 ,
         \25357 , \25358 , \25359 , \25360 , \25361 , \25362 , \25363 , \25364 , \25365 , \25366 ,
         \25367 , \25368 , \25369 , \25370 , \25371 , \25372 , \25373 , \25374 , \25375 , \25376 ,
         \25377 , \25378 , \25379 , \25380 , \25381 , \25382 , \25383 , \25384 , \25385 , \25386 ,
         \25387 , \25388 , \25389 , \25390 , \25391 , \25392 , \25393 , \25394 , \25395 , \25396 ,
         \25397 , \25398 , \25399 , \25400 , \25401 , \25402 , \25403 , \25404 , \25405 , \25406 ,
         \25407 , \25408 , \25409 , \25410 , \25411 , \25412 , \25413 , \25414 , \25415 , \25416 ,
         \25417 , \25418 , \25419 , \25420 , \25421 , \25422 , \25423 , \25424 , \25425 , \25426 ,
         \25427 , \25428 , \25429 , \25430 , \25431 , \25432 , \25433 , \25434 , \25435 , \25436 ,
         \25437 , \25438 , \25439 , \25440 , \25441 , \25442 , \25443 , \25444 , \25445 , \25446 ,
         \25447 , \25448 , \25449 , \25450 , \25451 , \25452 , \25453 , \25454 , \25455 , \25456 ,
         \25457 , \25458 , \25459 , \25460 , \25461 , \25462 , \25463 , \25464 , \25465 , \25466 ,
         \25467 , \25468 , \25469 , \25470 , \25471 , \25472 , \25473 , \25474 , \25475 , \25476 ,
         \25477 , \25478 , \25479 , \25480 , \25481 , \25482 , \25483 , \25484 , \25485 , \25486 ,
         \25487 , \25488 , \25489 , \25490 , \25491 , \25492 , \25493 , \25494 , \25495 , \25496 ,
         \25497 , \25498 , \25499 , \25500 , \25501 , \25502 , \25503 , \25504 , \25505 , \25506 ,
         \25507 , \25508 , \25509 , \25510 , \25511 , \25512 , \25513 , \25514 , \25515 , \25516 ,
         \25517 , \25518 , \25519 , \25520 , \25521 , \25522 , \25523 , \25524 , \25525 , \25526 ,
         \25527 , \25528 , \25529 , \25530 , \25531 , \25532 , \25533 , \25534 , \25535 , \25536 ,
         \25537 , \25538 , \25539 , \25540 , \25541 , \25542 , \25543 , \25544 , \25545 , \25546 ,
         \25547 , \25548 , \25549 , \25550 , \25551 , \25552 , \25553 , \25554 , \25555 , \25556 ,
         \25557 , \25558 , \25559 , \25560 , \25561 , \25562 , \25563 , \25564 , \25565 , \25566 ,
         \25567 , \25568 , \25569 , \25570 , \25571 , \25572 , \25573 , \25574 , \25575 , \25576 ,
         \25577 , \25578 , \25579 , \25580 , \25581 , \25582 , \25583 , \25584 , \25585 , \25586 ,
         \25587 , \25588 , \25589 , \25590 , \25591 , \25592 , \25593 , \25594 , \25595 , \25596 ,
         \25597 , \25598 , \25599 , \25600 , \25601 , \25602 , \25603 , \25604 , \25605 , \25606 ,
         \25607 , \25608 , \25609 , \25610 , \25611 , \25612 , \25613 , \25614 , \25615 , \25616 ,
         \25617 , \25618 , \25619 , \25620 , \25621 , \25622 , \25623 , \25624 , \25625 , \25626 ,
         \25627 , \25628 , \25629 , \25630 , \25631 , \25632 , \25633 , \25634 , \25635 , \25636 ,
         \25637 , \25638 , \25639 , \25640 , \25641 , \25642 , \25643 , \25644 , \25645 , \25646 ,
         \25647 , \25648 , \25649 , \25650 , \25651 , \25652 , \25653 , \25654 , \25655 , \25656 ,
         \25657 , \25658 , \25659 , \25660 , \25661 , \25662 , \25663 , \25664 , \25665 , \25666 ,
         \25667 , \25668 , \25669 , \25670 , \25671 , \25672 , \25673 , \25674 , \25675 , \25676 ,
         \25677 , \25678 , \25679 , \25680 , \25681 , \25682 , \25683 , \25684 , \25685 , \25686 ,
         \25687 , \25688 , \25689 , \25690 , \25691 , \25692 , \25693 , \25694 , \25695 , \25696 ,
         \25697 , \25698 , \25699 , \25700 , \25701 , \25702 , \25703 , \25704 , \25705 , \25706 ,
         \25707 , \25708 , \25709 , \25710 , \25711 , \25712 , \25713 , \25714 , \25715 , \25716 ,
         \25717 , \25718 , \25719 , \25720 , \25721 , \25722 , \25723 , \25724 , \25725 , \25726 ,
         \25727 , \25728 , \25729 , \25730 , \25731 , \25732 , \25733 , \25734 , \25735 , \25736 ,
         \25737 , \25738 , \25739 , \25740 , \25741 , \25742 , \25743 , \25744 , \25745 , \25746 ,
         \25747 , \25748 , \25749 , \25750 , \25751 , \25752 , \25753 , \25754 , \25755 , \25756 ,
         \25757 , \25758 , \25759 , \25760 , \25761 , \25762 , \25763 , \25764 , \25765 , \25766 ,
         \25767 , \25768 , \25769 , \25770 , \25771 , \25772 , \25773 , \25774 , \25775 , \25776 ,
         \25777 , \25778 , \25779 , \25780 , \25781 , \25782 , \25783 , \25784 , \25785 , \25786 ,
         \25787 , \25788 , \25789 , \25790 , \25791 , \25792 , \25793 , \25794 , \25795 , \25796 ,
         \25797 , \25798 , \25799 , \25800 , \25801 , \25802 , \25803 , \25804 , \25805 , \25806 ,
         \25807 , \25808 , \25809 , \25810 , \25811 , \25812 , \25813 , \25814 , \25815 , \25816 ,
         \25817 , \25818 , \25819 , \25820 , \25821 , \25822 , \25823 , \25824 , \25825 , \25826 ,
         \25827 , \25828 , \25829 , \25830 , \25831 , \25832 , \25833 , \25834 , \25835 , \25836 ,
         \25837 , \25838 , \25839 , \25840 , \25841 , \25842 , \25843 , \25844 , \25845 , \25846 ,
         \25847 , \25848 , \25849 , \25850 , \25851 , \25852 , \25853 , \25854 , \25855 , \25856 ,
         \25857 , \25858 , \25859 , \25860 , \25861 , \25862 , \25863 , \25864 , \25865 , \25866 ,
         \25867 , \25868 , \25869 , \25870 , \25871 , \25872 , \25873 , \25874 , \25875 , \25876 ,
         \25877 , \25878 , \25879 , \25880 , \25881 , \25882 , \25883 , \25884 , \25885 , \25886 ,
         \25887 , \25888 , \25889 , \25890 , \25891 , \25892 , \25893 , \25894 , \25895 , \25896 ,
         \25897 , \25898 , \25899 , \25900 , \25901 , \25902 , \25903 , \25904 , \25905 , \25906 ,
         \25907 , \25908 , \25909 , \25910 , \25911 , \25912 , \25913 , \25914 , \25915 , \25916 ,
         \25917 , \25918 , \25919 , \25920 , \25921 , \25922 , \25923 , \25924 , \25925 , \25926 ,
         \25927 , \25928 , \25929 , \25930 , \25931 , \25932 , \25933 , \25934 , \25935 , \25936 ,
         \25937 , \25938 , \25939 , \25940 , \25941 , \25942 , \25943 , \25944 , \25945 , \25946 ,
         \25947 , \25948 , \25949 , \25950 , \25951 , \25952 , \25953 , \25954 , \25955 , \25956 ,
         \25957 , \25958 , \25959 , \25960 , \25961 , \25962 , \25963 , \25964 , \25965 , \25966 ,
         \25967 , \25968 , \25969 , \25970 , \25971 , \25972 , \25973 , \25974 , \25975 , \25976 ,
         \25977 , \25978 , \25979 , \25980 , \25981 , \25982 , \25983 , \25984 , \25985 , \25986 ,
         \25987 , \25988 , \25989 , \25990 , \25991 , \25992 , \25993 , \25994 , \25995 , \25996 ,
         \25997 , \25998 , \25999 , \26000 , \26001 , \26002 , \26003 , \26004 , \26005 , \26006 ,
         \26007 , \26008 , \26009 , \26010 , \26011 , \26012 , \26013 , \26014 , \26015 , \26016 ,
         \26017 , \26018 , \26019 , \26020 , \26021 , \26022 , \26023 , \26024 , \26025 , \26026 ,
         \26027 , \26028 , \26029 , \26030 , \26031 , \26032 , \26033 , \26034 , \26035 , \26036 ,
         \26037 , \26038 , \26039 , \26040 , \26041 , \26042 , \26043 , \26044 , \26045 , \26046 ,
         \26047 , \26048 , \26049 , \26050 , \26051 , \26052 , \26053 , \26054 , \26055 , \26056 ,
         \26057 , \26058 , \26059 , \26060 , \26061 , \26062 , \26063 , \26064 , \26065 , \26066 ,
         \26067 , \26068 , \26069 , \26070 , \26071 , \26072 , \26073 , \26074 , \26075 , \26076 ,
         \26077 , \26078 , \26079 , \26080 , \26081 , \26082 , \26083 , \26084 , \26085 , \26086 ,
         \26087 , \26088 , \26089 , \26090 , \26091 , \26092 , \26093 , \26094 , \26095 , \26096 ,
         \26097 , \26098 , \26099 , \26100 , \26101 , \26102 , \26103 , \26104 , \26105 , \26106 ,
         \26107 , \26108 , \26109 , \26110 , \26111 , \26112 , \26113 , \26114 , \26115 , \26116 ,
         \26117 , \26118 , \26119 , \26120 , \26121 , \26122 , \26123 , \26124 , \26125 , \26126 ,
         \26127 , \26128 , \26129 , \26130 , \26131 , \26132 , \26133 , \26134 , \26135 , \26136 ,
         \26137 , \26138 , \26139 , \26140 , \26141 , \26142 , \26143 , \26144 , \26145 , \26146 ,
         \26147 , \26148 , \26149 , \26150 , \26151 , \26152 , \26153 , \26154 , \26155 , \26156 ,
         \26157 , \26158 , \26159 , \26160 , \26161 , \26162 , \26163 , \26164 , \26165 , \26166 ,
         \26167 , \26168 , \26169 , \26170 , \26171 , \26172 , \26173 , \26174 , \26175 , \26176 ,
         \26177 , \26178 , \26179 , \26180 , \26181 , \26182 , \26183 , \26184 , \26185 , \26186 ,
         \26187 , \26188 , \26189 , \26190 , \26191 , \26192 , \26193 , \26194 , \26195 , \26196 ,
         \26197 , \26198 , \26199 , \26200 , \26201 , \26202 , \26203 , \26204 , \26205 , \26206 ,
         \26207 , \26208 , \26209 , \26210 , \26211 , \26212 , \26213 , \26214 , \26215 , \26216 ,
         \26217 , \26218 , \26219 , \26220 , \26221 , \26222 , \26223 , \26224 , \26225 , \26226 ,
         \26227 , \26228 , \26229 , \26230 , \26231 , \26232 , \26233 , \26234 , \26235 , \26236 ,
         \26237 , \26238 , \26239 , \26240 , \26241 , \26242 , \26243 , \26244 , \26245 , \26246 ,
         \26247 , \26248 , \26249 , \26250 , \26251 , \26252 , \26253 , \26254 , \26255 , \26256 ,
         \26257 , \26258 , \26259 , \26260 , \26261 , \26262 , \26263 , \26264 , \26265 , \26266 ,
         \26267 , \26268 , \26269 , \26270 , \26271 , \26272 , \26273 , \26274 , \26275 , \26276 ,
         \26277 , \26278 , \26279 , \26280 , \26281 , \26282 , \26283 , \26284 , \26285 , \26286 ,
         \26287 , \26288 , \26289 , \26290 , \26291 , \26292 , \26293 , \26294 , \26295 , \26296 ,
         \26297 , \26298 , \26299 , \26300 , \26301 , \26302 , \26303 , \26304 , \26305 , \26306 ,
         \26307 , \26308 , \26309 , \26310 , \26311 , \26312 , \26313 , \26314 , \26315 , \26316 ,
         \26317 , \26318 , \26319 , \26320 , \26321 , \26322 , \26323 , \26324 , \26325 , \26326 ,
         \26327 , \26328 , \26329 , \26330 , \26331 , \26332 , \26333 , \26334 , \26335 , \26336 ,
         \26337 , \26338 , \26339 , \26340 , \26341 , \26342 , \26343 , \26344 , \26345 , \26346 ,
         \26347 , \26348 , \26349 , \26350 , \26351 , \26352 , \26353 , \26354 , \26355 , \26356 ,
         \26357 , \26358 , \26359 , \26360 , \26361 , \26362 , \26363 , \26364 , \26365 , \26366 ,
         \26367 , \26368 , \26369 , \26370 , \26371 , \26372 , \26373 , \26374 , \26375 , \26376 ,
         \26377 , \26378 , \26379 , \26380 , \26381 , \26382 , \26383 , \26384 , \26385 , \26386 ,
         \26387 , \26388 , \26389 , \26390 , \26391 , \26392 , \26393 , \26394 , \26395 , \26396 ,
         \26397 , \26398 , \26399 , \26400 , \26401 , \26402 , \26403 , \26404 , \26405 , \26406 ,
         \26407 , \26408 , \26409 , \26410 , \26411 , \26412 , \26413 , \26414 , \26415 , \26416 ,
         \26417 , \26418 , \26419 , \26420 , \26421 , \26422 , \26423 , \26424 , \26425 , \26426 ,
         \26427 , \26428 , \26429 , \26430 , \26431 , \26432 , \26433 , \26434 , \26435 , \26436 ,
         \26437 , \26438 , \26439 , \26440 , \26441 , \26442 , \26443 , \26444 , \26445 , \26446 ,
         \26447 , \26448 , \26449 , \26450 , \26451 , \26452 , \26453 , \26454 , \26455 , \26456 ,
         \26457 , \26458 , \26459 , \26460 , \26461 , \26462 , \26463 , \26464 , \26465 , \26466 ,
         \26467 , \26468 , \26469 , \26470 , \26471 , \26472 , \26473 , \26474 , \26475 , \26476 ,
         \26477 , \26478 , \26479 , \26480 , \26481 , \26482 , \26483 , \26484 , \26485 , \26486 ,
         \26487 , \26488 , \26489 , \26490 , \26491 , \26492 , \26493 , \26494 , \26495 , \26496 ,
         \26497 , \26498 , \26499 , \26500 , \26501 , \26502 , \26503 , \26504 , \26505 , \26506 ,
         \26507 , \26508 , \26509 , \26510 , \26511 , \26512 , \26513 , \26514 , \26515 , \26516 ,
         \26517 , \26518 , \26519 , \26520 , \26521 , \26522 , \26523 , \26524 , \26525 , \26526 ,
         \26527 , \26528 , \26529 , \26530 , \26531 , \26532 , \26533 , \26534 , \26535 , \26536 ,
         \26537 , \26538 , \26539 , \26540 , \26541 , \26542 , \26543 , \26544 , \26545 , \26546 ,
         \26547 , \26548 , \26549 , \26550 , \26551 , \26552 , \26553 , \26554 , \26555 , \26556 ,
         \26557 , \26558 , \26559 , \26560 , \26561 , \26562 , \26563 , \26564 , \26565 , \26566 ,
         \26567 , \26568 , \26569 , \26570 , \26571 , \26572 , \26573 , \26574 , \26575 , \26576 ,
         \26577 , \26578 , \26579 , \26580 , \26581 , \26582 , \26583 , \26584 , \26585 , \26586 ,
         \26587 , \26588 , \26589 , \26590 , \26591 , \26592 , \26593 , \26594 , \26595 , \26596 ,
         \26597 , \26598 , \26599 , \26600 , \26601 , \26602 , \26603 , \26604 , \26605 , \26606 ,
         \26607 , \26608 , \26609 , \26610 , \26611 , \26612 , \26613 , \26614 , \26615 , \26616 ,
         \26617 , \26618 , \26619 , \26620 , \26621 , \26622 , \26623 , \26624 , \26625 , \26626 ,
         \26627 , \26628 , \26629 , \26630 , \26631 , \26632 , \26633 , \26634 , \26635 , \26636 ,
         \26637 , \26638 , \26639 , \26640 , \26641 , \26642 , \26643 , \26644 , \26645 , \26646 ,
         \26647 , \26648 , \26649 , \26650 , \26651 , \26652 , \26653 , \26654 , \26655 , \26656 ,
         \26657 , \26658 , \26659 , \26660 , \26661 , \26662 , \26663 , \26664 , \26665 , \26666 ,
         \26667 , \26668 , \26669 , \26670 , \26671 , \26672 , \26673 , \26674 , \26675 , \26676 ,
         \26677 , \26678 , \26679 , \26680 , \26681 , \26682 , \26683 , \26684 , \26685 , \26686 ,
         \26687 , \26688 , \26689 , \26690 , \26691 , \26692 , \26693 , \26694 , \26695 , \26696 ,
         \26697 , \26698 , \26699 , \26700 , \26701 , \26702 , \26703 , \26704 , \26705 , \26706 ,
         \26707 , \26708 , \26709 , \26710 , \26711 , \26712 , \26713 , \26714 , \26715 , \26716 ,
         \26717 , \26718 , \26719 , \26720 , \26721 , \26722 , \26723 , \26724 , \26725 , \26726 ,
         \26727 , \26728 , \26729 , \26730 , \26731 , \26732 , \26733 , \26734 , \26735 , \26736 ,
         \26737 , \26738 , \26739 , \26740 , \26741 , \26742 , \26743 , \26744 , \26745 , \26746 ,
         \26747 , \26748 , \26749 , \26750 , \26751 , \26752 , \26753 , \26754 , \26755 , \26756 ,
         \26757 , \26758 , \26759 , \26760 , \26761 , \26762 , \26763 , \26764 , \26765 , \26766 ,
         \26767 , \26768 , \26769 , \26770 , \26771 , \26772 , \26773 , \26774 , \26775 , \26776 ,
         \26777 , \26778 , \26779 , \26780 , \26781 , \26782 , \26783 , \26784 , \26785 , \26786 ,
         \26787 , \26788 , \26789 , \26790 , \26791 , \26792 , \26793 , \26794 , \26795 , \26796 ,
         \26797 , \26798 , \26799 , \26800 , \26801 , \26802 , \26803 , \26804 , \26805 , \26806 ,
         \26807 , \26808 , \26809 , \26810 , \26811 , \26812 , \26813 , \26814 , \26815 , \26816 ,
         \26817 , \26818 , \26819 , \26820 , \26821 , \26822 , \26823 , \26824 , \26825 , \26826 ,
         \26827 , \26828 , \26829 , \26830 , \26831 , \26832 , \26833 , \26834 , \26835 , \26836 ,
         \26837 , \26838 , \26839 , \26840 , \26841 , \26842 , \26843 , \26844 , \26845 , \26846 ,
         \26847 , \26848 , \26849 , \26850 , \26851 , \26852 , \26853 , \26854 , \26855 , \26856 ,
         \26857 , \26858 , \26859 , \26860 , \26861 , \26862 , \26863 , \26864 , \26865 , \26866 ,
         \26867 , \26868 , \26869 , \26870 , \26871 , \26872 , \26873 , \26874 , \26875 , \26876 ,
         \26877 , \26878 , \26879 , \26880 , \26881 , \26882 , \26883 , \26884 , \26885 , \26886 ,
         \26887 , \26888 , \26889 , \26890 , \26891 , \26892 , \26893 , \26894 , \26895 , \26896 ,
         \26897 , \26898 , \26899 , \26900 , \26901 , \26902 , \26903 , \26904 , \26905 , \26906 ,
         \26907 , \26908 , \26909 , \26910 , \26911 , \26912 , \26913 , \26914 , \26915 , \26916 ,
         \26917 , \26918 , \26919 , \26920 , \26921 , \26922 , \26923 , \26924 , \26925 , \26926 ,
         \26927 , \26928 , \26929 , \26930 , \26931 , \26932 , \26933 , \26934 , \26935 , \26936 ,
         \26937 , \26938 , \26939 , \26940 , \26941 , \26942 , \26943 , \26944 , \26945 , \26946 ,
         \26947 , \26948 , \26949 , \26950 , \26951 , \26952 , \26953 , \26954 , \26955 , \26956 ,
         \26957 , \26958 , \26959 , \26960 , \26961 , \26962 , \26963 , \26964 , \26965 , \26966 ,
         \26967 , \26968 , \26969 , \26970 , \26971 , \26972 , \26973 , \26974 , \26975 , \26976 ,
         \26977 , \26978 , \26979 , \26980 , \26981 , \26982 , \26983 , \26984 , \26985 , \26986 ,
         \26987 , \26988 , \26989 , \26990 , \26991 , \26992 , \26993 , \26994 , \26995 , \26996 ,
         \26997 , \26998 , \26999 , \27000 , \27001 , \27002 , \27003 , \27004 , \27005 , \27006 ,
         \27007 , \27008 , \27009 , \27010 , \27011 , \27012 , \27013 , \27014 , \27015 , \27016 ,
         \27017 , \27018 , \27019 , \27020 , \27021 , \27022 , \27023 , \27024 , \27025 , \27026 ,
         \27027 , \27028 , \27029 , \27030 , \27031 , \27032 , \27033 , \27034 , \27035 , \27036 ,
         \27037 , \27038 , \27039 , \27040 , \27041 , \27042 , \27043 , \27044 , \27045 , \27046 ,
         \27047 , \27048 , \27049 , \27050 , \27051 , \27052 , \27053 , \27054 , \27055 , \27056 ,
         \27057 , \27058 , \27059 , \27060 , \27061 , \27062 , \27063 , \27064 , \27065 , \27066 ,
         \27067 , \27068 , \27069 , \27070 , \27071 , \27072 , \27073 , \27074 , \27075 , \27076 ,
         \27077 , \27078 , \27079 , \27080 , \27081 , \27082 , \27083 , \27084 , \27085 , \27086 ,
         \27087 , \27088 , \27089 , \27090 , \27091 , \27092 , \27093 , \27094 , \27095 , \27096 ,
         \27097 , \27098 , \27099 , \27100 , \27101 , \27102 , \27103 , \27104 , \27105 , \27106 ,
         \27107 , \27108 , \27109 , \27110 , \27111 , \27112 , \27113 , \27114 , \27115 , \27116 ,
         \27117 , \27118 , \27119 , \27120 , \27121 , \27122 , \27123 , \27124 , \27125 , \27126 ,
         \27127 , \27128 , \27129 , \27130 , \27131 , \27132 , \27133 , \27134 , \27135 , \27136 ,
         \27137 , \27138 , \27139 , \27140 , \27141 , \27142 , \27143 , \27144 , \27145 , \27146 ,
         \27147 , \27148 , \27149 , \27150 , \27151 , \27152 , \27153 , \27154 , \27155 , \27156 ,
         \27157 , \27158 , \27159 , \27160 , \27161 , \27162 , \27163 , \27164 , \27165 , \27166 ,
         \27167 , \27168 , \27169 , \27170 , \27171 , \27172 , \27173 , \27174 , \27175 , \27176 ,
         \27177 , \27178 , \27179 , \27180 , \27181 , \27182 , \27183 , \27184 , \27185 , \27186 ,
         \27187 , \27188 , \27189 , \27190 , \27191 , \27192 , \27193 , \27194 , \27195 , \27196 ,
         \27197 , \27198 , \27199 , \27200 , \27201 , \27202 , \27203 , \27204 , \27205 , \27206 ,
         \27207 , \27208 , \27209 , \27210 , \27211 , \27212 , \27213 , \27214 , \27215 , \27216 ,
         \27217 , \27218 , \27219 , \27220 , \27221 , \27222 , \27223 , \27224 , \27225 , \27226 ,
         \27227 , \27228 , \27229 , \27230 , \27231 , \27232 , \27233 , \27234 , \27235 , \27236 ,
         \27237 , \27238 , \27239 , \27240 , \27241 , \27242 , \27243 , \27244 , \27245 , \27246 ,
         \27247 , \27248 , \27249 , \27250 , \27251 , \27252 , \27253 , \27254 , \27255 , \27256 ,
         \27257 , \27258 , \27259 , \27260 , \27261 , \27262 , \27263 , \27264 , \27265 , \27266 ,
         \27267 , \27268 , \27269 , \27270 , \27271 , \27272 , \27273 , \27274 , \27275 , \27276 ,
         \27277 , \27278 , \27279 , \27280 , \27281 , \27282 , \27283 , \27284 , \27285 , \27286 ,
         \27287 , \27288 , \27289 , \27290 , \27291 , \27292 , \27293 , \27294 , \27295 , \27296 ,
         \27297 , \27298 , \27299 , \27300 , \27301 , \27302 , \27303 , \27304 , \27305 , \27306 ,
         \27307 , \27308 , \27309 , \27310 , \27311 , \27312 , \27313 , \27314 , \27315 , \27316 ,
         \27317 , \27318 , \27319 , \27320 , \27321 , \27322 , \27323 , \27324 , \27325 , \27326 ,
         \27327 , \27328 , \27329 , \27330 , \27331 , \27332 , \27333 , \27334 , \27335 , \27336 ,
         \27337 , \27338 , \27339 , \27340 , \27341 , \27342 , \27343 , \27344 , \27345 , \27346 ,
         \27347 , \27348 , \27349 , \27350 , \27351 , \27352 , \27353 , \27354 , \27355 , \27356 ,
         \27357 , \27358 , \27359 , \27360 , \27361 , \27362 , \27363 , \27364 , \27365 , \27366 ,
         \27367 , \27368 , \27369 , \27370 , \27371 , \27372 , \27373 , \27374 , \27375 , \27376 ,
         \27377 , \27378 , \27379 , \27380 , \27381 , \27382 , \27383 , \27384 , \27385 , \27386 ,
         \27387 , \27388 , \27389 , \27390 , \27391 , \27392 , \27393 , \27394 , \27395 , \27396 ,
         \27397 , \27398 , \27399 , \27400 , \27401 , \27402 , \27403 , \27404 , \27405 , \27406 ,
         \27407 , \27408 , \27409 , \27410 , \27411 , \27412 , \27413 , \27414 , \27415 , \27416 ,
         \27417 , \27418 , \27419 , \27420 , \27421 , \27422 , \27423 , \27424 , \27425 , \27426 ,
         \27427 , \27428 , \27429 , \27430 , \27431 , \27432 , \27433 , \27434 , \27435 , \27436 ,
         \27437 , \27438 , \27439 , \27440 , \27441 , \27442 , \27443 , \27444 , \27445 , \27446 ,
         \27447 , \27448 , \27449 , \27450 , \27451 , \27452 , \27453 , \27454 , \27455 , \27456 ,
         \27457 , \27458 , \27459 , \27460 , \27461 , \27462 , \27463 , \27464 , \27465 , \27466 ,
         \27467 , \27468 , \27469 , \27470 , \27471 , \27472 , \27473 , \27474 , \27475 , \27476 ,
         \27477 , \27478 , \27479 , \27480 , \27481 , \27482 , \27483 , \27484 , \27485 , \27486 ,
         \27487 , \27488 , \27489 , \27490 , \27491 , \27492 , \27493 , \27494 , \27495 , \27496 ,
         \27497 , \27498 , \27499 , \27500 , \27501 , \27502 , \27503 , \27504 , \27505 , \27506 ,
         \27507 , \27508 , \27509 , \27510 , \27511 , \27512 , \27513 , \27514 , \27515 , \27516 ,
         \27517 , \27518 , \27519 , \27520 , \27521 , \27522 , \27523 , \27524 , \27525 , \27526 ,
         \27527 , \27528 , \27529 , \27530 , \27531 , \27532 , \27533 , \27534 , \27535 , \27536 ,
         \27537 , \27538 , \27539 , \27540 , \27541 , \27542 , \27543 , \27544 , \27545 , \27546 ,
         \27547 , \27548 , \27549 , \27550 , \27551 , \27552 , \27553 , \27554 , \27555 , \27556 ,
         \27557 , \27558 , \27559 , \27560 , \27561 , \27562 , \27563 , \27564 , \27565 , \27566 ,
         \27567 , \27568 , \27569 , \27570 , \27571 , \27572 , \27573 , \27574 , \27575 , \27576 ,
         \27577 , \27578 , \27579 , \27580 , \27581 , \27582 , \27583 , \27584 , \27585 , \27586 ,
         \27587 , \27588 , \27589 , \27590 , \27591 , \27592 , \27593 , \27594 , \27595 , \27596 ,
         \27597 , \27598 , \27599 , \27600 , \27601 , \27602 , \27603 , \27604 , \27605 , \27606 ,
         \27607 , \27608 , \27609 , \27610 , \27611 , \27612 , \27613 , \27614 , \27615 , \27616 ,
         \27617 , \27618 , \27619 , \27620 , \27621 , \27622 , \27623 , \27624 , \27625 , \27626 ,
         \27627 , \27628 , \27629 , \27630 , \27631 , \27632 , \27633 , \27634 , \27635 , \27636 ,
         \27637 , \27638 , \27639 , \27640 , \27641 , \27642 , \27643 , \27644 , \27645 , \27646 ,
         \27647 , \27648 , \27649 , \27650 , \27651 , \27652 , \27653 , \27654 , \27655 , \27656 ,
         \27657 , \27658 , \27659 , \27660 , \27661 , \27662 , \27663 , \27664 , \27665 , \27666 ,
         \27667 , \27668 , \27669 , \27670 , \27671 , \27672 , \27673 , \27674 , \27675 , \27676 ,
         \27677 , \27678 , \27679 , \27680 , \27681 , \27682 , \27683 , \27684 , \27685 , \27686 ,
         \27687 , \27688 , \27689 , \27690 , \27691 , \27692 , \27693 , \27694 , \27695 , \27696 ,
         \27697 , \27698 , \27699 , \27700 , \27701 , \27702 , \27703 , \27704 , \27705 , \27706 ,
         \27707 , \27708 , \27709 , \27710 , \27711 , \27712 , \27713 , \27714 , \27715 , \27716 ,
         \27717 , \27718 , \27719 , \27720 , \27721 , \27722 , \27723 , \27724 , \27725 , \27726 ,
         \27727 , \27728 , \27729 , \27730 , \27731 , \27732 , \27733 , \27734 , \27735 , \27736 ,
         \27737 , \27738 , \27739 , \27740 , \27741 , \27742 , \27743 , \27744 , \27745 , \27746 ,
         \27747 , \27748 , \27749 , \27750 , \27751 , \27752 , \27753 , \27754 , \27755 , \27756 ,
         \27757 , \27758 , \27759 , \27760 , \27761 , \27762 , \27763 , \27764 , \27765 , \27766 ,
         \27767 , \27768 , \27769 , \27770 , \27771 , \27772 , \27773 , \27774 , \27775 , \27776 ,
         \27777 , \27778 , \27779 , \27780 , \27781 , \27782 , \27783 , \27784 , \27785 , \27786 ,
         \27787 , \27788 , \27789 , \27790 , \27791 , \27792 , \27793 , \27794 , \27795 , \27796 ,
         \27797 , \27798 , \27799 , \27800 , \27801 , \27802 , \27803 , \27804 , \27805 , \27806 ,
         \27807 , \27808 , \27809 , \27810 , \27811 , \27812 , \27813 , \27814 , \27815 , \27816 ,
         \27817 , \27818 , \27819 , \27820 , \27821 , \27822 , \27823 , \27824 , \27825 , \27826 ,
         \27827 , \27828 , \27829 , \27830 , \27831 , \27832 , \27833 , \27834 , \27835 , \27836 ,
         \27837 , \27838 , \27839 , \27840 , \27841 , \27842 , \27843 , \27844 , \27845 , \27846 ,
         \27847 , \27848 , \27849 , \27850 , \27851 , \27852 , \27853 , \27854 , \27855 , \27856 ,
         \27857 , \27858 , \27859 , \27860 , \27861 , \27862 , \27863 , \27864 , \27865 , \27866 ,
         \27867 , \27868 , \27869 , \27870 , \27871 , \27872 , \27873 , \27874 , \27875 , \27876 ,
         \27877 , \27878 , \27879 , \27880 , \27881 , \27882 , \27883 , \27884 , \27885 , \27886 ,
         \27887 , \27888 , \27889 , \27890 , \27891 , \27892 , \27893 , \27894 , \27895 , \27896 ,
         \27897 , \27898 , \27899 , \27900 , \27901 , \27902 , \27903 , \27904 , \27905 , \27906 ,
         \27907 , \27908 , \27909 , \27910 , \27911 , \27912 , \27913 , \27914 , \27915 , \27916 ,
         \27917 , \27918 , \27919 , \27920 , \27921 , \27922 , \27923 , \27924 , \27925 , \27926 ,
         \27927 , \27928 , \27929 , \27930 , \27931 , \27932 , \27933 , \27934 , \27935 , \27936 ,
         \27937 , \27938 , \27939 , \27940 , \27941 , \27942 , \27943 , \27944 , \27945 , \27946 ,
         \27947 , \27948 , \27949 , \27950 , \27951 , \27952 , \27953 , \27954 , \27955 , \27956 ,
         \27957 , \27958 , \27959 , \27960 , \27961 , \27962 , \27963 , \27964 , \27965 , \27966 ,
         \27967 , \27968 , \27969 , \27970 , \27971 , \27972 , \27973 , \27974 , \27975 , \27976 ,
         \27977 , \27978 , \27979 , \27980 , \27981 , \27982 , \27983 , \27984 , \27985 , \27986 ,
         \27987 , \27988 , \27989 , \27990 , \27991 , \27992 , \27993 , \27994 , \27995 , \27996 ,
         \27997 , \27998 , \27999 , \28000 , \28001 , \28002 , \28003 , \28004 , \28005 , \28006 ,
         \28007 , \28008 , \28009 , \28010 , \28011 , \28012 , \28013 , \28014 , \28015 , \28016 ,
         \28017 , \28018 , \28019 , \28020 , \28021 , \28022 , \28023 , \28024 , \28025 , \28026 ,
         \28027 , \28028 , \28029 , \28030 , \28031 , \28032 , \28033 , \28034 , \28035 , \28036 ,
         \28037 , \28038 , \28039 , \28040 , \28041 , \28042 , \28043 , \28044 , \28045 , \28046 ,
         \28047 , \28048 , \28049 , \28050 , \28051 , \28052 , \28053 , \28054 , \28055 , \28056 ,
         \28057 , \28058 , \28059 , \28060 , \28061 , \28062 , \28063 , \28064 , \28065 , \28066 ,
         \28067 , \28068 , \28069 , \28070 , \28071 , \28072 , \28073 , \28074 , \28075 , \28076 ,
         \28077 , \28078 , \28079 , \28080 , \28081 , \28082 , \28083 , \28084 , \28085 , \28086 ,
         \28087 , \28088 , \28089 , \28090 , \28091 , \28092 , \28093 , \28094 , \28095 , \28096 ,
         \28097 , \28098 , \28099 , \28100 , \28101 , \28102 , \28103 , \28104 , \28105 , \28106 ,
         \28107 , \28108 , \28109 , \28110 , \28111 , \28112 , \28113 , \28114 , \28115 , \28116 ,
         \28117 , \28118 , \28119 , \28120 , \28121 , \28122 , \28123 , \28124 , \28125 , \28126 ,
         \28127 , \28128 , \28129 , \28130 , \28131 , \28132 , \28133 , \28134 , \28135 , \28136 ,
         \28137 , \28138 , \28139 , \28140 , \28141 , \28142 , \28143 , \28144 , \28145 , \28146 ,
         \28147 , \28148 , \28149 , \28150 , \28151 , \28152 , \28153 , \28154 , \28155 , \28156 ,
         \28157 , \28158 , \28159 , \28160 , \28161 , \28162 , \28163 , \28164 , \28165 , \28166 ,
         \28167 , \28168 , \28169 , \28170 , \28171 , \28172 , \28173 , \28174 , \28175 , \28176 ,
         \28177 , \28178 , \28179 , \28180 , \28181 , \28182 , \28183 , \28184 , \28185 , \28186 ,
         \28187 , \28188 , \28189 , \28190 , \28191 , \28192 , \28193 , \28194 , \28195 , \28196 ,
         \28197 , \28198 , \28199 , \28200 , \28201 , \28202 , \28203 , \28204 , \28205 , \28206 ,
         \28207 , \28208 , \28209 , \28210 , \28211 , \28212 , \28213 , \28214 , \28215 , \28216 ,
         \28217 , \28218 , \28219 , \28220 , \28221 , \28222 , \28223 , \28224 , \28225 , \28226 ,
         \28227 , \28228 , \28229 , \28230 , \28231 , \28232 , \28233 , \28234 , \28235 , \28236 ,
         \28237 , \28238 , \28239 , \28240 , \28241 , \28242 , \28243 , \28244 , \28245 , \28246 ,
         \28247 , \28248 , \28249 , \28250 , \28251 , \28252 , \28253 , \28254 , \28255 , \28256 ,
         \28257 , \28258 , \28259 , \28260 , \28261 , \28262 , \28263 , \28264 , \28265 , \28266 ,
         \28267 , \28268 , \28269 , \28270 , \28271 , \28272 , \28273 , \28274 , \28275 , \28276 ,
         \28277 , \28278 , \28279 , \28280 , \28281 , \28282 , \28283 , \28284 , \28285 , \28286 ,
         \28287 , \28288 , \28289 , \28290 , \28291 , \28292 , \28293 , \28294 , \28295 , \28296 ,
         \28297 , \28298 , \28299 , \28300 , \28301 , \28302 , \28303 , \28304 , \28305 , \28306 ,
         \28307 , \28308 , \28309 , \28310 , \28311 , \28312 , \28313 , \28314 , \28315 , \28316 ,
         \28317 , \28318 , \28319 , \28320 , \28321 , \28322 , \28323 , \28324 , \28325 , \28326 ,
         \28327 , \28328 , \28329 , \28330 , \28331 , \28332 , \28333 , \28334 , \28335 , \28336 ,
         \28337 , \28338 , \28339 , \28340 , \28341 , \28342 , \28343 , \28344 , \28345 , \28346 ,
         \28347 , \28348 , \28349 , \28350 , \28351 , \28352 , \28353 , \28354 , \28355 , \28356 ,
         \28357 , \28358 , \28359 , \28360 , \28361 , \28362 , \28363 , \28364 , \28365 , \28366 ,
         \28367 , \28368 , \28369 , \28370 , \28371 , \28372 , \28373 , \28374 , \28375 , \28376 ,
         \28377 , \28378 , \28379 , \28380 , \28381 , \28382 , \28383 , \28384 , \28385 , \28386 ,
         \28387 , \28388 , \28389 , \28390 , \28391 , \28392 , \28393 , \28394 , \28395 , \28396 ,
         \28397 , \28398 , \28399 , \28400 , \28401 , \28402 , \28403 , \28404 , \28405 , \28406 ,
         \28407 , \28408 , \28409 , \28410 , \28411 , \28412 , \28413 , \28414 , \28415 , \28416 ,
         \28417 , \28418 , \28419 , \28420 , \28421 , \28422 , \28423 , \28424 , \28425 , \28426 ,
         \28427 , \28428 , \28429 , \28430 , \28431 , \28432 , \28433 , \28434 , \28435 , \28436 ,
         \28437 , \28438 , \28439 , \28440 , \28441 , \28442 , \28443 , \28444 , \28445 , \28446 ,
         \28447 , \28448 , \28449 , \28450 , \28451 , \28452 , \28453 , \28454 , \28455 , \28456 ,
         \28457 , \28458 , \28459 , \28460 , \28461 , \28462 , \28463 , \28464 , \28465 , \28466 ,
         \28467 , \28468 , \28469 , \28470 , \28471 , \28472 , \28473 , \28474 , \28475 , \28476 ,
         \28477 , \28478 , \28479 , \28480 , \28481 , \28482 , \28483 , \28484 , \28485 , \28486 ,
         \28487 , \28488 , \28489 , \28490 , \28491 , \28492 , \28493 , \28494 , \28495 , \28496 ,
         \28497 , \28498 , \28499 , \28500 , \28501 , \28502 , \28503 , \28504 , \28505 , \28506 ,
         \28507 , \28508 , \28509 , \28510 , \28511 , \28512 , \28513 , \28514 , \28515 , \28516 ,
         \28517 , \28518 , \28519 , \28520 , \28521 , \28522 , \28523 , \28524 , \28525 , \28526 ,
         \28527 , \28528 , \28529 , \28530 , \28531 , \28532 , \28533 , \28534 , \28535 , \28536 ,
         \28537 , \28538 , \28539 , \28540 , \28541 , \28542 , \28543 , \28544 , \28545 , \28546 ,
         \28547 , \28548 , \28549 , \28550 , \28551 , \28552 , \28553 , \28554 , \28555 , \28556 ,
         \28557 , \28558 , \28559 , \28560 , \28561 , \28562 , \28563 , \28564 , \28565 , \28566 ,
         \28567 , \28568 , \28569 , \28570 , \28571 , \28572 , \28573 , \28574 , \28575 , \28576 ,
         \28577 , \28578 , \28579 , \28580 , \28581 , \28582 , \28583 , \28584 , \28585 , \28586 ,
         \28587 , \28588 , \28589 , \28590 , \28591 , \28592 , \28593 , \28594 , \28595 , \28596 ,
         \28597 , \28598 , \28599 , \28600 , \28601 , \28602 , \28603 , \28604 , \28605 , \28606 ,
         \28607 , \28608 , \28609 , \28610 , \28611 , \28612 , \28613 , \28614 , \28615 , \28616 ,
         \28617 , \28618 , \28619 , \28620 , \28621 , \28622 , \28623 , \28624 , \28625 , \28626 ,
         \28627 , \28628 , \28629 , \28630 , \28631 , \28632 , \28633 , \28634 , \28635 , \28636 ,
         \28637 , \28638 , \28639 , \28640 , \28641 , \28642 , \28643 , \28644 , \28645 , \28646 ,
         \28647 , \28648 , \28649 , \28650 , \28651 , \28652 , \28653 , \28654 , \28655 , \28656 ,
         \28657 , \28658 , \28659 , \28660 , \28661 , \28662 , \28663 , \28664 , \28665 , \28666 ,
         \28667 , \28668 , \28669 , \28670 , \28671 , \28672 , \28673 , \28674 , \28675 , \28676 ,
         \28677 , \28678 , \28679 , \28680 , \28681 , \28682 , \28683 , \28684 , \28685 , \28686 ,
         \28687 , \28688 , \28689 , \28690 , \28691 , \28692 , \28693 , \28694 , \28695 , \28696 ,
         \28697 , \28698 , \28699 , \28700 , \28701 , \28702 , \28703 , \28704 , \28705 , \28706 ,
         \28707 , \28708 , \28709 , \28710 , \28711 , \28712 , \28713 , \28714 , \28715 , \28716 ,
         \28717 , \28718 , \28719 , \28720 , \28721 , \28722 , \28723 , \28724 , \28725 , \28726 ,
         \28727 , \28728 , \28729 , \28730 , \28731 , \28732 , \28733 , \28734 , \28735 , \28736 ,
         \28737 , \28738 , \28739 , \28740 , \28741 , \28742 , \28743 , \28744 , \28745 , \28746 ,
         \28747 , \28748 , \28749 , \28750 , \28751 , \28752 , \28753 , \28754 , \28755 , \28756 ,
         \28757 , \28758 , \28759 , \28760 , \28761 , \28762 , \28763 , \28764 , \28765 , \28766 ,
         \28767 , \28768 , \28769 , \28770 , \28771 , \28772 , \28773 , \28774 , \28775 , \28776 ,
         \28777 , \28778 , \28779 , \28780 , \28781 , \28782 , \28783 , \28784 , \28785 , \28786 ,
         \28787 , \28788 , \28789 , \28790 , \28791 , \28792 , \28793 , \28794 , \28795 , \28796 ,
         \28797 , \28798 , \28799 , \28800 , \28801 , \28802 , \28803 , \28804 , \28805 , \28806 ,
         \28807 , \28808 , \28809 , \28810 , \28811 , \28812 , \28813 , \28814 , \28815 , \28816 ,
         \28817 , \28818 , \28819 , \28820 , \28821 , \28822 , \28823 , \28824 , \28825 , \28826 ,
         \28827 , \28828 , \28829 , \28830 , \28831 , \28832 , \28833 , \28834 , \28835 , \28836 ,
         \28837 , \28838 , \28839 , \28840 , \28841 , \28842 , \28843 , \28844 , \28845 , \28846 ,
         \28847 , \28848 , \28849 , \28850 , \28851 , \28852 , \28853 , \28854 , \28855 , \28856 ,
         \28857 , \28858 , \28859 , \28860 , \28861 , \28862 , \28863 , \28864 , \28865 , \28866 ,
         \28867 , \28868 , \28869 , \28870 , \28871 , \28872 , \28873 , \28874 , \28875 , \28876 ,
         \28877 , \28878 , \28879 , \28880 , \28881 , \28882 , \28883 , \28884 , \28885 , \28886 ,
         \28887 , \28888 , \28889 , \28890 , \28891 , \28892 , \28893 , \28894 , \28895 , \28896 ,
         \28897 , \28898 , \28899 , \28900 , \28901 , \28902 , \28903 , \28904 , \28905 , \28906 ,
         \28907 , \28908 , \28909 , \28910 , \28911 , \28912 , \28913 , \28914 , \28915 , \28916 ,
         \28917 , \28918 , \28919 , \28920 , \28921 , \28922 , \28923 , \28924 , \28925 , \28926 ,
         \28927 , \28928 , \28929 , \28930 , \28931 , \28932 , \28933 , \28934 , \28935 , \28936 ,
         \28937 , \28938 , \28939 , \28940 , \28941 , \28942 , \28943 , \28944 , \28945 , \28946 ,
         \28947 , \28948 , \28949 , \28950 , \28951 , \28952 , \28953 , \28954 , \28955 , \28956 ,
         \28957 , \28958 , \28959 , \28960 , \28961 , \28962 , \28963 , \28964 , \28965 , \28966 ,
         \28967 , \28968 , \28969 , \28970 , \28971 , \28972 , \28973 , \28974 , \28975 , \28976 ,
         \28977 , \28978 , \28979 , \28980 , \28981 , \28982 , \28983 , \28984 , \28985 , \28986 ,
         \28987 , \28988 , \28989 , \28990 , \28991 , \28992 , \28993 , \28994 , \28995 , \28996 ,
         \28997 , \28998 , \28999 , \29000 , \29001 , \29002 , \29003 , \29004 , \29005 , \29006 ,
         \29007 , \29008 , \29009 , \29010 , \29011 , \29012 , \29013 , \29014 , \29015 , \29016 ,
         \29017 , \29018 , \29019 , \29020 , \29021 , \29022 , \29023 , \29024 , \29025 , \29026 ,
         \29027 , \29028 , \29029 , \29030 , \29031 , \29032 , \29033 , \29034 , \29035 , \29036 ,
         \29037 , \29038 , \29039 , \29040 , \29041 , \29042 , \29043 , \29044 , \29045 , \29046 ,
         \29047 , \29048 , \29049 , \29050 , \29051 , \29052 , \29053 , \29054 , \29055 , \29056 ,
         \29057 , \29058 , \29059 , \29060 , \29061 , \29062 , \29063 , \29064 , \29065 , \29066 ,
         \29067 , \29068 , \29069 , \29070 , \29071 , \29072 , \29073 , \29074 , \29075 , \29076 ,
         \29077 , \29078 , \29079 , \29080 , \29081 , \29082 , \29083 , \29084 , \29085 , \29086 ,
         \29087 , \29088 , \29089 , \29090 , \29091 , \29092 , \29093 , \29094 , \29095 , \29096 ,
         \29097 , \29098 , \29099 , \29100 , \29101 , \29102 , \29103 , \29104 , \29105 , \29106 ,
         \29107 , \29108 , \29109 , \29110 , \29111 , \29112 , \29113 , \29114 , \29115 , \29116 ,
         \29117 , \29118 , \29119 , \29120 , \29121 , \29122 , \29123 , \29124 , \29125 , \29126 ,
         \29127 , \29128 , \29129 , \29130 , \29131 , \29132 , \29133 , \29134 , \29135 , \29136 ,
         \29137 , \29138 , \29139 , \29140 , \29141 , \29142 , \29143 , \29144 , \29145 , \29146 ,
         \29147 , \29148 , \29149 , \29150 , \29151 , \29152 , \29153 , \29154 , \29155 , \29156 ,
         \29157 , \29158 , \29159 , \29160 , \29161 , \29162 , \29163 , \29164 , \29165 , \29166 ,
         \29167 , \29168 , \29169 , \29170 , \29171 , \29172 , \29173 , \29174 , \29175 , \29176 ,
         \29177 , \29178 , \29179 , \29180 , \29181 , \29182 , \29183 , \29184 , \29185 , \29186 ,
         \29187 , \29188 , \29189 , \29190 , \29191 , \29192 , \29193 , \29194 , \29195 , \29196 ,
         \29197 , \29198 , \29199 , \29200 , \29201 , \29202 , \29203 , \29204 , \29205 , \29206 ,
         \29207 , \29208 , \29209 , \29210 , \29211 , \29212 , \29213 , \29214 , \29215 , \29216 ,
         \29217 , \29218 , \29219 , \29220 , \29221 , \29222 , \29223 , \29224 , \29225 , \29226 ,
         \29227 , \29228 , \29229 , \29230 , \29231 , \29232 , \29233 , \29234 , \29235 , \29236 ,
         \29237 , \29238 , \29239 , \29240 , \29241 , \29242 , \29243 , \29244 , \29245 , \29246 ,
         \29247 , \29248 , \29249 , \29250 , \29251 , \29252 , \29253 , \29254 , \29255 , \29256 ,
         \29257 , \29258 , \29259 , \29260 , \29261 , \29262 , \29263 , \29264 , \29265 , \29266 ,
         \29267 , \29268 , \29269 , \29270 , \29271 , \29272 , \29273 , \29274 , \29275 , \29276 ,
         \29277 , \29278 , \29279 , \29280 , \29281 , \29282 , \29283 , \29284 , \29285 , \29286 ,
         \29287 , \29288 , \29289 , \29290 , \29291 , \29292 , \29293 , \29294 , \29295 , \29296 ,
         \29297 , \29298 , \29299 , \29300 , \29301 , \29302 , \29303 , \29304 , \29305 , \29306 ,
         \29307 , \29308 , \29309 , \29310 , \29311 , \29312 , \29313 , \29314 , \29315 , \29316 ,
         \29317 , \29318 , \29319 , \29320 , \29321 , \29322 , \29323 , \29324 , \29325 , \29326 ,
         \29327 , \29328 , \29329 , \29330 , \29331 , \29332 , \29333 , \29334 , \29335 , \29336 ,
         \29337 , \29338 , \29339 , \29340 , \29341 , \29342 , \29343 , \29344 , \29345 , \29346 ,
         \29347 , \29348 , \29349 , \29350 , \29351 , \29352 , \29353 , \29354 , \29355 , \29356 ,
         \29357 , \29358 , \29359 , \29360 , \29361 , \29362 , \29363 , \29364 , \29365 , \29366 ,
         \29367 , \29368 , \29369 , \29370 , \29371 , \29372 , \29373 , \29374 , \29375 , \29376 ,
         \29377 , \29378 , \29379 , \29380 , \29381 , \29382 , \29383 , \29384 , \29385 , \29386 ,
         \29387 , \29388 , \29389 , \29390 , \29391 , \29392 , \29393 , \29394 , \29395 , \29396 ,
         \29397 , \29398 , \29399 , \29400 , \29401 , \29402 , \29403 , \29404 , \29405 , \29406 ,
         \29407 , \29408 , \29409 , \29410 , \29411 , \29412 , \29413 , \29414 , \29415 , \29416 ,
         \29417 , \29418 , \29419 , \29420 , \29421 , \29422 , \29423 , \29424 , \29425 , \29426 ,
         \29427 , \29428 , \29429 , \29430 , \29431 , \29432 , \29433 , \29434 , \29435 , \29436 ,
         \29437 , \29438 , \29439 , \29440 , \29441 , \29442 , \29443 , \29444 , \29445 , \29446 ,
         \29447 , \29448 , \29449 , \29450 , \29451 , \29452 , \29453 , \29454 , \29455 , \29456 ,
         \29457 , \29458 , \29459 , \29460 , \29461 , \29462 , \29463 , \29464 , \29465 , \29466 ,
         \29467 , \29468 , \29469 , \29470 , \29471 , \29472 , \29473 , \29474 , \29475 , \29476 ,
         \29477 , \29478 , \29479 , \29480 , \29481 , \29482 , \29483 , \29484 , \29485 , \29486 ,
         \29487 , \29488 , \29489 , \29490 , \29491 , \29492 , \29493 , \29494 , \29495 , \29496 ,
         \29497 , \29498 , \29499 , \29500 , \29501 , \29502 , \29503 , \29504 , \29505 , \29506 ,
         \29507 , \29508 , \29509 , \29510 , \29511 , \29512 , \29513 , \29514 , \29515 , \29516 ,
         \29517 , \29518 , \29519 , \29520 , \29521 , \29522 , \29523 , \29524 , \29525 , \29526 ,
         \29527 , \29528 , \29529 , \29530 , \29531 , \29532 , \29533 , \29534 , \29535 , \29536 ,
         \29537 , \29538 , \29539 , \29540 , \29541 , \29542 , \29543 , \29544 , \29545 , \29546 ,
         \29547 , \29548 , \29549 , \29550 , \29551 , \29552 , \29553 , \29554 , \29555 , \29556 ,
         \29557 , \29558 , \29559 , \29560 , \29561 , \29562 , \29563 , \29564 , \29565 , \29566 ,
         \29567 , \29568 , \29569 , \29570 , \29571 , \29572 , \29573 , \29574 , \29575 , \29576 ,
         \29577 , \29578 , \29579 , \29580 , \29581 , \29582 , \29583 , \29584 , \29585 , \29586 ,
         \29587 , \29588 , \29589 , \29590 , \29591 , \29592 , \29593 , \29594 , \29595 , \29596 ,
         \29597 , \29598 , \29599 , \29600 , \29601 , \29602 , \29603 , \29604 , \29605 , \29606 ,
         \29607 , \29608 , \29609 , \29610 , \29611 , \29612 , \29613 , \29614 , \29615 , \29616 ,
         \29617 , \29618 , \29619 , \29620 , \29621 , \29622 , \29623 , \29624 , \29625 , \29626 ,
         \29627 , \29628 , \29629 , \29630 , \29631 , \29632 , \29633 , \29634 , \29635 , \29636 ,
         \29637 , \29638 , \29639 , \29640 , \29641 , \29642 , \29643 , \29644 , \29645 , \29646 ,
         \29647 , \29648 , \29649 , \29650 , \29651 , \29652 , \29653 , \29654 , \29655 , \29656 ,
         \29657 , \29658 , \29659 , \29660 , \29661 , \29662 , \29663 , \29664 , \29665 , \29666 ,
         \29667 , \29668 , \29669 , \29670 , \29671 , \29672 , \29673 , \29674 , \29675 , \29676 ,
         \29677 , \29678 , \29679 , \29680 , \29681 , \29682 , \29683 , \29684 , \29685 , \29686 ,
         \29687 , \29688 , \29689 , \29690 , \29691 , \29692 , \29693 , \29694 , \29695 , \29696 ,
         \29697 , \29698 , \29699 , \29700 , \29701 , \29702 , \29703 , \29704 , \29705 , \29706 ,
         \29707 , \29708 , \29709 , \29710 , \29711 , \29712 , \29713 , \29714 , \29715 , \29716 ,
         \29717 , \29718 , \29719 , \29720 , \29721 , \29722 , \29723 , \29724 , \29725 , \29726 ,
         \29727 , \29728 , \29729 , \29730 , \29731 , \29732 , \29733 , \29734 , \29735 , \29736 ,
         \29737 , \29738 , \29739 , \29740 , \29741 , \29742 , \29743 , \29744 , \29745 , \29746 ,
         \29747 , \29748 , \29749 , \29750 , \29751 , \29752 , \29753 , \29754 , \29755 , \29756 ,
         \29757 , \29758 , \29759 , \29760 , \29761 , \29762 , \29763 , \29764 , \29765 , \29766 ,
         \29767 , \29768 , \29769 , \29770 , \29771 , \29772 , \29773 , \29774 , \29775 , \29776 ,
         \29777 , \29778 , \29779 , \29780 , \29781 , \29782 , \29783 , \29784 , \29785 , \29786 ,
         \29787 , \29788 , \29789 , \29790 , \29791 , \29792 , \29793 , \29794 , \29795 , \29796 ,
         \29797 , \29798 , \29799 , \29800 , \29801 , \29802 , \29803 , \29804 , \29805 , \29806 ,
         \29807 , \29808 , \29809 , \29810 , \29811 , \29812 , \29813 , \29814 , \29815 , \29816 ,
         \29817 , \29818 , \29819 , \29820 , \29821 , \29822 , \29823 , \29824 , \29825 , \29826 ,
         \29827 , \29828 , \29829 , \29830 , \29831 , \29832 , \29833 , \29834 , \29835 , \29836 ,
         \29837 , \29838 , \29839 , \29840 , \29841 , \29842 , \29843 , \29844 , \29845 , \29846 ,
         \29847 , \29848 , \29849 , \29850 , \29851 , \29852 , \29853 , \29854 , \29855 , \29856 ,
         \29857 , \29858 , \29859 , \29860 , \29861 , \29862 , \29863 , \29864 , \29865 , \29866 ,
         \29867 , \29868 , \29869 , \29870 , \29871 , \29872 , \29873 , \29874 , \29875 , \29876 ,
         \29877 , \29878 , \29879 , \29880 , \29881 , \29882 , \29883 , \29884 , \29885 , \29886 ,
         \29887 , \29888 , \29889 , \29890 , \29891 , \29892 , \29893 , \29894 , \29895 , \29896 ,
         \29897 , \29898 , \29899 , \29900 , \29901 , \29902 , \29903 , \29904 , \29905 , \29906 ,
         \29907 , \29908 , \29909 , \29910 , \29911 , \29912 , \29913 , \29914 , \29915 , \29916 ,
         \29917 , \29918 , \29919 , \29920 , \29921 , \29922 , \29923 , \29924 , \29925 , \29926 ,
         \29927 , \29928 , \29929 , \29930 , \29931 , \29932 , \29933 , \29934 , \29935 , \29936 ,
         \29937 , \29938 , \29939 , \29940 , \29941 , \29942 , \29943 , \29944 , \29945 , \29946 ,
         \29947 , \29948 , \29949 , \29950 , \29951 , \29952 , \29953 , \29954 , \29955 , \29956 ,
         \29957 , \29958 , \29959 , \29960 , \29961 , \29962 , \29963 , \29964 , \29965 , \29966 ,
         \29967 , \29968 , \29969 , \29970 , \29971 , \29972 , \29973 , \29974 , \29975 , \29976 ,
         \29977 , \29978 , \29979 , \29980 , \29981 , \29982 , \29983 , \29984 , \29985 , \29986 ,
         \29987 , \29988 , \29989 , \29990 , \29991 , \29992 , \29993 , \29994 , \29995 , \29996 ,
         \29997 , \29998 , \29999 , \30000 , \30001 , \30002 , \30003 , \30004 , \30005 , \30006 ,
         \30007 , \30008 , \30009 , \30010 , \30011 , \30012 , \30013 , \30014 , \30015 , \30016 ,
         \30017 , \30018 , \30019 , \30020 , \30021 , \30022 , \30023 , \30024 , \30025 , \30026 ,
         \30027 , \30028 , \30029 , \30030 , \30031 , \30032 , \30033 , \30034 , \30035 , \30036 ,
         \30037 , \30038 , \30039 , \30040 , \30041 , \30042 , \30043 , \30044 , \30045 , \30046 ,
         \30047 , \30048 , \30049 , \30050 , \30051 , \30052 , \30053 , \30054 , \30055 , \30056 ,
         \30057 , \30058 , \30059 , \30060 , \30061 , \30062 , \30063 , \30064 , \30065 , \30066 ,
         \30067 , \30068 , \30069 , \30070 , \30071 , \30072 , \30073 , \30074 , \30075 , \30076 ,
         \30077 , \30078 , \30079 , \30080 , \30081 , \30082 , \30083 , \30084 , \30085 , \30086 ,
         \30087 , \30088 , \30089 , \30090 , \30091 , \30092 , \30093 , \30094 , \30095 , \30096 ,
         \30097 , \30098 , \30099 , \30100 , \30101 , \30102 , \30103 , \30104 , \30105 , \30106 ,
         \30107 , \30108 , \30109 , \30110 , \30111 , \30112 , \30113 , \30114 , \30115 , \30116 ,
         \30117 , \30118 , \30119 , \30120 , \30121 , \30122 , \30123 , \30124 , \30125 , \30126 ,
         \30127 , \30128 , \30129 , \30130 , \30131 , \30132 , \30133 , \30134 , \30135 , \30136 ,
         \30137 , \30138 , \30139 , \30140 , \30141 , \30142 , \30143 , \30144 , \30145 , \30146 ,
         \30147 , \30148 , \30149 , \30150 , \30151 , \30152 , \30153 , \30154 , \30155 , \30156 ,
         \30157 , \30158 , \30159 , \30160 , \30161 , \30162 , \30163 , \30164 , \30165 , \30166 ,
         \30167 , \30168 , \30169 , \30170 , \30171 , \30172 , \30173 , \30174 , \30175 , \30176 ,
         \30177 , \30178 , \30179 , \30180 , \30181 , \30182 , \30183 , \30184 , \30185 , \30186 ,
         \30187 , \30188 , \30189 , \30190 , \30191 , \30192 , \30193 , \30194 , \30195 , \30196 ,
         \30197 , \30198 , \30199 , \30200 , \30201 , \30202 , \30203 , \30204 , \30205 , \30206 ,
         \30207 , \30208 , \30209 , \30210 , \30211 , \30212 , \30213 , \30214 , \30215 , \30216 ,
         \30217 , \30218 , \30219 , \30220 , \30221 , \30222 , \30223 , \30224 , \30225 , \30226 ,
         \30227 , \30228 , \30229 , \30230 , \30231 , \30232 , \30233 , \30234 , \30235 , \30236 ,
         \30237 , \30238 , \30239 , \30240 , \30241 , \30242 , \30243 , \30244 , \30245 , \30246 ,
         \30247 , \30248 , \30249 , \30250 , \30251 , \30252 , \30253 , \30254 , \30255 , \30256 ,
         \30257 , \30258 , \30259 , \30260 , \30261 , \30262 , \30263 , \30264 , \30265 , \30266 ,
         \30267 , \30268 , \30269 , \30270 , \30271 , \30272 , \30273 , \30274 , \30275 , \30276 ,
         \30277 , \30278 , \30279 , \30280 , \30281 , \30282 , \30283 , \30284 , \30285 , \30286 ,
         \30287 , \30288 , \30289 , \30290 , \30291 , \30292 , \30293 , \30294 , \30295 , \30296 ,
         \30297 , \30298 , \30299 , \30300 , \30301 , \30302 , \30303 , \30304 , \30305 , \30306 ,
         \30307 , \30308 , \30309 , \30310 , \30311 , \30312 , \30313 , \30314 , \30315 , \30316 ,
         \30317 , \30318 , \30319 , \30320 , \30321 , \30322 , \30323 , \30324 , \30325 , \30326 ,
         \30327 , \30328 , \30329 , \30330 , \30331 , \30332 , \30333 , \30334 , \30335 , \30336 ,
         \30337 , \30338 , \30339 , \30340 , \30341 , \30342 , \30343 , \30344 , \30345 , \30346 ,
         \30347 , \30348 , \30349 , \30350 , \30351 , \30352 , \30353 , \30354 , \30355 , \30356 ,
         \30357 , \30358 , \30359 , \30360 , \30361 , \30362 , \30363 , \30364 , \30365 , \30366 ,
         \30367 , \30368 , \30369 , \30370 , \30371 , \30372 , \30373 , \30374 , \30375 , \30376 ,
         \30377 , \30378 , \30379 , \30380 , \30381 , \30382 , \30383 , \30384 , \30385 , \30386 ,
         \30387 , \30388 , \30389 , \30390 , \30391 , \30392 , \30393 , \30394 , \30395 , \30396 ,
         \30397 , \30398 , \30399 , \30400 , \30401 , \30402 , \30403 , \30404 , \30405 , \30406 ,
         \30407 , \30408 , \30409 , \30410 , \30411 , \30412 , \30413 , \30414 , \30415 , \30416 ,
         \30417 , \30418 , \30419 , \30420 , \30421 , \30422 , \30423 , \30424 , \30425 , \30426 ,
         \30427 , \30428 , \30429 , \30430 , \30431 , \30432 , \30433 , \30434 , \30435 , \30436 ,
         \30437 , \30438 , \30439 , \30440 , \30441 , \30442 , \30443 , \30444 , \30445 , \30446 ,
         \30447 , \30448 , \30449 , \30450 , \30451 , \30452 , \30453 , \30454 , \30455 , \30456 ,
         \30457 , \30458 , \30459 , \30460 , \30461 , \30462 , \30463 , \30464 , \30465 , \30466 ,
         \30467 , \30468 , \30469 , \30470 , \30471 , \30472 , \30473 , \30474 , \30475 , \30476 ,
         \30477 , \30478 , \30479 , \30480 , \30481 , \30482 , \30483 , \30484 , \30485 , \30486 ,
         \30487 , \30488 , \30489 , \30490 , \30491 , \30492 , \30493 , \30494 , \30495 , \30496 ,
         \30497 , \30498 , \30499 , \30500 , \30501 , \30502 , \30503 , \30504 , \30505 , \30506 ,
         \30507 , \30508 , \30509 , \30510 , \30511 , \30512 , \30513 , \30514 , \30515 , \30516 ,
         \30517 , \30518 , \30519 , \30520 , \30521 , \30522 , \30523 , \30524 , \30525 , \30526 ,
         \30527 , \30528 , \30529 , \30530 , \30531 , \30532 , \30533 , \30534 , \30535 , \30536 ,
         \30537 , \30538 , \30539 , \30540 , \30541 , \30542 , \30543 , \30544 , \30545 , \30546 ,
         \30547 , \30548 , \30549 , \30550 , \30551 , \30552 , \30553 , \30554 , \30555 , \30556 ,
         \30557 , \30558 , \30559 , \30560 , \30561 , \30562 , \30563 , \30564 , \30565 , \30566 ,
         \30567 , \30568 , \30569 , \30570 , \30571 , \30572 , \30573 , \30574 , \30575 , \30576 ,
         \30577 , \30578 , \30579 , \30580 , \30581 , \30582 , \30583 , \30584 , \30585 , \30586 ,
         \30587 , \30588 , \30589 , \30590 , \30591 , \30592 , \30593 , \30594 , \30595 , \30596 ,
         \30597 , \30598 , \30599 , \30600 , \30601 , \30602 , \30603 , \30604 , \30605 , \30606 ,
         \30607 , \30608 , \30609 , \30610 , \30611 , \30612 , \30613 , \30614 , \30615 , \30616 ,
         \30617 , \30618 , \30619 , \30620 , \30621 , \30622 , \30623 , \30624 , \30625 , \30626 ,
         \30627 , \30628 , \30629 , \30630 , \30631 , \30632 , \30633 , \30634 , \30635 , \30636 ,
         \30637 , \30638 , \30639 , \30640 , \30641 , \30642 , \30643 , \30644 , \30645 , \30646 ,
         \30647 , \30648 , \30649 , \30650 , \30651 , \30652 , \30653 , \30654 , \30655 , \30656 ,
         \30657 , \30658 , \30659 , \30660 , \30661 , \30662 , \30663 , \30664 , \30665 , \30666 ,
         \30667 , \30668 , \30669 , \30670 , \30671 , \30672 , \30673 , \30674 , \30675 , \30676 ,
         \30677 , \30678 , \30679 , \30680 , \30681 , \30682 , \30683 , \30684 , \30685 , \30686 ,
         \30687 , \30688 , \30689 , \30690 , \30691 , \30692 , \30693 , \30694 , \30695 , \30696 ,
         \30697 , \30698 , \30699 , \30700 , \30701 , \30702 , \30703 , \30704 , \30705 , \30706 ,
         \30707 , \30708 , \30709 , \30710 , \30711 , \30712 , \30713 , \30714 , \30715 , \30716 ,
         \30717 , \30718 , \30719 , \30720 , \30721 , \30722 , \30723 , \30724 , \30725 , \30726 ,
         \30727 , \30728 , \30729 , \30730 , \30731 , \30732 , \30733 , \30734 , \30735 , \30736 ,
         \30737 , \30738 , \30739 , \30740 , \30741 , \30742 , \30743 , \30744 , \30745 , \30746 ,
         \30747 , \30748 , \30749 , \30750 , \30751 , \30752 , \30753 , \30754 , \30755 , \30756 ,
         \30757 , \30758 , \30759 , \30760 , \30761 , \30762 , \30763 , \30764 , \30765 , \30766 ,
         \30767 , \30768 , \30769 , \30770 , \30771 , \30772 , \30773 , \30774 , \30775 , \30776 ,
         \30777 , \30778 , \30779 , \30780 , \30781 , \30782 , \30783 , \30784 , \30785 , \30786 ,
         \30787 , \30788 , \30789 , \30790 , \30791 , \30792 , \30793 , \30794 , \30795 , \30796 ,
         \30797 , \30798 , \30799 , \30800 , \30801 , \30802 , \30803 , \30804 , \30805 , \30806 ,
         \30807 , \30808 , \30809 , \30810 , \30811 , \30812 , \30813 , \30814 , \30815 , \30816 ,
         \30817 , \30818 , \30819 , \30820 , \30821 , \30822 , \30823 , \30824 , \30825 , \30826 ,
         \30827 , \30828 , \30829 , \30830 , \30831 , \30832 , \30833 , \30834 , \30835 , \30836 ,
         \30837 , \30838 , \30839 , \30840 , \30841 , \30842 , \30843 , \30844 , \30845 , \30846 ,
         \30847 , \30848 , \30849 , \30850 , \30851 , \30852 , \30853 , \30854 , \30855 , \30856 ,
         \30857 , \30858 , \30859 , \30860 , \30861 , \30862 , \30863 , \30864 , \30865 , \30866 ,
         \30867 , \30868 , \30869 , \30870 , \30871 , \30872 , \30873 , \30874 , \30875 , \30876 ,
         \30877 , \30878 , \30879 , \30880 , \30881 , \30882 , \30883 , \30884 , \30885 , \30886 ,
         \30887 , \30888 , \30889 , \30890 , \30891 , \30892 , \30893 , \30894 , \30895 , \30896 ,
         \30897 , \30898 , \30899 , \30900 , \30901 , \30902 , \30903 , \30904 , \30905 , \30906 ,
         \30907 , \30908 , \30909 , \30910 , \30911 , \30912 , \30913 , \30914 , \30915 , \30916 ,
         \30917 , \30918 , \30919 , \30920 , \30921 , \30922 , \30923 , \30924 , \30925 , \30926 ,
         \30927 , \30928 , \30929 , \30930 , \30931 , \30932 , \30933 , \30934 , \30935 , \30936 ,
         \30937 , \30938 , \30939 , \30940 , \30941 , \30942 , \30943 , \30944 , \30945 , \30946 ,
         \30947 , \30948 , \30949 , \30950 , \30951 , \30952 , \30953 , \30954 , \30955 , \30956 ,
         \30957 , \30958 , \30959 , \30960 , \30961 , \30962 , \30963 , \30964 , \30965 , \30966 ,
         \30967 , \30968 , \30969 , \30970 , \30971 , \30972 , \30973 , \30974 , \30975 , \30976 ,
         \30977 , \30978 , \30979 , \30980 , \30981 , \30982 , \30983 , \30984 , \30985 , \30986 ,
         \30987 , \30988 , \30989 , \30990 , \30991 , \30992 , \30993 , \30994 , \30995 , \30996 ,
         \30997 , \30998 , \30999 , \31000 , \31001 , \31002 , \31003 , \31004 , \31005 , \31006 ,
         \31007 , \31008 , \31009 , \31010 , \31011 , \31012 , \31013 , \31014 , \31015 , \31016 ,
         \31017 , \31018 , \31019 , \31020 , \31021 , \31022 , \31023 , \31024 , \31025 , \31026 ,
         \31027 , \31028 , \31029 , \31030 , \31031 , \31032 , \31033 , \31034 , \31035 , \31036 ,
         \31037 , \31038 , \31039 , \31040 , \31041 , \31042 , \31043 , \31044 , \31045 , \31046 ,
         \31047 , \31048 , \31049 , \31050 , \31051 , \31052 , \31053 , \31054 , \31055 , \31056 ,
         \31057 , \31058 , \31059 , \31060 , \31061 , \31062 , \31063 , \31064 , \31065 , \31066 ,
         \31067 , \31068 , \31069 , \31070 , \31071 , \31072 , \31073 , \31074 , \31075 , \31076 ,
         \31077 , \31078 , \31079 , \31080 , \31081 , \31082 , \31083 , \31084 , \31085 , \31086 ,
         \31087 , \31088 , \31089 , \31090 , \31091 , \31092 , \31093 , \31094 , \31095 , \31096 ,
         \31097 , \31098 , \31099 , \31100 , \31101 , \31102 , \31103 , \31104 , \31105 , \31106 ,
         \31107 , \31108 , \31109 , \31110 , \31111 , \31112 , \31113 , \31114 , \31115 , \31116 ,
         \31117 , \31118 , \31119 , \31120 , \31121 , \31122 , \31123 , \31124 , \31125 , \31126 ,
         \31127 , \31128 , \31129 , \31130 , \31131 , \31132 , \31133 , \31134 , \31135 , \31136 ,
         \31137 , \31138 , \31139 , \31140 , \31141 , \31142 , \31143 , \31144 , \31145 , \31146 ,
         \31147 , \31148 , \31149 , \31150 , \31151 , \31152 , \31153 , \31154 , \31155 , \31156 ,
         \31157 , \31158 , \31159 , \31160 , \31161 , \31162 , \31163 , \31164 , \31165 , \31166 ,
         \31167 , \31168 , \31169 , \31170 , \31171 , \31172 , \31173 , \31174 , \31175 , \31176 ,
         \31177 , \31178 , \31179 , \31180 , \31181 , \31182 , \31183 , \31184 , \31185 , \31186 ,
         \31187 , \31188 , \31189 , \31190 , \31191 , \31192 , \31193 , \31194 , \31195 , \31196 ,
         \31197 , \31198 , \31199 , \31200 , \31201 , \31202 , \31203 , \31204 , \31205 , \31206 ,
         \31207 , \31208 , \31209 , \31210 , \31211 , \31212 , \31213 , \31214 , \31215 , \31216 ,
         \31217 , \31218 , \31219 , \31220 , \31221 , \31222 , \31223 , \31224 , \31225 , \31226 ,
         \31227 , \31228 , \31229 , \31230 , \31231 , \31232 , \31233 , \31234 , \31235 , \31236 ,
         \31237 , \31238 , \31239 , \31240 , \31241 , \31242 , \31243 , \31244 , \31245 , \31246 ,
         \31247 , \31248 , \31249 , \31250 , \31251 , \31252 , \31253 , \31254 , \31255 , \31256 ,
         \31257 , \31258 , \31259 , \31260 , \31261 , \31262 , \31263 , \31264 , \31265 , \31266 ,
         \31267 , \31268 , \31269 , \31270 , \31271 , \31272 , \31273 , \31274 , \31275 , \31276 ,
         \31277 , \31278 , \31279 , \31280 , \31281 , \31282 , \31283 , \31284 , \31285 , \31286 ,
         \31287 , \31288 , \31289 , \31290 , \31291 , \31292 , \31293 , \31294 , \31295 , \31296 ,
         \31297 , \31298 , \31299 , \31300 , \31301 , \31302 , \31303 , \31304 , \31305 , \31306 ,
         \31307 , \31308 , \31309 , \31310 , \31311 , \31312 , \31313 , \31314 , \31315 , \31316 ,
         \31317 , \31318 , \31319 , \31320 , \31321 , \31322 , \31323 , \31324 , \31325 , \31326 ,
         \31327 , \31328 , \31329 , \31330 , \31331 , \31332 , \31333 , \31334 , \31335 , \31336 ,
         \31337 , \31338 , \31339 , \31340 , \31341 , \31342 , \31343 , \31344 , \31345 , \31346 ,
         \31347 , \31348 , \31349 , \31350 , \31351 , \31352 , \31353 , \31354 , \31355 , \31356 ,
         \31357 , \31358 , \31359 , \31360 , \31361 , \31362 , \31363 , \31364 , \31365 , \31366 ,
         \31367 , \31368 , \31369 , \31370 , \31371 , \31372 , \31373 , \31374 , \31375 , \31376 ,
         \31377 , \31378 , \31379 , \31380 , \31381 , \31382 , \31383 , \31384 , \31385 , \31386 ,
         \31387 , \31388 , \31389 , \31390 , \31391 , \31392 , \31393 , \31394 , \31395 , \31396 ,
         \31397 , \31398 , \31399 , \31400 , \31401 , \31402 , \31403 , \31404 , \31405 , \31406 ,
         \31407 , \31408 , \31409 , \31410 , \31411 , \31412 , \31413 , \31414 , \31415 , \31416 ,
         \31417 , \31418 , \31419 , \31420 , \31421 , \31422 , \31423 , \31424 , \31425 , \31426 ,
         \31427 , \31428 , \31429 , \31430 , \31431 , \31432 , \31433 , \31434 , \31435 , \31436 ,
         \31437 , \31438 , \31439 , \31440 , \31441 , \31442 , \31443 , \31444 , \31445 , \31446 ,
         \31447 , \31448 , \31449 , \31450 , \31451 , \31452 , \31453 , \31454 , \31455 , \31456 ,
         \31457 , \31458 , \31459 , \31460 , \31461 , \31462 , \31463 , \31464 , \31465 , \31466 ,
         \31467 , \31468 , \31469 , \31470 , \31471 , \31472 , \31473 , \31474 , \31475 , \31476 ,
         \31477 , \31478 , \31479 , \31480 , \31481 , \31482 , \31483 , \31484 , \31485 , \31486 ,
         \31487 , \31488 , \31489 , \31490 , \31491 , \31492 , \31493 , \31494 , \31495 , \31496 ,
         \31497 , \31498 , \31499 , \31500 , \31501 , \31502 , \31503 , \31504 , \31505 , \31506 ,
         \31507 , \31508 , \31509 , \31510 , \31511 , \31512 , \31513 , \31514 , \31515 , \31516 ,
         \31517 , \31518 , \31519 , \31520 , \31521 , \31522 , \31523 , \31524 , \31525 , \31526 ,
         \31527 , \31528 , \31529 , \31530 , \31531 , \31532 , \31533 , \31534 , \31535 , \31536 ,
         \31537 , \31538 , \31539 , \31540 , \31541 , \31542 , \31543 , \31544 , \31545 , \31546 ,
         \31547 , \31548 , \31549 , \31550 , \31551 , \31552 , \31553 , \31554 , \31555 , \31556 ,
         \31557 , \31558 , \31559 , \31560 , \31561 , \31562 , \31563 , \31564 , \31565 , \31566 ,
         \31567 , \31568 , \31569 , \31570 , \31571 , \31572 , \31573 , \31574 , \31575 , \31576 ,
         \31577 , \31578 , \31579 , \31580 , \31581 , \31582 , \31583 , \31584 , \31585 , \31586 ,
         \31587 , \31588 , \31589 , \31590 , \31591 , \31592 , \31593 , \31594 , \31595 , \31596 ,
         \31597 , \31598 , \31599 , \31600 , \31601 , \31602 , \31603 , \31604 , \31605 , \31606 ,
         \31607 , \31608 , \31609 , \31610 , \31611 , \31612 , \31613 , \31614 , \31615 , \31616 ,
         \31617 , \31618 , \31619 , \31620 , \31621 , \31622 , \31623 , \31624 , \31625 , \31626 ,
         \31627 , \31628 , \31629 , \31630 , \31631 , \31632 , \31633 , \31634 , \31635 , \31636 ,
         \31637 , \31638 , \31639 , \31640 , \31641 , \31642 , \31643 , \31644 , \31645 , \31646 ,
         \31647 , \31648 , \31649 , \31650 , \31651 , \31652 , \31653 , \31654 , \31655 , \31656 ,
         \31657 , \31658 , \31659 , \31660 , \31661 , \31662 , \31663 , \31664 , \31665 , \31666 ,
         \31667 , \31668 , \31669 , \31670 , \31671 , \31672 , \31673 , \31674 , \31675 , \31676 ,
         \31677 , \31678 , \31679 , \31680 , \31681 , \31682 , \31683 , \31684 , \31685 , \31686 ,
         \31687 , \31688 , \31689 , \31690 , \31691 , \31692 , \31693 , \31694 , \31695 , \31696 ,
         \31697 , \31698 , \31699 , \31700 , \31701 , \31702 , \31703 , \31704 , \31705 , \31706 ,
         \31707 , \31708 , \31709 , \31710 , \31711 , \31712 , \31713 , \31714 , \31715 , \31716 ,
         \31717 , \31718 , \31719 , \31720 , \31721 , \31722 , \31723 , \31724 , \31725 , \31726 ,
         \31727 , \31728 , \31729 , \31730 , \31731 , \31732 , \31733 , \31734 , \31735 , \31736 ,
         \31737 , \31738 , \31739 , \31740 , \31741 , \31742 , \31743 , \31744 , \31745 , \31746 ,
         \31747 , \31748 , \31749 , \31750 , \31751 , \31752 , \31753 , \31754 , \31755 , \31756 ,
         \31757 , \31758 , \31759 , \31760 , \31761 , \31762 , \31763 , \31764 , \31765 , \31766 ,
         \31767 , \31768 , \31769 , \31770 , \31771 , \31772 , \31773 , \31774 , \31775 , \31776 ,
         \31777 , \31778 , \31779 , \31780 , \31781 , \31782 , \31783 , \31784 , \31785 , \31786 ,
         \31787 , \31788 , \31789 , \31790 , \31791 , \31792 , \31793 , \31794 , \31795 , \31796 ,
         \31797 , \31798 , \31799 , \31800 , \31801 , \31802 , \31803 , \31804 , \31805 , \31806 ,
         \31807 , \31808 , \31809 , \31810 , \31811 , \31812 , \31813 , \31814 , \31815 , \31816 ,
         \31817 , \31818 , \31819 , \31820 , \31821 , \31822 , \31823 , \31824 , \31825 , \31826 ,
         \31827 , \31828 , \31829 , \31830 , \31831 , \31832 , \31833 , \31834 , \31835 , \31836 ,
         \31837 , \31838 , \31839 , \31840 , \31841 , \31842 , \31843 , \31844 , \31845 , \31846 ,
         \31847 , \31848 , \31849 , \31850 , \31851 , \31852 , \31853 , \31854 , \31855 , \31856 ,
         \31857 , \31858 , \31859 , \31860 , \31861 , \31862 , \31863 , \31864 , \31865 , \31866 ,
         \31867 , \31868 , \31869 , \31870 , \31871 , \31872 , \31873 , \31874 , \31875 , \31876 ,
         \31877 , \31878 , \31879 , \31880 , \31881 , \31882 , \31883 , \31884 , \31885 , \31886 ,
         \31887 , \31888 , \31889 , \31890 , \31891 , \31892 , \31893 , \31894 , \31895 , \31896 ,
         \31897 , \31898 , \31899 , \31900 , \31901 , \31902 , \31903 , \31904 , \31905 , \31906 ,
         \31907 , \31908 , \31909 , \31910 , \31911 , \31912 , \31913 , \31914 , \31915 , \31916 ,
         \31917 , \31918 , \31919 , \31920 , \31921 , \31922 , \31923 , \31924 , \31925 , \31926 ,
         \31927 , \31928 , \31929 , \31930 , \31931 , \31932 , \31933 , \31934 , \31935 , \31936 ,
         \31937 , \31938 , \31939 , \31940 , \31941 , \31942 , \31943 , \31944 , \31945 , \31946 ,
         \31947 , \31948 , \31949 , \31950 , \31951 , \31952 , \31953 , \31954 , \31955 , \31956 ,
         \31957 , \31958 , \31959 , \31960 , \31961 , \31962 , \31963 , \31964 , \31965 , \31966 ,
         \31967 , \31968 , \31969 , \31970 , \31971 , \31972 , \31973 , \31974 , \31975 , \31976 ,
         \31977 , \31978 , \31979 , \31980 , \31981 , \31982 , \31983 , \31984 , \31985 , \31986 ,
         \31987 , \31988 , \31989 , \31990 , \31991 , \31992 , \31993 , \31994 , \31995 , \31996 ,
         \31997 , \31998 , \31999 , \32000 , \32001 , \32002 , \32003 , \32004 , \32005 , \32006 ,
         \32007 , \32008 , \32009 , \32010 , \32011 , \32012 , \32013 , \32014 , \32015 , \32016 ,
         \32017 , \32018 , \32019 , \32020 , \32021 , \32022 , \32023 , \32024 , \32025 , \32026 ,
         \32027 , \32028 , \32029 , \32030 , \32031 , \32032 , \32033 , \32034 , \32035 , \32036 ,
         \32037 , \32038 , \32039 , \32040 , \32041 , \32042 , \32043 , \32044 , \32045 , \32046 ,
         \32047 , \32048 , \32049 , \32050 , \32051 , \32052 , \32053 , \32054 , \32055 , \32056 ,
         \32057 , \32058 , \32059 , \32060 , \32061 , \32062 , \32063 , \32064 , \32065 , \32066 ,
         \32067 , \32068 , \32069 , \32070 , \32071 , \32072 , \32073 , \32074 , \32075 , \32076 ,
         \32077 , \32078 , \32079 , \32080 , \32081 , \32082 , \32083 , \32084 , \32085 , \32086 ,
         \32087 , \32088 , \32089 , \32090 , \32091 , \32092 , \32093 , \32094 , \32095 , \32096 ,
         \32097 , \32098 , \32099 , \32100 , \32101 , \32102 , \32103 , \32104 , \32105 , \32106 ,
         \32107 , \32108 , \32109 , \32110 , \32111 , \32112 , \32113 , \32114 , \32115 , \32116 ,
         \32117 , \32118 , \32119 , \32120 , \32121 , \32122 , \32123 , \32124 , \32125 , \32126 ,
         \32127 , \32128 , \32129 , \32130 , \32131 , \32132 , \32133 , \32134 , \32135 , \32136 ,
         \32137 , \32138 , \32139 , \32140 , \32141 , \32142 , \32143 , \32144 , \32145 , \32146 ,
         \32147 , \32148 , \32149 , \32150 , \32151 , \32152 , \32153 , \32154 , \32155 , \32156 ,
         \32157 , \32158 , \32159 , \32160 , \32161 , \32162 , \32163 , \32164 , \32165 , \32166 ,
         \32167 , \32168 , \32169 , \32170 , \32171 , \32172 , \32173 , \32174 , \32175 , \32176 ,
         \32177 , \32178 , \32179 , \32180 , \32181 , \32182 , \32183 , \32184 , \32185 , \32186 ,
         \32187 , \32188 , \32189 , \32190 , \32191 , \32192 , \32193 , \32194 , \32195 , \32196 ,
         \32197 , \32198 , \32199 , \32200 , \32201 , \32202 , \32203 , \32204 , \32205 , \32206 ,
         \32207 , \32208 , \32209 , \32210 , \32211 , \32212 , \32213 , \32214 , \32215 , \32216 ,
         \32217 , \32218 , \32219 , \32220 , \32221 , \32222 , \32223 , \32224 , \32225 , \32226 ,
         \32227 , \32228 , \32229 , \32230 , \32231 , \32232 , \32233 , \32234 , \32235 , \32236 ,
         \32237 , \32238 , \32239 , \32240 , \32241 , \32242 , \32243 , \32244 , \32245 , \32246 ,
         \32247 , \32248 , \32249 , \32250 , \32251 , \32252 , \32253 , \32254 , \32255 , \32256 ,
         \32257 , \32258 , \32259 , \32260 , \32261 , \32262 , \32263 , \32264 , \32265 , \32266 ,
         \32267 , \32268 , \32269 , \32270 , \32271 , \32272 , \32273 , \32274 , \32275 , \32276 ,
         \32277 , \32278 , \32279 , \32280 , \32281 , \32282 , \32283 , \32284 , \32285 , \32286 ,
         \32287 , \32288 , \32289 , \32290 , \32291 , \32292 , \32293 , \32294 , \32295 , \32296 ,
         \32297 , \32298 , \32299 , \32300 , \32301 , \32302 , \32303 , \32304 , \32305 , \32306 ,
         \32307 , \32308 , \32309 , \32310 , \32311 , \32312 , \32313 , \32314 , \32315 , \32316 ,
         \32317 , \32318 , \32319 , \32320 , \32321 , \32322 , \32323 , \32324 , \32325 , \32326 ,
         \32327 , \32328 , \32329 , \32330 , \32331 , \32332 , \32333 , \32334 , \32335 , \32336 ,
         \32337 , \32338 , \32339 , \32340 , \32341 , \32342 , \32343 , \32344 , \32345 , \32346 ,
         \32347 , \32348 , \32349 , \32350 , \32351 , \32352 , \32353 , \32354 , \32355 , \32356 ,
         \32357 , \32358 , \32359 , \32360 , \32361 , \32362 , \32363 , \32364 , \32365 , \32366 ,
         \32367 , \32368 , \32369 , \32370 , \32371 , \32372 , \32373 , \32374 , \32375 , \32376 ,
         \32377 , \32378 , \32379 , \32380 , \32381 , \32382 , \32383 , \32384 , \32385 , \32386 ,
         \32387 , \32388 , \32389 , \32390 , \32391 , \32392 , \32393 , \32394 , \32395 , \32396 ,
         \32397 , \32398 , \32399 , \32400 , \32401 , \32402 , \32403 , \32404 , \32405 , \32406 ,
         \32407 , \32408 , \32409 , \32410 , \32411 , \32412 , \32413 , \32414 , \32415 , \32416 ,
         \32417 , \32418 , \32419 , \32420 , \32421 , \32422 , \32423 , \32424 , \32425 , \32426 ,
         \32427 , \32428 , \32429 , \32430 , \32431 , \32432 , \32433 , \32434 , \32435 , \32436 ,
         \32437 , \32438 , \32439 , \32440 , \32441 , \32442 , \32443 , \32444 , \32445 , \32446 ,
         \32447 , \32448 , \32449 , \32450 , \32451 , \32452 , \32453 , \32454 , \32455 , \32456 ,
         \32457 , \32458 , \32459 , \32460 , \32461 , \32462 , \32463 , \32464 , \32465 , \32466 ,
         \32467 , \32468 , \32469 , \32470 , \32471 , \32472 , \32473 , \32474 , \32475 , \32476 ,
         \32477 , \32478 , \32479 , \32480 , \32481 , \32482 , \32483 , \32484 , \32485 , \32486 ,
         \32487 , \32488 , \32489 , \32490 , \32491 , \32492 , \32493 , \32494 , \32495 , \32496 ,
         \32497 , \32498 , \32499 , \32500 , \32501 , \32502 , \32503 , \32504 , \32505 , \32506 ,
         \32507 , \32508 , \32509 , \32510 , \32511 , \32512 , \32513 , \32514 , \32515 , \32516 ,
         \32517 , \32518 , \32519 , \32520 , \32521 , \32522 , \32523 , \32524 , \32525 , \32526 ,
         \32527 , \32528 , \32529 , \32530 , \32531 , \32532 , \32533 , \32534 , \32535 , \32536 ,
         \32537 , \32538 , \32539 , \32540 , \32541 , \32542 , \32543 , \32544 , \32545 , \32546 ,
         \32547 , \32548 , \32549 , \32550 , \32551 , \32552 , \32553 , \32554 , \32555 , \32556 ,
         \32557 , \32558 , \32559 , \32560 , \32561 , \32562 , \32563 , \32564 , \32565 , \32566 ,
         \32567 , \32568 , \32569 , \32570 , \32571 , \32572 , \32573 , \32574 , \32575 , \32576 ,
         \32577 , \32578 , \32579 , \32580 , \32581 , \32582 , \32583 , \32584 , \32585 , \32586 ,
         \32587 , \32588 , \32589 , \32590 , \32591 , \32592 , \32593 , \32594 , \32595 , \32596 ,
         \32597 , \32598 , \32599 , \32600 , \32601 , \32602 , \32603 , \32604 , \32605 , \32606 ,
         \32607 , \32608 , \32609 , \32610 , \32611 , \32612 , \32613 , \32614 , \32615 , \32616 ,
         \32617 , \32618 , \32619 , \32620 , \32621 , \32622 , \32623 , \32624 , \32625 , \32626 ,
         \32627 , \32628 , \32629 , \32630 , \32631 , \32632 , \32633 , \32634 , \32635 , \32636 ,
         \32637 , \32638 , \32639 , \32640 , \32641 , \32642 , \32643 , \32644 , \32645 , \32646 ,
         \32647 , \32648 , \32649 , \32650 , \32651 , \32652 , \32653 , \32654 , \32655 , \32656 ,
         \32657 , \32658 , \32659 , \32660 , \32661 , \32662 , \32663 , \32664 , \32665 , \32666 ,
         \32667 , \32668 , \32669 , \32670 , \32671 , \32672 , \32673 , \32674 , \32675 , \32676 ,
         \32677 , \32678 , \32679 , \32680 , \32681 , \32682 , \32683 , \32684 , \32685 , \32686 ,
         \32687 , \32688 , \32689 , \32690 , \32691 , \32692 , \32693 , \32694 , \32695 , \32696 ,
         \32697 , \32698 , \32699 , \32700 , \32701 , \32702 , \32703 , \32704 , \32705 , \32706 ,
         \32707 , \32708 , \32709 , \32710 , \32711 , \32712 , \32713 , \32714 , \32715 , \32716 ,
         \32717 , \32718 , \32719 , \32720 , \32721 , \32722 , \32723 , \32724 , \32725 , \32726 ,
         \32727 , \32728 , \32729 , \32730 , \32731 , \32732 , \32733 , \32734 , \32735 , \32736 ,
         \32737 , \32738 , \32739 , \32740 , \32741 , \32742 , \32743 , \32744 , \32745 , \32746 ,
         \32747 , \32748 , \32749 , \32750 , \32751 , \32752 , \32753 , \32754 , \32755 , \32756 ,
         \32757 , \32758 , \32759 , \32760 , \32761 , \32762 , \32763 , \32764 , \32765 , \32766 ,
         \32767 , \32768 , \32769 , \32770 , \32771 , \32772 , \32773 , \32774 , \32775 , \32776 ,
         \32777 , \32778 , \32779 , \32780 , \32781 , \32782 , \32783 , \32784 , \32785 , \32786 ,
         \32787 , \32788 , \32789 , \32790 , \32791 , \32792 , \32793 , \32794 , \32795 , \32796 ,
         \32797 , \32798 , \32799 , \32800 , \32801 , \32802 , \32803 , \32804 , \32805 , \32806 ,
         \32807 , \32808 , \32809 , \32810 , \32811 , \32812 , \32813 , \32814 , \32815 , \32816 ,
         \32817 , \32818 , \32819 , \32820 , \32821 , \32822 , \32823 , \32824 , \32825 , \32826 ,
         \32827 , \32828 , \32829 , \32830 , \32831 , \32832 , \32833 , \32834 , \32835 , \32836 ,
         \32837 , \32838 , \32839 , \32840 , \32841 , \32842 , \32843 , \32844 , \32845 , \32846 ,
         \32847 , \32848 , \32849 , \32850 , \32851 , \32852 , \32853 , \32854 , \32855 , \32856 ,
         \32857 , \32858 , \32859 , \32860 , \32861 , \32862 , \32863 , \32864 , \32865 , \32866 ,
         \32867 , \32868 , \32869 , \32870 , \32871 , \32872 , \32873 , \32874 , \32875 , \32876 ,
         \32877 , \32878 , \32879 , \32880 , \32881 , \32882 , \32883 , \32884 , \32885 , \32886 ,
         \32887 , \32888 , \32889 , \32890 , \32891 , \32892 , \32893 , \32894 , \32895 , \32896 ,
         \32897 , \32898 , \32899 , \32900 , \32901 , \32902 , \32903 , \32904 , \32905 , \32906 ,
         \32907 , \32908 , \32909 , \32910 , \32911 , \32912 , \32913 , \32914 , \32915 , \32916 ,
         \32917 , \32918 , \32919 , \32920 , \32921 , \32922 , \32923 , \32924 , \32925 , \32926 ,
         \32927 , \32928 , \32929 , \32930 , \32931 , \32932 , \32933 , \32934 , \32935 , \32936 ,
         \32937 , \32938 , \32939 , \32940 , \32941 , \32942 , \32943 , \32944 , \32945 , \32946 ,
         \32947 , \32948 , \32949 , \32950 , \32951 , \32952 , \32953 , \32954 , \32955 , \32956 ,
         \32957 , \32958 , \32959 , \32960 , \32961 , \32962 , \32963 , \32964 , \32965 , \32966 ,
         \32967 , \32968 , \32969 , \32970 , \32971 , \32972 , \32973 , \32974 , \32975 , \32976 ,
         \32977 , \32978 , \32979 , \32980 , \32981 , \32982 , \32983 , \32984 , \32985 , \32986 ,
         \32987 , \32988 , \32989 , \32990 , \32991 , \32992 , \32993 , \32994 , \32995 , \32996 ,
         \32997 , \32998 , \32999 , \33000 , \33001 , \33002 , \33003 , \33004 , \33005 , \33006 ,
         \33007 , \33008 , \33009 , \33010 , \33011 , \33012 , \33013 , \33014 , \33015 , \33016 ,
         \33017 , \33018 , \33019 , \33020 , \33021 , \33022 , \33023 , \33024 , \33025 , \33026 ,
         \33027 , \33028 , \33029 , \33030 , \33031 , \33032 , \33033 , \33034 , \33035 , \33036 ,
         \33037 , \33038 , \33039 , \33040 , \33041 , \33042 , \33043 , \33044 , \33045 , \33046 ,
         \33047 , \33048 , \33049 , \33050 , \33051 , \33052 , \33053 , \33054 , \33055 , \33056 ,
         \33057 , \33058 , \33059 , \33060 , \33061 , \33062 , \33063 , \33064 , \33065 , \33066 ,
         \33067 , \33068 , \33069 , \33070 , \33071 , \33072 , \33073 , \33074 , \33075 , \33076 ,
         \33077 , \33078 , \33079 , \33080 , \33081 , \33082 , \33083 , \33084 , \33085 , \33086 ,
         \33087 , \33088 , \33089 , \33090 , \33091 , \33092 , \33093 , \33094 , \33095 , \33096 ,
         \33097 , \33098 , \33099 , \33100 , \33101 , \33102 , \33103 , \33104 , \33105 , \33106 ,
         \33107 , \33108 , \33109 , \33110 , \33111 , \33112 , \33113 , \33114 , \33115 , \33116 ,
         \33117 , \33118 , \33119 , \33120 , \33121 , \33122 , \33123 , \33124 , \33125 , \33126 ,
         \33127 , \33128 , \33129 , \33130 , \33131 , \33132 , \33133 , \33134 , \33135 , \33136 ,
         \33137 , \33138 , \33139 , \33140 , \33141 , \33142 , \33143 , \33144 , \33145 , \33146 ,
         \33147 , \33148 , \33149 , \33150 , \33151 , \33152 , \33153 , \33154 , \33155 , \33156 ,
         \33157 , \33158 , \33159 , \33160 , \33161 , \33162 , \33163 , \33164 , \33165 , \33166 ,
         \33167 , \33168 , \33169 , \33170 , \33171 , \33172 , \33173 , \33174 , \33175 , \33176 ,
         \33177 , \33178 , \33179 , \33180 , \33181 , \33182 , \33183 , \33184 , \33185 , \33186 ,
         \33187 , \33188 , \33189 , \33190 , \33191 , \33192 , \33193 , \33194 , \33195 , \33196 ,
         \33197 , \33198 , \33199 , \33200 , \33201 , \33202 , \33203 , \33204 , \33205 , \33206 ,
         \33207 , \33208 , \33209 , \33210 , \33211 , \33212 , \33213 , \33214 , \33215 , \33216 ,
         \33217 , \33218 , \33219 , \33220 , \33221 , \33222 , \33223 , \33224 , \33225 , \33226 ,
         \33227 , \33228 , \33229 , \33230 , \33231 , \33232 , \33233 , \33234 , \33235 , \33236 ,
         \33237 , \33238 , \33239 , \33240 , \33241 , \33242 , \33243 , \33244 , \33245 , \33246 ,
         \33247 , \33248 , \33249 , \33250 , \33251 , \33252 , \33253 , \33254 , \33255 , \33256 ,
         \33257 , \33258 , \33259 , \33260 , \33261 , \33262 , \33263 , \33264 , \33265 , \33266 ,
         \33267 , \33268 , \33269 , \33270 , \33271 , \33272 , \33273 , \33274 , \33275 , \33276 ,
         \33277 , \33278 , \33279 , \33280 , \33281 , \33282 , \33283 , \33284 , \33285 , \33286 ,
         \33287 , \33288 , \33289 , \33290 , \33291 , \33292 , \33293 , \33294 , \33295 , \33296 ,
         \33297 , \33298 , \33299 , \33300 , \33301 , \33302 , \33303 , \33304 , \33305 , \33306 ,
         \33307 , \33308 , \33309 , \33310 , \33311 , \33312 , \33313 , \33314 , \33315 , \33316 ,
         \33317 , \33318 , \33319 , \33320 , \33321 , \33322 , \33323 , \33324 , \33325 , \33326 ,
         \33327 , \33328 , \33329 , \33330 , \33331 , \33332 , \33333 , \33334 , \33335 , \33336 ,
         \33337 , \33338 , \33339 , \33340 , \33341 , \33342 , \33343 , \33344 , \33345 , \33346 ,
         \33347 , \33348 , \33349 , \33350 , \33351 , \33352 , \33353 , \33354 , \33355 , \33356 ,
         \33357 , \33358 , \33359 , \33360 , \33361 , \33362 , \33363 , \33364 , \33365 , \33366 ,
         \33367 , \33368 , \33369 , \33370 , \33371 , \33372 , \33373 , \33374 , \33375 , \33376 ,
         \33377 , \33378 , \33379 , \33380 , \33381 , \33382 , \33383 , \33384 , \33385 , \33386 ,
         \33387 , \33388 , \33389 , \33390 , \33391 , \33392 , \33393 , \33394 , \33395 , \33396 ,
         \33397 , \33398 , \33399 , \33400 , \33401 , \33402 , \33403 , \33404 , \33405 , \33406 ,
         \33407 , \33408 , \33409 , \33410 , \33411 , \33412 , \33413 , \33414 , \33415 , \33416 ,
         \33417 , \33418 , \33419 , \33420 , \33421 , \33422 , \33423 , \33424 , \33425 , \33426 ,
         \33427 , \33428 , \33429 , \33430 , \33431 , \33432 , \33433 , \33434 , \33435 , \33436 ,
         \33437 , \33438 , \33439 , \33440 , \33441 , \33442 , \33443 , \33444 , \33445 , \33446 ,
         \33447 , \33448 , \33449 , \33450 , \33451 , \33452 , \33453 , \33454 , \33455 , \33456 ,
         \33457 , \33458 , \33459 , \33460 , \33461 , \33462 , \33463 , \33464 , \33465 , \33466 ,
         \33467 , \33468 , \33469 , \33470 , \33471 , \33472 , \33473 , \33474 , \33475 , \33476 ,
         \33477 , \33478 , \33479 , \33480 , \33481 , \33482 , \33483 , \33484 , \33485 , \33486 ,
         \33487 , \33488 , \33489 , \33490 , \33491 , \33492 , \33493 , \33494 , \33495 , \33496 ,
         \33497 , \33498 , \33499 , \33500 , \33501 , \33502 , \33503 , \33504 , \33505 , \33506 ,
         \33507 , \33508 , \33509 , \33510 , \33511 , \33512 , \33513 , \33514 , \33515 , \33516 ,
         \33517 , \33518 , \33519 , \33520 , \33521 , \33522 , \33523 , \33524 , \33525 , \33526 ,
         \33527 , \33528 , \33529 , \33530 , \33531 , \33532 , \33533 , \33534 , \33535 , \33536 ,
         \33537 , \33538 , \33539 , \33540 , \33541 , \33542 , \33543 , \33544 , \33545 , \33546 ,
         \33547 , \33548 , \33549 , \33550 , \33551 , \33552 , \33553 , \33554 , \33555 , \33556 ,
         \33557 , \33558 , \33559 , \33560 , \33561 , \33562 , \33563 , \33564 , \33565 , \33566 ,
         \33567 , \33568 , \33569 , \33570 , \33571 , \33572 , \33573 , \33574 , \33575 , \33576 ,
         \33577 , \33578 , \33579 , \33580 , \33581 , \33582 , \33583 , \33584 , \33585 , \33586 ,
         \33587 , \33588 , \33589 , \33590 , \33591 , \33592 , \33593 , \33594 , \33595 , \33596 ,
         \33597 , \33598 , \33599 , \33600 , \33601 , \33602 , \33603 , \33604 , \33605 , \33606 ,
         \33607 , \33608 , \33609 , \33610 , \33611 , \33612 , \33613 , \33614 , \33615 , \33616 ,
         \33617 , \33618 , \33619 , \33620 , \33621 , \33622 , \33623 , \33624 , \33625 , \33626 ,
         \33627 , \33628 , \33629 , \33630 , \33631 , \33632 , \33633 , \33634 , \33635 , \33636 ,
         \33637 , \33638 , \33639 , \33640 , \33641 , \33642 , \33643 , \33644 , \33645 , \33646 ,
         \33647 , \33648 , \33649 , \33650 , \33651 , \33652 , \33653 , \33654 , \33655 , \33656 ,
         \33657 , \33658 , \33659 , \33660 , \33661 , \33662 , \33663 , \33664 , \33665 , \33666 ,
         \33667 , \33668 , \33669 , \33670 , \33671 , \33672 , \33673 , \33674 , \33675 , \33676 ,
         \33677 , \33678 , \33679 , \33680 , \33681 , \33682 , \33683 , \33684 , \33685 , \33686 ,
         \33687 , \33688 , \33689 , \33690 , \33691 , \33692 , \33693 , \33694 , \33695 , \33696 ,
         \33697 , \33698 , \33699 , \33700 , \33701 , \33702 , \33703 , \33704 , \33705 , \33706 ,
         \33707 , \33708 , \33709 , \33710 , \33711 , \33712 , \33713 , \33714 , \33715 , \33716 ,
         \33717 , \33718 , \33719 , \33720 , \33721 , \33722 , \33723 , \33724 , \33725 , \33726 ,
         \33727 , \33728 , \33729 , \33730 , \33731 , \33732 , \33733 , \33734 , \33735 , \33736 ,
         \33737 , \33738 , \33739 , \33740 , \33741 , \33742 , \33743 , \33744 , \33745 , \33746 ,
         \33747 , \33748 , \33749 , \33750 , \33751 , \33752 , \33753 , \33754 , \33755 , \33756 ,
         \33757 , \33758 , \33759 , \33760 , \33761 , \33762 , \33763 , \33764 , \33765 , \33766 ,
         \33767 , \33768 , \33769 , \33770 , \33771 , \33772 , \33773 , \33774 , \33775 , \33776 ,
         \33777 , \33778 , \33779 , \33780 , \33781 , \33782 , \33783 , \33784 , \33785 , \33786 ,
         \33787 , \33788 , \33789 , \33790 , \33791 , \33792 , \33793 , \33794 , \33795 , \33796 ,
         \33797 , \33798 , \33799 , \33800 , \33801 , \33802 , \33803 , \33804 , \33805 , \33806 ,
         \33807 , \33808 , \33809 , \33810 , \33811 , \33812 , \33813 , \33814 , \33815 , \33816 ,
         \33817 , \33818 , \33819 , \33820 , \33821 , \33822 , \33823 , \33824 , \33825 , \33826 ,
         \33827 , \33828 , \33829 , \33830 , \33831 , \33832 , \33833 , \33834 , \33835 , \33836 ,
         \33837 , \33838 , \33839 , \33840 , \33841 , \33842 , \33843 , \33844 , \33845 , \33846 ,
         \33847 , \33848 , \33849 , \33850 , \33851 , \33852 , \33853 , \33854 , \33855 , \33856 ,
         \33857 , \33858 , \33859 , \33860 , \33861 , \33862 , \33863 , \33864 , \33865 , \33866 ,
         \33867 , \33868 , \33869 , \33870 , \33871 , \33872 , \33873 , \33874 , \33875 , \33876 ,
         \33877 , \33878 , \33879 , \33880 , \33881 , \33882 , \33883 , \33884 , \33885 , \33886 ,
         \33887 , \33888 , \33889 , \33890 , \33891 , \33892 , \33893 , \33894 , \33895 , \33896 ,
         \33897 , \33898 , \33899 , \33900 , \33901 , \33902 , \33903 , \33904 , \33905 , \33906 ,
         \33907 , \33908 , \33909 , \33910 , \33911 , \33912 , \33913 , \33914 , \33915 , \33916 ,
         \33917 , \33918 , \33919 , \33920 , \33921 , \33922 , \33923 , \33924 , \33925 , \33926 ,
         \33927 , \33928 , \33929 , \33930 , \33931 , \33932 , \33933 , \33934 , \33935 , \33936 ,
         \33937 , \33938 , \33939 , \33940 , \33941 , \33942 , \33943 , \33944 , \33945 , \33946 ,
         \33947 , \33948 , \33949 , \33950 , \33951 , \33952 , \33953 , \33954 , \33955 , \33956 ,
         \33957 , \33958 , \33959 , \33960 , \33961 , \33962 , \33963 , \33964 , \33965 , \33966 ,
         \33967 , \33968 , \33969 , \33970 , \33971 , \33972 , \33973 , \33974 , \33975 , \33976 ,
         \33977 , \33978 , \33979 , \33980 , \33981 , \33982 , \33983 , \33984 , \33985 , \33986 ,
         \33987 , \33988 , \33989 , \33990 , \33991 , \33992 , \33993 , \33994 , \33995 , \33996 ,
         \33997 , \33998 , \33999 , \34000 , \34001 , \34002 , \34003 , \34004 , \34005 , \34006 ,
         \34007 , \34008 , \34009 , \34010 , \34011 , \34012 , \34013 , \34014 , \34015 , \34016 ,
         \34017 , \34018 , \34019 , \34020 , \34021 , \34022 , \34023 , \34024 , \34025 , \34026 ,
         \34027 , \34028 , \34029 , \34030 , \34031 , \34032 , \34033 , \34034 , \34035 , \34036 ,
         \34037 , \34038 , \34039 , \34040 , \34041 , \34042 , \34043 , \34044 , \34045 , \34046 ,
         \34047 , \34048 , \34049 , \34050 , \34051 , \34052 , \34053 , \34054 , \34055 , \34056 ,
         \34057 , \34058 , \34059 , \34060 , \34061 , \34062 , \34063 , \34064 , \34065 , \34066 ,
         \34067 , \34068 , \34069 , \34070 , \34071 , \34072 , \34073 , \34074 , \34075 , \34076 ,
         \34077 , \34078 , \34079 , \34080 , \34081 , \34082 , \34083 , \34084 , \34085 , \34086 ,
         \34087 , \34088 , \34089 , \34090 , \34091 , \34092 , \34093 , \34094 , \34095 , \34096 ,
         \34097 , \34098 , \34099 , \34100 , \34101 , \34102 , \34103 , \34104 , \34105 , \34106 ,
         \34107 , \34108 , \34109 , \34110 , \34111 , \34112 , \34113 , \34114 , \34115 , \34116 ,
         \34117 , \34118 , \34119 , \34120 , \34121 , \34122 , \34123 , \34124 , \34125 , \34126 ,
         \34127 , \34128 , \34129 , \34130 , \34131 , \34132 , \34133 , \34134 , \34135 , \34136 ,
         \34137 , \34138 , \34139 , \34140 , \34141 , \34142 , \34143 , \34144 , \34145 , \34146 ,
         \34147 , \34148 , \34149 , \34150 , \34151 , \34152 , \34153 , \34154 , \34155 , \34156 ,
         \34157 , \34158 , \34159 , \34160 , \34161 , \34162 , \34163 , \34164 , \34165 , \34166 ,
         \34167 , \34168 , \34169 , \34170 , \34171 , \34172 , \34173 , \34174 , \34175 , \34176 ,
         \34177 , \34178 , \34179 , \34180 , \34181 , \34182 , \34183 , \34184 , \34185 , \34186 ,
         \34187 , \34188 , \34189 , \34190 , \34191 , \34192 , \34193 , \34194 , \34195 , \34196 ,
         \34197 , \34198 , \34199 , \34200 , \34201 , \34202 , \34203 , \34204 , \34205 , \34206 ,
         \34207 , \34208 , \34209 , \34210 , \34211 , \34212 , \34213 , \34214 , \34215 , \34216 ,
         \34217 , \34218 , \34219 , \34220 , \34221 , \34222 , \34223 , \34224 , \34225 , \34226 ,
         \34227 , \34228 , \34229 , \34230 , \34231 , \34232 , \34233 , \34234 , \34235 , \34236 ,
         \34237 , \34238 , \34239 , \34240 , \34241 , \34242 , \34243 , \34244 , \34245 , \34246 ,
         \34247 , \34248 , \34249 , \34250 , \34251 , \34252 , \34253 , \34254 , \34255 , \34256 ,
         \34257 , \34258 , \34259 , \34260 , \34261 , \34262 , \34263 , \34264 , \34265 , \34266 ,
         \34267 , \34268 , \34269 , \34270 , \34271 , \34272 , \34273 , \34274 , \34275 , \34276 ,
         \34277 , \34278 , \34279 , \34280 , \34281 , \34282 , \34283 , \34284 , \34285 , \34286 ,
         \34287 , \34288 , \34289 , \34290 , \34291 , \34292 , \34293 , \34294 , \34295 , \34296 ,
         \34297 , \34298 , \34299 , \34300 , \34301 , \34302 , \34303 , \34304 , \34305 , \34306 ,
         \34307 , \34308 , \34309 , \34310 , \34311 , \34312 , \34313 , \34314 , \34315 , \34316 ,
         \34317 , \34318 , \34319 , \34320 , \34321 , \34322 , \34323 , \34324 , \34325 , \34326 ,
         \34327 , \34328 , \34329 , \34330 , \34331 , \34332 , \34333 , \34334 , \34335 , \34336 ,
         \34337 , \34338 , \34339 , \34340 , \34341 , \34342 , \34343 , \34344 , \34345 , \34346 ,
         \34347 , \34348 , \34349 , \34350 , \34351 , \34352 , \34353 , \34354 , \34355 , \34356 ,
         \34357 , \34358 , \34359 , \34360 , \34361 , \34362 , \34363 , \34364 , \34365 , \34366 ,
         \34367 , \34368 , \34369 , \34370 , \34371 , \34372 , \34373 , \34374 , \34375 , \34376 ,
         \34377 , \34378 , \34379 , \34380 , \34381 , \34382 , \34383 , \34384 , \34385 , \34386 ,
         \34387 , \34388 , \34389 , \34390 , \34391 , \34392 , \34393 , \34394 , \34395 , \34396 ,
         \34397 , \34398 , \34399 , \34400 , \34401 , \34402 , \34403 , \34404 , \34405 , \34406 ,
         \34407 , \34408 , \34409 , \34410 , \34411 , \34412 , \34413 , \34414 , \34415 , \34416 ,
         \34417 , \34418 , \34419 , \34420 , \34421 , \34422 , \34423 , \34424 , \34425 , \34426 ,
         \34427 , \34428 , \34429 , \34430 , \34431 , \34432 , \34433 , \34434 , \34435 , \34436 ,
         \34437 , \34438 , \34439 , \34440 , \34441 , \34442 , \34443 , \34444 , \34445 , \34446 ,
         \34447 , \34448 , \34449 , \34450 , \34451 , \34452 , \34453 , \34454 , \34455 , \34456 ,
         \34457 , \34458 , \34459 , \34460 , \34461 , \34462 , \34463 , \34464 , \34465 , \34466 ,
         \34467 , \34468 , \34469 , \34470 , \34471 , \34472 , \34473 , \34474 , \34475 , \34476 ,
         \34477 , \34478 , \34479 , \34480 , \34481 , \34482 , \34483 , \34484 , \34485 , \34486 ,
         \34487 , \34488 , \34489 , \34490 , \34491 , \34492 , \34493 , \34494 , \34495 , \34496 ,
         \34497 , \34498 , \34499 , \34500 , \34501 , \34502 , \34503 , \34504 , \34505 , \34506 ,
         \34507 , \34508 , \34509 , \34510 , \34511 , \34512 , \34513 , \34514 , \34515 , \34516 ,
         \34517 , \34518 , \34519 , \34520 , \34521 , \34522 , \34523 , \34524 , \34525 , \34526 ,
         \34527 , \34528 , \34529 , \34530 , \34531 , \34532 , \34533 , \34534 , \34535 , \34536 ,
         \34537 , \34538 , \34539 , \34540 , \34541 , \34542 , \34543 , \34544 , \34545 , \34546 ,
         \34547 , \34548 , \34549 , \34550 , \34551 , \34552 , \34553 , \34554 , \34555 , \34556 ,
         \34557 , \34558 , \34559 , \34560 , \34561 , \34562 , \34563 , \34564 , \34565 , \34566 ,
         \34567 , \34568 , \34569 , \34570 , \34571 , \34572 , \34573 , \34574 , \34575 , \34576 ,
         \34577 , \34578 , \34579 , \34580 , \34581 , \34582 , \34583 , \34584 , \34585 , \34586 ,
         \34587 , \34588 , \34589 , \34590 , \34591 , \34592 , \34593 , \34594 , \34595 , \34596 ,
         \34597 , \34598 , \34599 , \34600 , \34601 , \34602 , \34603 , \34604 , \34605 , \34606 ,
         \34607 , \34608 , \34609 , \34610 , \34611 , \34612 , \34613 , \34614 , \34615 , \34616 ,
         \34617 , \34618 , \34619 , \34620 , \34621 , \34622 , \34623 , \34624 , \34625 , \34626 ,
         \34627 , \34628 , \34629 , \34630 , \34631 , \34632 , \34633 , \34634 , \34635 , \34636 ,
         \34637 , \34638 , \34639 , \34640 , \34641 , \34642 , \34643 , \34644 , \34645 , \34646 ,
         \34647 , \34648 , \34649 , \34650 , \34651 , \34652 , \34653 , \34654 , \34655 , \34656 ,
         \34657 , \34658 , \34659 , \34660 , \34661 , \34662 , \34663 , \34664 , \34665 , \34666 ,
         \34667 , \34668 , \34669 , \34670 , \34671 , \34672 , \34673 , \34674 , \34675 , \34676 ,
         \34677 , \34678 , \34679 , \34680 , \34681 , \34682 , \34683 , \34684 , \34685 , \34686 ,
         \34687 , \34688 , \34689 , \34690 , \34691 , \34692 , \34693 , \34694 , \34695 , \34696 ,
         \34697 , \34698 , \34699 , \34700 , \34701 , \34702 , \34703 , \34704 , \34705 , \34706 ,
         \34707 , \34708 , \34709 , \34710 , \34711 , \34712 , \34713 , \34714 , \34715 , \34716 ,
         \34717 , \34718 , \34719 , \34720 , \34721 , \34722 , \34723 , \34724 , \34725 , \34726 ,
         \34727 , \34728 , \34729 , \34730 , \34731 , \34732 , \34733 , \34734 , \34735 , \34736 ,
         \34737 , \34738 , \34739 , \34740 , \34741 , \34742 , \34743 , \34744 , \34745 , \34746 ,
         \34747 , \34748 , \34749 , \34750 , \34751 , \34752 , \34753 , \34754 , \34755 , \34756 ,
         \34757 , \34758 , \34759 , \34760 , \34761 , \34762 , \34763 , \34764 , \34765 , \34766 ,
         \34767 , \34768 , \34769 , \34770 , \34771 , \34772 , \34773 , \34774 , \34775 , \34776 ,
         \34777 , \34778 , \34779 , \34780 , \34781 , \34782 , \34783 , \34784 , \34785 , \34786 ,
         \34787 , \34788 , \34789 , \34790 , \34791 , \34792 , \34793 , \34794 , \34795 , \34796 ,
         \34797 , \34798 , \34799 , \34800 , \34801 , \34802 , \34803 , \34804 , \34805 , \34806 ,
         \34807 , \34808 , \34809 , \34810 , \34811 , \34812 , \34813 , \34814 , \34815 , \34816 ,
         \34817 , \34818 , \34819 , \34820 , \34821 , \34822 , \34823 , \34824 , \34825 , \34826 ,
         \34827 , \34828 , \34829 , \34830 , \34831 , \34832 , \34833 , \34834 , \34835 , \34836 ,
         \34837 , \34838 , \34839 , \34840 , \34841 , \34842 , \34843 , \34844 , \34845 , \34846 ,
         \34847 , \34848 , \34849 , \34850 , \34851 , \34852 , \34853 , \34854 , \34855 , \34856 ,
         \34857 , \34858 , \34859 , \34860 , \34861 , \34862 , \34863 , \34864 , \34865 , \34866 ,
         \34867 , \34868 , \34869 , \34870 , \34871 , \34872 , \34873 , \34874 , \34875 , \34876 ,
         \34877 , \34878 , \34879 , \34880 , \34881 , \34882 , \34883 , \34884 , \34885 , \34886 ,
         \34887 , \34888 , \34889 , \34890 , \34891 , \34892 , \34893 , \34894 , \34895 , \34896 ,
         \34897 , \34898 , \34899 , \34900 , \34901 , \34902 , \34903 , \34904 , \34905 , \34906 ,
         \34907 , \34908 , \34909 , \34910 , \34911 , \34912 , \34913 , \34914 , \34915 , \34916 ,
         \34917 , \34918 , \34919 , \34920 , \34921 , \34922 , \34923 , \34924 , \34925 , \34926 ,
         \34927 , \34928 , \34929 , \34930 , \34931 , \34932 , \34933 , \34934 , \34935 , \34936 ,
         \34937 , \34938 , \34939 , \34940 , \34941 , \34942 , \34943 , \34944 , \34945 , \34946 ,
         \34947 , \34948 , \34949 , \34950 , \34951 , \34952 , \34953 , \34954 , \34955 , \34956 ,
         \34957 , \34958 , \34959 , \34960 , \34961 , \34962 , \34963 , \34964 , \34965 , \34966 ,
         \34967 , \34968 , \34969 , \34970 , \34971 , \34972 , \34973 , \34974 , \34975 , \34976 ,
         \34977 , \34978 , \34979 , \34980 , \34981 , \34982 , \34983 , \34984 , \34985 , \34986 ,
         \34987 , \34988 , \34989 , \34990 , \34991 , \34992 , \34993 , \34994 , \34995 , \34996 ,
         \34997 , \34998 , \34999 , \35000 , \35001 , \35002 , \35003 , \35004 , \35005 , \35006 ,
         \35007 , \35008 , \35009 , \35010 , \35011 , \35012 , \35013 , \35014 , \35015 , \35016 ,
         \35017 , \35018 , \35019 , \35020 , \35021 , \35022 , \35023 , \35024 , \35025 , \35026 ,
         \35027 , \35028 , \35029 , \35030 , \35031 , \35032 , \35033 , \35034 , \35035 , \35036 ,
         \35037 , \35038 , \35039 , \35040 , \35041 , \35042 , \35043 , \35044 , \35045 , \35046 ,
         \35047 , \35048 , \35049 , \35050 , \35051 , \35052 , \35053 , \35054 , \35055 , \35056 ,
         \35057 , \35058 , \35059 , \35060 , \35061 , \35062 , \35063 , \35064 , \35065 , \35066 ,
         \35067 , \35068 , \35069 , \35070 , \35071 , \35072 , \35073 , \35074 , \35075 , \35076 ,
         \35077 , \35078 , \35079 , \35080 , \35081 , \35082 , \35083 , \35084 , \35085 , \35086 ,
         \35087 , \35088 , \35089 , \35090 , \35091 , \35092 , \35093 , \35094 , \35095 , \35096 ,
         \35097 , \35098 , \35099 , \35100 , \35101 , \35102 , \35103 , \35104 , \35105 , \35106 ,
         \35107 , \35108 , \35109 , \35110 , \35111 , \35112 , \35113 , \35114 , \35115 , \35116 ,
         \35117 , \35118 , \35119 , \35120 , \35121 , \35122 , \35123 , \35124 , \35125 , \35126 ,
         \35127 , \35128 , \35129 , \35130 , \35131 , \35132 , \35133 , \35134 , \35135 , \35136 ,
         \35137 , \35138 , \35139 , \35140 , \35141 , \35142 , \35143 , \35144 , \35145 , \35146 ,
         \35147 , \35148 , \35149 , \35150 , \35151 , \35152 , \35153 , \35154 , \35155 , \35156 ,
         \35157 , \35158 , \35159 , \35160 , \35161 , \35162 , \35163 , \35164 , \35165 , \35166 ,
         \35167 , \35168 , \35169 , \35170 , \35171 , \35172 , \35173 , \35174 , \35175 , \35176 ,
         \35177 , \35178 , \35179 , \35180 , \35181 , \35182 , \35183 , \35184 , \35185 , \35186 ,
         \35187 , \35188 , \35189 , \35190 , \35191 , \35192 , \35193 , \35194 , \35195 , \35196 ,
         \35197 , \35198 , \35199 , \35200 , \35201 , \35202 , \35203 , \35204 , \35205 , \35206 ,
         \35207 , \35208 , \35209 , \35210 , \35211 , \35212 , \35213 , \35214 , \35215 , \35216 ,
         \35217 , \35218 , \35219 , \35220 , \35221 , \35222 , \35223 , \35224 , \35225 , \35226 ,
         \35227 , \35228 , \35229 , \35230 , \35231 , \35232 , \35233 , \35234 , \35235 , \35236 ,
         \35237 , \35238 , \35239 , \35240 , \35241 , \35242 , \35243 , \35244 , \35245 , \35246 ,
         \35247 , \35248 , \35249 , \35250 , \35251 , \35252 , \35253 , \35254 , \35255 , \35256 ,
         \35257 , \35258 , \35259 , \35260 , \35261 , \35262 , \35263 , \35264 , \35265 , \35266 ,
         \35267 , \35268 , \35269 , \35270 , \35271 , \35272 , \35273 , \35274 , \35275 , \35276 ,
         \35277 , \35278 , \35279 , \35280 , \35281 , \35282 , \35283 , \35284 , \35285 , \35286 ,
         \35287 , \35288 , \35289 , \35290 , \35291 , \35292 , \35293 , \35294 , \35295 , \35296 ,
         \35297 , \35298 , \35299 , \35300 , \35301 , \35302 , \35303 , \35304 , \35305 , \35306 ,
         \35307 , \35308 , \35309 , \35310 , \35311 , \35312 , \35313 , \35314 , \35315 , \35316 ,
         \35317 , \35318 , \35319 , \35320 , \35321 , \35322 , \35323 , \35324 , \35325 , \35326 ,
         \35327 , \35328 , \35329 , \35330 , \35331 , \35332 , \35333 , \35334 , \35335 , \35336 ,
         \35337 , \35338 , \35339 , \35340 , \35341 , \35342 , \35343 , \35344 , \35345 , \35346 ,
         \35347 , \35348 , \35349 , \35350 , \35351 , \35352 , \35353 , \35354 , \35355 , \35356 ,
         \35357 , \35358 , \35359 , \35360 , \35361 , \35362 , \35363 , \35364 , \35365 , \35366 ,
         \35367 , \35368 , \35369 , \35370 , \35371 , \35372 , \35373 , \35374 , \35375 , \35376 ,
         \35377 , \35378 , \35379 , \35380 , \35381 , \35382 , \35383 , \35384 , \35385 , \35386 ,
         \35387 , \35388 , \35389 , \35390 , \35391 , \35392 , \35393 , \35394 , \35395 , \35396 ,
         \35397 , \35398 , \35399 , \35400 , \35401 , \35402 , \35403 , \35404 , \35405 , \35406 ,
         \35407 , \35408 , \35409 , \35410 , \35411 , \35412 , \35413 , \35414 , \35415 , \35416 ,
         \35417 , \35418 , \35419 , \35420 , \35421 , \35422 , \35423 , \35424 , \35425 , \35426 ,
         \35427 , \35428 , \35429 , \35430 , \35431 , \35432 , \35433 , \35434 , \35435 , \35436 ,
         \35437 , \35438 , \35439 , \35440 , \35441 , \35442 , \35443 , \35444 , \35445 , \35446 ,
         \35447 , \35448 , \35449 , \35450 , \35451 , \35452 , \35453 , \35454 , \35455 , \35456 ,
         \35457 , \35458 , \35459 , \35460 , \35461 , \35462 , \35463 , \35464 , \35465 , \35466 ,
         \35467 , \35468 , \35469 , \35470 , \35471 , \35472 , \35473 , \35474 , \35475 , \35476 ,
         \35477 , \35478 , \35479 , \35480 , \35481 , \35482 , \35483 , \35484 , \35485 , \35486 ,
         \35487 , \35488 , \35489 , \35490 , \35491 , \35492 , \35493 , \35494 , \35495 , \35496 ,
         \35497 , \35498 , \35499 , \35500 , \35501 , \35502 , \35503 , \35504 , \35505 , \35506 ,
         \35507 , \35508 , \35509 , \35510 , \35511 , \35512 , \35513 , \35514 , \35515 , \35516 ,
         \35517 , \35518 , \35519 , \35520 , \35521 , \35522 , \35523 , \35524 , \35525 , \35526 ,
         \35527 , \35528 , \35529 , \35530 , \35531 , \35532 , \35533 , \35534 , \35535 , \35536 ,
         \35537 , \35538 , \35539 , \35540 , \35541 , \35542 , \35543 , \35544 , \35545 , \35546 ,
         \35547 , \35548 , \35549 , \35550 , \35551 , \35552 , \35553 , \35554 , \35555 , \35556 ,
         \35557 , \35558 , \35559 , \35560 , \35561 , \35562 , \35563 , \35564 , \35565 , \35566 ,
         \35567 , \35568 , \35569 , \35570 , \35571 , \35572 , \35573 , \35574 , \35575 , \35576 ,
         \35577 , \35578 , \35579 , \35580 , \35581 , \35582 , \35583 , \35584 , \35585 , \35586 ,
         \35587 , \35588 , \35589 , \35590 , \35591 , \35592 , \35593 , \35594 , \35595 , \35596 ,
         \35597 , \35598 , \35599 , \35600 , \35601 , \35602 , \35603 , \35604 , \35605 , \35606 ,
         \35607 , \35608 , \35609 , \35610 , \35611 , \35612 , \35613 , \35614 , \35615 , \35616 ,
         \35617 , \35618 , \35619 , \35620 , \35621 , \35622 , \35623 , \35624 , \35625 , \35626 ,
         \35627 , \35628 , \35629 , \35630 , \35631 , \35632 , \35633 , \35634 , \35635 , \35636 ,
         \35637 , \35638 , \35639 , \35640 , \35641 , \35642 , \35643 , \35644 , \35645 , \35646 ,
         \35647 , \35648 , \35649 , \35650 , \35651 , \35652 , \35653 , \35654 , \35655 , \35656 ,
         \35657 , \35658 , \35659 , \35660 , \35661 , \35662 , \35663 , \35664 , \35665 , \35666 ,
         \35667 , \35668 , \35669 , \35670 , \35671 , \35672 , \35673 , \35674 , \35675 , \35676 ,
         \35677 , \35678 , \35679 , \35680 , \35681 , \35682 , \35683 , \35684 , \35685 , \35686 ,
         \35687 , \35688 , \35689 , \35690 , \35691 , \35692 , \35693 , \35694 , \35695 , \35696 ,
         \35697 , \35698 , \35699 , \35700 , \35701 , \35702 , \35703 , \35704 , \35705 , \35706 ,
         \35707 , \35708 , \35709 , \35710 , \35711 , \35712 , \35713 , \35714 , \35715 , \35716 ,
         \35717 , \35718 , \35719 , \35720 , \35721 , \35722 , \35723 , \35724 , \35725 , \35726 ,
         \35727 , \35728 , \35729 , \35730 , \35731 , \35732 , \35733 , \35734 , \35735 , \35736 ,
         \35737 , \35738 , \35739 , \35740 , \35741 , \35742 , \35743 , \35744 , \35745 , \35746 ,
         \35747 , \35748 , \35749 , \35750 , \35751 , \35752 , \35753 , \35754 , \35755 , \35756 ,
         \35757 , \35758 , \35759 , \35760 , \35761 , \35762 , \35763 , \35764 , \35765 , \35766 ,
         \35767 , \35768 , \35769 , \35770 , \35771 , \35772 , \35773 , \35774 , \35775 , \35776 ,
         \35777 , \35778 , \35779 , \35780 , \35781 , \35782 , \35783 , \35784 , \35785 , \35786 ,
         \35787 , \35788 , \35789 , \35790 , \35791 , \35792 , \35793 , \35794 , \35795 , \35796 ,
         \35797 , \35798 , \35799 , \35800 , \35801 , \35802 , \35803 , \35804 , \35805 , \35806 ,
         \35807 , \35808 , \35809 , \35810 , \35811 , \35812 , \35813 , \35814 , \35815 , \35816 ,
         \35817 , \35818 , \35819 , \35820 , \35821 , \35822 , \35823 , \35824 , \35825 , \35826 ,
         \35827 , \35828 , \35829 , \35830 , \35831 , \35832 , \35833 , \35834 , \35835 , \35836 ,
         \35837 , \35838 , \35839 , \35840 , \35841 , \35842 , \35843 , \35844 , \35845 , \35846 ,
         \35847 , \35848 , \35849 , \35850 , \35851 , \35852 , \35853 , \35854 , \35855 , \35856 ,
         \35857 , \35858 , \35859 , \35860 , \35861 , \35862 , \35863 , \35864 , \35865 , \35866 ,
         \35867 , \35868 , \35869 , \35870 , \35871 , \35872 , \35873 , \35874 , \35875 , \35876 ,
         \35877 , \35878 , \35879 , \35880 , \35881 , \35882 , \35883 , \35884 , \35885 , \35886 ,
         \35887 , \35888 , \35889 , \35890 , \35891 , \35892 , \35893 , \35894 , \35895 , \35896 ,
         \35897 , \35898 , \35899 , \35900 , \35901 , \35902 , \35903 , \35904 , \35905 , \35906 ,
         \35907 , \35908 , \35909 , \35910 , \35911 , \35912 , \35913 , \35914 , \35915 , \35916 ,
         \35917 , \35918 , \35919 , \35920 , \35921 , \35922 , \35923 , \35924 , \35925 , \35926 ,
         \35927 , \35928 , \35929 , \35930 , \35931 , \35932 , \35933 , \35934 , \35935 , \35936 ,
         \35937 , \35938 , \35939 , \35940 , \35941 , \35942 , \35943 , \35944 , \35945 , \35946 ,
         \35947 , \35948 , \35949 , \35950 , \35951 , \35952 , \35953 , \35954 , \35955 , \35956 ,
         \35957 , \35958 , \35959 , \35960 , \35961 , \35962 , \35963 , \35964 , \35965 , \35966 ,
         \35967 , \35968 , \35969 , \35970 , \35971 , \35972 , \35973 , \35974 , \35975 , \35976 ,
         \35977 , \35978 , \35979 , \35980 , \35981 , \35982 , \35983 , \35984 , \35985 , \35986 ,
         \35987 , \35988 , \35989 , \35990 , \35991 , \35992 , \35993 , \35994 , \35995 , \35996 ,
         \35997 , \35998 , \35999 , \36000 , \36001 , \36002 , \36003 , \36004 , \36005 , \36006 ,
         \36007 , \36008 , \36009 , \36010 , \36011 , \36012 , \36013 , \36014 , \36015 , \36016 ,
         \36017 , \36018 , \36019 , \36020 , \36021 , \36022 , \36023 , \36024 , \36025 , \36026 ,
         \36027 , \36028 , \36029 , \36030 , \36031 , \36032 , \36033 , \36034 , \36035 , \36036 ,
         \36037 , \36038 , \36039 , \36040 , \36041 , \36042 , \36043 , \36044 , \36045 , \36046 ,
         \36047 , \36048 , \36049 , \36050 , \36051 , \36052 , \36053 , \36054 , \36055 , \36056 ,
         \36057 , \36058 , \36059 , \36060 , \36061 , \36062 , \36063 , \36064 , \36065 , \36066 ,
         \36067 , \36068 , \36069 , \36070 , \36071 , \36072 , \36073 , \36074 , \36075 , \36076 ,
         \36077 , \36078 , \36079 , \36080 , \36081 , \36082 , \36083 , \36084 , \36085 , \36086 ,
         \36087 , \36088 , \36089 , \36090 , \36091 , \36092 , \36093 , \36094 , \36095 , \36096 ,
         \36097 , \36098 , \36099 , \36100 , \36101 , \36102 , \36103 , \36104 , \36105 , \36106 ,
         \36107 , \36108 , \36109 , \36110 , \36111 , \36112 , \36113 , \36114 , \36115 , \36116 ,
         \36117 , \36118 , \36119 , \36120 , \36121 , \36122 , \36123 , \36124 , \36125 , \36126 ,
         \36127 , \36128 , \36129 , \36130 , \36131 , \36132 , \36133 , \36134 , \36135 , \36136 ,
         \36137 , \36138 , \36139 , \36140 , \36141 , \36142 , \36143 , \36144 , \36145 , \36146 ,
         \36147 , \36148 , \36149 , \36150 , \36151 , \36152 , \36153 , \36154 , \36155 , \36156 ,
         \36157 , \36158 , \36159 , \36160 , \36161 , \36162 , \36163 , \36164 , \36165 , \36166 ,
         \36167 , \36168 , \36169 , \36170 , \36171 , \36172 , \36173 , \36174 , \36175 , \36176 ,
         \36177 , \36178 , \36179 , \36180 , \36181 , \36182 , \36183 , \36184 , \36185 , \36186 ,
         \36187 , \36188 , \36189 , \36190 , \36191 , \36192 , \36193 , \36194 , \36195 , \36196 ,
         \36197 , \36198 , \36199 , \36200 , \36201 , \36202 , \36203 , \36204 , \36205 , \36206 ,
         \36207 , \36208 , \36209 , \36210 , \36211 , \36212 , \36213 , \36214 , \36215 , \36216 ,
         \36217 , \36218 , \36219 , \36220 , \36221 , \36222 , \36223 , \36224 , \36225 , \36226 ,
         \36227 , \36228 , \36229 , \36230 , \36231 , \36232 , \36233 , \36234 , \36235 , \36236 ,
         \36237 , \36238 , \36239 , \36240 , \36241 , \36242 , \36243 , \36244 , \36245 , \36246 ,
         \36247 , \36248 , \36249 , \36250 , \36251 , \36252 , \36253 , \36254 , \36255 , \36256 ,
         \36257 , \36258 , \36259 , \36260 , \36261 , \36262 , \36263 , \36264 , \36265 , \36266 ,
         \36267 , \36268 , \36269 , \36270 , \36271 , \36272 , \36273 , \36274 , \36275 , \36276 ,
         \36277 , \36278 , \36279 , \36280 , \36281 , \36282 , \36283 , \36284 , \36285 , \36286 ,
         \36287 , \36288 , \36289 , \36290 , \36291 , \36292 , \36293 , \36294 , \36295 , \36296 ,
         \36297 , \36298 , \36299 , \36300 , \36301 , \36302 , \36303 , \36304 , \36305 , \36306 ,
         \36307 , \36308 , \36309 , \36310 , \36311 , \36312 , \36313 , \36314 , \36315 , \36316 ,
         \36317 , \36318 , \36319 , \36320 , \36321 , \36322 , \36323 , \36324 , \36325 , \36326 ,
         \36327 , \36328 , \36329 , \36330 , \36331 , \36332 , \36333 , \36334 , \36335 , \36336 ,
         \36337 , \36338 , \36339 , \36340 , \36341 , \36342 , \36343 , \36344 , \36345 , \36346 ,
         \36347 , \36348 , \36349 , \36350 , \36351 , \36352 , \36353 , \36354 , \36355 , \36356 ,
         \36357 , \36358 , \36359 , \36360 , \36361 , \36362 , \36363 , \36364 , \36365 , \36366 ,
         \36367 , \36368 , \36369 , \36370 , \36371 , \36372 , \36373 , \36374 , \36375 , \36376 ,
         \36377 , \36378 , \36379 , \36380 , \36381 , \36382 , \36383 , \36384 , \36385 , \36386 ,
         \36387 , \36388 , \36389 , \36390 , \36391 , \36392 , \36393 , \36394 , \36395 , \36396 ,
         \36397 , \36398 , \36399 , \36400 , \36401 , \36402 , \36403 , \36404 , \36405 , \36406 ,
         \36407 , \36408 , \36409 , \36410 , \36411 , \36412 , \36413 , \36414 , \36415 , \36416 ,
         \36417 , \36418 , \36419 , \36420 , \36421 , \36422 , \36423 , \36424 , \36425 , \36426 ,
         \36427 , \36428 , \36429 , \36430 , \36431 , \36432 , \36433 , \36434 , \36435 , \36436 ,
         \36437 , \36438 , \36439 , \36440 , \36441 , \36442 , \36443 , \36444 , \36445 , \36446 ,
         \36447 , \36448 , \36449 , \36450 , \36451 , \36452 , \36453 , \36454 , \36455 , \36456 ,
         \36457 , \36458 , \36459 , \36460 , \36461 , \36462 , \36463 , \36464 , \36465 , \36466 ,
         \36467 , \36468 , \36469 , \36470 , \36471 , \36472 , \36473 , \36474 , \36475 , \36476 ,
         \36477 , \36478 , \36479 , \36480 , \36481 , \36482 , \36483 , \36484 , \36485 , \36486 ,
         \36487 , \36488 , \36489 , \36490 , \36491 , \36492 , \36493 , \36494 , \36495 , \36496 ,
         \36497 , \36498 , \36499 , \36500 , \36501 , \36502 , \36503 , \36504 , \36505 , \36506 ,
         \36507 , \36508 , \36509 , \36510 , \36511 , \36512 , \36513 , \36514 , \36515 , \36516 ,
         \36517 , \36518 , \36519 , \36520 , \36521 , \36522 , \36523 , \36524 , \36525 , \36526 ,
         \36527 , \36528 , \36529 , \36530 , \36531 , \36532 , \36533 , \36534 , \36535 , \36536 ,
         \36537 , \36538 , \36539 , \36540 , \36541 , \36542 , \36543 , \36544 , \36545 , \36546 ,
         \36547 , \36548 , \36549 , \36550 , \36551 , \36552 , \36553 , \36554 , \36555 , \36556 ,
         \36557 , \36558 , \36559 , \36560 , \36561 , \36562 , \36563 , \36564 , \36565 , \36566 ,
         \36567 , \36568 , \36569 , \36570 , \36571 , \36572 , \36573 , \36574 , \36575 , \36576 ,
         \36577 , \36578 , \36579 , \36580 , \36581 , \36582 , \36583 , \36584 , \36585 , \36586 ,
         \36587 , \36588 , \36589 , \36590 , \36591 , \36592 , \36593 , \36594 , \36595 , \36596 ,
         \36597 , \36598 , \36599 , \36600 , \36601 , \36602 , \36603 , \36604 , \36605 , \36606 ,
         \36607 , \36608 , \36609 , \36610 , \36611 , \36612 , \36613 , \36614 , \36615 , \36616 ,
         \36617 , \36618 , \36619 , \36620 , \36621 , \36622 , \36623 , \36624 , \36625 , \36626 ,
         \36627 , \36628 , \36629 , \36630 , \36631 , \36632 , \36633 , \36634 , \36635 , \36636 ,
         \36637 , \36638 , \36639 , \36640 , \36641 , \36642 , \36643 , \36644 , \36645 , \36646 ,
         \36647 , \36648 , \36649 , \36650 , \36651 , \36652 , \36653 , \36654 , \36655 , \36656 ,
         \36657 , \36658 , \36659 , \36660 , \36661 , \36662 , \36663 , \36664 , \36665 , \36666 ,
         \36667 , \36668 , \36669 , \36670 , \36671 , \36672 , \36673 , \36674 , \36675 , \36676 ,
         \36677 , \36678 , \36679 , \36680 , \36681 , \36682 , \36683 , \36684 , \36685 , \36686 ,
         \36687 , \36688 , \36689 , \36690 , \36691 , \36692 , \36693 , \36694 , \36695 , \36696 ,
         \36697 , \36698 , \36699 , \36700 , \36701 , \36702 , \36703 , \36704 , \36705 , \36706 ,
         \36707 , \36708 , \36709 , \36710 , \36711 , \36712 , \36713 , \36714 , \36715 , \36716 ,
         \36717 , \36718 , \36719 , \36720 , \36721 , \36722 , \36723 , \36724 , \36725 , \36726 ,
         \36727 , \36728 , \36729 , \36730 , \36731 , \36732 , \36733 , \36734 , \36735 , \36736 ,
         \36737 , \36738 , \36739 , \36740 , \36741 , \36742 , \36743 , \36744 , \36745 , \36746 ,
         \36747 , \36748 , \36749 , \36750 , \36751 , \36752 , \36753 , \36754 , \36755 , \36756 ,
         \36757 , \36758 , \36759 , \36760 , \36761 , \36762 , \36763 , \36764 , \36765 , \36766 ,
         \36767 , \36768 , \36769 , \36770 , \36771 , \36772 , \36773 , \36774 , \36775 , \36776 ,
         \36777 , \36778 , \36779 , \36780 , \36781 , \36782 , \36783 , \36784 , \36785 , \36786 ,
         \36787 , \36788 , \36789 , \36790 , \36791 , \36792 , \36793 , \36794 , \36795 , \36796 ,
         \36797 , \36798 , \36799 , \36800 , \36801 , \36802 , \36803 , \36804 , \36805 , \36806 ,
         \36807 , \36808 , \36809 , \36810 , \36811 , \36812 , \36813 , \36814 , \36815 , \36816 ,
         \36817 , \36818 , \36819 , \36820 , \36821 , \36822 , \36823 , \36824 , \36825 , \36826 ,
         \36827 , \36828 , \36829 , \36830 , \36831 , \36832 , \36833 , \36834 , \36835 , \36836 ,
         \36837 , \36838 , \36839 , \36840 , \36841 , \36842 , \36843 , \36844 , \36845 , \36846 ,
         \36847 , \36848 , \36849 , \36850 , \36851 , \36852 , \36853 , \36854 , \36855 , \36856 ,
         \36857 , \36858 , \36859 , \36860 , \36861 , \36862 , \36863 , \36864 , \36865 , \36866 ,
         \36867 , \36868 , \36869 , \36870 , \36871 , \36872 , \36873 , \36874 , \36875 , \36876 ,
         \36877 , \36878 , \36879 , \36880 , \36881 , \36882 , \36883 , \36884 , \36885 , \36886 ,
         \36887 , \36888 , \36889 , \36890 , \36891 , \36892 , \36893 , \36894 , \36895 , \36896 ,
         \36897 , \36898 , \36899 , \36900 , \36901 , \36902 , \36903 , \36904 , \36905 , \36906 ,
         \36907 , \36908 , \36909 , \36910 , \36911 , \36912 , \36913 , \36914 , \36915 , \36916 ,
         \36917 , \36918 , \36919 , \36920 , \36921 , \36922 , \36923 , \36924 , \36925 , \36926 ,
         \36927 , \36928 , \36929 , \36930 , \36931 , \36932 , \36933 , \36934 , \36935 , \36936 ,
         \36937 , \36938 , \36939 , \36940 , \36941 , \36942 , \36943 , \36944 , \36945 , \36946 ,
         \36947 , \36948 , \36949 , \36950 , \36951 , \36952 , \36953 , \36954 , \36955 , \36956 ,
         \36957 , \36958 , \36959 , \36960 , \36961 , \36962 , \36963 , \36964 , \36965 , \36966 ,
         \36967 , \36968 , \36969 , \36970 , \36971 , \36972 , \36973 , \36974 , \36975 , \36976 ,
         \36977 , \36978 , \36979 , \36980 , \36981 , \36982 , \36983 , \36984 , \36985 , \36986 ,
         \36987 , \36988 , \36989 , \36990 , \36991 , \36992 , \36993 , \36994 , \36995 , \36996 ,
         \36997 , \36998 , \36999 , \37000 , \37001 , \37002 , \37003 , \37004 , \37005 , \37006 ,
         \37007 , \37008 , \37009 , \37010 , \37011 , \37012 , \37013 , \37014 , \37015 , \37016 ,
         \37017 , \37018 , \37019 , \37020 , \37021 , \37022 , \37023 , \37024 , \37025 , \37026 ,
         \37027 , \37028 , \37029 , \37030 , \37031 , \37032 , \37033 , \37034 , \37035 , \37036 ,
         \37037 , \37038 , \37039 , \37040 , \37041 , \37042 , \37043 , \37044 , \37045 , \37046 ,
         \37047 , \37048 , \37049 , \37050 , \37051 , \37052 , \37053 , \37054 , \37055 , \37056 ,
         \37057 , \37058 , \37059 , \37060 , \37061 , \37062 , \37063 , \37064 , \37065 , \37066 ,
         \37067 , \37068 , \37069 , \37070 , \37071 , \37072 , \37073 , \37074 , \37075 , \37076 ,
         \37077 , \37078 , \37079 , \37080 , \37081 , \37082 , \37083 , \37084 , \37085 , \37086 ,
         \37087 , \37088 , \37089 , \37090 , \37091 , \37092 , \37093 , \37094 , \37095 , \37096 ,
         \37097 , \37098 , \37099 , \37100 , \37101 , \37102 , \37103 , \37104 , \37105 , \37106 ,
         \37107 , \37108 , \37109 , \37110 , \37111 , \37112 , \37113 , \37114 , \37115 , \37116 ,
         \37117 , \37118 , \37119 , \37120 , \37121 , \37122 , \37123 , \37124 , \37125 , \37126 ,
         \37127 , \37128 , \37129 , \37130 , \37131 , \37132 , \37133 , \37134 , \37135 , \37136 ,
         \37137 , \37138 , \37139 , \37140 , \37141 , \37142 , \37143 , \37144 , \37145 , \37146 ,
         \37147 , \37148 , \37149 , \37150 , \37151 , \37152 , \37153 , \37154 , \37155 , \37156 ,
         \37157 , \37158 , \37159 , \37160 , \37161 , \37162 , \37163 , \37164 , \37165 , \37166 ,
         \37167 , \37168 , \37169 , \37170 , \37171 , \37172 , \37173 , \37174 , \37175 , \37176 ,
         \37177 , \37178 , \37179 , \37180 , \37181 , \37182 , \37183 , \37184 , \37185 , \37186 ,
         \37187 , \37188 , \37189 , \37190 , \37191 , \37192 , \37193 , \37194 , \37195 , \37196 ,
         \37197 , \37198 , \37199 , \37200 , \37201 , \37202 , \37203 , \37204 , \37205 , \37206 ,
         \37207 , \37208 , \37209 , \37210 , \37211 , \37212 , \37213 , \37214 , \37215 , \37216 ,
         \37217 , \37218 , \37219 , \37220 , \37221 , \37222 , \37223 , \37224 , \37225 , \37226 ,
         \37227 , \37228 , \37229 , \37230 , \37231 , \37232 , \37233 , \37234 , \37235 , \37236 ,
         \37237 , \37238 , \37239 , \37240 , \37241 , \37242 , \37243 , \37244 , \37245 , \37246 ,
         \37247 , \37248 , \37249 , \37250 , \37251 , \37252 , \37253 , \37254 , \37255 , \37256 ,
         \37257 , \37258 , \37259 , \37260 , \37261 , \37262 , \37263 , \37264 , \37265 , \37266 ,
         \37267 , \37268 , \37269 , \37270 , \37271 , \37272 , \37273 , \37274 , \37275 , \37276 ,
         \37277 , \37278 , \37279 , \37280 , \37281 , \37282 , \37283 , \37284 , \37285 , \37286 ,
         \37287 , \37288 , \37289 , \37290 , \37291 , \37292 , \37293 , \37294 , \37295 , \37296 ,
         \37297 , \37298 , \37299 , \37300 , \37301 , \37302 , \37303 , \37304 , \37305 , \37306 ,
         \37307 , \37308 , \37309 , \37310 , \37311 , \37312 , \37313 , \37314 , \37315 , \37316 ,
         \37317 , \37318 , \37319 , \37320 , \37321 , \37322 , \37323 , \37324 , \37325 , \37326 ,
         \37327 , \37328 , \37329 , \37330 , \37331 , \37332 , \37333 , \37334 , \37335 , \37336 ,
         \37337 , \37338 , \37339 , \37340 , \37341 , \37342 , \37343 , \37344 , \37345 , \37346 ,
         \37347 , \37348 , \37349 , \37350 , \37351 , \37352 , \37353 , \37354 , \37355 , \37356 ,
         \37357 , \37358 , \37359 , \37360 , \37361 , \37362 , \37363 , \37364 , \37365 , \37366 ,
         \37367 , \37368 , \37369 , \37370 , \37371 , \37372 , \37373 , \37374 , \37375 , \37376 ,
         \37377 , \37378 , \37379 , \37380 , \37381 , \37382 , \37383 , \37384 , \37385 , \37386 ,
         \37387 , \37388 , \37389 , \37390 , \37391 , \37392 , \37393 , \37394 , \37395 , \37396 ,
         \37397 , \37398 , \37399 , \37400 , \37401 , \37402 , \37403 , \37404 , \37405 , \37406 ,
         \37407 , \37408 , \37409 , \37410 , \37411 , \37412 , \37413 , \37414 , \37415 , \37416 ,
         \37417 , \37418 , \37419 , \37420 , \37421 , \37422 , \37423 , \37424 , \37425 , \37426 ,
         \37427 , \37428 , \37429 , \37430 , \37431 , \37432 , \37433 , \37434 , \37435 , \37436 ,
         \37437 , \37438 , \37439 , \37440 , \37441 , \37442 , \37443 , \37444 , \37445 , \37446 ,
         \37447 , \37448 , \37449 , \37450 , \37451 , \37452 , \37453 , \37454 , \37455 , \37456 ,
         \37457 , \37458 , \37459 , \37460 , \37461 , \37462 , \37463 , \37464 , \37465 , \37466 ,
         \37467 , \37468 , \37469 , \37470 , \37471 , \37472 , \37473 , \37474 , \37475 , \37476 ,
         \37477 , \37478 , \37479 , \37480 , \37481 , \37482 , \37483 , \37484 , \37485 , \37486 ,
         \37487 , \37488 , \37489 , \37490 , \37491 , \37492 , \37493 , \37494 , \37495 , \37496 ,
         \37497 , \37498 , \37499 , \37500 , \37501 , \37502 , \37503 , \37504 , \37505 , \37506 ,
         \37507 , \37508 , \37509 , \37510 , \37511 , \37512 , \37513 , \37514 , \37515 , \37516 ,
         \37517 , \37518 , \37519 , \37520 , \37521 , \37522 , \37523 , \37524 , \37525 , \37526 ,
         \37527 , \37528 , \37529 , \37530 , \37531 , \37532 , \37533 , \37534 , \37535 , \37536 ,
         \37537 , \37538 , \37539 , \37540 , \37541 , \37542 , \37543 , \37544 , \37545 , \37546 ,
         \37547 , \37548 , \37549 , \37550 , \37551 , \37552 , \37553 , \37554 , \37555 , \37556 ,
         \37557 , \37558 , \37559 , \37560 , \37561 , \37562 , \37563 , \37564 , \37565 , \37566 ,
         \37567 , \37568 , \37569 , \37570 , \37571 , \37572 , \37573 , \37574 , \37575 , \37576 ,
         \37577 , \37578 , \37579 , \37580 , \37581 , \37582 , \37583 , \37584 , \37585 , \37586 ,
         \37587 , \37588 , \37589 , \37590 , \37591 , \37592 , \37593 , \37594 , \37595 , \37596 ,
         \37597 , \37598 , \37599 , \37600 , \37601 , \37602 , \37603 , \37604 , \37605 , \37606 ,
         \37607 , \37608 , \37609 , \37610 , \37611 , \37612 , \37613 , \37614 , \37615 , \37616 ,
         \37617 , \37618 , \37619 , \37620 , \37621 , \37622 , \37623 , \37624 , \37625 , \37626 ,
         \37627 , \37628 , \37629 , \37630 , \37631 , \37632 , \37633 , \37634 , \37635 , \37636 ,
         \37637 , \37638 , \37639 , \37640 , \37641 , \37642 , \37643 , \37644 , \37645 , \37646 ,
         \37647 , \37648 , \37649 , \37650 , \37651 , \37652 , \37653 , \37654 , \37655 , \37656 ,
         \37657 , \37658 , \37659 , \37660 , \37661 , \37662 , \37663 , \37664 , \37665 , \37666 ,
         \37667 , \37668 , \37669 , \37670 , \37671 , \37672 , \37673 , \37674 , \37675 , \37676 ,
         \37677 , \37678 , \37679 , \37680 , \37681 , \37682 , \37683 , \37684 , \37685 , \37686 ,
         \37687 , \37688 , \37689 , \37690 , \37691 , \37692 , \37693 , \37694 , \37695 , \37696 ,
         \37697 , \37698 , \37699 , \37700 , \37701 , \37702 , \37703 , \37704 , \37705 , \37706 ,
         \37707 , \37708 , \37709 , \37710 , \37711 , \37712 , \37713 , \37714 , \37715 , \37716 ,
         \37717 , \37718 , \37719 , \37720 , \37721 , \37722 , \37723 , \37724 , \37725 , \37726 ,
         \37727 , \37728 , \37729 , \37730 , \37731 , \37732 , \37733 , \37734 , \37735 , \37736 ,
         \37737 , \37738 , \37739 , \37740 , \37741 , \37742 , \37743 , \37744 , \37745 , \37746 ,
         \37747 , \37748 , \37749 , \37750 , \37751 , \37752 , \37753 , \37754 , \37755 , \37756 ,
         \37757 , \37758 , \37759 , \37760 , \37761 , \37762 , \37763 , \37764 , \37765 , \37766 ,
         \37767 , \37768 , \37769 , \37770 , \37771 , \37772 , \37773 , \37774 , \37775 , \37776 ,
         \37777 , \37778 , \37779 , \37780 , \37781 , \37782 , \37783 , \37784 , \37785 , \37786 ,
         \37787 , \37788 , \37789 , \37790 , \37791 , \37792 , \37793 , \37794 , \37795 , \37796 ,
         \37797 , \37798 , \37799 , \37800 , \37801 , \37802 , \37803 , \37804 , \37805 , \37806 ,
         \37807 , \37808 , \37809 , \37810 , \37811 , \37812 , \37813 , \37814 , \37815 , \37816 ,
         \37817 , \37818 , \37819 , \37820 , \37821 , \37822 , \37823 , \37824 , \37825 , \37826 ,
         \37827 , \37828 , \37829 , \37830 , \37831 , \37832 , \37833 , \37834 , \37835 , \37836 ,
         \37837 , \37838 , \37839 , \37840 , \37841 , \37842 , \37843 , \37844 , \37845 , \37846 ,
         \37847 , \37848 , \37849 , \37850 , \37851 , \37852 , \37853 , \37854 , \37855 , \37856 ,
         \37857 , \37858 , \37859 , \37860 , \37861 , \37862 , \37863 , \37864 , \37865 , \37866 ,
         \37867 , \37868 , \37869 , \37870 , \37871 , \37872 , \37873 , \37874 , \37875 , \37876 ,
         \37877 , \37878 , \37879 , \37880 , \37881 , \37882 , \37883 , \37884 , \37885 , \37886 ,
         \37887 , \37888 , \37889 , \37890 , \37891 , \37892 , \37893 , \37894 , \37895 , \37896 ,
         \37897 , \37898 , \37899 , \37900 , \37901 , \37902 , \37903 , \37904 , \37905 , \37906 ,
         \37907 , \37908 , \37909 , \37910 , \37911 , \37912 , \37913 , \37914 , \37915 , \37916 ,
         \37917 , \37918 , \37919 , \37920 , \37921 , \37922 , \37923 , \37924 , \37925 , \37926 ,
         \37927 , \37928 , \37929 , \37930 , \37931 , \37932 , \37933 , \37934 , \37935 , \37936 ,
         \37937 , \37938 , \37939 , \37940 , \37941 , \37942 , \37943 , \37944 , \37945 , \37946 ,
         \37947 , \37948 , \37949 , \37950 , \37951 , \37952 , \37953 , \37954 , \37955 , \37956 ,
         \37957 , \37958 , \37959 , \37960 , \37961 , \37962 , \37963 , \37964 , \37965 , \37966 ,
         \37967 , \37968 , \37969 , \37970 , \37971 , \37972 , \37973 , \37974 , \37975 , \37976 ,
         \37977 , \37978 , \37979 , \37980 , \37981 , \37982 , \37983 , \37984 , \37985 , \37986 ,
         \37987 , \37988 , \37989 , \37990 , \37991 , \37992 , \37993 , \37994 , \37995 , \37996 ,
         \37997 , \37998 , \37999 , \38000 , \38001 , \38002 , \38003 , \38004 , \38005 , \38006 ,
         \38007 , \38008 , \38009 , \38010 , \38011 , \38012 , \38013 , \38014 , \38015 , \38016 ,
         \38017 , \38018 , \38019 , \38020 , \38021 , \38022 , \38023 , \38024 , \38025 , \38026 ,
         \38027 , \38028 , \38029 , \38030 , \38031 , \38032 , \38033 , \38034 , \38035 , \38036 ,
         \38037 , \38038 , \38039 , \38040 , \38041 , \38042 , \38043 , \38044 , \38045 , \38046 ,
         \38047 , \38048 , \38049 , \38050 , \38051 , \38052 , \38053 , \38054 , \38055 , \38056 ,
         \38057 , \38058 , \38059 , \38060 , \38061 , \38062 , \38063 , \38064 , \38065 , \38066 ,
         \38067 , \38068 , \38069 , \38070 , \38071 , \38072 , \38073 , \38074 , \38075 , \38076 ,
         \38077 , \38078 , \38079 , \38080 , \38081 , \38082 , \38083 , \38084 , \38085 , \38086 ,
         \38087 , \38088 , \38089 , \38090 , \38091 , \38092 , \38093 , \38094 , \38095 , \38096 ,
         \38097 , \38098 , \38099 , \38100 , \38101 , \38102 , \38103 , \38104 , \38105 , \38106 ,
         \38107 , \38108 , \38109 , \38110 , \38111 , \38112 , \38113 , \38114 , \38115 , \38116 ,
         \38117 , \38118 , \38119 , \38120 , \38121 , \38122 , \38123 , \38124 , \38125 , \38126 ,
         \38127 , \38128 , \38129 , \38130 , \38131 , \38132 , \38133 , \38134 , \38135 , \38136 ,
         \38137 , \38138 , \38139 , \38140 , \38141 , \38142 , \38143 , \38144 , \38145 , \38146 ,
         \38147 , \38148 , \38149 , \38150 , \38151 , \38152 , \38153 , \38154 , \38155 , \38156 ,
         \38157 , \38158 , \38159 , \38160 , \38161 , \38162 , \38163 , \38164 , \38165 , \38166 ,
         \38167 , \38168 , \38169 , \38170 , \38171 , \38172 , \38173 , \38174 , \38175 , \38176 ,
         \38177 , \38178 , \38179 , \38180 , \38181 , \38182 , \38183 , \38184 , \38185 , \38186 ,
         \38187 , \38188 , \38189 , \38190 , \38191 , \38192 , \38193 , \38194 , \38195 , \38196 ,
         \38197 , \38198 , \38199 , \38200 , \38201 , \38202 , \38203 , \38204 , \38205 , \38206 ,
         \38207 , \38208 , \38209 , \38210 , \38211 , \38212 , \38213 , \38214 , \38215 , \38216 ,
         \38217 , \38218 , \38219 , \38220 , \38221 , \38222 , \38223 , \38224 , \38225 , \38226 ,
         \38227 , \38228 , \38229 , \38230 , \38231 , \38232 , \38233 , \38234 , \38235 , \38236 ,
         \38237 , \38238 , \38239 , \38240 , \38241 , \38242 , \38243 , \38244 , \38245 , \38246 ,
         \38247 , \38248 , \38249 , \38250 , \38251 , \38252 , \38253 , \38254 , \38255 , \38256 ,
         \38257 , \38258 , \38259 , \38260 , \38261 , \38262 , \38263 , \38264 , \38265 , \38266 ,
         \38267 , \38268 , \38269 , \38270 , \38271 , \38272 , \38273 , \38274 , \38275 , \38276 ,
         \38277 , \38278 , \38279 , \38280 , \38281 , \38282 , \38283 , \38284 , \38285 , \38286 ,
         \38287 , \38288 , \38289 , \38290 , \38291 , \38292 , \38293 , \38294 , \38295 , \38296 ,
         \38297 , \38298 , \38299 , \38300 , \38301 , \38302 , \38303 , \38304 , \38305 , \38306 ,
         \38307 , \38308 , \38309 , \38310 , \38311 , \38312 , \38313 , \38314 , \38315 , \38316 ,
         \38317 , \38318 , \38319 , \38320 , \38321 , \38322 , \38323 , \38324 , \38325 , \38326 ,
         \38327 , \38328 , \38329 , \38330 , \38331 , \38332 , \38333 , \38334 , \38335 , \38336 ,
         \38337 , \38338 , \38339 , \38340 , \38341 , \38342 , \38343 , \38344 , \38345 , \38346 ,
         \38347 , \38348 , \38349 , \38350 , \38351 , \38352 , \38353 , \38354 , \38355 , \38356 ,
         \38357 , \38358 , \38359 , \38360 , \38361 , \38362 , \38363 , \38364 , \38365 , \38366 ,
         \38367 , \38368 , \38369 , \38370 , \38371 , \38372 , \38373 , \38374 , \38375 , \38376 ,
         \38377 , \38378 , \38379 , \38380 , \38381 , \38382 , \38383 , \38384 , \38385 , \38386 ,
         \38387 , \38388 , \38389 , \38390 , \38391 , \38392 , \38393 , \38394 , \38395 , \38396 ,
         \38397 , \38398 , \38399 , \38400 , \38401 , \38402 , \38403 , \38404 , \38405 , \38406 ,
         \38407 , \38408 , \38409 , \38410 , \38411 , \38412 , \38413 , \38414 , \38415 , \38416 ,
         \38417 , \38418 , \38419 , \38420 , \38421 , \38422 , \38423 , \38424 , \38425 , \38426 ,
         \38427 , \38428 , \38429 , \38430 , \38431 , \38432 , \38433 , \38434 , \38435 , \38436 ,
         \38437 , \38438 , \38439 , \38440 , \38441 , \38442 , \38443 , \38444 , \38445 , \38446 ,
         \38447 , \38448 , \38449 , \38450 , \38451 , \38452 , \38453 , \38454 , \38455 , \38456 ,
         \38457 , \38458 , \38459 , \38460 , \38461 , \38462 , \38463 , \38464 , \38465 , \38466 ,
         \38467 , \38468 , \38469 , \38470 , \38471 , \38472 , \38473 , \38474 , \38475 , \38476 ,
         \38477 , \38478 , \38479 , \38480 , \38481 , \38482 , \38483 , \38484 , \38485 , \38486 ,
         \38487 , \38488 , \38489 , \38490 , \38491 , \38492 , \38493 , \38494 , \38495 , \38496 ,
         \38497 , \38498 , \38499 , \38500 , \38501 , \38502 , \38503 , \38504 , \38505 , \38506 ,
         \38507 , \38508 , \38509 , \38510 , \38511 , \38512 , \38513 , \38514 , \38515 , \38516 ,
         \38517 , \38518 , \38519 , \38520 , \38521 , \38522 , \38523 , \38524 , \38525 , \38526 ,
         \38527 , \38528 , \38529 , \38530 , \38531 , \38532 , \38533 , \38534 , \38535 , \38536 ,
         \38537 , \38538 , \38539 , \38540 , \38541 , \38542 , \38543 , \38544 , \38545 , \38546 ,
         \38547 , \38548 , \38549 , \38550 , \38551 , \38552 , \38553 , \38554 , \38555 , \38556 ,
         \38557 , \38558 , \38559 , \38560 , \38561 , \38562 , \38563 , \38564 , \38565 , \38566 ,
         \38567 , \38568 , \38569 , \38570 , \38571 , \38572 , \38573 , \38574 , \38575 , \38576 ,
         \38577 , \38578 , \38579 , \38580 , \38581 , \38582 , \38583 , \38584 , \38585 , \38586 ,
         \38587 , \38588 , \38589 , \38590 , \38591 , \38592 , \38593 , \38594 , \38595 , \38596 ,
         \38597 , \38598 , \38599 , \38600 , \38601 , \38602 , \38603 , \38604 , \38605 , \38606 ,
         \38607 , \38608 , \38609 , \38610 , \38611 , \38612 , \38613 , \38614 , \38615 , \38616 ,
         \38617 , \38618 , \38619 , \38620 , \38621 , \38622 , \38623 , \38624 , \38625 , \38626 ,
         \38627 , \38628 , \38629 , \38630 , \38631 , \38632 , \38633 , \38634 , \38635 , \38636 ,
         \38637 , \38638 , \38639 , \38640 , \38641 , \38642 , \38643 , \38644 , \38645 , \38646 ,
         \38647 , \38648 , \38649 , \38650 , \38651 , \38652 , \38653 , \38654 , \38655 , \38656 ,
         \38657 , \38658 , \38659 , \38660 , \38661 , \38662 , \38663 , \38664 , \38665 , \38666 ,
         \38667 , \38668 , \38669 , \38670 , \38671 , \38672 , \38673 , \38674 , \38675 , \38676 ,
         \38677 , \38678 , \38679 , \38680 , \38681 , \38682 , \38683 , \38684 , \38685 , \38686 ,
         \38687 , \38688 , \38689 , \38690 , \38691 , \38692 , \38693 , \38694 , \38695 , \38696 ,
         \38697 , \38698 , \38699 , \38700 , \38701 , \38702 , \38703 , \38704 , \38705 , \38706 ,
         \38707 , \38708 , \38709 , \38710 , \38711 , \38712 , \38713 , \38714 , \38715 , \38716 ,
         \38717 , \38718 , \38719 , \38720 , \38721 , \38722 , \38723 , \38724 , \38725 , \38726 ,
         \38727 , \38728 , \38729 , \38730 , \38731 , \38732 , \38733 , \38734 , \38735 , \38736 ,
         \38737 , \38738 , \38739 , \38740 , \38741 , \38742 , \38743 , \38744 , \38745 , \38746 ,
         \38747 , \38748 , \38749 , \38750 , \38751 , \38752 , \38753 , \38754 , \38755 , \38756 ,
         \38757 , \38758 , \38759 , \38760 , \38761 , \38762 , \38763 , \38764 , \38765 , \38766 ,
         \38767 , \38768 , \38769 , \38770 , \38771 , \38772 , \38773 , \38774 , \38775 , \38776 ,
         \38777 , \38778 , \38779 , \38780 , \38781 , \38782 , \38783 , \38784 , \38785 , \38786 ,
         \38787 , \38788 , \38789 , \38790 , \38791 , \38792 , \38793 , \38794 , \38795 , \38796 ,
         \38797 , \38798 , \38799 , \38800 , \38801 , \38802 , \38803 , \38804 , \38805 , \38806 ,
         \38807 , \38808 , \38809 , \38810 , \38811 , \38812 , \38813 , \38814 , \38815 , \38816 ,
         \38817 , \38818 , \38819 , \38820 , \38821 , \38822 , \38823 , \38824 , \38825 , \38826 ,
         \38827 , \38828 , \38829 , \38830 , \38831 , \38832 , \38833 , \38834 , \38835 , \38836 ,
         \38837 , \38838 , \38839 , \38840 , \38841 , \38842 , \38843 , \38844 , \38845 , \38846 ,
         \38847 , \38848 , \38849 , \38850 , \38851 , \38852 , \38853 , \38854 , \38855 , \38856 ,
         \38857 , \38858 , \38859 , \38860 , \38861 , \38862 , \38863 , \38864 , \38865 , \38866 ,
         \38867 , \38868 , \38869 , \38870 , \38871 , \38872 , \38873 , \38874 , \38875 , \38876 ,
         \38877 , \38878 , \38879 , \38880 , \38881 , \38882 , \38883 , \38884 , \38885 , \38886 ,
         \38887 , \38888 , \38889 , \38890 , \38891 , \38892 , \38893 , \38894 , \38895 , \38896 ,
         \38897 , \38898 , \38899 , \38900 , \38901 , \38902 , \38903 , \38904 , \38905 , \38906 ,
         \38907 , \38908 , \38909 , \38910 , \38911 , \38912 , \38913 , \38914 , \38915 , \38916 ,
         \38917 , \38918 , \38919 , \38920 , \38921 , \38922 , \38923 , \38924 , \38925 , \38926 ,
         \38927 , \38928 , \38929 , \38930 , \38931 , \38932 , \38933 , \38934 , \38935 , \38936 ,
         \38937 , \38938 , \38939 , \38940 , \38941 , \38942 , \38943 , \38944 , \38945 , \38946 ,
         \38947 , \38948 , \38949 , \38950 , \38951 , \38952 , \38953 , \38954 , \38955 , \38956 ,
         \38957 , \38958 , \38959 , \38960 , \38961 , \38962 , \38963 , \38964 , \38965 , \38966 ,
         \38967 , \38968 , \38969 , \38970 , \38971 , \38972 , \38973 , \38974 , \38975 , \38976 ,
         \38977 , \38978 , \38979 , \38980 , \38981 , \38982 , \38983 , \38984 , \38985 , \38986 ,
         \38987 , \38988 , \38989 , \38990 , \38991 , \38992 , \38993 , \38994 , \38995 , \38996 ,
         \38997 , \38998 , \38999 , \39000 , \39001 , \39002 , \39003 , \39004 , \39005 , \39006 ,
         \39007 , \39008 , \39009 , \39010 , \39011 , \39012 , \39013 , \39014 , \39015 , \39016 ,
         \39017 , \39018 , \39019 , \39020 , \39021 , \39022 , \39023 , \39024 , \39025 , \39026 ,
         \39027 , \39028 , \39029 , \39030 , \39031 , \39032 , \39033 , \39034 , \39035 , \39036 ,
         \39037 , \39038 , \39039 , \39040 , \39041 , \39042 , \39043 , \39044 , \39045 , \39046 ,
         \39047 , \39048 , \39049 , \39050 , \39051 , \39052 , \39053 , \39054 , \39055 , \39056 ,
         \39057 , \39058 , \39059 , \39060 , \39061 , \39062 , \39063 , \39064 , \39065 , \39066 ,
         \39067 , \39068 , \39069 , \39070 , \39071 , \39072 , \39073 , \39074 , \39075 , \39076 ,
         \39077 , \39078 , \39079 , \39080 , \39081 , \39082 , \39083 , \39084 , \39085 , \39086 ,
         \39087 , \39088 , \39089 , \39090 , \39091 , \39092 , \39093 , \39094 , \39095 , \39096 ,
         \39097 , \39098 , \39099 , \39100 , \39101 , \39102 , \39103 , \39104 , \39105 , \39106 ,
         \39107 , \39108 , \39109 , \39110 , \39111 , \39112 , \39113 , \39114 , \39115 , \39116 ,
         \39117 , \39118 , \39119 , \39120 , \39121 , \39122 , \39123 , \39124 , \39125 , \39126 ,
         \39127 , \39128 , \39129 , \39130 , \39131 , \39132 , \39133 , \39134 , \39135 , \39136 ,
         \39137 , \39138 , \39139 , \39140 , \39141 , \39142 , \39143 , \39144 , \39145 , \39146 ,
         \39147 , \39148 , \39149 , \39150 , \39151 , \39152 , \39153 , \39154 , \39155 , \39156 ,
         \39157 , \39158 , \39159 , \39160 , \39161 , \39162 , \39163 , \39164 , \39165 , \39166 ,
         \39167 , \39168 , \39169 , \39170 , \39171 , \39172 , \39173 , \39174 , \39175 , \39176 ,
         \39177 , \39178 , \39179 , \39180 , \39181 , \39182 , \39183 , \39184 , \39185 , \39186 ,
         \39187 , \39188 , \39189 , \39190 , \39191 , \39192 , \39193 , \39194 , \39195 , \39196 ,
         \39197 , \39198 , \39199 , \39200 , \39201 , \39202 , \39203 , \39204 , \39205 , \39206 ,
         \39207 , \39208 , \39209 , \39210 , \39211 , \39212 , \39213 , \39214 , \39215 , \39216 ,
         \39217 , \39218 , \39219 , \39220 , \39221 , \39222 , \39223 , \39224 , \39225 , \39226 ,
         \39227 , \39228 , \39229 , \39230 , \39231 , \39232 , \39233 , \39234 , \39235 , \39236 ,
         \39237 , \39238 , \39239 , \39240 , \39241 , \39242 , \39243 , \39244 , \39245 , \39246 ,
         \39247 , \39248 , \39249 , \39250 , \39251 , \39252 , \39253 , \39254 , \39255 , \39256 ,
         \39257 , \39258 , \39259 , \39260 , \39261 , \39262 , \39263 , \39264 , \39265 , \39266 ,
         \39267 , \39268 , \39269 , \39270 , \39271 , \39272 , \39273 , \39274 , \39275 , \39276 ,
         \39277 , \39278 , \39279 , \39280 , \39281 , \39282 , \39283 , \39284 , \39285 , \39286 ,
         \39287 , \39288 , \39289 , \39290 , \39291 , \39292 , \39293 , \39294 , \39295 , \39296 ,
         \39297 , \39298 , \39299 , \39300 , \39301 , \39302 , \39303 , \39304 , \39305 , \39306 ,
         \39307 , \39308 , \39309 , \39310 , \39311 , \39312 , \39313 , \39314 , \39315 , \39316 ,
         \39317 , \39318 , \39319 , \39320 , \39321 , \39322 , \39323 , \39324 , \39325 , \39326 ,
         \39327 , \39328 , \39329 , \39330 , \39331 , \39332 , \39333 , \39334 , \39335 , \39336 ,
         \39337 , \39338 , \39339 , \39340 , \39341 , \39342 , \39343 , \39344 , \39345 , \39346 ,
         \39347 , \39348 , \39349 , \39350 , \39351 , \39352 , \39353 , \39354 , \39355 , \39356 ,
         \39357 , \39358 , \39359 , \39360 , \39361 , \39362 , \39363 , \39364 , \39365 , \39366 ,
         \39367 , \39368 , \39369 , \39370 , \39371 , \39372 , \39373 , \39374 , \39375 , \39376 ,
         \39377 , \39378 , \39379 , \39380 , \39381 , \39382 , \39383 , \39384 , \39385 , \39386 ,
         \39387 , \39388 , \39389 , \39390 , \39391 , \39392 , \39393 , \39394 , \39395 , \39396 ,
         \39397 , \39398 , \39399 , \39400 , \39401 , \39402 , \39403 , \39404 , \39405 , \39406 ,
         \39407 , \39408 , \39409 , \39410 , \39411 , \39412 , \39413 , \39414 , \39415 , \39416 ,
         \39417 , \39418 , \39419 , \39420 , \39421 , \39422 , \39423 , \39424 , \39425 , \39426 ,
         \39427 , \39428 , \39429 , \39430 , \39431 , \39432 , \39433 , \39434 , \39435 , \39436 ,
         \39437 , \39438 , \39439 , \39440 , \39441 , \39442 , \39443 , \39444 , \39445 , \39446 ,
         \39447 , \39448 , \39449 , \39450 , \39451 , \39452 , \39453 , \39454 , \39455 , \39456 ,
         \39457 , \39458 , \39459 , \39460 , \39461 , \39462 , \39463 , \39464 , \39465 , \39466 ,
         \39467 , \39468 , \39469 , \39470 , \39471 , \39472 , \39473 , \39474 , \39475 , \39476 ,
         \39477 , \39478 , \39479 , \39480 , \39481 , \39482 , \39483 , \39484 , \39485 , \39486 ,
         \39487 , \39488 , \39489 , \39490 , \39491 , \39492 , \39493 , \39494 , \39495 , \39496 ,
         \39497 , \39498 , \39499 , \39500 , \39501 , \39502 , \39503 , \39504 , \39505 , \39506 ,
         \39507 , \39508 , \39509 , \39510 , \39511 , \39512 , \39513 , \39514 , \39515 , \39516 ,
         \39517 , \39518 , \39519 , \39520 , \39521 , \39522 , \39523 , \39524 , \39525 , \39526 ,
         \39527 , \39528 , \39529 , \39530 , \39531 , \39532 , \39533 , \39534 , \39535 , \39536 ,
         \39537 , \39538 , \39539 , \39540 , \39541 , \39542 , \39543 , \39544 , \39545 , \39546 ,
         \39547 , \39548 , \39549 , \39550 , \39551 , \39552 , \39553 , \39554 , \39555 , \39556 ,
         \39557 , \39558 , \39559 , \39560 , \39561 , \39562 , \39563 , \39564 , \39565 , \39566 ,
         \39567 , \39568 , \39569 , \39570 , \39571 , \39572 , \39573 , \39574 , \39575 , \39576 ,
         \39577 , \39578 , \39579 , \39580 , \39581 , \39582 , \39583 , \39584 , \39585 , \39586 ,
         \39587 , \39588 , \39589 , \39590 , \39591 , \39592 , \39593 , \39594 , \39595 , \39596 ,
         \39597 , \39598 , \39599 , \39600 , \39601 , \39602 , \39603 , \39604 , \39605 , \39606 ,
         \39607 , \39608 , \39609 , \39610 , \39611 , \39612 , \39613 , \39614 , \39615 , \39616 ,
         \39617 , \39618 , \39619 , \39620 , \39621 , \39622 , \39623 , \39624 , \39625 , \39626 ,
         \39627 , \39628 , \39629 , \39630 , \39631 , \39632 , \39633 , \39634 , \39635 , \39636 ,
         \39637 , \39638 , \39639 , \39640 , \39641 , \39642 , \39643 , \39644 , \39645 , \39646 ,
         \39647 , \39648 , \39649 , \39650 , \39651 , \39652 , \39653 , \39654 , \39655 , \39656 ,
         \39657 , \39658 , \39659 , \39660 , \39661 , \39662 , \39663 , \39664 , \39665 , \39666 ,
         \39667 , \39668 , \39669 , \39670 , \39671 , \39672 , \39673 , \39674 , \39675 , \39676 ,
         \39677 , \39678 , \39679 , \39680 , \39681 , \39682 , \39683 , \39684 , \39685 , \39686 ,
         \39687 , \39688 , \39689 , \39690 , \39691 , \39692 , \39693 , \39694 , \39695 , \39696 ,
         \39697 , \39698 , \39699 , \39700 , \39701 , \39702 , \39703 , \39704 , \39705 , \39706 ,
         \39707 , \39708 , \39709 , \39710 , \39711 , \39712 , \39713 , \39714 , \39715 , \39716 ,
         \39717 , \39718 , \39719 , \39720 , \39721 , \39722 , \39723 , \39724 , \39725 , \39726 ,
         \39727 , \39728 , \39729 , \39730 , \39731 , \39732 , \39733 , \39734 , \39735 , \39736 ,
         \39737 , \39738 , \39739 , \39740 , \39741 , \39742 , \39743 , \39744 , \39745 , \39746 ,
         \39747 , \39748 , \39749 , \39750 , \39751 , \39752 , \39753 , \39754 , \39755 , \39756 ,
         \39757 , \39758 , \39759 , \39760 , \39761 , \39762 , \39763 , \39764 , \39765 , \39766 ,
         \39767 , \39768 , \39769 , \39770 , \39771 , \39772 , \39773 , \39774 , \39775 , \39776 ,
         \39777 , \39778 , \39779 , \39780 , \39781 , \39782 , \39783 , \39784 , \39785 , \39786 ,
         \39787 , \39788 , \39789 , \39790 , \39791 , \39792 , \39793 , \39794 , \39795 , \39796 ,
         \39797 , \39798 , \39799 , \39800 , \39801 , \39802 , \39803 , \39804 , \39805 , \39806 ,
         \39807 , \39808 , \39809 , \39810 , \39811 , \39812 , \39813 , \39814 , \39815 , \39816 ,
         \39817 , \39818 , \39819 , \39820 , \39821 , \39822 , \39823 , \39824 , \39825 , \39826 ,
         \39827 , \39828 , \39829 , \39830 , \39831 , \39832 , \39833 , \39834 , \39835 , \39836 ,
         \39837 , \39838 , \39839 , \39840 , \39841 , \39842 , \39843 , \39844 , \39845 , \39846 ,
         \39847 , \39848 , \39849 , \39850 , \39851 , \39852 , \39853 , \39854 , \39855 , \39856 ,
         \39857 , \39858 , \39859 , \39860 , \39861 , \39862 , \39863 , \39864 , \39865 , \39866 ,
         \39867 , \39868 , \39869 , \39870 , \39871 , \39872 , \39873 , \39874 , \39875 , \39876 ,
         \39877 , \39878 , \39879 , \39880 , \39881 , \39882 , \39883 , \39884 , \39885 , \39886 ,
         \39887 , \39888 , \39889 , \39890 , \39891 , \39892 , \39893 , \39894 , \39895 , \39896 ,
         \39897 , \39898 , \39899 , \39900 , \39901 , \39902 , \39903 , \39904 , \39905 , \39906 ,
         \39907 , \39908 , \39909 , \39910 , \39911 , \39912 , \39913 , \39914 , \39915 , \39916 ,
         \39917 , \39918 , \39919 , \39920 , \39921 , \39922 , \39923 , \39924 , \39925 , \39926 ,
         \39927 , \39928 , \39929 , \39930 , \39931 , \39932 , \39933 , \39934 , \39935 , \39936 ,
         \39937 , \39938 , \39939 , \39940 , \39941 , \39942 , \39943 , \39944 , \39945 , \39946 ,
         \39947 , \39948 , \39949 , \39950 , \39951 , \39952 , \39953 , \39954 , \39955 , \39956 ,
         \39957 , \39958 , \39959 , \39960 , \39961 , \39962 , \39963 , \39964 , \39965 , \39966 ,
         \39967 , \39968 , \39969 , \39970 , \39971 , \39972 , \39973 , \39974 , \39975 , \39976 ,
         \39977 , \39978 , \39979 , \39980 , \39981 , \39982 , \39983 , \39984 , \39985 , \39986 ,
         \39987 , \39988 , \39989 , \39990 , \39991 , \39992 , \39993 , \39994 , \39995 , \39996 ,
         \39997 , \39998 , \39999 , \40000 , \40001 , \40002 , \40003 , \40004 , \40005 , \40006 ,
         \40007 , \40008 , \40009 , \40010 , \40011 , \40012 , \40013 , \40014 , \40015 , \40016 ,
         \40017 , \40018 , \40019 , \40020 , \40021 , \40022 , \40023 , \40024 , \40025 , \40026 ,
         \40027 , \40028 , \40029 , \40030 , \40031 , \40032 , \40033 , \40034 , \40035 , \40036 ,
         \40037 , \40038 , \40039 , \40040 , \40041 , \40042 , \40043 , \40044 , \40045 , \40046 ,
         \40047 , \40048 , \40049 , \40050 , \40051 , \40052 , \40053 , \40054 , \40055 , \40056 ,
         \40057 , \40058 , \40059 , \40060 , \40061 , \40062 , \40063 , \40064 , \40065 , \40066 ,
         \40067 , \40068 , \40069 , \40070 , \40071 , \40072 , \40073 , \40074 , \40075 , \40076 ,
         \40077 , \40078 , \40079 , \40080 , \40081 , \40082 , \40083 , \40084 , \40085 , \40086 ,
         \40087 , \40088 , \40089 , \40090 , \40091 , \40092 , \40093 , \40094 , \40095 , \40096 ,
         \40097 , \40098 , \40099 , \40100 , \40101 , \40102 , \40103 , \40104 , \40105 , \40106 ,
         \40107 , \40108 , \40109 , \40110 , \40111 , \40112 , \40113 , \40114 , \40115 , \40116 ,
         \40117 , \40118 , \40119 , \40120 , \40121 , \40122 , \40123 , \40124 , \40125 , \40126 ,
         \40127 , \40128 , \40129 , \40130 , \40131 , \40132 , \40133 , \40134 , \40135 , \40136 ,
         \40137 , \40138 , \40139 , \40140 , \40141 , \40142 , \40143 , \40144 , \40145 , \40146 ,
         \40147 , \40148 , \40149 , \40150 , \40151 , \40152 , \40153 , \40154 , \40155 , \40156 ,
         \40157 , \40158 , \40159 , \40160 , \40161 , \40162 , \40163 , \40164 , \40165 , \40166 ,
         \40167 , \40168 , \40169 , \40170 , \40171 , \40172 , \40173 , \40174 , \40175 , \40176 ,
         \40177 , \40178 , \40179 , \40180 , \40181 , \40182 , \40183 , \40184 , \40185 , \40186 ,
         \40187 , \40188 , \40189 , \40190 , \40191 , \40192 , \40193 , \40194 , \40195 , \40196 ,
         \40197 , \40198 , \40199 , \40200 , \40201 , \40202 , \40203 , \40204 , \40205 , \40206 ,
         \40207 , \40208 , \40209 , \40210 , \40211 , \40212 , \40213 , \40214 , \40215 , \40216 ,
         \40217 , \40218 , \40219 , \40220 , \40221 , \40222 , \40223 , \40224 , \40225 , \40226 ,
         \40227 , \40228 , \40229 , \40230 , \40231 , \40232 , \40233 , \40234 , \40235 , \40236 ,
         \40237 , \40238 , \40239 , \40240 , \40241 , \40242 , \40243 , \40244 , \40245 , \40246 ,
         \40247 , \40248 , \40249 , \40250 , \40251 , \40252 , \40253 , \40254 , \40255 , \40256 ,
         \40257 , \40258 , \40259 , \40260 , \40261 , \40262 , \40263 , \40264 , \40265 , \40266 ,
         \40267 , \40268 , \40269 , \40270 , \40271 , \40272 , \40273 , \40274 , \40275 , \40276 ,
         \40277 , \40278 , \40279 , \40280 , \40281 , \40282 , \40283 , \40284 , \40285 , \40286 ,
         \40287 , \40288 , \40289 , \40290 , \40291 , \40292 , \40293 , \40294 , \40295 , \40296 ,
         \40297 , \40298 , \40299 , \40300 , \40301 , \40302 , \40303 , \40304 , \40305 , \40306 ,
         \40307 , \40308 , \40309 , \40310 , \40311 , \40312 , \40313 , \40314 , \40315 , \40316 ,
         \40317 , \40318 , \40319 , \40320 , \40321 , \40322 , \40323 , \40324 , \40325 , \40326 ,
         \40327 , \40328 , \40329 , \40330 , \40331 , \40332 , \40333 , \40334 , \40335 , \40336 ,
         \40337 , \40338 , \40339 , \40340 , \40341 , \40342 , \40343 , \40344 , \40345 , \40346 ,
         \40347 , \40348 , \40349 , \40350 , \40351 , \40352 , \40353 , \40354 , \40355 , \40356 ,
         \40357 , \40358 , \40359 , \40360 , \40361 , \40362 , \40363 , \40364 , \40365 , \40366 ,
         \40367 , \40368 , \40369 , \40370 , \40371 , \40372 , \40373 , \40374 , \40375 , \40376 ,
         \40377 , \40378 , \40379 , \40380 , \40381 , \40382 , \40383 , \40384 , \40385 , \40386 ,
         \40387 , \40388 , \40389 , \40390 , \40391 , \40392 , \40393 , \40394 , \40395 , \40396 ,
         \40397 , \40398 , \40399 , \40400 , \40401 , \40402 , \40403 , \40404 , \40405 , \40406 ,
         \40407 , \40408 , \40409 , \40410 , \40411 , \40412 , \40413 , \40414 , \40415 , \40416 ,
         \40417 , \40418 , \40419 , \40420 , \40421 , \40422 , \40423 , \40424 , \40425 , \40426 ,
         \40427 , \40428 , \40429 , \40430 , \40431 , \40432 , \40433 , \40434 , \40435 , \40436 ,
         \40437 , \40438 , \40439 , \40440 , \40441 , \40442 , \40443 , \40444 , \40445 , \40446 ,
         \40447 , \40448 , \40449 , \40450 , \40451 , \40452 , \40453 , \40454 , \40455 , \40456 ,
         \40457 , \40458 , \40459 , \40460 , \40461 , \40462 , \40463 , \40464 , \40465 , \40466 ,
         \40467 , \40468 , \40469 , \40470 , \40471 , \40472 , \40473 , \40474 , \40475 , \40476 ,
         \40477 , \40478 , \40479 , \40480 , \40481 , \40482 , \40483 , \40484 , \40485 , \40486 ,
         \40487 , \40488 , \40489 , \40490 , \40491 , \40492 , \40493 , \40494 , \40495 , \40496 ,
         \40497 , \40498 , \40499 , \40500 , \40501 , \40502 , \40503 , \40504 , \40505 , \40506 ,
         \40507 , \40508 , \40509 , \40510 , \40511 , \40512 , \40513 , \40514 , \40515 , \40516 ,
         \40517 , \40518 , \40519 , \40520 , \40521 , \40522 , \40523 , \40524 , \40525 , \40526 ,
         \40527 , \40528 , \40529 , \40530 , \40531 , \40532 , \40533 , \40534 , \40535 , \40536 ,
         \40537 , \40538 , \40539 , \40540 , \40541 , \40542 , \40543 , \40544 , \40545 , \40546 ,
         \40547 , \40548 , \40549 , \40550 , \40551 , \40552 , \40553 , \40554 , \40555 , \40556 ,
         \40557 , \40558 , \40559 , \40560 , \40561 , \40562 , \40563 , \40564 , \40565 , \40566 ,
         \40567 , \40568 , \40569 , \40570 , \40571 , \40572 , \40573 , \40574 , \40575 , \40576 ,
         \40577 , \40578 , \40579 , \40580 , \40581 , \40582 , \40583 , \40584 , \40585 , \40586 ,
         \40587 , \40588 , \40589 , \40590 , \40591 , \40592 , \40593 , \40594 , \40595 , \40596 ,
         \40597 , \40598 , \40599 , \40600 , \40601 , \40602 , \40603 , \40604 , \40605 , \40606 ,
         \40607 , \40608 , \40609 , \40610 , \40611 , \40612 , \40613 , \40614 , \40615 , \40616 ,
         \40617 , \40618 , \40619 , \40620 , \40621 , \40622 , \40623 , \40624 , \40625 , \40626 ,
         \40627 , \40628 , \40629 , \40630 , \40631 , \40632 , \40633 , \40634 , \40635 , \40636 ,
         \40637 , \40638 , \40639 , \40640 , \40641 , \40642 , \40643 , \40644 , \40645 , \40646 ,
         \40647 , \40648 , \40649 , \40650 , \40651 , \40652 , \40653 , \40654 , \40655 , \40656 ,
         \40657 , \40658 , \40659 , \40660 , \40661 , \40662 , \40663 , \40664 , \40665 , \40666 ,
         \40667 , \40668 , \40669 , \40670 , \40671 , \40672 , \40673 , \40674 , \40675 , \40676 ,
         \40677 , \40678 , \40679 , \40680 , \40681 , \40682 , \40683 , \40684 , \40685 , \40686 ,
         \40687 , \40688 , \40689 , \40690 , \40691 , \40692 , \40693 , \40694 , \40695 , \40696 ,
         \40697 , \40698 , \40699 , \40700 , \40701 , \40702 , \40703 , \40704 , \40705 , \40706 ,
         \40707 , \40708 , \40709 , \40710 , \40711 , \40712 , \40713 , \40714 , \40715 , \40716 ,
         \40717 , \40718 , \40719 , \40720 , \40721 , \40722 , \40723 , \40724 , \40725 , \40726 ,
         \40727 , \40728 , \40729 , \40730 , \40731 , \40732 , \40733 , \40734 , \40735 , \40736 ,
         \40737 , \40738 , \40739 , \40740 , \40741 , \40742 , \40743 , \40744 , \40745 , \40746 ,
         \40747 , \40748 , \40749 , \40750 , \40751 , \40752 , \40753 , \40754 , \40755 , \40756 ,
         \40757 , \40758 , \40759 , \40760 , \40761 , \40762 , \40763 , \40764 , \40765 , \40766 ,
         \40767 , \40768 , \40769 , \40770 , \40771 , \40772 , \40773 , \40774 , \40775 , \40776 ,
         \40777 , \40778 , \40779 , \40780 , \40781 , \40782 , \40783 , \40784 , \40785 , \40786 ,
         \40787 , \40788 , \40789 , \40790 , \40791 , \40792 , \40793 , \40794 , \40795 , \40796 ,
         \40797 , \40798 , \40799 , \40800 , \40801 , \40802 , \40803 , \40804 , \40805 , \40806 ,
         \40807 , \40808 , \40809 , \40810 , \40811 , \40812 , \40813 , \40814 , \40815 , \40816 ,
         \40817 , \40818 , \40819 , \40820 , \40821 , \40822 , \40823 , \40824 , \40825 , \40826 ,
         \40827 , \40828 , \40829 , \40830 , \40831 , \40832 , \40833 , \40834 , \40835 , \40836 ,
         \40837 , \40838 , \40839 , \40840 , \40841 , \40842 , \40843 , \40844 , \40845 , \40846 ,
         \40847 , \40848 , \40849 , \40850 , \40851 , \40852 , \40853 , \40854 , \40855 , \40856 ,
         \40857 , \40858 , \40859 , \40860 , \40861 , \40862 , \40863 , \40864 , \40865 , \40866 ,
         \40867 , \40868 , \40869 , \40870 , \40871 , \40872 , \40873 , \40874 , \40875 , \40876 ,
         \40877 , \40878 , \40879 , \40880 , \40881 , \40882 , \40883 , \40884 , \40885 , \40886 ,
         \40887 , \40888 , \40889 , \40890 , \40891 , \40892 , \40893 , \40894 , \40895 , \40896 ,
         \40897 , \40898 , \40899 , \40900 , \40901 , \40902 , \40903 , \40904 , \40905 , \40906 ,
         \40907 , \40908 , \40909 , \40910 , \40911 , \40912 , \40913 , \40914 , \40915 , \40916 ,
         \40917 , \40918 , \40919 , \40920 , \40921 , \40922 , \40923 , \40924 , \40925 , \40926 ,
         \40927 , \40928 , \40929 , \40930 , \40931 , \40932 , \40933 , \40934 , \40935 , \40936 ,
         \40937 , \40938 , \40939 , \40940 , \40941 , \40942 , \40943 , \40944 , \40945 , \40946 ,
         \40947 , \40948 , \40949 , \40950 , \40951 , \40952 , \40953 , \40954 , \40955 , \40956 ,
         \40957 , \40958 , \40959 , \40960 , \40961 , \40962 , \40963 , \40964 , \40965 , \40966 ,
         \40967 , \40968 , \40969 , \40970 , \40971 , \40972 , \40973 , \40974 , \40975 , \40976 ,
         \40977 , \40978 , \40979 , \40980 , \40981 , \40982 , \40983 , \40984 , \40985 , \40986 ,
         \40987 , \40988 , \40989 , \40990 , \40991 , \40992 , \40993 , \40994 , \40995 , \40996 ,
         \40997 , \40998 , \40999 , \41000 , \41001 , \41002 , \41003 , \41004 , \41005 , \41006 ,
         \41007 , \41008 , \41009 , \41010 , \41011 , \41012 , \41013 , \41014 , \41015 , \41016 ,
         \41017 , \41018 , \41019 , \41020 , \41021 , \41022 , \41023 , \41024 , \41025 , \41026 ,
         \41027 , \41028 , \41029 , \41030 , \41031 , \41032 , \41033 , \41034 , \41035 , \41036 ,
         \41037 , \41038 , \41039 , \41040 , \41041 , \41042 , \41043 , \41044 , \41045 , \41046 ,
         \41047 , \41048 , \41049 , \41050 , \41051 , \41052 , \41053 , \41054 , \41055 , \41056 ,
         \41057 , \41058 , \41059 , \41060 , \41061 , \41062 , \41063 , \41064 , \41065 , \41066 ,
         \41067 , \41068 , \41069 , \41070 , \41071 , \41072 , \41073 , \41074 , \41075 , \41076 ,
         \41077 , \41078 , \41079 , \41080 , \41081 , \41082 , \41083 , \41084 , \41085 , \41086 ,
         \41087 , \41088 , \41089 , \41090 , \41091 , \41092 , \41093 , \41094 , \41095 , \41096 ,
         \41097 , \41098 , \41099 , \41100 , \41101 , \41102 , \41103 , \41104 , \41105 , \41106 ,
         \41107 , \41108 , \41109 , \41110 , \41111 , \41112 , \41113 , \41114 , \41115 , \41116 ,
         \41117 , \41118 , \41119 , \41120 , \41121 , \41122 , \41123 , \41124 , \41125 , \41126 ,
         \41127 , \41128 , \41129 , \41130 , \41131 , \41132 , \41133 , \41134 , \41135 , \41136 ,
         \41137 , \41138 , \41139 , \41140 , \41141 , \41142 , \41143 , \41144 , \41145 , \41146 ,
         \41147 , \41148 , \41149 , \41150 , \41151 , \41152 , \41153 , \41154 , \41155 , \41156 ,
         \41157 , \41158 , \41159 , \41160 , \41161 , \41162 , \41163 , \41164 , \41165 , \41166 ,
         \41167 , \41168 , \41169 , \41170 , \41171 , \41172 , \41173 , \41174 , \41175 , \41176 ,
         \41177 , \41178 , \41179 , \41180 , \41181 , \41182 , \41183 , \41184 , \41185 , \41186 ,
         \41187 , \41188 , \41189 , \41190 , \41191 , \41192 , \41193 , \41194 , \41195 , \41196 ,
         \41197 , \41198 , \41199 , \41200 , \41201 , \41202 , \41203 , \41204 , \41205 , \41206 ,
         \41207 , \41208 , \41209 , \41210 , \41211 , \41212 , \41213 , \41214 , \41215 , \41216 ,
         \41217 , \41218 , \41219 , \41220 , \41221 , \41222 , \41223 , \41224 , \41225 , \41226 ,
         \41227 , \41228 , \41229 , \41230 , \41231 , \41232 , \41233 , \41234 , \41235 , \41236 ,
         \41237 , \41238 , \41239 , \41240 , \41241 , \41242 , \41243 , \41244 , \41245 , \41246 ,
         \41247 , \41248 , \41249 , \41250 , \41251 , \41252 , \41253 , \41254 , \41255 , \41256 ,
         \41257 , \41258 , \41259 , \41260 , \41261 , \41262 , \41263 , \41264 , \41265 , \41266 ,
         \41267 , \41268 , \41269 , \41270 , \41271 , \41272 , \41273 , \41274 , \41275 , \41276 ,
         \41277 , \41278 , \41279 , \41280 , \41281 , \41282 , \41283 , \41284 , \41285 , \41286 ,
         \41287 , \41288 , \41289 , \41290 , \41291 , \41292 , \41293 , \41294 , \41295 , \41296 ,
         \41297 , \41298 , \41299 , \41300 , \41301 , \41302 , \41303 , \41304 , \41305 , \41306 ,
         \41307 , \41308 , \41309 , \41310 , \41311 , \41312 , \41313 , \41314 , \41315 , \41316 ,
         \41317 , \41318 , \41319 , \41320 , \41321 , \41322 , \41323 , \41324 , \41325 , \41326 ,
         \41327 , \41328 , \41329 , \41330 , \41331 , \41332 , \41333 , \41334 , \41335 , \41336 ,
         \41337 , \41338 , \41339 , \41340 , \41341 , \41342 , \41343 , \41344 , \41345 , \41346 ,
         \41347 , \41348 , \41349 , \41350 , \41351 , \41352 , \41353 , \41354 , \41355 , \41356 ,
         \41357 , \41358 , \41359 , \41360 , \41361 , \41362 , \41363 , \41364 , \41365 , \41366 ,
         \41367 , \41368 , \41369 , \41370 , \41371 , \41372 , \41373 , \41374 , \41375 , \41376 ,
         \41377 , \41378 , \41379 , \41380 , \41381 , \41382 , \41383 , \41384 , \41385 , \41386 ,
         \41387 , \41388 , \41389 , \41390 , \41391 , \41392 , \41393 , \41394 , \41395 , \41396 ,
         \41397 , \41398 , \41399 , \41400 , \41401 , \41402 , \41403 , \41404 , \41405 , \41406 ,
         \41407 , \41408 , \41409 , \41410 , \41411 , \41412 , \41413 , \41414 , \41415 , \41416 ,
         \41417 , \41418 , \41419 , \41420 , \41421 , \41422 , \41423 , \41424 , \41425 , \41426 ,
         \41427 , \41428 , \41429 , \41430 , \41431 , \41432 , \41433 , \41434 , \41435 , \41436 ,
         \41437 , \41438 , \41439 , \41440 , \41441 , \41442 , \41443 , \41444 , \41445 , \41446 ,
         \41447 , \41448 , \41449 , \41450 , \41451 , \41452 , \41453 , \41454 , \41455 , \41456 ,
         \41457 , \41458 , \41459 , \41460 , \41461 , \41462 , \41463 , \41464 , \41465 , \41466 ,
         \41467 , \41468 , \41469 , \41470 , \41471 , \41472 , \41473 , \41474 , \41475 , \41476 ,
         \41477 , \41478 , \41479 , \41480 , \41481 , \41482 , \41483 , \41484 , \41485 , \41486 ,
         \41487 , \41488 , \41489 , \41490 , \41491 , \41492 , \41493 , \41494 , \41495 , \41496 ,
         \41497 , \41498 , \41499 , \41500 , \41501 , \41502 , \41503 , \41504 , \41505 , \41506 ,
         \41507 , \41508 , \41509 , \41510 , \41511 , \41512 , \41513 , \41514 , \41515 , \41516 ,
         \41517 , \41518 , \41519 , \41520 , \41521 , \41522 , \41523 , \41524 , \41525 , \41526 ,
         \41527 , \41528 , \41529 , \41530 , \41531 , \41532 , \41533 , \41534 , \41535 , \41536 ,
         \41537 , \41538 , \41539 , \41540 , \41541 , \41542 , \41543 , \41544 , \41545 , \41546 ,
         \41547 , \41548 , \41549 , \41550 , \41551 , \41552 , \41553 , \41554 , \41555 , \41556 ,
         \41557 , \41558 , \41559 , \41560 , \41561 , \41562 , \41563 , \41564 , \41565 , \41566 ,
         \41567 , \41568 , \41569 , \41570 , \41571 , \41572 , \41573 , \41574 , \41575 , \41576 ,
         \41577 , \41578 , \41579 , \41580 , \41581 , \41582 , \41583 , \41584 , \41585 , \41586 ,
         \41587 , \41588 , \41589 , \41590 , \41591 , \41592 , \41593 , \41594 , \41595 , \41596 ,
         \41597 , \41598 , \41599 , \41600 , \41601 , \41602 , \41603 , \41604 , \41605 , \41606 ,
         \41607 , \41608 , \41609 , \41610 , \41611 , \41612 , \41613 , \41614 , \41615 , \41616 ,
         \41617 , \41618 , \41619 , \41620 , \41621 , \41622 , \41623 , \41624 , \41625 , \41626 ,
         \41627 , \41628 , \41629 , \41630 , \41631 , \41632 , \41633 , \41634 , \41635 , \41636 ,
         \41637 , \41638 , \41639 , \41640 , \41641 , \41642 , \41643 , \41644 , \41645 , \41646 ,
         \41647 , \41648 , \41649 , \41650 , \41651 , \41652 , \41653 , \41654 , \41655 , \41656 ,
         \41657 , \41658 , \41659 , \41660 , \41661 , \41662 , \41663 , \41664 , \41665 , \41666 ,
         \41667 , \41668 , \41669 , \41670 , \41671 , \41672 , \41673 , \41674 , \41675 , \41676 ,
         \41677 , \41678 , \41679 , \41680 , \41681 , \41682 , \41683 , \41684 , \41685 , \41686 ,
         \41687 , \41688 , \41689 , \41690 , \41691 , \41692 , \41693 , \41694 , \41695 , \41696 ,
         \41697 , \41698 , \41699 , \41700 , \41701 , \41702 , \41703 , \41704 , \41705 , \41706 ,
         \41707 , \41708 , \41709 , \41710 , \41711 , \41712 , \41713 , \41714 , \41715 , \41716 ,
         \41717 , \41718 , \41719 , \41720 , \41721 , \41722 , \41723 , \41724 , \41725 , \41726 ,
         \41727 , \41728 , \41729 , \41730 , \41731 , \41732 , \41733 , \41734 , \41735 , \41736 ,
         \41737 , \41738 , \41739 , \41740 , \41741 , \41742 , \41743 , \41744 , \41745 , \41746 ,
         \41747 , \41748 , \41749 , \41750 , \41751 , \41752 , \41753 , \41754 , \41755 , \41756 ,
         \41757 , \41758 , \41759 , \41760 , \41761 , \41762 , \41763 , \41764 , \41765 , \41766 ,
         \41767 , \41768 , \41769 , \41770 , \41771 , \41772 , \41773 , \41774 , \41775 , \41776 ,
         \41777 , \41778 , \41779 , \41780 , \41781 , \41782 , \41783 , \41784 , \41785 , \41786 ,
         \41787 , \41788 , \41789 , \41790 , \41791 , \41792 , \41793 , \41794 , \41795 , \41796 ,
         \41797 , \41798 , \41799 , \41800 , \41801 , \41802 , \41803 , \41804 , \41805 , \41806 ,
         \41807 , \41808 , \41809 , \41810 , \41811 , \41812 , \41813 , \41814 , \41815 , \41816 ,
         \41817 , \41818 , \41819 , \41820 , \41821 , \41822 , \41823 , \41824 , \41825 , \41826 ,
         \41827 , \41828 , \41829 , \41830 , \41831 , \41832 , \41833 , \41834 , \41835 , \41836 ,
         \41837 , \41838 , \41839 , \41840 , \41841 , \41842 , \41843 , \41844 , \41845 , \41846 ,
         \41847 , \41848 , \41849 , \41850 , \41851 , \41852 , \41853 , \41854 , \41855 , \41856 ,
         \41857 , \41858 , \41859 , \41860 , \41861 , \41862 , \41863 , \41864 , \41865 , \41866 ,
         \41867 , \41868 , \41869 , \41870 , \41871 , \41872 , \41873 , \41874 , \41875 , \41876 ,
         \41877 , \41878 , \41879 , \41880 , \41881 , \41882 , \41883 , \41884 , \41885 , \41886 ,
         \41887 , \41888 , \41889 , \41890 , \41891 , \41892 , \41893 , \41894 , \41895 , \41896 ,
         \41897 , \41898 , \41899 , \41900 , \41901 , \41902 , \41903 , \41904 , \41905 , \41906 ,
         \41907 , \41908 , \41909 , \41910 , \41911 , \41912 , \41913 , \41914 , \41915 , \41916 ,
         \41917 , \41918 , \41919 , \41920 , \41921 , \41922 , \41923 , \41924 , \41925 , \41926 ,
         \41927 , \41928 , \41929 , \41930 , \41931 , \41932 , \41933 , \41934 , \41935 , \41936 ,
         \41937 , \41938 , \41939 , \41940 , \41941 , \41942 , \41943 , \41944 , \41945 , \41946 ,
         \41947 , \41948 , \41949 , \41950 , \41951 , \41952 , \41953 , \41954 , \41955 , \41956 ,
         \41957 , \41958 , \41959 , \41960 , \41961 , \41962 , \41963 , \41964 , \41965 , \41966 ,
         \41967 , \41968 , \41969 , \41970 , \41971 , \41972 , \41973 , \41974 , \41975 , \41976 ,
         \41977 , \41978 , \41979 , \41980 , \41981 , \41982 , \41983 , \41984 , \41985 , \41986 ,
         \41987 , \41988 , \41989 , \41990 , \41991 , \41992 , \41993 , \41994 , \41995 , \41996 ,
         \41997 , \41998 , \41999 , \42000 , \42001 , \42002 , \42003 , \42004 , \42005 , \42006 ,
         \42007 , \42008 , \42009 , \42010 , \42011 , \42012 , \42013 , \42014 , \42015 , \42016 ,
         \42017 , \42018 , \42019 , \42020 , \42021 , \42022 , \42023 , \42024 , \42025 , \42026 ,
         \42027 , \42028 , \42029 , \42030 , \42031 , \42032 , \42033 , \42034 , \42035 , \42036 ,
         \42037 , \42038 , \42039 , \42040 , \42041 , \42042 , \42043 , \42044 , \42045 , \42046 ,
         \42047 , \42048 , \42049 , \42050 , \42051 , \42052 , \42053 , \42054 , \42055 , \42056 ,
         \42057 , \42058 , \42059 , \42060 , \42061 , \42062 , \42063 , \42064 , \42065 , \42066 ,
         \42067 , \42068 , \42069 , \42070 , \42071 , \42072 , \42073 , \42074 , \42075 , \42076 ,
         \42077 , \42078 , \42079 , \42080 , \42081 , \42082 , \42083 , \42084 , \42085 , \42086 ,
         \42087 , \42088 , \42089 , \42090 , \42091 , \42092 , \42093 , \42094 , \42095 , \42096 ,
         \42097 , \42098 , \42099 , \42100 , \42101 , \42102 , \42103 , \42104 , \42105 , \42106 ,
         \42107 , \42108 , \42109 , \42110 , \42111 , \42112 , \42113 , \42114 , \42115 , \42116 ,
         \42117 , \42118 , \42119 , \42120 , \42121 , \42122 , \42123 , \42124 , \42125 , \42126 ,
         \42127 , \42128 , \42129 , \42130 , \42131 , \42132 , \42133 , \42134 , \42135 , \42136 ,
         \42137 , \42138 , \42139 , \42140 , \42141 , \42142 , \42143 , \42144 , \42145 , \42146 ,
         \42147 , \42148 , \42149 , \42150 , \42151 , \42152 , \42153 , \42154 , \42155 , \42156 ,
         \42157 , \42158 , \42159 , \42160 , \42161 , \42162 , \42163 , \42164 , \42165 , \42166 ,
         \42167 , \42168 , \42169 , \42170 , \42171 , \42172 , \42173 , \42174 , \42175 , \42176 ,
         \42177 , \42178 , \42179 , \42180 , \42181 , \42182 , \42183 , \42184 , \42185 , \42186 ,
         \42187 , \42188 , \42189 , \42190 , \42191 , \42192 , \42193 , \42194 , \42195 , \42196 ,
         \42197 , \42198 , \42199 , \42200 , \42201 , \42202 , \42203 , \42204 , \42205 , \42206 ,
         \42207 , \42208 , \42209 , \42210 , \42211 , \42212 , \42213 , \42214 , \42215 , \42216 ,
         \42217 , \42218 , \42219 , \42220 , \42221 , \42222 , \42223 , \42224 , \42225 , \42226 ,
         \42227 , \42228 , \42229 , \42230 , \42231 , \42232 , \42233 , \42234 , \42235 , \42236 ,
         \42237 , \42238 , \42239 , \42240 , \42241 , \42242 , \42243 , \42244 , \42245 , \42246 ,
         \42247 , \42248 , \42249 , \42250 , \42251 , \42252 , \42253 , \42254 , \42255 , \42256 ,
         \42257 , \42258 , \42259 , \42260 , \42261 , \42262 , \42263 , \42264 , \42265 , \42266 ,
         \42267 , \42268 , \42269 , \42270 , \42271 , \42272 , \42273 , \42274 , \42275 , \42276 ,
         \42277 , \42278 , \42279 , \42280 , \42281 , \42282 , \42283 , \42284 , \42285 , \42286 ,
         \42287 , \42288 , \42289 , \42290 , \42291 , \42292 , \42293 , \42294 , \42295 , \42296 ,
         \42297 , \42298 , \42299 , \42300 , \42301 , \42302 , \42303 , \42304 , \42305 , \42306 ,
         \42307 , \42308 , \42309 , \42310 , \42311 , \42312 , \42313 , \42314 , \42315 , \42316 ,
         \42317 , \42318 , \42319 , \42320 , \42321 , \42322 , \42323 , \42324 , \42325 , \42326 ,
         \42327 , \42328 , \42329 , \42330 , \42331 , \42332 , \42333 , \42334 , \42335 , \42336 ,
         \42337 , \42338 , \42339 , \42340 , \42341 , \42342 , \42343 , \42344 , \42345 , \42346 ,
         \42347 , \42348 , \42349 , \42350 , \42351 , \42352 , \42353 , \42354 , \42355 , \42356 ,
         \42357 , \42358 , \42359 , \42360 , \42361 , \42362 , \42363 , \42364 , \42365 , \42366 ,
         \42367 , \42368 , \42369 , \42370 , \42371 , \42372 , \42373 , \42374 , \42375 , \42376 ,
         \42377 , \42378 , \42379 , \42380 , \42381 , \42382 , \42383 , \42384 , \42385 , \42386 ,
         \42387 , \42388 , \42389 , \42390 , \42391 , \42392 , \42393 , \42394 , \42395 , \42396 ,
         \42397 , \42398 , \42399 , \42400 , \42401 , \42402 , \42403 , \42404 , \42405 , \42406 ,
         \42407 , \42408 , \42409 , \42410 , \42411 , \42412 , \42413 , \42414 , \42415 , \42416 ,
         \42417 , \42418 , \42419 , \42420 , \42421 , \42422 , \42423 , \42424 , \42425 , \42426 ,
         \42427 , \42428 , \42429 , \42430 , \42431 , \42432 , \42433 , \42434 , \42435 , \42436 ,
         \42437 , \42438 , \42439 , \42440 , \42441 , \42442 , \42443 , \42444 , \42445 , \42446 ,
         \42447 , \42448 , \42449 , \42450 , \42451 , \42452 , \42453 , \42454 , \42455 , \42456 ,
         \42457 , \42458 , \42459 , \42460 , \42461 , \42462 , \42463 , \42464 , \42465 , \42466 ,
         \42467 , \42468 , \42469 , \42470 , \42471 , \42472 , \42473 , \42474 , \42475 , \42476 ,
         \42477 , \42478 , \42479 , \42480 , \42481 , \42482 , \42483 , \42484 , \42485 , \42486 ,
         \42487 , \42488 , \42489 , \42490 , \42491 , \42492 , \42493 , \42494 , \42495 , \42496 ,
         \42497 , \42498 , \42499 , \42500 , \42501 , \42502 , \42503 , \42504 , \42505 , \42506 ,
         \42507 , \42508 , \42509 , \42510 , \42511 , \42512 , \42513 , \42514 , \42515 , \42516 ,
         \42517 , \42518 , \42519 , \42520 , \42521 , \42522 , \42523 , \42524 , \42525 , \42526 ,
         \42527 , \42528 , \42529 , \42530 , \42531 , \42532 , \42533 , \42534 , \42535 , \42536 ,
         \42537 , \42538 , \42539 , \42540 , \42541 , \42542 , \42543 , \42544 , \42545 , \42546 ,
         \42547 , \42548 , \42549 , \42550 , \42551 , \42552 , \42553 , \42554 , \42555 , \42556 ,
         \42557 , \42558 , \42559 , \42560 , \42561 , \42562 , \42563 , \42564 , \42565 , \42566 ,
         \42567 , \42568 , \42569 , \42570 , \42571 , \42572 , \42573 , \42574 , \42575 , \42576 ,
         \42577 , \42578 , \42579 , \42580 , \42581 , \42582 , \42583 , \42584 , \42585 , \42586 ,
         \42587 , \42588 , \42589 , \42590 , \42591 , \42592 , \42593 , \42594 , \42595 , \42596 ,
         \42597 , \42598 , \42599 , \42600 , \42601 , \42602 , \42603 , \42604 , \42605 , \42606 ,
         \42607 , \42608 , \42609 , \42610 , \42611 , \42612 , \42613 , \42614 , \42615 , \42616 ,
         \42617 , \42618 , \42619 , \42620 , \42621 , \42622 , \42623 , \42624 , \42625 , \42626 ,
         \42627 , \42628 , \42629 , \42630 , \42631 , \42632 , \42633 , \42634 , \42635 , \42636 ,
         \42637 , \42638 , \42639 , \42640 , \42641 , \42642 , \42643 , \42644 , \42645 , \42646 ,
         \42647 , \42648 , \42649 , \42650 , \42651 , \42652 , \42653 , \42654 , \42655 , \42656 ,
         \42657 , \42658 , \42659 , \42660 , \42661 , \42662 , \42663 , \42664 , \42665 , \42666 ,
         \42667 , \42668 , \42669 , \42670 , \42671 , \42672 , \42673 , \42674 , \42675 , \42676 ,
         \42677 , \42678 , \42679 , \42680 , \42681 , \42682 , \42683 , \42684 , \42685 , \42686 ,
         \42687 , \42688 , \42689 , \42690 , \42691 , \42692 , \42693 , \42694 , \42695 , \42696 ,
         \42697 , \42698 , \42699 , \42700 , \42701 , \42702 , \42703 , \42704 , \42705 , \42706 ,
         \42707 , \42708 , \42709 , \42710 , \42711 , \42712 , \42713 , \42714 , \42715 , \42716 ,
         \42717 , \42718 , \42719 , \42720 , \42721 , \42722 , \42723 , \42724 , \42725 , \42726 ,
         \42727 , \42728 , \42729 , \42730 , \42731 , \42732 , \42733 , \42734 , \42735 , \42736 ,
         \42737 , \42738 , \42739 , \42740 , \42741 , \42742 , \42743 , \42744 , \42745 , \42746 ,
         \42747 , \42748 , \42749 , \42750 , \42751 , \42752 , \42753 , \42754 , \42755 , \42756 ,
         \42757 , \42758 , \42759 , \42760 , \42761 , \42762 , \42763 , \42764 , \42765 , \42766 ,
         \42767 , \42768 , \42769 , \42770 , \42771 , \42772 , \42773 , \42774 , \42775 , \42776 ,
         \42777 , \42778 , \42779 , \42780 , \42781 , \42782 , \42783 , \42784 , \42785 , \42786 ,
         \42787 , \42788 , \42789 , \42790 , \42791 , \42792 , \42793 , \42794 , \42795 , \42796 ,
         \42797 , \42798 , \42799 , \42800 , \42801 , \42802 , \42803 , \42804 , \42805 , \42806 ,
         \42807 , \42808 , \42809 , \42810 , \42811 , \42812 , \42813 , \42814 , \42815 , \42816 ,
         \42817 , \42818 , \42819 , \42820 , \42821 , \42822 , \42823 , \42824 , \42825 , \42826 ,
         \42827 , \42828 , \42829 , \42830 , \42831 , \42832 , \42833 , \42834 , \42835 , \42836 ,
         \42837 , \42838 , \42839 , \42840 , \42841 , \42842 , \42843 , \42844 , \42845 , \42846 ,
         \42847 , \42848 , \42849 , \42850 , \42851 , \42852 , \42853 , \42854 , \42855 , \42856 ,
         \42857 , \42858 , \42859 , \42860 , \42861 , \42862 , \42863 , \42864 , \42865 , \42866 ,
         \42867 , \42868 , \42869 , \42870 , \42871 , \42872 , \42873 , \42874 , \42875 , \42876 ,
         \42877 , \42878 , \42879 , \42880 , \42881 , \42882 , \42883 , \42884 , \42885 , \42886 ,
         \42887 , \42888 , \42889 , \42890 , \42891 , \42892 , \42893 , \42894 , \42895 , \42896 ,
         \42897 , \42898 , \42899 , \42900 , \42901 , \42902 , \42903 , \42904 , \42905 , \42906 ,
         \42907 , \42908 , \42909 , \42910 , \42911 , \42912 , \42913 , \42914 , \42915 , \42916 ,
         \42917 , \42918 , \42919 , \42920 , \42921 , \42922 , \42923 , \42924 , \42925 , \42926 ,
         \42927 , \42928 , \42929 , \42930 , \42931 , \42932 , \42933 , \42934 , \42935 , \42936 ,
         \42937 , \42938 , \42939 , \42940 , \42941 , \42942 , \42943 , \42944 , \42945 , \42946 ,
         \42947 , \42948 , \42949 , \42950 , \42951 , \42952 , \42953 , \42954 , \42955 , \42956 ,
         \42957 , \42958 , \42959 , \42960 , \42961 , \42962 , \42963 , \42964 , \42965 , \42966 ,
         \42967 , \42968 , \42969 , \42970 , \42971 , \42972 , \42973 , \42974 , \42975 , \42976 ,
         \42977 , \42978 , \42979 , \42980 , \42981 , \42982 , \42983 , \42984 , \42985 , \42986 ,
         \42987 , \42988 , \42989 , \42990 , \42991 , \42992 , \42993 , \42994 , \42995 , \42996 ,
         \42997 , \42998 , \42999 , \43000 , \43001 , \43002 , \43003 , \43004 , \43005 , \43006 ,
         \43007 , \43008 , \43009 , \43010 , \43011 , \43012 , \43013 , \43014 , \43015 , \43016 ,
         \43017 , \43018 , \43019 , \43020 , \43021 , \43022 , \43023 , \43024 , \43025 , \43026 ,
         \43027 , \43028 , \43029 , \43030 , \43031 , \43032 , \43033 , \43034 , \43035 , \43036 ,
         \43037 , \43038 , \43039 , \43040 , \43041 , \43042 , \43043 , \43044 , \43045 , \43046 ,
         \43047 , \43048 , \43049 , \43050 , \43051 , \43052 , \43053 , \43054 , \43055 , \43056 ,
         \43057 , \43058 , \43059 , \43060 , \43061 , \43062 , \43063 , \43064 , \43065 , \43066 ,
         \43067 , \43068 , \43069 , \43070 , \43071 , \43072 , \43073 , \43074 , \43075 , \43076 ,
         \43077 , \43078 , \43079 , \43080 , \43081 , \43082 , \43083 , \43084 , \43085 , \43086 ,
         \43087 , \43088 , \43089 , \43090 , \43091 , \43092 , \43093 , \43094 , \43095 , \43096 ,
         \43097 , \43098 , \43099 , \43100 , \43101 , \43102 , \43103 , \43104 , \43105 , \43106 ,
         \43107 , \43108 , \43109 , \43110 , \43111 , \43112 , \43113 , \43114 , \43115 , \43116 ,
         \43117 , \43118 , \43119 , \43120 , \43121 , \43122 , \43123 , \43124 , \43125 , \43126 ,
         \43127 , \43128 , \43129 , \43130 , \43131 , \43132 , \43133 , \43134 , \43135 , \43136 ,
         \43137 , \43138 , \43139 , \43140 , \43141 , \43142 , \43143 , \43144 , \43145 , \43146 ,
         \43147 , \43148 , \43149 , \43150 , \43151 , \43152 , \43153 , \43154 , \43155 , \43156 ,
         \43157 , \43158 , \43159 , \43160 , \43161 , \43162 , \43163 , \43164 , \43165 , \43166 ,
         \43167 , \43168 , \43169 , \43170 , \43171 , \43172 , \43173 , \43174 , \43175 , \43176 ,
         \43177 , \43178 , \43179 , \43180 , \43181 , \43182 , \43183 , \43184 , \43185 , \43186 ,
         \43187 , \43188 , \43189 , \43190 , \43191 , \43192 , \43193 , \43194 , \43195 , \43196 ,
         \43197 , \43198 , \43199 , \43200 , \43201 , \43202 , \43203 , \43204 , \43205 , \43206 ,
         \43207 , \43208 , \43209 , \43210 , \43211 , \43212 , \43213 , \43214 , \43215 , \43216 ,
         \43217 , \43218 , \43219 , \43220 , \43221 , \43222 , \43223 , \43224 , \43225 , \43226 ,
         \43227 , \43228 , \43229 , \43230 , \43231 , \43232 , \43233 , \43234 , \43235 , \43236 ,
         \43237 , \43238 , \43239 , \43240 , \43241 , \43242 , \43243 , \43244 , \43245 , \43246 ,
         \43247 , \43248 , \43249 , \43250 , \43251 , \43252 , \43253 , \43254 , \43255 , \43256 ,
         \43257 , \43258 , \43259 , \43260 , \43261 , \43262 , \43263 , \43264 , \43265 , \43266 ,
         \43267 , \43268 , \43269 , \43270 , \43271 , \43272 , \43273 , \43274 , \43275 , \43276 ,
         \43277 , \43278 , \43279 , \43280 , \43281 , \43282 , \43283 , \43284 , \43285 , \43286 ,
         \43287 , \43288 , \43289 , \43290 , \43291 , \43292 , \43293 , \43294 , \43295 , \43296 ,
         \43297 , \43298 , \43299 , \43300 , \43301 , \43302 , \43303 , \43304 , \43305 , \43306 ,
         \43307 , \43308 , \43309 , \43310 , \43311 , \43312 , \43313 , \43314 , \43315 , \43316 ,
         \43317 , \43318 , \43319 , \43320 , \43321 , \43322 , \43323 , \43324 , \43325 , \43326 ,
         \43327 , \43328 , \43329 , \43330 , \43331 , \43332 , \43333 , \43334 , \43335 , \43336 ,
         \43337 , \43338 , \43339 , \43340 , \43341 , \43342 , \43343 , \43344 , \43345 , \43346 ,
         \43347 , \43348 , \43349 , \43350 , \43351 , \43352 , \43353 , \43354 , \43355 , \43356 ,
         \43357 , \43358 , \43359 , \43360 , \43361 , \43362 , \43363 , \43364 , \43365 , \43366 ,
         \43367 , \43368 , \43369 , \43370 , \43371 , \43372 , \43373 , \43374 , \43375 , \43376 ,
         \43377 , \43378 , \43379 , \43380 , \43381 , \43382 , \43383 , \43384 , \43385 , \43386 ,
         \43387 , \43388 , \43389 , \43390 , \43391 , \43392 , \43393 , \43394 , \43395 , \43396 ,
         \43397 , \43398 , \43399 , \43400 , \43401 , \43402 , \43403 , \43404 , \43405 , \43406 ,
         \43407 , \43408 , \43409 , \43410 , \43411 , \43412 , \43413 , \43414 , \43415 , \43416 ,
         \43417 , \43418 , \43419 , \43420 , \43421 , \43422 , \43423 , \43424 , \43425 , \43426 ,
         \43427 , \43428 , \43429 , \43430 , \43431 , \43432 , \43433 , \43434 , \43435 , \43436 ,
         \43437 , \43438 , \43439 , \43440 , \43441 , \43442 , \43443 , \43444 , \43445 , \43446 ,
         \43447 , \43448 , \43449 , \43450 , \43451 , \43452 , \43453 , \43454 , \43455 , \43456 ,
         \43457 , \43458 , \43459 , \43460 , \43461 , \43462 , \43463 , \43464 , \43465 , \43466 ,
         \43467 , \43468 , \43469 , \43470 , \43471 , \43472 , \43473 , \43474 , \43475 , \43476 ,
         \43477 , \43478 , \43479 , \43480 , \43481 , \43482 , \43483 , \43484 , \43485 , \43486 ,
         \43487 , \43488 , \43489 , \43490 , \43491 , \43492 , \43493 , \43494 , \43495 , \43496 ,
         \43497 , \43498 , \43499 , \43500 , \43501 , \43502 , \43503 , \43504 , \43505 , \43506 ,
         \43507 , \43508 , \43509 , \43510 , \43511 , \43512 , \43513 , \43514 , \43515 , \43516 ,
         \43517 , \43518 , \43519 , \43520 , \43521 , \43522 , \43523 , \43524 , \43525 , \43526 ,
         \43527 , \43528 , \43529 , \43530 , \43531 , \43532 , \43533 , \43534 , \43535 , \43536 ,
         \43537 , \43538 , \43539 , \43540 , \43541 , \43542 , \43543 , \43544 , \43545 , \43546 ,
         \43547 , \43548 , \43549 , \43550 , \43551 , \43552 , \43553 , \43554 , \43555 , \43556 ,
         \43557 , \43558 , \43559 , \43560 , \43561 , \43562 , \43563 , \43564 , \43565 , \43566 ,
         \43567 , \43568 , \43569 , \43570 , \43571 , \43572 , \43573 , \43574 , \43575 , \43576 ,
         \43577 , \43578 , \43579 , \43580 , \43581 , \43582 , \43583 , \43584 , \43585 , \43586 ,
         \43587 , \43588 , \43589 , \43590 , \43591 , \43592 , \43593 , \43594 , \43595 , \43596 ,
         \43597 , \43598 , \43599 , \43600 , \43601 , \43602 , \43603 , \43604 , \43605 , \43606 ,
         \43607 , \43608 , \43609 , \43610 , \43611 , \43612 , \43613 , \43614 , \43615 , \43616 ,
         \43617 , \43618 , \43619 , \43620 , \43621 , \43622 , \43623 , \43624 , \43625 , \43626 ,
         \43627 , \43628 , \43629 , \43630 , \43631 , \43632 , \43633 , \43634 , \43635 , \43636 ,
         \43637 , \43638 , \43639 , \43640 , \43641 , \43642 , \43643 , \43644 , \43645 , \43646 ,
         \43647 , \43648 , \43649 , \43650 , \43651 , \43652 , \43653 , \43654 , \43655 , \43656 ,
         \43657 , \43658 , \43659 , \43660 , \43661 , \43662 , \43663 , \43664 , \43665 , \43666 ,
         \43667 , \43668 , \43669 , \43670 , \43671 , \43672 , \43673 , \43674 , \43675 , \43676 ,
         \43677 , \43678 , \43679 , \43680 , \43681 , \43682 , \43683 , \43684 , \43685 , \43686 ,
         \43687 , \43688 , \43689 , \43690 , \43691 , \43692 , \43693 , \43694 , \43695 , \43696 ,
         \43697 , \43698 , \43699 , \43700 , \43701 , \43702 , \43703 , \43704 , \43705 , \43706 ,
         \43707 , \43708 , \43709 , \43710 , \43711 , \43712 , \43713 , \43714 , \43715 , \43716 ,
         \43717 , \43718 , \43719 , \43720 , \43721 , \43722 , \43723 , \43724 , \43725 , \43726 ,
         \43727 , \43728 , \43729 , \43730 , \43731 , \43732 , \43733 , \43734 , \43735 , \43736 ,
         \43737 , \43738 , \43739 , \43740 , \43741 , \43742 , \43743 , \43744 , \43745 , \43746 ,
         \43747 , \43748 , \43749 , \43750 , \43751 , \43752 , \43753 , \43754 , \43755 , \43756 ,
         \43757 , \43758 , \43759 , \43760 , \43761 , \43762 , \43763 , \43764 , \43765 , \43766 ,
         \43767 , \43768 , \43769 , \43770 , \43771 , \43772 , \43773 , \43774 , \43775 , \43776 ,
         \43777 , \43778 , \43779 , \43780 , \43781 , \43782 , \43783 , \43784 , \43785 , \43786 ,
         \43787 , \43788 , \43789 , \43790 , \43791 , \43792 , \43793 , \43794 , \43795 , \43796 ,
         \43797 , \43798 , \43799 , \43800 , \43801 , \43802 , \43803 , \43804 , \43805 , \43806 ,
         \43807 , \43808 , \43809 , \43810 , \43811 , \43812 , \43813 , \43814 , \43815 , \43816 ,
         \43817 , \43818 , \43819 , \43820 , \43821 , \43822 , \43823 , \43824 , \43825 , \43826 ,
         \43827 , \43828 , \43829 , \43830 , \43831 , \43832 , \43833 , \43834 , \43835 , \43836 ,
         \43837 , \43838 , \43839 , \43840 , \43841 , \43842 , \43843 , \43844 , \43845 , \43846 ,
         \43847 , \43848 , \43849 , \43850 , \43851 , \43852 , \43853 , \43854 , \43855 , \43856 ,
         \43857 , \43858 , \43859 , \43860 , \43861 , \43862 , \43863 , \43864 , \43865 , \43866 ,
         \43867 , \43868 , \43869 , \43870 , \43871 , \43872 , \43873 , \43874 , \43875 , \43876 ,
         \43877 , \43878 , \43879 , \43880 , \43881 , \43882 , \43883 , \43884 , \43885 , \43886 ,
         \43887 , \43888 , \43889 , \43890 , \43891 , \43892 , \43893 , \43894 , \43895 , \43896 ,
         \43897 , \43898 , \43899 , \43900 , \43901 , \43902 , \43903 , \43904 , \43905 , \43906 ,
         \43907 , \43908 , \43909 , \43910 , \43911 , \43912 , \43913 , \43914 , \43915 , \43916 ,
         \43917 , \43918 , \43919 , \43920 , \43921 , \43922 , \43923 , \43924 , \43925 , \43926 ,
         \43927 , \43928 , \43929 , \43930 , \43931 , \43932 , \43933 , \43934 , \43935 , \43936 ,
         \43937 , \43938 , \43939 , \43940 , \43941 , \43942 , \43943 , \43944 , \43945 , \43946 ,
         \43947 , \43948 , \43949 , \43950 , \43951 , \43952 , \43953 , \43954 , \43955 , \43956 ,
         \43957 , \43958 , \43959 , \43960 , \43961 , \43962 , \43963 , \43964 , \43965 , \43966 ,
         \43967 , \43968 , \43969 , \43970 , \43971 , \43972 , \43973 , \43974 , \43975 , \43976 ,
         \43977 , \43978 , \43979 , \43980 , \43981 , \43982 , \43983 , \43984 , \43985 , \43986 ,
         \43987 , \43988 , \43989 , \43990 , \43991 , \43992 , \43993 , \43994 , \43995 , \43996 ,
         \43997 , \43998 , \43999 , \44000 , \44001 , \44002 , \44003 , \44004 , \44005 , \44006 ,
         \44007 , \44008 , \44009 , \44010 , \44011 , \44012 , \44013 , \44014 , \44015 , \44016 ,
         \44017 , \44018 , \44019 , \44020 , \44021 , \44022 , \44023 , \44024 , \44025 , \44026 ,
         \44027 , \44028 , \44029 , \44030 , \44031 , \44032 , \44033 , \44034 , \44035 , \44036 ,
         \44037 , \44038 , \44039 , \44040 , \44041 , \44042 , \44043 , \44044 , \44045 , \44046 ,
         \44047 , \44048 , \44049 , \44050 , \44051 , \44052 , \44053 , \44054 , \44055 , \44056 ,
         \44057 , \44058 , \44059 , \44060 , \44061 , \44062 , \44063 , \44064 , \44065 , \44066 ,
         \44067 , \44068 , \44069 , \44070 , \44071 , \44072 , \44073 , \44074 , \44075 , \44076 ,
         \44077 , \44078 , \44079 , \44080 , \44081 , \44082 , \44083 , \44084 , \44085 , \44086 ,
         \44087 , \44088 , \44089 , \44090 , \44091 , \44092 , \44093 , \44094 , \44095 , \44096 ,
         \44097 , \44098 , \44099 , \44100 , \44101 , \44102 , \44103 , \44104 , \44105 , \44106 ,
         \44107 , \44108 , \44109 , \44110 , \44111 , \44112 , \44113 , \44114 , \44115 , \44116 ,
         \44117 , \44118 , \44119 , \44120 , \44121 , \44122 , \44123 , \44124 , \44125 , \44126 ,
         \44127 , \44128 , \44129 , \44130 , \44131 , \44132 , \44133 , \44134 , \44135 , \44136 ,
         \44137 , \44138 , \44139 , \44140 , \44141 , \44142 , \44143 , \44144 , \44145 , \44146 ,
         \44147 , \44148 , \44149 , \44150 , \44151 , \44152 , \44153 , \44154 , \44155 , \44156 ,
         \44157 , \44158 , \44159 , \44160 , \44161 , \44162 , \44163 , \44164 , \44165 , \44166 ,
         \44167 , \44168 , \44169 , \44170 , \44171 , \44172 , \44173 , \44174 , \44175 , \44176 ,
         \44177 , \44178 , \44179 , \44180 , \44181 , \44182 , \44183 , \44184 , \44185 , \44186 ,
         \44187 , \44188 , \44189 , \44190 , \44191 , \44192 , \44193 , \44194 , \44195 , \44196 ,
         \44197 , \44198 , \44199 , \44200 , \44201 , \44202 , \44203 , \44204 , \44205 , \44206 ,
         \44207 , \44208 , \44209 , \44210 , \44211 , \44212 , \44213 , \44214 , \44215 , \44216 ,
         \44217 , \44218 , \44219 , \44220 , \44221 , \44222 , \44223 , \44224 , \44225 , \44226 ,
         \44227 , \44228 , \44229 , \44230 , \44231 , \44232 , \44233 , \44234 , \44235 , \44236 ,
         \44237 , \44238 , \44239 , \44240 , \44241 , \44242 , \44243 , \44244 , \44245 , \44246 ,
         \44247 , \44248 , \44249 , \44250 , \44251 , \44252 , \44253 , \44254 , \44255 , \44256 ,
         \44257 , \44258 , \44259 , \44260 , \44261 , \44262 , \44263 , \44264 , \44265 , \44266 ,
         \44267 , \44268 , \44269 , \44270 , \44271 , \44272 , \44273 , \44274 , \44275 , \44276 ,
         \44277 , \44278 , \44279 , \44280 , \44281 , \44282 , \44283 , \44284 , \44285 , \44286 ,
         \44287 , \44288 , \44289 , \44290 , \44291 , \44292 , \44293 , \44294 , \44295 , \44296 ,
         \44297 , \44298 , \44299 , \44300 , \44301 , \44302 , \44303 , \44304 , \44305 , \44306 ,
         \44307 , \44308 , \44309 , \44310 , \44311 , \44312 , \44313 , \44314 , \44315 , \44316 ,
         \44317 , \44318 , \44319 , \44320 , \44321 , \44322 , \44323 , \44324 , \44325 , \44326 ,
         \44327 , \44328 , \44329 , \44330 , \44331 , \44332 , \44333 , \44334 , \44335 , \44336 ,
         \44337 , \44338 , \44339 , \44340 , \44341 , \44342 , \44343 , \44344 , \44345 , \44346 ,
         \44347 , \44348 , \44349 , \44350 , \44351 , \44352 , \44353 , \44354 , \44355 , \44356 ,
         \44357 , \44358 , \44359 , \44360 , \44361 , \44362 , \44363 , \44364 , \44365 , \44366 ,
         \44367 , \44368 , \44369 , \44370 , \44371 , \44372 , \44373 , \44374 , \44375 , \44376 ,
         \44377 , \44378 , \44379 , \44380 , \44381 , \44382 , \44383 , \44384 , \44385 , \44386 ,
         \44387 , \44388 , \44389 , \44390 , \44391 , \44392 , \44393 , \44394 , \44395 , \44396 ,
         \44397 , \44398 , \44399 , \44400 , \44401 , \44402 , \44403 , \44404 , \44405 , \44406 ,
         \44407 , \44408 , \44409 , \44410 , \44411 , \44412 , \44413 , \44414 , \44415 , \44416 ,
         \44417 , \44418 , \44419 , \44420 , \44421 , \44422 , \44423 , \44424 , \44425 , \44426 ,
         \44427 , \44428 , \44429 , \44430 , \44431 , \44432 , \44433 , \44434 , \44435 , \44436 ,
         \44437 , \44438 , \44439 , \44440 , \44441 , \44442 , \44443 , \44444 , \44445 , \44446 ,
         \44447 , \44448 , \44449 , \44450 , \44451 , \44452 , \44453 , \44454 , \44455 , \44456 ,
         \44457 , \44458 , \44459 , \44460 , \44461 , \44462 , \44463 , \44464 , \44465 , \44466 ,
         \44467 , \44468 , \44469 , \44470 , \44471 , \44472 , \44473 , \44474 , \44475 , \44476 ,
         \44477 , \44478 , \44479 , \44480 , \44481 , \44482 , \44483 , \44484 , \44485 , \44486 ,
         \44487 , \44488 , \44489 , \44490 , \44491 , \44492 , \44493 , \44494 , \44495 , \44496 ,
         \44497 , \44498 , \44499 , \44500 , \44501 , \44502 , \44503 , \44504 , \44505 , \44506 ,
         \44507 , \44508 , \44509 , \44510 , \44511 , \44512 , \44513 , \44514 , \44515 , \44516 ,
         \44517 , \44518 , \44519 , \44520 , \44521 , \44522 , \44523 , \44524 , \44525 , \44526 ,
         \44527 , \44528 , \44529 , \44530 , \44531 , \44532 , \44533 , \44534 , \44535 , \44536 ,
         \44537 , \44538 , \44539 , \44540 , \44541 , \44542 , \44543 , \44544 , \44545 , \44546 ,
         \44547 , \44548 , \44549 , \44550 , \44551 , \44552 , \44553 , \44554 , \44555 , \44556 ,
         \44557 , \44558 , \44559 , \44560 , \44561 , \44562 , \44563 , \44564 , \44565 , \44566 ,
         \44567 , \44568 , \44569 , \44570 , \44571 , \44572 , \44573 , \44574 , \44575 , \44576 ,
         \44577 , \44578 , \44579 , \44580 , \44581 , \44582 , \44583 , \44584 , \44585 , \44586 ,
         \44587 , \44588 , \44589 , \44590 , \44591 , \44592 , \44593 , \44594 , \44595 , \44596 ,
         \44597 , \44598 , \44599 , \44600 , \44601 , \44602 , \44603 , \44604 , \44605 , \44606 ,
         \44607 , \44608 , \44609 , \44610 , \44611 , \44612 , \44613 , \44614 , \44615 , \44616 ,
         \44617 , \44618 , \44619 , \44620 , \44621 , \44622 , \44623 , \44624 , \44625 , \44626 ,
         \44627 , \44628 , \44629 , \44630 , \44631 , \44632 , \44633 , \44634 , \44635 , \44636 ,
         \44637 , \44638 , \44639 , \44640 , \44641 , \44642 , \44643 , \44644 , \44645 , \44646 ,
         \44647 , \44648 , \44649 , \44650 , \44651 , \44652 , \44653 , \44654 , \44655 , \44656 ,
         \44657 , \44658 , \44659 , \44660 , \44661 , \44662 , \44663 , \44664 , \44665 , \44666 ,
         \44667 , \44668 , \44669 , \44670 , \44671 , \44672 , \44673 , \44674 , \44675 , \44676 ,
         \44677 , \44678 , \44679 , \44680 , \44681 , \44682 , \44683 , \44684 , \44685 , \44686 ,
         \44687 , \44688 , \44689 , \44690 , \44691 , \44692 , \44693 , \44694 , \44695 , \44696 ,
         \44697 , \44698 , \44699 , \44700 , \44701 , \44702 , \44703 , \44704 , \44705 , \44706 ,
         \44707 , \44708 , \44709 , \44710 , \44711 , \44712 , \44713 , \44714 , \44715 , \44716 ,
         \44717 , \44718 , \44719 , \44720 , \44721 , \44722 , \44723 , \44724 , \44725 , \44726 ,
         \44727 , \44728 , \44729 , \44730 , \44731 , \44732 , \44733 , \44734 , \44735 , \44736 ,
         \44737 , \44738 , \44739 , \44740 , \44741 , \44742 , \44743 , \44744 , \44745 , \44746 ,
         \44747 , \44748 , \44749 , \44750 , \44751 , \44752 , \44753 , \44754 , \44755 , \44756 ,
         \44757 , \44758 , \44759 , \44760 , \44761 , \44762 , \44763 , \44764 , \44765 , \44766 ,
         \44767 , \44768 , \44769 , \44770 , \44771 , \44772 , \44773 , \44774 , \44775 , \44776 ,
         \44777 , \44778 , \44779 , \44780 , \44781 , \44782 , \44783 , \44784 , \44785 , \44786 ,
         \44787 , \44788 , \44789 , \44790 , \44791 , \44792 , \44793 , \44794 , \44795 , \44796 ,
         \44797 , \44798 , \44799 , \44800 , \44801 , \44802 , \44803 , \44804 , \44805 , \44806 ,
         \44807 , \44808 , \44809 , \44810 , \44811 , \44812 , \44813 , \44814 , \44815 , \44816 ,
         \44817 , \44818 , \44819 , \44820 , \44821 , \44822 , \44823 , \44824 , \44825 , \44826 ,
         \44827 , \44828 , \44829 , \44830 , \44831 , \44832 , \44833 , \44834 , \44835 , \44836 ,
         \44837 , \44838 , \44839 , \44840 , \44841 , \44842 , \44843 , \44844 , \44845 , \44846 ,
         \44847 , \44848 , \44849 , \44850 , \44851 , \44852 , \44853 , \44854 , \44855 , \44856 ,
         \44857 , \44858 , \44859 , \44860 , \44861 , \44862 , \44863 , \44864 , \44865 , \44866 ,
         \44867 , \44868 , \44869 , \44870 , \44871 , \44872 , \44873 , \44874 , \44875 , \44876 ,
         \44877 , \44878 , \44879 , \44880 , \44881 , \44882 , \44883 , \44884 , \44885 , \44886 ,
         \44887 , \44888 , \44889 , \44890 , \44891 , \44892 , \44893 , \44894 , \44895 , \44896 ,
         \44897 , \44898 , \44899 , \44900 , \44901 , \44902 , \44903 , \44904 , \44905 , \44906 ,
         \44907 , \44908 , \44909 , \44910 , \44911 , \44912 , \44913 , \44914 , \44915 , \44916 ,
         \44917 , \44918 , \44919 , \44920 , \44921 , \44922 , \44923 , \44924 , \44925 , \44926 ,
         \44927 , \44928 , \44929 , \44930 , \44931 , \44932 , \44933 , \44934 , \44935 , \44936 ,
         \44937 , \44938 , \44939 , \44940 , \44941 , \44942 , \44943 , \44944 , \44945 , \44946 ,
         \44947 , \44948 , \44949 , \44950 , \44951 , \44952 , \44953 , \44954 , \44955 , \44956 ,
         \44957 , \44958 , \44959 , \44960 , \44961 , \44962 , \44963 , \44964 , \44965 , \44966 ,
         \44967 , \44968 , \44969 , \44970 , \44971 , \44972 , \44973 , \44974 , \44975 , \44976 ,
         \44977 , \44978 , \44979 , \44980 , \44981 , \44982 , \44983 , \44984 , \44985 , \44986 ,
         \44987 , \44988 , \44989 , \44990 , \44991 , \44992 , \44993 , \44994 , \44995 , \44996 ,
         \44997 , \44998 , \44999 , \45000 , \45001 , \45002 , \45003 , \45004 , \45005 , \45006 ,
         \45007 , \45008 , \45009 , \45010 , \45011 , \45012 , \45013 , \45014 , \45015 , \45016 ,
         \45017 , \45018 , \45019 , \45020 , \45021 , \45022 , \45023 , \45024 , \45025 , \45026 ,
         \45027 , \45028 , \45029 , \45030 , \45031 , \45032 , \45033 , \45034 , \45035 , \45036 ,
         \45037 , \45038 , \45039 , \45040 , \45041 , \45042 , \45043 , \45044 , \45045 , \45046 ,
         \45047 , \45048 , \45049 , \45050 , \45051 , \45052 , \45053 , \45054 , \45055 , \45056 ,
         \45057 , \45058 , \45059 , \45060 , \45061 , \45062 , \45063 , \45064 , \45065 , \45066 ,
         \45067 , \45068 , \45069 , \45070 , \45071 , \45072 , \45073 , \45074 , \45075 , \45076 ,
         \45077 , \45078 , \45079 , \45080 , \45081 , \45082 , \45083 , \45084 , \45085 , \45086 ,
         \45087 , \45088 , \45089 , \45090 , \45091 , \45092 , \45093 , \45094 , \45095 , \45096 ,
         \45097 , \45098 , \45099 , \45100 , \45101 , \45102 , \45103 , \45104 , \45105 , \45106 ,
         \45107 , \45108 , \45109 , \45110 , \45111 , \45112 , \45113 , \45114 , \45115 , \45116 ,
         \45117 , \45118 , \45119 , \45120 , \45121 , \45122 , \45123 , \45124 , \45125 , \45126 ,
         \45127 , \45128 , \45129 , \45130 , \45131 , \45132 , \45133 , \45134 , \45135 , \45136 ,
         \45137 , \45138 , \45139 , \45140 , \45141 , \45142 , \45143 , \45144 , \45145 , \45146 ,
         \45147 , \45148 , \45149 , \45150 , \45151 , \45152 , \45153 , \45154 , \45155 , \45156 ,
         \45157 , \45158 , \45159 , \45160 , \45161 , \45162 , \45163 , \45164 , \45165 , \45166 ,
         \45167 , \45168 , \45169 , \45170 , \45171 , \45172 , \45173 , \45174 , \45175 , \45176 ,
         \45177 , \45178 , \45179 , \45180 , \45181 , \45182 , \45183 , \45184 , \45185 , \45186 ,
         \45187 , \45188 , \45189 , \45190 , \45191 , \45192 , \45193 , \45194 , \45195 , \45196 ,
         \45197 , \45198 , \45199 , \45200 , \45201 , \45202 , \45203 , \45204 , \45205 , \45206 ,
         \45207 , \45208 , \45209 , \45210 , \45211 , \45212 , \45213 , \45214 , \45215 , \45216 ,
         \45217 , \45218 , \45219 , \45220 , \45221 , \45222 , \45223 , \45224 , \45225 , \45226 ,
         \45227 , \45228 , \45229 , \45230 , \45231 , \45232 , \45233 , \45234 , \45235 , \45236 ,
         \45237 , \45238 , \45239 , \45240 , \45241 , \45242 , \45243 , \45244 , \45245 , \45246 ,
         \45247 , \45248 , \45249 , \45250 , \45251 , \45252 , \45253 , \45254 , \45255 , \45256 ,
         \45257 , \45258 , \45259 , \45260 , \45261 , \45262 , \45263 , \45264 , \45265 , \45266 ,
         \45267 , \45268 , \45269 , \45270 , \45271 , \45272 , \45273 , \45274 , \45275 , \45276 ,
         \45277 , \45278 , \45279 , \45280 , \45281 , \45282 , \45283 , \45284 , \45285 , \45286 ,
         \45287 , \45288 , \45289 , \45290 , \45291 , \45292 , \45293 , \45294 , \45295 , \45296 ,
         \45297 , \45298 , \45299 , \45300 , \45301 , \45302 , \45303 , \45304 , \45305 , \45306 ,
         \45307 , \45308 , \45309 , \45310 , \45311 , \45312 , \45313 , \45314 , \45315 , \45316 ,
         \45317 , \45318 , \45319 , \45320 , \45321 , \45322 , \45323 , \45324 , \45325 , \45326 ,
         \45327 , \45328 , \45329 , \45330 , \45331 , \45332 , \45333 , \45334 , \45335 , \45336 ,
         \45337 , \45338 , \45339 , \45340 , \45341 , \45342 , \45343 , \45344 , \45345 , \45346 ,
         \45347 , \45348 , \45349 , \45350 , \45351 , \45352 , \45353 , \45354 , \45355 , \45356 ,
         \45357 , \45358 , \45359 , \45360 , \45361 , \45362 , \45363 , \45364 , \45365 , \45366 ,
         \45367 , \45368 , \45369 , \45370 , \45371 , \45372 , \45373 , \45374 , \45375 , \45376 ,
         \45377 , \45378 , \45379 , \45380 , \45381 , \45382 , \45383 , \45384 , \45385 , \45386 ,
         \45387 , \45388 , \45389 , \45390 , \45391 , \45392 , \45393 , \45394 , \45395 , \45396 ,
         \45397 , \45398 , \45399 , \45400 , \45401 , \45402 , \45403 , \45404 , \45405 , \45406 ,
         \45407 , \45408 , \45409 , \45410 , \45411 , \45412 , \45413 , \45414 , \45415 , \45416 ,
         \45417 , \45418 , \45419 , \45420 , \45421 , \45422 , \45423 , \45424 , \45425 , \45426 ,
         \45427 , \45428 , \45429 , \45430 , \45431 , \45432 , \45433 , \45434 , \45435 , \45436 ,
         \45437 , \45438 , \45439 , \45440 , \45441 , \45442 , \45443 , \45444 , \45445 , \45446 ,
         \45447 , \45448 , \45449 , \45450 , \45451 , \45452 , \45453 , \45454 , \45455 , \45456 ,
         \45457 , \45458 , \45459 , \45460 , \45461 , \45462 , \45463 , \45464 , \45465 , \45466 ,
         \45467 , \45468 , \45469 , \45470 , \45471 , \45472 , \45473 , \45474 , \45475 , \45476 ,
         \45477 , \45478 , \45479 , \45480 , \45481 , \45482 , \45483 , \45484 , \45485 , \45486 ,
         \45487 , \45488 , \45489 , \45490 , \45491 , \45492 , \45493 , \45494 , \45495 , \45496 ,
         \45497 , \45498 , \45499 , \45500 , \45501 , \45502 , \45503 , \45504 , \45505 , \45506 ,
         \45507 , \45508 , \45509 , \45510 , \45511 , \45512 , \45513 , \45514 , \45515 , \45516 ,
         \45517 , \45518 , \45519 , \45520 , \45521 , \45522 , \45523 , \45524 , \45525 , \45526 ,
         \45527 , \45528 , \45529 , \45530 , \45531 , \45532 , \45533 , \45534 , \45535 , \45536 ,
         \45537 , \45538 , \45539 , \45540 , \45541 , \45542 , \45543 , \45544 , \45545 , \45546 ,
         \45547 , \45548 , \45549 , \45550 , \45551 , \45552 , \45553 , \45554 , \45555 , \45556 ,
         \45557 , \45558 , \45559 , \45560 , \45561 , \45562 , \45563 , \45564 , \45565 , \45566 ,
         \45567 , \45568 , \45569 , \45570 , \45571 , \45572 , \45573 , \45574 , \45575 , \45576 ,
         \45577 , \45578 , \45579 , \45580 , \45581 , \45582 , \45583 , \45584 , \45585 , \45586 ,
         \45587 , \45588 , \45589 , \45590 , \45591 , \45592 , \45593 , \45594 , \45595 , \45596 ,
         \45597 , \45598 , \45599 , \45600 , \45601 , \45602 , \45603 , \45604 , \45605 , \45606 ,
         \45607 , \45608 , \45609 , \45610 , \45611 , \45612 , \45613 , \45614 , \45615 , \45616 ,
         \45617 , \45618 , \45619 , \45620 , \45621 , \45622 , \45623 , \45624 , \45625 , \45626 ,
         \45627 , \45628 , \45629 , \45630 , \45631 , \45632 , \45633 , \45634 , \45635 , \45636 ,
         \45637 , \45638 , \45639 , \45640 , \45641 , \45642 , \45643 , \45644 , \45645 , \45646 ,
         \45647 , \45648 , \45649 , \45650 , \45651 , \45652 , \45653 , \45654 , \45655 , \45656 ,
         \45657 , \45658 , \45659 , \45660 , \45661 , \45662 , \45663 , \45664 , \45665 , \45666 ,
         \45667 , \45668 , \45669 , \45670 , \45671 , \45672 , \45673 , \45674 , \45675 , \45676 ,
         \45677 , \45678 , \45679 , \45680 , \45681 , \45682 , \45683 , \45684 , \45685 , \45686 ,
         \45687 , \45688 , \45689 , \45690 , \45691 , \45692 , \45693 , \45694 , \45695 , \45696 ,
         \45697 , \45698 , \45699 , \45700 , \45701 , \45702 , \45703 , \45704 , \45705 , \45706 ,
         \45707 , \45708 , \45709 , \45710 , \45711 , \45712 , \45713 , \45714 , \45715 , \45716 ,
         \45717 , \45718 , \45719 , \45720 , \45721 , \45722 , \45723 , \45724 , \45725 , \45726 ,
         \45727 , \45728 , \45729 , \45730 , \45731 , \45732 , \45733 , \45734 , \45735 , \45736 ,
         \45737 , \45738 , \45739 , \45740 , \45741 , \45742 , \45743 , \45744 , \45745 , \45746 ,
         \45747 , \45748 , \45749 , \45750 , \45751 , \45752 , \45753 , \45754 , \45755 , \45756 ,
         \45757 , \45758 , \45759 , \45760 , \45761 , \45762 , \45763 , \45764 , \45765 , \45766 ,
         \45767 , \45768 , \45769 , \45770 , \45771 , \45772 , \45773 , \45774 , \45775 , \45776 ,
         \45777 , \45778 , \45779 , \45780 , \45781 , \45782 , \45783 , \45784 , \45785 , \45786 ,
         \45787 , \45788 , \45789 , \45790 , \45791 , \45792 , \45793 , \45794 , \45795 , \45796 ,
         \45797 , \45798 , \45799 , \45800 , \45801 , \45802 , \45803 , \45804 , \45805 , \45806 ,
         \45807 , \45808 , \45809 , \45810 , \45811 , \45812 , \45813 , \45814 , \45815 , \45816 ,
         \45817 , \45818 , \45819 , \45820 , \45821 , \45822 , \45823 , \45824 , \45825 , \45826 ,
         \45827 , \45828 , \45829 , \45830 , \45831 , \45832 , \45833 , \45834 , \45835 , \45836 ,
         \45837 , \45838 , \45839 , \45840 , \45841 , \45842 , \45843 , \45844 , \45845 , \45846 ,
         \45847 , \45848 , \45849 , \45850 , \45851 , \45852 , \45853 , \45854 , \45855 , \45856 ,
         \45857 , \45858 , \45859 , \45860 , \45861 , \45862 , \45863 , \45864 , \45865 , \45866 ,
         \45867 , \45868 , \45869 , \45870 , \45871 , \45872 , \45873 , \45874 , \45875 , \45876 ,
         \45877 , \45878 , \45879 , \45880 , \45881 , \45882 , \45883 , \45884 , \45885 , \45886 ,
         \45887 , \45888 , \45889 , \45890 , \45891 , \45892 , \45893 , \45894 , \45895 , \45896 ,
         \45897 , \45898 , \45899 , \45900 , \45901 , \45902 , \45903 , \45904 , \45905 , \45906 ,
         \45907 , \45908 , \45909 , \45910 , \45911 , \45912 , \45913 , \45914 , \45915 , \45916 ,
         \45917 , \45918 , \45919 , \45920 , \45921 , \45922 , \45923 , \45924 , \45925 , \45926 ,
         \45927 , \45928 , \45929 , \45930 , \45931 , \45932 , \45933 , \45934 , \45935 , \45936 ,
         \45937 , \45938 , \45939 , \45940 , \45941 , \45942 , \45943 , \45944 , \45945 , \45946 ,
         \45947 , \45948 , \45949 , \45950 , \45951 , \45952 , \45953 , \45954 , \45955 , \45956 ,
         \45957 , \45958 , \45959 , \45960 , \45961 , \45962 , \45963 , \45964 , \45965 , \45966 ,
         \45967 , \45968 , \45969 , \45970 , \45971 , \45972 , \45973 , \45974 , \45975 , \45976 ,
         \45977 , \45978 , \45979 , \45980 , \45981 , \45982 , \45983 , \45984 , \45985 , \45986 ,
         \45987 , \45988 , \45989 , \45990 , \45991 , \45992 , \45993 , \45994 , \45995 , \45996 ,
         \45997 , \45998 , \45999 , \46000 , \46001 , \46002 , \46003 , \46004 , \46005 , \46006 ,
         \46007 , \46008 , \46009 , \46010 , \46011 , \46012 , \46013 , \46014 , \46015 , \46016 ,
         \46017 , \46018 , \46019 , \46020 , \46021 , \46022 , \46023 , \46024 , \46025 , \46026 ,
         \46027 , \46028 , \46029 , \46030 , \46031 , \46032 , \46033 , \46034 , \46035 , \46036 ,
         \46037 , \46038 , \46039 , \46040 , \46041 , \46042 , \46043 , \46044 , \46045 , \46046 ,
         \46047 , \46048 , \46049 , \46050 , \46051 , \46052 , \46053 , \46054 , \46055 , \46056 ,
         \46057 , \46058 , \46059 , \46060 , \46061 , \46062 , \46063 , \46064 , \46065 , \46066 ,
         \46067 , \46068 , \46069 , \46070 , \46071 , \46072 , \46073 , \46074 , \46075 , \46076 ,
         \46077 , \46078 , \46079 , \46080 , \46081 , \46082 , \46083 , \46084 , \46085 , \46086 ,
         \46087 , \46088 , \46089 , \46090 , \46091 , \46092 , \46093 , \46094 , \46095 , \46096 ,
         \46097 , \46098 , \46099 , \46100 , \46101 , \46102 , \46103 , \46104 , \46105 , \46106 ,
         \46107 , \46108 , \46109 , \46110 , \46111 , \46112 , \46113 , \46114 , \46115 , \46116 ,
         \46117 , \46118 , \46119 , \46120 , \46121 , \46122 , \46123 , \46124 , \46125 , \46126 ,
         \46127 , \46128 , \46129 , \46130 , \46131 , \46132 , \46133 , \46134 , \46135 , \46136 ,
         \46137 , \46138 , \46139 , \46140 , \46141 , \46142 , \46143 , \46144 , \46145 , \46146 ,
         \46147 , \46148 , \46149 , \46150 , \46151 , \46152 , \46153 , \46154 , \46155 , \46156 ,
         \46157 , \46158 , \46159 , \46160 , \46161 , \46162 , \46163 , \46164 , \46165 , \46166 ,
         \46167 , \46168 , \46169 , \46170 , \46171 , \46172 , \46173 , \46174 , \46175 , \46176 ,
         \46177 , \46178 , \46179 , \46180 , \46181 , \46182 , \46183 , \46184 , \46185 , \46186 ,
         \46187 , \46188 , \46189 , \46190 , \46191 , \46192 , \46193 , \46194 , \46195 , \46196 ,
         \46197 , \46198 , \46199 , \46200 , \46201 , \46202 , \46203 , \46204 , \46205 , \46206 ,
         \46207 , \46208 , \46209 , \46210 , \46211 , \46212 , \46213 , \46214 , \46215 , \46216 ,
         \46217 , \46218 , \46219 , \46220 , \46221 , \46222 , \46223 , \46224 , \46225 , \46226 ,
         \46227 , \46228 , \46229 , \46230 , \46231 , \46232 , \46233 , \46234 , \46235 , \46236 ,
         \46237 , \46238 , \46239 , \46240 , \46241 , \46242 , \46243 , \46244 , \46245 , \46246 ,
         \46247 , \46248 , \46249 , \46250 , \46251 , \46252 , \46253 , \46254 , \46255 , \46256 ,
         \46257 , \46258 , \46259 , \46260 , \46261 , \46262 , \46263 , \46264 , \46265 , \46266 ,
         \46267 , \46268 , \46269 , \46270 , \46271 , \46272 , \46273 , \46274 , \46275 , \46276 ,
         \46277 , \46278 , \46279 , \46280 , \46281 , \46282 , \46283 , \46284 , \46285 , \46286 ,
         \46287 , \46288 , \46289 , \46290 , \46291 , \46292 , \46293 , \46294 , \46295 , \46296 ,
         \46297 , \46298 , \46299 , \46300 , \46301 , \46302 , \46303 , \46304 , \46305 , \46306 ,
         \46307 , \46308 , \46309 , \46310 , \46311 , \46312 , \46313 , \46314 , \46315 , \46316 ,
         \46317 , \46318 , \46319 , \46320 , \46321 , \46322 , \46323 , \46324 , \46325 , \46326 ,
         \46327 , \46328 , \46329 , \46330 , \46331 , \46332 , \46333 , \46334 , \46335 , \46336 ,
         \46337 , \46338 , \46339 , \46340 , \46341 , \46342 , \46343 , \46344 , \46345 , \46346 ,
         \46347 , \46348 , \46349 , \46350 , \46351 , \46352 , \46353 , \46354 , \46355 , \46356 ,
         \46357 , \46358 , \46359 , \46360 , \46361 , \46362 , \46363 , \46364 , \46365 , \46366 ,
         \46367 , \46368 , \46369 , \46370 , \46371 , \46372 , \46373 , \46374 , \46375 , \46376 ,
         \46377 , \46378 , \46379 , \46380 , \46381 , \46382 , \46383 , \46384 , \46385 , \46386 ,
         \46387 , \46388 , \46389 , \46390 , \46391 , \46392 , \46393 , \46394 , \46395 , \46396 ,
         \46397 , \46398 , \46399 , \46400 , \46401 , \46402 , \46403 , \46404 , \46405 , \46406 ,
         \46407 , \46408 , \46409 , \46410 , \46411 , \46412 , \46413 , \46414 , \46415 , \46416 ,
         \46417 , \46418 , \46419 , \46420 , \46421 , \46422 , \46423 , \46424 , \46425 , \46426 ,
         \46427 , \46428 , \46429 , \46430 , \46431 , \46432 , \46433 , \46434 , \46435 , \46436 ,
         \46437 , \46438 , \46439 , \46440 , \46441 , \46442 , \46443 , \46444 , \46445 , \46446 ,
         \46447 , \46448 , \46449 , \46450 , \46451 , \46452 , \46453 , \46454 , \46455 , \46456 ,
         \46457 , \46458 , \46459 , \46460 , \46461 , \46462 , \46463 , \46464 , \46465 , \46466 ,
         \46467 , \46468 , \46469 , \46470 , \46471 , \46472 , \46473 , \46474 , \46475 , \46476 ,
         \46477 , \46478 , \46479 , \46480 , \46481 , \46482 , \46483 , \46484 , \46485 , \46486 ,
         \46487 , \46488 , \46489 , \46490 , \46491 , \46492 , \46493 , \46494 , \46495 , \46496 ,
         \46497 , \46498 , \46499 , \46500 , \46501 , \46502 , \46503 , \46504 , \46505 , \46506 ,
         \46507 , \46508 , \46509 , \46510 , \46511 , \46512 , \46513 , \46514 , \46515 , \46516 ,
         \46517 , \46518 , \46519 , \46520 , \46521 , \46522 , \46523 , \46524 , \46525 , \46526 ,
         \46527 , \46528 , \46529 , \46530 , \46531 , \46532 , \46533 , \46534 , \46535 , \46536 ,
         \46537 , \46538 , \46539 , \46540 , \46541 , \46542 , \46543 , \46544 , \46545 , \46546 ,
         \46547 , \46548 , \46549 , \46550 , \46551 , \46552 , \46553 , \46554 , \46555 , \46556 ,
         \46557 , \46558 , \46559 , \46560 , \46561 , \46562 , \46563 , \46564 , \46565 , \46566 ,
         \46567 , \46568 , \46569 , \46570 , \46571 , \46572 , \46573 , \46574 , \46575 , \46576 ,
         \46577 , \46578 , \46579 , \46580 , \46581 , \46582 , \46583 , \46584 , \46585 , \46586 ,
         \46587 , \46588 , \46589 , \46590 , \46591 , \46592 , \46593 , \46594 , \46595 , \46596 ,
         \46597 , \46598 , \46599 , \46600 , \46601 , \46602 , \46603 , \46604 , \46605 , \46606 ,
         \46607 , \46608 , \46609 , \46610 , \46611 , \46612 , \46613 , \46614 , \46615 , \46616 ,
         \46617 , \46618 , \46619 , \46620 , \46621 , \46622 , \46623 , \46624 , \46625 , \46626 ,
         \46627 , \46628 , \46629 , \46630 , \46631 , \46632 , \46633 , \46634 , \46635 , \46636 ,
         \46637 , \46638 , \46639 , \46640 , \46641 , \46642 , \46643 , \46644 , \46645 , \46646 ,
         \46647 , \46648 , \46649 , \46650 , \46651 , \46652 , \46653 , \46654 , \46655 , \46656 ,
         \46657 , \46658 , \46659 , \46660 , \46661 , \46662 , \46663 , \46664 , \46665 , \46666 ,
         \46667 , \46668 , \46669 , \46670 , \46671 , \46672 , \46673 , \46674 , \46675 , \46676 ,
         \46677 , \46678 , \46679 , \46680 , \46681 , \46682 , \46683 , \46684 , \46685 , \46686 ,
         \46687 , \46688 , \46689 , \46690 , \46691 , \46692 , \46693 , \46694 , \46695 , \46696 ,
         \46697 , \46698 , \46699 , \46700 , \46701 , \46702 , \46703 , \46704 , \46705 , \46706 ,
         \46707 , \46708 , \46709 , \46710 , \46711 , \46712 , \46713 , \46714 , \46715 , \46716 ,
         \46717 , \46718 , \46719 , \46720 , \46721 , \46722 , \46723 , \46724 , \46725 , \46726 ,
         \46727 , \46728 , \46729 , \46730 , \46731 , \46732 , \46733 , \46734 , \46735 , \46736 ,
         \46737 , \46738 , \46739 , \46740 , \46741 , \46742 , \46743 , \46744 , \46745 , \46746 ,
         \46747 , \46748 , \46749 , \46750 , \46751 , \46752 , \46753 , \46754 , \46755 , \46756 ,
         \46757 , \46758 , \46759 , \46760 , \46761 , \46762 , \46763 , \46764 , \46765 , \46766 ,
         \46767 , \46768 , \46769 , \46770 , \46771 , \46772 , \46773 , \46774 , \46775 , \46776 ,
         \46777 , \46778 , \46779 , \46780 , \46781 , \46782 , \46783 , \46784 , \46785 , \46786 ,
         \46787 , \46788 , \46789 , \46790 , \46791 , \46792 , \46793 , \46794 , \46795 , \46796 ,
         \46797 , \46798 , \46799 , \46800 , \46801 , \46802 , \46803 , \46804 , \46805 , \46806 ,
         \46807 , \46808 , \46809 , \46810 , \46811 , \46812 , \46813 , \46814 , \46815 , \46816 ,
         \46817 , \46818 , \46819 , \46820 , \46821 , \46822 , \46823 , \46824 , \46825 , \46826 ,
         \46827 , \46828 , \46829 , \46830 , \46831 , \46832 , \46833 , \46834 , \46835 , \46836 ,
         \46837 , \46838 , \46839 , \46840 , \46841 , \46842 , \46843 , \46844 , \46845 , \46846 ,
         \46847 , \46848 , \46849 , \46850 , \46851 , \46852 , \46853 , \46854 , \46855 , \46856 ,
         \46857 , \46858 , \46859 , \46860 , \46861 , \46862 , \46863 , \46864 , \46865 , \46866 ,
         \46867 , \46868 , \46869 , \46870 , \46871 , \46872 , \46873 , \46874 , \46875 , \46876 ,
         \46877 , \46878 , \46879 , \46880 , \46881 , \46882 , \46883 , \46884 , \46885 , \46886 ,
         \46887 , \46888 , \46889 , \46890 , \46891 , \46892 , \46893 , \46894 , \46895 , \46896 ,
         \46897 , \46898 , \46899 , \46900 , \46901 , \46902 , \46903 , \46904 , \46905 , \46906 ,
         \46907 , \46908 , \46909 , \46910 , \46911 , \46912 , \46913 , \46914 , \46915 , \46916 ,
         \46917 , \46918 , \46919 , \46920 , \46921 , \46922 , \46923 , \46924 , \46925 , \46926 ,
         \46927 , \46928 , \46929 , \46930 , \46931 , \46932 , \46933 , \46934 , \46935 , \46936 ,
         \46937 , \46938 , \46939 , \46940 , \46941 , \46942 , \46943 , \46944 , \46945 , \46946 ,
         \46947 , \46948 , \46949 , \46950 , \46951 , \46952 , \46953 , \46954 , \46955 , \46956 ,
         \46957 , \46958 , \46959 , \46960 , \46961 , \46962 , \46963 , \46964 , \46965 , \46966 ,
         \46967 , \46968 , \46969 , \46970 , \46971 , \46972 , \46973 , \46974 , \46975 , \46976 ,
         \46977 , \46978 , \46979 , \46980 , \46981 , \46982 , \46983 , \46984 , \46985 , \46986 ,
         \46987 , \46988 , \46989 , \46990 , \46991 , \46992 , \46993 , \46994 , \46995 , \46996 ,
         \46997 , \46998 , \46999 , \47000 , \47001 , \47002 , \47003 , \47004 , \47005 , \47006 ,
         \47007 , \47008 , \47009 , \47010 , \47011 , \47012 , \47013 , \47014 , \47015 , \47016 ,
         \47017 , \47018 , \47019 , \47020 , \47021 , \47022 , \47023 , \47024 , \47025 , \47026 ,
         \47027 , \47028 , \47029 , \47030 , \47031 , \47032 , \47033 , \47034 , \47035 , \47036 ,
         \47037 , \47038 , \47039 , \47040 , \47041 , \47042 , \47043 , \47044 , \47045 , \47046 ,
         \47047 , \47048 , \47049 , \47050 , \47051 , \47052 , \47053 , \47054 , \47055 , \47056 ,
         \47057 , \47058 , \47059 , \47060 , \47061 , \47062 , \47063 , \47064 , \47065 , \47066 ,
         \47067 , \47068 , \47069 , \47070 , \47071 , \47072 , \47073 , \47074 , \47075 , \47076 ,
         \47077 , \47078 , \47079 , \47080 , \47081 , \47082 , \47083 , \47084 , \47085 , \47086 ,
         \47087 , \47088 , \47089 , \47090 , \47091 , \47092 , \47093 , \47094 , \47095 , \47096 ,
         \47097 , \47098 , \47099 , \47100 , \47101 , \47102 , \47103 , \47104 , \47105 , \47106 ,
         \47107 , \47108 , \47109 , \47110 , \47111 , \47112 , \47113 , \47114 , \47115 , \47116 ,
         \47117 , \47118 , \47119 , \47120 , \47121 , \47122 , \47123 , \47124 , \47125 , \47126 ,
         \47127 , \47128 , \47129 , \47130 , \47131 , \47132 , \47133 , \47134 , \47135 , \47136 ,
         \47137 , \47138 , \47139 , \47140 , \47141 , \47142 , \47143 , \47144 , \47145 , \47146 ,
         \47147 , \47148 , \47149 , \47150 , \47151 , \47152 , \47153 , \47154 , \47155 , \47156 ,
         \47157 , \47158 , \47159 , \47160 , \47161 , \47162 , \47163 , \47164 , \47165 , \47166 ,
         \47167 , \47168 , \47169 , \47170 , \47171 , \47172 , \47173 , \47174 , \47175 , \47176 ,
         \47177 , \47178 , \47179 , \47180 , \47181 , \47182 , \47183 , \47184 , \47185 , \47186 ,
         \47187 , \47188 , \47189 , \47190 , \47191 , \47192 , \47193 , \47194 , \47195 , \47196 ,
         \47197 , \47198 , \47199 , \47200 , \47201 , \47202 , \47203 , \47204 , \47205 , \47206 ,
         \47207 , \47208 , \47209 , \47210 , \47211 , \47212 , \47213 , \47214 , \47215 , \47216 ,
         \47217 , \47218 , \47219 , \47220 , \47221 , \47222 , \47223 , \47224 , \47225 , \47226 ,
         \47227 , \47228 , \47229 , \47230 , \47231 , \47232 , \47233 , \47234 , \47235 , \47236 ,
         \47237 , \47238 , \47239 , \47240 , \47241 , \47242 , \47243 , \47244 , \47245 , \47246 ,
         \47247 , \47248 , \47249 , \47250 , \47251 , \47252 , \47253 , \47254 , \47255 , \47256 ,
         \47257 , \47258 , \47259 , \47260 , \47261 , \47262 , \47263 , \47264 , \47265 , \47266 ,
         \47267 , \47268 , \47269 , \47270 , \47271 , \47272 , \47273 , \47274 , \47275 , \47276 ,
         \47277 , \47278 , \47279 , \47280 , \47281 , \47282 , \47283 , \47284 , \47285 , \47286 ,
         \47287 , \47288 , \47289 , \47290 , \47291 , \47292 , \47293 , \47294 , \47295 , \47296 ,
         \47297 , \47298 , \47299 , \47300 , \47301 , \47302 , \47303 , \47304 , \47305 , \47306 ,
         \47307 , \47308 , \47309 , \47310 , \47311 , \47312 , \47313 , \47314 , \47315 , \47316 ,
         \47317 , \47318 , \47319 , \47320 , \47321 , \47322 , \47323 , \47324 , \47325 , \47326 ,
         \47327 , \47328 , \47329 , \47330 , \47331 , \47332 , \47333 , \47334 , \47335 , \47336 ,
         \47337 , \47338 , \47339 , \47340 , \47341 , \47342 , \47343 , \47344 , \47345 , \47346 ,
         \47347 , \47348 , \47349 , \47350 , \47351 , \47352 , \47353 , \47354 , \47355 , \47356 ,
         \47357 , \47358 , \47359 , \47360 , \47361 , \47362 , \47363 , \47364 , \47365 , \47366 ,
         \47367 , \47368 , \47369 , \47370 , \47371 , \47372 , \47373 , \47374 , \47375 , \47376 ,
         \47377 , \47378 , \47379 , \47380 , \47381 , \47382 , \47383 , \47384 , \47385 , \47386 ,
         \47387 , \47388 , \47389 , \47390 , \47391 , \47392 , \47393 , \47394 , \47395 , \47396 ,
         \47397 , \47398 , \47399 , \47400 , \47401 , \47402 , \47403 , \47404 , \47405 , \47406 ,
         \47407 , \47408 , \47409 , \47410 , \47411 , \47412 , \47413 , \47414 , \47415 , \47416 ,
         \47417 , \47418 , \47419 , \47420 , \47421 , \47422 , \47423 , \47424 , \47425 , \47426 ,
         \47427 , \47428 , \47429 , \47430 , \47431 , \47432 , \47433 , \47434 , \47435 , \47436 ,
         \47437 , \47438 , \47439 , \47440 , \47441 , \47442 , \47443 , \47444 , \47445 , \47446 ,
         \47447 , \47448 , \47449 , \47450 , \47451 , \47452 , \47453 , \47454 , \47455 , \47456 ,
         \47457 , \47458 , \47459 , \47460 , \47461 , \47462 , \47463 , \47464 , \47465 , \47466 ,
         \47467 , \47468 , \47469 , \47470 , \47471 , \47472 , \47473 , \47474 , \47475 , \47476 ,
         \47477 , \47478 , \47479 , \47480 , \47481 , \47482 , \47483 , \47484 , \47485 , \47486 ,
         \47487 , \47488 , \47489 , \47490 , \47491 , \47492 , \47493 , \47494 , \47495 , \47496 ,
         \47497 , \47498 , \47499 , \47500 , \47501 , \47502 , \47503 , \47504 , \47505 , \47506 ,
         \47507 , \47508 , \47509 , \47510 , \47511 , \47512 , \47513 , \47514 , \47515 , \47516 ,
         \47517 , \47518 , \47519 , \47520 , \47521 , \47522 , \47523 , \47524 , \47525 , \47526 ,
         \47527 , \47528 , \47529 , \47530 , \47531 , \47532 , \47533 , \47534 , \47535 , \47536 ,
         \47537 , \47538 , \47539 , \47540 , \47541 , \47542 , \47543 , \47544 , \47545 , \47546 ,
         \47547 , \47548 , \47549 , \47550 , \47551 , \47552 , \47553 , \47554 , \47555 , \47556 ,
         \47557 , \47558 , \47559 , \47560 , \47561 , \47562 , \47563 , \47564 , \47565 , \47566 ,
         \47567 , \47568 , \47569 , \47570 , \47571 , \47572 , \47573 , \47574 , \47575 , \47576 ,
         \47577 , \47578 , \47579 , \47580 , \47581 , \47582 , \47583 , \47584 , \47585 , \47586 ,
         \47587 , \47588 , \47589 , \47590 , \47591 , \47592 , \47593 , \47594 , \47595 , \47596 ,
         \47597 , \47598 , \47599 , \47600 , \47601 , \47602 , \47603 , \47604 , \47605 , \47606 ,
         \47607 , \47608 , \47609 , \47610 , \47611 , \47612 , \47613 , \47614 , \47615 , \47616 ,
         \47617 , \47618 , \47619 , \47620 , \47621 , \47622 , \47623 , \47624 , \47625 , \47626 ,
         \47627 , \47628 , \47629 , \47630 , \47631 , \47632 , \47633 , \47634 , \47635 , \47636 ,
         \47637 , \47638 , \47639 , \47640 , \47641 , \47642 , \47643 , \47644 , \47645 , \47646 ,
         \47647 , \47648 , \47649 , \47650 , \47651 , \47652 , \47653 , \47654 , \47655 , \47656 ,
         \47657 , \47658 , \47659 , \47660 , \47661 , \47662 , \47663 , \47664 , \47665 , \47666 ,
         \47667 , \47668 , \47669 , \47670 , \47671 , \47672 , \47673 , \47674 , \47675 , \47676 ,
         \47677 , \47678 , \47679 , \47680 , \47681 , \47682 , \47683 , \47684 , \47685 , \47686 ,
         \47687 , \47688 , \47689 , \47690 , \47691 , \47692 , \47693 , \47694 , \47695 , \47696 ,
         \47697 , \47698 , \47699 , \47700 , \47701 , \47702 , \47703 , \47704 , \47705 , \47706 ,
         \47707 , \47708 , \47709 , \47710 , \47711 , \47712 , \47713 , \47714 , \47715 , \47716 ,
         \47717 , \47718 , \47719 , \47720 , \47721 , \47722 , \47723 , \47724 , \47725 , \47726 ,
         \47727 , \47728 , \47729 , \47730 , \47731 , \47732 , \47733 , \47734 , \47735 , \47736 ,
         \47737 , \47738 , \47739 , \47740 , \47741 , \47742 , \47743 , \47744 , \47745 , \47746 ,
         \47747 , \47748 , \47749 , \47750 , \47751 , \47752 , \47753 , \47754 , \47755 , \47756 ,
         \47757 , \47758 , \47759 , \47760 , \47761 , \47762 , \47763 , \47764 , \47765 , \47766 ,
         \47767 , \47768 , \47769 , \47770 , \47771 , \47772 , \47773 , \47774 , \47775 , \47776 ,
         \47777 , \47778 , \47779 , \47780 , \47781 , \47782 , \47783 , \47784 , \47785 , \47786 ,
         \47787 , \47788 , \47789 , \47790 , \47791 , \47792 , \47793 , \47794 , \47795 , \47796 ,
         \47797 , \47798 , \47799 , \47800 , \47801 , \47802 , \47803 , \47804 , \47805 , \47806 ,
         \47807 , \47808 , \47809 , \47810 , \47811 , \47812 , \47813 , \47814 , \47815 , \47816 ,
         \47817 , \47818 , \47819 , \47820 , \47821 , \47822 , \47823 , \47824 , \47825 , \47826 ,
         \47827 , \47828 , \47829 , \47830 , \47831 , \47832 , \47833 , \47834 , \47835 , \47836 ,
         \47837 , \47838 , \47839 , \47840 , \47841 , \47842 , \47843 , \47844 , \47845 , \47846 ,
         \47847 , \47848 , \47849 , \47850 , \47851 , \47852 , \47853 , \47854 , \47855 , \47856 ,
         \47857 , \47858 , \47859 , \47860 , \47861 , \47862 , \47863 , \47864 , \47865 , \47866 ,
         \47867 , \47868 , \47869 , \47870 , \47871 , \47872 , \47873 , \47874 , \47875 , \47876 ,
         \47877 , \47878 , \47879 , \47880 , \47881 , \47882 , \47883 , \47884 , \47885 , \47886 ,
         \47887 , \47888 , \47889 , \47890 , \47891 , \47892 , \47893 , \47894 , \47895 , \47896 ,
         \47897 , \47898 , \47899 , \47900 , \47901 , \47902 , \47903 , \47904 , \47905 , \47906 ,
         \47907 , \47908 , \47909 , \47910 , \47911 , \47912 , \47913 , \47914 , \47915 , \47916 ,
         \47917 , \47918 , \47919 , \47920 , \47921 , \47922 , \47923 , \47924 , \47925 , \47926 ,
         \47927 , \47928 , \47929 , \47930 , \47931 , \47932 , \47933 , \47934 , \47935 , \47936 ,
         \47937 , \47938 , \47939 , \47940 , \47941 , \47942 , \47943 , \47944 , \47945 , \47946 ,
         \47947 , \47948 , \47949 , \47950 , \47951 , \47952 , \47953 , \47954 , \47955 , \47956 ,
         \47957 , \47958 , \47959 , \47960 , \47961 , \47962 , \47963 , \47964 , \47965 , \47966 ,
         \47967 , \47968 , \47969 , \47970 , \47971 , \47972 , \47973 , \47974 , \47975 , \47976 ,
         \47977 , \47978 , \47979 , \47980 , \47981 , \47982 , \47983 , \47984 , \47985 , \47986 ,
         \47987 , \47988 , \47989 , \47990 , \47991 , \47992 , \47993 , \47994 , \47995 , \47996 ,
         \47997 , \47998 , \47999 , \48000 , \48001 , \48002 , \48003 , \48004 , \48005 , \48006 ,
         \48007 , \48008 , \48009 , \48010 , \48011 , \48012 , \48013 , \48014 , \48015 , \48016 ,
         \48017 , \48018 , \48019 , \48020 , \48021 , \48022 , \48023 , \48024 , \48025 , \48026 ,
         \48027 , \48028 , \48029 , \48030 , \48031 , \48032 , \48033 , \48034 , \48035 , \48036 ,
         \48037 , \48038 , \48039 , \48040 , \48041 , \48042 , \48043 , \48044 , \48045 , \48046 ,
         \48047 , \48048 , \48049 , \48050 , \48051 , \48052 , \48053 , \48054 , \48055 , \48056 ,
         \48057 , \48058 , \48059 , \48060 , \48061 , \48062 , \48063 , \48064 , \48065 , \48066 ,
         \48067 , \48068 , \48069 , \48070 , \48071 , \48072 , \48073 , \48074 , \48075 , \48076 ,
         \48077 , \48078 , \48079 , \48080 , \48081 , \48082 , \48083 , \48084 , \48085 , \48086 ,
         \48087 , \48088 , \48089 , \48090 , \48091 , \48092 , \48093 , \48094 , \48095 , \48096 ,
         \48097 , \48098 , \48099 , \48100 , \48101 , \48102 , \48103 , \48104 , \48105 , \48106 ,
         \48107 , \48108 , \48109 , \48110 , \48111 , \48112 , \48113 , \48114 , \48115 , \48116 ,
         \48117 , \48118 , \48119 , \48120 , \48121 , \48122 , \48123 , \48124 , \48125 , \48126 ,
         \48127 , \48128 , \48129 , \48130 , \48131 , \48132 , \48133 , \48134 , \48135 , \48136 ,
         \48137 , \48138 , \48139 , \48140 , \48141 , \48142 , \48143 , \48144 , \48145 , \48146 ,
         \48147 , \48148 , \48149 , \48150 , \48151 , \48152 , \48153 , \48154 , \48155 , \48156 ,
         \48157 , \48158 , \48159 , \48160 , \48161 , \48162 , \48163 , \48164 , \48165 , \48166 ,
         \48167 , \48168 , \48169 , \48170 , \48171 , \48172 , \48173 , \48174 , \48175 , \48176 ,
         \48177 , \48178 , \48179 , \48180 , \48181 , \48182 , \48183 , \48184 , \48185 , \48186 ,
         \48187 , \48188 , \48189 , \48190 , \48191 , \48192 , \48193 , \48194 , \48195 , \48196 ,
         \48197 , \48198 , \48199 , \48200 , \48201 , \48202 , \48203 , \48204 , \48205 , \48206 ,
         \48207 , \48208 , \48209 , \48210 , \48211 , \48212 , \48213 , \48214 , \48215 , \48216 ,
         \48217 , \48218 , \48219 , \48220 , \48221 , \48222 , \48223 , \48224 , \48225 , \48226 ,
         \48227 , \48228 , \48229 , \48230 , \48231 , \48232 , \48233 , \48234 , \48235 , \48236 ,
         \48237 , \48238 , \48239 , \48240 , \48241 , \48242 , \48243 , \48244 , \48245 , \48246 ,
         \48247 , \48248 , \48249 , \48250 , \48251 , \48252 , \48253 , \48254 , \48255 , \48256 ,
         \48257 , \48258 , \48259 , \48260 , \48261 , \48262 , \48263 , \48264 , \48265 , \48266 ,
         \48267 , \48268 , \48269 , \48270 , \48271 , \48272 , \48273 , \48274 , \48275 , \48276 ,
         \48277 , \48278 , \48279 , \48280 , \48281 , \48282 , \48283 , \48284 , \48285 , \48286 ,
         \48287 , \48288 , \48289 , \48290 , \48291 , \48292 , \48293 , \48294 , \48295 , \48296 ,
         \48297 , \48298 , \48299 , \48300 , \48301 , \48302 , \48303 , \48304 , \48305 , \48306 ,
         \48307 , \48308 , \48309 , \48310 , \48311 , \48312 , \48313 , \48314 , \48315 , \48316 ,
         \48317 , \48318 , \48319 , \48320 , \48321 , \48322 , \48323 , \48324 , \48325 , \48326 ,
         \48327 , \48328 , \48329 , \48330 , \48331 , \48332 , \48333 , \48334 , \48335 , \48336 ,
         \48337 , \48338 , \48339 , \48340 , \48341 , \48342 , \48343 , \48344 , \48345 , \48346 ,
         \48347 , \48348 , \48349 , \48350 , \48351 , \48352 , \48353 , \48354 , \48355 , \48356 ,
         \48357 , \48358 , \48359 , \48360 , \48361 , \48362 , \48363 , \48364 , \48365 , \48366 ,
         \48367 , \48368 , \48369 , \48370 , \48371 , \48372 , \48373 , \48374 , \48375 , \48376 ,
         \48377 , \48378 , \48379 , \48380 , \48381 , \48382 , \48383 , \48384 , \48385 , \48386 ,
         \48387 , \48388 , \48389 , \48390 , \48391 , \48392 , \48393 , \48394 , \48395 , \48396 ,
         \48397 , \48398 , \48399 , \48400 , \48401 , \48402 , \48403 , \48404 , \48405 , \48406 ,
         \48407 , \48408 , \48409 , \48410 , \48411 , \48412 , \48413 , \48414 , \48415 , \48416 ,
         \48417 , \48418 , \48419 , \48420 , \48421 , \48422 , \48423 , \48424 , \48425 , \48426 ,
         \48427 , \48428 , \48429 , \48430 , \48431 , \48432 , \48433 , \48434 , \48435 , \48436 ,
         \48437 , \48438 , \48439 , \48440 , \48441 , \48442 , \48443 , \48444 , \48445 , \48446 ,
         \48447 , \48448 , \48449 , \48450 , \48451 , \48452 , \48453 , \48454 , \48455 , \48456 ,
         \48457 , \48458 , \48459 , \48460 , \48461 , \48462 , \48463 , \48464 , \48465 , \48466 ,
         \48467 , \48468 , \48469 , \48470 , \48471 , \48472 , \48473 , \48474 , \48475 , \48476 ,
         \48477 , \48478 , \48479 , \48480 , \48481 , \48482 , \48483 , \48484 , \48485 , \48486 ,
         \48487 , \48488 , \48489 , \48490 , \48491 , \48492 , \48493 , \48494 , \48495 , \48496 ,
         \48497 , \48498 , \48499 , \48500 , \48501 , \48502 , \48503 , \48504 , \48505 , \48506 ,
         \48507 , \48508 , \48509 , \48510 , \48511 , \48512 , \48513 , \48514 , \48515 , \48516 ,
         \48517 , \48518 , \48519 , \48520 , \48521 , \48522 , \48523 , \48524 , \48525 , \48526 ,
         \48527 , \48528 , \48529 , \48530 , \48531 , \48532 , \48533 , \48534 , \48535 , \48536 ,
         \48537 , \48538 , \48539 , \48540 , \48541 , \48542 , \48543 , \48544 , \48545 , \48546 ,
         \48547 , \48548 , \48549 , \48550 , \48551 , \48552 , \48553 , \48554 , \48555 , \48556 ,
         \48557 , \48558 , \48559 , \48560 , \48561 , \48562 , \48563 , \48564 , \48565 , \48566 ,
         \48567 , \48568 , \48569 , \48570 , \48571 , \48572 , \48573 , \48574 , \48575 , \48576 ,
         \48577 , \48578 , \48579 , \48580 , \48581 , \48582 , \48583 , \48584 , \48585 , \48586 ,
         \48587 , \48588 , \48589 , \48590 , \48591 , \48592 , \48593 , \48594 , \48595 , \48596 ,
         \48597 , \48598 , \48599 , \48600 , \48601 , \48602 , \48603 , \48604 , \48605 , \48606 ,
         \48607 , \48608 , \48609 , \48610 , \48611 , \48612 , \48613 , \48614 , \48615 , \48616 ,
         \48617 , \48618 , \48619 , \48620 , \48621 , \48622 , \48623 , \48624 , \48625 , \48626 ,
         \48627 , \48628 , \48629 , \48630 , \48631 , \48632 , \48633 , \48634 , \48635 , \48636 ,
         \48637 , \48638 , \48639 , \48640 , \48641 , \48642 , \48643 , \48644 , \48645 , \48646 ,
         \48647 , \48648 , \48649 , \48650 , \48651 , \48652 , \48653 , \48654 , \48655 , \48656 ,
         \48657 , \48658 , \48659 , \48660 , \48661 , \48662 , \48663 , \48664 , \48665 , \48666 ,
         \48667 , \48668 , \48669 , \48670 , \48671 , \48672 , \48673 , \48674 , \48675 , \48676 ,
         \48677 , \48678 , \48679 , \48680 , \48681 , \48682 , \48683 , \48684 , \48685 , \48686 ,
         \48687 , \48688 , \48689 , \48690 , \48691 , \48692 , \48693 , \48694 , \48695 , \48696 ,
         \48697 , \48698 , \48699 , \48700 , \48701 , \48702 , \48703 , \48704 , \48705 , \48706 ,
         \48707 , \48708 , \48709 , \48710 , \48711 , \48712 , \48713 , \48714 , \48715 , \48716 ,
         \48717 , \48718 , \48719 , \48720 , \48721 , \48722 , \48723 , \48724 , \48725 , \48726 ,
         \48727 , \48728 , \48729 , \48730 , \48731 , \48732 , \48733 , \48734 , \48735 , \48736 ,
         \48737 , \48738 , \48739 , \48740 , \48741 , \48742 , \48743 , \48744 , \48745 , \48746 ,
         \48747 , \48748 , \48749 , \48750 , \48751 , \48752 , \48753 , \48754 , \48755 , \48756 ,
         \48757 , \48758 , \48759 , \48760 , \48761 , \48762 , \48763 , \48764 , \48765 , \48766 ,
         \48767 , \48768 , \48769 , \48770 , \48771 , \48772 , \48773 , \48774 , \48775 , \48776 ,
         \48777 , \48778 , \48779 , \48780 , \48781 , \48782 , \48783 , \48784 , \48785 , \48786 ,
         \48787 , \48788 , \48789 , \48790 , \48791 , \48792 , \48793 , \48794 , \48795 , \48796 ,
         \48797 , \48798 , \48799 , \48800 , \48801 , \48802 , \48803 , \48804 , \48805 , \48806 ,
         \48807 , \48808 , \48809 , \48810 , \48811 , \48812 , \48813 , \48814 , \48815 , \48816 ,
         \48817 , \48818 , \48819 , \48820 , \48821 , \48822 , \48823 , \48824 , \48825 , \48826 ,
         \48827 , \48828 , \48829 , \48830 , \48831 , \48832 , \48833 , \48834 , \48835 , \48836 ,
         \48837 , \48838 , \48839 , \48840 , \48841 , \48842 , \48843 , \48844 , \48845 , \48846 ,
         \48847 , \48848 , \48849 , \48850 , \48851 , \48852 , \48853 , \48854 , \48855 , \48856 ,
         \48857 , \48858 , \48859 , \48860 , \48861 , \48862 , \48863 , \48864 , \48865 , \48866 ,
         \48867 , \48868 , \48869 , \48870 , \48871 , \48872 , \48873 , \48874 , \48875 , \48876 ,
         \48877 , \48878 , \48879 , \48880 , \48881 , \48882 , \48883 , \48884 , \48885 , \48886 ,
         \48887 , \48888 , \48889 , \48890 , \48891 , \48892 , \48893 , \48894 , \48895 , \48896 ,
         \48897 , \48898 , \48899 , \48900 , \48901 , \48902 , \48903 , \48904 , \48905 , \48906 ,
         \48907 , \48908 , \48909 , \48910 , \48911 , \48912 , \48913 , \48914 , \48915 , \48916 ,
         \48917 , \48918 , \48919 , \48920 , \48921 , \48922 , \48923 , \48924 , \48925 , \48926 ,
         \48927 , \48928 , \48929 , \48930 , \48931 , \48932 , \48933 , \48934 , \48935 , \48936 ,
         \48937 , \48938 , \48939 , \48940 , \48941 , \48942 , \48943 , \48944 , \48945 , \48946 ,
         \48947 , \48948 , \48949 , \48950 , \48951 , \48952 , \48953 , \48954 , \48955 , \48956 ,
         \48957 , \48958 , \48959 , \48960 , \48961 , \48962 , \48963 , \48964 , \48965 , \48966 ,
         \48967 , \48968 , \48969 , \48970 , \48971 , \48972 , \48973 , \48974 , \48975 , \48976 ,
         \48977 , \48978 , \48979 , \48980 , \48981 , \48982 , \48983 , \48984 , \48985 , \48986 ,
         \48987 , \48988 , \48989 , \48990 , \48991 , \48992 , \48993 , \48994 , \48995 , \48996 ,
         \48997 , \48998 , \48999 , \49000 , \49001 , \49002 , \49003 , \49004 , \49005 , \49006 ,
         \49007 , \49008 , \49009 , \49010 , \49011 , \49012 , \49013 , \49014 , \49015 , \49016 ,
         \49017 , \49018 , \49019 , \49020 , \49021 , \49022 , \49023 , \49024 , \49025 , \49026 ,
         \49027 , \49028 , \49029 , \49030 , \49031 , \49032 , \49033 , \49034 , \49035 , \49036 ,
         \49037 , \49038 , \49039 , \49040 , \49041 , \49042 , \49043 , \49044 , \49045 , \49046 ,
         \49047 , \49048 , \49049 , \49050 , \49051 , \49052 , \49053 , \49054 , \49055 , \49056 ,
         \49057 , \49058 , \49059 , \49060 , \49061 , \49062 , \49063 , \49064 , \49065 , \49066 ,
         \49067 , \49068 , \49069 , \49070 , \49071 , \49072 , \49073 , \49074 , \49075 , \49076 ,
         \49077 , \49078 , \49079 , \49080 , \49081 , \49082 , \49083 , \49084 , \49085 , \49086 ,
         \49087 , \49088 , \49089 , \49090 , \49091 , \49092 , \49093 , \49094 , \49095 , \49096 ,
         \49097 , \49098 , \49099 , \49100 , \49101 , \49102 , \49103 , \49104 , \49105 , \49106 ,
         \49107 , \49108 , \49109 , \49110 , \49111 , \49112 , \49113 , \49114 , \49115 , \49116 ,
         \49117 , \49118 , \49119 , \49120 , \49121 , \49122 , \49123 , \49124 , \49125 , \49126 ,
         \49127 , \49128 , \49129 , \49130 , \49131 , \49132 , \49133 , \49134 , \49135 , \49136 ,
         \49137 , \49138 , \49139 , \49140 , \49141 , \49142 , \49143 , \49144 , \49145 , \49146 ,
         \49147 , \49148 , \49149 , \49150 , \49151 , \49152 , \49153 , \49154 , \49155 , \49156 ,
         \49157 , \49158 , \49159 , \49160 , \49161 , \49162 , \49163 , \49164 , \49165 , \49166 ,
         \49167 , \49168 , \49169 , \49170 , \49171 , \49172 , \49173 , \49174 , \49175 , \49176 ,
         \49177 , \49178 , \49179 , \49180 , \49181 , \49182 , \49183 , \49184 , \49185 , \49186 ,
         \49187 , \49188 , \49189 , \49190 , \49191 , \49192 , \49193 , \49194 , \49195 , \49196 ,
         \49197 , \49198 , \49199 , \49200 , \49201 , \49202 , \49203 , \49204 , \49205 , \49206 ,
         \49207 , \49208 , \49209 , \49210 , \49211 , \49212 , \49213 , \49214 , \49215 , \49216 ,
         \49217 , \49218 , \49219 , \49220 , \49221 , \49222 , \49223 , \49224 , \49225 , \49226 ,
         \49227 , \49228 , \49229 , \49230 , \49231 , \49232 , \49233 , \49234 , \49235 , \49236 ,
         \49237 , \49238 , \49239 , \49240 , \49241 , \49242 , \49243 , \49244 , \49245 , \49246 ,
         \49247 , \49248 , \49249 , \49250 , \49251 , \49252 , \49253 , \49254 , \49255 , \49256 ,
         \49257 , \49258 , \49259 , \49260 , \49261 , \49262 , \49263 , \49264 , \49265 , \49266 ,
         \49267 , \49268 , \49269 , \49270 , \49271 , \49272 , \49273 , \49274 , \49275 , \49276 ,
         \49277 , \49278 , \49279 , \49280 , \49281 , \49282 , \49283 , \49284 , \49285 , \49286 ,
         \49287 , \49288 , \49289 , \49290 , \49291 , \49292 , \49293 , \49294 , \49295 , \49296 ,
         \49297 , \49298 , \49299 , \49300 , \49301 , \49302 , \49303 , \49304 , \49305 , \49306 ,
         \49307 , \49308 , \49309 , \49310 , \49311 , \49312 , \49313 , \49314 , \49315 , \49316 ,
         \49317 , \49318 , \49319 , \49320 , \49321 , \49322 , \49323 , \49324 , \49325 , \49326 ,
         \49327 , \49328 , \49329 , \49330 , \49331 , \49332 , \49333 , \49334 , \49335 , \49336 ,
         \49337 , \49338 , \49339 , \49340 , \49341 , \49342 , \49343 , \49344 , \49345 , \49346 ,
         \49347 , \49348 , \49349 , \49350 , \49351 , \49352 , \49353 , \49354 , \49355 , \49356 ,
         \49357 , \49358 , \49359 , \49360 , \49361 , \49362 , \49363 , \49364 , \49365 , \49366 ,
         \49367 , \49368 , \49369 , \49370 , \49371 , \49372 , \49373 , \49374 , \49375 , \49376 ,
         \49377 , \49378 , \49379 , \49380 , \49381 , \49382 , \49383 , \49384 , \49385 , \49386 ,
         \49387 , \49388 , \49389 , \49390 , \49391 , \49392 , \49393 , \49394 , \49395 , \49396 ,
         \49397 , \49398 , \49399 , \49400 , \49401 , \49402 , \49403 , \49404 , \49405 , \49406 ,
         \49407 , \49408 , \49409 , \49410 , \49411 , \49412 , \49413 , \49414 , \49415 , \49416 ,
         \49417 , \49418 , \49419 , \49420 , \49421 , \49422 , \49423 , \49424 , \49425 , \49426 ,
         \49427 , \49428 , \49429 , \49430 , \49431 , \49432 , \49433 , \49434 , \49435 , \49436 ,
         \49437 , \49438 , \49439 , \49440 , \49441 , \49442 , \49443 , \49444 , \49445 , \49446 ,
         \49447 , \49448 , \49449 , \49450 , \49451 , \49452 , \49453 , \49454 , \49455 , \49456 ,
         \49457 , \49458 , \49459 , \49460 , \49461 , \49462 , \49463 , \49464 , \49465 , \49466 ,
         \49467 , \49468 , \49469 , \49470 , \49471 , \49472 , \49473 , \49474 , \49475 , \49476 ,
         \49477 , \49478 , \49479 , \49480 , \49481 , \49482 , \49483 , \49484 , \49485 , \49486 ,
         \49487 , \49488 , \49489 , \49490 , \49491 , \49492 , \49493 , \49494 , \49495 , \49496 ,
         \49497 , \49498 , \49499 , \49500 , \49501 , \49502 , \49503 , \49504 , \49505 , \49506 ,
         \49507 , \49508 , \49509 , \49510 , \49511 , \49512 , \49513 , \49514 , \49515 , \49516 ,
         \49517 , \49518 , \49519 , \49520 , \49521 , \49522 , \49523 , \49524 , \49525 , \49526 ,
         \49527 , \49528 , \49529 , \49530 , \49531 , \49532 , \49533 , \49534 , \49535 , \49536 ,
         \49537 , \49538 , \49539 , \49540 , \49541 , \49542 , \49543 , \49544 , \49545 , \49546 ,
         \49547 , \49548 , \49549 , \49550 , \49551 , \49552 , \49553 , \49554 , \49555 , \49556 ,
         \49557 , \49558 , \49559 , \49560 , \49561 , \49562 , \49563 , \49564 , \49565 , \49566 ,
         \49567 , \49568 , \49569 , \49570 , \49571 , \49572 , \49573 , \49574 , \49575 , \49576 ,
         \49577 , \49578 , \49579 , \49580 , \49581 , \49582 , \49583 , \49584 , \49585 , \49586 ,
         \49587 , \49588 , \49589 , \49590 , \49591 , \49592 , \49593 , \49594 , \49595 , \49596 ,
         \49597 , \49598 , \49599 , \49600 , \49601 , \49602 , \49603 , \49604 , \49605 , \49606 ,
         \49607 , \49608 , \49609 , \49610 , \49611 , \49612 , \49613 , \49614 , \49615 , \49616 ,
         \49617 , \49618 , \49619 , \49620 , \49621 , \49622 , \49623 , \49624 , \49625 , \49626 ,
         \49627 , \49628 , \49629 , \49630 , \49631 , \49632 , \49633 , \49634 , \49635 , \49636 ,
         \49637 , \49638 , \49639 , \49640 , \49641 , \49642 , \49643 , \49644 , \49645 , \49646 ,
         \49647 , \49648 , \49649 , \49650 , \49651 , \49652 , \49653 , \49654 , \49655 , \49656 ,
         \49657 , \49658 , \49659 , \49660 , \49661 , \49662 , \49663 , \49664 , \49665 , \49666 ,
         \49667 , \49668 , \49669 , \49670 , \49671 , \49672 , \49673 , \49674 , \49675 , \49676 ,
         \49677 , \49678 , \49679 , \49680 , \49681 , \49682 , \49683 , \49684 , \49685 , \49686 ,
         \49687 , \49688 , \49689 , \49690 , \49691 , \49692 , \49693 , \49694 , \49695 , \49696 ,
         \49697 , \49698 , \49699 , \49700 , \49701 , \49702 , \49703 , \49704 , \49705 , \49706 ,
         \49707 , \49708 , \49709 , \49710 , \49711 , \49712 , \49713 , \49714 , \49715 , \49716 ,
         \49717 , \49718 , \49719 , \49720 , \49721 , \49722 , \49723 , \49724 , \49725 , \49726 ,
         \49727 , \49728 , \49729 , \49730 , \49731 , \49732 , \49733 , \49734 , \49735 , \49736 ,
         \49737 , \49738 , \49739 , \49740 , \49741 , \49742 , \49743 , \49744 , \49745 , \49746 ,
         \49747 , \49748 , \49749 , \49750 , \49751 , \49752 , \49753 , \49754 , \49755 , \49756 ,
         \49757 , \49758 , \49759 , \49760 , \49761 , \49762 , \49763 , \49764 , \49765 , \49766 ,
         \49767 , \49768 , \49769 , \49770 , \49771 , \49772 , \49773 , \49774 , \49775 , \49776 ,
         \49777 , \49778 , \49779 , \49780 , \49781 , \49782 , \49783 , \49784 , \49785 , \49786 ,
         \49787 , \49788 , \49789 , \49790 , \49791 , \49792 , \49793 , \49794 , \49795 , \49796 ,
         \49797 , \49798 , \49799 , \49800 , \49801 , \49802 , \49803 , \49804 , \49805 , \49806 ,
         \49807 , \49808 , \49809 , \49810 , \49811 , \49812 , \49813 , \49814 , \49815 , \49816 ,
         \49817 , \49818 , \49819 , \49820 , \49821 , \49822 , \49823 , \49824 , \49825 , \49826 ,
         \49827 , \49828 , \49829 , \49830 , \49831 , \49832 , \49833 , \49834 , \49835 , \49836 ,
         \49837 , \49838 , \49839 , \49840 , \49841 , \49842 , \49843 , \49844 , \49845 , \49846 ,
         \49847 , \49848 , \49849 , \49850 , \49851 , \49852 , \49853 , \49854 , \49855 , \49856 ,
         \49857 , \49858 , \49859 , \49860 , \49861 , \49862 , \49863 , \49864 , \49865 , \49866 ,
         \49867 , \49868 , \49869 , \49870 , \49871 , \49872 , \49873 , \49874 , \49875 , \49876 ,
         \49877 , \49878 , \49879 , \49880 , \49881 , \49882 , \49883 , \49884 , \49885 , \49886 ,
         \49887 , \49888 , \49889 , \49890 , \49891 , \49892 , \49893 , \49894 , \49895 , \49896 ,
         \49897 , \49898 , \49899 , \49900 , \49901 , \49902 , \49903 , \49904 , \49905 , \49906 ,
         \49907 , \49908 , \49909 , \49910 , \49911 , \49912 , \49913 , \49914 , \49915 , \49916 ,
         \49917 , \49918 , \49919 , \49920 , \49921 , \49922 , \49923 , \49924 , \49925 , \49926 ,
         \49927 , \49928 , \49929 , \49930 , \49931 , \49932 , \49933 , \49934 , \49935 , \49936 ,
         \49937 , \49938 , \49939 , \49940 , \49941 , \49942 , \49943 , \49944 , \49945 , \49946 ,
         \49947 , \49948 , \49949 , \49950 , \49951 , \49952 , \49953 , \49954 , \49955 , \49956 ,
         \49957 , \49958 , \49959 , \49960 , \49961 , \49962 , \49963 , \49964 , \49965 , \49966 ,
         \49967 , \49968 , \49969 , \49970 , \49971 , \49972 , \49973 , \49974 , \49975 , \49976 ,
         \49977 , \49978 , \49979 , \49980 , \49981 , \49982 , \49983 , \49984 , \49985 , \49986 ,
         \49987 , \49988 , \49989 , \49990 , \49991 , \49992 , \49993 , \49994 , \49995 , \49996 ,
         \49997 , \49998 , \49999 , \50000 , \50001 , \50002 , \50003 , \50004 , \50005 , \50006 ,
         \50007 , \50008 , \50009 , \50010 , \50011 , \50012 , \50013 , \50014 , \50015 , \50016 ,
         \50017 , \50018 , \50019 , \50020 , \50021 , \50022 , \50023 , \50024 , \50025 , \50026 ,
         \50027 , \50028 , \50029 , \50030 , \50031 , \50032 , \50033 , \50034 , \50035 , \50036 ,
         \50037 , \50038 , \50039 , \50040 , \50041 , \50042 , \50043 , \50044 , \50045 , \50046 ,
         \50047 , \50048 , \50049 , \50050 , \50051 , \50052 , \50053 , \50054 , \50055 , \50056 ,
         \50057 , \50058 , \50059 , \50060 , \50061 , \50062 , \50063 , \50064 , \50065 , \50066 ,
         \50067 , \50068 , \50069 , \50070 , \50071 , \50072 , \50073 , \50074 , \50075 , \50076 ,
         \50077 , \50078 , \50079 , \50080 , \50081 , \50082 , \50083 , \50084 , \50085 , \50086 ,
         \50087 , \50088 , \50089 , \50090 , \50091 , \50092 , \50093 , \50094 , \50095 , \50096 ,
         \50097 , \50098 , \50099 , \50100 , \50101 , \50102 , \50103 , \50104 , \50105 , \50106 ,
         \50107 , \50108 , \50109 , \50110 , \50111 , \50112 , \50113 , \50114 , \50115 , \50116 ,
         \50117 , \50118 , \50119 , \50120 , \50121 , \50122 , \50123 , \50124 , \50125 , \50126 ,
         \50127 , \50128 , \50129 , \50130 , \50131 , \50132 , \50133 , \50134 , \50135 , \50136 ,
         \50137 , \50138 , \50139 , \50140 , \50141 , \50142 , \50143 , \50144 , \50145 , \50146 ,
         \50147 , \50148 , \50149 , \50150 , \50151 , \50152 , \50153 , \50154 , \50155 , \50156 ,
         \50157 , \50158 , \50159 , \50160 , \50161 , \50162 , \50163 , \50164 , \50165 , \50166 ,
         \50167 , \50168 , \50169 , \50170 , \50171 , \50172 , \50173 , \50174 , \50175 , \50176 ,
         \50177 , \50178 , \50179 , \50180 , \50181 , \50182 , \50183 , \50184 , \50185 , \50186 ,
         \50187 , \50188 , \50189 , \50190 , \50191 , \50192 , \50193 , \50194 , \50195 , \50196 ,
         \50197 , \50198 , \50199 , \50200 , \50201 , \50202 , \50203 , \50204 , \50205 , \50206 ,
         \50207 , \50208 , \50209 , \50210 , \50211 , \50212 , \50213 , \50214 , \50215 , \50216 ,
         \50217 , \50218 , \50219 , \50220 , \50221 , \50222 , \50223 , \50224 , \50225 , \50226 ,
         \50227 , \50228 , \50229 , \50230 , \50231 , \50232 , \50233 , \50234 , \50235 , \50236 ,
         \50237 , \50238 , \50239 , \50240 , \50241 , \50242 , \50243 , \50244 , \50245 , \50246 ,
         \50247 , \50248 , \50249 , \50250 , \50251 , \50252 , \50253 , \50254 , \50255 , \50256 ,
         \50257 , \50258 , \50259 , \50260 , \50261 , \50262 , \50263 , \50264 , \50265 , \50266 ,
         \50267 , \50268 , \50269 , \50270 , \50271 , \50272 , \50273 , \50274 , \50275 , \50276 ,
         \50277 , \50278 , \50279 , \50280 , \50281 , \50282 , \50283 , \50284 , \50285 , \50286 ,
         \50287 , \50288 , \50289 , \50290 , \50291 , \50292 , \50293 , \50294 , \50295 , \50296 ,
         \50297 , \50298 , \50299 , \50300 , \50301 , \50302 , \50303 , \50304 , \50305 , \50306 ,
         \50307 , \50308 , \50309 , \50310 , \50311 , \50312 , \50313 , \50314 , \50315 , \50316 ,
         \50317 , \50318 , \50319 , \50320 , \50321 , \50322 , \50323 , \50324 , \50325 , \50326 ,
         \50327 , \50328 , \50329 , \50330 , \50331 , \50332 , \50333 , \50334 , \50335 , \50336 ,
         \50337 , \50338 , \50339 , \50340 , \50341 , \50342 , \50343 , \50344 , \50345 , \50346 ,
         \50347 , \50348 , \50349 , \50350 , \50351 , \50352 , \50353 , \50354 , \50355 , \50356 ,
         \50357 , \50358 , \50359 , \50360 , \50361 , \50362 , \50363 , \50364 , \50365 , \50366 ,
         \50367 , \50368 , \50369 , \50370 , \50371 , \50372 , \50373 , \50374 , \50375 , \50376 ,
         \50377 , \50378 , \50379 , \50380 , \50381 , \50382 , \50383 , \50384 , \50385 , \50386 ,
         \50387 , \50388 , \50389 , \50390 , \50391 , \50392 , \50393 , \50394 , \50395 , \50396 ,
         \50397 , \50398 , \50399 , \50400 , \50401 , \50402 , \50403 , \50404 , \50405 , \50406 ,
         \50407 , \50408 , \50409 , \50410 , \50411 , \50412 , \50413 , \50414 , \50415 , \50416 ,
         \50417 , \50418 , \50419 , \50420 , \50421 , \50422 , \50423 , \50424 , \50425 , \50426 ,
         \50427 , \50428 , \50429 , \50430 , \50431 , \50432 , \50433 , \50434 , \50435 , \50436 ,
         \50437 , \50438 , \50439 , \50440 , \50441 , \50442 , \50443 , \50444 , \50445 , \50446 ,
         \50447 , \50448 , \50449 , \50450 , \50451 , \50452 , \50453 , \50454 , \50455 , \50456 ,
         \50457 , \50458 , \50459 , \50460 , \50461 , \50462 , \50463 , \50464 , \50465 , \50466 ,
         \50467 , \50468 , \50469 , \50470 , \50471 , \50472 , \50473 , \50474 , \50475 , \50476 ,
         \50477 , \50478 , \50479 , \50480 , \50481 , \50482 , \50483 , \50484 , \50485 , \50486 ,
         \50487 , \50488 , \50489 , \50490 , \50491 , \50492 , \50493 , \50494 , \50495 , \50496 ,
         \50497 , \50498 , \50499 , \50500 , \50501 , \50502 , \50503 , \50504 , \50505 , \50506 ,
         \50507 , \50508 , \50509 , \50510 , \50511 , \50512 , \50513 , \50514 , \50515 , \50516 ,
         \50517 , \50518 , \50519 , \50520 , \50521 , \50522 , \50523 , \50524 , \50525 , \50526 ,
         \50527 , \50528 , \50529 , \50530 , \50531 , \50532 , \50533 , \50534 , \50535 , \50536 ,
         \50537 , \50538 , \50539 , \50540 , \50541 , \50542 , \50543 , \50544 , \50545 , \50546 ,
         \50547 , \50548 , \50549 , \50550 , \50551 , \50552 , \50553 , \50554 , \50555 , \50556 ,
         \50557 , \50558 , \50559 , \50560 , \50561 , \50562 , \50563 , \50564 , \50565 , \50566 ,
         \50567 , \50568 , \50569 , \50570 , \50571 , \50572 , \50573 , \50574 , \50575 , \50576 ,
         \50577 , \50578 , \50579 , \50580 , \50581 , \50582 , \50583 , \50584 , \50585 , \50586 ,
         \50587 , \50588 , \50589 , \50590 , \50591 , \50592 , \50593 , \50594 , \50595 , \50596 ,
         \50597 , \50598 , \50599 , \50600 , \50601 , \50602 , \50603 , \50604 , \50605 , \50606 ,
         \50607 , \50608 , \50609 , \50610 , \50611 , \50612 , \50613 , \50614 , \50615 , \50616 ,
         \50617 , \50618 , \50619 , \50620 , \50621 , \50622 , \50623 , \50624 , \50625 , \50626 ,
         \50627 , \50628 , \50629 , \50630 , \50631 , \50632 , \50633 , \50634 , \50635 , \50636 ,
         \50637 , \50638 , \50639 , \50640 , \50641 , \50642 , \50643 , \50644 , \50645 , \50646 ,
         \50647 , \50648 , \50649 , \50650 , \50651 , \50652 , \50653 , \50654 , \50655 , \50656 ,
         \50657 , \50658 , \50659 , \50660 , \50661 , \50662 , \50663 , \50664 , \50665 , \50666 ,
         \50667 , \50668 , \50669 , \50670 , \50671 , \50672 , \50673 , \50674 , \50675 , \50676 ,
         \50677 , \50678 , \50679 , \50680 , \50681 , \50682 , \50683 , \50684 , \50685 , \50686 ,
         \50687 , \50688 , \50689 , \50690 , \50691 , \50692 , \50693 , \50694 , \50695 , \50696 ,
         \50697 , \50698 , \50699 , \50700 , \50701 , \50702 , \50703 , \50704 , \50705 , \50706 ,
         \50707 , \50708 , \50709 , \50710 , \50711 , \50712 , \50713 , \50714 , \50715 , \50716 ,
         \50717 , \50718 , \50719 , \50720 , \50721 , \50722 , \50723 , \50724 , \50725 , \50726 ,
         \50727 , \50728 , \50729 , \50730 , \50731 , \50732 , \50733 , \50734 , \50735 , \50736 ,
         \50737 , \50738 , \50739 , \50740 , \50741 , \50742 , \50743 , \50744 , \50745 , \50746 ,
         \50747 , \50748 , \50749 , \50750 , \50751 , \50752 , \50753 , \50754 , \50755 , \50756 ,
         \50757 , \50758 , \50759 , \50760 , \50761 , \50762 , \50763 , \50764 , \50765 , \50766 ,
         \50767 , \50768 , \50769 , \50770 , \50771 , \50772 , \50773 , \50774 , \50775 , \50776 ,
         \50777 , \50778 , \50779 , \50780 , \50781 , \50782 , \50783 , \50784 , \50785 , \50786 ,
         \50787 , \50788 , \50789 , \50790 , \50791 , \50792 , \50793 , \50794 , \50795 , \50796 ,
         \50797 , \50798 , \50799 , \50800 , \50801 , \50802 , \50803 , \50804 , \50805 , \50806 ,
         \50807 , \50808 , \50809 , \50810 , \50811 , \50812 , \50813 , \50814 , \50815 , \50816 ,
         \50817 , \50818 , \50819 , \50820 , \50821 , \50822 , \50823 , \50824 , \50825 , \50826 ,
         \50827 , \50828 , \50829 , \50830 , \50831 , \50832 , \50833 , \50834 , \50835 , \50836 ,
         \50837 , \50838 , \50839 , \50840 , \50841 , \50842 , \50843 , \50844 , \50845 , \50846 ,
         \50847 , \50848 , \50849 , \50850 , \50851 , \50852 , \50853 , \50854 , \50855 , \50856 ,
         \50857 , \50858 , \50859 , \50860 , \50861 , \50862 , \50863 , \50864 , \50865 , \50866 ,
         \50867 , \50868 , \50869 , \50870 , \50871 , \50872 , \50873 , \50874 , \50875 , \50876 ,
         \50877 , \50878 , \50879 , \50880 , \50881 , \50882 , \50883 , \50884 , \50885 , \50886 ,
         \50887 , \50888 , \50889 , \50890 , \50891 , \50892 , \50893 , \50894 , \50895 , \50896 ,
         \50897 , \50898 , \50899 , \50900 , \50901 , \50902 , \50903 , \50904 , \50905 , \50906 ,
         \50907 , \50908 , \50909 , \50910 , \50911 , \50912 , \50913 , \50914 , \50915 , \50916 ,
         \50917 , \50918 , \50919 , \50920 , \50921 , \50922 , \50923 , \50924 , \50925 , \50926 ,
         \50927 , \50928 , \50929 , \50930 , \50931 , \50932 , \50933 , \50934 , \50935 , \50936 ,
         \50937 , \50938 , \50939 , \50940 , \50941 , \50942 , \50943 , \50944 , \50945 , \50946 ,
         \50947 , \50948 , \50949 , \50950 , \50951 , \50952 , \50953 , \50954 , \50955 , \50956 ,
         \50957 , \50958 , \50959 , \50960 , \50961 , \50962 , \50963 , \50964 , \50965 , \50966 ,
         \50967 , \50968 , \50969 , \50970 , \50971 , \50972 , \50973 , \50974 , \50975 , \50976 ,
         \50977 , \50978 , \50979 , \50980 , \50981 , \50982 , \50983 , \50984 , \50985 , \50986 ,
         \50987 , \50988 , \50989 , \50990 , \50991 , \50992 , \50993 , \50994 , \50995 , \50996 ,
         \50997 , \50998 , \50999 , \51000 , \51001 , \51002 , \51003 , \51004 , \51005 , \51006 ,
         \51007 , \51008 , \51009 , \51010 , \51011 , \51012 , \51013 , \51014 , \51015 , \51016 ,
         \51017 , \51018 , \51019 , \51020 , \51021 , \51022 , \51023 , \51024 , \51025 , \51026 ,
         \51027 , \51028 , \51029 , \51030 , \51031 , \51032 , \51033 , \51034 , \51035 , \51036 ,
         \51037 , \51038 , \51039 , \51040 , \51041 , \51042 , \51043 , \51044 , \51045 , \51046 ,
         \51047 , \51048 , \51049 , \51050 , \51051 , \51052 , \51053 , \51054 , \51055 , \51056 ,
         \51057 , \51058 , \51059 , \51060 , \51061 , \51062 , \51063 , \51064 , \51065 , \51066 ,
         \51067 , \51068 , \51069 , \51070 , \51071 , \51072 , \51073 , \51074 , \51075 , \51076 ,
         \51077 , \51078 , \51079 , \51080 , \51081 , \51082 , \51083 , \51084 , \51085 , \51086 ,
         \51087 , \51088 , \51089 , \51090 , \51091 , \51092 , \51093 , \51094 , \51095 , \51096 ,
         \51097 , \51098 , \51099 , \51100 , \51101 , \51102 , \51103 , \51104 , \51105 , \51106 ,
         \51107 , \51108 , \51109 , \51110 , \51111 , \51112 , \51113 , \51114 , \51115 , \51116 ,
         \51117 , \51118 , \51119 , \51120 , \51121 , \51122 , \51123 , \51124 , \51125 , \51126 ,
         \51127 , \51128 , \51129 , \51130 , \51131 , \51132 , \51133 , \51134 , \51135 , \51136 ,
         \51137 , \51138 , \51139 , \51140 , \51141 , \51142 , \51143 , \51144 , \51145 , \51146 ,
         \51147 , \51148 , \51149 , \51150 , \51151 , \51152 , \51153 , \51154 , \51155 , \51156 ,
         \51157 , \51158 , \51159 , \51160 , \51161 , \51162 , \51163 , \51164 , \51165 , \51166 ,
         \51167 , \51168 , \51169 , \51170 , \51171 , \51172 , \51173 , \51174 , \51175 , \51176 ,
         \51177 , \51178 , \51179 , \51180 , \51181 , \51182 , \51183 , \51184 , \51185 , \51186 ,
         \51187 , \51188 , \51189 , \51190 , \51191 , \51192 , \51193 , \51194 , \51195 , \51196 ,
         \51197 , \51198 , \51199 , \51200 , \51201 , \51202 , \51203 , \51204 , \51205 , \51206 ,
         \51207 , \51208 , \51209 , \51210 , \51211 , \51212 , \51213 , \51214 , \51215 , \51216 ,
         \51217 , \51218 , \51219 , \51220 , \51221 , \51222 , \51223 , \51224 , \51225 , \51226 ,
         \51227 , \51228 , \51229 , \51230 , \51231 , \51232 , \51233 , \51234 , \51235 , \51236 ,
         \51237 , \51238 , \51239 , \51240 , \51241 , \51242 , \51243 , \51244 , \51245 , \51246 ,
         \51247 , \51248 , \51249 , \51250 , \51251 , \51252 , \51253 , \51254 , \51255 , \51256 ,
         \51257 , \51258 , \51259 , \51260 , \51261 , \51262 , \51263 , \51264 , \51265 , \51266 ,
         \51267 , \51268 , \51269 , \51270 , \51271 , \51272 , \51273 , \51274 , \51275 , \51276 ,
         \51277 , \51278 , \51279 , \51280 , \51281 , \51282 , \51283 , \51284 , \51285 , \51286 ,
         \51287 , \51288 , \51289 , \51290 , \51291 , \51292 , \51293 , \51294 , \51295 , \51296 ,
         \51297 , \51298 , \51299 , \51300 , \51301 , \51302 , \51303 , \51304 , \51305 , \51306 ,
         \51307 , \51308 , \51309 , \51310 , \51311 , \51312 , \51313 , \51314 , \51315 , \51316 ,
         \51317 , \51318 , \51319 , \51320 , \51321 , \51322 , \51323 , \51324 , \51325 , \51326 ,
         \51327 , \51328 , \51329 , \51330 , \51331 , \51332 , \51333 , \51334 , \51335 , \51336 ,
         \51337 , \51338 , \51339 , \51340 , \51341 , \51342 , \51343 , \51344 , \51345 , \51346 ,
         \51347 , \51348 , \51349 , \51350 , \51351 , \51352 , \51353 , \51354 , \51355 , \51356 ,
         \51357 , \51358 , \51359 , \51360 , \51361 , \51362 , \51363 , \51364 , \51365 , \51366 ,
         \51367 , \51368 , \51369 , \51370 , \51371 , \51372 , \51373 , \51374 , \51375 , \51376 ,
         \51377 , \51378 , \51379 , \51380 , \51381 , \51382 , \51383 , \51384 , \51385 , \51386 ,
         \51387 , \51388 , \51389 , \51390 , \51391 , \51392 , \51393 , \51394 , \51395 , \51396 ,
         \51397 , \51398 , \51399 , \51400 , \51401 , \51402 , \51403 , \51404 , \51405 , \51406 ,
         \51407 , \51408 , \51409 , \51410 , \51411 , \51412 , \51413 , \51414 , \51415 , \51416 ,
         \51417 , \51418 , \51419 , \51420 , \51421 , \51422 , \51423 , \51424 , \51425 , \51426 ,
         \51427 , \51428 , \51429 , \51430 , \51431 , \51432 , \51433 , \51434 , \51435 , \51436 ,
         \51437 , \51438 , \51439 , \51440 , \51441 , \51442 , \51443 , \51444 , \51445 , \51446 ,
         \51447 , \51448 , \51449 , \51450 , \51451 , \51452 , \51453 , \51454 , \51455 , \51456 ,
         \51457 , \51458 , \51459 , \51460 , \51461 , \51462 , \51463 , \51464 , \51465 , \51466 ,
         \51467 , \51468 , \51469 , \51470 , \51471 , \51472 , \51473 , \51474 , \51475 , \51476 ,
         \51477 , \51478 , \51479 , \51480 , \51481 , \51482 , \51483 , \51484 , \51485 , \51486 ,
         \51487 , \51488 , \51489 , \51490 , \51491 , \51492 , \51493 , \51494 , \51495 , \51496 ,
         \51497 , \51498 , \51499 , \51500 , \51501 , \51502 , \51503 , \51504 , \51505 , \51506 ,
         \51507 , \51508 , \51509 , \51510 , \51511 , \51512 , \51513 , \51514 , \51515 , \51516 ,
         \51517 , \51518 , \51519 , \51520 , \51521 , \51522 , \51523 , \51524 , \51525 , \51526 ,
         \51527 , \51528 , \51529 , \51530 , \51531 , \51532 , \51533 , \51534 , \51535 , \51536 ,
         \51537 , \51538 , \51539 , \51540 , \51541 , \51542 , \51543 , \51544 , \51545 , \51546 ,
         \51547 , \51548 , \51549 , \51550 , \51551 , \51552 , \51553 , \51554 , \51555 , \51556 ,
         \51557 , \51558 , \51559 , \51560 , \51561 , \51562 , \51563 , \51564 , \51565 , \51566 ,
         \51567 , \51568 , \51569 , \51570 , \51571 , \51572 , \51573 , \51574 , \51575 , \51576 ,
         \51577 , \51578 , \51579 , \51580 , \51581 , \51582 , \51583 , \51584 , \51585 , \51586 ,
         \51587 , \51588 , \51589 , \51590 , \51591 , \51592 , \51593 , \51594 , \51595 , \51596 ,
         \51597 , \51598 , \51599 , \51600 , \51601 , \51602 , \51603 , \51604 , \51605 , \51606 ,
         \51607 , \51608 , \51609 , \51610 , \51611 , \51612 , \51613 , \51614 , \51615 , \51616 ,
         \51617 , \51618 , \51619 , \51620 , \51621 , \51622 , \51623 , \51624 , \51625 , \51626 ,
         \51627 , \51628 , \51629 , \51630 , \51631 , \51632 , \51633 , \51634 , \51635 , \51636 ,
         \51637 , \51638 , \51639 , \51640 , \51641 , \51642 , \51643 , \51644 , \51645 , \51646 ,
         \51647 , \51648 , \51649 , \51650 , \51651 , \51652 , \51653 , \51654 , \51655 , \51656 ,
         \51657 , \51658 , \51659 , \51660 , \51661 , \51662 , \51663 , \51664 , \51665 , \51666 ,
         \51667 , \51668 , \51669 , \51670 , \51671 , \51672 , \51673 , \51674 , \51675 , \51676 ,
         \51677 , \51678 , \51679 , \51680 , \51681 , \51682 , \51683 , \51684 , \51685 , \51686 ,
         \51687 , \51688 , \51689 , \51690 , \51691 , \51692 , \51693 , \51694 , \51695 , \51696 ,
         \51697 , \51698 , \51699 , \51700 , \51701 , \51702 , \51703 , \51704 , \51705 , \51706 ,
         \51707 , \51708 , \51709 , \51710 , \51711 , \51712 , \51713 , \51714 , \51715 , \51716 ,
         \51717 , \51718 , \51719 , \51720 , \51721 , \51722 , \51723 , \51724 , \51725 , \51726 ,
         \51727 , \51728 , \51729 , \51730 , \51731 , \51732 , \51733 , \51734 , \51735 , \51736 ,
         \51737 , \51738 , \51739 , \51740 , \51741 , \51742 , \51743 , \51744 , \51745 , \51746 ,
         \51747 , \51748 , \51749 , \51750 , \51751 , \51752 , \51753 , \51754 , \51755 , \51756 ,
         \51757 , \51758 , \51759 , \51760 , \51761 , \51762 , \51763 , \51764 , \51765 , \51766 ,
         \51767 , \51768 , \51769 , \51770 , \51771 , \51772 , \51773 , \51774 , \51775 , \51776 ,
         \51777 , \51778 , \51779 , \51780 , \51781 , \51782 , \51783 , \51784 , \51785 , \51786 ,
         \51787 , \51788 , \51789 , \51790 , \51791 , \51792 , \51793 , \51794 , \51795 , \51796 ,
         \51797 , \51798 , \51799 , \51800 , \51801 , \51802 , \51803 , \51804 , \51805 , \51806 ,
         \51807 , \51808 , \51809 , \51810 , \51811 , \51812 , \51813 , \51814 , \51815 , \51816 ,
         \51817 , \51818 , \51819 , \51820 , \51821 , \51822 , \51823 , \51824 , \51825 , \51826 ,
         \51827 , \51828 , \51829 , \51830 , \51831 , \51832 , \51833 , \51834 , \51835 , \51836 ,
         \51837 , \51838 , \51839 , \51840 , \51841 , \51842 , \51843 , \51844 , \51845 , \51846 ,
         \51847 , \51848 , \51849 , \51850 , \51851 , \51852 , \51853 , \51854 , \51855 , \51856 ,
         \51857 , \51858 , \51859 , \51860 , \51861 , \51862 , \51863 , \51864 , \51865 , \51866 ,
         \51867 , \51868 , \51869 , \51870 , \51871 , \51872 , \51873 , \51874 , \51875 , \51876 ,
         \51877 , \51878 , \51879 , \51880 , \51881 , \51882 , \51883 , \51884 , \51885 , \51886 ,
         \51887 , \51888 , \51889 , \51890 , \51891 , \51892 , \51893 , \51894 , \51895 , \51896 ,
         \51897 , \51898 , \51899 , \51900 , \51901 , \51902 , \51903 , \51904 , \51905 , \51906 ,
         \51907 , \51908 , \51909 , \51910 , \51911 , \51912 , \51913 , \51914 , \51915 , \51916 ,
         \51917 , \51918 , \51919 , \51920 , \51921 , \51922 , \51923 , \51924 , \51925 , \51926 ,
         \51927 , \51928 , \51929 , \51930 , \51931 , \51932 , \51933 , \51934 , \51935 , \51936 ,
         \51937 , \51938 , \51939 , \51940 , \51941 , \51942 , \51943 , \51944 , \51945 , \51946 ,
         \51947 , \51948 , \51949 , \51950 , \51951 , \51952 , \51953 , \51954 , \51955 , \51956 ,
         \51957 , \51958 , \51959 , \51960 , \51961 , \51962 , \51963 , \51964 , \51965 , \51966 ,
         \51967 , \51968 , \51969 , \51970 , \51971 , \51972 , \51973 , \51974 , \51975 , \51976 ,
         \51977 , \51978 , \51979 , \51980 , \51981 , \51982 , \51983 , \51984 , \51985 , \51986 ,
         \51987 , \51988 , \51989 , \51990 , \51991 , \51992 , \51993 , \51994 , \51995 , \51996 ,
         \51997 , \51998 , \51999 , \52000 , \52001 , \52002 , \52003 , \52004 , \52005 , \52006 ,
         \52007 , \52008 , \52009 , \52010 , \52011 , \52012 , \52013 , \52014 , \52015 , \52016 ,
         \52017 , \52018 , \52019 , \52020 , \52021 , \52022 , \52023 , \52024 , \52025 , \52026 ,
         \52027 , \52028 , \52029 , \52030 , \52031 , \52032 , \52033 , \52034 , \52035 , \52036 ,
         \52037 , \52038 , \52039 , \52040 , \52041 , \52042 , \52043 , \52044 , \52045 , \52046 ,
         \52047 , \52048 , \52049 , \52050 , \52051 , \52052 , \52053 , \52054 , \52055 , \52056 ,
         \52057 , \52058 , \52059 , \52060 , \52061 , \52062 , \52063 , \52064 , \52065 , \52066 ,
         \52067 , \52068 , \52069 , \52070 , \52071 , \52072 , \52073 , \52074 , \52075 , \52076 ,
         \52077 , \52078 , \52079 , \52080 , \52081 , \52082 , \52083 , \52084 , \52085 , \52086 ,
         \52087 , \52088 , \52089 , \52090 , \52091 , \52092 , \52093 , \52094 , \52095 , \52096 ,
         \52097 , \52098 , \52099 , \52100 , \52101 , \52102 , \52103 , \52104 , \52105 , \52106 ,
         \52107 , \52108 , \52109 , \52110 , \52111 , \52112 , \52113 , \52114 , \52115 , \52116 ,
         \52117 , \52118 , \52119 , \52120 , \52121 , \52122 , \52123 , \52124 , \52125 , \52126 ,
         \52127 , \52128 , \52129 , \52130 , \52131 , \52132 , \52133 , \52134 , \52135 , \52136 ,
         \52137 , \52138 , \52139 , \52140 , \52141 , \52142 , \52143 , \52144 , \52145 , \52146 ,
         \52147 , \52148 , \52149 , \52150 , \52151 , \52152 , \52153 , \52154 , \52155 , \52156 ,
         \52157 , \52158 , \52159 , \52160 , \52161 , \52162 , \52163 , \52164 , \52165 , \52166 ,
         \52167 , \52168 , \52169 , \52170 , \52171 , \52172 , \52173 , \52174 , \52175 , \52176 ,
         \52177 , \52178 , \52179 , \52180 , \52181 , \52182 , \52183 , \52184 , \52185 , \52186 ,
         \52187 , \52188 , \52189 , \52190 , \52191 , \52192 , \52193 , \52194 , \52195 , \52196 ,
         \52197 , \52198 , \52199 , \52200 , \52201 , \52202 , \52203 , \52204 , \52205 , \52206 ,
         \52207 , \52208 , \52209 , \52210 , \52211 , \52212 , \52213 , \52214 , \52215 , \52216 ,
         \52217 , \52218 , \52219 , \52220 , \52221 , \52222 , \52223 , \52224 , \52225 , \52226 ,
         \52227 , \52228 , \52229 , \52230 , \52231 , \52232 , \52233 , \52234 , \52235 , \52236 ,
         \52237 , \52238 , \52239 , \52240 , \52241 , \52242 , \52243 , \52244 , \52245 , \52246 ,
         \52247 , \52248 , \52249 , \52250 , \52251 , \52252 , \52253 , \52254 , \52255 , \52256 ,
         \52257 , \52258 , \52259 , \52260 , \52261 , \52262 , \52263 , \52264 , \52265 , \52266 ,
         \52267 , \52268 , \52269 , \52270 , \52271 , \52272 , \52273 , \52274 , \52275 , \52276 ,
         \52277 , \52278 , \52279 , \52280 , \52281 , \52282 , \52283 , \52284 , \52285 , \52286 ,
         \52287 , \52288 , \52289 , \52290 , \52291 , \52292 , \52293 , \52294 , \52295 , \52296 ,
         \52297 , \52298 , \52299 , \52300 , \52301 , \52302 , \52303 , \52304 , \52305 , \52306 ,
         \52307 , \52308 , \52309 , \52310 , \52311 , \52312 , \52313 , \52314 , \52315 , \52316 ,
         \52317 , \52318 , \52319 , \52320 , \52321 , \52322 , \52323 , \52324 , \52325 , \52326 ,
         \52327 , \52328 , \52329 , \52330 , \52331 , \52332 , \52333 , \52334 , \52335 , \52336 ,
         \52337 , \52338 , \52339 , \52340 , \52341 , \52342 , \52343 , \52344 , \52345 , \52346 ,
         \52347 , \52348 , \52349 , \52350 , \52351 , \52352 , \52353 , \52354 , \52355 , \52356 ,
         \52357 , \52358 , \52359 , \52360 , \52361 , \52362 , \52363 , \52364 , \52365 , \52366 ,
         \52367 , \52368 , \52369 , \52370 , \52371 , \52372 , \52373 , \52374 , \52375 , \52376 ,
         \52377 , \52378 , \52379 , \52380 , \52381 , \52382 , \52383 , \52384 , \52385 , \52386 ,
         \52387 , \52388 , \52389 , \52390 , \52391 , \52392 , \52393 , \52394 , \52395 , \52396 ,
         \52397 , \52398 , \52399 , \52400 , \52401 , \52402 , \52403 , \52404 , \52405 , \52406 ,
         \52407 , \52408 , \52409 , \52410 , \52411 , \52412 , \52413 , \52414 , \52415 , \52416 ,
         \52417 , \52418 , \52419 , \52420 , \52421 , \52422 , \52423 , \52424 , \52425 , \52426 ,
         \52427 , \52428 , \52429 , \52430 , \52431 , \52432 , \52433 , \52434 , \52435 , \52436 ,
         \52437 , \52438 , \52439 , \52440 , \52441 , \52442 , \52443 , \52444 , \52445 , \52446 ,
         \52447 , \52448 , \52449 , \52450 , \52451 , \52452 , \52453 , \52454 , \52455 , \52456 ,
         \52457 , \52458 , \52459 , \52460 , \52461 , \52462 , \52463 , \52464 , \52465 , \52466 ,
         \52467 , \52468 , \52469 , \52470 , \52471 , \52472 , \52473 , \52474 , \52475 , \52476 ,
         \52477 , \52478 , \52479 , \52480 , \52481 , \52482 , \52483 , \52484 , \52485 , \52486 ,
         \52487 , \52488 , \52489 , \52490 , \52491 , \52492 , \52493 , \52494 , \52495 , \52496 ,
         \52497 , \52498 , \52499 , \52500 , \52501 , \52502 , \52503 , \52504 , \52505 , \52506 ,
         \52507 , \52508 , \52509 , \52510 , \52511 , \52512 , \52513 , \52514 , \52515 , \52516 ,
         \52517 , \52518 , \52519 , \52520 , \52521 , \52522 , \52523 , \52524 , \52525 , \52526 ,
         \52527 , \52528 , \52529 , \52530 , \52531 , \52532 , \52533 , \52534 , \52535 , \52536 ,
         \52537 , \52538 , \52539 , \52540 , \52541 , \52542 , \52543 , \52544 , \52545 , \52546 ,
         \52547 , \52548 , \52549 , \52550 , \52551 , \52552 , \52553 , \52554 , \52555 , \52556 ,
         \52557 , \52558 , \52559 , \52560 , \52561 , \52562 , \52563 , \52564 , \52565 , \52566 ,
         \52567 , \52568 , \52569 , \52570 , \52571 , \52572 , \52573 , \52574 , \52575 , \52576 ,
         \52577 , \52578 , \52579 , \52580 , \52581 , \52582 , \52583 , \52584 , \52585 , \52586 ,
         \52587 , \52588 , \52589 , \52590 , \52591 , \52592 , \52593 , \52594 , \52595 , \52596 ,
         \52597 , \52598 , \52599 , \52600 , \52601 , \52602 , \52603 , \52604 , \52605 , \52606 ,
         \52607 , \52608 , \52609 , \52610 , \52611 , \52612 , \52613 , \52614 , \52615 , \52616 ,
         \52617 , \52618 , \52619 , \52620 , \52621 , \52622 , \52623 , \52624 , \52625 , \52626 ,
         \52627 , \52628 , \52629 , \52630 , \52631 , \52632 , \52633 , \52634 , \52635 , \52636 ,
         \52637 , \52638 , \52639 , \52640 , \52641 , \52642 , \52643 , \52644 , \52645 , \52646 ,
         \52647 , \52648 , \52649 , \52650 , \52651 , \52652 , \52653 , \52654 , \52655 , \52656 ,
         \52657 , \52658 , \52659 , \52660 , \52661 , \52662 , \52663 , \52664 , \52665 , \52666 ,
         \52667 , \52668 , \52669 , \52670 , \52671 , \52672 , \52673 , \52674 , \52675 , \52676 ,
         \52677 , \52678 , \52679 , \52680 , \52681 , \52682 , \52683 , \52684 , \52685 , \52686 ,
         \52687 , \52688 , \52689 , \52690 , \52691 , \52692 , \52693 , \52694 , \52695 , \52696 ,
         \52697 , \52698 , \52699 , \52700 , \52701 , \52702 , \52703 , \52704 , \52705 , \52706 ,
         \52707 , \52708 , \52709 , \52710 , \52711 , \52712 , \52713 , \52714 , \52715 , \52716 ,
         \52717 , \52718 , \52719 , \52720 , \52721 , \52722 , \52723 , \52724 , \52725 , \52726 ,
         \52727 , \52728 , \52729 , \52730 , \52731 , \52732 , \52733 , \52734 , \52735 , \52736 ,
         \52737 , \52738 , \52739 , \52740 , \52741 , \52742 , \52743 , \52744 , \52745 , \52746 ,
         \52747 , \52748 , \52749 , \52750 , \52751 , \52752 , \52753 , \52754 , \52755 , \52756 ,
         \52757 , \52758 , \52759 , \52760 , \52761 , \52762 , \52763 , \52764 , \52765 , \52766 ,
         \52767 , \52768 , \52769 , \52770 , \52771 , \52772 , \52773 , \52774 , \52775 , \52776 ,
         \52777 , \52778 , \52779 , \52780 , \52781 , \52782 , \52783 , \52784 , \52785 , \52786 ,
         \52787 , \52788 , \52789 , \52790 , \52791 , \52792 , \52793 , \52794 , \52795 , \52796 ,
         \52797 , \52798 , \52799 , \52800 , \52801 , \52802 , \52803 , \52804 , \52805 , \52806 ,
         \52807 , \52808 , \52809 , \52810 , \52811 , \52812 , \52813 , \52814 , \52815 , \52816 ,
         \52817 , \52818 , \52819 , \52820 , \52821 , \52822 , \52823 , \52824 , \52825 , \52826 ,
         \52827 , \52828 , \52829 , \52830 , \52831 , \52832 , \52833 , \52834 , \52835 , \52836 ,
         \52837 , \52838 , \52839 , \52840 , \52841 , \52842 , \52843 , \52844 , \52845 , \52846 ,
         \52847 , \52848 , \52849 , \52850 , \52851 , \52852 , \52853 , \52854 , \52855 , \52856 ,
         \52857 , \52858 , \52859 , \52860 , \52861 , \52862 , \52863 , \52864 , \52865 , \52866 ,
         \52867 , \52868 , \52869 , \52870 , \52871 , \52872 , \52873 , \52874 , \52875 , \52876 ,
         \52877 , \52878 , \52879 , \52880 , \52881 , \52882 , \52883 , \52884 , \52885 , \52886 ,
         \52887 , \52888 , \52889 , \52890 , \52891 , \52892 , \52893 , \52894 , \52895 , \52896 ,
         \52897 , \52898 , \52899 , \52900 , \52901 , \52902 , \52903 , \52904 , \52905 , \52906 ,
         \52907 , \52908 , \52909 , \52910 , \52911 , \52912 , \52913 , \52914 , \52915 , \52916 ,
         \52917 , \52918 , \52919 , \52920 , \52921 , \52922 , \52923 , \52924 , \52925 , \52926 ,
         \52927 , \52928 , \52929 , \52930 , \52931 , \52932 , \52933 , \52934 , \52935 , \52936 ,
         \52937 , \52938 , \52939 , \52940 , \52941 , \52942 , \52943 , \52944 , \52945 , \52946 ,
         \52947 , \52948 , \52949 , \52950 , \52951 , \52952 , \52953 , \52954 , \52955 , \52956 ,
         \52957 , \52958 , \52959 , \52960 , \52961 , \52962 , \52963 , \52964 , \52965 , \52966 ,
         \52967 , \52968 , \52969 , \52970 , \52971 , \52972 , \52973 , \52974 , \52975 , \52976 ,
         \52977 , \52978 , \52979 , \52980 , \52981 , \52982 , \52983 , \52984 , \52985 , \52986 ,
         \52987 , \52988 , \52989 , \52990 , \52991 , \52992 , \52993 , \52994 , \52995 , \52996 ,
         \52997 , \52998 , \52999 , \53000 , \53001 , \53002 , \53003 , \53004 , \53005 , \53006 ,
         \53007 , \53008 , \53009 , \53010 , \53011 , \53012 , \53013 , \53014 , \53015 , \53016 ,
         \53017 , \53018 , \53019 , \53020 , \53021 , \53022 , \53023 , \53024 , \53025 , \53026 ,
         \53027 , \53028 , \53029 , \53030 , \53031 , \53032 , \53033 , \53034 , \53035 , \53036 ,
         \53037 , \53038 , \53039 , \53040 , \53041 , \53042 , \53043 , \53044 , \53045 , \53046 ,
         \53047 , \53048 , \53049 , \53050 , \53051 , \53052 , \53053 , \53054 , \53055 , \53056 ,
         \53057 , \53058 , \53059 , \53060 , \53061 , \53062 , \53063 , \53064 , \53065 , \53066 ,
         \53067 , \53068 , \53069 , \53070 , \53071 , \53072 , \53073 , \53074 , \53075 , \53076 ,
         \53077 , \53078 , \53079 , \53080 , \53081 , \53082 , \53083 , \53084 , \53085 , \53086 ,
         \53087 , \53088 , \53089 , \53090 , \53091 , \53092 , \53093 , \53094 , \53095 , \53096 ,
         \53097 , \53098 , \53099 , \53100 , \53101 , \53102 , \53103 , \53104 , \53105 , \53106 ,
         \53107 , \53108 , \53109 , \53110 , \53111 , \53112 , \53113 , \53114 , \53115 , \53116 ,
         \53117 , \53118 , \53119 , \53120 , \53121 , \53122 , \53123 , \53124 , \53125 , \53126 ,
         \53127 , \53128 , \53129 , \53130 , \53131 , \53132 , \53133 , \53134 , \53135 , \53136 ,
         \53137 , \53138 , \53139 , \53140 , \53141 , \53142 , \53143 , \53144 , \53145 , \53146 ,
         \53147 , \53148 , \53149 , \53150 , \53151 , \53152 , \53153 , \53154 , \53155 , \53156 ,
         \53157 , \53158 , \53159 , \53160 , \53161 , \53162 , \53163 , \53164 , \53165 , \53166 ,
         \53167 , \53168 , \53169 , \53170 , \53171 , \53172 , \53173 , \53174 , \53175 , \53176 ,
         \53177 , \53178 , \53179 , \53180 , \53181 , \53182 , \53183 , \53184 , \53185 , \53186 ,
         \53187 , \53188 , \53189 , \53190 , \53191 , \53192 , \53193 , \53194 , \53195 , \53196 ,
         \53197 , \53198 , \53199 , \53200 , \53201 , \53202 , \53203 , \53204 , \53205 , \53206 ,
         \53207 , \53208 , \53209 , \53210 , \53211 , \53212 , \53213 , \53214 , \53215 , \53216 ,
         \53217 , \53218 , \53219 , \53220 , \53221 , \53222 , \53223 , \53224 , \53225 , \53226 ,
         \53227 , \53228 , \53229 , \53230 , \53231 , \53232 , \53233 , \53234 , \53235 , \53236 ,
         \53237 , \53238 , \53239 , \53240 , \53241 , \53242 , \53243 , \53244 , \53245 , \53246 ,
         \53247 , \53248 , \53249 , \53250 , \53251 , \53252 , \53253 , \53254 , \53255 , \53256 ,
         \53257 , \53258 , \53259 , \53260 , \53261 , \53262 , \53263 , \53264 , \53265 , \53266 ,
         \53267 , \53268 , \53269 , \53270 , \53271 , \53272 , \53273 , \53274 , \53275 , \53276 ,
         \53277 , \53278 , \53279 , \53280 , \53281 , \53282 , \53283 , \53284 , \53285 , \53286 ,
         \53287 , \53288 , \53289 , \53290 , \53291 , \53292 , \53293 , \53294 , \53295 , \53296 ,
         \53297 , \53298 , \53299 , \53300 , \53301 , \53302 , \53303 , \53304 , \53305 , \53306 ,
         \53307 , \53308 , \53309 , \53310 , \53311 , \53312 , \53313 , \53314 , \53315 , \53316 ,
         \53317 , \53318 , \53319 , \53320 , \53321 , \53322 , \53323 , \53324 , \53325 , \53326 ,
         \53327 , \53328 , \53329 , \53330 , \53331 , \53332 , \53333 , \53334 , \53335 , \53336 ,
         \53337 , \53338 , \53339 , \53340 , \53341 , \53342 , \53343 , \53344 , \53345 , \53346 ,
         \53347 , \53348 , \53349 , \53350 , \53351 , \53352 , \53353 , \53354 , \53355 , \53356 ,
         \53357 , \53358 , \53359 , \53360 , \53361 , \53362 , \53363 , \53364 , \53365 , \53366 ,
         \53367 , \53368 , \53369 , \53370 , \53371 , \53372 , \53373 , \53374 , \53375 , \53376 ,
         \53377 , \53378 , \53379 , \53380 , \53381 , \53382 , \53383 , \53384 , \53385 , \53386 ,
         \53387 , \53388 , \53389 , \53390 , \53391 , \53392 , \53393 , \53394 , \53395 , \53396 ,
         \53397 , \53398 , \53399 , \53400 , \53401 , \53402 , \53403 , \53404 , \53405 , \53406 ,
         \53407 , \53408 , \53409 , \53410 , \53411 , \53412 , \53413 , \53414 , \53415 , \53416 ,
         \53417 , \53418 , \53419 , \53420 , \53421 , \53422 , \53423 , \53424 , \53425 , \53426 ,
         \53427 , \53428 , \53429 , \53430 , \53431 , \53432 , \53433 , \53434 , \53435 , \53436 ,
         \53437 , \53438 , \53439 , \53440 , \53441 , \53442 , \53443 , \53444 , \53445 , \53446 ,
         \53447 , \53448 , \53449 , \53450 , \53451 , \53452 , \53453 , \53454 , \53455 , \53456 ,
         \53457 , \53458 , \53459 , \53460 , \53461 , \53462 , \53463 , \53464 , \53465 , \53466 ,
         \53467 , \53468 , \53469 , \53470 , \53471 , \53472 , \53473 , \53474 , \53475 , \53476 ,
         \53477 , \53478 , \53479 , \53480 , \53481 , \53482 , \53483 , \53484 , \53485 , \53486 ,
         \53487 , \53488 , \53489 , \53490 , \53491 , \53492 , \53493 , \53494 , \53495 , \53496 ,
         \53497 , \53498 , \53499 , \53500 , \53501 , \53502 , \53503 , \53504 , \53505 , \53506 ,
         \53507 , \53508 , \53509 , \53510 , \53511 , \53512 , \53513 , \53514 , \53515 , \53516 ,
         \53517 , \53518 , \53519 , \53520 , \53521 , \53522 , \53523 , \53524 , \53525 , \53526 ,
         \53527 , \53528 , \53529 , \53530 , \53531 , \53532 , \53533 , \53534 , \53535 , \53536 ,
         \53537 , \53538 , \53539 , \53540 , \53541 , \53542 , \53543 , \53544 , \53545 , \53546 ,
         \53547 , \53548 , \53549 , \53550 , \53551 , \53552 , \53553 , \53554 , \53555 , \53556 ,
         \53557 , \53558 , \53559 , \53560 , \53561 , \53562 , \53563 , \53564 , \53565 , \53566 ,
         \53567 , \53568 , \53569 , \53570 , \53571 , \53572 , \53573 , \53574 , \53575 , \53576 ,
         \53577 , \53578 , \53579 , \53580 , \53581 , \53582 , \53583 , \53584 , \53585 , \53586 ,
         \53587 , \53588 , \53589 , \53590 , \53591 , \53592 , \53593 , \53594 , \53595 , \53596 ,
         \53597 , \53598 , \53599 , \53600 , \53601 , \53602 , \53603 , \53604 , \53605 , \53606 ,
         \53607 , \53608 , \53609 , \53610 , \53611 , \53612 , \53613 , \53614 , \53615 , \53616 ,
         \53617 , \53618 , \53619 , \53620 , \53621 , \53622 , \53623 , \53624 , \53625 , \53626 ,
         \53627 , \53628 , \53629 , \53630 , \53631 , \53632 , \53633 , \53634 , \53635 , \53636 ,
         \53637 , \53638 , \53639 , \53640 , \53641 , \53642 , \53643 , \53644 , \53645 , \53646 ,
         \53647 , \53648 , \53649 , \53650 , \53651 , \53652 , \53653 , \53654 , \53655 , \53656 ,
         \53657 , \53658 , \53659 , \53660 , \53661 , \53662 , \53663 , \53664 , \53665 , \53666 ,
         \53667 , \53668 , \53669 , \53670 , \53671 , \53672 , \53673 , \53674 , \53675 , \53676 ,
         \53677 , \53678 , \53679 , \53680 , \53681 , \53682 , \53683 , \53684 , \53685 , \53686 ,
         \53687 , \53688 , \53689 , \53690 , \53691 , \53692 , \53693 , \53694 , \53695 , \53696 ,
         \53697 , \53698 , \53699 , \53700 , \53701 , \53702 , \53703 , \53704 , \53705 , \53706 ,
         \53707 , \53708 , \53709 , \53710 , \53711 , \53712 , \53713 , \53714 , \53715 , \53716 ,
         \53717 , \53718 , \53719 , \53720 , \53721 , \53722 , \53723 , \53724 , \53725 , \53726 ,
         \53727 , \53728 , \53729 , \53730 , \53731 , \53732 , \53733 , \53734 , \53735 , \53736 ,
         \53737 , \53738 , \53739 , \53740 , \53741 , \53742 , \53743 , \53744 , \53745 , \53746 ,
         \53747 , \53748 , \53749 , \53750 , \53751 , \53752 , \53753 , \53754 , \53755 , \53756 ,
         \53757 , \53758 , \53759 , \53760 , \53761 , \53762 , \53763 , \53764 , \53765 , \53766 ,
         \53767 , \53768 , \53769 , \53770 , \53771 , \53772 , \53773 , \53774 , \53775 , \53776 ,
         \53777 , \53778 , \53779 , \53780 , \53781 , \53782 , \53783 , \53784 , \53785 , \53786 ,
         \53787 , \53788 , \53789 , \53790 , \53791 , \53792 , \53793 , \53794 , \53795 , \53796 ,
         \53797 , \53798 , \53799 , \53800 , \53801 , \53802 , \53803 , \53804 , \53805 , \53806 ,
         \53807 , \53808 , \53809 , \53810 , \53811 , \53812 , \53813 , \53814 , \53815 , \53816 ,
         \53817 , \53818 , \53819 , \53820 , \53821 , \53822 , \53823 , \53824 , \53825 , \53826 ,
         \53827 , \53828 , \53829 , \53830 , \53831 , \53832 , \53833 , \53834 , \53835 , \53836 ,
         \53837 , \53838 , \53839 , \53840 , \53841 , \53842 , \53843 , \53844 , \53845 , \53846 ,
         \53847 , \53848 , \53849 , \53850 , \53851 , \53852 , \53853 , \53854 , \53855 , \53856 ,
         \53857 , \53858 , \53859 , \53860 , \53861 , \53862 , \53863 , \53864 , \53865 , \53866 ,
         \53867 , \53868 , \53869 , \53870 , \53871 , \53872 , \53873 , \53874 , \53875 , \53876 ,
         \53877 , \53878 , \53879 , \53880 , \53881 , \53882 , \53883 , \53884 , \53885 , \53886 ,
         \53887 , \53888 , \53889 , \53890 , \53891 , \53892 , \53893 , \53894 , \53895 , \53896 ,
         \53897 , \53898 , \53899 , \53900 , \53901 , \53902 , \53903 , \53904 , \53905 , \53906 ,
         \53907 , \53908 , \53909 , \53910 , \53911 , \53912 , \53913 , \53914 , \53915 , \53916 ,
         \53917 , \53918 , \53919 , \53920 , \53921 , \53922 , \53923 , \53924 , \53925 , \53926 ,
         \53927 , \53928 , \53929 , \53930 , \53931 , \53932 , \53933 , \53934 , \53935 , \53936 ,
         \53937 , \53938 , \53939 , \53940 , \53941 , \53942 , \53943 , \53944 , \53945 , \53946 ,
         \53947 , \53948 , \53949 , \53950 , \53951 , \53952 , \53953 , \53954 , \53955 , \53956 ,
         \53957 , \53958 , \53959 , \53960 , \53961 , \53962 , \53963 , \53964 , \53965 , \53966 ,
         \53967 , \53968 , \53969 , \53970 , \53971 , \53972 , \53973 , \53974 , \53975 , \53976 ,
         \53977 , \53978 , \53979 , \53980 , \53981 , \53982 , \53983 , \53984 , \53985 , \53986 ,
         \53987 , \53988 , \53989 , \53990 , \53991 , \53992 , \53993 , \53994 , \53995 , \53996 ,
         \53997 , \53998 , \53999 , \54000 , \54001 , \54002 , \54003 , \54004 , \54005 , \54006 ,
         \54007 , \54008 , \54009 , \54010 , \54011 , \54012 , \54013 , \54014 , \54015 , \54016 ,
         \54017 , \54018 , \54019 , \54020 , \54021 , \54022 , \54023 , \54024 , \54025 , \54026 ,
         \54027 , \54028 , \54029 , \54030 , \54031 , \54032 , \54033 , \54034 , \54035 , \54036 ,
         \54037 , \54038 , \54039 , \54040 , \54041 , \54042 , \54043 , \54044 , \54045 , \54046 ,
         \54047 , \54048 , \54049 , \54050 , \54051 , \54052 , \54053 , \54054 , \54055 , \54056 ,
         \54057 , \54058 , \54059 , \54060 , \54061 , \54062 , \54063 , \54064 , \54065 , \54066 ,
         \54067 , \54068 , \54069 , \54070 , \54071 , \54072 , \54073 , \54074 , \54075 , \54076 ,
         \54077 , \54078 , \54079 , \54080 , \54081 , \54082 , \54083 , \54084 , \54085 , \54086 ,
         \54087 , \54088 , \54089 , \54090 , \54091 , \54092 , \54093 , \54094 , \54095 , \54096 ,
         \54097 , \54098 , \54099 , \54100 , \54101 , \54102 , \54103 , \54104 , \54105 , \54106 ,
         \54107 , \54108 , \54109 , \54110 , \54111 , \54112 , \54113 , \54114 , \54115 , \54116 ,
         \54117 , \54118 , \54119 , \54120 , \54121 , \54122 , \54123 , \54124 , \54125 , \54126 ,
         \54127 , \54128 , \54129 , \54130 , \54131 , \54132 , \54133 , \54134 , \54135 , \54136 ,
         \54137 , \54138 , \54139 , \54140 , \54141 , \54142 , \54143 , \54144 , \54145 , \54146 ,
         \54147 , \54148 , \54149 , \54150 , \54151 , \54152 , \54153 , \54154 , \54155 , \54156 ,
         \54157 , \54158 , \54159 , \54160 , \54161 , \54162 , \54163 , \54164 , \54165 , \54166 ,
         \54167 , \54168 , \54169 , \54170 , \54171 , \54172 , \54173 , \54174 , \54175 , \54176 ,
         \54177 , \54178 , \54179 , \54180 , \54181 , \54182 , \54183 , \54184 , \54185 , \54186 ,
         \54187 , \54188 , \54189 , \54190 , \54191 , \54192 , \54193 , \54194 , \54195 , \54196 ,
         \54197 , \54198 , \54199 , \54200 , \54201 , \54202 , \54203 , \54204 , \54205 , \54206 ,
         \54207 , \54208 , \54209 , \54210 , \54211 , \54212 , \54213 , \54214 , \54215 , \54216 ,
         \54217 , \54218 , \54219 , \54220 , \54221 , \54222 , \54223 , \54224 , \54225 , \54226 ,
         \54227 , \54228 , \54229 , \54230 , \54231 , \54232 , \54233 , \54234 , \54235 , \54236 ,
         \54237 , \54238 , \54239 , \54240 , \54241 , \54242 , \54243 , \54244 , \54245 , \54246 ,
         \54247 , \54248 , \54249 , \54250 , \54251 , \54252 , \54253 , \54254 , \54255 , \54256 ,
         \54257 , \54258 , \54259 , \54260 , \54261 , \54262 , \54263 , \54264 , \54265 , \54266 ,
         \54267 , \54268 , \54269 , \54270 , \54271 , \54272 , \54273 , \54274 , \54275 , \54276 ,
         \54277 , \54278 , \54279 , \54280 , \54281 , \54282 , \54283 , \54284 , \54285 , \54286 ,
         \54287 , \54288 , \54289 , \54290 , \54291 , \54292 , \54293 , \54294 , \54295 , \54296 ,
         \54297 , \54298 , \54299 , \54300 , \54301 , \54302 , \54303 , \54304 , \54305 , \54306 ,
         \54307 , \54308 , \54309 , \54310 , \54311 , \54312 , \54313 , \54314 , \54315 , \54316 ,
         \54317 , \54318 , \54319 , \54320 , \54321 , \54322 , \54323 , \54324 , \54325 , \54326 ,
         \54327 , \54328 , \54329 , \54330 , \54331 , \54332 , \54333 , \54334 , \54335 , \54336 ,
         \54337 , \54338 , \54339 , \54340 , \54341 , \54342 , \54343 , \54344 , \54345 , \54346 ,
         \54347 , \54348 , \54349 , \54350 , \54351 , \54352 , \54353 , \54354 , \54355 , \54356 ,
         \54357 , \54358 , \54359 , \54360 , \54361 , \54362 , \54363 , \54364 , \54365 , \54366 ,
         \54367 , \54368 , \54369 , \54370 , \54371 , \54372 , \54373 , \54374 , \54375 , \54376 ,
         \54377 , \54378 , \54379 , \54380 , \54381 , \54382 , \54383 , \54384 , \54385 , \54386 ,
         \54387 , \54388 , \54389 , \54390 , \54391 , \54392 , \54393 , \54394 , \54395 , \54396 ,
         \54397 , \54398 , \54399 , \54400 , \54401 , \54402 , \54403 , \54404 , \54405 , \54406 ,
         \54407 , \54408 , \54409 , \54410 , \54411 , \54412 , \54413 , \54414 , \54415 , \54416 ,
         \54417 , \54418 , \54419 , \54420 , \54421 , \54422 , \54423 , \54424 , \54425 , \54426 ,
         \54427 , \54428 , \54429 , \54430 , \54431 , \54432 , \54433 , \54434 , \54435 , \54436 ,
         \54437 , \54438 , \54439 , \54440 , \54441 , \54442 , \54443 , \54444 , \54445 , \54446 ,
         \54447 , \54448 , \54449 , \54450 , \54451 , \54452 , \54453 , \54454 , \54455 , \54456 ,
         \54457 , \54458 , \54459 , \54460 , \54461 , \54462 , \54463 , \54464 , \54465 , \54466 ,
         \54467 , \54468 , \54469 , \54470 , \54471 , \54472 , \54473 , \54474 , \54475 , \54476 ,
         \54477 , \54478 , \54479 , \54480 , \54481 , \54482 , \54483 , \54484 , \54485 , \54486 ,
         \54487 , \54488 , \54489 , \54490 , \54491 , \54492 , \54493 , \54494 , \54495 , \54496 ,
         \54497 , \54498 , \54499 , \54500 , \54501 , \54502 , \54503 , \54504 , \54505 , \54506 ,
         \54507 , \54508 , \54509 , \54510 , \54511 , \54512 , \54513 , \54514 , \54515 , \54516 ,
         \54517 , \54518 , \54519 , \54520 , \54521 , \54522 , \54523 , \54524 , \54525 , \54526 ,
         \54527 , \54528 , \54529 , \54530 , \54531 , \54532 , \54533 , \54534 , \54535 , \54536 ,
         \54537 , \54538 , \54539 , \54540 , \54541 , \54542 , \54543 , \54544 , \54545 , \54546 ,
         \54547 , \54548 , \54549 , \54550 , \54551 , \54552 , \54553 , \54554 , \54555 , \54556 ,
         \54557 , \54558 , \54559 , \54560 , \54561 , \54562 , \54563 , \54564 , \54565 , \54566 ,
         \54567 , \54568 , \54569 , \54570 , \54571 , \54572 , \54573 , \54574 , \54575 , \54576 ,
         \54577 , \54578 , \54579 , \54580 , \54581 , \54582 , \54583 , \54584 , \54585 , \54586 ,
         \54587 , \54588 , \54589 , \54590 , \54591 , \54592 , \54593 , \54594 , \54595 , \54596 ,
         \54597 , \54598 , \54599 , \54600 , \54601 , \54602 , \54603 , \54604 , \54605 , \54606 ,
         \54607 , \54608 , \54609 , \54610 , \54611 , \54612 , \54613 , \54614 , \54615 , \54616 ,
         \54617 , \54618 , \54619 , \54620 , \54621 , \54622 , \54623 , \54624 , \54625 , \54626 ,
         \54627 , \54628 , \54629 , \54630 , \54631 , \54632 , \54633 , \54634 , \54635 , \54636 ,
         \54637 , \54638 , \54639 , \54640 , \54641 , \54642 , \54643 , \54644 , \54645 , \54646 ,
         \54647 , \54648 , \54649 , \54650 , \54651 , \54652 , \54653 , \54654 , \54655 , \54656 ,
         \54657 , \54658 , \54659 , \54660 , \54661 , \54662 , \54663 , \54664 , \54665 , \54666 ,
         \54667 , \54668 , \54669 , \54670 , \54671 , \54672 , \54673 , \54674 , \54675 , \54676 ,
         \54677 , \54678 , \54679 , \54680 , \54681 , \54682 , \54683 , \54684 , \54685 , \54686 ,
         \54687 , \54688 , \54689 , \54690 , \54691 , \54692 , \54693 , \54694 , \54695 , \54696 ,
         \54697 , \54698 , \54699 , \54700 , \54701 , \54702 , \54703 , \54704 , \54705 , \54706 ,
         \54707 , \54708 , \54709 , \54710 , \54711 , \54712 , \54713 , \54714 , \54715 , \54716 ,
         \54717 , \54718 , \54719 , \54720 , \54721 , \54722 , \54723 , \54724 , \54725 , \54726 ,
         \54727 , \54728 , \54729 , \54730 , \54731 , \54732 , \54733 , \54734 , \54735 , \54736 ,
         \54737 , \54738 , \54739 , \54740 , \54741 , \54742 , \54743 , \54744 , \54745 , \54746 ,
         \54747 , \54748 , \54749 , \54750 , \54751 , \54752 , \54753 , \54754 , \54755 , \54756 ,
         \54757 , \54758 , \54759 , \54760 , \54761 , \54762 , \54763 , \54764 , \54765 , \54766 ,
         \54767 , \54768 , \54769 , \54770 , \54771 , \54772 , \54773 , \54774 , \54775 , \54776 ,
         \54777 , \54778 , \54779 , \54780 , \54781 , \54782 , \54783 , \54784 , \54785 , \54786 ,
         \54787 , \54788 , \54789 , \54790 , \54791 , \54792 , \54793 , \54794 , \54795 , \54796 ,
         \54797 , \54798 , \54799 , \54800 , \54801 , \54802 , \54803 , \54804 , \54805 , \54806 ,
         \54807 , \54808 , \54809 , \54810 , \54811 , \54812 , \54813 , \54814 , \54815 , \54816 ,
         \54817 , \54818 , \54819 , \54820 , \54821 , \54822 , \54823 , \54824 , \54825 , \54826 ,
         \54827 , \54828 , \54829 , \54830 , \54831 , \54832 , \54833 , \54834 , \54835 , \54836 ,
         \54837 , \54838 , \54839 , \54840 , \54841 , \54842 , \54843 , \54844 , \54845 , \54846 ,
         \54847 , \54848 , \54849 , \54850 , \54851 , \54852 , \54853 , \54854 , \54855 , \54856 ,
         \54857 , \54858 , \54859 , \54860 , \54861 , \54862 , \54863 , \54864 , \54865 , \54866 ,
         \54867 , \54868 , \54869 , \54870 , \54871 , \54872 , \54873 , \54874 , \54875 , \54876 ,
         \54877 , \54878 , \54879 , \54880 , \54881 , \54882 , \54883 , \54884 , \54885 , \54886 ,
         \54887 , \54888 , \54889 , \54890 , \54891 , \54892 , \54893 , \54894 , \54895 , \54896 ,
         \54897 , \54898 , \54899 , \54900 , \54901 , \54902 , \54903 , \54904 , \54905 , \54906 ,
         \54907 , \54908 , \54909 , \54910 , \54911 , \54912 , \54913 , \54914 , \54915 , \54916 ,
         \54917 , \54918 , \54919 , \54920 , \54921 , \54922 , \54923 , \54924 , \54925 , \54926 ,
         \54927 , \54928 , \54929 , \54930 , \54931 , \54932 , \54933 , \54934 , \54935 , \54936 ,
         \54937 , \54938 , \54939 , \54940 , \54941 , \54942 , \54943 , \54944 , \54945 , \54946 ,
         \54947 , \54948 , \54949 , \54950 , \54951 , \54952 , \54953 , \54954 , \54955 , \54956 ,
         \54957 , \54958 , \54959 , \54960 , \54961 , \54962 , \54963 , \54964 , \54965 , \54966 ,
         \54967 , \54968 , \54969 , \54970 , \54971 , \54972 , \54973 , \54974 , \54975 , \54976 ,
         \54977 , \54978 , \54979 , \54980 , \54981 , \54982 , \54983 , \54984 , \54985 , \54986 ,
         \54987 , \54988 , \54989 , \54990 , \54991 , \54992 , \54993 , \54994 , \54995 , \54996 ,
         \54997 , \54998 , \54999 , \55000 , \55001 , \55002 , \55003 , \55004 , \55005 , \55006 ,
         \55007 , \55008 , \55009 , \55010 , \55011 , \55012 , \55013 , \55014 , \55015 , \55016 ,
         \55017 , \55018 , \55019 , \55020 , \55021 , \55022 , \55023 , \55024 , \55025 , \55026 ,
         \55027 , \55028 , \55029 , \55030 , \55031 , \55032 , \55033 , \55034 , \55035 , \55036 ,
         \55037 , \55038 , \55039 , \55040 , \55041 , \55042 , \55043 , \55044 , \55045 , \55046 ,
         \55047 , \55048 , \55049 , \55050 , \55051 , \55052 , \55053 , \55054 , \55055 , \55056 ,
         \55057 , \55058 , \55059 , \55060 , \55061 , \55062 , \55063 , \55064 , \55065 , \55066 ,
         \55067 , \55068 , \55069 , \55070 , \55071 , \55072 , \55073 , \55074 , \55075 , \55076 ,
         \55077 , \55078 , \55079 , \55080 , \55081 , \55082 , \55083 , \55084 , \55085 , \55086 ,
         \55087 , \55088 , \55089 , \55090 , \55091 , \55092 , \55093 , \55094 , \55095 , \55096 ,
         \55097 , \55098 , \55099 , \55100 , \55101 , \55102 , \55103 , \55104 , \55105 , \55106 ,
         \55107 , \55108 , \55109 , \55110 , \55111 , \55112 , \55113 , \55114 , \55115 , \55116 ,
         \55117 , \55118 , \55119 , \55120 , \55121 , \55122 , \55123 , \55124 , \55125 , \55126 ,
         \55127 , \55128 , \55129 , \55130 , \55131 , \55132 , \55133 , \55134 , \55135 , \55136 ,
         \55137 , \55138 , \55139 , \55140 , \55141 , \55142 , \55143 , \55144 , \55145 , \55146 ,
         \55147 , \55148 , \55149 , \55150 , \55151 , \55152 , \55153 , \55154 , \55155 , \55156 ,
         \55157 , \55158 , \55159 , \55160 , \55161 , \55162 , \55163 , \55164 , \55165 , \55166 ,
         \55167 , \55168 , \55169 , \55170 , \55171 , \55172 , \55173 , \55174 , \55175 , \55176 ,
         \55177 , \55178 , \55179 , \55180 , \55181 , \55182 , \55183 , \55184 , \55185 , \55186 ,
         \55187 , \55188 , \55189 , \55190 , \55191 , \55192 , \55193 , \55194 , \55195 , \55196 ,
         \55197 , \55198 , \55199 , \55200 , \55201 , \55202 , \55203 , \55204 , \55205 , \55206 ,
         \55207 , \55208 , \55209 , \55210 , \55211 , \55212 , \55213 , \55214 , \55215 , \55216 ,
         \55217 , \55218 , \55219 , \55220 , \55221 , \55222 , \55223 , \55224 , \55225 , \55226 ,
         \55227 , \55228 , \55229 , \55230 , \55231 , \55232 , \55233 , \55234 , \55235 , \55236 ,
         \55237 , \55238 , \55239 , \55240 , \55241 , \55242 , \55243 , \55244 , \55245 , \55246 ,
         \55247 , \55248 , \55249 , \55250 , \55251 , \55252 , \55253 , \55254 , \55255 , \55256 ,
         \55257 , \55258 , \55259 , \55260 , \55261 , \55262 , \55263 , \55264 , \55265 , \55266 ,
         \55267 , \55268 , \55269 , \55270 , \55271 , \55272 , \55273 , \55274 , \55275 , \55276 ,
         \55277 , \55278 , \55279 , \55280 , \55281 , \55282 , \55283 , \55284 , \55285 , \55286 ,
         \55287 , \55288 , \55289 , \55290 , \55291 , \55292 , \55293 , \55294 , \55295 , \55296 ,
         \55297 , \55298 , \55299 , \55300 , \55301 , \55302 , \55303 , \55304 , \55305 , \55306 ,
         \55307 , \55308 , \55309 , \55310 , \55311 , \55312 , \55313 , \55314 , \55315 , \55316 ,
         \55317 , \55318 , \55319 , \55320 , \55321 , \55322 , \55323 , \55324 , \55325 , \55326 ,
         \55327 , \55328 , \55329 , \55330 , \55331 , \55332 , \55333 , \55334 , \55335 , \55336 ,
         \55337 , \55338 , \55339 , \55340 , \55341 , \55342 , \55343 , \55344 , \55345 , \55346 ,
         \55347 , \55348 , \55349 , \55350 , \55351 , \55352 , \55353 , \55354 , \55355 , \55356 ,
         \55357 , \55358 , \55359 , \55360 , \55361 , \55362 , \55363 , \55364 , \55365 , \55366 ,
         \55367 , \55368 , \55369 , \55370 , \55371 , \55372 , \55373 , \55374 , \55375 , \55376 ,
         \55377 , \55378 , \55379 , \55380 , \55381 , \55382 , \55383 , \55384 , \55385 , \55386 ,
         \55387 , \55388 , \55389 , \55390 , \55391 , \55392 , \55393 , \55394 , \55395 , \55396 ,
         \55397 , \55398 , \55399 , \55400 , \55401 , \55402 , \55403 , \55404 , \55405 , \55406 ,
         \55407 , \55408 , \55409 , \55410 , \55411 , \55412 , \55413 , \55414 , \55415 , \55416 ,
         \55417 , \55418 , \55419 , \55420 , \55421 , \55422 , \55423 , \55424 , \55425 , \55426 ,
         \55427 , \55428 , \55429 , \55430 , \55431 , \55432 , \55433 , \55434 , \55435 , \55436 ,
         \55437 , \55438 , \55439 , \55440 , \55441 , \55442 , \55443 , \55444 , \55445 , \55446 ,
         \55447 , \55448 , \55449 , \55450 , \55451 , \55452 , \55453 , \55454 , \55455 , \55456 ,
         \55457 , \55458 , \55459 , \55460 , \55461 , \55462 , \55463 , \55464 , \55465 , \55466 ,
         \55467 , \55468 , \55469 , \55470 , \55471 , \55472 , \55473 , \55474 , \55475 , \55476 ,
         \55477 , \55478 , \55479 , \55480 , \55481 , \55482 , \55483 , \55484 , \55485 , \55486 ,
         \55487 , \55488 , \55489 , \55490 , \55491 , \55492 , \55493 , \55494 , \55495 , \55496 ,
         \55497 , \55498 , \55499 , \55500 , \55501 , \55502 , \55503 , \55504 , \55505 , \55506 ,
         \55507 , \55508 , \55509 , \55510 , \55511 , \55512 , \55513 , \55514 , \55515 , \55516 ,
         \55517 , \55518 , \55519 , \55520 , \55521 , \55522 , \55523 , \55524 , \55525 , \55526 ,
         \55527 , \55528 , \55529 , \55530 , \55531 , \55532 , \55533 , \55534 , \55535 , \55536 ,
         \55537 , \55538 , \55539 , \55540 , \55541 , \55542 , \55543 , \55544 , \55545 , \55546 ,
         \55547 , \55548 , \55549 , \55550 , \55551 , \55552 , \55553 , \55554 , \55555 , \55556 ,
         \55557 , \55558 , \55559 , \55560 , \55561 , \55562 , \55563 , \55564 , \55565 , \55566 ,
         \55567 , \55568 , \55569 , \55570 , \55571 , \55572 , \55573 , \55574 , \55575 , \55576 ,
         \55577 , \55578 , \55579 , \55580 , \55581 , \55582 , \55583 , \55584 , \55585 , \55586 ,
         \55587 , \55588 , \55589 , \55590 , \55591 , \55592 , \55593 , \55594 , \55595 , \55596 ,
         \55597 , \55598 , \55599 , \55600 , \55601 , \55602 , \55603 , \55604 , \55605 , \55606 ,
         \55607 , \55608 , \55609 , \55610 , \55611 , \55612 , \55613 , \55614 , \55615 , \55616 ,
         \55617 , \55618 , \55619 , \55620 , \55621 , \55622 , \55623 , \55624 , \55625 , \55626 ,
         \55627 , \55628 , \55629 , \55630 , \55631 , \55632 , \55633 , \55634 , \55635 , \55636 ,
         \55637 , \55638 , \55639 , \55640 , \55641 , \55642 , \55643 , \55644 , \55645 , \55646 ,
         \55647 , \55648 , \55649 , \55650 , \55651 , \55652 , \55653 , \55654 , \55655 , \55656 ,
         \55657 , \55658 , \55659 , \55660 , \55661 , \55662 , \55663 , \55664 , \55665 , \55666 ,
         \55667 , \55668 , \55669 , \55670 , \55671 , \55672 , \55673 , \55674 , \55675 , \55676 ,
         \55677 , \55678 , \55679 , \55680 , \55681 , \55682 , \55683 , \55684 , \55685 , \55686 ,
         \55687 , \55688 , \55689 , \55690 , \55691 , \55692 , \55693 , \55694 , \55695 , \55696 ,
         \55697 , \55698 , \55699 , \55700 , \55701 , \55702 , \55703 , \55704 , \55705 , \55706 ,
         \55707 , \55708 , \55709 , \55710 , \55711 , \55712 , \55713 , \55714 , \55715 , \55716 ,
         \55717 , \55718 , \55719 , \55720 , \55721 , \55722 , \55723 , \55724 , \55725 , \55726 ,
         \55727 , \55728 , \55729 , \55730 , \55731 , \55732 , \55733 , \55734 , \55735 , \55736 ,
         \55737 , \55738 , \55739 , \55740 , \55741 , \55742 , \55743 , \55744 , \55745 , \55746 ,
         \55747 , \55748 , \55749 , \55750 , \55751 , \55752 , \55753 , \55754 , \55755 , \55756 ,
         \55757 , \55758 , \55759 , \55760 , \55761 , \55762 , \55763 , \55764 , \55765 , \55766 ,
         \55767 , \55768 , \55769 , \55770 , \55771 , \55772 , \55773 , \55774 , \55775 , \55776 ,
         \55777 , \55778 , \55779 , \55780 , \55781 , \55782 , \55783 , \55784 , \55785 , \55786 ,
         \55787 , \55788 , \55789 , \55790 , \55791 , \55792 , \55793 , \55794 , \55795 , \55796 ,
         \55797 , \55798 , \55799 , \55800 , \55801 , \55802 , \55803 , \55804 , \55805 , \55806 ,
         \55807 , \55808 , \55809 , \55810 , \55811 , \55812 , \55813 , \55814 , \55815 , \55816 ,
         \55817 , \55818 , \55819 , \55820 , \55821 , \55822 , \55823 , \55824 , \55825 , \55826 ,
         \55827 , \55828 , \55829 , \55830 , \55831 , \55832 , \55833 , \55834 , \55835 , \55836 ,
         \55837 , \55838 , \55839 , \55840 , \55841 , \55842 , \55843 , \55844 , \55845 , \55846 ,
         \55847 , \55848 , \55849 , \55850 , \55851 , \55852 , \55853 , \55854 , \55855 , \55856 ,
         \55857 , \55858 , \55859 , \55860 , \55861 , \55862 , \55863 , \55864 , \55865 , \55866 ,
         \55867 , \55868 , \55869 , \55870 , \55871 , \55872 , \55873 , \55874 , \55875 , \55876 ,
         \55877 , \55878 , \55879 , \55880 , \55881 , \55882 , \55883 , \55884 , \55885 , \55886 ,
         \55887 , \55888 , \55889 , \55890 , \55891 , \55892 , \55893 , \55894 , \55895 , \55896 ,
         \55897 , \55898 , \55899 , \55900 , \55901 , \55902 , \55903 , \55904 , \55905 , \55906 ,
         \55907 , \55908 , \55909 , \55910 , \55911 , \55912 , \55913 , \55914 , \55915 , \55916 ,
         \55917 , \55918 , \55919 , \55920 , \55921 , \55922 , \55923 , \55924 , \55925 , \55926 ,
         \55927 , \55928 , \55929 , \55930 , \55931 , \55932 , \55933 , \55934 , \55935 , \55936 ,
         \55937 , \55938 , \55939 , \55940 , \55941 , \55942 , \55943 , \55944 , \55945 , \55946 ,
         \55947 , \55948 , \55949 , \55950 , \55951 , \55952 , \55953 , \55954 , \55955 , \55956 ,
         \55957 , \55958 , \55959 , \55960 , \55961 , \55962 , \55963 , \55964 , \55965 , \55966 ,
         \55967 , \55968 , \55969 , \55970 , \55971 , \55972 , \55973 , \55974 , \55975 , \55976 ,
         \55977 , \55978 , \55979 , \55980 , \55981 , \55982 , \55983 , \55984 , \55985 , \55986 ,
         \55987 , \55988 , \55989 , \55990 , \55991 , \55992 , \55993 , \55994 , \55995 , \55996 ,
         \55997 , \55998 , \55999 , \56000 , \56001 , \56002 , \56003 , \56004 , \56005 , \56006 ,
         \56007 , \56008 , \56009 , \56010 , \56011 , \56012 , \56013 , \56014 , \56015 , \56016 ,
         \56017 , \56018 , \56019 , \56020 , \56021 , \56022 , \56023 , \56024 , \56025 , \56026 ,
         \56027 , \56028 , \56029 , \56030 , \56031 , \56032 , \56033 , \56034 , \56035 , \56036 ,
         \56037 , \56038 , \56039 , \56040 , \56041 , \56042 , \56043 , \56044 , \56045 , \56046 ,
         \56047 , \56048 , \56049 , \56050 , \56051 , \56052 , \56053 , \56054 , \56055 , \56056 ,
         \56057 , \56058 , \56059 , \56060 , \56061 , \56062 , \56063 , \56064 , \56065 , \56066 ,
         \56067 , \56068 , \56069 , \56070 , \56071 , \56072 , \56073 , \56074 , \56075 , \56076 ,
         \56077 , \56078 , \56079 , \56080 , \56081 , \56082 , \56083 , \56084 , \56085 , \56086 ,
         \56087 , \56088 , \56089 , \56090 , \56091 , \56092 , \56093 , \56094 , \56095 , \56096 ,
         \56097 , \56098 , \56099 , \56100 , \56101 , \56102 , \56103 , \56104 , \56105 , \56106 ,
         \56107 , \56108 , \56109 , \56110 , \56111 , \56112 , \56113 , \56114 , \56115 , \56116 ,
         \56117 , \56118 , \56119 , \56120 , \56121 , \56122 , \56123 , \56124 , \56125 , \56126 ,
         \56127 , \56128 , \56129 , \56130 , \56131 , \56132 , \56133 , \56134 , \56135 , \56136 ,
         \56137 , \56138 , \56139 , \56140 , \56141 , \56142 , \56143 , \56144 , \56145 , \56146 ,
         \56147 , \56148 , \56149 , \56150 , \56151 , \56152 , \56153 , \56154 , \56155 , \56156 ,
         \56157 , \56158 , \56159 , \56160 , \56161 , \56162 , \56163 , \56164 , \56165 , \56166 ,
         \56167 , \56168 , \56169 , \56170 , \56171 , \56172 , \56173 , \56174 , \56175 , \56176 ,
         \56177 , \56178 , \56179 , \56180 , \56181 , \56182 , \56183 , \56184 , \56185 , \56186 ,
         \56187 , \56188 , \56189 , \56190 , \56191 , \56192 , \56193 , \56194 , \56195 , \56196 ,
         \56197 , \56198 , \56199 , \56200 , \56201 , \56202 , \56203 , \56204 , \56205 , \56206 ,
         \56207 , \56208 , \56209 , \56210 , \56211 , \56212 , \56213 , \56214 , \56215 , \56216 ,
         \56217 , \56218 , \56219 , \56220 , \56221 , \56222 , \56223 , \56224 , \56225 , \56226 ,
         \56227 , \56228 , \56229 , \56230 , \56231 , \56232 , \56233 , \56234 , \56235 , \56236 ,
         \56237 , \56238 , \56239 , \56240 , \56241 , \56242 , \56243 , \56244 , \56245 , \56246 ,
         \56247 , \56248 , \56249 , \56250 , \56251 , \56252 , \56253 , \56254 , \56255 , \56256 ,
         \56257 , \56258 , \56259 , \56260 , \56261 , \56262 , \56263 , \56264 , \56265 , \56266 ,
         \56267 , \56268 , \56269 , \56270 , \56271 , \56272 , \56273 , \56274 , \56275 , \56276 ,
         \56277 , \56278 , \56279 , \56280 , \56281 , \56282 , \56283 , \56284 , \56285 , \56286 ,
         \56287 , \56288 , \56289 , \56290 , \56291 , \56292 , \56293 , \56294 , \56295 , \56296 ,
         \56297 , \56298 , \56299 , \56300 , \56301 , \56302 , \56303 , \56304 , \56305 , \56306 ,
         \56307 , \56308 , \56309 , \56310 , \56311 , \56312 , \56313 , \56314 , \56315 , \56316 ,
         \56317 , \56318 , \56319 , \56320 , \56321 , \56322 , \56323 , \56324 , \56325 , \56326 ,
         \56327 , \56328 , \56329 , \56330 , \56331 , \56332 , \56333 , \56334 , \56335 , \56336 ,
         \56337 , \56338 , \56339 , \56340 , \56341 , \56342 , \56343 , \56344 , \56345 , \56346 ,
         \56347 , \56348 , \56349 , \56350 , \56351 , \56352 , \56353 , \56354 , \56355 , \56356 ,
         \56357 , \56358 , \56359 , \56360 , \56361 , \56362 , \56363 , \56364 , \56365 , \56366 ,
         \56367 , \56368 , \56369 , \56370 , \56371 , \56372 , \56373 , \56374 , \56375 , \56376 ,
         \56377 , \56378 , \56379 , \56380 , \56381 , \56382 , \56383 , \56384 , \56385 , \56386 ,
         \56387 , \56388 , \56389 , \56390 , \56391 , \56392 , \56393 , \56394 , \56395 , \56396 ,
         \56397 , \56398 , \56399 , \56400 , \56401 , \56402 , \56403 , \56404 , \56405 , \56406 ,
         \56407 , \56408 , \56409 , \56410 , \56411 , \56412 , \56413 , \56414 , \56415 , \56416 ,
         \56417 , \56418 , \56419 , \56420 , \56421 , \56422 , \56423 , \56424 , \56425 , \56426 ,
         \56427 , \56428 , \56429 , \56430 , \56431 , \56432 , \56433 , \56434 , \56435 , \56436 ,
         \56437 , \56438 , \56439 , \56440 , \56441 , \56442 , \56443 , \56444 , \56445 , \56446 ,
         \56447 , \56448 , \56449 , \56450 , \56451 , \56452 , \56453 , \56454 , \56455 , \56456 ,
         \56457 , \56458 , \56459 , \56460 , \56461 , \56462 , \56463 , \56464 , \56465 , \56466 ,
         \56467 , \56468 , \56469 , \56470 , \56471 , \56472 , \56473 , \56474 , \56475 , \56476 ,
         \56477 , \56478 , \56479 , \56480 , \56481 , \56482 , \56483 , \56484 , \56485 , \56486 ,
         \56487 , \56488 , \56489 , \56490 , \56491 , \56492 , \56493 , \56494 , \56495 , \56496 ,
         \56497 , \56498 , \56499 , \56500 , \56501 , \56502 , \56503 , \56504 , \56505 , \56506 ,
         \56507 , \56508 , \56509 , \56510 , \56511 , \56512 , \56513 , \56514 , \56515 , \56516 ,
         \56517 , \56518 , \56519 , \56520 , \56521 , \56522 , \56523 , \56524 , \56525 , \56526 ,
         \56527 , \56528 , \56529 , \56530 , \56531 , \56532 , \56533 , \56534 , \56535 , \56536 ,
         \56537 , \56538 , \56539 , \56540 , \56541 , \56542 , \56543 , \56544 , \56545 , \56546 ,
         \56547 , \56548 , \56549 , \56550 , \56551 , \56552 , \56553 , \56554 , \56555 , \56556 ,
         \56557 , \56558 , \56559 , \56560 , \56561 , \56562 , \56563 , \56564 , \56565 , \56566 ,
         \56567 , \56568 , \56569 , \56570 , \56571 , \56572 , \56573 , \56574 , \56575 , \56576 ,
         \56577 , \56578 , \56579 , \56580 , \56581 , \56582 , \56583 , \56584 , \56585 , \56586 ,
         \56587 , \56588 , \56589 , \56590 , \56591 , \56592 , \56593 , \56594 , \56595 , \56596 ,
         \56597 , \56598 , \56599 , \56600 , \56601 , \56602 , \56603 , \56604 , \56605 , \56606 ,
         \56607 , \56608 , \56609 , \56610 , \56611 , \56612 , \56613 , \56614 , \56615 , \56616 ,
         \56617 , \56618 , \56619 , \56620 , \56621 , \56622 , \56623 , \56624 , \56625 , \56626 ,
         \56627 , \56628 , \56629 , \56630 , \56631 , \56632 , \56633 , \56634 , \56635 , \56636 ,
         \56637 , \56638 , \56639 , \56640 , \56641 , \56642 , \56643 , \56644 , \56645 , \56646 ,
         \56647 , \56648 , \56649 , \56650 , \56651 , \56652 , \56653 , \56654 , \56655 , \56656 ,
         \56657 , \56658 , \56659 , \56660 , \56661 , \56662 , \56663 , \56664 , \56665 , \56666 ,
         \56667 , \56668 , \56669 , \56670 , \56671 , \56672 , \56673 , \56674 , \56675 , \56676 ,
         \56677 , \56678 , \56679 , \56680 , \56681 , \56682 , \56683 , \56684 , \56685 , \56686 ,
         \56687 , \56688 , \56689 , \56690 , \56691 , \56692 , \56693 , \56694 , \56695 , \56696 ,
         \56697 , \56698 , \56699 , \56700 , \56701 , \56702 , \56703 , \56704 , \56705 , \56706 ,
         \56707 , \56708 , \56709 , \56710 , \56711 , \56712 , \56713 , \56714 , \56715 , \56716 ,
         \56717 , \56718 , \56719 , \56720 , \56721 , \56722 , \56723 , \56724 , \56725 , \56726 ,
         \56727 , \56728 , \56729 , \56730 , \56731 , \56732 , \56733 , \56734 , \56735 , \56736 ,
         \56737 , \56738 , \56739 , \56740 , \56741 , \56742 , \56743 , \56744 , \56745 , \56746 ,
         \56747 , \56748 , \56749 , \56750 , \56751 , \56752 , \56753 , \56754 , \56755 , \56756 ,
         \56757 , \56758 , \56759 , \56760 , \56761 , \56762 , \56763 , \56764 , \56765 , \56766 ,
         \56767 , \56768 , \56769 , \56770 , \56771 , \56772 , \56773 , \56774 , \56775 , \56776 ,
         \56777 , \56778 , \56779 , \56780 , \56781 , \56782 , \56783 , \56784 , \56785 , \56786 ,
         \56787 , \56788 , \56789 , \56790 , \56791 , \56792 , \56793 , \56794 , \56795 , \56796 ,
         \56797 , \56798 , \56799 , \56800 , \56801 , \56802 , \56803 , \56804 , \56805 , \56806 ,
         \56807 , \56808 , \56809 , \56810 , \56811 , \56812 , \56813 , \56814 , \56815 , \56816 ,
         \56817 , \56818 , \56819 , \56820 , \56821 , \56822 , \56823 , \56824 , \56825 , \56826 ,
         \56827 , \56828 , \56829 , \56830 , \56831 , \56832 , \56833 , \56834 , \56835 , \56836 ,
         \56837 , \56838 , \56839 , \56840 , \56841 , \56842 , \56843 , \56844 , \56845 , \56846 ,
         \56847 , \56848 , \56849 , \56850 , \56851 , \56852 , \56853 , \56854 , \56855 , \56856 ,
         \56857 , \56858 , \56859 , \56860 , \56861 , \56862 , \56863 , \56864 , \56865 , \56866 ,
         \56867 , \56868 , \56869 , \56870 , \56871 , \56872 , \56873 , \56874 , \56875 , \56876 ,
         \56877 , \56878 , \56879 , \56880 , \56881 , \56882 , \56883 , \56884 , \56885 , \56886 ,
         \56887 , \56888 , \56889 , \56890 , \56891 , \56892 , \56893 , \56894 , \56895 , \56896 ,
         \56897 , \56898 , \56899 , \56900 , \56901 , \56902 , \56903 , \56904 , \56905 , \56906 ,
         \56907 , \56908 , \56909 , \56910 , \56911 , \56912 , \56913 , \56914 , \56915 , \56916 ,
         \56917 , \56918 , \56919 , \56920 , \56921 , \56922 , \56923 , \56924 , \56925 , \56926 ,
         \56927 , \56928 , \56929 , \56930 , \56931 , \56932 , \56933 , \56934 , \56935 , \56936 ,
         \56937 , \56938 , \56939 , \56940 , \56941 , \56942 , \56943 , \56944 , \56945 , \56946 ,
         \56947 , \56948 , \56949 , \56950 , \56951 , \56952 , \56953 , \56954 , \56955 , \56956 ,
         \56957 , \56958 , \56959 , \56960 , \56961 , \56962 , \56963 , \56964 , \56965 , \56966 ,
         \56967 , \56968 , \56969 , \56970 , \56971 , \56972 , \56973 , \56974 , \56975 , \56976 ,
         \56977 , \56978 , \56979 , \56980 , \56981 , \56982 , \56983 , \56984 , \56985 , \56986 ,
         \56987 , \56988 , \56989 , \56990 , \56991 , \56992 , \56993 , \56994 , \56995 , \56996 ,
         \56997 , \56998 , \56999 , \57000 , \57001 , \57002 , \57003 , \57004 , \57005 , \57006 ,
         \57007 , \57008 , \57009 , \57010 , \57011 , \57012 , \57013 , \57014 , \57015 , \57016 ,
         \57017 , \57018 , \57019 , \57020 , \57021 , \57022 , \57023 , \57024 , \57025 , \57026 ,
         \57027 , \57028 , \57029 , \57030 , \57031 , \57032 , \57033 , \57034 , \57035 , \57036 ,
         \57037 , \57038 , \57039 , \57040 , \57041 , \57042 , \57043 , \57044 , \57045 , \57046 ,
         \57047 , \57048 , \57049 , \57050 , \57051 , \57052 , \57053 , \57054 , \57055 , \57056 ,
         \57057 , \57058 , \57059 , \57060 , \57061 , \57062 , \57063 , \57064 , \57065 , \57066 ,
         \57067 , \57068 , \57069 , \57070 , \57071 , \57072 , \57073 , \57074 , \57075 , \57076 ,
         \57077 , \57078 , \57079 , \57080 , \57081 , \57082 , \57083 , \57084 , \57085 , \57086 ,
         \57087 , \57088 , \57089 , \57090 , \57091 , \57092 , \57093 , \57094 , \57095 , \57096 ,
         \57097 , \57098 , \57099 , \57100 , \57101 , \57102 , \57103 , \57104 , \57105 , \57106 ,
         \57107 , \57108 , \57109 , \57110 , \57111 , \57112 , \57113 , \57114 , \57115 , \57116 ,
         \57117 , \57118 , \57119 , \57120 , \57121 , \57122 , \57123 , \57124 , \57125 , \57126 ,
         \57127 , \57128 , \57129 , \57130 , \57131 , \57132 , \57133 , \57134 , \57135 , \57136 ,
         \57137 , \57138 , \57139 , \57140 , \57141 , \57142 , \57143 , \57144 , \57145 , \57146 ,
         \57147 , \57148 , \57149 , \57150 , \57151 , \57152 , \57153 , \57154 , \57155 , \57156 ,
         \57157 , \57158 , \57159 , \57160 , \57161 , \57162 , \57163 , \57164 , \57165 , \57166 ,
         \57167 , \57168 , \57169 , \57170 , \57171 , \57172 , \57173 , \57174 , \57175 , \57176 ,
         \57177 , \57178 , \57179 , \57180 , \57181 , \57182 , \57183 , \57184 , \57185 , \57186 ,
         \57187 , \57188 , \57189 , \57190 , \57191 , \57192 , \57193 , \57194 , \57195 , \57196 ,
         \57197 , \57198 , \57199 , \57200 , \57201 , \57202 , \57203 , \57204 , \57205 , \57206 ,
         \57207 , \57208 , \57209 , \57210 , \57211 , \57212 , \57213 , \57214 , \57215 , \57216 ,
         \57217 , \57218 , \57219 , \57220 , \57221 , \57222 , \57223 , \57224 , \57225 , \57226 ,
         \57227 , \57228 , \57229 , \57230 , \57231 , \57232 , \57233 , \57234 , \57235 , \57236 ,
         \57237 , \57238 , \57239 , \57240 , \57241 , \57242 , \57243 , \57244 , \57245 , \57246 ,
         \57247 , \57248 , \57249 , \57250 , \57251 , \57252 , \57253 , \57254 , \57255 , \57256 ,
         \57257 , \57258 , \57259 , \57260 , \57261 , \57262 , \57263 , \57264 , \57265 , \57266 ,
         \57267 , \57268 , \57269 , \57270 , \57271 , \57272 , \57273 , \57274 , \57275 , \57276 ,
         \57277 , \57278 , \57279 , \57280 , \57281 , \57282 , \57283 , \57284 , \57285 , \57286 ,
         \57287 , \57288 , \57289 , \57290 , \57291 , \57292 , \57293 , \57294 , \57295 , \57296 ,
         \57297 , \57298 , \57299 , \57300 , \57301 , \57302 , \57303 , \57304 , \57305 , \57306 ,
         \57307 , \57308 , \57309 , \57310 , \57311 , \57312 , \57313 , \57314 , \57315 , \57316 ,
         \57317 , \57318 , \57319 , \57320 , \57321 , \57322 , \57323 , \57324 , \57325 , \57326 ,
         \57327 , \57328 , \57329 , \57330 , \57331 , \57332 , \57333 , \57334 , \57335 , \57336 ,
         \57337 , \57338 , \57339 , \57340 , \57341 , \57342 , \57343 , \57344 , \57345 , \57346 ,
         \57347 , \57348 , \57349 , \57350 , \57351 , \57352 , \57353 , \57354 , \57355 , \57356 ,
         \57357 , \57358 , \57359 , \57360 , \57361 , \57362 , \57363 , \57364 , \57365 , \57366 ,
         \57367 , \57368 , \57369 , \57370 , \57371 , \57372 , \57373 , \57374 , \57375 , \57376 ,
         \57377 , \57378 , \57379 , \57380 , \57381 , \57382 , \57383 , \57384 , \57385 , \57386 ,
         \57387 , \57388 , \57389 , \57390 , \57391 , \57392 , \57393 , \57394 , \57395 , \57396 ,
         \57397 , \57398 , \57399 , \57400 , \57401 , \57402 , \57403 , \57404 , \57405 , \57406 ,
         \57407 , \57408 , \57409 , \57410 , \57411 , \57412 , \57413 , \57414 , \57415 , \57416 ,
         \57417 , \57418 , \57419 , \57420 , \57421 , \57422 , \57423 , \57424 , \57425 , \57426 ,
         \57427 , \57428 , \57429 , \57430 , \57431 , \57432 , \57433 , \57434 , \57435 , \57436 ,
         \57437 , \57438 , \57439 , \57440 , \57441 , \57442 , \57443 , \57444 , \57445 , \57446 ,
         \57447 , \57448 , \57449 , \57450 , \57451 , \57452 , \57453 , \57454 , \57455 , \57456 ,
         \57457 , \57458 , \57459 , \57460 , \57461 , \57462 , \57463 , \57464 , \57465 , \57466 ,
         \57467 , \57468 , \57469 , \57470 , \57471 , \57472 , \57473 , \57474 , \57475 , \57476 ,
         \57477 , \57478 , \57479 , \57480 , \57481 , \57482 , \57483 , \57484 , \57485 , \57486 ,
         \57487 , \57488 , \57489 , \57490 , \57491 , \57492 , \57493 , \57494 , \57495 , \57496 ,
         \57497 , \57498 , \57499 , \57500 , \57501 , \57502 , \57503 , \57504 , \57505 , \57506 ,
         \57507 , \57508 , \57509 , \57510 , \57511 , \57512 , \57513 , \57514 , \57515 , \57516 ,
         \57517 , \57518 , \57519 , \57520 , \57521 , \57522 , \57523 , \57524 , \57525 , \57526 ,
         \57527 , \57528 , \57529 , \57530 , \57531 , \57532 , \57533 , \57534 , \57535 , \57536 ,
         \57537 , \57538 , \57539 , \57540 , \57541 , \57542 , \57543 , \57544 , \57545 , \57546 ,
         \57547 , \57548 , \57549 , \57550 , \57551 , \57552 , \57553 , \57554 , \57555 , \57556 ,
         \57557 , \57558 , \57559 , \57560 , \57561 , \57562 , \57563 , \57564 , \57565 , \57566 ,
         \57567 , \57568 , \57569 , \57570 , \57571 , \57572 , \57573 , \57574 , \57575 , \57576 ,
         \57577 , \57578 , \57579 , \57580 , \57581 , \57582 , \57583 , \57584 , \57585 , \57586 ,
         \57587 , \57588 , \57589 , \57590 , \57591 , \57592 , \57593 , \57594 , \57595 , \57596 ,
         \57597 , \57598 , \57599 , \57600 , \57601 , \57602 , \57603 , \57604 , \57605 , \57606 ,
         \57607 , \57608 , \57609 , \57610 , \57611 , \57612 , \57613 , \57614 , \57615 , \57616 ,
         \57617 , \57618 , \57619 , \57620 , \57621 , \57622 , \57623 , \57624 , \57625 , \57626 ,
         \57627 , \57628 , \57629 , \57630 , \57631 , \57632 , \57633 , \57634 , \57635 , \57636 ,
         \57637 , \57638 , \57639 , \57640 , \57641 , \57642 , \57643 , \57644 , \57645 , \57646 ,
         \57647 , \57648 , \57649 , \57650 , \57651 , \57652 , \57653 , \57654 , \57655 , \57656 ,
         \57657 , \57658 , \57659 , \57660 , \57661 , \57662 , \57663 , \57664 , \57665 , \57666 ,
         \57667 , \57668 , \57669 , \57670 , \57671 , \57672 , \57673 , \57674 , \57675 , \57676 ,
         \57677 , \57678 , \57679 , \57680 , \57681 , \57682 , \57683 , \57684 , \57685 , \57686 ,
         \57687 , \57688 , \57689 , \57690 , \57691 , \57692 , \57693 , \57694 , \57695 , \57696 ,
         \57697 , \57698 , \57699 , \57700 , \57701 , \57702 , \57703 , \57704 , \57705 , \57706 ,
         \57707 , \57708 , \57709 , \57710 , \57711 , \57712 , \57713 , \57714 , \57715 , \57716 ,
         \57717 , \57718 , \57719 , \57720 , \57721 , \57722 , \57723 , \57724 , \57725 , \57726 ,
         \57727 , \57728 , \57729 , \57730 , \57731 , \57732 , \57733 , \57734 , \57735 , \57736 ,
         \57737 , \57738 , \57739 , \57740 , \57741 , \57742 , \57743 , \57744 , \57745 , \57746 ,
         \57747 , \57748 , \57749 , \57750 , \57751 , \57752 , \57753 , \57754 , \57755 , \57756 ,
         \57757 , \57758 , \57759 , \57760 , \57761 , \57762 , \57763 , \57764 , \57765 , \57766 ,
         \57767 , \57768 , \57769 , \57770 , \57771 , \57772 , \57773 , \57774 , \57775 , \57776 ,
         \57777 , \57778 , \57779 , \57780 , \57781 , \57782 , \57783 , \57784 , \57785 , \57786 ,
         \57787 , \57788 , \57789 , \57790 , \57791 , \57792 , \57793 , \57794 , \57795 , \57796 ,
         \57797 , \57798 , \57799 , \57800 , \57801 , \57802 , \57803 , \57804 , \57805 , \57806 ,
         \57807 , \57808 , \57809 , \57810 , \57811 , \57812 , \57813 , \57814 , \57815 , \57816 ,
         \57817 , \57818 , \57819 , \57820 , \57821 , \57822 , \57823 , \57824 , \57825 , \57826 ,
         \57827 , \57828 , \57829 , \57830 , \57831 , \57832 , \57833 , \57834 , \57835 , \57836 ,
         \57837 , \57838 , \57839 , \57840 , \57841 , \57842 , \57843 , \57844 , \57845 , \57846 ,
         \57847 , \57848 , \57849 , \57850 , \57851 , \57852 , \57853 , \57854 , \57855 , \57856 ,
         \57857 , \57858 , \57859 , \57860 , \57861 , \57862 , \57863 , \57864 , \57865 , \57866 ,
         \57867 , \57868 , \57869 , \57870 , \57871 , \57872 , \57873 , \57874 , \57875 , \57876 ,
         \57877 , \57878 , \57879 , \57880 , \57881 , \57882 , \57883 , \57884 , \57885 , \57886 ,
         \57887 , \57888 , \57889 , \57890 , \57891 , \57892 , \57893 , \57894 , \57895 , \57896 ,
         \57897 , \57898 , \57899 , \57900 , \57901 , \57902 , \57903 , \57904 , \57905 , \57906 ,
         \57907 , \57908 , \57909 , \57910 , \57911 , \57912 , \57913 , \57914 , \57915 , \57916 ,
         \57917 , \57918 , \57919 , \57920 , \57921 , \57922 , \57923 , \57924 , \57925 , \57926 ,
         \57927 , \57928 , \57929 , \57930 , \57931 , \57932 , \57933 , \57934 , \57935 , \57936 ,
         \57937 , \57938 , \57939 , \57940 , \57941 , \57942 , \57943 , \57944 , \57945 , \57946 ,
         \57947 , \57948 , \57949 , \57950 , \57951 , \57952 , \57953 , \57954 , \57955 , \57956 ,
         \57957 , \57958 , \57959 , \57960 , \57961 , \57962 , \57963 , \57964 , \57965 , \57966 ,
         \57967 , \57968 , \57969 , \57970 , \57971 , \57972 , \57973 , \57974 , \57975 , \57976 ,
         \57977 , \57978 , \57979 , \57980 , \57981 , \57982 , \57983 , \57984 , \57985 , \57986 ,
         \57987 , \57988 , \57989 , \57990 , \57991 , \57992 , \57993 , \57994 , \57995 , \57996 ,
         \57997 , \57998 , \57999 , \58000 , \58001 , \58002 , \58003 , \58004 , \58005 , \58006 ,
         \58007 , \58008 , \58009 , \58010 , \58011 , \58012 , \58013 , \58014 , \58015 , \58016 ,
         \58017 , \58018 , \58019 , \58020 , \58021 , \58022 , \58023 , \58024 , \58025 , \58026 ,
         \58027 , \58028 , \58029 , \58030 , \58031 , \58032 , \58033 , \58034 , \58035 , \58036 ,
         \58037 , \58038 , \58039 , \58040 , \58041 , \58042 , \58043 , \58044 , \58045 , \58046 ,
         \58047 , \58048 , \58049 , \58050 , \58051 , \58052 , \58053 , \58054 , \58055 , \58056 ,
         \58057 , \58058 , \58059 , \58060 , \58061 , \58062 , \58063 , \58064 , \58065 , \58066 ,
         \58067 , \58068 , \58069 , \58070 , \58071 , \58072 , \58073 , \58074 , \58075 , \58076 ,
         \58077 , \58078 , \58079 , \58080 , \58081 , \58082 , \58083 , \58084 , \58085 , \58086 ,
         \58087 , \58088 , \58089 , \58090 , \58091 , \58092 , \58093 , \58094 , \58095 , \58096 ,
         \58097 , \58098 , \58099 , \58100 , \58101 , \58102 , \58103 , \58104 , \58105 , \58106 ,
         \58107 , \58108 , \58109 , \58110 , \58111 , \58112 , \58113 , \58114 , \58115 , \58116 ,
         \58117 , \58118 , \58119 , \58120 , \58121 , \58122 , \58123 , \58124 , \58125 , \58126 ,
         \58127 , \58128 , \58129 , \58130 , \58131 , \58132 , \58133 , \58134 , \58135 , \58136 ,
         \58137 , \58138 , \58139 , \58140 , \58141 , \58142 , \58143 , \58144 , \58145 , \58146 ,
         \58147 , \58148 , \58149 , \58150 , \58151 , \58152 , \58153 , \58154 , \58155 , \58156 ,
         \58157 , \58158 , \58159 , \58160 , \58161 , \58162 , \58163 , \58164 , \58165 , \58166 ,
         \58167 , \58168 , \58169 , \58170 , \58171 , \58172 , \58173 , \58174 , \58175 , \58176 ,
         \58177 , \58178 , \58179 , \58180 , \58181 , \58182 , \58183 , \58184 , \58185 , \58186 ,
         \58187 , \58188 , \58189 , \58190 , \58191 , \58192 , \58193 , \58194 , \58195 , \58196 ,
         \58197 , \58198 , \58199 , \58200 , \58201 , \58202 , \58203 , \58204 , \58205 , \58206 ,
         \58207 , \58208 , \58209 , \58210 , \58211 , \58212 , \58213 , \58214 , \58215 , \58216 ,
         \58217 , \58218 , \58219 , \58220 , \58221 , \58222 , \58223 , \58224 , \58225 , \58226 ,
         \58227 , \58228 , \58229 , \58230 , \58231 , \58232 , \58233 , \58234 , \58235 , \58236 ,
         \58237 , \58238 , \58239 , \58240 , \58241 , \58242 , \58243 , \58244 , \58245 , \58246 ,
         \58247 , \58248 , \58249 , \58250 , \58251 , \58252 , \58253 , \58254 , \58255 , \58256 ,
         \58257 , \58258 , \58259 , \58260 , \58261 , \58262 , \58263 , \58264 , \58265 , \58266 ,
         \58267 , \58268 , \58269 , \58270 , \58271 , \58272 , \58273 , \58274 , \58275 , \58276 ,
         \58277 , \58278 , \58279 , \58280 , \58281 , \58282 , \58283 , \58284 , \58285 , \58286 ,
         \58287 , \58288 , \58289 , \58290 , \58291 , \58292 , \58293 , \58294 , \58295 , \58296 ,
         \58297 , \58298 , \58299 , \58300 , \58301 , \58302 , \58303 , \58304 , \58305 , \58306 ,
         \58307 , \58308 , \58309 , \58310 , \58311 , \58312 , \58313 , \58314 , \58315 , \58316 ,
         \58317 , \58318 , \58319 , \58320 , \58321 , \58322 , \58323 , \58324 , \58325 , \58326 ,
         \58327 , \58328 , \58329 , \58330 , \58331 , \58332 , \58333 , \58334 , \58335 , \58336 ,
         \58337 , \58338 , \58339 , \58340 , \58341 , \58342 , \58343 , \58344 , \58345 , \58346 ,
         \58347 , \58348 , \58349 , \58350 , \58351 , \58352 , \58353 , \58354 , \58355 , \58356 ,
         \58357 , \58358 , \58359 , \58360 , \58361 , \58362 , \58363 , \58364 , \58365 , \58366 ,
         \58367 , \58368 , \58369 , \58370 , \58371 , \58372 , \58373 , \58374 , \58375 , \58376 ,
         \58377 , \58378 , \58379 , \58380 , \58381 , \58382 , \58383 , \58384 , \58385 , \58386 ,
         \58387 , \58388 , \58389 , \58390 , \58391 , \58392 , \58393 , \58394 , \58395 , \58396 ,
         \58397 , \58398 , \58399 , \58400 , \58401 , \58402 , \58403 , \58404 , \58405 , \58406 ,
         \58407 , \58408 , \58409 , \58410 , \58411 , \58412 , \58413 , \58414 , \58415 , \58416 ,
         \58417 , \58418 , \58419 , \58420 , \58421 , \58422 , \58423 , \58424 , \58425 , \58426 ,
         \58427 , \58428 , \58429 , \58430 , \58431 , \58432 , \58433 , \58434 , \58435 , \58436 ,
         \58437 , \58438 , \58439 , \58440 , \58441 , \58442 , \58443 , \58444 , \58445 , \58446 ,
         \58447 , \58448 , \58449 , \58450 , \58451 , \58452 , \58453 , \58454 , \58455 , \58456 ,
         \58457 , \58458 , \58459 , \58460 , \58461 , \58462 , \58463 , \58464 , \58465 , \58466 ,
         \58467 , \58468 , \58469 , \58470 , \58471 , \58472 , \58473 , \58474 , \58475 , \58476 ,
         \58477 , \58478 , \58479 , \58480 , \58481 , \58482 , \58483 , \58484 , \58485 , \58486 ,
         \58487 , \58488 , \58489 , \58490 , \58491 , \58492 , \58493 , \58494 , \58495 , \58496 ,
         \58497 , \58498 , \58499 , \58500 , \58501 , \58502 , \58503 , \58504 , \58505 , \58506 ,
         \58507 , \58508 , \58509 , \58510 , \58511 , \58512 , \58513 , \58514 , \58515 , \58516 ,
         \58517 , \58518 , \58519 , \58520 , \58521 , \58522 , \58523 , \58524 , \58525 , \58526 ,
         \58527 , \58528 , \58529 , \58530 , \58531 , \58532 , \58533 , \58534 , \58535 , \58536 ,
         \58537 , \58538 , \58539 , \58540 , \58541 , \58542 , \58543 , \58544 , \58545 , \58546 ,
         \58547 , \58548 , \58549 , \58550 , \58551 , \58552 , \58553 , \58554 , \58555 , \58556 ,
         \58557 , \58558 , \58559 , \58560 , \58561 , \58562 , \58563 , \58564 , \58565 , \58566 ,
         \58567 , \58568 , \58569 , \58570 , \58571 , \58572 , \58573 , \58574 , \58575 , \58576 ,
         \58577 , \58578 , \58579 , \58580 , \58581 , \58582 , \58583 , \58584 , \58585 , \58586 ,
         \58587 , \58588 , \58589 , \58590 , \58591 , \58592 , \58593 , \58594 , \58595 , \58596 ,
         \58597 , \58598 , \58599 , \58600 , \58601 , \58602 , \58603 , \58604 , \58605 , \58606 ,
         \58607 , \58608 , \58609 , \58610 , \58611 , \58612 , \58613 , \58614 , \58615 , \58616 ,
         \58617 , \58618 , \58619 , \58620 , \58621 , \58622 , \58623 , \58624 , \58625 , \58626 ,
         \58627 , \58628 , \58629 , \58630 , \58631 , \58632 , \58633 , \58634 , \58635 , \58636 ,
         \58637 , \58638 , \58639 , \58640 , \58641 , \58642 , \58643 , \58644 , \58645 , \58646 ,
         \58647 , \58648 , \58649 , \58650 , \58651 , \58652 , \58653 , \58654 , \58655 , \58656 ,
         \58657 , \58658 , \58659 , \58660 , \58661 , \58662 , \58663 , \58664 , \58665 , \58666 ,
         \58667 , \58668 , \58669 , \58670 , \58671 , \58672 , \58673 , \58674 , \58675 , \58676 ,
         \58677 , \58678 , \58679 , \58680 , \58681 , \58682 , \58683 , \58684 , \58685 , \58686 ,
         \58687 , \58688 , \58689 , \58690 , \58691 , \58692 , \58693 , \58694 , \58695 , \58696 ,
         \58697 , \58698 , \58699 , \58700 , \58701 , \58702 , \58703 , \58704 , \58705 , \58706 ,
         \58707 , \58708 , \58709 , \58710 , \58711 , \58712 , \58713 , \58714 , \58715 , \58716 ,
         \58717 , \58718 , \58719 , \58720 , \58721 , \58722 , \58723 , \58724 , \58725 , \58726 ,
         \58727 , \58728 , \58729 , \58730 , \58731 , \58732 , \58733 , \58734 , \58735 , \58736 ,
         \58737 , \58738 , \58739 , \58740 , \58741 , \58742 , \58743 , \58744 , \58745 , \58746 ,
         \58747 , \58748 , \58749 , \58750 , \58751 , \58752 , \58753 , \58754 , \58755 , \58756 ,
         \58757 , \58758 , \58759 , \58760 , \58761 , \58762 , \58763 , \58764 , \58765 , \58766 ,
         \58767 , \58768 , \58769 , \58770 , \58771 , \58772 , \58773 , \58774 , \58775 , \58776 ,
         \58777 , \58778 , \58779 , \58780 , \58781 , \58782 , \58783 , \58784 , \58785 , \58786 ,
         \58787 , \58788 , \58789 , \58790 , \58791 , \58792 , \58793 , \58794 , \58795 , \58796 ,
         \58797 , \58798 , \58799 , \58800 , \58801 , \58802 , \58803 , \58804 , \58805 , \58806 ,
         \58807 , \58808 , \58809 , \58810 , \58811 , \58812 , \58813 , \58814 , \58815 , \58816 ,
         \58817 , \58818 , \58819 , \58820 , \58821 , \58822 , \58823 , \58824 , \58825 , \58826 ,
         \58827 , \58828 , \58829 , \58830 , \58831 , \58832 , \58833 , \58834 , \58835 , \58836 ,
         \58837 , \58838 , \58839 , \58840 , \58841 , \58842 , \58843 , \58844 , \58845 , \58846 ,
         \58847 , \58848 , \58849 , \58850 , \58851 , \58852 , \58853 , \58854 , \58855 , \58856 ,
         \58857 , \58858 , \58859 , \58860 , \58861 , \58862 , \58863 , \58864 , \58865 , \58866 ,
         \58867 , \58868 , \58869 , \58870 , \58871 , \58872 , \58873 , \58874 , \58875 , \58876 ,
         \58877 , \58878 , \58879 , \58880 , \58881 , \58882 , \58883 , \58884 , \58885 , \58886 ,
         \58887 , \58888 , \58889 , \58890 , \58891 , \58892 , \58893 , \58894 , \58895 , \58896 ,
         \58897 , \58898 , \58899 , \58900 , \58901 , \58902 , \58903 , \58904 , \58905 , \58906 ,
         \58907 , \58908 , \58909 , \58910 , \58911 , \58912 , \58913 , \58914 , \58915 , \58916 ,
         \58917 , \58918 , \58919 , \58920 , \58921 , \58922 , \58923 , \58924 , \58925 , \58926 ,
         \58927 , \58928 , \58929 , \58930 , \58931 , \58932 , \58933 , \58934 , \58935 , \58936 ,
         \58937 , \58938 , \58939 , \58940 , \58941 , \58942 , \58943 , \58944 , \58945 , \58946 ,
         \58947 , \58948 , \58949 , \58950 , \58951 , \58952 , \58953 , \58954 , \58955 , \58956 ,
         \58957 , \58958 , \58959 , \58960 , \58961 , \58962 , \58963 , \58964 , \58965 , \58966 ,
         \58967 , \58968 , \58969 , \58970 , \58971 , \58972 , \58973 , \58974 , \58975 , \58976 ,
         \58977 , \58978 , \58979 , \58980 , \58981 , \58982 , \58983 , \58984 , \58985 , \58986 ,
         \58987 , \58988 , \58989 , \58990 , \58991 , \58992 , \58993 , \58994 , \58995 , \58996 ,
         \58997 , \58998 , \58999 , \59000 , \59001 , \59002 , \59003 , \59004 , \59005 , \59006 ,
         \59007 , \59008 , \59009 , \59010 , \59011 , \59012 , \59013 , \59014 , \59015 , \59016 ,
         \59017 , \59018 , \59019 , \59020 , \59021 , \59022 , \59023 , \59024 , \59025 , \59026 ,
         \59027 , \59028 , \59029 , \59030 , \59031 , \59032 , \59033 , \59034 , \59035 , \59036 ,
         \59037 , \59038 , \59039 , \59040 , \59041 , \59042 , \59043 , \59044 , \59045 , \59046 ,
         \59047 , \59048 , \59049 , \59050 , \59051 , \59052 , \59053 , \59054 , \59055 , \59056 ,
         \59057 , \59058 , \59059 , \59060 , \59061 , \59062 , \59063 , \59064 , \59065 , \59066 ,
         \59067 , \59068 , \59069 , \59070 , \59071 , \59072 , \59073 , \59074 , \59075 , \59076 ,
         \59077 , \59078 , \59079 , \59080 , \59081 , \59082 , \59083 , \59084 , \59085 , \59086 ,
         \59087 , \59088 , \59089 , \59090 , \59091 , \59092 , \59093 , \59094 , \59095 , \59096 ,
         \59097 , \59098 , \59099 , \59100 , \59101 , \59102 , \59103 , \59104 , \59105 , \59106 ,
         \59107 , \59108 , \59109 , \59110 , \59111 , \59112 , \59113 , \59114 , \59115 , \59116 ,
         \59117 , \59118 , \59119 , \59120 , \59121 , \59122 , \59123 , \59124 , \59125 , \59126 ,
         \59127 , \59128 , \59129 , \59130 , \59131 , \59132 , \59133 , \59134 , \59135 , \59136 ,
         \59137 , \59138 , \59139 , \59140 , \59141 , \59142 , \59143 , \59144 , \59145 , \59146 ,
         \59147 , \59148 , \59149 , \59150 , \59151 , \59152 , \59153 , \59154 , \59155 , \59156 ,
         \59157 , \59158 , \59159 , \59160 , \59161 , \59162 , \59163 , \59164 , \59165 , \59166 ,
         \59167 , \59168 , \59169 , \59170 , \59171 , \59172 , \59173 , \59174 , \59175 , \59176 ,
         \59177 , \59178 , \59179 , \59180 , \59181 , \59182 , \59183 , \59184 , \59185 , \59186 ,
         \59187 , \59188 , \59189 , \59190 , \59191 , \59192 , \59193 , \59194 , \59195 , \59196 ,
         \59197 , \59198 , \59199 , \59200 , \59201 , \59202 , \59203 , \59204 , \59205 , \59206 ,
         \59207 , \59208 , \59209 , \59210 , \59211 , \59212 , \59213 , \59214 , \59215 , \59216 ,
         \59217 , \59218 , \59219 , \59220 , \59221 , \59222 , \59223 , \59224 , \59225 , \59226 ,
         \59227 , \59228 , \59229 , \59230 , \59231 , \59232 , \59233 , \59234 , \59235 , \59236 ,
         \59237 , \59238 , \59239 , \59240 , \59241 , \59242 , \59243 , \59244 , \59245 , \59246 ,
         \59247 , \59248 , \59249 , \59250 , \59251 , \59252 , \59253 , \59254 , \59255 , \59256 ,
         \59257 , \59258 , \59259 , \59260 , \59261 , \59262 , \59263 , \59264 , \59265 , \59266 ,
         \59267 , \59268 , \59269 , \59270 , \59271 , \59272 , \59273 , \59274 , \59275 , \59276 ,
         \59277 , \59278 , \59279 , \59280 , \59281 , \59282 , \59283 , \59284 , \59285 , \59286 ,
         \59287 , \59288 , \59289 , \59290 , \59291 , \59292 , \59293 , \59294 , \59295 , \59296 ,
         \59297 , \59298 , \59299 , \59300 , \59301 , \59302 , \59303 , \59304 , \59305 , \59306 ,
         \59307 , \59308 , \59309 , \59310 , \59311 , \59312 , \59313 , \59314 , \59315 , \59316 ,
         \59317 , \59318 , \59319 , \59320 , \59321 , \59322 , \59323 , \59324 , \59325 , \59326 ,
         \59327 , \59328 , \59329 , \59330 , \59331 , \59332 , \59333 , \59334 , \59335 , \59336 ,
         \59337 , \59338 , \59339 , \59340 , \59341 , \59342 , \59343 , \59344 , \59345 , \59346 ,
         \59347 , \59348 , \59349 , \59350 , \59351 , \59352 , \59353 , \59354 , \59355 , \59356 ,
         \59357 , \59358 , \59359 , \59360 , \59361 , \59362 , \59363 , \59364 , \59365 , \59366 ,
         \59367 , \59368 , \59369 , \59370 , \59371 , \59372 , \59373 , \59374 , \59375 , \59376 ,
         \59377 , \59378 , \59379 , \59380 , \59381 , \59382 , \59383 , \59384 , \59385 , \59386 ,
         \59387 , \59388 , \59389 , \59390 , \59391 , \59392 , \59393 , \59394 , \59395 , \59396 ,
         \59397 , \59398 , \59399 , \59400 , \59401 , \59402 , \59403 , \59404 , \59405 , \59406 ,
         \59407 , \59408 , \59409 , \59410 , \59411 , \59412 , \59413 , \59414 , \59415 , \59416 ,
         \59417 , \59418 , \59419 , \59420 , \59421 , \59422 , \59423 , \59424 , \59425 , \59426 ,
         \59427 , \59428 , \59429 , \59430 , \59431 , \59432 , \59433 , \59434 , \59435 , \59436 ,
         \59437 , \59438 , \59439 , \59440 , \59441 , \59442 , \59443 , \59444 , \59445 , \59446 ,
         \59447 , \59448 , \59449 , \59450 , \59451 , \59452 , \59453 , \59454 , \59455 , \59456 ,
         \59457 , \59458 , \59459 , \59460 , \59461 , \59462 , \59463 , \59464 , \59465 , \59466 ,
         \59467 , \59468 , \59469 , \59470 , \59471 , \59472 , \59473 , \59474 , \59475 , \59476 ,
         \59477 , \59478 , \59479 , \59480 , \59481 , \59482 , \59483 , \59484 , \59485 , \59486 ,
         \59487 , \59488 , \59489 , \59490 , \59491 , \59492 , \59493 , \59494 , \59495 , \59496 ,
         \59497 , \59498 , \59499 , \59500 , \59501 , \59502 , \59503 , \59504 , \59505 , \59506 ,
         \59507 , \59508 , \59509 , \59510 , \59511 , \59512 , \59513 , \59514 , \59515 , \59516 ,
         \59517 , \59518 , \59519 , \59520 , \59521 , \59522 , \59523 , \59524 , \59525 , \59526 ,
         \59527 , \59528 , \59529 , \59530 , \59531 , \59532 , \59533 , \59534 , \59535 , \59536 ,
         \59537 , \59538 , \59539 , \59540 , \59541 , \59542 , \59543 , \59544 , \59545 , \59546 ,
         \59547 , \59548 , \59549 , \59550 , \59551 , \59552 , \59553 , \59554 , \59555 , \59556 ,
         \59557 , \59558 , \59559 , \59560 , \59561 , \59562 , \59563 , \59564 , \59565 , \59566 ,
         \59567 , \59568 , \59569 , \59570 , \59571 , \59572 , \59573 , \59574 , \59575 , \59576 ,
         \59577 , \59578 , \59579 , \59580 , \59581 , \59582 , \59583 , \59584 , \59585 , \59586 ,
         \59587 , \59588 , \59589 , \59590 , \59591 , \59592 , \59593 , \59594 , \59595 , \59596 ,
         \59597 , \59598 , \59599 , \59600 , \59601 , \59602 , \59603 , \59604 , \59605 , \59606 ,
         \59607 , \59608 , \59609 , \59610 , \59611 , \59612 , \59613 , \59614 , \59615 , \59616 ,
         \59617 , \59618 , \59619 , \59620 , \59621 , \59622 , \59623 , \59624 , \59625 , \59626 ,
         \59627 , \59628 , \59629 , \59630 , \59631 , \59632 , \59633 , \59634 , \59635 , \59636 ,
         \59637 , \59638 , \59639 , \59640 , \59641 , \59642 , \59643 , \59644 , \59645 , \59646 ,
         \59647 , \59648 , \59649 , \59650 , \59651 , \59652 , \59653 , \59654 , \59655 , \59656 ,
         \59657 , \59658 , \59659 , \59660 , \59661 , \59662 , \59663 , \59664 , \59665 , \59666 ,
         \59667 , \59668 , \59669 , \59670 , \59671 , \59672 , \59673 , \59674 , \59675 , \59676 ,
         \59677 , \59678 , \59679 , \59680 , \59681 , \59682 , \59683 , \59684 , \59685 , \59686 ,
         \59687 , \59688 , \59689 , \59690 , \59691 , \59692 , \59693 , \59694 , \59695 , \59696 ,
         \59697 , \59698 , \59699 , \59700 , \59701 , \59702 , \59703 , \59704 , \59705 , \59706 ,
         \59707 , \59708 , \59709 , \59710 , \59711 , \59712 , \59713 , \59714 , \59715 , \59716 ,
         \59717 , \59718 , \59719 , \59720 , \59721 , \59722 , \59723 , \59724 , \59725 , \59726 ,
         \59727 , \59728 , \59729 , \59730 , \59731 , \59732 , \59733 , \59734 , \59735 , \59736 ,
         \59737 , \59738 , \59739 , \59740 , \59741 , \59742 , \59743 , \59744 , \59745 , \59746 ,
         \59747 , \59748 , \59749 , \59750 , \59751 , \59752 , \59753 , \59754 , \59755 , \59756 ,
         \59757 , \59758 , \59759 , \59760 , \59761 , \59762 , \59763 , \59764 , \59765 , \59766 ,
         \59767 , \59768 , \59769 , \59770 , \59771 , \59772 , \59773 , \59774 , \59775 , \59776 ,
         \59777 , \59778 , \59779 , \59780 , \59781 , \59782 , \59783 , \59784 , \59785 , \59786 ,
         \59787 , \59788 , \59789 , \59790 , \59791 , \59792 , \59793 , \59794 , \59795 , \59796 ,
         \59797 , \59798 , \59799 , \59800 , \59801 , \59802 , \59803 , \59804 , \59805 , \59806 ,
         \59807 , \59808 , \59809 , \59810 , \59811 , \59812 , \59813 , \59814 , \59815 , \59816 ,
         \59817 , \59818 , \59819 , \59820 , \59821 , \59822 , \59823 , \59824 , \59825 , \59826 ,
         \59827 , \59828 , \59829 , \59830 , \59831 , \59832 , \59833 , \59834 , \59835 , \59836 ,
         \59837 , \59838 , \59839 , \59840 , \59841 , \59842 , \59843 , \59844 , \59845 , \59846 ,
         \59847 , \59848 , \59849 , \59850 , \59851 , \59852 , \59853 , \59854 , \59855 , \59856 ,
         \59857 , \59858 , \59859 , \59860 , \59861 , \59862 , \59863 , \59864 , \59865 , \59866 ,
         \59867 , \59868 , \59869 , \59870 , \59871 , \59872 , \59873 , \59874 , \59875 , \59876 ,
         \59877 , \59878 , \59879 , \59880 , \59881 , \59882 , \59883 , \59884 , \59885 , \59886 ,
         \59887 , \59888 , \59889 , \59890 , \59891 , \59892 , \59893 , \59894 , \59895 , \59896 ,
         \59897 , \59898 , \59899 , \59900 , \59901 , \59902 , \59903 , \59904 , \59905 , \59906 ,
         \59907 , \59908 , \59909 , \59910 , \59911 , \59912 , \59913 , \59914 , \59915 , \59916 ,
         \59917 , \59918 , \59919 , \59920 , \59921 , \59922 , \59923 , \59924 , \59925 , \59926 ,
         \59927 , \59928 , \59929 , \59930 , \59931 , \59932 , \59933 , \59934 , \59935 , \59936 ,
         \59937 , \59938 , \59939 , \59940 , \59941 , \59942 , \59943 , \59944 , \59945 , \59946 ,
         \59947 , \59948 , \59949 , \59950 , \59951 , \59952 , \59953 , \59954 , \59955 , \59956 ,
         \59957 , \59958 , \59959 , \59960 , \59961 , \59962 , \59963 , \59964 , \59965 , \59966 ,
         \59967 , \59968 , \59969 , \59970 , \59971 , \59972 , \59973 , \59974 , \59975 , \59976 ,
         \59977 , \59978 , \59979 , \59980 , \59981 , \59982 , \59983 , \59984 , \59985 , \59986 ,
         \59987 , \59988 , \59989 , \59990 , \59991 , \59992 , \59993 , \59994 , \59995 , \59996 ,
         \59997 , \59998 , \59999 , \60000 , \60001 , \60002 , \60003 , \60004 , \60005 , \60006 ,
         \60007 , \60008 , \60009 , \60010 , \60011 , \60012 , \60013 , \60014 , \60015 , \60016 ,
         \60017 , \60018 , \60019 , \60020 , \60021 , \60022 , \60023 , \60024 , \60025 , \60026 ,
         \60027 , \60028 , \60029 , \60030 , \60031 , \60032 , \60033 , \60034 , \60035 , \60036 ,
         \60037 , \60038 , \60039 , \60040 , \60041 , \60042 , \60043 , \60044 , \60045 , \60046 ,
         \60047 , \60048 , \60049 , \60050 , \60051 , \60052 , \60053 , \60054 , \60055 , \60056 ,
         \60057 , \60058 , \60059 , \60060 , \60061 , \60062 , \60063 , \60064 , \60065 , \60066 ,
         \60067 , \60068 , \60069 , \60070 , \60071 , \60072 , \60073 , \60074 , \60075 , \60076 ,
         \60077 , \60078 , \60079 , \60080 , \60081 , \60082 , \60083 , \60084 , \60085 , \60086 ,
         \60087 , \60088 , \60089 , \60090 , \60091 , \60092 , \60093 , \60094 , \60095 , \60096 ,
         \60097 , \60098 , \60099 , \60100 , \60101 , \60102 , \60103 , \60104 , \60105 , \60106 ,
         \60107 , \60108 , \60109 , \60110 , \60111 , \60112 , \60113 , \60114 , \60115 , \60116 ,
         \60117 , \60118 , \60119 , \60120 , \60121 , \60122 , \60123 , \60124 , \60125 , \60126 ,
         \60127 , \60128 , \60129 , \60130 , \60131 , \60132 , \60133 , \60134 , \60135 , \60136 ,
         \60137 , \60138 , \60139 , \60140 , \60141 , \60142 , \60143 , \60144 , \60145 , \60146 ,
         \60147 , \60148 , \60149 , \60150 , \60151 , \60152 , \60153 , \60154 , \60155 , \60156 ,
         \60157 , \60158 , \60159 , \60160 , \60161 , \60162 , \60163 , \60164 , \60165 , \60166 ,
         \60167 , \60168 , \60169 , \60170 , \60171 , \60172 , \60173 , \60174 , \60175 , \60176 ,
         \60177 , \60178 , \60179 , \60180 , \60181 , \60182 , \60183 , \60184 , \60185 , \60186 ,
         \60187 , \60188 , \60189 , \60190 , \60191 , \60192 , \60193 , \60194 , \60195 , \60196 ,
         \60197 , \60198 , \60199 , \60200 , \60201 , \60202 , \60203 , \60204 , \60205 , \60206 ,
         \60207 , \60208 , \60209 , \60210 , \60211 , \60212 , \60213 , \60214 , \60215 , \60216 ,
         \60217 , \60218 , \60219 , \60220 , \60221 , \60222 , \60223 , \60224 , \60225 , \60226 ,
         \60227 , \60228 , \60229 , \60230 , \60231 , \60232 , \60233 , \60234 , \60235 , \60236 ,
         \60237 , \60238 , \60239 , \60240 , \60241 , \60242 , \60243 , \60244 , \60245 , \60246 ,
         \60247 , \60248 , \60249 , \60250 , \60251 , \60252 , \60253 , \60254 , \60255 , \60256 ,
         \60257 , \60258 , \60259 , \60260 , \60261 , \60262 , \60263 , \60264 , \60265 , \60266 ,
         \60267 , \60268 , \60269 , \60270 , \60271 , \60272 , \60273 , \60274 , \60275 , \60276 ,
         \60277 , \60278 , \60279 , \60280 , \60281 , \60282 , \60283 , \60284 , \60285 , \60286 ,
         \60287 , \60288 , \60289 , \60290 , \60291 , \60292 , \60293 , \60294 , \60295 , \60296 ,
         \60297 , \60298 , \60299 , \60300 , \60301 , \60302 , \60303 , \60304 , \60305 , \60306 ,
         \60307 , \60308 , \60309 , \60310 , \60311 , \60312 , \60313 , \60314 , \60315 , \60316 ,
         \60317 , \60318 , \60319 , \60320 , \60321 , \60322 , \60323 , \60324 , \60325 , \60326 ,
         \60327 , \60328 , \60329 , \60330 , \60331 , \60332 , \60333 , \60334 , \60335 , \60336 ,
         \60337 , \60338 , \60339 , \60340 , \60341 , \60342 , \60343 , \60344 , \60345 , \60346 ,
         \60347 , \60348 , \60349 , \60350 , \60351 , \60352 , \60353 , \60354 , \60355 , \60356 ,
         \60357 , \60358 , \60359 , \60360 , \60361 , \60362 , \60363 , \60364 , \60365 , \60366 ,
         \60367 , \60368 , \60369 , \60370 , \60371 , \60372 , \60373 , \60374 , \60375 , \60376 ,
         \60377 , \60378 , \60379 , \60380 , \60381 , \60382 , \60383 , \60384 , \60385 , \60386 ,
         \60387 , \60388 , \60389 , \60390 , \60391 , \60392 , \60393 , \60394 , \60395 , \60396 ,
         \60397 , \60398 , \60399 , \60400 , \60401 , \60402 , \60403 , \60404 , \60405 , \60406 ,
         \60407 , \60408 , \60409 , \60410 , \60411 , \60412 , \60413 , \60414 , \60415 , \60416 ,
         \60417 , \60418 , \60419 , \60420 , \60421 , \60422 , \60423 , \60424 , \60425 , \60426 ,
         \60427 , \60428 , \60429 , \60430 , \60431 , \60432 , \60433 , \60434 , \60435 , \60436 ,
         \60437 , \60438 , \60439 , \60440 , \60441 , \60442 , \60443 , \60444 , \60445 , \60446 ,
         \60447 , \60448 , \60449 , \60450 , \60451 , \60452 , \60453 , \60454 , \60455 , \60456 ,
         \60457 , \60458 , \60459 , \60460 , \60461 , \60462 , \60463 , \60464 , \60465 , \60466 ,
         \60467 , \60468 , \60469 , \60470 , \60471 , \60472 , \60473 , \60474 , \60475 , \60476 ,
         \60477 , \60478 , \60479 , \60480 , \60481 , \60482 , \60483 , \60484 , \60485 , \60486 ,
         \60487 , \60488 , \60489 , \60490 , \60491 , \60492 , \60493 , \60494 , \60495 , \60496 ,
         \60497 , \60498 , \60499 , \60500 , \60501 , \60502 , \60503 , \60504 , \60505 , \60506 ,
         \60507 , \60508 , \60509 , \60510 , \60511 , \60512 , \60513 , \60514 , \60515 , \60516 ,
         \60517 , \60518 , \60519 , \60520 , \60521 , \60522 , \60523 , \60524 , \60525 , \60526 ,
         \60527 , \60528 , \60529 , \60530 , \60531 , \60532 , \60533 , \60534 , \60535 , \60536 ,
         \60537 , \60538 , \60539 , \60540 , \60541 , \60542 , \60543 , \60544 , \60545 , \60546 ,
         \60547 , \60548 , \60549 , \60550 , \60551 , \60552 , \60553 , \60554 , \60555 , \60556 ,
         \60557 , \60558 , \60559 , \60560 , \60561 , \60562 , \60563 , \60564 , \60565 , \60566 ,
         \60567 , \60568 , \60569 , \60570 , \60571 , \60572 , \60573 , \60574 , \60575 , \60576 ,
         \60577 , \60578 , \60579 , \60580 , \60581 , \60582 , \60583 , \60584 , \60585 , \60586 ,
         \60587 , \60588 , \60589 , \60590 , \60591 , \60592 , \60593 , \60594 , \60595 , \60596 ,
         \60597 , \60598 , \60599 , \60600 , \60601 , \60602 , \60603 , \60604 , \60605 , \60606 ,
         \60607 , \60608 , \60609 , \60610 , \60611 , \60612 , \60613 , \60614 , \60615 , \60616 ,
         \60617 , \60618 , \60619 , \60620 , \60621 , \60622 , \60623 , \60624 , \60625 , \60626 ,
         \60627 , \60628 , \60629 , \60630 , \60631 , \60632 , \60633 , \60634 , \60635 , \60636 ,
         \60637 , \60638 , \60639 , \60640 , \60641 , \60642 , \60643 , \60644 , \60645 , \60646 ,
         \60647 , \60648 , \60649 , \60650 , \60651 , \60652 , \60653 , \60654 , \60655 , \60656 ,
         \60657 , \60658 , \60659 , \60660 , \60661 , \60662 , \60663 , \60664 , \60665 , \60666 ,
         \60667 , \60668 , \60669 , \60670 , \60671 , \60672 , \60673 , \60674 , \60675 , \60676 ,
         \60677 , \60678 , \60679 , \60680 , \60681 , \60682 , \60683 , \60684 , \60685 , \60686 ,
         \60687 , \60688 , \60689 , \60690 , \60691 , \60692 , \60693 , \60694 , \60695 , \60696 ,
         \60697 , \60698 , \60699 , \60700 , \60701 , \60702 , \60703 , \60704 , \60705 , \60706 ,
         \60707 , \60708 , \60709 , \60710 , \60711 , \60712 , \60713 , \60714 , \60715 , \60716 ,
         \60717 , \60718 , \60719 , \60720 , \60721 , \60722 , \60723 , \60724 , \60725 , \60726 ,
         \60727 , \60728 , \60729 , \60730 , \60731 , \60732 , \60733 , \60734 , \60735 , \60736 ,
         \60737 , \60738 , \60739 , \60740 , \60741 , \60742 , \60743 , \60744 , \60745 , \60746 ,
         \60747 , \60748 , \60749 , \60750 , \60751 , \60752 , \60753 , \60754 , \60755 , \60756 ,
         \60757 , \60758 , \60759 , \60760 , \60761 , \60762 , \60763 , \60764 , \60765 , \60766 ,
         \60767 , \60768 , \60769 , \60770 , \60771 , \60772 , \60773 , \60774 , \60775 , \60776 ,
         \60777 , \60778 , \60779 , \60780 , \60781 , \60782 , \60783 , \60784 , \60785 , \60786 ,
         \60787 , \60788 , \60789 , \60790 , \60791 , \60792 , \60793 , \60794 , \60795 , \60796 ,
         \60797 , \60798 , \60799 , \60800 , \60801 , \60802 , \60803 , \60804 , \60805 , \60806 ,
         \60807 , \60808 , \60809 , \60810 , \60811 , \60812 , \60813 , \60814 , \60815 , \60816 ,
         \60817 , \60818 , \60819 , \60820 , \60821 , \60822 , \60823 , \60824 , \60825 , \60826 ,
         \60827 , \60828 , \60829 , \60830 , \60831 , \60832 , \60833 , \60834 , \60835 , \60836 ,
         \60837 , \60838 , \60839 , \60840 , \60841 , \60842 , \60843 , \60844 , \60845 , \60846 ,
         \60847 , \60848 , \60849 , \60850 , \60851 , \60852 , \60853 , \60854 , \60855 , \60856 ,
         \60857 , \60858 , \60859 , \60860 , \60861 , \60862 , \60863 , \60864 , \60865 , \60866 ,
         \60867 , \60868 , \60869 , \60870 , \60871 , \60872 , \60873 , \60874 , \60875 , \60876 ,
         \60877 , \60878 , \60879 , \60880 , \60881 , \60882 , \60883 , \60884 , \60885 , \60886 ,
         \60887 , \60888 , \60889 , \60890 , \60891 , \60892 , \60893 , \60894 , \60895 , \60896 ,
         \60897 , \60898 , \60899 , \60900 , \60901 , \60902 , \60903 , \60904 , \60905 , \60906 ,
         \60907 , \60908 , \60909 , \60910 , \60911 , \60912 , \60913 , \60914 , \60915 , \60916 ,
         \60917 , \60918 , \60919 , \60920 , \60921 , \60922 , \60923 , \60924 , \60925 , \60926 ,
         \60927 , \60928 , \60929 , \60930 , \60931 , \60932 , \60933 , \60934 , \60935 , \60936 ,
         \60937 , \60938 , \60939 , \60940 , \60941 , \60942 , \60943 , \60944 , \60945 , \60946 ,
         \60947 , \60948 , \60949 , \60950 , \60951 , \60952 , \60953 , \60954 , \60955 , \60956 ,
         \60957 , \60958 , \60959 , \60960 , \60961 , \60962 , \60963 , \60964 , \60965 , \60966 ,
         \60967 , \60968 , \60969 , \60970 , \60971 , \60972 , \60973 , \60974 , \60975 , \60976 ,
         \60977 , \60978 , \60979 , \60980 , \60981 , \60982 , \60983 , \60984 , \60985 , \60986 ,
         \60987 , \60988 , \60989 , \60990 , \60991 , \60992 , \60993 , \60994 , \60995 , \60996 ,
         \60997 , \60998 , \60999 , \61000 , \61001 , \61002 , \61003 , \61004 , \61005 , \61006 ,
         \61007 , \61008 , \61009 , \61010 , \61011 , \61012 , \61013 , \61014 , \61015 , \61016 ,
         \61017 , \61018 , \61019 , \61020 , \61021 , \61022 , \61023 , \61024 , \61025 , \61026 ,
         \61027 , \61028 , \61029 , \61030 , \61031 , \61032 , \61033 , \61034 , \61035 , \61036 ,
         \61037 , \61038 , \61039 , \61040 , \61041 , \61042 , \61043 , \61044 , \61045 , \61046 ,
         \61047 , \61048 , \61049 , \61050 , \61051 , \61052 , \61053 , \61054 , \61055 , \61056 ,
         \61057 , \61058 , \61059 , \61060 , \61061 , \61062 , \61063 , \61064 , \61065 , \61066 ,
         \61067 , \61068 , \61069 , \61070 , \61071 , \61072 , \61073 , \61074 , \61075 , \61076 ,
         \61077 , \61078 , \61079 , \61080 , \61081 , \61082 , \61083 , \61084 , \61085 , \61086 ,
         \61087 , \61088 , \61089 , \61090 , \61091 , \61092 , \61093 , \61094 , \61095 , \61096 ,
         \61097 , \61098 , \61099 , \61100 , \61101 , \61102 , \61103 , \61104 , \61105 , \61106 ,
         \61107 , \61108 , \61109 , \61110 , \61111 , \61112 , \61113 , \61114 , \61115 , \61116 ,
         \61117 , \61118 , \61119 , \61120 , \61121 , \61122 , \61123 , \61124 , \61125 , \61126 ,
         \61127 , \61128 , \61129 , \61130 , \61131 , \61132 , \61133 , \61134 , \61135 , \61136 ,
         \61137 , \61138 , \61139 , \61140 , \61141 , \61142 , \61143 , \61144 , \61145 , \61146 ,
         \61147 , \61148 , \61149 , \61150 , \61151 , \61152 , \61153 , \61154 , \61155 , \61156 ,
         \61157 , \61158 , \61159 , \61160 , \61161 , \61162 , \61163 , \61164 , \61165 , \61166 ,
         \61167 , \61168 , \61169 , \61170 , \61171 , \61172 , \61173 , \61174 , \61175 , \61176 ,
         \61177 , \61178 , \61179 , \61180 , \61181 , \61182 , \61183 , \61184 , \61185 , \61186 ,
         \61187 , \61188 , \61189 , \61190 , \61191 , \61192 , \61193 , \61194 , \61195 , \61196 ,
         \61197 , \61198 , \61199 , \61200 , \61201 , \61202 , \61203 , \61204 , \61205 , \61206 ,
         \61207 , \61208 , \61209 , \61210 , \61211 , \61212 , \61213 , \61214 , \61215 , \61216 ,
         \61217 , \61218 , \61219 , \61220 , \61221 , \61222 , \61223 , \61224 , \61225 , \61226 ,
         \61227 , \61228 , \61229 , \61230 , \61231 , \61232 , \61233 , \61234 , \61235 , \61236 ,
         \61237 , \61238 , \61239 , \61240 , \61241 , \61242 , \61243 , \61244 , \61245 , \61246 ,
         \61247 , \61248 , \61249 , \61250 , \61251 , \61252 , \61253 , \61254 , \61255 , \61256 ,
         \61257 , \61258 , \61259 , \61260 , \61261 , \61262 , \61263 , \61264 , \61265 , \61266 ,
         \61267 , \61268 , \61269 , \61270 , \61271 , \61272 , \61273 , \61274 , \61275 , \61276 ,
         \61277 , \61278 , \61279 , \61280 , \61281 , \61282 , \61283 , \61284 , \61285 , \61286 ,
         \61287 , \61288 , \61289 , \61290 , \61291 , \61292 , \61293 , \61294 , \61295 , \61296 ,
         \61297 , \61298 , \61299 , \61300 , \61301 , \61302 , \61303 , \61304 , \61305 , \61306 ,
         \61307 , \61308 , \61309 , \61310 , \61311 , \61312 , \61313 , \61314 , \61315 , \61316 ,
         \61317 , \61318 , \61319 , \61320 , \61321 , \61322 , \61323 , \61324 , \61325 , \61326 ,
         \61327 , \61328 , \61329 , \61330 , \61331 , \61332 , \61333 , \61334 , \61335 , \61336 ,
         \61337 , \61338 , \61339 , \61340 , \61341 , \61342 , \61343 , \61344 , \61345 , \61346 ,
         \61347 , \61348 , \61349 , \61350 , \61351 , \61352 , \61353 , \61354 , \61355 , \61356 ,
         \61357 , \61358 , \61359 , \61360 , \61361 , \61362 , \61363 , \61364 , \61365 , \61366 ,
         \61367 , \61368 , \61369 , \61370 , \61371 , \61372 , \61373 , \61374 , \61375 , \61376 ,
         \61377 , \61378 , \61379 , \61380 , \61381 , \61382 , \61383 , \61384 , \61385 , \61386 ,
         \61387 , \61388 , \61389 , \61390 , \61391 , \61392 , \61393 , \61394 , \61395 , \61396 ,
         \61397 , \61398 , \61399 , \61400 , \61401 , \61402 , \61403 , \61404 , \61405 , \61406 ,
         \61407 , \61408 , \61409 , \61410 , \61411 , \61412 , \61413 , \61414 , \61415 , \61416 ,
         \61417 , \61418 , \61419 , \61420 , \61421 , \61422 , \61423 , \61424 , \61425 , \61426 ,
         \61427 , \61428 , \61429 , \61430 , \61431 , \61432 , \61433 , \61434 , \61435 , \61436 ,
         \61437 , \61438 , \61439 , \61440 , \61441 , \61442 , \61443 , \61444 , \61445 , \61446 ,
         \61447 , \61448 , \61449 , \61450 , \61451 , \61452 , \61453 , \61454 , \61455 , \61456 ,
         \61457 , \61458 , \61459 , \61460 , \61461 , \61462 , \61463 , \61464 , \61465 , \61466 ,
         \61467 , \61468 , \61469 , \61470 , \61471 , \61472 , \61473 , \61474 , \61475 , \61476 ,
         \61477 , \61478 , \61479 , \61480 , \61481 , \61482 , \61483 , \61484 , \61485 , \61486 ,
         \61487 , \61488 , \61489 , \61490 , \61491 , \61492 , \61493 , \61494 , \61495 , \61496 ,
         \61497 , \61498 , \61499 , \61500 , \61501 , \61502 , \61503 , \61504 , \61505 , \61506 ,
         \61507 , \61508 , \61509 , \61510 , \61511 , \61512 , \61513 , \61514 , \61515 , \61516 ,
         \61517 , \61518 , \61519 , \61520 , \61521 , \61522 , \61523 , \61524 , \61525 , \61526 ,
         \61527 , \61528 , \61529 , \61530 , \61531 , \61532 , \61533 , \61534 , \61535 , \61536 ,
         \61537 , \61538 , \61539 , \61540 , \61541 , \61542 , \61543 , \61544 , \61545 , \61546 ,
         \61547 , \61548 , \61549 , \61550 , \61551 , \61552 , \61553 , \61554 , \61555 , \61556 ,
         \61557 , \61558 , \61559 , \61560 , \61561 , \61562 , \61563 , \61564 , \61565 , \61566 ,
         \61567 , \61568 , \61569 , \61570 , \61571 , \61572 , \61573 , \61574 , \61575 , \61576 ,
         \61577 , \61578 , \61579 , \61580 , \61581 , \61582 , \61583 , \61584 , \61585 , \61586 ,
         \61587 , \61588 , \61589 , \61590 , \61591 , \61592 , \61593 , \61594 , \61595 , \61596 ,
         \61597 , \61598 , \61599 , \61600 , \61601 , \61602 , \61603 , \61604 , \61605 , \61606 ,
         \61607 , \61608 , \61609 , \61610 , \61611 , \61612 , \61613 , \61614 , \61615 , \61616 ,
         \61617 , \61618 , \61619 , \61620 , \61621 , \61622 , \61623 , \61624 , \61625 , \61626 ,
         \61627 , \61628 , \61629 , \61630 , \61631 , \61632 , \61633 , \61634 , \61635 , \61636 ,
         \61637 , \61638 , \61639 , \61640 , \61641 , \61642 , \61643 , \61644 , \61645 , \61646 ,
         \61647 , \61648 , \61649 , \61650 , \61651 , \61652 , \61653 , \61654 , \61655 , \61656 ,
         \61657 , \61658 , \61659 , \61660 , \61661 , \61662 , \61663 , \61664 , \61665 , \61666 ,
         \61667 , \61668 , \61669 , \61670 , \61671 , \61672 , \61673 , \61674 , \61675 , \61676 ,
         \61677 , \61678 , \61679 , \61680 , \61681 , \61682 , \61683 , \61684 , \61685 , \61686 ,
         \61687 , \61688 , \61689 , \61690 , \61691 , \61692 , \61693 , \61694 , \61695 , \61696 ,
         \61697 , \61698 , \61699 , \61700 , \61701 , \61702 , \61703 , \61704 , \61705 , \61706 ,
         \61707 , \61708 , \61709 , \61710 , \61711 , \61712 , \61713 , \61714 , \61715 , \61716 ,
         \61717 , \61718 , \61719 , \61720 , \61721 , \61722 , \61723 , \61724 , \61725 , \61726 ,
         \61727 , \61728 , \61729 , \61730 , \61731 , \61732 , \61733 , \61734 , \61735 , \61736 ,
         \61737 , \61738 , \61739 , \61740 , \61741 , \61742 , \61743 , \61744 , \61745 , \61746 ,
         \61747 , \61748 , \61749 , \61750 , \61751 , \61752 , \61753 , \61754 , \61755 , \61756 ,
         \61757 , \61758 , \61759 , \61760 , \61761 , \61762 , \61763 , \61764 , \61765 , \61766 ,
         \61767 , \61768 , \61769 , \61770 , \61771 , \61772 , \61773 , \61774 , \61775 , \61776 ,
         \61777 , \61778 , \61779 , \61780 , \61781 , \61782 , \61783 , \61784 , \61785 , \61786 ,
         \61787 , \61788 , \61789 , \61790 , \61791 , \61792 , \61793 , \61794 , \61795 , \61796 ,
         \61797 , \61798 , \61799 , \61800 , \61801 , \61802 , \61803 , \61804 , \61805 , \61806 ,
         \61807 , \61808 , \61809 , \61810 , \61811 , \61812 , \61813 , \61814 , \61815 , \61816 ,
         \61817 , \61818 , \61819 , \61820 , \61821 , \61822 , \61823 , \61824 , \61825 , \61826 ,
         \61827 , \61828 , \61829 , \61830 , \61831 , \61832 , \61833 , \61834 , \61835 , \61836 ,
         \61837 , \61838 , \61839 , \61840 , \61841 , \61842 , \61843 , \61844 , \61845 , \61846 ,
         \61847 , \61848 , \61849 , \61850 , \61851 , \61852 , \61853 , \61854 , \61855 , \61856 ,
         \61857 , \61858 , \61859 , \61860 , \61861 , \61862 , \61863 , \61864 , \61865 , \61866 ,
         \61867 , \61868 , \61869 , \61870 , \61871 , \61872 , \61873 , \61874 , \61875 , \61876 ,
         \61877 , \61878 , \61879 , \61880 , \61881 , \61882 , \61883 , \61884 , \61885 , \61886 ,
         \61887 , \61888 , \61889 , \61890 , \61891 , \61892 , \61893 , \61894 , \61895 , \61896 ,
         \61897 , \61898 , \61899 , \61900 , \61901 , \61902 , \61903 , \61904 , \61905 , \61906 ,
         \61907 , \61908 , \61909 , \61910 , \61911 , \61912 , \61913 , \61914 , \61915 , \61916 ,
         \61917 , \61918 , \61919 , \61920 , \61921 , \61922 , \61923 , \61924 , \61925 , \61926 ,
         \61927 , \61928 , \61929 , \61930 , \61931 , \61932 , \61933 , \61934 , \61935 , \61936 ,
         \61937 , \61938 , \61939 , \61940 , \61941 , \61942 , \61943 , \61944 , \61945 , \61946 ,
         \61947 , \61948 , \61949 , \61950 , \61951 , \61952 , \61953 , \61954 , \61955 , \61956 ,
         \61957 , \61958 , \61959 , \61960 , \61961 , \61962 , \61963 , \61964 , \61965 , \61966 ,
         \61967 , \61968 , \61969 , \61970 , \61971 , \61972 , \61973 , \61974 , \61975 , \61976 ,
         \61977 , \61978 , \61979 , \61980 , \61981 , \61982 , \61983 , \61984 , \61985 , \61986 ,
         \61987 , \61988 , \61989 , \61990 , \61991 , \61992 , \61993 , \61994 , \61995 , \61996 ,
         \61997 , \61998 , \61999 , \62000 , \62001 , \62002 , \62003 , \62004 , \62005 , \62006 ,
         \62007 , \62008 , \62009 , \62010 , \62011 , \62012 , \62013 , \62014 , \62015 , \62016 ,
         \62017 , \62018 , \62019 , \62020 , \62021 , \62022 , \62023 , \62024 , \62025 , \62026 ,
         \62027 , \62028 , \62029 , \62030 , \62031 , \62032 , \62033 , \62034 , \62035 , \62036 ,
         \62037 , \62038 , \62039 , \62040 , \62041 , \62042 , \62043 , \62044 , \62045 , \62046 ,
         \62047 , \62048 , \62049 , \62050 , \62051 , \62052 , \62053 , \62054 , \62055 , \62056 ,
         \62057 , \62058 , \62059 , \62060 , \62061 , \62062 , \62063 , \62064 , \62065 , \62066 ,
         \62067 , \62068 , \62069 , \62070 , \62071 , \62072 , \62073 , \62074 , \62075 , \62076 ,
         \62077 , \62078 , \62079 , \62080 , \62081 , \62082 , \62083 , \62084 , \62085 , \62086 ,
         \62087 , \62088 , \62089 , \62090 , \62091 , \62092 , \62093 , \62094 , \62095 , \62096 ,
         \62097 , \62098 , \62099 , \62100 , \62101 , \62102 , \62103 , \62104 , \62105 , \62106 ,
         \62107 , \62108 , \62109 , \62110 , \62111 , \62112 , \62113 , \62114 , \62115 , \62116 ,
         \62117 , \62118 , \62119 , \62120 , \62121 , \62122 , \62123 , \62124 , \62125 , \62126 ,
         \62127 , \62128 , \62129 , \62130 , \62131 , \62132 , \62133 , \62134 , \62135 , \62136 ,
         \62137 , \62138 , \62139 , \62140 , \62141 , \62142 , \62143 , \62144 , \62145 , \62146 ,
         \62147 , \62148 , \62149 , \62150 , \62151 , \62152 , \62153 , \62154 , \62155 , \62156 ,
         \62157 , \62158 , \62159 , \62160 , \62161 , \62162 , \62163 , \62164 , \62165 , \62166 ,
         \62167 , \62168 , \62169 , \62170 , \62171 , \62172 , \62173 , \62174 , \62175 , \62176 ,
         \62177 , \62178 , \62179 , \62180 , \62181 , \62182 , \62183 , \62184 , \62185 , \62186 ,
         \62187 , \62188 , \62189 , \62190 , \62191 , \62192 , \62193 , \62194 , \62195 , \62196 ,
         \62197 , \62198 , \62199 , \62200 , \62201 , \62202 , \62203 , \62204 , \62205 , \62206 ,
         \62207 , \62208 , \62209 , \62210 , \62211 , \62212 , \62213 , \62214 , \62215 , \62216 ,
         \62217 , \62218 , \62219 , \62220 , \62221 , \62222 , \62223 , \62224 , \62225 , \62226 ,
         \62227 , \62228 , \62229 , \62230 , \62231 , \62232 , \62233 , \62234 , \62235 , \62236 ,
         \62237 , \62238 , \62239 , \62240 , \62241 , \62242 , \62243 , \62244 , \62245 , \62246 ,
         \62247 , \62248 , \62249 , \62250 , \62251 , \62252 , \62253 , \62254 , \62255 , \62256 ,
         \62257 , \62258 , \62259 , \62260 , \62261 , \62262 , \62263 , \62264 , \62265 , \62266 ,
         \62267 , \62268 , \62269 , \62270 , \62271 , \62272 , \62273 , \62274 , \62275 , \62276 ,
         \62277 , \62278 , \62279 , \62280 , \62281 , \62282 , \62283 , \62284 , \62285 , \62286 ,
         \62287 , \62288 , \62289 , \62290 , \62291 , \62292 , \62293 , \62294 , \62295 , \62296 ,
         \62297 , \62298 , \62299 , \62300 , \62301 , \62302 , \62303 , \62304 , \62305 , \62306 ,
         \62307 , \62308 , \62309 , \62310 , \62311 , \62312 , \62313 , \62314 , \62315 , \62316 ,
         \62317 , \62318 , \62319 , \62320 , \62321 , \62322 , \62323 , \62324 , \62325 , \62326 ,
         \62327 , \62328 , \62329 , \62330 , \62331 , \62332 , \62333 , \62334 , \62335 , \62336 ,
         \62337 , \62338 , \62339 , \62340 , \62341 , \62342 , \62343 , \62344 , \62345 , \62346 ,
         \62347 , \62348 , \62349 , \62350 , \62351 , \62352 , \62353 , \62354 , \62355 , \62356 ,
         \62357 , \62358 , \62359 , \62360 , \62361 , \62362 , \62363 , \62364 , \62365 , \62366 ,
         \62367 , \62368 , \62369 , \62370 , \62371 , \62372 , \62373 , \62374 , \62375 , \62376 ,
         \62377 , \62378 , \62379 , \62380 , \62381 , \62382 , \62383 , \62384 , \62385 , \62386 ,
         \62387 , \62388 , \62389 , \62390 , \62391 , \62392 , \62393 , \62394 , \62395 , \62396 ,
         \62397 , \62398 , \62399 , \62400 , \62401 , \62402 , \62403 , \62404 , \62405 , \62406 ,
         \62407 , \62408 , \62409 , \62410 , \62411 , \62412 , \62413 , \62414 , \62415 , \62416 ,
         \62417 , \62418 , \62419 , \62420 , \62421 , \62422 , \62423 , \62424 , \62425 , \62426 ,
         \62427 , \62428 , \62429 , \62430 , \62431 , \62432 , \62433 , \62434 , \62435 , \62436 ,
         \62437 , \62438 , \62439 , \62440 , \62441 , \62442 , \62443 , \62444 , \62445 , \62446 ,
         \62447 , \62448 , \62449 , \62450 , \62451 , \62452 , \62453 , \62454 , \62455 , \62456 ,
         \62457 , \62458 , \62459 , \62460 , \62461 , \62462 , \62463 , \62464 , \62465 , \62466 ,
         \62467 , \62468 , \62469 , \62470 , \62471 , \62472 , \62473 , \62474 , \62475 , \62476 ,
         \62477 , \62478 , \62479 , \62480 , \62481 , \62482 , \62483 , \62484 , \62485 , \62486 ,
         \62487 , \62488 , \62489 , \62490 , \62491 , \62492 , \62493 , \62494 , \62495 , \62496 ,
         \62497 , \62498 , \62499 , \62500 , \62501 , \62502 , \62503 , \62504 , \62505 , \62506 ,
         \62507 , \62508 , \62509 , \62510 , \62511 , \62512 , \62513 , \62514 , \62515 , \62516 ,
         \62517 , \62518 , \62519 , \62520 , \62521 , \62522 , \62523 , \62524 , \62525 , \62526 ,
         \62527 , \62528 , \62529 , \62530 , \62531 , \62532 , \62533 , \62534 , \62535 , \62536 ,
         \62537 , \62538 , \62539 , \62540 , \62541 , \62542 , \62543 , \62544 , \62545 , \62546 ,
         \62547 , \62548 , \62549 , \62550 , \62551 , \62552 , \62553 , \62554 , \62555 , \62556 ,
         \62557 , \62558 , \62559 , \62560 , \62561 , \62562 , \62563 , \62564 , \62565 , \62566 ,
         \62567 , \62568 , \62569 , \62570 , \62571 , \62572 , \62573 , \62574 , \62575 , \62576 ,
         \62577 , \62578 , \62579 , \62580 , \62581 , \62582 , \62583 , \62584 , \62585 , \62586 ,
         \62587 , \62588 , \62589 , \62590 , \62591 , \62592 , \62593 , \62594 , \62595 , \62596 ,
         \62597 , \62598 , \62599 , \62600 , \62601 , \62602 , \62603 , \62604 , \62605 , \62606 ,
         \62607 , \62608 , \62609 , \62610 , \62611 , \62612 , \62613 , \62614 , \62615 , \62616 ,
         \62617 , \62618 , \62619 , \62620 , \62621 , \62622 , \62623 , \62624 , \62625 , \62626 ,
         \62627 , \62628 , \62629 , \62630 , \62631 , \62632 , \62633 , \62634 , \62635 , \62636 ,
         \62637 , \62638 , \62639 , \62640 , \62641 , \62642 , \62643 , \62644 , \62645 , \62646 ,
         \62647 , \62648 , \62649 , \62650 , \62651 , \62652 , \62653 , \62654 , \62655 , \62656 ,
         \62657 , \62658 , \62659 , \62660 , \62661 , \62662 , \62663 , \62664 , \62665 , \62666 ,
         \62667 , \62668 , \62669 , \62670 , \62671 , \62672 , \62673 , \62674 , \62675 , \62676 ,
         \62677 , \62678 , \62679 , \62680 , \62681 , \62682 , \62683 , \62684 , \62685 , \62686 ,
         \62687 , \62688 , \62689 , \62690 , \62691 , \62692 , \62693 , \62694 , \62695 , \62696 ,
         \62697 , \62698 , \62699 , \62700 , \62701 , \62702 , \62703 , \62704 , \62705 , \62706 ,
         \62707 , \62708 , \62709 , \62710 , \62711 , \62712 , \62713 , \62714 , \62715 , \62716 ,
         \62717 , \62718 , \62719 , \62720 , \62721 , \62722 , \62723 , \62724 , \62725 , \62726 ,
         \62727 , \62728 , \62729 , \62730 , \62731 , \62732 , \62733 , \62734 , \62735 , \62736 ,
         \62737 , \62738 , \62739 , \62740 , \62741 , \62742 , \62743 , \62744 , \62745 , \62746 ,
         \62747 , \62748 , \62749 , \62750 , \62751 , \62752 , \62753 , \62754 , \62755 , \62756 ,
         \62757 , \62758 , \62759 , \62760 , \62761 , \62762 , \62763 , \62764 , \62765 , \62766 ,
         \62767 , \62768 , \62769 , \62770 , \62771 , \62772 , \62773 , \62774 , \62775 , \62776 ,
         \62777 , \62778 , \62779 , \62780 , \62781 , \62782 , \62783 , \62784 , \62785 , \62786 ,
         \62787 , \62788 , \62789 , \62790 , \62791 , \62792 , \62793 , \62794 , \62795 , \62796 ,
         \62797 , \62798 , \62799 , \62800 , \62801 , \62802 , \62803 , \62804 , \62805 , \62806 ,
         \62807 , \62808 , \62809 , \62810 , \62811 , \62812 , \62813 , \62814 , \62815 , \62816 ,
         \62817 , \62818 , \62819 , \62820 , \62821 , \62822 , \62823 , \62824 , \62825 , \62826 ,
         \62827 , \62828 , \62829 , \62830 , \62831 , \62832 , \62833 , \62834 , \62835 , \62836 ,
         \62837 , \62838 , \62839 , \62840 , \62841 , \62842 , \62843 , \62844 , \62845 , \62846 ,
         \62847 , \62848 , \62849 , \62850 , \62851 , \62852 , \62853 , \62854 , \62855 , \62856 ,
         \62857 , \62858 , \62859 , \62860 , \62861 , \62862 , \62863 , \62864 , \62865 , \62866 ,
         \62867 , \62868 , \62869 , \62870 , \62871 , \62872 , \62873 , \62874 , \62875 , \62876 ,
         \62877 , \62878 , \62879 , \62880 , \62881 , \62882 , \62883 , \62884 , \62885 , \62886 ,
         \62887 , \62888 , \62889 , \62890 , \62891 , \62892 , \62893 , \62894 , \62895 , \62896 ,
         \62897 , \62898 , \62899 , \62900 , \62901 , \62902 , \62903 , \62904 , \62905 , \62906 ,
         \62907 , \62908 , \62909 , \62910 , \62911 , \62912 , \62913 , \62914 , \62915 , \62916 ,
         \62917 , \62918 , \62919 , \62920 , \62921 , \62922 , \62923 , \62924 , \62925 , \62926 ,
         \62927 , \62928 , \62929 , \62930 , \62931 , \62932 , \62933 , \62934 , \62935 , \62936 ,
         \62937 , \62938 , \62939 , \62940 , \62941 , \62942 , \62943 , \62944 , \62945 , \62946 ,
         \62947 , \62948 , \62949 , \62950 , \62951 , \62952 , \62953 , \62954 , \62955 , \62956 ,
         \62957 , \62958 , \62959 , \62960 , \62961 , \62962 , \62963 , \62964 , \62965 , \62966 ,
         \62967 , \62968 , \62969 , \62970 , \62971 , \62972 , \62973 , \62974 , \62975 , \62976 ,
         \62977 , \62978 , \62979 , \62980 , \62981 , \62982 , \62983 , \62984 , \62985 , \62986 ,
         \62987 , \62988 , \62989 , \62990 , \62991 , \62992 , \62993 , \62994 , \62995 , \62996 ,
         \62997 , \62998 , \62999 , \63000 , \63001 , \63002 , \63003 , \63004 , \63005 , \63006 ,
         \63007 , \63008 , \63009 , \63010 , \63011 , \63012 , \63013 , \63014 , \63015 , \63016 ,
         \63017 , \63018 , \63019 , \63020 , \63021 , \63022 , \63023 , \63024 , \63025 , \63026 ,
         \63027 , \63028 , \63029 , \63030 , \63031 , \63032 , \63033 , \63034 , \63035 , \63036 ,
         \63037 , \63038 , \63039 , \63040 , \63041 , \63042 , \63043 , \63044 , \63045 , \63046 ,
         \63047 , \63048 , \63049 , \63050 , \63051 , \63052 , \63053 , \63054 , \63055 , \63056 ,
         \63057 , \63058 , \63059 , \63060 , \63061 , \63062 , \63063 , \63064 , \63065 , \63066 ,
         \63067 , \63068 , \63069 , \63070 , \63071 , \63072 , \63073 , \63074 , \63075 , \63076 ,
         \63077 , \63078 , \63079 , \63080 , \63081 , \63082 , \63083 , \63084 , \63085 , \63086 ,
         \63087 , \63088 , \63089 , \63090 , \63091 , \63092 , \63093 , \63094 , \63095 , \63096 ,
         \63097 , \63098 , \63099 , \63100 , \63101 , \63102 , \63103 , \63104 , \63105 , \63106 ,
         \63107 , \63108 , \63109 , \63110 , \63111 , \63112 , \63113 , \63114 , \63115 , \63116 ,
         \63117 , \63118 , \63119 , \63120 , \63121 , \63122 , \63123 , \63124 , \63125 , \63126 ,
         \63127 , \63128 , \63129 , \63130 , \63131 , \63132 , \63133 , \63134 , \63135 , \63136 ,
         \63137 , \63138 , \63139 , \63140 , \63141 , \63142 , \63143 , \63144 , \63145 , \63146 ,
         \63147 , \63148 , \63149 , \63150 , \63151 , \63152 , \63153 , \63154 , \63155 , \63156 ,
         \63157 , \63158 , \63159 , \63160 , \63161 , \63162 , \63163 , \63164 , \63165 , \63166 ,
         \63167 , \63168 , \63169 , \63170 , \63171 , \63172 , \63173 , \63174 , \63175 , \63176 ,
         \63177 , \63178 , \63179 , \63180 , \63181 , \63182 , \63183 , \63184 , \63185 , \63186 ,
         \63187 , \63188 , \63189 , \63190 , \63191 , \63192 , \63193 , \63194 , \63195 , \63196 ,
         \63197 , \63198 , \63199 , \63200 , \63201 , \63202 , \63203 , \63204 , \63205 , \63206 ,
         \63207 , \63208 , \63209 , \63210 , \63211 , \63212 , \63213 , \63214 , \63215 , \63216 ,
         \63217 , \63218 , \63219 , \63220 , \63221 , \63222 , \63223 , \63224 , \63225 , \63226 ,
         \63227 , \63228 , \63229 , \63230 , \63231 , \63232 , \63233 , \63234 , \63235 , \63236 ,
         \63237 , \63238 , \63239 , \63240 , \63241 , \63242 , \63243 , \63244 , \63245 , \63246 ,
         \63247 , \63248 , \63249 , \63250 , \63251 , \63252 , \63253 , \63254 , \63255 , \63256 ,
         \63257 , \63258 , \63259 , \63260 , \63261 , \63262 , \63263 , \63264 , \63265 , \63266 ,
         \63267 , \63268 , \63269 , \63270 , \63271 , \63272 , \63273 , \63274 , \63275 , \63276 ,
         \63277 , \63278 , \63279 , \63280 , \63281 , \63282 , \63283 , \63284 , \63285 , \63286 ,
         \63287 , \63288 , \63289 , \63290 , \63291 , \63292 , \63293 , \63294 , \63295 , \63296 ,
         \63297 , \63298 , \63299 , \63300 , \63301 , \63302 , \63303 , \63304 , \63305 , \63306 ,
         \63307 , \63308 , \63309 , \63310 , \63311 , \63312 , \63313 , \63314 , \63315 , \63316 ,
         \63317 , \63318 , \63319 , \63320 , \63321 , \63322 , \63323 , \63324 , \63325 , \63326 ,
         \63327 , \63328 , \63329 , \63330 , \63331 , \63332 , \63333 , \63334 , \63335 , \63336 ,
         \63337 , \63338 , \63339 , \63340 , \63341 , \63342 , \63343 , \63344 , \63345 , \63346 ,
         \63347 , \63348 , \63349 , \63350 , \63351 , \63352 , \63353 , \63354 , \63355 , \63356 ,
         \63357 , \63358 , \63359 , \63360 , \63361 , \63362 , \63363 , \63364 , \63365 , \63366 ,
         \63367 , \63368 , \63369 , \63370 , \63371 , \63372 , \63373 , \63374 , \63375 , \63376 ,
         \63377 , \63378 , \63379 , \63380 , \63381 , \63382 , \63383 , \63384 , \63385 , \63386 ,
         \63387 , \63388 , \63389 , \63390 , \63391 , \63392 , \63393 , \63394 , \63395 , \63396 ,
         \63397 , \63398 , \63399 , \63400 , \63401 , \63402 , \63403 , \63404 , \63405 , \63406 ,
         \63407 , \63408 , \63409 , \63410 , \63411 , \63412 , \63413 , \63414 , \63415 , \63416 ,
         \63417 , \63418 , \63419 , \63420 , \63421 , \63422 , \63423 , \63424 , \63425 , \63426 ,
         \63427 , \63428 , \63429 , \63430 , \63431 , \63432 , \63433 , \63434 , \63435 , \63436 ,
         \63437 , \63438 , \63439 , \63440 , \63441 , \63442 , \63443 , \63444 , \63445 , \63446 ,
         \63447 , \63448 , \63449 , \63450 , \63451 , \63452 , \63453 , \63454 , \63455 , \63456 ,
         \63457 , \63458 , \63459 , \63460 , \63461 , \63462 , \63463 , \63464 , \63465 , \63466 ,
         \63467 , \63468 , \63469 , \63470 , \63471 , \63472 , \63473 , \63474 , \63475 , \63476 ,
         \63477 , \63478 , \63479 , \63480 , \63481 , \63482 , \63483 , \63484 , \63485 , \63486 ,
         \63487 , \63488 , \63489 , \63490 , \63491 , \63492 , \63493 , \63494 , \63495 , \63496 ,
         \63497 , \63498 , \63499 , \63500 , \63501 , \63502 , \63503 , \63504 , \63505 , \63506 ,
         \63507 , \63508 , \63509 , \63510 , \63511 , \63512 , \63513 , \63514 , \63515 , \63516 ,
         \63517 , \63518 , \63519 , \63520 , \63521 , \63522 , \63523 , \63524 , \63525 , \63526 ,
         \63527 , \63528 , \63529 , \63530 , \63531 , \63532 , \63533 , \63534 , \63535 , \63536 ,
         \63537 , \63538 , \63539 , \63540 , \63541 , \63542 , \63543 , \63544 , \63545 , \63546 ,
         \63547 , \63548 , \63549 , \63550 , \63551 , \63552 , \63553 , \63554 , \63555 , \63556 ,
         \63557 , \63558 , \63559 , \63560 , \63561 , \63562 , \63563 , \63564 , \63565 , \63566 ,
         \63567 , \63568 , \63569 , \63570 , \63571 , \63572 , \63573 , \63574 , \63575 , \63576 ,
         \63577 , \63578 , \63579 , \63580 , \63581 , \63582 , \63583 , \63584 , \63585 , \63586 ,
         \63587 , \63588 , \63589 , \63590 , \63591 , \63592 , \63593 , \63594 , \63595 , \63596 ,
         \63597 , \63598 , \63599 , \63600 , \63601 , \63602 , \63603 , \63604 , \63605 , \63606 ,
         \63607 , \63608 , \63609 , \63610 , \63611 , \63612 , \63613 , \63614 , \63615 , \63616 ,
         \63617 , \63618 , \63619 , \63620 , \63621 , \63622 , \63623 , \63624 , \63625 , \63626 ,
         \63627 , \63628 , \63629 , \63630 , \63631 , \63632 , \63633 , \63634 , \63635 , \63636 ,
         \63637 , \63638 , \63639 , \63640 , \63641 , \63642 , \63643 , \63644 , \63645 , \63646 ,
         \63647 , \63648 , \63649 , \63650 , \63651 , \63652 , \63653 , \63654 , \63655 , \63656 ,
         \63657 , \63658 , \63659 , \63660 , \63661 , \63662 , \63663 , \63664 , \63665 , \63666 ,
         \63667 , \63668 , \63669 , \63670 , \63671 , \63672 , \63673 , \63674 , \63675 , \63676 ,
         \63677 , \63678 , \63679 , \63680 , \63681 , \63682 , \63683 , \63684 , \63685 , \63686 ,
         \63687 , \63688 , \63689 , \63690 , \63691 , \63692 , \63693 , \63694 , \63695 , \63696 ,
         \63697 , \63698 , \63699 , \63700 , \63701 , \63702 , \63703 , \63704 , \63705 , \63706 ,
         \63707 , \63708 , \63709 , \63710 , \63711 , \63712 , \63713 , \63714 , \63715 , \63716 ,
         \63717 , \63718 , \63719 , \63720 , \63721 , \63722 , \63723 , \63724 , \63725 , \63726 ,
         \63727 , \63728 , \63729 , \63730 , \63731 , \63732 , \63733 , \63734 , \63735 , \63736 ,
         \63737 , \63738 , \63739 , \63740 , \63741 , \63742 , \63743 , \63744 , \63745 , \63746 ,
         \63747 , \63748 , \63749 , \63750 , \63751 , \63752 , \63753 , \63754 , \63755 , \63756 ,
         \63757 , \63758 , \63759 , \63760 , \63761 , \63762 , \63763 , \63764 , \63765 , \63766 ,
         \63767 , \63768 , \63769 , \63770 , \63771 , \63772 , \63773 , \63774 , \63775 , \63776 ,
         \63777 , \63778 , \63779 , \63780 , \63781 , \63782 , \63783 , \63784 , \63785 , \63786 ,
         \63787 , \63788 , \63789 , \63790 , \63791 , \63792 , \63793 , \63794 , \63795 , \63796 ,
         \63797 , \63798 , \63799 , \63800 , \63801 , \63802 , \63803 , \63804 , \63805 , \63806 ,
         \63807 , \63808 , \63809 , \63810 , \63811 , \63812 , \63813 , \63814 , \63815 , \63816 ,
         \63817 , \63818 , \63819 , \63820 , \63821 , \63822 , \63823 , \63824 , \63825 , \63826 ,
         \63827 , \63828 , \63829 , \63830 , \63831 , \63832 , \63833 , \63834 , \63835 , \63836 ,
         \63837 , \63838 , \63839 , \63840 , \63841 , \63842 , \63843 , \63844 , \63845 , \63846 ,
         \63847 , \63848 , \63849 , \63850 , \63851 , \63852 , \63853 , \63854 , \63855 , \63856 ,
         \63857 , \63858 , \63859 , \63860 , \63861 , \63862 , \63863 , \63864 , \63865 , \63866 ,
         \63867 , \63868 , \63869 , \63870 , \63871 , \63872 , \63873 , \63874 , \63875 , \63876 ,
         \63877 , \63878 , \63879 , \63880 , \63881 , \63882 , \63883 , \63884 , \63885 , \63886 ,
         \63887 , \63888 , \63889 , \63890 , \63891 , \63892 , \63893 , \63894 , \63895 , \63896 ,
         \63897 , \63898 , \63899 , \63900 , \63901 , \63902 , \63903 , \63904 , \63905 , \63906 ,
         \63907 , \63908 , \63909 , \63910 , \63911 , \63912 , \63913 , \63914 , \63915 , \63916 ,
         \63917 , \63918 , \63919 , \63920 , \63921 , \63922 , \63923 , \63924 , \63925 , \63926 ,
         \63927 , \63928 , \63929 , \63930 , \63931 , \63932 , \63933 , \63934 , \63935 , \63936 ,
         \63937 , \63938 , \63939 , \63940 , \63941 , \63942 , \63943 , \63944 , \63945 , \63946 ,
         \63947 , \63948 , \63949 , \63950 , \63951 , \63952 , \63953 , \63954 , \63955 , \63956 ,
         \63957 , \63958 , \63959 , \63960 , \63961 , \63962 , \63963 , \63964 , \63965 , \63966 ,
         \63967 , \63968 , \63969 , \63970 , \63971 , \63972 , \63973 , \63974 , \63975 , \63976 ,
         \63977 , \63978 , \63979 , \63980 , \63981 , \63982 , \63983 , \63984 , \63985 , \63986 ,
         \63987 , \63988 , \63989 , \63990 , \63991 , \63992 , \63993 , \63994 , \63995 , \63996 ,
         \63997 , \63998 , \63999 , \64000 , \64001 , \64002 , \64003 , \64004 , \64005 , \64006 ,
         \64007 , \64008 , \64009 , \64010 , \64011 , \64012 , \64013 , \64014 , \64015 , \64016 ,
         \64017 , \64018 , \64019 , \64020 , \64021 , \64022 , \64023 , \64024 , \64025 , \64026 ,
         \64027 , \64028 , \64029 , \64030 , \64031 , \64032 , \64033 , \64034 , \64035 , \64036 ,
         \64037 , \64038 , \64039 , \64040 , \64041 , \64042 , \64043 , \64044 , \64045 , \64046 ,
         \64047 , \64048 , \64049 , \64050 , \64051 , \64052 , \64053 , \64054 , \64055 , \64056 ,
         \64057 , \64058 , \64059 , \64060 , \64061 , \64062 , \64063 , \64064 , \64065 , \64066 ,
         \64067 , \64068 , \64069 , \64070 , \64071 , \64072 , \64073 , \64074 , \64075 , \64076 ,
         \64077 , \64078 , \64079 , \64080 , \64081 , \64082 , \64083 , \64084 , \64085 , \64086 ,
         \64087 , \64088 , \64089 , \64090 , \64091 , \64092 , \64093 , \64094 , \64095 , \64096 ,
         \64097 , \64098 , \64099 , \64100 , \64101 , \64102 , \64103 , \64104 , \64105 , \64106 ,
         \64107 , \64108 , \64109 , \64110 , \64111 , \64112 , \64113 , \64114 , \64115 , \64116 ,
         \64117 , \64118 , \64119 , \64120 , \64121 , \64122 , \64123 , \64124 , \64125 , \64126 ,
         \64127 , \64128 , \64129 , \64130 , \64131 , \64132 , \64133 , \64134 , \64135 , \64136 ,
         \64137 , \64138 , \64139 , \64140 , \64141 , \64142 , \64143 , \64144 , \64145 , \64146 ,
         \64147 , \64148 , \64149 , \64150 , \64151 , \64152 , \64153 , \64154 , \64155 , \64156 ,
         \64157 , \64158 , \64159 , \64160 , \64161 , \64162 , \64163 , \64164 , \64165 , \64166 ,
         \64167 , \64168 , \64169 , \64170 , \64171 , \64172 , \64173 , \64174 , \64175 , \64176 ,
         \64177 , \64178 , \64179 , \64180 , \64181 , \64182 , \64183 , \64184 , \64185 , \64186 ,
         \64187 , \64188 , \64189 , \64190 , \64191 , \64192 , \64193 , \64194 , \64195 , \64196 ,
         \64197 , \64198 , \64199 , \64200 , \64201 , \64202 , \64203 , \64204 , \64205 , \64206 ,
         \64207 , \64208 , \64209 , \64210 , \64211 , \64212 , \64213 , \64214 , \64215 , \64216 ,
         \64217 , \64218 , \64219 , \64220 , \64221 , \64222 , \64223 , \64224 , \64225 , \64226 ,
         \64227 , \64228 , \64229 , \64230 , \64231 , \64232 , \64233 , \64234 , \64235 , \64236 ,
         \64237 , \64238 , \64239 , \64240 , \64241 , \64242 , \64243 , \64244 , \64245 , \64246 ,
         \64247 , \64248 , \64249 , \64250 , \64251 , \64252 , \64253 , \64254 , \64255 , \64256 ,
         \64257 , \64258 , \64259 , \64260 , \64261 , \64262 , \64263 , \64264 , \64265 , \64266 ,
         \64267 , \64268 , \64269 , \64270 , \64271 , \64272 , \64273 , \64274 , \64275 , \64276 ,
         \64277 , \64278 , \64279 , \64280 , \64281 , \64282 , \64283 , \64284 , \64285 , \64286 ,
         \64287 , \64288 , \64289 , \64290 , \64291 , \64292 , \64293 , \64294 , \64295 , \64296 ,
         \64297 , \64298 , \64299 , \64300 , \64301 , \64302 , \64303 , \64304 , \64305 , \64306 ,
         \64307 , \64308 , \64309 , \64310 , \64311 , \64312 , \64313 , \64314 , \64315 , \64316 ,
         \64317 , \64318 , \64319 , \64320 , \64321 , \64322 , \64323 , \64324 , \64325 , \64326 ,
         \64327 , \64328 , \64329 , \64330 , \64331 , \64332 , \64333 , \64334 , \64335 , \64336 ,
         \64337 , \64338 , \64339 , \64340 , \64341 , \64342 , \64343 , \64344 , \64345 , \64346 ,
         \64347 , \64348 , \64349 , \64350 , \64351 , \64352 , \64353 , \64354 , \64355 , \64356 ,
         \64357 , \64358 , \64359 , \64360 , \64361 , \64362 , \64363 , \64364 , \64365 , \64366 ,
         \64367 , \64368 , \64369 , \64370 , \64371 , \64372 , \64373 , \64374 , \64375 , \64376 ,
         \64377 , \64378 , \64379 , \64380 , \64381 , \64382 , \64383 , \64384 , \64385 , \64386 ,
         \64387 , \64388 , \64389 , \64390 , \64391 , \64392 , \64393 , \64394 , \64395 , \64396 ,
         \64397 , \64398 , \64399 , \64400 , \64401 , \64402 , \64403 , \64404 , \64405 , \64406 ,
         \64407 , \64408 , \64409 , \64410 , \64411 , \64412 , \64413 , \64414 , \64415 , \64416 ,
         \64417 , \64418 , \64419 , \64420 , \64421 , \64422 , \64423 , \64424 , \64425 , \64426 ,
         \64427 , \64428 , \64429 , \64430 , \64431 , \64432 , \64433 , \64434 , \64435 , \64436 ,
         \64437 , \64438 , \64439 , \64440 , \64441 , \64442 , \64443 , \64444 , \64445 , \64446 ,
         \64447 , \64448 , \64449 , \64450 , \64451 , \64452 , \64453 , \64454 , \64455 , \64456 ,
         \64457 , \64458 , \64459 , \64460 , \64461 , \64462 , \64463 , \64464 , \64465 , \64466 ,
         \64467 , \64468 , \64469 , \64470 , \64471 , \64472 , \64473 , \64474 , \64475 , \64476 ,
         \64477 , \64478 , \64479 , \64480 , \64481 , \64482 , \64483 , \64484 , \64485 , \64486 ,
         \64487 , \64488 , \64489 , \64490 , \64491 , \64492 , \64493 , \64494 , \64495 , \64496 ,
         \64497 , \64498 , \64499 , \64500 , \64501 , \64502 , \64503 , \64504 , \64505 , \64506 ,
         \64507 , \64508 , \64509 , \64510 , \64511 , \64512 , \64513 , \64514 , \64515 , \64516 ,
         \64517 , \64518 , \64519 , \64520 , \64521 , \64522 , \64523 , \64524 , \64525 , \64526 ,
         \64527 , \64528 , \64529 , \64530 , \64531 , \64532 , \64533 , \64534 , \64535 , \64536 ,
         \64537 , \64538 , \64539 , \64540 , \64541 , \64542 , \64543 , \64544 , \64545 , \64546 ,
         \64547 , \64548 , \64549 , \64550 , \64551 , \64552 , \64553 , \64554 , \64555 , \64556 ,
         \64557 , \64558 , \64559 , \64560 , \64561 , \64562 , \64563 , \64564 , \64565 , \64566 ,
         \64567 , \64568 , \64569 , \64570 , \64571 , \64572 , \64573 , \64574 , \64575 , \64576 ,
         \64577 , \64578 , \64579 , \64580 , \64581 , \64582 , \64583 , \64584 , \64585 , \64586 ,
         \64587 , \64588 , \64589 , \64590 , \64591 , \64592 , \64593 , \64594 , \64595 , \64596 ,
         \64597 , \64598 , \64599 , \64600 , \64601 , \64602 , \64603 , \64604 , \64605 , \64606 ,
         \64607 , \64608 , \64609 , \64610 , \64611 , \64612 , \64613 , \64614 , \64615 , \64616 ,
         \64617 , \64618 , \64619 , \64620 , \64621 , \64622 , \64623 , \64624 , \64625 , \64626 ,
         \64627 , \64628 , \64629 , \64630 , \64631 , \64632 , \64633 , \64634 , \64635 , \64636 ,
         \64637 , \64638 , \64639 , \64640 , \64641 , \64642 , \64643 , \64644 , \64645 , \64646 ,
         \64647 , \64648 , \64649 , \64650 , \64651 , \64652 , \64653 , \64654 , \64655 , \64656 ,
         \64657 , \64658 , \64659 , \64660 , \64661 , \64662 , \64663 , \64664 , \64665 , \64666 ,
         \64667 , \64668 , \64669 , \64670 , \64671 , \64672 , \64673 , \64674 , \64675 , \64676 ,
         \64677 , \64678 , \64679 , \64680 , \64681 , \64682 , \64683 , \64684 , \64685 , \64686 ,
         \64687 , \64688 , \64689 , \64690 , \64691 , \64692 , \64693 , \64694 , \64695 , \64696 ,
         \64697 , \64698 , \64699 , \64700 , \64701 , \64702 , \64703 , \64704 , \64705 , \64706 ,
         \64707 , \64708 , \64709 , \64710 , \64711 , \64712 , \64713 , \64714 , \64715 , \64716 ,
         \64717 , \64718 , \64719 , \64720 , \64721 , \64722 , \64723 , \64724 , \64725 , \64726 ,
         \64727 , \64728 , \64729 , \64730 , \64731 , \64732 , \64733 , \64734 , \64735 , \64736 ,
         \64737 , \64738 , \64739 , \64740 , \64741 , \64742 , \64743 , \64744 , \64745 , \64746 ,
         \64747 , \64748 , \64749 , \64750 , \64751 , \64752 , \64753 , \64754 , \64755 , \64756 ,
         \64757 , \64758 , \64759 , \64760 , \64761 , \64762 , \64763 , \64764 , \64765 , \64766 ,
         \64767 , \64768 , \64769 , \64770 , \64771 , \64772 , \64773 , \64774 , \64775 , \64776 ,
         \64777 , \64778 , \64779 , \64780 , \64781 , \64782 , \64783 , \64784 , \64785 , \64786 ,
         \64787 , \64788 , \64789 , \64790 , \64791 , \64792 , \64793 , \64794 , \64795 , \64796 ,
         \64797 , \64798 , \64799 , \64800 , \64801 , \64802 , \64803 , \64804 , \64805 , \64806 ,
         \64807 , \64808 , \64809 , \64810 , \64811 , \64812 , \64813 , \64814 , \64815 , \64816 ,
         \64817 , \64818 , \64819 , \64820 , \64821 , \64822 , \64823 , \64824 , \64825 , \64826 ,
         \64827 , \64828 , \64829 , \64830 , \64831 , \64832 , \64833 , \64834 , \64835 , \64836 ,
         \64837 , \64838 , \64839 , \64840 , \64841 , \64842 , \64843 , \64844 , \64845 , \64846 ,
         \64847 , \64848 , \64849 , \64850 , \64851 , \64852 , \64853 , \64854 , \64855 , \64856 ,
         \64857 , \64858 , \64859 , \64860 , \64861 , \64862 , \64863 , \64864 , \64865 , \64866 ,
         \64867 , \64868 , \64869 , \64870 , \64871 , \64872 , \64873 , \64874 , \64875 , \64876 ,
         \64877 , \64878 , \64879 , \64880 , \64881 , \64882 , \64883 , \64884 , \64885 , \64886 ,
         \64887 , \64888 , \64889 , \64890 , \64891 , \64892 , \64893 , \64894 , \64895 , \64896 ,
         \64897 , \64898 , \64899 , \64900 , \64901 , \64902 , \64903 , \64904 , \64905 , \64906 ,
         \64907 , \64908 , \64909 , \64910 , \64911 , \64912 , \64913 , \64914 , \64915 , \64916 ,
         \64917 , \64918 , \64919 , \64920 , \64921 , \64922 , \64923 , \64924 , \64925 , \64926 ,
         \64927 , \64928 , \64929 , \64930 , \64931 , \64932 , \64933 , \64934 , \64935 , \64936 ,
         \64937 , \64938 , \64939 , \64940 , \64941 , \64942 , \64943 , \64944 , \64945 , \64946 ,
         \64947 , \64948 , \64949 , \64950 , \64951 , \64952 , \64953 , \64954 , \64955 , \64956 ,
         \64957 , \64958 , \64959 , \64960 , \64961 , \64962 , \64963 , \64964 , \64965 , \64966 ,
         \64967 , \64968 , \64969 , \64970 , \64971 , \64972 , \64973 , \64974 , \64975 , \64976 ,
         \64977 , \64978 , \64979 , \64980 , \64981 , \64982 , \64983 , \64984 , \64985 , \64986 ,
         \64987 , \64988 , \64989 , \64990 , \64991 , \64992 , \64993 , \64994 , \64995 , \64996 ,
         \64997 , \64998 , \64999 , \65000 , \65001 , \65002 , \65003 , \65004 , \65005 , \65006 ,
         \65007 , \65008 , \65009 , \65010 , \65011 , \65012 , \65013 , \65014 , \65015 , \65016 ,
         \65017 , \65018 , \65019 , \65020 , \65021 , \65022 , \65023 , \65024 , \65025 , \65026 ,
         \65027 , \65028 , \65029 , \65030 , \65031 , \65032 , \65033 , \65034 , \65035 , \65036 ,
         \65037 , \65038 , \65039 , \65040 , \65041 , \65042 , \65043 , \65044 , \65045 , \65046 ,
         \65047 , \65048 , \65049 , \65050 , \65051 , \65052 , \65053 , \65054 , \65055 , \65056 ,
         \65057 , \65058 , \65059 , \65060 , \65061 , \65062 , \65063 , \65064 , \65065 , \65066 ,
         \65067 , \65068 , \65069 , \65070 , \65071 , \65072 , \65073 , \65074 , \65075 , \65076 ,
         \65077 , \65078 , \65079 , \65080 , \65081 , \65082 , \65083 , \65084 , \65085 , \65086 ,
         \65087 , \65088 , \65089 , \65090 , \65091 , \65092 , \65093 , \65094 , \65095 , \65096 ,
         \65097 , \65098 , \65099 , \65100 , \65101 , \65102 , \65103 , \65104 , \65105 , \65106 ,
         \65107 , \65108 , \65109 , \65110 , \65111 , \65112 , \65113 , \65114 , \65115 , \65116 ,
         \65117 , \65118 , \65119 , \65120 , \65121 , \65122 , \65123 , \65124 , \65125 , \65126 ,
         \65127 , \65128 , \65129 , \65130 , \65131 , \65132 , \65133 , \65134 , \65135 , \65136 ,
         \65137 , \65138 , \65139 , \65140 , \65141 , \65142 , \65143 , \65144 , \65145 , \65146 ,
         \65147 , \65148 , \65149 , \65150 , \65151 , \65152 , \65153 , \65154 , \65155 , \65156 ,
         \65157 , \65158 , \65159 , \65160 , \65161 , \65162 , \65163 , \65164 , \65165 , \65166 ,
         \65167 , \65168 , \65169 , \65170 , \65171 , \65172 , \65173 , \65174 , \65175 , \65176 ,
         \65177 , \65178 , \65179 , \65180 , \65181 , \65182 , \65183 , \65184 , \65185 , \65186 ,
         \65187 , \65188 , \65189 , \65190 , \65191 , \65192 , \65193 , \65194 , \65195 , \65196 ,
         \65197 , \65198 , \65199 , \65200 , \65201 , \65202 , \65203 , \65204 , \65205 , \65206 ,
         \65207 , \65208 , \65209 , \65210 , \65211 , \65212 , \65213 , \65214 , \65215 , \65216 ,
         \65217 , \65218 , \65219 , \65220 , \65221 , \65222 , \65223 , \65224 , \65225 ;
buf \U$labajz7360 ( R_58_102f1b78, \65057 );
buf \U$labajz7361 ( R_59_be1fc68, \65063 );
buf \U$labajz7362 ( R_5a_10279198, \65064 );
buf \U$labajz7363 ( R_5b_102299e8, \65065 );
buf \U$labajz7364 ( R_5c_101d0448, \65066 );
buf \U$labajz7365 ( R_5d_f7f82f0, \65067 );
buf \U$labajz7366 ( R_5e_be21600, \65068 );
buf \U$labajz7367 ( R_5f_f7fa5b8, \65069 );
buf \U$labajz7368 ( R_60_1027d530, \65070 );
buf \U$labajz7369 ( R_61_10205ae8, \65071 );
buf \U$labajz7370 ( R_62_10283510, \65072 );
buf \U$labajz7371 ( R_63_f82b578, \65073 );
buf \U$labajz7372 ( R_64_ace4e68, \65074 );
buf \U$labajz7373 ( R_65_f8204e0, \65075 );
buf \U$labajz7374 ( R_66_1027a0b0, \65080 );
buf \U$labajz7375 ( R_67_1022dc30, \65081 );
buf \U$labajz7376 ( R_68_102478a8, \65082 );
buf \U$labajz7377 ( R_69_10286f78, \65083 );
buf \U$labajz7378 ( R_6a_f7edd80, \65084 );
buf \U$labajz7379 ( R_6b_101c3628, \65085 );
buf \U$labajz7380 ( R_6c_f7fbe00, \65086 );
buf \U$labajz7381 ( R_6d_f7ce9f8, \65087 );
buf \U$labajz7382 ( R_6e_f7c8830, \65088 );
buf \U$labajz7383 ( R_6f_101ffc68, \65089 );
buf \U$labajz7384 ( R_70_f7d4000, \65090 );
buf \U$labajz7385 ( R_71_acee958, \65091 );
buf \U$labajz7386 ( R_72_94046c0, \65092 );
buf \U$labajz7387 ( R_73_101ee420, \65093 );
buf \U$labajz7388 ( R_74_102eb268, \65094 );
buf \U$labajz7389 ( R_75_b320c50, \65095 );
buf \U$labajz7390 ( R_76_ad80a90, \65096 );
buf \U$labajz7391 ( R_77_1027fd48, \65097 );
buf \U$labajz7392 ( R_78_f7ce4b8, \65098 );
buf \U$labajz7393 ( R_79_ad77048, \65099 );
buf \U$labajz7394 ( R_7a_102a6ae0, \65100 );
buf \U$labajz7395 ( R_7b_f7e4c78, \65101 );
buf \U$labajz7396 ( R_7c_e2a6ce0, \65102 );
buf \U$labajz7397 ( R_7d_101e86e0, \65103 );
buf \U$labajz7398 ( R_7e_e2a9cc8, \65108 );
buf \U$labajz7399 ( R_7f_10292be0, \65109 );
buf \U$labajz7400 ( R_80_b33cde8, \65110 );
buf \U$labajz7401 ( R_81_101e2908, \65111 );
buf \U$labajz7402 ( R_82_102e9780, \65112 );
buf \U$labajz7403 ( R_83_f8157a0, \65113 );
buf \U$labajz7404 ( R_84_f819358, \65114 );
buf \U$labajz7405 ( R_85_ace8b70, \65115 );
buf \U$labajz7406 ( R_86_be142b0, \65116 );
buf \U$labajz7407 ( R_87_f81b770, \65117 );
buf \U$labajz7408 ( R_88_b330278, \65118 );
buf \U$labajz7409 ( R_89_f7fe9f8, \65119 );
buf \U$labajz7410 ( R_8a_101cf488, \65124 );
buf \U$labajz7411 ( R_8b_f8225c0, \65125 );
buf \U$labajz7412 ( R_8c_101d4738, \65126 );
buf \U$labajz7413 ( R_8d_101c4000, \65127 );
buf \U$labajz7414 ( R_8e_101fe960, \65132 );
buf \U$labajz7415 ( R_8f_102a0330, \65137 );
buf \U$labajz7416 ( R_90_f7f4bd0, \65142 );
buf \U$labajz7417 ( R_91_1023e5a8, \65143 );
buf \U$labajz7418 ( R_92_10248da8, \65148 );
buf \U$labajz7419 ( R_93_be2c938, \65149 );
buf \U$labajz7420 ( R_94_f7f5458, \65154 );
buf \U$labajz7421 ( R_95_f7c6808, \65158 );
buf \U$labajz7422 ( R_96_be316a8, \65197 );
buf \U$labajz7423 ( R_97_e2a0328, \65201 );
buf \U$labajz7424 ( R_98_be2d850, \65163 );
buf \U$labajz7425 ( R_99_10217db0, \65165 );
buf \U$labajz7426 ( R_9a_f7ec340, \65166 );
buf \U$labajz7427 ( R_9b_be23ec0, \65205 );
buf \U$labajz7428 ( R_9c_101d4540, \65167 );
buf \U$labajz7429 ( R_9d_f800828, \65209 );
buf \U$labajz7430 ( R_9e_102970c8, \65168 );
buf \U$labajz7431 ( R_9f_10221de0, \65213 );
buf \U$labajz7432 ( R_a0_ad8d568, \65169 );
buf \U$labajz7433 ( R_a1_be4eb58, \65217 );
buf \U$labajz7434 ( R_a2_f7c5500, \65170 );
buf \U$labajz7435 ( R_a3_ad88f30, \65221 );
buf \U$labajz7436 ( R_a4_f82f088, \65171 );
buf \U$labajz7437 ( R_a5_f7dcbc8, \65225 );
buf \U$labajz7438 ( R_a6_10292940, \65172 );
buf \U$labajz7439 ( R_a7_be138d8, \65174 );
buf \U$labajz7440 ( R_a8_acee418, \65175 );
buf \U$labajz7441 ( R_a9_ad84450, \65177 );
buf \U$labajz7442 ( R_aa_be10838, \65178 );
buf \U$labajz7443 ( R_ab_be31fd8, \65180 );
buf \U$labajz7444 ( R_ac_acdaef0, \65181 );
buf \U$labajz7445 ( R_ad_acea908, \65183 );
buf \U$labajz7446 ( R_ae_101f8830, \65184 );
buf \U$labajz7447 ( R_af_f7dec98, \65186 );
buf \U$labajz7448 ( R_b0_101e2c50, \65187 );
buf \U$labajz7449 ( R_b1_f801b30, \65189 );
buf \U$labajz7450 ( R_b2_be16e00, \65190 );
buf \U$labajz7451 ( R_b3_102e3cf0, \65192 );
buf \U$labajz7452 ( R_b4_10291788, \65193 );
not \g455721/U$2 ( \8311 , RIbc62af0_23);
nor \g455721/U$1 ( \8312 , \8311 , RIbc62a78_22);
buf \g455719/U$1 ( \8313 , \8312 );
not \g455723/U$1 ( \8314 , RIbc62a00_21);
not \g455725/U$1 ( \8315 , RIbc62988_20);
and \g455694/U$1 ( \8316 , \8314 , \8315 );
and \g455554/U$1 ( \8317 , \8313 , \8316 );
not \drc_bufs455883/U$1 ( \8318 , \8317 );
not \drc_bufs455882/U$1 ( \8319 , \8318 );
and \g449061/U$2 ( \8320 , RIe14a150_2220, \8319 );
not \g455697/U$2 ( \8321 , RIbc62a78_22);
nor \g455697/U$1 ( \8322 , \8321 , RIbc62af0_23);
buf \g455695/U$1 ( \8323 , \8322 );
and \g455545/U$1 ( \8324 , \8323 , \8316 );
not \drc_bufs455818/U$1 ( \8325 , \8324 );
not \drc_bufs455815/U$1 ( \8326 , \8325 );
and \g449061/U$3 ( \8327 , \8326 , RIe14ce50_2252);
nand \g455687/U$1 ( \8328 , RIbc62a00_21, RIbc62988_20);
not \g455685/U$1 ( \8329 , \8328 );
and \g455559/U$1 ( \8330 , \8323 , \8329 );
and \g449061/U$4 ( \8331 , RIe163650_2508, \8330 );
nor \g449061/U$1 ( \8332 , \8320 , \8327 , \8331 );
nor \g455684/U$1 ( \8333 , RIbc62af0_23, RIbc62a78_22);
and \g455478/U$1 ( \8334 , \8316 , \8333 );
buf \g455477/U$1 ( \8335 , \8334 );
and \g452459/U$2 ( \8336 , \8335 , RIe147450_2188);
not \g2/U$2 ( \8337 , \8316 );
nand \g455700/U$1 ( \8338 , RIbc62a78_22, RIbc62af0_23);
nor \g2/U$1 ( \8339 , \8337 , \8338 );
buf \g455431/U$1 ( \8340 , \8339 );
and \g452459/U$3 ( \8341 , RIfc62f30_6148, \8340 );
nor \g452459/U$1 ( \8342 , \8336 , \8341 );
and \g454863/U$2 ( \8343 , \8313 , RIee35638_5066);
and \g454863/U$3 ( \8344 , RIe152850_2316, \8323 );
nor \g454863/U$1 ( \8345 , \8343 , \8344 );
not \g450075/U$3 ( \8346 , \8345 );
or \g455714/U$1 ( \8347 , \8314 , RIbc62988_20);
not \g450075/U$4 ( \8348 , \8347 );
and \g450075/U$2 ( \8349 , \8346 , \8348 );
nor \g455456/U$1 ( \8350 , \8328 , \8338 );
buf \g455455/U$1 ( \8351 , \8350 );
and \g450075/U$5 ( \8352 , \8351 , RIe166350_2540);
nor \g450075/U$1 ( \8353 , \8349 , \8352 );
not \g455467/U$2 ( \8354 , \8333 );
nor \g455467/U$1 ( \8355 , \8354 , \8347 );
buf \g455466/U$1 ( \8356 , \8355 );
and \g452456/U$2 ( \8357 , \8356 , RIe14fb50_2284);
nor \g455438/U$1 ( \8358 , \8347 , \8338 );
buf \g455437/U$1 ( \8359 , \8358 );
and \g452456/U$3 ( \8360 , RIfea3ba8_8207, \8359 );
nor \g452456/U$1 ( \8361 , \8357 , \8360 );
nand \g447758/U$1 ( \8362 , \8332 , \8342 , \8353 , \8361 );
or \g455681/U$1 ( \8363 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
not \g454133/U$2 ( \8364 , \8363 );
nand \g454133/U$1 ( \8365 , \8364 , RIbc62820_17);
not \g450543/U$2 ( \8366 , \8365 );
nand \g450543/U$1 ( \8367 , \8366 , RIbc62910_19);
or \g448476/U$1 ( \8368 , \8367 , RIbc62898_18);
not \g448475/U$1 ( \8369 , \8368 );
and \g444779/U$2 ( \8370 , \8362 , \8369 );
and \g455568/U$1 ( \8371 , \8313 , \8329 );
not \drc_bufs455896/U$1 ( \8372 , \8371 );
not \drc_bufs455893/U$1 ( \8373 , \8372 );
and \g446144/U$2 ( \8374 , RIfc8f558_6653, \8373 );
not \g455422/U$2 ( \8375 , \8333 );
or \g455692/U$1 ( \8376 , \8315 , RIbc62a00_21);
nor \g455422/U$1 ( \8377 , \8375 , \8376 );
buf \g455421/U$1 ( \8378 , \8377 );
and \g446144/U$3 ( \8379 , RIdf3b308_2050, \8378 );
and \g449063/U$2 ( \8380 , RIfea3a40_8206, \8319 );
and \g449063/U$3 ( \8381 , \8324 , RIfea38d8_8205);
not \drc_bufs455779/U$1 ( \8382 , \8330 );
not \drc_bufs455778/U$1 ( \8383 , \8382 );
and \g449063/U$4 ( \8384 , RIfc89888_6587, \8383 );
nor \g449063/U$1 ( \8385 , \8380 , \8381 , \8384 );
and \g452465/U$2 ( \8386 , \8335 , RIdf2ff08_1922);
and \g452465/U$3 ( \8387 , RIdf365b0_1995, \8340 );
nor \g452465/U$1 ( \8388 , \8386 , \8387 );
and \g454866/U$2 ( \8389 , \8313 , RIee2e9f0_4989);
and \g454866/U$3 ( \8390 , RIfc568e8_6007, \8323 );
nor \g454866/U$1 ( \8391 , \8389 , \8390 );
not \g450078/U$3 ( \8392 , \8391 );
not \g450078/U$4 ( \8393 , \8347 );
and \g450078/U$2 ( \8394 , \8392 , \8393 );
and \g450078/U$5 ( \8395 , \8351 , RIfc97f28_6751);
nor \g450078/U$1 ( \8396 , \8394 , \8395 );
and \g452464/U$2 ( \8397 , \8356 , RIee2dbe0_4979);
and \g452464/U$3 ( \8398 , RIee30a48_5012, \8359 );
nor \g452464/U$1 ( \8399 , \8397 , \8398 );
nand \g447759/U$1 ( \8400 , \8385 , \8388 , \8396 , \8399 );
nor \g446144/U$1 ( \8401 , \8374 , \8379 , \8400 );
not \g455449/U$2 ( \8402 , \8333 );
nor \g455449/U$1 ( \8403 , \8402 , \8328 );
buf \g455448/U$1 ( \8404 , \8403 );
and \g452463/U$2 ( \8405 , \8404 , RIfc52838_5961);
not \g455690/U$1 ( \8406 , \8376 );
and \g455669/U$1 ( \8407 , \8323 , \8406 );
not \drc_bufs455909/U$1 ( \8408 , \8407 );
not \drc_bufs455907/U$1 ( \8409 , \8408 );
and \g452463/U$3 ( \8410 , RIe13f890_2100, \8409 );
nor \g452463/U$1 ( \8411 , \8405 , \8410 );
and \g455661/U$1 ( \8412 , \8313 , \8406 );
not \drc_bufs455922/U$1 ( \8413 , \8412 );
not \drc_bufs455921/U$1 ( \8414 , \8413 );
and \g452462/U$2 ( \8415 , \8414 , RIdf3d798_2076);
nor \g455488/U$1 ( \8416 , \8376 , \8338 );
buf \g455487/U$1 ( \8417 , \8416 );
and \g452462/U$3 ( \8418 , RIe141bb8_2125, \8417 );
nor \g452462/U$1 ( \8419 , \8415 , \8418 );
and \g445254/U$2 ( \8420 , \8401 , \8411 , \8419 );
or \g450538/U$1 ( \8421 , \8365 , RIbc62910_19);
or \g448464/U$1 ( \8422 , \8421 , RIbc62898_18);
nor \g445254/U$1 ( \8423 , \8420 , \8422 );
nor \g444779/U$1 ( \8424 , \8370 , \8423 );
not \g455440/U$1 ( \8425 , \8403 );
nor \g448398/U$1 ( \8426 , \8368 , \8425 );
and \g446916/U$2 ( \8427 , \8426 , RIe160950_2476);
nor \g448395/U$1 ( \8428 , \8368 , \8372 );
and \g446916/U$3 ( \8429 , RIee37d98_5094, \8428 );
nor \g446916/U$1 ( \8430 , \8427 , \8429 );
nor \g448397/U$1 ( \8431 , \8368 , \8408 );
and \g446915/U$2 ( \8432 , \8431 , RIe15dc50_2444);
not \g455486/U$1 ( \8433 , \8417 );
nor \g448318/U$1 ( \8434 , \8368 , \8433 );
and \g446915/U$3 ( \8435 , RIfcaa678_6961, \8434 );
nor \g446915/U$1 ( \8436 , \8432 , \8435 );
not \g455413/U$1 ( \8437 , \8377 );
nor \g448400/U$1 ( \8438 , \8368 , \8437 );
and \g446917/U$2 ( \8439 , \8438 , RIe155550_2348);
nor \g448399/U$1 ( \8440 , \8368 , \8413 );
and \g446917/U$3 ( \8441 , RIe158250_2380, \8440 );
nor \g446917/U$1 ( \8442 , \8439 , \8441 );
nand \g444503/U$1 ( \8443 , \8424 , \8430 , \8436 , \8442 );
and \g452475/U$2 ( \8444 , \8404 , RIdf0f820_1553);
and \g452475/U$3 ( \8445 , RIdf09e20_1489, \8407 );
nor \g452475/U$1 ( \8446 , \8444 , \8445 );
and \g446146/U$2 ( \8447 , RIdf12520_1585, \8373 );
and \g446146/U$3 ( \8448 , RIdf04420_1425, \8378 );
and \g449067/U$2 ( \8449 , RIdeedc20_1169, \8319 );
and \g449067/U$3 ( \8450 , \8326 , RIdef0920_1201);
and \g449067/U$4 ( \8451 , RIdf15220_1617, \8383 );
nor \g449067/U$1 ( \8452 , \8449 , \8450 , \8451 );
and \g452478/U$2 ( \8453 , \8335 , RIdeeaf20_1137);
and \g452478/U$3 ( \8454 , RIdef3620_1233, \8340 );
nor \g452478/U$1 ( \8455 , \8453 , \8454 );
and \g454874/U$2 ( \8456 , \8313 , RIdef9020_1297);
and \g454874/U$3 ( \8457 , RIdefbd20_1329, \8323 );
nor \g454874/U$1 ( \8458 , \8456 , \8457 );
not \g450081/U$3 ( \8459 , \8458 );
not \g450081/U$4 ( \8460 , \8347 );
and \g450081/U$2 ( \8461 , \8459 , \8460 );
and \g450081/U$5 ( \8462 , \8351 , RIdf17f20_1649);
nor \g450081/U$1 ( \8463 , \8461 , \8462 );
and \g452477/U$2 ( \8464 , \8356 , RIdef6320_1265);
and \g452477/U$3 ( \8465 , RIdefea20_1361, \8359 );
nor \g452477/U$1 ( \8466 , \8464 , \8465 );
nand \g447762/U$1 ( \8467 , \8452 , \8455 , \8463 , \8466 );
nor \g446146/U$1 ( \8468 , \8447 , \8448 , \8467 );
and \g452473/U$2 ( \8469 , \8412 , RIdf07120_1457);
and \g452473/U$3 ( \8470 , RIdf0cb20_1521, \8417 );
nor \g452473/U$1 ( \8471 , \8469 , \8470 );
nand \g445611/U$1 ( \8472 , \8446 , \8468 , \8471 );
not \g450537/U$2 ( \8473 , RIbc62910_19);
nor \g454135/U$1 ( \8474 , \8363 , RIbc62820_17);
nand \g450537/U$1 ( \8475 , \8473 , \8474 );
not \g455722/U$1 ( \8476 , RIbc62898_18);
or \g448474/U$1 ( \8477 , \8475 , \8476 );
not \g448473/U$1 ( \8478 , \8477 );
and \g444780/U$2 ( \8479 , \8472 , \8478 );
nand \g450542/U$1 ( \8480 , RIbc62910_19, \8474 );
or \g448468/U$1 ( \8481 , \8480 , RIbc62898_18);
not \g448467/U$1 ( \8482 , \8481 );
and \g449065/U$2 ( \8483 , RIdee15d8_1028, \8412 );
and \g449065/U$3 ( \8484 , \8409 , RIdee3798_1052);
not \g455712/U$1 ( \8485 , \8347 );
and \g455652/U$1 ( \8486 , \8323 , \8485 );
not \drc_bufs455740/U$1 ( \8487 , \8486 );
not \drc_bufs455738/U$1 ( \8488 , \8487 );
and \g449065/U$4 ( \8489 , RIfc72ae8_6327, \8488 );
nor \g449065/U$1 ( \8490 , \8483 , \8484 , \8489 );
and \g454234/U$2 ( \8491 , \8313 , RIfc5beb0_6068);
and \g454234/U$3 ( \8492 , RIfc7c598_6437, \8323 );
nor \g454234/U$1 ( \8493 , \8491 , \8492 );
not \g450079/U$3 ( \8494 , \8493 );
not \g450079/U$4 ( \8495 , \8328 );
and \g450079/U$2 ( \8496 , \8494 , \8495 );
and \g450079/U$5 ( \8497 , \8359 , RIfcb3048_7059);
nor \g450079/U$1 ( \8498 , \8496 , \8497 );
and \g452467/U$2 ( \8499 , \8404 , RIfc58ee0_6034);
and \g452467/U$3 ( \8500 , RIfcab8c0_6974, \8351 );
nor \g452467/U$1 ( \8501 , \8499 , \8500 );
and \g452469/U$2 ( \8502 , \8378 , RIdedf580_1005);
and \g452469/U$3 ( \8503 , RIdee5688_1074, \8417 );
nor \g452469/U$1 ( \8504 , \8502 , \8503 );
nand \g447761/U$1 ( \8505 , \8490 , \8498 , \8501 , \8504 );
and \g444780/U$3 ( \8506 , \8482 , \8505 );
nor \g444780/U$1 ( \8507 , \8479 , \8506 );
not \g455469/U$1 ( \8508 , \8334 );
nor \g448290/U$1 ( \8509 , \8481 , \8508 );
and \g446923/U$2 ( \8510 , \8509 , RIded3a78_872);
nor \g448289/U$1 ( \8511 , \8481 , \8318 );
and \g446923/U$3 ( \8512 , RIfea3068_8199, \8511 );
nor \g446923/U$1 ( \8513 , \8510 , \8512 );
nor \g448288/U$1 ( \8514 , \8481 , \8325 );
and \g446922/U$2 ( \8515 , \8514 , RIded7f60_921);
not \g455425/U$1 ( \8516 , \8339 );
nor \g448260/U$1 ( \8517 , \8481 , \8516 );
and \g446922/U$3 ( \8518 , RIdeda558_948, \8517 );
nor \g446922/U$1 ( \8519 , \8515 , \8518 );
not \g455458/U$1 ( \8520 , \8355 );
nor \g448305/U$1 ( \8521 , \8481 , \8520 );
and \g446924/U$2 ( \8522 , \8521 , RIfcb6450_7096);
and \g455645/U$1 ( \8523 , \8313 , \8485 );
not \drc_bufs455857/U$1 ( \8524 , \8523 );
nor \g448306/U$1 ( \8525 , \8481 , \8524 );
and \g446924/U$3 ( \8526 , RIfca3d00_6886, \8525 );
nor \g446924/U$1 ( \8527 , \8522 , \8526 );
nand \g444504/U$1 ( \8528 , \8507 , \8513 , \8519 , \8527 );
and \g446139/U$2 ( \8529 , RIfcc6440_7278, \8373 );
and \g446139/U$3 ( \8530 , RIfea3338_8201, \8378 );
not \drc_bufs455855/U$1 ( \8531 , \8524 );
and \g449056/U$2 ( \8532 , RIfc9dd60_6818, \8531 );
and \g449056/U$3 ( \8533 , \8488 , RIfcb6888_7099);
and \g449056/U$4 ( \8534 , RIfcda648_7507, \8330 );
nor \g449056/U$1 ( \8535 , \8532 , \8533 , \8534 );
and \g452444/U$2 ( \8536 , \8335 , RIfec62e8_8375);
and \g452444/U$3 ( \8537 , RIfc50c18_5941, \8340 );
nor \g452444/U$1 ( \8538 , \8536 , \8537 );
and \g454263/U$2 ( \8539 , \8313 , RIfc80a80_6486);
and \g454263/U$3 ( \8540 , RIe16c458_2609, \8323 );
nor \g454263/U$1 ( \8541 , \8539 , \8540 );
not \g454262/U$1 ( \8542 , \8541 );
and \g450071/U$2 ( \8543 , \8542 , \8316 );
and \g450071/U$3 ( \8544 , RIee1d4e8_4792, \8351 );
nor \g450071/U$1 ( \8545 , \8543 , \8544 );
and \g452443/U$2 ( \8546 , \8356 , RIee19708_4748);
and \g452443/U$3 ( \8547 , RIfcb6b58_7101, \8359 );
nor \g452443/U$1 ( \8548 , \8546 , \8547 );
nand \g448201/U$1 ( \8549 , \8535 , \8538 , \8545 , \8548 );
nor \g446139/U$1 ( \8550 , \8529 , \8530 , \8549 );
and \g452442/U$2 ( \8551 , \8404 , RIfcd5620_7450);
and \g452442/U$3 ( \8552 , RIfea34a0_8202, \8409 );
nor \g452442/U$1 ( \8553 , \8551 , \8552 );
and \g452440/U$2 ( \8554 , \8414 , RIfea31d0_8200);
and \g452440/U$3 ( \8555 , RIde92ac8_305, \8417 );
nor \g452440/U$1 ( \8556 , \8554 , \8555 );
and \g445250/U$2 ( \8557 , \8550 , \8553 , \8556 );
or \g448466/U$1 ( \8558 , \8421 , \8476 );
nor \g445250/U$1 ( \8559 , \8557 , \8558 );
and \g446141/U$2 ( \8560 , RIfcaf3d0_7016, \8373 );
and \g446141/U$3 ( \8561 , RIdebaf50_591, \8414 );
and \g449059/U$2 ( \8562 , RIdea5f38_399, \8319 );
and \g449059/U$3 ( \8563 , \8326 , RIdeac838_431);
and \g449059/U$4 ( \8564 , RIdec3650_687, \8383 );
nor \g449059/U$1 ( \8565 , \8562 , \8563 , \8564 );
and \g452453/U$2 ( \8566 , \8335 , RIde9f638_367);
and \g452453/U$3 ( \8567 , RIfc8c6f0_6620, \8340 );
nor \g452453/U$1 ( \8568 , \8566 , \8567 );
and \g454256/U$2 ( \8569 , \8313 , RIfc981f8_6753);
and \g454256/U$3 ( \8570 , RIdeb2850_495, \8323 );
nor \g454256/U$1 ( \8571 , \8569 , \8570 );
not \g450073/U$3 ( \8572 , \8571 );
not \g450073/U$4 ( \8573 , \8347 );
and \g450073/U$2 ( \8574 , \8572 , \8573 );
and \g450073/U$5 ( \8575 , \8351 , RIdec6350_719);
nor \g450073/U$1 ( \8576 , \8574 , \8575 );
and \g452451/U$2 ( \8577 , \8356 , RIdeafb50_463);
and \g452451/U$3 ( \8578 , RIfc42f50_5784, \8359 );
nor \g452451/U$1 ( \8579 , \8577 , \8578 );
nand \g447756/U$1 ( \8580 , \8565 , \8568 , \8576 , \8579 );
nor \g446141/U$1 ( \8581 , \8560 , \8561 , \8580 );
and \g452449/U$2 ( \8582 , \8404 , RIdec0950_655);
and \g452449/U$3 ( \8583 , RIfc6a280_6230, \8417 );
nor \g452449/U$1 ( \8584 , \8582 , \8583 );
and \g452450/U$2 ( \8585 , \8378 , RIdeb8250_559);
and \g452450/U$3 ( \8586 , RIdebdc50_623, \8407 );
nor \g452450/U$1 ( \8587 , \8585 , \8586 );
and \g445252/U$2 ( \8588 , \8581 , \8584 , \8587 );
or \g448482/U$1 ( \8589 , \8367 , \8476 );
nor \g445252/U$1 ( \8590 , \8588 , \8589 );
or \g444399/U$1 ( \8591 , \8443 , \8528 , \8559 , \8590 );
and \g446137/U$2 ( \8592 , RIfca50b0_6900, \8531 );
and \g446137/U$3 ( \8593 , RIfc73628_6335, \8319 );
and \g449053/U$2 ( \8594 , RIee29590_4929, \8373 );
and \g449053/U$3 ( \8595 , \8383 , RIee2ac10_4945);
and \g449053/U$4 ( \8596 , RIfc75c20_6362, \8488 );
nor \g449053/U$1 ( \8597 , \8594 , \8595 , \8596 );
and \g454853/U$2 ( \8598 , \8313 , RIfea3608_8203);
and \g454853/U$3 ( \8599 , RIdf28e88_1842, \8323 );
nor \g454853/U$1 ( \8600 , \8598 , \8599 );
not \g450067/U$3 ( \8601 , \8600 );
not \g450067/U$4 ( \8602 , \8376 );
and \g450067/U$2 ( \8603 , \8601 , \8602 );
and \g450067/U$5 ( \8604 , \8359 , RIfcc0d10_7216);
nor \g450067/U$1 ( \8605 , \8603 , \8604 );
and \g452427/U$2 ( \8606 , \8404 , RIee28348_4916);
and \g452427/U$3 ( \8607 , RIee2c6c8_4964, \8351 );
nor \g452427/U$1 ( \8608 , \8606 , \8607 );
and \g452429/U$2 ( \8609 , \8378 , RIfea3770_8204);
and \g452429/U$3 ( \8610 , RIdf2ad78_1864, \8417 );
nor \g452429/U$1 ( \8611 , \8609 , \8610 );
nand \g447753/U$1 ( \8612 , \8597 , \8605 , \8608 , \8611 );
nor \g446137/U$1 ( \8613 , \8592 , \8593 , \8612 );
and \g452425/U$2 ( \8614 , \8335 , RIdf1a0e0_1673);
and \g452425/U$3 ( \8615 , RIfcc9410_7312, \8340 );
nor \g452425/U$1 ( \8616 , \8614 , \8615 );
and \g452424/U$2 ( \8617 , \8326 , RIdf20620_1745);
and \g452424/U$3 ( \8618 , RIfc74e10_6352, \8356 );
nor \g452424/U$1 ( \8619 , \8617 , \8618 );
and \g445247/U$2 ( \8620 , \8613 , \8616 , \8619 );
or \g448470/U$1 ( \8621 , \8480 , \8476 );
nor \g445247/U$1 ( \8622 , \8620 , \8621 );
and \g446138/U$2 ( \8623 , RIdeb5550_527, \8417 );
and \g446138/U$3 ( \8624 , RIdec9050_751, \8404 );
and \g449055/U$2 ( \8625 , RIdf2d7a8_1894, \8531 );
and \g449055/U$3 ( \8626 , \8488 , RIdf39148_2026);
and \g449055/U$4 ( \8627 , RIdecea50_815, \8383 );
nor \g449055/U$1 ( \8628 , \8625 , \8626 , \8627 );
and \g452437/U$2 ( \8629 , \8335 , RIde7ec80_208);
and \g452437/U$3 ( \8630 , RIdf01720_1393, \8340 );
nor \g452437/U$1 ( \8631 , \8629 , \8630 );
and \g454858/U$2 ( \8632 , \8313 , RIdedcf88_978);
and \g454858/U$3 ( \8633 , RIdee8220_1105, \8323 );
nor \g454858/U$1 ( \8634 , \8632 , \8633 );
not \g454857/U$1 ( \8635 , \8634 );
and \g450070/U$2 ( \8636 , \8635 , \8316 );
and \g450070/U$3 ( \8637 , RIded1750_847, \8351 );
nor \g450070/U$1 ( \8638 , \8636 , \8637 );
and \g452436/U$2 ( \8639 , \8356 , RIdf1e028_1718);
and \g452436/U$3 ( \8640 , RIe144750_2156, \8359 );
nor \g452436/U$1 ( \8641 , \8639 , \8640 );
nand \g448200/U$1 ( \8642 , \8628 , \8631 , \8638 , \8641 );
nor \g446138/U$1 ( \8643 , \8623 , \8624 , \8642 );
and \g452434/U$2 ( \8644 , \8378 , RIe15af50_2412);
and \g452434/U$3 ( \8645 , RIdecbd50_783, \8373 );
nor \g452434/U$1 ( \8646 , \8644 , \8645 );
and \g452433/U$2 ( \8647 , \8414 , RIe16f158_2641);
and \g452433/U$3 ( \8648 , RIde98d38_335, \8409 );
nor \g452433/U$1 ( \8649 , \8647 , \8648 );
and \g445248/U$2 ( \8650 , \8643 , \8646 , \8649 );
or \g448488/U$1 ( \8651 , \8475 , RIbc62898_18);
nor \g445248/U$1 ( \8652 , \8650 , \8651 );
or \g444191/U$1 ( \8653 , \8591 , \8622 , \8652 );
buf \g455927/U$1 ( \8654 , \8363 );
_DC \g2235/U$1 ( \8655 , \8653 , \8654 );
and \g449093/U$2 ( \8656 , RIe1580e8_2379, \8414 );
and \g449093/U$3 ( \8657 , \8409 , RIe15dae8_2443);
and \g449093/U$4 ( \8658 , RIe1526e8_2315, \8488 );
nor \g449093/U$1 ( \8659 , \8656 , \8657 , \8658 );
and \g454909/U$2 ( \8660 , \8313 , RIee37c30_5093);
and \g454909/U$3 ( \8661 , RIe1634e8_2507, \8323 );
nor \g454909/U$1 ( \8662 , \8660 , \8661 );
not \g450108/U$3 ( \8663 , \8662 );
not \g450108/U$4 ( \8664 , \8328 );
and \g450108/U$2 ( \8665 , \8663 , \8664 );
and \g450108/U$5 ( \8666 , \8359 , RIfc3f698_5747);
nor \g450108/U$1 ( \8667 , \8665 , \8666 );
and \g452571/U$2 ( \8668 , \8404 , RIe1607e8_2475);
and \g452571/U$3 ( \8669 , RIe1661e8_2539, \8351 );
nor \g452571/U$1 ( \8670 , \8668 , \8669 );
and \g452574/U$2 ( \8671 , \8378 , RIe1553e8_2347);
and \g452574/U$3 ( \8672 , RIfce7500_7654, \8417 );
nor \g452574/U$1 ( \8673 , \8671 , \8672 );
nand \g447777/U$1 ( \8674 , \8659 , \8667 , \8670 , \8673 );
and \g444782/U$2 ( \8675 , \8674 , \8369 );
and \g446169/U$2 ( \8676 , RIfc88a78_6577, \8531 );
and \g446169/U$3 ( \8677 , RIdf31df8_1944, \8319 );
and \g449095/U$2 ( \8678 , RIfc695d8_6221, \8373 );
and \g449095/U$3 ( \8679 , \8330 , RIfcb7ad0_7112);
and \g449095/U$4 ( \8680 , RIee2fda0_5003, \8488 );
nor \g449095/U$1 ( \8681 , \8678 , \8679 , \8680 );
and \g454146/U$2 ( \8682 , \8313 , RIdf3d630_2075);
and \g454146/U$3 ( \8683 , RIe13f728_2099, \8323 );
nor \g454146/U$1 ( \8684 , \8682 , \8683 );
not \g450111/U$3 ( \8685 , \8684 );
not \g450111/U$4 ( \8686 , \8376 );
and \g450111/U$2 ( \8687 , \8685 , \8686 );
and \g450111/U$5 ( \8688 , \8359 , RIfca9e08_6955);
nor \g450111/U$1 ( \8689 , \8687 , \8688 );
and \g452580/U$2 ( \8690 , \8404 , RIfc51a28_5951);
and \g452580/U$3 ( \8691 , RIfcea4d0_7688, \8351 );
nor \g452580/U$1 ( \8692 , \8690 , \8691 );
and \g452581/U$2 ( \8693 , \8378 , RIdf3b1a0_2049);
and \g452581/U$3 ( \8694 , RIe141a50_2124, \8417 );
nor \g452581/U$1 ( \8695 , \8693 , \8694 );
nand \g447778/U$1 ( \8696 , \8681 , \8689 , \8692 , \8695 );
nor \g446169/U$1 ( \8697 , \8676 , \8677 , \8696 );
and \g452579/U$2 ( \8698 , \8335 , RIfea2258_8189);
and \g452579/U$3 ( \8699 , RIdf36448_1994, \8340 );
nor \g452579/U$1 ( \8700 , \8698 , \8699 );
and \g452578/U$2 ( \8701 , \8326 , RIdf33fb8_1968);
and \g452578/U$3 ( \8702 , RIee2da78_4978, \8356 );
nor \g452578/U$1 ( \8703 , \8701 , \8702 );
and \g445271/U$2 ( \8704 , \8697 , \8700 , \8703 );
nor \g445271/U$1 ( \8705 , \8704 , \8422 );
nor \g444782/U$1 ( \8706 , \8675 , \8705 );
nor \g448404/U$1 ( \8707 , \8368 , \8508 );
and \g446943/U$2 ( \8708 , \8707 , RIe1472e8_2187);
nor \g448403/U$1 ( \8709 , \8368 , \8318 );
and \g446943/U$3 ( \8710 , RIe149fe8_2219, \8709 );
nor \g446943/U$1 ( \8711 , \8708 , \8710 );
nor \g448402/U$1 ( \8712 , \8368 , \8325 );
and \g446942/U$2 ( \8713 , \8712 , RIe14cce8_2251);
nor \g448319/U$1 ( \8714 , \8368 , \8516 );
and \g446942/U$3 ( \8715 , RIfc83e88_6523, \8714 );
nor \g446942/U$1 ( \8716 , \8713 , \8715 );
nor \g448406/U$1 ( \8717 , \8368 , \8520 );
and \g446944/U$2 ( \8718 , \8717 , RIe14f9e8_2283);
nor \g448405/U$1 ( \8719 , \8368 , \8524 );
and \g446944/U$3 ( \8720 , RIee354d0_5065, \8719 );
nor \g446944/U$1 ( \8721 , \8718 , \8720 );
nand \g444507/U$1 ( \8722 , \8706 , \8711 , \8716 , \8721 );
and \g452592/U$2 ( \8723 , \8404 , RIee281e0_4915);
and \g452592/U$3 ( \8724 , RIdf28d20_1841, \8409 );
nor \g452592/U$1 ( \8725 , \8723 , \8724 );
and \g446170/U$2 ( \8726 , RIee29428_4928, \8373 );
and \g446170/U$3 ( \8727 , RIfea2960_8194, \8378 );
and \g449099/U$2 ( \8728 , RIfc99cb0_6772, \8319 );
and \g449099/U$3 ( \8729 , \8324 , RIdf204b8_1744);
and \g449099/U$4 ( \8730 , RIee2aaa8_4944, \8383 );
nor \g449099/U$1 ( \8731 , \8728 , \8729 , \8730 );
and \g452596/U$2 ( \8732 , \8335 , RIdf19f78_1672);
and \g452596/U$3 ( \8733 , RIfca0a60_6850, \8340 );
nor \g452596/U$1 ( \8734 , \8732 , \8733 );
and \g454921/U$2 ( \8735 , \8313 , RIfc8b1d8_6605);
and \g454921/U$3 ( \8736 , RIfca08f8_6849, \8323 );
nor \g454921/U$1 ( \8737 , \8735 , \8736 );
not \g450114/U$3 ( \8738 , \8737 );
not \g450114/U$4 ( \8739 , \8347 );
and \g450114/U$2 ( \8740 , \8738 , \8739 );
and \g450114/U$5 ( \8741 , \8351 , RIee2c560_4963);
nor \g450114/U$1 ( \8742 , \8740 , \8741 );
and \g452594/U$2 ( \8743 , \8356 , RIfc49058_5853);
and \g452594/U$3 ( \8744 , RIfcdabe8_7511, \8359 );
nor \g452594/U$1 ( \8745 , \8743 , \8744 );
nand \g447781/U$1 ( \8746 , \8731 , \8734 , \8742 , \8745 );
nor \g446170/U$1 ( \8747 , \8726 , \8727 , \8746 );
and \g452591/U$2 ( \8748 , \8414 , RIfea27f8_8193);
and \g452591/U$3 ( \8749 , RIdf2ac10_1863, \8417 );
nor \g452591/U$1 ( \8750 , \8748 , \8749 );
nand \g445616/U$1 ( \8751 , \8725 , \8747 , \8750 );
not \g448469/U$1 ( \8752 , \8621 );
and \g444725/U$2 ( \8753 , \8751 , \8752 );
and \g449097/U$2 ( \8754 , RIdf06fb8_1456, \8412 );
and \g449097/U$3 ( \8755 , \8409 , RIdf09cb8_1488);
and \g449097/U$4 ( \8756 , RIdefbbb8_1328, \8488 );
nor \g449097/U$1 ( \8757 , \8754 , \8755 , \8756 );
and \g454917/U$2 ( \8758 , \8313 , RIdf123b8_1584);
and \g454917/U$3 ( \8759 , RIdf150b8_1616, \8323 );
nor \g454917/U$1 ( \8760 , \8758 , \8759 );
not \g450112/U$3 ( \8761 , \8760 );
not \g450112/U$4 ( \8762 , \8328 );
and \g450112/U$2 ( \8763 , \8761 , \8762 );
and \g450112/U$5 ( \8764 , \8359 , RIdefe8b8_1360);
nor \g450112/U$1 ( \8765 , \8763 , \8764 );
and \g452584/U$2 ( \8766 , \8404 , RIdf0f6b8_1552);
and \g452584/U$3 ( \8767 , RIdf17db8_1648, \8351 );
nor \g452584/U$1 ( \8768 , \8766 , \8767 );
and \g452585/U$2 ( \8769 , \8378 , RIdf042b8_1424);
and \g452585/U$3 ( \8770 , RIdf0c9b8_1520, \8417 );
nor \g452585/U$1 ( \8771 , \8769 , \8770 );
nand \g447779/U$1 ( \8772 , \8757 , \8765 , \8768 , \8771 );
and \g444725/U$3 ( \8773 , \8478 , \8772 );
nor \g444725/U$1 ( \8774 , \8753 , \8773 );
nor \g448309/U$1 ( \8775 , \8477 , \8520 );
and \g446946/U$2 ( \8776 , \8775 , RIdef61b8_1264);
nor \g448351/U$1 ( \8777 , \8477 , \8524 );
and \g446946/U$3 ( \8778 , RIdef8eb8_1296, \8777 );
nor \g446946/U$1 ( \8779 , \8776 , \8778 );
nor \g448340/U$1 ( \8780 , \8477 , \8325 );
and \g446947/U$2 ( \8781 , \8780 , RIdef07b8_1200);
nor \g448352/U$1 ( \8782 , \8477 , \8516 );
and \g446947/U$3 ( \8783 , RIdef34b8_1232, \8782 );
nor \g446947/U$1 ( \8784 , \8781 , \8783 );
nor \g448311/U$1 ( \8785 , \8477 , \8508 );
and \g446949/U$2 ( \8786 , \8785 , RIdeeadb8_1136);
nor \g448338/U$1 ( \8787 , \8477 , \8318 );
and \g446949/U$3 ( \8788 , RIdeedab8_1168, \8787 );
nor \g446949/U$1 ( \8789 , \8786 , \8788 );
nand \g444624/U$1 ( \8790 , \8774 , \8779 , \8784 , \8789 );
and \g446164/U$2 ( \8791 , RIfc87830_6564, \8531 );
and \g446164/U$3 ( \8792 , RIdea5bf0_398, \8319 );
and \g449089/U$2 ( \8793 , RIee20620_4827, \8371 );
and \g449089/U$3 ( \8794 , \8330 , RIdec34e8_686);
and \g449089/U$4 ( \8795 , RIdeb26e8_494, \8488 );
nor \g449089/U$1 ( \8796 , \8793 , \8794 , \8795 );
and \g454903/U$2 ( \8797 , \8313 , RIdebade8_590);
and \g454903/U$3 ( \8798 , RIdebdae8_622, \8323 );
nor \g454903/U$1 ( \8799 , \8797 , \8798 );
not \g450104/U$3 ( \8800 , \8799 );
not \g450104/U$4 ( \8801 , \8376 );
and \g450104/U$2 ( \8802 , \8800 , \8801 );
and \g450104/U$5 ( \8803 , \8359 , RIfc41150_5766);
nor \g450104/U$1 ( \8804 , \8802 , \8803 );
and \g452559/U$2 ( \8805 , \8404 , RIdec07e8_654);
and \g452559/U$3 ( \8806 , RIdec61e8_718, \8351 );
nor \g452559/U$1 ( \8807 , \8805 , \8806 );
and \g452561/U$2 ( \8808 , \8378 , RIdeb80e8_558);
and \g452561/U$3 ( \8809 , RIfc4b7b8_5881, \8417 );
nor \g452561/U$1 ( \8810 , \8808 , \8809 );
nand \g447774/U$1 ( \8811 , \8796 , \8804 , \8807 , \8810 );
nor \g446164/U$1 ( \8812 , \8791 , \8792 , \8811 );
and \g452558/U$2 ( \8813 , \8335 , RIde9f2f0_366);
and \g452558/U$3 ( \8814 , RIee1dec0_4799, \8340 );
nor \g452558/U$1 ( \8815 , \8813 , \8814 );
and \g452557/U$2 ( \8816 , \8326 , RIdeac4f0_430);
and \g452557/U$3 ( \8817 , RIdeaf9e8_462, \8356 );
nor \g452557/U$1 ( \8818 , \8816 , \8817 );
and \g445266/U$2 ( \8819 , \8812 , \8815 , \8818 );
nor \g445266/U$1 ( \8820 , \8819 , \8589 );
and \g446166/U$2 ( \8821 , RIfc84f68_6535, \8373 );
and \g446166/U$3 ( \8822 , RIde86c78_247, \8378 );
and \g449091/U$2 ( \8823 , RIee388d8_5102, \8319 );
and \g449091/U$3 ( \8824 , \8326 , RIe16c2f0_2608);
and \g449091/U$4 ( \8825 , RIfc77c78_6385, \8330 );
nor \g449091/U$1 ( \8826 , \8823 , \8824 , \8825 );
and \g452566/U$2 ( \8827 , \8335 , RIfea20f0_8188);
and \g452566/U$3 ( \8828 , RIfc76328_6367, \8340 );
nor \g452566/U$1 ( \8829 , \8827 , \8828 );
and \g454161/U$2 ( \8830 , \8313 , RIfcd7240_7470);
and \g454161/U$3 ( \8831 , RIee19f78_4754, \8323 );
nor \g454161/U$1 ( \8832 , \8830 , \8831 );
not \g450106/U$3 ( \8833 , \8832 );
not \g450106/U$4 ( \8834 , \8347 );
and \g450106/U$2 ( \8835 , \8833 , \8834 );
and \g450106/U$5 ( \8836 , \8351 , RIee1d380_4791);
nor \g450106/U$1 ( \8837 , \8835 , \8836 );
and \g452565/U$2 ( \8838 , \8356 , RIfcbeb50_7192);
and \g452565/U$3 ( \8839 , RIee1a680_4759, \8359 );
nor \g452565/U$1 ( \8840 , \8838 , \8839 );
nand \g447775/U$1 ( \8841 , \8826 , \8829 , \8837 , \8840 );
nor \g446166/U$1 ( \8842 , \8821 , \8822 , \8841 );
and \g452564/U$2 ( \8843 , \8404 , RIfc6ff50_6296);
and \g452564/U$3 ( \8844 , RIde8efb8_287, \8409 );
nor \g452564/U$1 ( \8845 , \8843 , \8844 );
and \g452563/U$2 ( \8846 , \8414 , RIde8ae18_267);
and \g452563/U$3 ( \8847 , RIde92780_304, \8417 );
nor \g452563/U$1 ( \8848 , \8846 , \8847 );
and \g445268/U$2 ( \8849 , \8842 , \8845 , \8848 );
nor \g445268/U$1 ( \8850 , \8849 , \8558 );
or \g444401/U$1 ( \8851 , \8722 , \8790 , \8820 , \8850 );
and \g446161/U$2 ( \8852 , RIfcbd7a0_7178, \8531 );
and \g446161/U$3 ( \8853 , RIded3910_871, \8335 );
and \g449084/U$2 ( \8854 , RIfcbe2e0_7186, \8373 );
and \g449084/U$3 ( \8855 , \8383 , RIfc57f68_6023);
and \g449084/U$4 ( \8856 , RIfcb35e8_7063, \8488 );
nor \g449084/U$1 ( \8857 , \8854 , \8855 , \8856 );
and \g454899/U$2 ( \8858 , \8313 , RIdee1470_1027);
and \g454899/U$3 ( \8859 , RIfea2690_8192, \8323 );
nor \g454899/U$1 ( \8860 , \8858 , \8859 );
not \g450099/U$3 ( \8861 , \8860 );
not \g450099/U$4 ( \8862 , \8376 );
and \g450099/U$2 ( \8863 , \8861 , \8862 );
and \g450099/U$5 ( \8864 , \8359 , RIfc57b30_6020);
nor \g450099/U$1 ( \8865 , \8863 , \8864 );
and \g452543/U$2 ( \8866 , \8404 , RIfcd8fc8_7491);
and \g452543/U$3 ( \8867 , RIfcd1f48_7411, \8351 );
nor \g452543/U$1 ( \8868 , \8866 , \8867 );
and \g452546/U$2 ( \8869 , \8378 , RIdedf418_1004);
and \g452546/U$3 ( \8870 , RIdee5520_1073, \8417 );
nor \g452546/U$1 ( \8871 , \8869 , \8870 );
nand \g447771/U$1 ( \8872 , \8857 , \8865 , \8868 , \8871 );
nor \g446161/U$1 ( \8873 , \8852 , \8853 , \8872 );
and \g452541/U$2 ( \8874 , \8356 , RIfc91178_6673);
and \g452541/U$3 ( \8875 , RIfea2528_8191, \8340 );
nor \g452541/U$1 ( \8876 , \8874 , \8875 );
and \g452542/U$2 ( \8877 , \8319 , RIfea23c0_8190);
and \g452542/U$3 ( \8878 , RIded7df8_920, \8326 );
nor \g452542/U$1 ( \8879 , \8877 , \8878 );
and \g445264/U$2 ( \8880 , \8873 , \8876 , \8879 );
nor \g445264/U$1 ( \8881 , \8880 , \8481 );
and \g446163/U$2 ( \8882 , RIdeb53e8_526, \8417 );
and \g446163/U$3 ( \8883 , RIdec8ee8_750, \8404 );
and \g449086/U$2 ( \8884 , RIdedce20_977, \8319 );
and \g449086/U$3 ( \8885 , \8324 , RIdee80b8_1104);
and \g449086/U$4 ( \8886 , RIdece8e8_814, \8383 );
nor \g449086/U$1 ( \8887 , \8884 , \8885 , \8886 );
and \g452554/U$2 ( \8888 , \8335 , RIde7e938_207);
and \g452554/U$3 ( \8889 , RIdf015b8_1392, \8340 );
nor \g452554/U$1 ( \8890 , \8888 , \8889 );
and \g454173/U$2 ( \8891 , \8313 , RIdf2d640_1893);
and \g454173/U$3 ( \8892 , RIdf38fe0_2025, \8323 );
nor \g454173/U$1 ( \8893 , \8891 , \8892 );
not \g450102/U$3 ( \8894 , \8893 );
not \g450102/U$4 ( \8895 , \8347 );
and \g450102/U$2 ( \8896 , \8894 , \8895 );
and \g450102/U$5 ( \8897 , \8351 , RIded15e8_846);
nor \g450102/U$1 ( \8898 , \8896 , \8897 );
and \g452553/U$2 ( \8899 , \8356 , RIdf1dec0_1717);
and \g452553/U$3 ( \8900 , RIe1445e8_2155, \8359 );
nor \g452553/U$1 ( \8901 , \8899 , \8900 );
nand \g447772/U$1 ( \8902 , \8887 , \8890 , \8898 , \8901 );
nor \g446163/U$1 ( \8903 , \8882 , \8883 , \8902 );
and \g452552/U$2 ( \8904 , \8378 , RIe15ade8_2411);
and \g452552/U$3 ( \8905 , RIdecbbe8_782, \8373 );
nor \g452552/U$1 ( \8906 , \8904 , \8905 );
and \g452551/U$2 ( \8907 , \8414 , RIe16eff0_2640);
and \g452551/U$3 ( \8908 , RIde989f0_334, \8407 );
nor \g452551/U$1 ( \8909 , \8907 , \8908 );
and \g445265/U$2 ( \8910 , \8903 , \8906 , \8909 );
nor \g445265/U$1 ( \8911 , \8910 , \8651 );
or \g444171/U$1 ( \8912 , \8851 , \8881 , \8911 );
_DC \g22ba/U$1 ( \8913 , \8912 , \8654 );
and \g451668/U$2 ( \8914 , \8378 , RIdf03fe8_1422);
and \g451668/U$3 ( \8915 , RIdf099e8_1486, \8409 );
nor \g451668/U$1 ( \8916 , \8914 , \8915 );
and \g445952/U$2 ( \8917 , RIdf120e8_1582, \8373 );
and \g445952/U$3 ( \8918 , RIdf06ce8_1454, \8414 );
and \g448817/U$2 ( \8919 , RIdeed7e8_1166, \8317 );
and \g448817/U$3 ( \8920 , \8326 , RIdef04e8_1198);
and \g448817/U$4 ( \8921 , RIdf14de8_1614, \8383 );
nor \g448817/U$1 ( \8922 , \8919 , \8920 , \8921 );
and \g451674/U$2 ( \8923 , \8335 , RIdeeaae8_1134);
and \g451674/U$3 ( \8924 , RIdef31e8_1230, \8340 );
nor \g451674/U$1 ( \8925 , \8923 , \8924 );
and \g454163/U$2 ( \8926 , \8313 , RIdef8be8_1294);
and \g454163/U$3 ( \8927 , RIdefb8e8_1326, \8323 );
nor \g454163/U$1 ( \8928 , \8926 , \8927 );
not \g449843/U$3 ( \8929 , \8928 );
not \g449843/U$4 ( \8930 , \8347 );
and \g449843/U$2 ( \8931 , \8929 , \8930 );
and \g449843/U$5 ( \8932 , \8351 , RIdf17ae8_1646);
nor \g449843/U$1 ( \8933 , \8931 , \8932 );
and \g451673/U$2 ( \8934 , \8356 , RIdef5ee8_1262);
and \g451673/U$3 ( \8935 , RIdefe5e8_1358, \8359 );
nor \g451673/U$1 ( \8936 , \8934 , \8935 );
nand \g447630/U$1 ( \8937 , \8922 , \8925 , \8933 , \8936 );
nor \g445952/U$1 ( \8938 , \8917 , \8918 , \8937 );
and \g451667/U$2 ( \8939 , \8404 , RIdf0f3e8_1550);
and \g451667/U$3 ( \8940 , RIdf0c6e8_1518, \8417 );
nor \g451667/U$1 ( \8941 , \8939 , \8940 );
nand \g445566/U$1 ( \8942 , \8916 , \8938 , \8941 );
and \g444768/U$2 ( \8943 , \8942 , \8478 );
and \g448813/U$2 ( \8944 , RIfc74870_6348, \8531 );
and \g448813/U$3 ( \8945 , \8488 , RIfc4b0b0_5876);
and \g448813/U$4 ( \8946 , RIfcc54c8_7267, \8330 );
nor \g448813/U$1 ( \8947 , \8944 , \8945 , \8946 );
and \g451661/U$2 ( \8948 , \8335 , RIded3640_869);
and \g451661/U$3 ( \8949 , RIdeda288_946, \8340 );
nor \g451661/U$1 ( \8950 , \8948 , \8949 );
and \g454626/U$2 ( \8951 , \8313 , RIded5da0_897);
and \g454626/U$3 ( \8952 , RIded7c90_919, \8323 );
nor \g454626/U$1 ( \8953 , \8951 , \8952 );
not \g454625/U$1 ( \8954 , \8953 );
and \g449840/U$2 ( \8955 , \8954 , \8316 );
and \g449840/U$3 ( \8956 , RIfc89018_6581, \8351 );
nor \g449840/U$1 ( \8957 , \8955 , \8956 );
and \g452136/U$2 ( \8958 , \8356 , RIfce4968_7623);
and \g452136/U$3 ( \8959 , RIfcae188_7003, \8359 );
nor \g452136/U$1 ( \8960 , \8958 , \8959 );
nand \g448168/U$1 ( \8961 , \8947 , \8950 , \8957 , \8960 );
and \g444768/U$3 ( \8962 , \8482 , \8961 );
nor \g444768/U$1 ( \8963 , \8943 , \8962 );
nor \g448296/U$1 ( \8964 , \8481 , \8408 );
and \g446735/U$2 ( \8965 , \8964 , RIdee34c8_1050);
nor \g448259/U$1 ( \8966 , \8481 , \8433 );
and \g446735/U$3 ( \8967 , RIdee53b8_1072, \8966 );
nor \g446735/U$1 ( \8968 , \8965 , \8967 );
nor \g448297/U$1 ( \8969 , \8481 , \8425 );
and \g446737/U$2 ( \8970 , \8969 , RIfc4b380_5878);
nor \g448274/U$1 ( \8971 , \8481 , \8372 );
and \g446737/U$3 ( \8972 , RIfc89180_6582, \8971 );
nor \g446737/U$1 ( \8973 , \8970 , \8972 );
nor \g448299/U$1 ( \8974 , \8481 , \8437 );
and \g446739/U$2 ( \8975 , \8974 , RIdedf148_1002);
nor \g448298/U$1 ( \8976 , \8481 , \8413 );
and \g446739/U$3 ( \8977 , RIfea3d10_8208, \8976 );
nor \g446739/U$1 ( \8978 , \8975 , \8977 );
nand \g444478/U$1 ( \8979 , \8963 , \8968 , \8973 , \8978 );
and \g451075/U$2 ( \8980 , \8324 , RIdf201e8_1742);
and \g451075/U$3 ( \8981 , RIfc86318_6549, \8356 );
nor \g451075/U$1 ( \8982 , \8980 , \8981 );
and \g445956/U$2 ( \8983 , RIdf23320_1777, \8531 );
and \g445956/U$3 ( \8984 , RIdf1b5f8_1688, \8319 );
and \g448826/U$2 ( \8985 , RIdf26b60_1817, \8412 );
and \g448826/U$3 ( \8986 , \8409 , RIdf28a50_1839);
and \g448826/U$4 ( \8987 , RIfcb9df8_7137, \8488 );
nor \g448826/U$1 ( \8988 , \8985 , \8986 , \8987 );
and \g454645/U$2 ( \8989 , \8313 , RIfc572c0_6014);
and \g454645/U$3 ( \8990 , RIfc4cfa0_5898, \8323 );
nor \g454645/U$1 ( \8991 , \8989 , \8990 );
not \g449853/U$3 ( \8992 , \8991 );
not \g449853/U$4 ( \8993 , \8328 );
and \g449853/U$2 ( \8994 , \8992 , \8993 );
and \g449853/U$5 ( \8995 , \8359 , RIfc9b600_6790);
nor \g449853/U$1 ( \8996 , \8994 , \8995 );
and \g451693/U$2 ( \8997 , \8404 , RIfc4f430_5924);
and \g451693/U$3 ( \8998 , RIee2c3f8_4962, \8351 );
nor \g451693/U$1 ( \8999 , \8997 , \8998 );
and \g451696/U$2 ( \9000 , \8378 , RIdf250a8_1798);
and \g451696/U$3 ( \9001 , RIfea3e78_8209, \8417 );
nor \g451696/U$1 ( \9002 , \9000 , \9001 );
nand \g447633/U$1 ( \9003 , \8988 , \8996 , \8999 , \9002 );
nor \g445956/U$1 ( \9004 , \8983 , \8984 , \9003 );
and \g451689/U$2 ( \9005 , \8335 , RIdf19ca8_1670);
and \g451689/U$3 ( \9006 , RIfeabfd8_8273, \8340 );
nor \g451689/U$1 ( \9007 , \9005 , \9006 );
nand \g445568/U$1 ( \9008 , \8982 , \9004 , \9007 );
and \g444843/U$2 ( \9009 , \9008 , \8752 );
not \g448487/U$1 ( \9010 , \8651 );
and \g448821/U$2 ( \9011 , RIdf2d370_1891, \8531 );
and \g448821/U$3 ( \9012 , \8488 , RIdf38d10_2023);
and \g448821/U$4 ( \9013 , RIdece618_812, \8383 );
nor \g448821/U$1 ( \9014 , \9011 , \9012 , \9013 );
and \g451684/U$2 ( \9015 , \8335 , RIde7e2a8_205);
and \g451684/U$3 ( \9016 , RIdf012e8_1390, \8340 );
nor \g451684/U$1 ( \9017 , \9015 , \9016 );
and \g454369/U$2 ( \9018 , \8313 , RIdedcb50_975);
and \g454369/U$3 ( \9019 , RIdee7de8_1102, \8323 );
nor \g454369/U$1 ( \9020 , \9018 , \9019 );
not \g454368/U$1 ( \9021 , \9020 );
and \g449713/U$2 ( \9022 , \9021 , \8316 );
and \g449713/U$3 ( \9023 , RIded1318_844, \8351 );
nor \g449713/U$1 ( \9024 , \9022 , \9023 );
and \g451683/U$2 ( \9025 , \8356 , RIdf1dbf0_1715);
and \g451683/U$3 ( \9026 , RIe144318_2153, \8359 );
nor \g451683/U$1 ( \9027 , \9025 , \9026 );
nand \g448169/U$1 ( \9028 , \9014 , \9017 , \9024 , \9027 );
and \g444843/U$3 ( \9029 , \9010 , \9028 );
nor \g444843/U$1 ( \9030 , \9009 , \9029 );
nor \g448388/U$1 ( \9031 , \8651 , \8437 );
and \g446745/U$2 ( \9032 , \9031 , RIe15ab18_2409);
nor \g448387/U$1 ( \9033 , \8651 , \8413 );
and \g446745/U$3 ( \9034 , RIe16ed20_2638, \9033 );
nor \g446745/U$1 ( \9035 , \9032 , \9034 );
nor \g448381/U$1 ( \9036 , \8651 , \8408 );
and \g446744/U$2 ( \9037 , \9036 , RIde98360_332);
nor \g448315/U$1 ( \9038 , \8651 , \8433 );
and \g446744/U$3 ( \9039 , RIdeb5118_524, \9038 );
nor \g446744/U$1 ( \9040 , \9037 , \9039 );
nor \g448380/U$1 ( \9041 , \8651 , \8425 );
and \g446746/U$2 ( \9042 , \9041 , RIdec8c18_748);
nor \g448374/U$1 ( \9043 , \8651 , \8372 );
and \g446746/U$3 ( \9044 , RIdecb918_780, \9043 );
nor \g446746/U$1 ( \9045 , \9042 , \9044 );
nand \g444588/U$1 ( \9046 , \9030 , \9035 , \9040 , \9045 );
and \g445941/U$2 ( \9047 , RIfcadd50_7000, \8371 );
and \g445941/U$3 ( \9048 , RIe155118_2345, \8378 );
and \g448804/U$2 ( \9049 , RIe149d18_2217, \8319 );
and \g448804/U$3 ( \9050 , \8326 , RIe14ca18_2249);
and \g448804/U$4 ( \9051 , RIe163218_2505, \8330 );
nor \g448804/U$1 ( \9052 , \9049 , \9050 , \9051 );
and \g451632/U$2 ( \9053 , \8335 , RIe147018_2185);
and \g451632/U$3 ( \9054 , RIfcbda70_7180, \8340 );
nor \g451632/U$1 ( \9055 , \9053 , \9054 );
and \g455151/U$2 ( \9056 , \8313 , RIfc498c8_5859);
and \g455151/U$3 ( \9057 , RIe152418_2313, \8323 );
nor \g455151/U$1 ( \9058 , \9056 , \9057 );
not \g449831/U$3 ( \9059 , \9058 );
not \g449831/U$4 ( \9060 , \8347 );
and \g449831/U$2 ( \9061 , \9059 , \9060 );
and \g449831/U$5 ( \9062 , \8351 , RIe165f18_2537);
nor \g449831/U$1 ( \9063 , \9061 , \9062 );
and \g453088/U$2 ( \9064 , \8356 , RIe14f718_2281);
and \g453088/U$3 ( \9065 , RIfc45548_5811, \8359 );
nor \g453088/U$1 ( \9066 , \9064 , \9065 );
nand \g447627/U$1 ( \9067 , \9052 , \9055 , \9063 , \9066 );
nor \g445941/U$1 ( \9068 , \9047 , \9048 , \9067 );
and \g451626/U$2 ( \9069 , \8404 , RIe160518_2473);
and \g451626/U$3 ( \9070 , RIe15d818_2441, \8407 );
nor \g451626/U$1 ( \9071 , \9069 , \9070 );
and \g451623/U$2 ( \9072 , \8414 , RIe157e18_2377);
and \g451623/U$3 ( \9073 , RIfc55268_5991, \8417 );
nor \g451623/U$1 ( \9074 , \9072 , \9073 );
and \g445107/U$2 ( \9075 , \9068 , \9071 , \9074 );
nor \g445107/U$1 ( \9076 , \9075 , \8368 );
and \g445945/U$2 ( \9077 , RIfcb7260_7106, \8356 );
and \g445945/U$3 ( \9078 , RIfea42b0_8212, \8340 );
and \g448810/U$2 ( \9079 , RIee32668_5032, \8373 );
and \g448810/U$3 ( \9080 , \8330 , RIee33748_5044);
and \g448810/U$4 ( \9081 , RIfc42848_5779, \8488 );
nor \g448810/U$1 ( \9082 , \9079 , \9080 , \9081 );
and \g454274/U$2 ( \9083 , \8313 , RIdf3d360_2073);
and \g454274/U$3 ( \9084 , RIe13f458_2097, \8323 );
nor \g454274/U$1 ( \9085 , \9083 , \9084 );
not \g449836/U$3 ( \9086 , \9085 );
not \g449836/U$4 ( \9087 , \8376 );
and \g449836/U$2 ( \9088 , \9086 , \9087 );
and \g449836/U$5 ( \9089 , \8359 , RIfc526d0_5960);
nor \g449836/U$1 ( \9090 , \9088 , \9089 );
and \g451643/U$2 ( \9091 , \8404 , RIee31588_5020);
and \g451643/U$3 ( \9092 , RIee34828_5056, \8351 );
nor \g451643/U$1 ( \9093 , \9091 , \9092 );
and \g451645/U$2 ( \9094 , \8378 , RIdf3aed0_2047);
and \g451645/U$3 ( \9095 , RIe1418e8_2123, \8417 );
nor \g451645/U$1 ( \9096 , \9094 , \9095 );
nand \g447628/U$1 ( \9097 , \9082 , \9090 , \9093 , \9096 );
nor \g445945/U$1 ( \9098 , \9077 , \9078 , \9097 );
and \g451640/U$2 ( \9099 , \8335 , RIdf2fc38_1920);
and \g451640/U$3 ( \9100 , RIfcae9f8_7009, \8531 );
nor \g451640/U$1 ( \9101 , \9099 , \9100 );
and \g451638/U$2 ( \9102 , \8317 , RIdf31b28_1942);
and \g451638/U$3 ( \9103 , RIdf33ce8_1966, \8326 );
nor \g451638/U$1 ( \9104 , \9102 , \9103 );
and \g445109/U$2 ( \9105 , \9098 , \9101 , \9104 );
nor \g445109/U$1 ( \9106 , \9105 , \8422 );
or \g444364/U$1 ( \9107 , \8979 , \9046 , \9076 , \9106 );
and \g445933/U$2 ( \9108 , RIdeaf718_460, \8356 );
and \g445933/U$3 ( \9109 , RIfce20a0_7594, \8340 );
and \g448794/U$2 ( \9110 , RIee20350_4825, \8373 );
and \g448794/U$3 ( \9111 , \8330 , RIdec3218_684);
and \g448794/U$4 ( \9112 , RIdeb2418_492, \8488 );
nor \g448794/U$1 ( \9113 , \9110 , \9111 , \9112 );
and \g455027/U$2 ( \9114 , \8313 , RIdebab18_588);
and \g455027/U$3 ( \9115 , RIdebd818_620, \8323 );
nor \g455027/U$1 ( \9116 , \9114 , \9115 );
not \g449822/U$3 ( \9117 , \9116 );
not \g449822/U$4 ( \9118 , \8376 );
and \g449822/U$2 ( \9119 , \9117 , \9118 );
and \g449822/U$5 ( \9120 , \8359 , RIfce4da0_7626);
nor \g449822/U$1 ( \9121 , \9119 , \9120 );
and \g454010/U$2 ( \9122 , \8404 , RIdec0518_652);
and \g454010/U$3 ( \9123 , RIdec5f18_716, \8351 );
nor \g454010/U$1 ( \9124 , \9122 , \9123 );
and \g451598/U$2 ( \9125 , \8378 , RIdeb7e18_556);
and \g451598/U$3 ( \9126 , RIee1f6a8_4816, \8417 );
nor \g451598/U$1 ( \9127 , \9125 , \9126 );
nand \g447622/U$1 ( \9128 , \9113 , \9121 , \9124 , \9127 );
nor \g445933/U$1 ( \9129 , \9108 , \9109 , \9128 );
and \g454128/U$2 ( \9130 , \8335 , RIde9ec60_364);
and \g454128/U$3 ( \9131 , RIfcea908_7691, \8523 );
nor \g454128/U$1 ( \9132 , \9130 , \9131 );
and \g451590/U$2 ( \9133 , \8319 , RIdea5560_396);
and \g451590/U$3 ( \9134 , RIdeabe60_428, \8324 );
nor \g451590/U$1 ( \9135 , \9133 , \9134 );
and \g445100/U$2 ( \9136 , \9129 , \9132 , \9135 );
nor \g445100/U$1 ( \9137 , \9136 , \8589 );
and \g445936/U$2 ( \9138 , RIde920f0_302, \8417 );
and \g445936/U$3 ( \9139 , RIee1ad88_4764, \8404 );
and \g448799/U$2 ( \9140 , RIe16a130_2584, \8319 );
and \g448799/U$3 ( \9141 , \8324 , RIe16c020_2606);
and \g448799/U$4 ( \9142 , RIee1c2a0_4779, \8330 );
nor \g448799/U$1 ( \9143 , \9140 , \9141 , \9142 );
and \g453519/U$2 ( \9144 , \8335 , RIe1687e0_2566);
and \g453519/U$3 ( \9145 , RIfcae2f0_7004, \8340 );
nor \g453519/U$1 ( \9146 , \9144 , \9145 );
and \g454727/U$2 ( \9147 , \8313 , RIfc5dc38_6089);
and \g454727/U$3 ( \9148 , RIfc6f848_6291, \8323 );
nor \g454727/U$1 ( \9149 , \9147 , \9148 );
not \g450350/U$3 ( \9150 , \9149 );
not \g450350/U$4 ( \9151 , \8347 );
and \g450350/U$2 ( \9152 , \9150 , \9151 );
and \g450350/U$5 ( \9153 , \8351 , RIfce6420_7642);
nor \g450350/U$1 ( \9154 , \9152 , \9153 );
and \g451613/U$2 ( \9155 , \8356 , RIfc76b98_6373);
and \g451613/U$3 ( \9156 , RIde82790_226, \8359 );
nor \g451613/U$1 ( \9157 , \9155 , \9156 );
nand \g447625/U$1 ( \9158 , \9143 , \9146 , \9154 , \9157 );
nor \g445936/U$1 ( \9159 , \9138 , \9139 , \9158 );
and \g451608/U$2 ( \9160 , \8378 , RIfea3fe0_8210);
and \g451608/U$3 ( \9161 , RIfc75950_6360, \8373 );
nor \g451608/U$1 ( \9162 , \9160 , \9161 );
and \g451605/U$2 ( \9163 , \8412 , RIfeaa688_8255);
and \g451605/U$3 ( \9164 , RIfea4148_8211, \8409 );
nor \g451605/U$1 ( \9165 , \9163 , \9164 );
and \g445101/U$2 ( \9166 , \9159 , \9162 , \9165 );
nor \g445101/U$1 ( \9167 , \9166 , \8558 );
or \g444274/U$1 ( \9168 , \9107 , \9137 , \9167 );
_DC \g233f/U$1 ( \9169 , \9168 , \8654 );
nor \g448307/U$1 ( \9170 , \8589 , \8437 );
and \g446796/U$2 ( \9171 , \9170 , RIdeb7cb0_555);
nor \g448349/U$1 ( \9172 , \8589 , \8413 );
and \g446796/U$3 ( \9173 , RIdeba9b0_587, \9172 );
nor \g446796/U$1 ( \9174 , \9171 , \9173 );
and \g446007/U$2 ( \9175 , RIdeb22b0_491, \8488 );
and \g446007/U$3 ( \9176 , RIfc40fe8_5765, \8359 );
and \g448891/U$2 ( \9177 , RIdebd6b0_619, \8409 );
and \g448891/U$3 ( \9178 , \8373 , RIee201e8_4824);
and \g448891/U$4 ( \9179 , RIdec30b0_683, \8383 );
nor \g448891/U$1 ( \9180 , \9177 , \9178 , \9179 );
and \g451894/U$2 ( \9181 , \8335 , RIde9e918_363);
and \g451894/U$3 ( \9182 , RIee1dd58_4798, \8340 );
nor \g451894/U$1 ( \9183 , \9181 , \9182 );
and \g451891/U$2 ( \9184 , \8404 , RIdec03b0_651);
and \g451891/U$3 ( \9185 , RIdec5db0_715, \8351 );
nor \g451891/U$1 ( \9186 , \9184 , \9185 );
and \g454907/U$2 ( \9187 , \8313 , RIdea5218_395);
and \g454907/U$3 ( \9188 , RIdeabb18_427, \8323 );
nor \g454907/U$1 ( \9189 , \9187 , \9188 );
not \g454906/U$1 ( \9190 , \9189 );
and \g449913/U$2 ( \9191 , \9190 , \8316 );
and \g449913/U$3 ( \9192 , RIfcaf538_7017, \8417 );
nor \g449913/U$1 ( \9193 , \9191 , \9192 );
nand \g448180/U$1 ( \9194 , \9180 , \9183 , \9186 , \9193 );
nor \g446007/U$1 ( \9195 , \9175 , \9176 , \9194 );
not \g444816/U$3 ( \9196 , \9195 );
not \g444816/U$4 ( \9197 , \8589 );
and \g444816/U$2 ( \9198 , \9196 , \9197 );
and \g446011/U$2 ( \9199 , RIde865e8_245, \8378 );
and \g446011/U$3 ( \9200 , RIde82448_225, \8359 );
and \g448897/U$2 ( \9201 , RIe169fc8_2583, \8317 );
and \g448897/U$3 ( \9202 , \8326 , RIfec5eb0_8372);
and \g448897/U$4 ( \9203 , RIde8e928_285, \8409 );
nor \g448897/U$1 ( \9204 , \9201 , \9202 , \9203 );
and \g451909/U$2 ( \9205 , \8335 , RIe168678_2565);
and \g451909/U$3 ( \9206 , RIfced8d8_7725, \8340 );
nor \g451909/U$1 ( \9207 , \9205 , \9206 );
and \g451907/U$2 ( \9208 , \8404 , RIfcc92a8_7311);
and \g451907/U$3 ( \9209 , RIee1d218_4790, \8351 );
nor \g451907/U$1 ( \9210 , \9208 , \9209 );
and \g454209/U$2 ( \9211 , \8313 , RIfce62b8_7641);
and \g454209/U$3 ( \9212 , RIfcedd10_7728, \8323 );
nor \g454209/U$1 ( \9213 , \9211 , \9212 );
not \g449918/U$3 ( \9214 , \9213 );
not \g449918/U$4 ( \9215 , \8328 );
and \g449918/U$2 ( \9216 , \9214 , \9215 );
and \g449918/U$5 ( \9217 , \8417 , RIde91da8_301);
nor \g449918/U$1 ( \9218 , \9216 , \9217 );
nand \g447667/U$1 ( \9219 , \9204 , \9207 , \9210 , \9218 );
nor \g446011/U$1 ( \9220 , \9199 , \9200 , \9219 );
and \g451903/U$2 ( \9221 , \8356 , RIfcc19b8_7225);
and \g451903/U$3 ( \9222 , RIde8a788_265, \8414 );
nor \g451903/U$1 ( \9223 , \9221 , \9222 );
and \g451901/U$2 ( \9224 , \8531 , RIfc750e0_6354);
and \g451901/U$3 ( \9225 , RIfea1448_8179, \8488 );
nor \g451901/U$1 ( \9226 , \9224 , \9225 );
and \g445158/U$2 ( \9227 , \9220 , \9223 , \9226 );
nor \g445158/U$1 ( \9228 , \9227 , \8558 );
nor \g444816/U$1 ( \9229 , \9198 , \9228 );
nor \g448310/U$1 ( \9230 , \8589 , \8520 );
and \g446793/U$2 ( \9231 , \9230 , RIdeaf5b0_459);
nor \g448368/U$1 ( \9232 , \8589 , \8524 );
and \g446793/U$3 ( \9233 , RIfcd08c8_7395, \9232 );
nor \g446793/U$1 ( \9234 , \9231 , \9233 );
nand \g444425/U$1 ( \9235 , \9174 , \9229 , \9234 );
and \g451944/U$2 ( \9236 , \8531 , RIee35200_5063);
and \g451944/U$3 ( \9237 , RIe1522b0_2312, \8486 );
nor \g451944/U$1 ( \9238 , \9236 , \9237 );
and \g446020/U$2 ( \9239 , RIe154fb0_2344, \8378 );
and \g446020/U$3 ( \9240 , RIfea1718_8181, \8359 );
and \g448908/U$2 ( \9241 , RIe149bb0_2216, \8319 );
and \g448908/U$3 ( \9242 , \8326 , RIe14c8b0_2248);
and \g448908/U$4 ( \9243 , RIe15d6b0_2440, \8409 );
nor \g448908/U$1 ( \9244 , \9241 , \9242 , \9243 );
and \g451935/U$2 ( \9245 , \8335 , RIe146eb0_2184);
and \g451935/U$3 ( \9246 , RIfcb0348_7027, \8340 );
nor \g451935/U$1 ( \9247 , \9245 , \9246 );
and \g451783/U$2 ( \9248 , \8404 , RIe1603b0_2472);
and \g451783/U$3 ( \9249 , RIe165db0_2536, \8351 );
nor \g451783/U$1 ( \9250 , \9248 , \9249 );
and \g455086/U$2 ( \9251 , \8313 , RIfccfc20_7386);
and \g455086/U$3 ( \9252 , RIe1630b0_2504, \8323 );
nor \g455086/U$1 ( \9253 , \9251 , \9252 );
not \g449927/U$3 ( \9254 , \9253 );
not \g449927/U$4 ( \9255 , \8328 );
and \g449927/U$2 ( \9256 , \9254 , \9255 );
and \g449927/U$5 ( \9257 , \8417 , RIee365b0_5077);
nor \g449927/U$1 ( \9258 , \9256 , \9257 );
nand \g447670/U$1 ( \9259 , \9244 , \9247 , \9250 , \9258 );
nor \g446020/U$1 ( \9260 , \9239 , \9240 , \9259 );
and \g451932/U$2 ( \9261 , \8356 , RIe14f5b0_2280);
and \g451932/U$3 ( \9262 , RIe157cb0_2376, \8412 );
nor \g451932/U$1 ( \9263 , \9261 , \9262 );
nand \g445580/U$1 ( \9264 , \9238 , \9260 , \9263 );
and \g444851/U$2 ( \9265 , \9264 , \8369 );
not \g448463/U$1 ( \9266 , \8422 );
and \g448901/U$2 ( \9267 , RIfec5be0_8370, \8414 );
and \g448901/U$3 ( \9268 , \8407 , RIe13f2f0_2096);
and \g448901/U$4 ( \9269 , RIdf33b80_1965, \8326 );
nor \g448901/U$1 ( \9270 , \9267 , \9268 , \9269 );
and \g451927/U$2 ( \9271 , \8356 , RIfc74438_6345);
and \g451927/U$3 ( \9272 , RIfea15b0_8180, \8359 );
nor \g451927/U$1 ( \9273 , \9271 , \9272 );
and \g454714/U$2 ( \9274 , \8313 , RIfcae728_7007);
and \g454714/U$3 ( \9275 , RIfc5fb28_6111, \8323 );
nor \g454714/U$1 ( \9276 , \9274 , \9275 );
not \g449922/U$3 ( \9277 , \9276 );
not \g449922/U$4 ( \9278 , \8347 );
and \g449922/U$2 ( \9279 , \9277 , \9278 );
and \g449922/U$5 ( \9280 , \8340 , RIdf36178_1992);
nor \g449922/U$1 ( \9281 , \9279 , \9280 );
and \g451924/U$2 ( \9282 , \8378 , RIdf3ad68_2046);
and \g451924/U$3 ( \9283 , RIe141780_2122, \8417 );
nor \g451924/U$1 ( \9284 , \9282 , \9283 );
nand \g447669/U$1 ( \9285 , \9270 , \9273 , \9281 , \9284 );
and \g444851/U$3 ( \9286 , \9266 , \9285 );
nor \g444851/U$1 ( \9287 , \9265 , \9286 );
nor \g448410/U$1 ( \9288 , \8422 , \8425 );
and \g446800/U$2 ( \9289 , \9288 , RIfc94f58_6717);
nor \g448439/U$1 ( \9290 , \8422 , \8372 );
and \g446800/U$3 ( \9291 , RIee32500_5031, \9290 );
nor \g446800/U$1 ( \9292 , \9289 , \9291 );
nor \g448437/U$1 ( \9293 , \8422 , \8382 );
and \g446801/U$2 ( \9294 , \9293 , RIfcdf238_7561);
not \g455453/U$1 ( \9295 , \8351 );
nor \g448436/U$1 ( \9296 , \8422 , \9295 );
and \g446801/U$3 ( \9297 , RIfc73790_6336, \9296 );
nor \g446801/U$1 ( \9298 , \9294 , \9297 );
nor \g448409/U$1 ( \9299 , \8422 , \8508 );
and \g446802/U$2 ( \9300 , \9299 , RIdf2fad0_1919);
nor \g448417/U$1 ( \9301 , \8422 , \8318 );
and \g446802/U$3 ( \9302 , RIdf319c0_1941, \9301 );
nor \g446802/U$1 ( \9303 , \9300 , \9302 );
nand \g444601/U$1 ( \9304 , \9287 , \9292 , \9298 , \9303 );
and \g445999/U$2 ( \9305 , RIdf03e80_1421, \8378 );
and \g445999/U$3 ( \9306 , RIdefe480_1357, \8359 );
and \g448881/U$2 ( \9307 , RIdf09880_1485, \8409 );
and \g448881/U$3 ( \9308 , \8373 , RIdf11f80_1581);
and \g448881/U$4 ( \9309 , RIdf14c80_1613, \8330 );
nor \g448881/U$1 ( \9310 , \9307 , \9308 , \9309 );
and \g451865/U$2 ( \9311 , \8335 , RIdeea980_1133);
and \g451865/U$3 ( \9312 , RIdef3080_1229, \8340 );
nor \g451865/U$1 ( \9313 , \9311 , \9312 );
and \g451864/U$2 ( \9314 , \8404 , RIdf0f280_1549);
and \g451864/U$3 ( \9315 , RIdf17980_1645, \8351 );
nor \g451864/U$1 ( \9316 , \9314 , \9315 );
and \g454208/U$2 ( \9317 , \8313 , RIdeed680_1165);
and \g454208/U$3 ( \9318 , RIdef0380_1197, \8323 );
nor \g454208/U$1 ( \9319 , \9317 , \9318 );
not \g454207/U$1 ( \9320 , \9319 );
and \g449902/U$2 ( \9321 , \9320 , \8316 );
and \g449902/U$3 ( \9322 , RIdf0c580_1517, \8417 );
nor \g449902/U$1 ( \9323 , \9321 , \9322 );
nand \g448177/U$1 ( \9324 , \9310 , \9313 , \9316 , \9323 );
nor \g445999/U$1 ( \9325 , \9305 , \9306 , \9324 );
and \g451859/U$2 ( \9326 , \8356 , RIdef5d80_1261);
and \g451859/U$3 ( \9327 , RIdf06b80_1453, \8414 );
nor \g451859/U$1 ( \9328 , \9326 , \9327 );
and \g453423/U$2 ( \9329 , \8531 , RIdef8a80_1293);
and \g453423/U$3 ( \9330 , RIdefb780_1325, \8488 );
nor \g453423/U$1 ( \9331 , \9329 , \9330 );
and \g445150/U$2 ( \9332 , \9325 , \9328 , \9331 );
nor \g445150/U$1 ( \9333 , \9332 , \8477 );
and \g446004/U$2 ( \9334 , RIfea12e0_8178, \8378 );
and \g446004/U$3 ( \9335 , RIfc679b8_6201, \8359 );
and \g448885/U$2 ( \9336 , RIfea7f28_8227, \8409 );
and \g448885/U$3 ( \9337 , \8371 , RIfcccf20_7354);
and \g448885/U$4 ( \9338 , RIfcac568_6983, \8383 );
nor \g448885/U$1 ( \9339 , \9336 , \9337 , \9338 );
and \g451881/U$2 ( \9340 , \8335 , RIfec5d48_8371);
and \g451881/U$3 ( \9341 , RIdeda120_945, \8340 );
nor \g451881/U$1 ( \9342 , \9340 , \9341 );
and \g453667/U$2 ( \9343 , \8404 , RIfccd358_7357);
and \g453667/U$3 ( \9344 , RIfc595e8_6039, \8351 );
nor \g453667/U$1 ( \9345 , \9343 , \9344 );
and \g454807/U$2 ( \9346 , \8313 , RIded5c38_896);
and \g454807/U$3 ( \9347 , RIded7b28_918, \8323 );
nor \g454807/U$1 ( \9348 , \9346 , \9347 );
not \g454806/U$1 ( \9349 , \9348 );
and \g449908/U$2 ( \9350 , \9349 , \8316 );
and \g449908/U$3 ( \9351 , RIdee5250_1071, \8417 );
nor \g449908/U$1 ( \9352 , \9350 , \9351 );
nand \g448178/U$1 ( \9353 , \9339 , \9342 , \9345 , \9352 );
nor \g446004/U$1 ( \9354 , \9334 , \9335 , \9353 );
and \g451877/U$2 ( \9355 , \8356 , RIfc6cb48_6259);
and \g451877/U$3 ( \9356 , RIdee11a0_1025, \8414 );
nor \g451877/U$1 ( \9357 , \9355 , \9356 );
and \g451874/U$2 ( \9358 , \8523 , RIfc6dd90_6272);
and \g451874/U$3 ( \9359 , RIee22510_4849, \8486 );
nor \g451874/U$1 ( \9360 , \9358 , \9359 );
and \g445152/U$2 ( \9361 , \9354 , \9357 , \9360 );
nor \g445152/U$1 ( \9362 , \9361 , \8481 );
or \g444294/U$1 ( \9363 , \9235 , \9304 , \9333 , \9362 );
and \g445992/U$2 ( \9364 , RIdf24f40_1797, \8378 );
and \g445992/U$3 ( \9365 , RIfc64b50_6168, \8359 );
and \g448870/U$2 ( \9366 , RIdf1b490_1687, \8319 );
and \g448870/U$3 ( \9367 , \8326 , RIfeaad90_8260);
and \g448870/U$4 ( \9368 , RIdf288e8_1838, \8409 );
nor \g448870/U$1 ( \9369 , \9366 , \9367 , \9368 );
and \g451839/U$2 ( \9370 , \8335 , RIdf19b40_1669);
and \g451839/U$3 ( \9371 , RIdf21ca0_1761, \8340 );
nor \g451839/U$1 ( \9372 , \9370 , \9371 );
and \g451317/U$2 ( \9373 , \8404 , RIfc704f0_6300);
and \g451317/U$3 ( \9374 , RIee2c290_4961, \8351 );
nor \g451317/U$1 ( \9375 , \9373 , \9374 );
and \g455095/U$2 ( \9376 , \8313 , RIfc70658_6301);
and \g455095/U$3 ( \9377 , RIee2a940_4943, \8323 );
nor \g455095/U$1 ( \9378 , \9376 , \9377 );
not \g449892/U$3 ( \9379 , \9378 );
not \g449892/U$4 ( \9380 , \8328 );
and \g449892/U$2 ( \9381 , \9379 , \9380 );
and \g449892/U$5 ( \9382 , \8417 , RIdf2aaa8_1862);
nor \g449892/U$1 ( \9383 , \9381 , \9382 );
nand \g447654/U$1 ( \9384 , \9369 , \9372 , \9375 , \9383 );
nor \g445992/U$1 ( \9385 , \9364 , \9365 , \9384 );
and \g451832/U$2 ( \9386 , \8356 , RIfcad4e0_6994);
and \g451832/U$3 ( \9387 , RIdf269f8_1816, \8414 );
nor \g451832/U$1 ( \9388 , \9386 , \9387 );
and \g451831/U$2 ( \9389 , \8531 , RIdf231b8_1776);
and \g451831/U$3 ( \9390 , RIfccaa90_7328, \8488 );
nor \g451831/U$1 ( \9391 , \9389 , \9390 );
and \g445144/U$2 ( \9392 , \9385 , \9388 , \9391 );
nor \g445144/U$1 ( \9393 , \9392 , \8621 );
and \g445997/U$2 ( \9394 , RIded11b0_843, \8351 );
and \g445997/U$3 ( \9395 , RIde7df60_204, \8335 );
and \g448875/U$2 ( \9396 , RIdee7c80_1101, \8326 );
and \g448875/U$3 ( \9397 , \8531 , RIdf2d208_1890);
and \g448875/U$4 ( \9398 , RIdf38ba8_2022, \8488 );
nor \g448875/U$1 ( \9399 , \9396 , \9397 , \9398 );
and \g451853/U$2 ( \9400 , \8356 , RIdf1da88_1714);
and \g451853/U$3 ( \9401 , RIe1441b0_2152, \8359 );
nor \g451853/U$1 ( \9402 , \9400 , \9401 );
and \g454224/U$2 ( \9403 , \8313 , RIe16ebb8_2637);
and \g454224/U$3 ( \9404 , RIde98018_331, \8323 );
nor \g454224/U$1 ( \9405 , \9403 , \9404 );
not \g449898/U$3 ( \9406 , \9405 );
not \g449898/U$4 ( \9407 , \8376 );
and \g449898/U$2 ( \9408 , \9406 , \9407 );
and \g449898/U$5 ( \9409 , \8340 , RIdf01180_1389);
nor \g449898/U$1 ( \9410 , \9408 , \9409 );
and \g451850/U$2 ( \9411 , \8378 , RIe15a9b0_2408);
and \g451850/U$3 ( \9412 , RIdeb4fb0_523, \8417 );
nor \g451850/U$1 ( \9413 , \9411 , \9412 );
nand \g447655/U$1 ( \9414 , \9399 , \9402 , \9410 , \9413 );
nor \g445997/U$1 ( \9415 , \9394 , \9395 , \9414 );
and \g451849/U$2 ( \9416 , \8319 , RIdedc9e8_974);
and \g451849/U$3 ( \9417 , RIdec8ab0_747, \8404 );
nor \g451849/U$1 ( \9418 , \9416 , \9417 );
and \g451847/U$2 ( \9419 , \8373 , RIdecb7b0_779);
and \g451847/U$3 ( \9420 , RIdece4b0_811, \8383 );
nor \g451847/U$1 ( \9421 , \9419 , \9420 );
and \g445146/U$2 ( \9422 , \9415 , \9418 , \9421 );
nor \g445146/U$1 ( \9423 , \9422 , \8651 );
or \g444163/U$1 ( \9424 , \9363 , \9393 , \9423 );
_DC \g23c4/U$1 ( \9425 , \9424 , \8654 );
and \g450710/U$2 ( \9426 , \8326 , RIdf20080_1741);
and \g450710/U$3 ( \9427 , RIee28078_4914, \8404 );
nor \g450710/U$1 ( \9428 , \9426 , \9427 );
and \g445736/U$2 ( \9429 , RIee292c0_4927, \8373 );
and \g445736/U$3 ( \9430 , RIdf1b328_1686, \8319 );
and \g448538/U$2 ( \9431 , RIdf23050_1775, \8523 );
and \g448538/U$3 ( \9432 , \8486 , RIfca0628_6847);
and \g448538/U$4 ( \9433 , RIee2a7d8_4942, \8383 );
nor \g448538/U$1 ( \9434 , \9431 , \9432 , \9433 );
and \g450717/U$2 ( \9435 , \8356 , RIfcd3190_7424);
and \g450717/U$3 ( \9436 , RIfcd4f18_7445, \8359 );
nor \g450717/U$1 ( \9437 , \9435 , \9436 );
and \g454222/U$2 ( \9438 , \8313 , RIfea0a70_8172);
and \g454222/U$3 ( \9439 , RIdf28780_1837, \8323 );
nor \g454222/U$1 ( \9440 , \9438 , \9439 );
not \g449560/U$3 ( \9441 , \9440 );
not \g449560/U$4 ( \9442 , \8376 );
and \g449560/U$2 ( \9443 , \9441 , \9442 );
and \g449560/U$5 ( \9444 , \8351 , RIee2c128_4960);
nor \g449560/U$1 ( \9445 , \9443 , \9444 );
and \g450714/U$2 ( \9446 , \8378 , RIfea0908_8171);
and \g450714/U$3 ( \9447 , RIdf2a940_1861, \8417 );
nor \g450714/U$1 ( \9448 , \9446 , \9447 );
nand \g447476/U$1 ( \9449 , \9434 , \9437 , \9445 , \9448 );
nor \g445736/U$1 ( \9450 , \9429 , \9430 , \9449 );
and \g450712/U$2 ( \9451 , \8335 , RIdf199d8_1668);
and \g450712/U$3 ( \9452 , RIdf21b38_1760, \8340 );
nor \g450712/U$1 ( \9453 , \9451 , \9452 );
nand \g445514/U$1 ( \9454 , \9428 , \9450 , \9453 );
and \g444721/U$2 ( \9455 , \9454 , \8752 );
and \g448533/U$2 ( \9456 , RIdf06a18_1452, \8414 );
and \g448533/U$3 ( \9457 , \8407 , RIdf09718_1484);
and \g448533/U$4 ( \9458 , RIdf14b18_1612, \8383 );
nor \g448533/U$1 ( \9459 , \9456 , \9457 , \9458 );
and \g450703/U$2 ( \9460 , \8356 , RIdef5c18_1260);
and \g450703/U$3 ( \9461 , RIdefe318_1356, \8359 );
nor \g450703/U$1 ( \9462 , \9460 , \9461 );
and \g454268/U$2 ( \9463 , \8313 , RIdef8918_1292);
and \g454268/U$3 ( \9464 , RIdefb618_1324, \8323 );
nor \g454268/U$1 ( \9465 , \9463 , \9464 );
not \g449553/U$3 ( \9466 , \9465 );
not \g449553/U$4 ( \9467 , \8347 );
and \g449553/U$2 ( \9468 , \9466 , \9467 );
and \g449553/U$5 ( \9469 , \8351 , RIdf17818_1644);
nor \g449553/U$1 ( \9470 , \9468 , \9469 );
and \g450701/U$2 ( \9471 , \8378 , RIdf03d18_1420);
and \g450701/U$3 ( \9472 , RIdf0c418_1516, \8417 );
nor \g450701/U$1 ( \9473 , \9471 , \9472 );
nand \g447475/U$1 ( \9474 , \9459 , \9462 , \9470 , \9473 );
and \g444721/U$3 ( \9475 , \8478 , \9474 );
nor \g444721/U$1 ( \9476 , \9455 , \9475 );
and \g446533/U$2 ( \9477 , \8780 , RIdef0218_1196);
and \g446533/U$3 ( \9478 , RIdef2f18_1228, \8782 );
nor \g446533/U$1 ( \9479 , \9477 , \9478 );
nor \g448314/U$1 ( \9480 , \8477 , \8425 );
and \g446532/U$2 ( \9481 , \9480 , RIdf0f118_1548);
nor \g448366/U$1 ( \9482 , \8477 , \8372 );
and \g446532/U$3 ( \9483 , RIdf11e18_1580, \9482 );
nor \g446532/U$1 ( \9484 , \9481 , \9483 );
and \g446534/U$2 ( \9485 , \8785 , RIdeea818_1132);
and \g446534/U$3 ( \9486 , RIdeed518_1164, \8787 );
nor \g446534/U$1 ( \9487 , \9485 , \9486 );
nand \g444552/U$1 ( \9488 , \9476 , \9479 , \9484 , \9487 );
and \g450735/U$2 ( \9489 , \8324 , RIdee7b18_1100);
and \g450735/U$3 ( \9490 , RIdec8948_746, \8404 );
nor \g450735/U$1 ( \9491 , \9489 , \9490 );
and \g445741/U$2 ( \9492 , RIdecb648_778, \8373 );
and \g445741/U$3 ( \9493 , RIdedc880_973, \8317 );
and \g448545/U$2 ( \9494 , RIe16ea50_2636, \8414 );
and \g448545/U$3 ( \9495 , \8407 , RIde97cd0_330);
and \g448545/U$4 ( \9496 , RIdece348_810, \8330 );
nor \g448545/U$1 ( \9497 , \9494 , \9495 , \9496 );
and \g450742/U$2 ( \9498 , \8356 , RIdf1d920_1713);
and \g450742/U$3 ( \9499 , RIe144048_2151, \8359 );
nor \g450742/U$1 ( \9500 , \9498 , \9499 );
and \g454235/U$2 ( \9501 , \8313 , RIdf2d0a0_1889);
and \g454235/U$3 ( \9502 , RIdf38a40_2021, \8323 );
nor \g454235/U$1 ( \9503 , \9501 , \9502 );
not \g449568/U$3 ( \9504 , \9503 );
not \g449568/U$4 ( \9505 , \8347 );
and \g449568/U$2 ( \9506 , \9504 , \9505 );
and \g449568/U$5 ( \9507 , \8351 , RIded1048_842);
nor \g449568/U$1 ( \9508 , \9506 , \9507 );
and \g450740/U$2 ( \9509 , \8378 , RIe15a848_2407);
and \g450740/U$3 ( \9510 , RIdeb4e48_522, \8417 );
nor \g450740/U$1 ( \9511 , \9509 , \9510 );
nand \g447480/U$1 ( \9512 , \9497 , \9500 , \9508 , \9511 );
nor \g445741/U$1 ( \9513 , \9492 , \9493 , \9512 );
and \g450737/U$2 ( \9514 , \8335 , RIde7dc18_203);
and \g450737/U$3 ( \9515 , RIdf01018_1388, \8340 );
nor \g450737/U$1 ( \9516 , \9514 , \9515 );
nand \g445516/U$1 ( \9517 , \9491 , \9513 , \9516 );
and \g444871/U$2 ( \9518 , \9517 , \9010 );
and \g448541/U$2 ( \9519 , RIded5ad0_895, \8319 );
and \g448541/U$3 ( \9520 , \8326 , RIded79c0_917);
and \g448541/U$4 ( \9521 , RIfcd4978_7441, \8486 );
nor \g448541/U$1 ( \9522 , \9519 , \9520 , \9521 );
and \g450731/U$2 ( \9523 , \8335 , RIfeab498_8265);
and \g450731/U$3 ( \9524 , RIded9fb8_944, \8340 );
nor \g450731/U$1 ( \9525 , \9523 , \9524 );
and \g450726/U$2 ( \9526 , \8404 , RIfcdc6a0_7530);
and \g450726/U$3 ( \9527 , RIfcdf3a0_7562, \8351 );
nor \g450726/U$1 ( \9528 , \9526 , \9527 );
and \g454840/U$2 ( \9529 , \8313 , RIfcdc538_7529);
and \g454840/U$3 ( \9530 , RIfca5218_6901, \8323 );
nor \g454840/U$1 ( \9531 , \9529 , \9530 );
not \g449564/U$3 ( \9532 , \9531 );
not \g449564/U$4 ( \9533 , \8328 );
and \g449564/U$2 ( \9534 , \9532 , \9533 );
and \g449564/U$5 ( \9535 , \8359 , RIfcb0d20_7034);
nor \g449564/U$1 ( \9536 , \9534 , \9535 );
nand \g447479/U$1 ( \9537 , \9522 , \9525 , \9528 , \9536 );
and \g444871/U$3 ( \9538 , \8482 , \9537 );
nor \g444871/U$1 ( \9539 , \9518 , \9538 );
and \g446538/U$2 ( \9540 , \8964 , RIdee3360_1049);
and \g446538/U$3 ( \9541 , RIdee50e8_1070, \8966 );
nor \g446538/U$1 ( \9542 , \9540 , \9541 );
and \g446539/U$2 ( \9543 , \8521 , RIfca1708_6859);
and \g446539/U$3 ( \9544 , RIfca49a8_6895, \8525 );
nor \g446539/U$1 ( \9545 , \9543 , \9544 );
and \g446540/U$2 ( \9546 , \8974 , RIdedefe0_1001);
and \g446540/U$3 ( \9547 , RIfea07a0_8170, \8976 );
nor \g446540/U$1 ( \9548 , \9546 , \9547 );
nand \g444553/U$1 ( \9549 , \9539 , \9542 , \9545 , \9548 );
and \g445724/U$2 ( \9550 , RIde8e5e0_284, \8409 );
and \g445724/U$3 ( \9551 , RIfea0bd8_8173, \8378 );
and \g448525/U$2 ( \9552 , RIfcdbb60_7522, \8373 );
and \g448525/U$3 ( \9553 , \8383 , RIfc5b0a0_6058);
and \g448525/U$4 ( \9554 , RIfcb1b30_7044, \8488 );
nor \g448525/U$1 ( \9555 , \9552 , \9553 , \9554 );
and \g450667/U$2 ( \9556 , \8335 , RIe168510_2564);
and \g450667/U$3 ( \9557 , RIfc77b10_6384, \8340 );
nor \g450667/U$1 ( \9558 , \9556 , \9557 );
and \g450665/U$2 ( \9559 , \8404 , RIfc78650_6392);
and \g450665/U$3 ( \9560 , RIfc41e70_5772, \8351 );
nor \g450665/U$1 ( \9561 , \9559 , \9560 );
and \g454205/U$2 ( \9562 , \8313 , RIe169e60_2582);
and \g454205/U$3 ( \9563 , RIe16beb8_2605, \8323 );
nor \g454205/U$1 ( \9564 , \9562 , \9563 );
not \g454204/U$1 ( \9565 , \9564 );
and \g449545/U$2 ( \9566 , \9565 , \8316 );
and \g449545/U$3 ( \9567 , RIfcdf508_7563, \8359 );
nor \g449545/U$1 ( \9568 , \9566 , \9567 );
nand \g448134/U$1 ( \9569 , \9555 , \9558 , \9561 , \9568 );
nor \g445724/U$1 ( \9570 , \9550 , \9551 , \9569 );
and \g450657/U$2 ( \9571 , \8356 , RIfcb16f8_7041);
and \g450657/U$3 ( \9572 , RIfea92d8_8241, \8417 );
nor \g450657/U$1 ( \9573 , \9571 , \9572 );
and \g450656/U$2 ( \9574 , \8531 , RIfc5ccc0_6078);
and \g450656/U$3 ( \9575 , RIfea0d40_8174, \8414 );
nor \g450656/U$1 ( \9576 , \9574 , \9575 );
and \g444945/U$2 ( \9577 , \9570 , \9573 , \9576 );
nor \g444945/U$1 ( \9578 , \9577 , \8558 );
and \g445727/U$2 ( \9579 , RIfca38c8_6883, \8340 );
and \g445727/U$3 ( \9580 , RIdec0248_650, \8404 );
and \g448530/U$2 ( \9581 , RIfce7aa0_7658, \8531 );
and \g448530/U$3 ( \9582 , \8486 , RIdeb2148_490);
and \g448530/U$4 ( \9583 , RIdec2f48_682, \8330 );
nor \g448530/U$1 ( \9584 , \9581 , \9582 , \9583 );
and \g450685/U$2 ( \9585 , \8356 , RIdeaf448_458);
and \g450685/U$3 ( \9586 , RIfce7c08_7659, \8359 );
nor \g450685/U$1 ( \9587 , \9585 , \9586 );
and \g454214/U$2 ( \9588 , \8313 , RIdeba848_586);
and \g454214/U$3 ( \9589 , RIdebd548_618, \8323 );
nor \g454214/U$1 ( \9590 , \9588 , \9589 );
not \g449550/U$3 ( \9591 , \9590 );
not \g449550/U$4 ( \9592 , \8376 );
and \g449550/U$2 ( \9593 , \9591 , \9592 );
and \g449550/U$5 ( \9594 , \8351 , RIdec5c48_714);
nor \g449550/U$1 ( \9595 , \9593 , \9594 );
and \g450683/U$2 ( \9596 , \8378 , RIdeb7b48_554);
and \g450683/U$3 ( \9597 , RIfcb38b8_7065, \8417 );
nor \g450683/U$1 ( \9598 , \9596 , \9597 );
nand \g447472/U$1 ( \9599 , \9584 , \9587 , \9595 , \9598 );
nor \g445727/U$1 ( \9600 , \9579 , \9580 , \9599 );
and \g450676/U$2 ( \9601 , \8335 , RIde9e5d0_362);
and \g450676/U$3 ( \9602 , RIfc7c160_6434, \8373 );
nor \g450676/U$1 ( \9603 , \9601 , \9602 );
and \g450678/U$2 ( \9604 , \8317 , RIdea4ed0_394);
and \g450678/U$3 ( \9605 , RIdeab7d0_426, \8326 );
nor \g450678/U$1 ( \9606 , \9604 , \9605 );
and \g444949/U$2 ( \9607 , \9600 , \9603 , \9606 );
nor \g444949/U$1 ( \9608 , \9607 , \8589 );
or \g444381/U$1 ( \9609 , \9488 , \9549 , \9578 , \9608 );
and \g445717/U$2 ( \9610 , RIfea0ea8_8175, \8407 );
and \g445717/U$3 ( \9611 , RIdf3ac00_2045, \8378 );
and \g448515/U$2 ( \9612 , RIfcc5630_7268, \8371 );
and \g448515/U$3 ( \9613 , \8383 , RIfc9ecd8_6829);
and \g448515/U$4 ( \9614 , RIfcd3cd0_7432, \8486 );
nor \g448515/U$1 ( \9615 , \9612 , \9613 , \9614 );
and \g450630/U$2 ( \9616 , \8335 , RIdf2f968_1918);
and \g450630/U$3 ( \9617 , RIdf36010_1991, \8340 );
nor \g450630/U$1 ( \9618 , \9616 , \9617 );
and \g450629/U$2 ( \9619 , \8404 , RIfc83bb8_6521);
and \g450629/U$3 ( \9620 , RIfc9eb70_6828, \8351 );
nor \g450629/U$1 ( \9621 , \9619 , \9620 );
and \g454448/U$2 ( \9622 , \8313 , RIdf31858_1940);
and \g454448/U$3 ( \9623 , RIdf33a18_1964, \8323 );
nor \g454448/U$1 ( \9624 , \9622 , \9623 );
not \g454447/U$1 ( \9625 , \9624 );
and \g449535/U$2 ( \9626 , \9625 , \8316 );
and \g449535/U$3 ( \9627 , RIee308e0_5011, \8359 );
nor \g449535/U$1 ( \9628 , \9626 , \9627 );
nand \g448133/U$1 ( \9629 , \9615 , \9618 , \9621 , \9628 );
nor \g445717/U$1 ( \9630 , \9610 , \9611 , \9629 );
and \g450624/U$2 ( \9631 , \8356 , RIfc834b0_6516);
and \g450624/U$3 ( \9632 , RIe141618_2121, \8417 );
nor \g450624/U$1 ( \9633 , \9631 , \9632 );
and \g450623/U$2 ( \9634 , \8531 , RIfc84e00_6534);
and \g450623/U$3 ( \9635 , RIdf3d1f8_2072, \8414 );
nor \g450623/U$1 ( \9636 , \9634 , \9635 );
and \g444940/U$2 ( \9637 , \9630 , \9633 , \9636 );
nor \g444940/U$1 ( \9638 , \9637 , \8422 );
and \g445719/U$2 ( \9639 , RIe15d548_2439, \8409 );
and \g445719/U$3 ( \9640 , RIe154e48_2343, \8378 );
and \g448519/U$2 ( \9641 , RIe149a48_2215, \8319 );
and \g448519/U$3 ( \9642 , \8326 , RIe14c748_2247);
and \g448519/U$4 ( \9643 , RIe152148_2311, \8488 );
nor \g448519/U$1 ( \9644 , \9641 , \9642 , \9643 );
and \g450647/U$2 ( \9645 , \8335 , RIe146d48_2183);
and \g450647/U$3 ( \9646 , RIfc865e8_6551, \8340 );
nor \g450647/U$1 ( \9647 , \9645 , \9646 );
and \g450644/U$2 ( \9648 , \8404 , RIe160248_2471);
and \g450644/U$3 ( \9649 , RIe165c48_2535, \8351 );
nor \g450644/U$1 ( \9650 , \9648 , \9649 );
and \g454197/U$2 ( \9651 , \8313 , RIfc4f9d0_5928);
and \g454197/U$3 ( \9652 , RIe162f48_2503, \8323 );
nor \g454197/U$1 ( \9653 , \9651 , \9652 );
not \g449541/U$3 ( \9654 , \9653 );
not \g449541/U$4 ( \9655 , \8328 );
and \g449541/U$2 ( \9656 , \9654 , \9655 );
and \g449541/U$5 ( \9657 , \8359 , RIfc4e1e8_5911);
nor \g449541/U$1 ( \9658 , \9656 , \9657 );
nand \g447470/U$1 ( \9659 , \9644 , \9647 , \9650 , \9658 );
nor \g445719/U$1 ( \9660 , \9639 , \9640 , \9659 );
and \g450641/U$2 ( \9661 , \8356 , RIe14f448_2279);
and \g450641/U$3 ( \9662 , RIfc4e8f0_5916, \8417 );
nor \g450641/U$1 ( \9663 , \9661 , \9662 );
and \g450637/U$2 ( \9664 , \8531 , RIfc868b8_6553);
and \g450637/U$3 ( \9665 , RIe157b48_2375, \8412 );
nor \g450637/U$1 ( \9666 , \9664 , \9665 );
and \g444941/U$2 ( \9667 , \9660 , \9663 , \9666 );
nor \g444941/U$1 ( \9668 , \9667 , \8368 );
or \g444239/U$1 ( \9669 , \9609 , \9638 , \9668 );
_DC \g2449/U$1 ( \9670 , \9669 , \8654 );
and \g450969/U$2 ( \9671 , \8319 , RIfc68930_6212);
and \g450969/U$3 ( \9672 , RIe16bd50_2604, \8324 );
nor \g450969/U$1 ( \9673 , \9671 , \9672 );
and \g445790/U$2 ( \9674 , RIfcd0e68_7399, \8373 );
and \g445790/U$3 ( \9675 , RIe1683a8_2563, \8335 );
and \g448611/U$2 ( \9676 , RIfc52dd8_5965, \8523 );
and \g448611/U$3 ( \9677 , \8488 , RIfc4d810_5904);
and \g448611/U$4 ( \9678 , RIee1c138_4778, \8383 );
nor \g448611/U$1 ( \9679 , \9676 , \9677 , \9678 );
and \g450977/U$2 ( \9680 , \8356 , RIfcde590_7552);
and \g450977/U$3 ( \9681 , RIfcda7b0_7508, \8359 );
nor \g450977/U$1 ( \9682 , \9680 , \9681 );
and \g454323/U$2 ( \9683 , \8313 , RIfe88ec0_7902);
and \g454323/U$3 ( \9684 , RIfe88d58_7901, \8323 );
nor \g454323/U$1 ( \9685 , \9683 , \9684 );
not \g449638/U$3 ( \9686 , \9685 );
not \g449638/U$4 ( \9687 , \8376 );
and \g449638/U$2 ( \9688 , \9686 , \9687 );
and \g449638/U$5 ( \9689 , \8351 , RIee1d0b0_4789);
nor \g449638/U$1 ( \9690 , \9688 , \9689 );
and \g450974/U$2 ( \9691 , \8378 , RIfe88bf0_7900);
and \g450974/U$3 ( \9692 , RIfe89028_7903, \8417 );
nor \g450974/U$1 ( \9693 , \9691 , \9692 );
nand \g447516/U$1 ( \9694 , \9679 , \9682 , \9690 , \9693 );
nor \g445790/U$1 ( \9695 , \9674 , \9675 , \9694 );
and \g450968/U$2 ( \9696 , \8340 , RIfc4f868_5927);
and \g450968/U$3 ( \9697 , RIfc76d00_6374, \8404 );
nor \g450968/U$1 ( \9698 , \9696 , \9697 );
nand \g445527/U$1 ( \9699 , \9673 , \9695 , \9698 );
not \g448465/U$1 ( \9700 , \8558 );
and \g444691/U$2 ( \9701 , \9699 , \9700 );
not \g448481/U$1 ( \9702 , \8589 );
and \g448607/U$2 ( \9703 , RIfc9efa8_6831, \8531 );
and \g448607/U$3 ( \9704 , \8488 , RIdeb1fe0_489);
and \g448607/U$4 ( \9705 , RIdec2de0_681, \8383 );
nor \g448607/U$1 ( \9706 , \9703 , \9704 , \9705 );
and \g450962/U$2 ( \9707 , \8356 , RIdeaf2e0_457);
and \g450962/U$3 ( \9708 , RIfcb9858_7133, \8359 );
nor \g450962/U$1 ( \9709 , \9707 , \9708 );
and \g455287/U$2 ( \9710 , \8313 , RIdeba6e0_585);
and \g455287/U$3 ( \9711 , RIdebd3e0_617, \8323 );
nor \g455287/U$1 ( \9712 , \9710 , \9711 );
not \g449633/U$3 ( \9713 , \9712 );
not \g449633/U$4 ( \9714 , \8376 );
and \g449633/U$2 ( \9715 , \9713 , \9714 );
and \g449633/U$5 ( \9716 , \8351 , RIdec5ae0_713);
nor \g449633/U$1 ( \9717 , \9715 , \9716 );
and \g450959/U$2 ( \9718 , \8378 , RIdeb79e0_553);
and \g450959/U$3 ( \9719 , RIfcb8d18_7125, \8417 );
nor \g450959/U$1 ( \9720 , \9718 , \9719 );
nand \g447515/U$1 ( \9721 , \9706 , \9709 , \9717 , \9720 );
and \g444691/U$3 ( \9722 , \9702 , \9721 );
nor \g444691/U$1 ( \9723 , \9701 , \9722 );
nor \g448313/U$1 ( \9724 , \8589 , \8425 );
and \g446588/U$2 ( \9725 , \9724 , RIdec00e0_649);
nor \g448350/U$1 ( \9726 , \8589 , \8372 );
and \g446588/U$3 ( \9727 , RIfc82268_6503, \9726 );
nor \g446588/U$1 ( \9728 , \9725 , \9727 );
nor \g448312/U$1 ( \9729 , \8589 , \8508 );
and \g446587/U$2 ( \9730 , \9729 , RIde9e288_361);
nor \g448339/U$1 ( \9731 , \8589 , \8318 );
and \g446587/U$3 ( \9732 , RIdea4b88_393, \9731 );
nor \g446587/U$1 ( \9733 , \9730 , \9732 );
nor \g448341/U$1 ( \9734 , \8589 , \8325 );
and \g446586/U$2 ( \9735 , \9734 , RIdeab488_425);
nor \g448369/U$1 ( \9736 , \8589 , \8516 );
and \g446586/U$3 ( \9737 , RIfce0750_7576, \9736 );
nor \g446586/U$1 ( \9738 , \9735 , \9737 );
nand \g444458/U$1 ( \9739 , \9723 , \9728 , \9733 , \9738 );
and \g450997/U$2 ( \9740 , \8319 , RIdedc718_972);
and \g450997/U$3 ( \9741 , RIdee79b0_1099, \8324 );
nor \g450997/U$1 ( \9742 , \9740 , \9741 );
and \g445796/U$2 ( \9743 , RIdecb4e0_777, \8371 );
and \g445796/U$3 ( \9744 , RIde7d8d0_202, \8335 );
and \g448619/U$2 ( \9745 , RIe16e8e8_2635, \8414 );
and \g448619/U$3 ( \9746 , \8407 , RIde97988_329);
and \g448619/U$4 ( \9747 , RIdece1e0_809, \8383 );
nor \g448619/U$1 ( \9748 , \9745 , \9746 , \9747 );
and \g451004/U$2 ( \9749 , \8356 , RIdf1d7b8_1712);
and \g451004/U$3 ( \9750 , RIe143ee0_2150, \8359 );
nor \g451004/U$1 ( \9751 , \9749 , \9750 );
and \g454441/U$2 ( \9752 , \8313 , RIdf2cf38_1888);
and \g454441/U$3 ( \9753 , RIdf388d8_2020, \8323 );
nor \g454441/U$1 ( \9754 , \9752 , \9753 );
not \g449646/U$3 ( \9755 , \9754 );
not \g449646/U$4 ( \9756 , \8347 );
and \g449646/U$2 ( \9757 , \9755 , \9756 );
and \g449646/U$5 ( \9758 , \8351 , RIded0ee0_841);
nor \g449646/U$1 ( \9759 , \9757 , \9758 );
and \g451002/U$2 ( \9760 , \8378 , RIe15a6e0_2406);
and \g451002/U$3 ( \9761 , RIdeb4ce0_521, \8417 );
nor \g451002/U$1 ( \9762 , \9760 , \9761 );
nand \g447522/U$1 ( \9763 , \9748 , \9751 , \9759 , \9762 );
nor \g445796/U$1 ( \9764 , \9743 , \9744 , \9763 );
and \g450996/U$2 ( \9765 , \8340 , RIdf00eb0_1387);
and \g450996/U$3 ( \9766 , RIdec87e0_745, \8404 );
nor \g450996/U$1 ( \9767 , \9765 , \9766 );
nand \g445531/U$1 ( \9768 , \9742 , \9764 , \9767 );
and \g444873/U$2 ( \9769 , \9768 , \9010 );
and \g448615/U$2 ( \9770 , RIfcacc70_6988, \8373 );
and \g448615/U$3 ( \9771 , \8383 , RIfc69a10_6224);
and \g448615/U$4 ( \9772 , RIfc9bba0_6794, \8488 );
nor \g448615/U$1 ( \9773 , \9770 , \9771 , \9772 );
and \g450988/U$2 ( \9774 , \8335 , RIded34d8_868);
and \g450988/U$3 ( \9775 , RIded9e50_943, \8340 );
nor \g450988/U$1 ( \9776 , \9774 , \9775 );
and \g450986/U$2 ( \9777 , \8404 , RIfccbfa8_7343);
and \g450986/U$3 ( \9778 , RIfcc9848_7315, \8351 );
nor \g450986/U$1 ( \9779 , \9777 , \9778 );
and \g454559/U$2 ( \9780 , \8313 , RIfe887b8_7897);
and \g454559/U$3 ( \9781 , RIded7858_916, \8323 );
nor \g454559/U$1 ( \9782 , \9780 , \9781 );
not \g454558/U$1 ( \9783 , \9782 );
and \g449641/U$2 ( \9784 , \9783 , \8316 );
and \g449641/U$3 ( \9785 , RIfc84590_6528, \8359 );
nor \g449641/U$1 ( \9786 , \9784 , \9785 );
nand \g448148/U$1 ( \9787 , \9773 , \9776 , \9779 , \9786 );
and \g444873/U$3 ( \9788 , \8482 , \9787 );
nor \g444873/U$1 ( \9789 , \9769 , \9788 );
and \g446595/U$2 ( \9790 , \8964 , RIdee31f8_1048);
and \g446595/U$3 ( \9791 , RIdee4f80_1069, \8966 );
nor \g446595/U$1 ( \9792 , \9790 , \9791 );
and \g446596/U$2 ( \9793 , \8521 , RIfc47168_5831);
and \g446596/U$3 ( \9794 , RIee21b38_4842, \8525 );
nor \g446596/U$1 ( \9795 , \9793 , \9794 );
and \g446597/U$2 ( \9796 , \8974 , RIdedee78_1000);
and \g446597/U$3 ( \9797 , RIdee1038_1024, \8976 );
nor \g446597/U$1 ( \9798 , \9796 , \9797 );
nand \g444561/U$1 ( \9799 , \9789 , \9792 , \9795 , \9798 );
and \g445781/U$2 ( \9800 , RIee29158_4926, \8373 );
and \g445781/U$3 ( \9801 , RIdf19870_1667, \8335 );
and \g448600/U$2 ( \9802 , RIfc63368_6151, \8523 );
and \g448600/U$3 ( \9803 , \8488 , RIfc69fb0_6228);
and \g448600/U$4 ( \9804 , RIee2a670_4941, \8383 );
nor \g448600/U$1 ( \9805 , \9802 , \9803 , \9804 );
and \g450929/U$2 ( \9806 , \8356 , RIfc623f0_6140);
and \g450929/U$3 ( \9807 , RIfcad918_6997, \8359 );
nor \g450929/U$1 ( \9808 , \9806 , \9807 );
and \g454699/U$2 ( \9809 , \8313 , RIdf26890_1815);
and \g454699/U$3 ( \9810 , RIdf28618_1836, \8323 );
nor \g454699/U$1 ( \9811 , \9809 , \9810 );
not \g449626/U$3 ( \9812 , \9811 );
not \g449626/U$4 ( \9813 , \8376 );
and \g449626/U$2 ( \9814 , \9812 , \9813 );
and \g449626/U$5 ( \9815 , \8351 , RIee2bfc0_4959);
nor \g449626/U$1 ( \9816 , \9814 , \9815 );
and \g450928/U$2 ( \9817 , \8378 , RIdf24dd8_1796);
and \g450928/U$3 ( \9818 , RIdf2a7d8_1860, \8417 );
nor \g450928/U$1 ( \9819 , \9817 , \9818 );
nand \g447505/U$1 ( \9820 , \9805 , \9808 , \9816 , \9819 );
nor \g445781/U$1 ( \9821 , \9800 , \9801 , \9820 );
and \g450921/U$2 ( \9822 , \8340 , RIfc60938_6121);
and \g450921/U$3 ( \9823 , RIee27f10_4913, \8404 );
nor \g450921/U$1 ( \9824 , \9822 , \9823 );
and \g450922/U$2 ( \9825 , \8317 , RIfcba500_7142);
and \g450922/U$3 ( \9826 , RIdf1ff18_1740, \8326 );
nor \g450922/U$1 ( \9827 , \9825 , \9826 );
and \g444987/U$2 ( \9828 , \9821 , \9824 , \9827 );
nor \g444987/U$1 ( \9829 , \9828 , \8621 );
and \g445784/U$2 ( \9830 , RIdf11cb0_1579, \8371 );
and \g445784/U$3 ( \9831 , RIdeea6b0_1131, \8335 );
and \g448604/U$2 ( \9832 , RIdef87b0_1291, \8523 );
and \g448604/U$3 ( \9833 , \8486 , RIdefb4b0_1323);
and \g448604/U$4 ( \9834 , RIdf149b0_1611, \8383 );
nor \g448604/U$1 ( \9835 , \9832 , \9833 , \9834 );
and \g450945/U$2 ( \9836 , \8356 , RIdef5ab0_1259);
and \g450945/U$3 ( \9837 , RIdefe1b0_1355, \8359 );
nor \g450945/U$1 ( \9838 , \9836 , \9837 );
and \g455277/U$2 ( \9839 , \8313 , RIdf068b0_1451);
and \g455277/U$3 ( \9840 , RIdf095b0_1483, \8323 );
nor \g455277/U$1 ( \9841 , \9839 , \9840 );
not \g449630/U$3 ( \9842 , \9841 );
not \g449630/U$4 ( \9843 , \8376 );
and \g449630/U$2 ( \9844 , \9842 , \9843 );
and \g449630/U$5 ( \9845 , \8351 , RIdf176b0_1643);
nor \g449630/U$1 ( \9846 , \9844 , \9845 );
and \g450943/U$2 ( \9847 , \8378 , RIdf03bb0_1419);
and \g450943/U$3 ( \9848 , RIdf0c2b0_1515, \8417 );
nor \g450943/U$1 ( \9849 , \9847 , \9848 );
nand \g447508/U$1 ( \9850 , \9835 , \9838 , \9846 , \9849 );
nor \g445784/U$1 ( \9851 , \9830 , \9831 , \9850 );
and \g450937/U$2 ( \9852 , \8340 , RIdef2db0_1227);
and \g450937/U$3 ( \9853 , RIdf0efb0_1547, \8404 );
nor \g450937/U$1 ( \9854 , \9852 , \9853 );
and \g450938/U$2 ( \9855 , \8319 , RIdeed3b0_1163);
and \g450938/U$3 ( \9856 , RIdef00b0_1195, \8326 );
nor \g450938/U$1 ( \9857 , \9855 , \9856 );
and \g444988/U$2 ( \9858 , \9851 , \9854 , \9857 );
nor \g444988/U$1 ( \9859 , \9858 , \8477 );
or \g444375/U$1 ( \9860 , \9739 , \9799 , \9829 , \9859 );
and \g445774/U$2 ( \9861 , RIe15d3e0_2438, \8407 );
and \g445774/U$3 ( \9862 , RIe154ce0_2342, \8378 );
and \g448589/U$2 ( \9863 , RIe1498e0_2214, \8319 );
and \g448589/U$3 ( \9864 , \8326 , RIe14c5e0_2246);
and \g448589/U$4 ( \9865 , RIe151fe0_2310, \8488 );
nor \g448589/U$1 ( \9866 , \9863 , \9864 , \9865 );
and \g450898/U$2 ( \9867 , \8335 , RIe146be0_2182);
and \g450898/U$3 ( \9868 , RIfcc0338_7209, \8340 );
nor \g450898/U$1 ( \9869 , \9867 , \9868 );
and \g450896/U$2 ( \9870 , \8404 , RIe1600e0_2470);
and \g450896/U$3 ( \9871 , RIe165ae0_2534, \8351 );
nor \g450896/U$1 ( \9872 , \9870 , \9871 );
and \g455324/U$2 ( \9873 , \8313 , RIfe88a88_7899);
and \g455324/U$3 ( \9874 , RIe162de0_2502, \8323 );
nor \g455324/U$1 ( \9875 , \9873 , \9874 );
not \g449615/U$3 ( \9876 , \9875 );
not \g449615/U$4 ( \9877 , \8328 );
and \g449615/U$2 ( \9878 , \9876 , \9877 );
and \g449615/U$5 ( \9879 , \8359 , RIfc698a8_6223);
nor \g449615/U$1 ( \9880 , \9878 , \9879 );
nand \g447497/U$1 ( \9881 , \9866 , \9869 , \9872 , \9880 );
nor \g445774/U$1 ( \9882 , \9861 , \9862 , \9881 );
and \g450890/U$2 ( \9883 , \8356 , RIe14f2e0_2278);
and \g450890/U$3 ( \9884 , RIfcc9140_7310, \8417 );
nor \g450890/U$1 ( \9885 , \9883 , \9884 );
and \g450887/U$2 ( \9886 , \8531 , RIee35098_5062);
and \g450887/U$3 ( \9887 , RIe1579e0_2374, \8412 );
nor \g450887/U$1 ( \9888 , \9886 , \9887 );
and \g444982/U$2 ( \9889 , \9882 , \9885 , \9888 );
nor \g444982/U$1 ( \9890 , \9889 , \8368 );
and \g445778/U$2 ( \9891 , RIdf3d090_2071, \8414 );
and \g445778/U$3 ( \9892 , RIe1414b0_2120, \8417 );
and \g448595/U$2 ( \9893 , RIfe88920_7898, \8319 );
and \g448595/U$3 ( \9894 , \8326 , RIdf338b0_1963);
and \g448595/U$4 ( \9895 , RIfc7d7e0_6450, \8488 );
nor \g448595/U$1 ( \9896 , \9893 , \9894 , \9895 );
and \g450913/U$2 ( \9897 , \8335 , RIdf2f800_1917);
and \g450913/U$3 ( \9898 , RIdf35ea8_1990, \8340 );
nor \g450913/U$1 ( \9899 , \9897 , \9898 );
and \g450911/U$2 ( \9900 , \8404 , RIfcc4f28_7263);
and \g450911/U$3 ( \9901 , RIfc88208_6571, \8351 );
nor \g450911/U$1 ( \9902 , \9900 , \9901 );
and \g454569/U$2 ( \9903 , \8313 , RIfc81f98_6501);
and \g454569/U$3 ( \9904 , RIfc85670_6540, \8323 );
nor \g454569/U$1 ( \9905 , \9903 , \9904 );
not \g449622/U$3 ( \9906 , \9905 );
not \g449622/U$4 ( \9907 , \8328 );
and \g449622/U$2 ( \9908 , \9906 , \9907 );
and \g449622/U$5 ( \9909 , \8359 , RIfcd2920_7418);
nor \g449622/U$1 ( \9910 , \9908 , \9909 );
nand \g447501/U$1 ( \9911 , \9896 , \9899 , \9902 , \9910 );
nor \g445778/U$1 ( \9912 , \9891 , \9892 , \9911 );
and \g450906/U$2 ( \9913 , \8378 , RIdf3aa98_2044);
and \g450906/U$3 ( \9914 , RIfc49760_5858, \8531 );
nor \g450906/U$1 ( \9915 , \9913 , \9914 );
and \g450908/U$2 ( \9916 , \8356 , RIfce5a48_7635);
and \g450908/U$3 ( \9917 , RIe13f188_2095, \8407 );
nor \g450908/U$1 ( \9918 , \9916 , \9917 );
and \g444986/U$2 ( \9919 , \9912 , \9915 , \9918 );
nor \g444986/U$1 ( \9920 , \9919 , \8422 );
or \g444240/U$1 ( \9921 , \9860 , \9890 , \9920 );
_DC \g24ce/U$1 ( \9922 , \9921 , \8654 );
and \g453255/U$2 ( \9923 , \8326 , RIdee7848_1098);
and \g453255/U$3 ( \9924 , RIdec8678_744, \8404 );
nor \g453255/U$1 ( \9925 , \9923 , \9924 );
and \g446308/U$2 ( \9926 , RIdecb378_776, \8373 );
and \g446308/U$3 ( \9927 , RIdedc5b0_971, \8319 );
and \g449280/U$2 ( \9928 , RIdf2cdd0_1887, \8531 );
and \g449280/U$3 ( \9929 , \8488 , RIdf38770_2019);
and \g449280/U$4 ( \9930 , RIdece078_808, \8330 );
nor \g449280/U$1 ( \9931 , \9928 , \9929 , \9930 );
and \g453264/U$2 ( \9932 , \8356 , RIdf1d650_1711);
and \g453264/U$3 ( \9933 , RIe143d78_2149, \8359 );
nor \g453264/U$1 ( \9934 , \9932 , \9933 );
and \g455303/U$2 ( \9935 , \8313 , RIe16e780_2634);
and \g455303/U$3 ( \9936 , RIde97640_328, \8323 );
nor \g455303/U$1 ( \9937 , \9935 , \9936 );
not \g450296/U$3 ( \9938 , \9937 );
not \g450296/U$4 ( \9939 , \8376 );
and \g450296/U$2 ( \9940 , \9938 , \9939 );
and \g450296/U$5 ( \9941 , \8351 , RIded0d78_840);
nor \g450296/U$1 ( \9942 , \9940 , \9941 );
and \g453262/U$2 ( \9943 , \8378 , RIe15a578_2405);
and \g453262/U$3 ( \9944 , RIdeb4b78_520, \8417 );
nor \g453262/U$1 ( \9945 , \9943 , \9944 );
nand \g447873/U$1 ( \9946 , \9931 , \9934 , \9942 , \9945 );
nor \g446308/U$1 ( \9947 , \9926 , \9927 , \9946 );
and \g453259/U$2 ( \9948 , \8335 , RIde7d588_201);
and \g453259/U$3 ( \9949 , RIdf00d48_1386, \8340 );
nor \g453259/U$1 ( \9950 , \9948 , \9949 );
nand \g445654/U$1 ( \9951 , \9925 , \9947 , \9950 );
and \g444883/U$2 ( \9952 , \9951 , \9010 );
and \g449275/U$2 ( \9953 , RIfc97af0_6748, \8371 );
and \g449275/U$3 ( \9954 , \8383 , RIfc7cb38_6441);
and \g449275/U$4 ( \9955 , RIfcc2930_7236, \8486 );
nor \g449275/U$1 ( \9956 , \9953 , \9954 , \9955 );
and \g453248/U$2 ( \9957 , \8335 , RIded3370_867);
and \g453248/U$3 ( \9958 , RIded9ce8_942, \8340 );
nor \g453248/U$1 ( \9959 , \9957 , \9958 );
and \g453247/U$2 ( \9960 , \8404 , RIfcb3e58_7069);
and \g453247/U$3 ( \9961 , RIfcd9130_7492, \8351 );
nor \g453247/U$1 ( \9962 , \9960 , \9961 );
and \g454508/U$2 ( \9963 , \8313 , RIded5968_894);
and \g454508/U$3 ( \9964 , RIded76f0_915, \8323 );
nor \g454508/U$1 ( \9965 , \9963 , \9964 );
not \g454507/U$1 ( \9966 , \9965 );
and \g450292/U$2 ( \9967 , \9966 , \8316 );
and \g450292/U$3 ( \9968 , RIfc97dc0_6750, \8359 );
nor \g450292/U$1 ( \9969 , \9967 , \9968 );
nand \g448222/U$1 ( \9970 , \9956 , \9959 , \9962 , \9969 );
and \g444883/U$3 ( \9971 , \8482 , \9970 );
nor \g444883/U$1 ( \9972 , \9952 , \9971 );
and \g447076/U$2 ( \9973 , \8964 , RIdee3090_1047);
and \g447076/U$3 ( \9974 , RIdee4e18_1068, \8966 );
nor \g447076/U$1 ( \9975 , \9973 , \9974 );
and \g447077/U$2 ( \9976 , \8521 , RIfc7c868_6439);
and \g447077/U$3 ( \9977 , RIfcd9298_7493, \8525 );
nor \g447077/U$1 ( \9978 , \9976 , \9977 );
and \g447078/U$2 ( \9979 , \8974 , RIfe88380_7894);
and \g447078/U$3 ( \9980 , RIdee0ed0_1023, \8976 );
nor \g447078/U$1 ( \9981 , \9979 , \9980 );
nand \g444647/U$1 ( \9982 , \9972 , \9975 , \9978 , \9981 );
and \g449266/U$2 ( \9983 , RIfc8c150_6616, \8531 );
and \g449266/U$3 ( \9984 , \8488 , RIfcbbb80_7158);
and \g449266/U$4 ( \9985 , RIfcc38a8_7247, \8383 );
nor \g449266/U$1 ( \9986 , \9983 , \9984 , \9985 );
and \g453218/U$2 ( \9987 , \8356 , RIfcbbfb8_7161);
and \g453218/U$3 ( \9988 , RIde82100_224, \8359 );
nor \g453218/U$1 ( \9989 , \9987 , \9988 );
and \g455282/U$2 ( \9990 , \8313 , RIde8a440_264);
and \g455282/U$3 ( \9991 , RIde8e298_283, \8323 );
nor \g455282/U$1 ( \9992 , \9990 , \9991 );
not \g450283/U$3 ( \9993 , \9992 );
not \g450283/U$4 ( \9994 , \8376 );
and \g450283/U$2 ( \9995 , \9993 , \9994 );
and \g450283/U$5 ( \9996 , \8351 , RIfc8b070_6604);
nor \g450283/U$1 ( \9997 , \9995 , \9996 );
and \g453216/U$2 ( \9998 , \8378 , RIde862a0_244);
and \g453216/U$3 ( \9999 , RIde91a60_300, \8417 );
nor \g453216/U$1 ( \10000 , \9998 , \9999 );
nand \g447866/U$1 ( \10001 , \9986 , \9989 , \9997 , \10000 );
and \g444688/U$2 ( \10002 , \10001 , \9700 );
and \g446302/U$2 ( \10003 , RIfc8aad0_6600, \8371 );
and \g446302/U$3 ( \10004 , RIdea4840_392, \8319 );
and \g449270/U$2 ( \10005 , RIdeba578_584, \8414 );
and \g449270/U$3 ( \10006 , \8407 , RIdebd278_616);
and \g449270/U$4 ( \10007 , RIdec2c78_680, \8383 );
nor \g449270/U$1 ( \10008 , \10005 , \10006 , \10007 );
and \g453235/U$2 ( \10009 , \8356 , RIdeaf178_456);
and \g453235/U$3 ( \10010 , RIfc40e80_5764, \8359 );
nor \g453235/U$1 ( \10011 , \10009 , \10010 );
and \g455298/U$2 ( \10012 , \8313 , RIfcdaeb8_7513);
and \g455298/U$3 ( \10013 , RIdeb1e78_488, \8323 );
nor \g455298/U$1 ( \10014 , \10012 , \10013 );
not \g450288/U$3 ( \10015 , \10014 );
not \g450288/U$4 ( \10016 , \8347 );
and \g450288/U$2 ( \10017 , \10015 , \10016 );
and \g450288/U$5 ( \10018 , \8351 , RIdec5978_712);
nor \g450288/U$1 ( \10019 , \10017 , \10018 );
and \g453234/U$2 ( \10020 , \8378 , RIdeb7878_552);
and \g453234/U$3 ( \10021 , RIfc8ac38_6601, \8417 );
nor \g453234/U$1 ( \10022 , \10020 , \10021 );
nand \g447868/U$1 ( \10023 , \10008 , \10011 , \10019 , \10022 );
nor \g446302/U$1 ( \10024 , \10003 , \10004 , \10023 );
and \g453227/U$2 ( \10025 , \8335 , RIde9df40_360);
and \g453227/U$3 ( \10026 , RIee1dbf0_4797, \8340 );
nor \g453227/U$1 ( \10027 , \10025 , \10026 );
and \g453224/U$2 ( \10028 , \8326 , RIdeab140_424);
and \g453224/U$3 ( \10029 , RIdebff78_648, \8404 );
nor \g453224/U$1 ( \10030 , \10028 , \10029 );
and \g445364/U$2 ( \10031 , \10024 , \10027 , \10030 );
nor \g445364/U$1 ( \10032 , \10031 , \8589 );
nor \g444688/U$1 ( \10033 , \10002 , \10032 );
nor \g448275/U$1 ( \10034 , \8558 , \8325 );
and \g447070/U$2 ( \10035 , \10034 , RIe16bbe8_2603);
nor \g448291/U$1 ( \10036 , \8558 , \8516 );
and \g447070/U$3 ( \10037 , RIfc54458_5981, \10036 );
nor \g447070/U$1 ( \10038 , \10035 , \10037 );
nor \g448258/U$1 ( \10039 , \8558 , \8425 );
and \g447069/U$2 ( \10040 , \10039 , RIfcbb8b0_7156);
nor \g448303/U$1 ( \10041 , \8558 , \8372 );
and \g447069/U$3 ( \10042 , RIfc807b0_6484, \10041 );
nor \g447069/U$1 ( \10043 , \10040 , \10042 );
nor \g448257/U$1 ( \10044 , \8558 , \8508 );
and \g447072/U$2 ( \10045 , \10044 , RIe168240_2562);
nor \g448273/U$1 ( \10046 , \8558 , \8318 );
and \g447072/U$3 ( \10047 , RIfc8c2b8_6617, \10046 );
nor \g447072/U$1 ( \10048 , \10045 , \10047 );
nand \g444524/U$1 ( \10049 , \10033 , \10038 , \10043 , \10048 );
and \g446292/U$2 ( \10050 , RIe15d278_2437, \8407 );
and \g446292/U$3 ( \10051 , RIe154b78_2341, \8378 );
and \g449258/U$2 ( \10052 , RIee37960_5091, \8373 );
and \g449258/U$3 ( \10053 , \8330 , RIe162c78_2501);
and \g449258/U$4 ( \10054 , RIe151e78_2309, \8486 );
nor \g449258/U$1 ( \10055 , \10052 , \10053 , \10054 );
and \g453185/U$2 ( \10056 , \8335 , RIe146a78_2181);
and \g453185/U$3 ( \10057 , RIfc56ff0_6012, \8340 );
nor \g453185/U$1 ( \10058 , \10056 , \10057 );
and \g453184/U$2 ( \10059 , \8404 , RIe15ff78_2469);
and \g453184/U$3 ( \10060 , RIe165978_2533, \8351 );
nor \g453184/U$1 ( \10061 , \10059 , \10060 );
and \g455281/U$2 ( \10062 , \8313 , RIe149778_2213);
and \g455281/U$3 ( \10063 , RIe14c478_2245, \8323 );
nor \g455281/U$1 ( \10064 , \10062 , \10063 );
not \g455280/U$1 ( \10065 , \10064 );
and \g450274/U$2 ( \10066 , \10065 , \8316 );
and \g450274/U$3 ( \10067 , RIfc8e5e0_6642, \8359 );
nor \g450274/U$1 ( \10068 , \10066 , \10067 );
nand \g448221/U$1 ( \10069 , \10055 , \10058 , \10061 , \10068 );
nor \g446292/U$1 ( \10070 , \10050 , \10051 , \10069 );
and \g453178/U$2 ( \10071 , \8356 , RIe14f178_2277);
and \g453178/U$3 ( \10072 , RIfcd6b38_7465, \8417 );
nor \g453178/U$1 ( \10073 , \10071 , \10072 );
and \g453175/U$2 ( \10074 , \8523 , RIfcb4290_7072);
and \g453175/U$3 ( \10075 , RIe157878_2373, \8414 );
nor \g453175/U$1 ( \10076 , \10074 , \10075 );
and \g445358/U$2 ( \10077 , \10070 , \10073 , \10076 );
nor \g445358/U$1 ( \10078 , \10077 , \8368 );
and \g446296/U$2 ( \10079 , RIe13f020_2094, \8407 );
and \g446296/U$3 ( \10080 , RIdf3a930_2043, \8378 );
and \g449262/U$2 ( \10081 , RIdf316f0_1939, \8319 );
and \g449262/U$3 ( \10082 , \8326 , RIfe88218_7893);
and \g449262/U$4 ( \10083 , RIfc56780_6006, \8486 );
nor \g449262/U$1 ( \10084 , \10081 , \10082 , \10083 );
and \g453205/U$2 ( \10085 , \8335 , RIdf2f698_1916);
and \g453205/U$3 ( \10086 , RIdf35d40_1989, \8340 );
nor \g453205/U$1 ( \10087 , \10085 , \10086 );
and \g453204/U$2 ( \10088 , \8404 , RIee31420_5019);
and \g453204/U$3 ( \10089 , RIee346c0_5055, \8351 );
nor \g453204/U$1 ( \10090 , \10088 , \10089 );
and \g454612/U$2 ( \10091 , \8313 , RIee32398_5030);
and \g454612/U$3 ( \10092 , RIee335e0_5043, \8323 );
nor \g454612/U$1 ( \10093 , \10091 , \10092 );
not \g450279/U$3 ( \10094 , \10093 );
not \g450279/U$4 ( \10095 , \8328 );
and \g450279/U$2 ( \10096 , \10094 , \10095 );
and \g450279/U$5 ( \10097 , \8359 , RIfce3e28_7615);
nor \g450279/U$1 ( \10098 , \10096 , \10097 );
nand \g447863/U$1 ( \10099 , \10084 , \10087 , \10090 , \10098 );
nor \g446296/U$1 ( \10100 , \10079 , \10080 , \10099 );
and \g453200/U$2 ( \10101 , \8356 , RIfce2eb0_7604);
and \g453200/U$3 ( \10102 , RIe141348_2119, \8417 );
nor \g453200/U$1 ( \10103 , \10101 , \10102 );
and \g453196/U$2 ( \10104 , \8531 , RIfcb4128_7071);
and \g453196/U$3 ( \10105 , RIfec16f8_8321, \8414 );
nor \g453196/U$1 ( \10106 , \10104 , \10105 );
and \g445362/U$2 ( \10107 , \10100 , \10103 , \10106 );
nor \g445362/U$1 ( \10108 , \10107 , \8422 );
or \g444372/U$1 ( \10109 , \9982 , \10049 , \10078 , \10108 );
and \g446286/U$2 ( \10110 , RIdf284b0_1835, \8409 );
and \g446286/U$3 ( \10111 , RIdf24c70_1795, \8378 );
and \g449249/U$2 ( \10112 , RIfcd62c8_7459, \8371 );
and \g449249/U$3 ( \10113 , \8383 , RIfce4260_7618);
and \g449249/U$4 ( \10114 , RIfcc31a0_7242, \8488 );
nor \g449249/U$1 ( \10115 , \10112 , \10113 , \10114 );
and \g451869/U$2 ( \10116 , \8335 , RIdf19708_1666);
and \g451869/U$3 ( \10117 , RIfce2a78_7601, \8340 );
nor \g451869/U$1 ( \10118 , \10116 , \10117 );
and \g453148/U$2 ( \10119 , \8404 , RIfce9990_7680);
and \g453148/U$3 ( \10120 , RIfc7f9a0_6474, \8351 );
nor \g453148/U$1 ( \10121 , \10119 , \10120 );
and \g455262/U$2 ( \10122 , \8313 , RIfcc6e18_7285);
and \g455262/U$3 ( \10123 , RIdf1fdb0_1739, \8323 );
nor \g455262/U$1 ( \10124 , \10122 , \10123 );
not \g455261/U$1 ( \10125 , \10124 );
and \g450264/U$2 ( \10126 , \10125 , \8316 );
and \g450264/U$3 ( \10127 , RIfc7ecf8_6465, \8359 );
nor \g450264/U$1 ( \10128 , \10126 , \10127 );
nand \g448220/U$1 ( \10129 , \10115 , \10118 , \10121 , \10128 );
nor \g446286/U$1 ( \10130 , \10110 , \10111 , \10129 );
and \g453143/U$2 ( \10131 , \8356 , RIfc46e98_5829);
and \g453143/U$3 ( \10132 , RIdf2a670_1859, \8417 );
nor \g453143/U$1 ( \10133 , \10131 , \10132 );
and \g453142/U$2 ( \10134 , \8531 , RIfc99008_6763);
and \g453142/U$3 ( \10135 , RIdf26728_1814, \8412 );
nor \g453142/U$1 ( \10136 , \10134 , \10135 );
and \g445355/U$2 ( \10137 , \10130 , \10133 , \10136 );
nor \g445355/U$1 ( \10138 , \10137 , \8621 );
and \g446289/U$2 ( \10139 , RIdf06748_1450, \8412 );
and \g446289/U$3 ( \10140 , RIdf0c148_1514, \8417 );
and \g449254/U$2 ( \10141 , RIdeeff48_1194, \8326 );
and \g449254/U$3 ( \10142 , \8523 , RIdef8648_1290);
and \g449254/U$4 ( \10143 , RIdefb348_1322, \8488 );
nor \g449254/U$1 ( \10144 , \10141 , \10142 , \10143 );
and \g454660/U$2 ( \10145 , \8313 , RIdf11b48_1578);
and \g454660/U$3 ( \10146 , RIdf14848_1610, \8323 );
nor \g454660/U$1 ( \10147 , \10145 , \10146 );
not \g450270/U$3 ( \10148 , \10147 );
not \g450270/U$4 ( \10149 , \8328 );
and \g450270/U$2 ( \10150 , \10148 , \10149 );
and \g450270/U$5 ( \10151 , \8340 , RIdef2c48_1226);
nor \g450270/U$1 ( \10152 , \10150 , \10151 );
and \g453164/U$2 ( \10153 , \8404 , RIdf0ee48_1546);
and \g453164/U$3 ( \10154 , RIdf17548_1642, \8351 );
nor \g453164/U$1 ( \10155 , \10153 , \10154 );
and \g453166/U$2 ( \10156 , \8356 , RIdef5948_1258);
and \g453166/U$3 ( \10157 , RIdefe048_1354, \8359 );
nor \g453166/U$1 ( \10158 , \10156 , \10157 );
nand \g447860/U$1 ( \10159 , \10144 , \10152 , \10155 , \10158 );
nor \g446289/U$1 ( \10160 , \10139 , \10140 , \10159 );
and \g453159/U$2 ( \10161 , \8335 , RIdeea548_1130);
and \g453159/U$3 ( \10162 , RIdf09448_1482, \8407 );
nor \g453159/U$1 ( \10163 , \10161 , \10162 );
and \g453158/U$2 ( \10164 , \8319 , RIdeed248_1162);
and \g453158/U$3 ( \10165 , RIdf03a48_1418, \8378 );
nor \g453158/U$1 ( \10166 , \10164 , \10165 );
and \g445356/U$2 ( \10167 , \10160 , \10163 , \10166 );
nor \g445356/U$1 ( \10168 , \10167 , \8477 );
or \g444254/U$1 ( \10169 , \10109 , \10138 , \10168 );
_DC \g2553/U$1 ( \10170 , \10169 , \8654 );
and \g447116/U$2 ( \10171 , \9299 , RIdf2f530_1915);
and \g447116/U$3 ( \10172 , RIdf31588_1938, \9301 );
nor \g447116/U$1 ( \10173 , \10171 , \10172 );
and \g446357/U$2 ( \10174 , RIfccf0e0_7378, \8486 );
and \g446357/U$3 ( \10175 , RIfcc99b0_7316, \8359 );
and \g449341/U$2 ( \10176 , RIdf3cf28_2070, \8414 );
and \g449341/U$3 ( \10177 , \8409 , RIfe87570_7884);
and \g449341/U$4 ( \10178 , RIdf33748_1962, \8326 );
nor \g449341/U$1 ( \10179 , \10176 , \10177 , \10178 );
and \g455337/U$2 ( \10180 , \8313 , RIfc71b70_6316);
and \g455337/U$3 ( \10181 , RIee33478_5042, \8323 );
nor \g455337/U$1 ( \10182 , \10180 , \10181 );
not \g450360/U$3 ( \10183 , \10182 );
not \g450360/U$4 ( \10184 , \8328 );
and \g450360/U$2 ( \10185 , \10183 , \10184 );
and \g450360/U$5 ( \10186 , \8340 , RIdf35bd8_1988);
nor \g450360/U$1 ( \10187 , \10185 , \10186 );
and \g453485/U$2 ( \10188 , \8404 , RIee312b8_5018);
and \g453485/U$3 ( \10189 , RIfc62288_6139, \8351 );
nor \g453485/U$1 ( \10190 , \10188 , \10189 );
and \g453488/U$2 ( \10191 , \8378 , RIfe87408_7883);
and \g453488/U$3 ( \10192 , RIe1411e0_2118, \8417 );
nor \g453488/U$1 ( \10193 , \10191 , \10192 );
nand \g447910/U$1 ( \10194 , \10179 , \10187 , \10190 , \10193 );
nor \g446357/U$1 ( \10195 , \10174 , \10175 , \10194 );
not \g444870/U$3 ( \10196 , \10195 );
not \g444870/U$4 ( \10197 , \8422 );
and \g444870/U$2 ( \10198 , \10196 , \10197 );
and \g446365/U$2 ( \10199 , RIfc3f3c8_5745, \8359 );
and \g446365/U$3 ( \10200 , RIe146910_2180, \8335 );
and \g449345/U$2 ( \10201 , RIe14c310_2244, \8326 );
and \g449345/U$3 ( \10202 , \8371 , RIee377f8_5090);
and \g449345/U$4 ( \10203 , RIe162b10_2500, \8330 );
nor \g449345/U$1 ( \10204 , \10201 , \10202 , \10203 );
and \g454935/U$2 ( \10205 , \8313 , RIe157710_2372);
and \g454935/U$3 ( \10206 , RIe15d110_2436, \8323 );
nor \g454935/U$1 ( \10207 , \10205 , \10206 );
not \g450364/U$3 ( \10208 , \10207 );
not \g450364/U$4 ( \10209 , \8376 );
and \g450364/U$2 ( \10210 , \10208 , \10209 );
and \g450364/U$5 ( \10211 , \8340 , RIfc4a2a0_5866);
nor \g450364/U$1 ( \10212 , \10210 , \10211 );
and \g453508/U$2 ( \10213 , \8404 , RIe15fe10_2468);
and \g453508/U$3 ( \10214 , RIe165810_2532, \8351 );
nor \g453508/U$1 ( \10215 , \10213 , \10214 );
and \g453509/U$2 ( \10216 , \8378 , RIe154a10_2340);
and \g453509/U$3 ( \10217 , RIee36448_5076, \8417 );
nor \g453509/U$1 ( \10218 , \10216 , \10217 );
nand \g447914/U$1 ( \10219 , \10204 , \10212 , \10215 , \10218 );
nor \g446365/U$1 ( \10220 , \10199 , \10200 , \10219 );
and \g453499/U$2 ( \10221 , \8317 , RIe149610_2212);
and \g453499/U$3 ( \10222 , RIe14f010_2276, \8356 );
nor \g453499/U$1 ( \10223 , \10221 , \10222 );
and \g453497/U$2 ( \10224 , \8523 , RIfcde9c8_7555);
and \g453497/U$3 ( \10225 , RIe151d10_2308, \8488 );
nor \g453497/U$1 ( \10226 , \10224 , \10225 );
and \g445402/U$2 ( \10227 , \10220 , \10223 , \10226 );
nor \g445402/U$1 ( \10228 , \10227 , \8368 );
nor \g444870/U$1 ( \10229 , \10198 , \10228 );
nor \g448408/U$1 ( \10230 , \8422 , \8520 );
and \g447117/U$2 ( \10231 , \10230 , RIfcca220_7322);
nor \g448435/U$1 ( \10232 , \8422 , \8524 );
and \g447117/U$3 ( \10233 , RIfcaeb60_7010, \10232 );
nor \g447117/U$1 ( \10234 , \10231 , \10233 );
nand \g444433/U$1 ( \10235 , \10173 , \10229 , \10234 );
and \g453540/U$2 ( \10236 , \8404 , RIdf0ece0_1545);
and \g453540/U$3 ( \10237 , RIdf065e0_1449, \8412 );
nor \g453540/U$1 ( \10238 , \10236 , \10237 );
and \g446370/U$2 ( \10239 , RIdf119e0_1577, \8373 );
and \g446370/U$3 ( \10240 , RIdf146e0_1609, \8383 );
and \g449356/U$2 ( \10241 , RIdeed0e0_1161, \8317 );
and \g449356/U$3 ( \10242 , \8326 , RIdeefde0_1193);
and \g449356/U$4 ( \10243 , RIdf092e0_1481, \8407 );
nor \g449356/U$1 ( \10244 , \10241 , \10242 , \10243 );
and \g454547/U$2 ( \10245 , \8313 , RIdef84e0_1289);
and \g454547/U$3 ( \10246 , RIdefb1e0_1321, \8323 );
nor \g454547/U$1 ( \10247 , \10245 , \10246 );
not \g450377/U$3 ( \10248 , \10247 );
not \g450377/U$4 ( \10249 , \8347 );
and \g450377/U$2 ( \10250 , \10248 , \10249 );
and \g450377/U$5 ( \10251 , \8417 , RIdf0bfe0_1513);
nor \g450377/U$1 ( \10252 , \10250 , \10251 );
and \g453548/U$2 ( \10253 , \8335 , RIdeea3e0_1129);
and \g453548/U$3 ( \10254 , RIdef2ae0_1225, \8340 );
nor \g453548/U$1 ( \10255 , \10253 , \10254 );
and \g453545/U$2 ( \10256 , \8356 , RIdef57e0_1257);
and \g453545/U$3 ( \10257 , RIdefdee0_1353, \8359 );
nor \g453545/U$1 ( \10258 , \10256 , \10257 );
nand \g447920/U$1 ( \10259 , \10244 , \10252 , \10255 , \10258 );
nor \g446370/U$1 ( \10260 , \10239 , \10240 , \10259 );
and \g453536/U$2 ( \10261 , \8378 , RIdf038e0_1417);
and \g453536/U$3 ( \10262 , RIdf173e0_1641, \8351 );
nor \g453536/U$1 ( \10263 , \10261 , \10262 );
nand \g445672/U$1 ( \10264 , \10238 , \10260 , \10263 );
and \g444799/U$2 ( \10265 , \10264 , \8478 );
and \g449352/U$2 ( \10266 , RIfeaaac0_8258, \8326 );
and \g449352/U$3 ( \10267 , \8371 , RIee23e60_4867);
and \g449352/U$4 ( \10268 , RIfca73d8_6925, \8330 );
nor \g449352/U$1 ( \10269 , \10266 , \10267 , \10268 );
and \g454782/U$2 ( \10270 , \8313 , RIdee0d68_1022);
and \g454782/U$3 ( \10271 , RIdee2f28_1046, \8323 );
nor \g454782/U$1 ( \10272 , \10270 , \10271 );
not \g450370/U$3 ( \10273 , \10272 );
not \g450370/U$4 ( \10274 , \8376 );
and \g450370/U$2 ( \10275 , \10273 , \10274 );
and \g450370/U$5 ( \10276 , \8340 , RIded9b80_941);
nor \g450370/U$1 ( \10277 , \10275 , \10276 );
and \g453524/U$2 ( \10278 , \8404 , RIfce66f0_7644);
and \g453524/U$3 ( \10279 , RIee257b0_4885, \8351 );
nor \g453524/U$1 ( \10280 , \10278 , \10279 );
and \g453525/U$2 ( \10281 , \8378 , RIdeded10_999);
and \g453525/U$3 ( \10282 , RIdee4cb0_1067, \8417 );
nor \g453525/U$1 ( \10283 , \10281 , \10282 );
nand \g447917/U$1 ( \10284 , \10269 , \10277 , \10280 , \10283 );
and \g444799/U$3 ( \10285 , \8482 , \10284 );
nor \g444799/U$1 ( \10286 , \10265 , \10285 );
and \g447120/U$2 ( \10287 , \8509 , RIded3208_866);
and \g447120/U$3 ( \10288 , RIded5800_893, \8511 );
nor \g447120/U$1 ( \10289 , \10287 , \10288 );
nor \g448304/U$1 ( \10290 , \8481 , \8487 );
and \g447121/U$2 ( \10291 , \10290 , RIfce6858_7645);
not \g455434/U$1 ( \10292 , \8359 );
nor \g448261/U$1 ( \10293 , \8481 , \10292 );
and \g447121/U$3 ( \10294 , RIfcca388_7323, \10293 );
nor \g447121/U$1 ( \10295 , \10291 , \10294 );
and \g447122/U$2 ( \10296 , \8521 , RIfcdc970_7532);
and \g447122/U$3 ( \10297 , RIfcceca8_7375, \8525 );
nor \g447122/U$1 ( \10298 , \10296 , \10297 );
nand \g444530/U$1 ( \10299 , \10286 , \10289 , \10295 , \10298 );
and \g446348/U$2 ( \10300 , RIee28ff0_4925, \8371 );
and \g446348/U$3 ( \10301 , RIee2a508_4940, \8383 );
and \g449330/U$2 ( \10302 , RIfcaff10_7024, \8319 );
and \g449330/U$3 ( \10303 , \8326 , RIdf1fc48_1738);
and \g449330/U$4 ( \10304 , RIdf28348_1834, \8409 );
nor \g449330/U$1 ( \10305 , \10302 , \10303 , \10304 );
and \g455203/U$2 ( \10306 , \8313 , RIfc43388_5787);
and \g455203/U$3 ( \10307 , RIfc42578_5777, \8323 );
nor \g455203/U$1 ( \10308 , \10306 , \10307 );
not \g450347/U$3 ( \10309 , \10308 );
not \g450347/U$4 ( \10310 , \8347 );
and \g450347/U$2 ( \10311 , \10309 , \10310 );
and \g450347/U$5 ( \10312 , \8417 , RIdf2a508_1858);
nor \g450347/U$1 ( \10313 , \10311 , \10312 );
and \g453452/U$2 ( \10314 , \8335 , RIdf195a0_1665);
and \g453452/U$3 ( \10315 , RIfcb0078_7025, \8340 );
nor \g453452/U$1 ( \10316 , \10314 , \10315 );
and \g453451/U$2 ( \10317 , \8356 , RIfc745a0_6346);
and \g453451/U$3 ( \10318 , RIfc74708_6347, \8359 );
nor \g453451/U$1 ( \10319 , \10317 , \10318 );
nand \g447902/U$1 ( \10320 , \10305 , \10313 , \10316 , \10319 );
nor \g446348/U$1 ( \10321 , \10300 , \10301 , \10320 );
and \g453446/U$2 ( \10322 , \8378 , RIdf24b08_1794);
and \g453446/U$3 ( \10323 , RIee2be58_4958, \8351 );
nor \g453446/U$1 ( \10324 , \10322 , \10323 );
and \g453447/U$2 ( \10325 , \8404 , RIee27da8_4912);
and \g453447/U$3 ( \10326 , RIdf265c0_1813, \8414 );
nor \g453447/U$1 ( \10327 , \10325 , \10326 );
and \g445398/U$2 ( \10328 , \10321 , \10324 , \10327 );
nor \g445398/U$1 ( \10329 , \10328 , \8621 );
and \g446352/U$2 ( \10330 , RIdf1d4e8_1710, \8356 );
and \g446352/U$3 ( \10331 , RIe143c10_2148, \8359 );
and \g449335/U$2 ( \10332 , RIdee76e0_1097, \8326 );
and \g449335/U$3 ( \10333 , \8373 , RIdecb210_775);
and \g449335/U$4 ( \10334 , RIdecdf10_807, \8330 );
nor \g449335/U$1 ( \10335 , \10332 , \10333 , \10334 );
and \g454210/U$2 ( \10336 , \8313 , RIe16e618_2633);
and \g454210/U$3 ( \10337 , RIde972f8_327, \8323 );
nor \g454210/U$1 ( \10338 , \10336 , \10337 );
not \g450353/U$3 ( \10339 , \10338 );
not \g450353/U$4 ( \10340 , \8376 );
and \g450353/U$2 ( \10341 , \10339 , \10340 );
and \g450353/U$5 ( \10342 , \8340 , RIdf00be0_1385);
nor \g450353/U$1 ( \10343 , \10341 , \10342 );
and \g453468/U$2 ( \10344 , \8404 , RIdec8510_743);
and \g453468/U$3 ( \10345 , RIded0c10_839, \8351 );
nor \g453468/U$1 ( \10346 , \10344 , \10345 );
and \g453472/U$2 ( \10347 , \8378 , RIe15a410_2404);
and \g453472/U$3 ( \10348 , RIdeb4a10_519, \8417 );
nor \g453472/U$1 ( \10349 , \10347 , \10348 );
nand \g447905/U$1 ( \10350 , \10335 , \10343 , \10346 , \10349 );
nor \g446352/U$1 ( \10351 , \10330 , \10331 , \10350 );
and \g453464/U$2 ( \10352 , \8335 , RIde7d240_200);
and \g453464/U$3 ( \10353 , RIdf38608_2018, \8486 );
nor \g453464/U$1 ( \10354 , \10352 , \10353 );
and \g453460/U$2 ( \10355 , \8319 , RIdedc448_970);
and \g453460/U$3 ( \10356 , RIdf2cc68_1886, \8523 );
nor \g453460/U$1 ( \10357 , \10355 , \10356 );
and \g445399/U$2 ( \10358 , \10351 , \10354 , \10357 );
nor \g445399/U$1 ( \10359 , \10358 , \8651 );
or \g444293/U$1 ( \10360 , \10235 , \10299 , \10329 , \10359 );
and \g446340/U$2 ( \10361 , RIfcc16e8_7223, \8523 );
and \g446340/U$3 ( \10362 , RIdeb1d10_487, \8488 );
and \g449320/U$2 ( \10363 , RIdeaadf8_423, \8326 );
and \g449320/U$3 ( \10364 , \8371 , RIfce6f60_7650);
and \g449320/U$4 ( \10365 , RIdec2b10_679, \8383 );
nor \g449320/U$1 ( \10366 , \10363 , \10364 , \10365 );
and \g454178/U$2 ( \10367 , \8313 , RIdeba410_583);
and \g454178/U$3 ( \10368 , RIdebd110_615, \8323 );
nor \g454178/U$1 ( \10369 , \10367 , \10368 );
not \g450339/U$3 ( \10370 , \10369 );
not \g450339/U$4 ( \10371 , \8376 );
and \g450339/U$2 ( \10372 , \10370 , \10371 );
and \g450339/U$5 ( \10373 , \8340 , RIfca4f48_6899);
nor \g450339/U$1 ( \10374 , \10372 , \10373 );
and \g453412/U$2 ( \10375 , \8404 , RIdebfe10_647);
and \g453412/U$3 ( \10376 , RIdec5810_711, \8351 );
nor \g453412/U$1 ( \10377 , \10375 , \10376 );
and \g453413/U$2 ( \10378 , \8378 , RIdeb7710_551);
and \g453413/U$3 ( \10379 , RIfc95228_6719, \8417 );
nor \g453413/U$1 ( \10380 , \10378 , \10379 );
nand \g447894/U$1 ( \10381 , \10366 , \10374 , \10377 , \10380 );
nor \g446340/U$1 ( \10382 , \10361 , \10362 , \10381 );
and \g453405/U$2 ( \10383 , \8335 , RIde9dbf8_359);
and \g453405/U$3 ( \10384 , RIfe879a8_7887, \8359 );
nor \g453405/U$1 ( \10385 , \10383 , \10384 );
and \g453406/U$2 ( \10386 , \8319 , RIdea44f8_391);
and \g453406/U$3 ( \10387 , RIdeaf010_455, \8356 );
nor \g453406/U$1 ( \10388 , \10386 , \10387 );
and \g445390/U$2 ( \10389 , \10382 , \10385 , \10388 );
nor \g445390/U$1 ( \10390 , \10389 , \8589 );
and \g446345/U$2 ( \10391 , RIfcdee00_7558, \8356 );
and \g446345/U$3 ( \10392 , RIfcb0780_7030, \8359 );
and \g449325/U$2 ( \10393 , RIde8a0f8_263, \8412 );
and \g449325/U$3 ( \10394 , \8409 , RIfe876d8_7885);
and \g449325/U$4 ( \10395 , RIe16ba80_2602, \8326 );
nor \g449325/U$1 ( \10396 , \10393 , \10394 , \10395 );
and \g454987/U$2 ( \10397 , \8313 , RIfc95660_6722);
and \g454987/U$3 ( \10398 , RIee1bfd0_4777, \8323 );
nor \g454987/U$1 ( \10399 , \10397 , \10398 );
not \g450342/U$3 ( \10400 , \10399 );
not \g450342/U$4 ( \10401 , \8328 );
and \g450342/U$2 ( \10402 , \10400 , \10401 );
and \g450342/U$5 ( \10403 , \8340 , RIfcd8050_7480);
nor \g450342/U$1 ( \10404 , \10402 , \10403 );
and \g453433/U$2 ( \10405 , \8404 , RIfcee148_7731);
and \g453433/U$3 ( \10406 , RIee1cf48_4788, \8351 );
nor \g453433/U$1 ( \10407 , \10405 , \10406 );
and \g453434/U$2 ( \10408 , \8378 , RIde85f58_243);
and \g453434/U$3 ( \10409 , RIfe87840_7886, \8417 );
nor \g453434/U$1 ( \10410 , \10408 , \10409 );
nand \g447899/U$1 ( \10411 , \10396 , \10404 , \10407 , \10410 );
nor \g446345/U$1 ( \10412 , \10391 , \10392 , \10411 );
and \g453427/U$2 ( \10413 , \8335 , RIe1680d8_2561);
and \g453427/U$3 ( \10414 , RIfcee9b8_7737, \8488 );
nor \g453427/U$1 ( \10415 , \10413 , \10414 );
and \g453426/U$2 ( \10416 , \8319 , RIfca5380_6902);
and \g453426/U$3 ( \10417 , RIfc5f150_6104, \8531 );
nor \g453426/U$1 ( \10418 , \10416 , \10417 );
and \g445393/U$2 ( \10419 , \10412 , \10415 , \10418 );
nor \g445393/U$1 ( \10420 , \10419 , \8558 );
or \g444235/U$1 ( \10421 , \10360 , \10390 , \10420 );
_DC \g25d8/U$1 ( \10422 , \10421 , \8654 );
and \g452222/U$2 ( \10423 , \8326 , RIdee7578_1096);
and \g452222/U$3 ( \10424 , RIdec83a8_742, \8404 );
nor \g452222/U$1 ( \10425 , \10423 , \10424 );
and \g446093/U$2 ( \10426 , RIdecb0a8_774, \8373 );
and \g446093/U$3 ( \10427 , RIdedc2e0_969, \8319 );
and \g448997/U$2 ( \10428 , RIdf2cb00_1885, \8531 );
and \g448997/U$3 ( \10429 , \8488 , RIdf384a0_2017);
and \g448997/U$4 ( \10430 , RIdecdda8_806, \8383 );
nor \g448997/U$1 ( \10431 , \10428 , \10429 , \10430 );
and \g452234/U$2 ( \10432 , \8356 , RIdf1d380_1709);
and \g452234/U$3 ( \10433 , RIe143aa8_2147, \8359 );
nor \g452234/U$1 ( \10434 , \10432 , \10433 );
and \g454761/U$2 ( \10435 , \8313 , RIe16e4b0_2632);
and \g454761/U$3 ( \10436 , RIde96fb0_326, \8323 );
nor \g454761/U$1 ( \10437 , \10435 , \10436 );
not \g450010/U$3 ( \10438 , \10437 );
not \g450010/U$4 ( \10439 , \8376 );
and \g450010/U$2 ( \10440 , \10438 , \10439 );
and \g450010/U$5 ( \10441 , \8351 , RIded0aa8_838);
nor \g450010/U$1 ( \10442 , \10440 , \10441 );
and \g452231/U$2 ( \10443 , \8378 , RIe15a2a8_2403);
and \g452231/U$3 ( \10444 , RIdeb48a8_518, \8417 );
nor \g452231/U$1 ( \10445 , \10443 , \10444 );
nand \g447729/U$1 ( \10446 , \10431 , \10434 , \10442 , \10445 );
nor \g446093/U$1 ( \10447 , \10426 , \10427 , \10446 );
and \g452225/U$2 ( \10448 , \8335 , RIde7cef8_199);
and \g452225/U$3 ( \10449 , RIdf00a78_1384, \8340 );
nor \g452225/U$1 ( \10450 , \10448 , \10449 );
nand \g445598/U$1 ( \10451 , \10425 , \10447 , \10450 );
and \g444877/U$2 ( \10452 , \10451 , \9010 );
and \g448993/U$2 ( \10453 , RIdee0c00_1021, \8414 );
and \g448993/U$3 ( \10454 , \8409 , RIdee2dc0_1045);
and \g448993/U$4 ( \10455 , RIfc61a18_6133, \8383 );
nor \g448993/U$1 ( \10456 , \10453 , \10454 , \10455 );
and \g452214/U$2 ( \10457 , \8356 , RIee21430_4837);
and \g452214/U$3 ( \10458 , RIfc626c0_6142, \8359 );
nor \g452214/U$1 ( \10459 , \10457 , \10458 );
and \g454756/U$2 ( \10460 , \8313 , RIfcb31b0_7060);
and \g454756/U$3 ( \10461 , RIfc738f8_6337, \8323 );
nor \g454756/U$1 ( \10462 , \10460 , \10461 );
not \g450006/U$3 ( \10463 , \10462 );
not \g450006/U$4 ( \10464 , \8347 );
and \g450006/U$2 ( \10465 , \10463 , \10464 );
and \g450006/U$5 ( \10466 , \8351 , RIfc611a8_6127);
nor \g450006/U$1 ( \10467 , \10465 , \10466 );
and \g452211/U$2 ( \10468 , \8378 , RIdedeba8_998);
and \g452211/U$3 ( \10469 , RIdee4b48_1066, \8417 );
nor \g452211/U$1 ( \10470 , \10468 , \10469 );
nand \g447722/U$1 ( \10471 , \10456 , \10459 , \10467 , \10470 );
and \g444877/U$3 ( \10472 , \8482 , \10471 );
nor \g444877/U$1 ( \10473 , \10452 , \10472 );
and \g446864/U$2 ( \10474 , \8509 , RIded30a0_865);
and \g446864/U$3 ( \10475 , RIded5698_892, \8511 );
nor \g446864/U$1 ( \10476 , \10474 , \10475 );
and \g446863/U$2 ( \10477 , \8514 , RIded7588_914);
and \g446863/U$3 ( \10478 , RIded9a18_940, \8517 );
nor \g446863/U$1 ( \10479 , \10477 , \10478 );
and \g446865/U$2 ( \10480 , \8969 , RIfca6b68_6919);
and \g446865/U$3 ( \10481 , RIfca65c8_6915, \8971 );
nor \g446865/U$1 ( \10482 , \10480 , \10481 );
nand \g444609/U$1 ( \10483 , \10473 , \10476 , \10479 , \10482 );
and \g452186/U$2 ( \10484 , \8326 , RIdf1fae0_1737);
and \g452186/U$3 ( \10485 , RIfc61fb8_6137, \8404 );
nor \g452186/U$1 ( \10486 , \10484 , \10485 );
and \g446087/U$2 ( \10487 , RIfc62558_6141, \8373 );
and \g446087/U$3 ( \10488 , RIdf1b1c0_1685, \8319 );
and \g448988/U$2 ( \10489 , RIfe81cd8_7821, \8412 );
and \g448988/U$3 ( \10490 , \8407 , RIdf281e0_1833);
and \g448988/U$4 ( \10491 , RIfca6fa0_6922, \8383 );
nor \g448988/U$1 ( \10492 , \10489 , \10490 , \10491 );
and \g452196/U$2 ( \10493 , \8356 , RIfcaac18_6965);
and \g452196/U$3 ( \10494 , RIfc44300_5798, \8359 );
nor \g452196/U$1 ( \10495 , \10493 , \10494 );
and \g454748/U$2 ( \10496 , \8313 , RIdf22ee8_1774);
and \g454748/U$3 ( \10497 , RIfcafc40_7022, \8323 );
nor \g454748/U$1 ( \10498 , \10496 , \10497 );
not \g450000/U$3 ( \10499 , \10498 );
not \g450000/U$4 ( \10500 , \8347 );
and \g450000/U$2 ( \10501 , \10499 , \10500 );
and \g450000/U$5 ( \10502 , \8351 , RIfccef78_7377);
nor \g450000/U$1 ( \10503 , \10501 , \10502 );
and \g452192/U$2 ( \10504 , \8378 , RIdf249a0_1793);
and \g452192/U$3 ( \10505 , RIfe81b70_7820, \8417 );
nor \g452192/U$1 ( \10506 , \10504 , \10505 );
nand \g447721/U$1 ( \10507 , \10492 , \10495 , \10503 , \10506 );
nor \g446087/U$1 ( \10508 , \10487 , \10488 , \10507 );
and \g452189/U$2 ( \10509 , \8335 , RIdf19438_1664);
and \g452189/U$3 ( \10510 , RIdf219d0_1759, \8340 );
nor \g452189/U$1 ( \10511 , \10509 , \10510 );
nand \g445595/U$1 ( \10512 , \10486 , \10508 , \10511 );
and \g444826/U$2 ( \10513 , \10512 , \8752 );
and \g448983/U$2 ( \10514 , RIdf11878_1576, \8373 );
and \g448983/U$3 ( \10515 , \8383 , RIdf14578_1608);
and \g448983/U$4 ( \10516 , RIdefb078_1320, \8488 );
nor \g448983/U$1 ( \10517 , \10514 , \10515 , \10516 );
and \g452175/U$2 ( \10518 , \8335 , RIdeea278_1128);
and \g452175/U$3 ( \10519 , RIdef2978_1224, \8340 );
nor \g452175/U$1 ( \10520 , \10518 , \10519 );
and \g452173/U$2 ( \10521 , \8404 , RIdf0eb78_1544);
and \g452173/U$3 ( \10522 , RIdf17278_1640, \8351 );
nor \g452173/U$1 ( \10523 , \10521 , \10522 );
and \g454746/U$2 ( \10524 , \8313 , RIdeecf78_1160);
and \g454746/U$3 ( \10525 , RIdeefc78_1192, \8323 );
nor \g454746/U$1 ( \10526 , \10524 , \10525 );
not \g454745/U$1 ( \10527 , \10526 );
and \g449995/U$2 ( \10528 , \10527 , \8316 );
and \g449995/U$3 ( \10529 , RIdefdd78_1352, \8359 );
nor \g449995/U$1 ( \10530 , \10528 , \10529 );
nand \g448187/U$1 ( \10531 , \10517 , \10520 , \10523 , \10530 );
and \g444826/U$3 ( \10532 , \8478 , \10531 );
nor \g444826/U$1 ( \10533 , \10513 , \10532 );
nor \g448365/U$1 ( \10534 , \8477 , \8408 );
and \g446854/U$2 ( \10535 , \10534 , RIdf09178_1480);
nor \g448364/U$1 ( \10536 , \8477 , \8433 );
and \g446854/U$3 ( \10537 , RIdf0be78_1512, \10536 );
nor \g446854/U$1 ( \10538 , \10535 , \10537 );
nor \g448308/U$1 ( \10539 , \8477 , \8437 );
and \g446855/U$2 ( \10540 , \10539 , RIdf03778_1416);
nor \g448367/U$1 ( \10541 , \8477 , \8413 );
and \g446855/U$3 ( \10542 , RIdf06478_1448, \10541 );
nor \g446855/U$1 ( \10543 , \10540 , \10542 );
and \g446859/U$2 ( \10544 , \8775 , RIdef5678_1256);
and \g446859/U$3 ( \10545 , RIdef8378_1288, \8777 );
nor \g446859/U$1 ( \10546 , \10544 , \10545 );
nand \g444608/U$1 ( \10547 , \10533 , \10538 , \10543 , \10546 );
and \g446065/U$2 ( \10548 , RIfc54020_5978, \8373 );
and \g446065/U$3 ( \10549 , RIdea41b0_390, \8317 );
and \g448966/U$2 ( \10550 , RIfc6b630_6244, \8531 );
and \g448966/U$3 ( \10551 , \8488 , RIdeb1ba8_486);
and \g448966/U$4 ( \10552 , RIdec29a8_678, \8383 );
nor \g448966/U$1 ( \10553 , \10550 , \10551 , \10552 );
and \g453534/U$2 ( \10554 , \8356 , RIdeaeea8_454);
and \g453534/U$3 ( \10555 , RIfc4fe08_5931, \8359 );
nor \g453534/U$1 ( \10556 , \10554 , \10555 );
and \g455223/U$2 ( \10557 , \8313 , RIdeba2a8_582);
and \g455223/U$3 ( \10558 , RIdebcfa8_614, \8323 );
nor \g455223/U$1 ( \10559 , \10557 , \10558 );
not \g449978/U$3 ( \10560 , \10559 );
not \g449978/U$4 ( \10561 , \8376 );
and \g449978/U$2 ( \10562 , \10560 , \10561 );
and \g449978/U$5 ( \10563 , \8351 , RIdec56a8_710);
nor \g449978/U$1 ( \10564 , \10562 , \10563 );
and \g452114/U$2 ( \10565 , \8378 , RIdeb75a8_550);
and \g452114/U$3 ( \10566 , RIee1f540_4815, \8417 );
nor \g452114/U$1 ( \10567 , \10565 , \10566 );
nand \g447708/U$1 ( \10568 , \10553 , \10556 , \10564 , \10567 );
nor \g446065/U$1 ( \10569 , \10548 , \10549 , \10568 );
and \g452108/U$2 ( \10570 , \8335 , RIde9d8b0_358);
and \g452108/U$3 ( \10571 , RIfc6a118_6229, \8340 );
nor \g452108/U$1 ( \10572 , \10570 , \10571 );
and \g452102/U$2 ( \10573 , \8324 , RIdeaaab0_422);
and \g452102/U$3 ( \10574 , RIdebfca8_646, \8404 );
nor \g452102/U$1 ( \10575 , \10573 , \10574 );
and \g445199/U$2 ( \10576 , \10569 , \10572 , \10575 );
nor \g445199/U$1 ( \10577 , \10576 , \8589 );
and \g446074/U$2 ( \10578 , RIfc653c0_6174, \8373 );
and \g446074/U$3 ( \10579 , RIe169cf8_2581, \8317 );
and \g448975/U$2 ( \10580 , RIfcca4f0_7324, \8531 );
and \g448975/U$3 ( \10581 , \8488 , RIfca76a8_6927);
and \g448975/U$4 ( \10582 , RIee1be68_4776, \8383 );
nor \g448975/U$1 ( \10583 , \10580 , \10581 , \10582 );
and \g453435/U$2 ( \10584 , \8356 , RIfc4ce38_5897);
and \g453435/U$3 ( \10585 , RIde81db8_223, \8359 );
nor \g453435/U$1 ( \10586 , \10584 , \10585 );
and \g454634/U$2 ( \10587 , \8313 , RIde89db0_262);
and \g454634/U$3 ( \10588 , RIde8df50_282, \8323 );
nor \g454634/U$1 ( \10589 , \10587 , \10588 );
not \g449985/U$3 ( \10590 , \10589 );
not \g449985/U$4 ( \10591 , \8376 );
and \g449985/U$2 ( \10592 , \10590 , \10591 );
and \g449985/U$5 ( \10593 , \8351 , RIfc69ce0_6226);
nor \g449985/U$1 ( \10594 , \10592 , \10593 );
and \g453560/U$2 ( \10595 , \8378 , RIde85c10_242);
and \g453560/U$3 ( \10596 , RIde91718_299, \8417 );
nor \g453560/U$1 ( \10597 , \10595 , \10596 );
nand \g447714/U$1 ( \10598 , \10583 , \10586 , \10594 , \10597 );
nor \g446074/U$1 ( \10599 , \10578 , \10579 , \10598 );
and \g452133/U$2 ( \10600 , \8335 , RIe167f70_2560);
and \g452133/U$3 ( \10601 , RIfc6b360_6242, \8340 );
nor \g452133/U$1 ( \10602 , \10600 , \10601 );
and \g451213/U$2 ( \10603 , \8324 , RIe16b918_2601);
and \g451213/U$3 ( \10604 , RIee1ac20_4763, \8404 );
nor \g451213/U$1 ( \10605 , \10603 , \10604 );
and \g445207/U$2 ( \10606 , \10599 , \10602 , \10605 );
nor \g445207/U$1 ( \10607 , \10606 , \8558 );
or \g444393/U$1 ( \10608 , \10483 , \10547 , \10577 , \10607 );
and \g446050/U$2 ( \10609 , RIee37690_5089, \8373 );
and \g446050/U$3 ( \10610 , RIe1494a8_2211, \8319 );
and \g448949/U$2 ( \10611 , RIe1575a8_2371, \8414 );
and \g448949/U$3 ( \10612 , \8409 , RIe15cfa8_2435);
and \g448949/U$4 ( \10613 , RIe1629a8_2499, \8383 );
nor \g448949/U$1 ( \10614 , \10611 , \10612 , \10613 );
and \g451711/U$2 ( \10615 , \8356 , RIe14eea8_2275);
and \g451711/U$3 ( \10616 , RIee35908_5068, \8359 );
nor \g451711/U$1 ( \10617 , \10615 , \10616 );
and \g454712/U$2 ( \10618 , \8313 , RIee34f30_5061);
and \g454712/U$3 ( \10619 , RIe151ba8_2307, \8323 );
nor \g454712/U$1 ( \10620 , \10618 , \10619 );
not \g449963/U$3 ( \10621 , \10620 );
not \g449963/U$4 ( \10622 , \8347 );
and \g449963/U$2 ( \10623 , \10621 , \10622 );
and \g449963/U$5 ( \10624 , \8351 , RIe1656a8_2531);
nor \g449963/U$1 ( \10625 , \10623 , \10624 );
and \g452053/U$2 ( \10626 , \8378 , RIe1548a8_2339);
and \g452053/U$3 ( \10627 , RIfce93f0_7676, \8417 );
nor \g452053/U$1 ( \10628 , \10626 , \10627 );
nand \g447699/U$1 ( \10629 , \10614 , \10617 , \10625 , \10628 );
nor \g446050/U$1 ( \10630 , \10609 , \10610 , \10629 );
and \g452050/U$2 ( \10631 , \8335 , RIe1467a8_2179);
and \g452050/U$3 ( \10632 , RIfce32e8_7607, \8340 );
nor \g452050/U$1 ( \10633 , \10631 , \10632 );
and \g452045/U$2 ( \10634 , \8326 , RIe14c1a8_2243);
and \g452045/U$3 ( \10635 , RIe15fca8_2467, \8404 );
nor \g452045/U$1 ( \10636 , \10634 , \10635 );
and \g445186/U$2 ( \10637 , \10630 , \10633 , \10636 );
nor \g445186/U$1 ( \10638 , \10637 , \8368 );
and \g446058/U$2 ( \10639 , RIfca9160_6946, \8373 );
and \g446058/U$3 ( \10640 , RIdf2f3c8_1914, \8335 );
and \g448956/U$2 ( \10641 , RIdf3cdc0_2069, \8412 );
and \g448956/U$3 ( \10642 , \8409 , RIdf3ef80_2093);
and \g448956/U$4 ( \10643 , RIfc687c8_6211, \8383 );
nor \g448956/U$1 ( \10644 , \10641 , \10642 , \10643 );
and \g452496/U$2 ( \10645 , \8356 , RIfc676e8_6199);
and \g452496/U$3 ( \10646 , RIfc64448_6163, \8359 );
nor \g452496/U$1 ( \10647 , \10645 , \10646 );
and \g454715/U$2 ( \10648 , \8313 , RIfca7978_6929);
and \g454715/U$3 ( \10649 , RIee2fad0_5001, \8323 );
nor \g454715/U$1 ( \10650 , \10648 , \10649 );
not \g449971/U$3 ( \10651 , \10650 );
not \g449971/U$4 ( \10652 , \8347 );
and \g449971/U$2 ( \10653 , \10651 , \10652 );
and \g449971/U$5 ( \10654 , \8351 , RIfcde2c0_7550);
nor \g449971/U$1 ( \10655 , \10653 , \10654 );
and \g452083/U$2 ( \10656 , \8378 , RIfebeb60_8290);
and \g452083/U$3 ( \10657 , RIe141078_2117, \8417 );
nor \g452083/U$1 ( \10658 , \10656 , \10657 );
nand \g447703/U$1 ( \10659 , \10644 , \10647 , \10655 , \10658 );
nor \g446058/U$1 ( \10660 , \10639 , \10640 , \10659 );
and \g452073/U$2 ( \10661 , \8340 , RIdf35a70_1987);
and \g452073/U$3 ( \10662 , RIfcb1590_7040, \8404 );
nor \g452073/U$1 ( \10663 , \10661 , \10662 );
and \g452078/U$2 ( \10664 , \8317 , RIdf31420_1937);
and \g452078/U$3 ( \10665 , RIdf335e0_1961, \8326 );
nor \g452078/U$1 ( \10666 , \10664 , \10665 );
and \g445190/U$2 ( \10667 , \10660 , \10663 , \10666 );
nor \g445190/U$1 ( \10668 , \10667 , \8422 );
or \g444242/U$1 ( \10669 , \10608 , \10638 , \10668 );
_DC \g265d/U$1 ( \10670 , \10669 , \8654 );
and \g452454/U$2 ( \10671 , \8326 , RIdf1f978_1736);
and \g452454/U$3 ( \10672 , RIfcd3fa0_7434, \8404 );
nor \g452454/U$1 ( \10673 , \10671 , \10672 );
and \g446143/U$2 ( \10674 , RIfc51050_5944, \8373 );
and \g446143/U$3 ( \10675 , RIdf1b058_1684, \8319 );
and \g449062/U$2 ( \10676 , RIdf22d80_1773, \8531 );
and \g449062/U$3 ( \10677 , \8488 , RIfce7ed8_7661);
and \g449062/U$4 ( \10678 , RIee2a3a0_4939, \8383 );
nor \g449062/U$1 ( \10679 , \10676 , \10677 , \10678 );
and \g452460/U$2 ( \10680 , \8356 , RIfc515f0_5948);
and \g452460/U$3 ( \10681 , RIfc84428_6527, \8359 );
nor \g452460/U$1 ( \10682 , \10680 , \10681 );
and \g454245/U$2 ( \10683 , \8313 , RIfe81198_7813);
and \g454245/U$3 ( \10684 , RIdf28078_1832, \8323 );
nor \g454245/U$1 ( \10685 , \10683 , \10684 );
not \g450076/U$3 ( \10686 , \10685 );
not \g450076/U$4 ( \10687 , \8376 );
and \g450076/U$2 ( \10688 , \10686 , \10687 );
and \g450076/U$5 ( \10689 , \8351 , RIfcb7968_7111);
nor \g450076/U$1 ( \10690 , \10688 , \10689 );
and \g452457/U$2 ( \10691 , \8378 , RIdf24838_1792);
and \g452457/U$3 ( \10692 , RIdf2a3a0_1857, \8417 );
nor \g452457/U$1 ( \10693 , \10691 , \10692 );
nand \g447757/U$1 ( \10694 , \10679 , \10682 , \10690 , \10693 );
nor \g446143/U$1 ( \10695 , \10674 , \10675 , \10694 );
and \g452455/U$2 ( \10696 , \8335 , RIdf192d0_1663);
and \g452455/U$3 ( \10697 , RIdf21868_1758, \8340 );
nor \g452455/U$1 ( \10698 , \10696 , \10697 );
nand \g445609/U$1 ( \10699 , \10673 , \10695 , \10698 );
and \g444724/U$2 ( \10700 , \10699 , \8752 );
and \g449058/U$2 ( \10701 , RIdef8210_1287, \8523 );
and \g449058/U$3 ( \10702 , \8486 , RIdefaf10_1319);
and \g449058/U$4 ( \10703 , RIdf14410_1607, \8383 );
nor \g449058/U$1 ( \10704 , \10701 , \10702 , \10703 );
and \g452446/U$2 ( \10705 , \8356 , RIdef5510_1255);
and \g452446/U$3 ( \10706 , RIdefdc10_1351, \8359 );
nor \g452446/U$1 ( \10707 , \10705 , \10706 );
and \g454260/U$2 ( \10708 , \8313 , RIdf06310_1447);
and \g454260/U$3 ( \10709 , RIdf09010_1479, \8323 );
nor \g454260/U$1 ( \10710 , \10708 , \10709 );
not \g450072/U$3 ( \10711 , \10710 );
not \g450072/U$4 ( \10712 , \8376 );
and \g450072/U$2 ( \10713 , \10711 , \10712 );
and \g450072/U$5 ( \10714 , \8351 , RIdf17110_1639);
nor \g450072/U$1 ( \10715 , \10713 , \10714 );
and \g452445/U$2 ( \10716 , \8378 , RIdf03610_1415);
and \g452445/U$3 ( \10717 , RIdf0bd10_1511, \8417 );
nor \g452445/U$1 ( \10718 , \10716 , \10717 );
nand \g447755/U$1 ( \10719 , \10704 , \10707 , \10715 , \10718 );
and \g444724/U$3 ( \10720 , \8478 , \10719 );
nor \g444724/U$1 ( \10721 , \10700 , \10720 );
and \g446913/U$2 ( \10722 , \8780 , RIdeefb10_1191);
and \g446913/U$3 ( \10723 , RIdef2810_1223, \8782 );
nor \g446913/U$1 ( \10724 , \10722 , \10723 );
and \g446912/U$2 ( \10725 , \9480 , RIdf0ea10_1543);
and \g446912/U$3 ( \10726 , RIdf11710_1575, \9482 );
nor \g446912/U$1 ( \10727 , \10725 , \10726 );
and \g446914/U$2 ( \10728 , \8785 , RIdeea110_1127);
and \g446914/U$3 ( \10729 , RIdeece10_1159, \8787 );
nor \g446914/U$1 ( \10730 , \10728 , \10729 );
nand \g444618/U$1 ( \10731 , \10721 , \10724 , \10727 , \10730 );
and \g452479/U$2 ( \10732 , \8326 , RIdee7410_1095);
and \g452479/U$3 ( \10733 , RIdec8240_741, \8404 );
nor \g452479/U$1 ( \10734 , \10732 , \10733 );
and \g446148/U$2 ( \10735 , RIdecaf40_773, \8373 );
and \g446148/U$3 ( \10736 , RIdedc178_968, \8319 );
and \g449069/U$2 ( \10737 , RIdf2c998_1884, \8531 );
and \g449069/U$3 ( \10738 , \8488 , RIdf38338_2016);
and \g449069/U$4 ( \10739 , RIdecdc40_805, \8383 );
nor \g449069/U$1 ( \10740 , \10737 , \10738 , \10739 );
and \g452488/U$2 ( \10741 , \8356 , RIdf1d218_1708);
and \g452488/U$3 ( \10742 , RIe143940_2146, \8359 );
nor \g452488/U$1 ( \10743 , \10741 , \10742 );
and \g454223/U$2 ( \10744 , \8313 , RIe16e348_2631);
and \g454223/U$3 ( \10745 , RIde96c68_325, \8323 );
nor \g454223/U$1 ( \10746 , \10744 , \10745 );
not \g450083/U$3 ( \10747 , \10746 );
not \g450083/U$4 ( \10748 , \8376 );
and \g450083/U$2 ( \10749 , \10747 , \10748 );
and \g450083/U$5 ( \10750 , \8351 , RIded0940_837);
nor \g450083/U$1 ( \10751 , \10749 , \10750 );
and \g452485/U$2 ( \10752 , \8378 , RIe15a140_2402);
and \g452485/U$3 ( \10753 , RIdeb4740_517, \8417 );
nor \g452485/U$1 ( \10754 , \10752 , \10753 );
nand \g447763/U$1 ( \10755 , \10740 , \10743 , \10751 , \10754 );
nor \g446148/U$1 ( \10756 , \10735 , \10736 , \10755 );
and \g452480/U$2 ( \10757 , \8335 , RIde7cbb0_198);
and \g452480/U$3 ( \10758 , RIdf00910_1383, \8340 );
nor \g452480/U$1 ( \10759 , \10757 , \10758 );
nand \g445612/U$1 ( \10760 , \10734 , \10756 , \10759 );
and \g444879/U$2 ( \10761 , \10760 , \9010 );
and \g449066/U$2 ( \10762 , RIfe80ec8_7811, \8319 );
and \g449066/U$3 ( \10763 , \8324 , RIded7420_913);
and \g449066/U$4 ( \10764 , RIfce9f30_7684, \8488 );
nor \g449066/U$1 ( \10765 , \10762 , \10763 , \10764 );
and \g452470/U$2 ( \10766 , \8335 , RIded2f38_864);
and \g452470/U$3 ( \10767 , RIfe81030_7812, \8340 );
nor \g452470/U$1 ( \10768 , \10766 , \10767 );
and \g452468/U$2 ( \10769 , \8404 , RIfc7e488_6459);
and \g452468/U$3 ( \10770 , RIfc7e1b8_6457, \8351 );
nor \g452468/U$1 ( \10771 , \10769 , \10770 );
and \g454233/U$2 ( \10772 , \8313 , RIfc7dab0_6452);
and \g454233/U$3 ( \10773 , RIfca19d8_6861, \8323 );
nor \g454233/U$1 ( \10774 , \10772 , \10773 );
not \g450080/U$3 ( \10775 , \10774 );
not \g450080/U$4 ( \10776 , \8328 );
and \g450080/U$2 ( \10777 , \10775 , \10776 );
and \g450080/U$5 ( \10778 , \8359 , RIfcb3750_7064);
nor \g450080/U$1 ( \10779 , \10777 , \10778 );
nand \g447760/U$1 ( \10780 , \10765 , \10768 , \10771 , \10779 );
and \g444879/U$3 ( \10781 , \8482 , \10780 );
nor \g444879/U$1 ( \10782 , \10761 , \10781 );
and \g446919/U$2 ( \10783 , \8964 , RIfe80d60_7810);
and \g446919/U$3 ( \10784 , RIdee49e0_1065, \8966 );
nor \g446919/U$1 ( \10785 , \10783 , \10784 );
and \g446920/U$2 ( \10786 , \8521 , RIfc56a50_6008);
and \g446920/U$3 ( \10787 , RIfc7e5f0_6460, \8525 );
nor \g446920/U$1 ( \10788 , \10786 , \10787 );
and \g446921/U$2 ( \10789 , \8974 , RIfe80bf8_7809);
and \g446921/U$3 ( \10790 , RIfeabba0_8270, \8976 );
nor \g446921/U$1 ( \10791 , \10789 , \10790 );
nand \g444619/U$1 ( \10792 , \10782 , \10785 , \10788 , \10791 );
and \g446133/U$2 ( \10793 , RIde8dc08_281, \8409 );
and \g446133/U$3 ( \10794 , RIde858c8_241, \8378 );
and \g449051/U$2 ( \10795 , RIfc9dec8_6819, \8373 );
and \g449051/U$3 ( \10796 , \8330 , RIfc507e0_5938);
and \g449051/U$4 ( \10797 , RIfc84860_6530, \8488 );
nor \g449051/U$1 ( \10798 , \10795 , \10796 , \10797 );
and \g452415/U$2 ( \10799 , \8335 , RIe167e08_2559);
and \g452415/U$3 ( \10800 , RIfcb7da0_7114, \8340 );
nor \g452415/U$1 ( \10801 , \10799 , \10800 );
and \g452414/U$2 ( \10802 , \8404 , RIfc853a0_6538);
and \g452414/U$3 ( \10803 , RIfc50678_5937, \8351 );
nor \g452414/U$1 ( \10804 , \10802 , \10803 );
and \g454276/U$2 ( \10805 , \8313 , RIe169b90_2580);
and \g454276/U$3 ( \10806 , RIe16b7b0_2600, \8323 );
nor \g454276/U$1 ( \10807 , \10805 , \10806 );
not \g454275/U$1 ( \10808 , \10807 );
and \g450065/U$2 ( \10809 , \10808 , \8316 );
and \g450065/U$3 ( \10810 , RIde81a70_222, \8359 );
nor \g450065/U$1 ( \10811 , \10809 , \10810 );
nand \g448199/U$1 ( \10812 , \10798 , \10801 , \10804 , \10811 );
nor \g446133/U$1 ( \10813 , \10793 , \10794 , \10812 );
and \g452411/U$2 ( \10814 , \8356 , RIfc84c98_6533);
and \g452411/U$3 ( \10815 , RIde913d0_298, \8417 );
nor \g452411/U$1 ( \10816 , \10814 , \10815 );
and \g452410/U$2 ( \10817 , \8531 , RIfc50948_5939);
and \g452410/U$3 ( \10818 , RIde89a68_261, \8414 );
nor \g452410/U$1 ( \10819 , \10817 , \10818 );
and \g445244/U$2 ( \10820 , \10813 , \10816 , \10819 );
nor \g445244/U$1 ( \10821 , \10820 , \8558 );
and \g446136/U$2 ( \10822 , RIfcc4dc0_7262, \8373 );
and \g446136/U$3 ( \10823 , RIdea3e68_389, \8319 );
and \g449054/U$2 ( \10824 , RIdeba140_581, \8414 );
and \g449054/U$3 ( \10825 , \8407 , RIdebce40_613);
and \g449054/U$4 ( \10826 , RIdec2840_677, \8330 );
nor \g449054/U$1 ( \10827 , \10824 , \10825 , \10826 );
and \g452431/U$2 ( \10828 , \8356 , RIdeaed40_453);
and \g452431/U$3 ( \10829 , RIfc4d978_5905, \8359 );
nor \g452431/U$1 ( \10830 , \10828 , \10829 );
and \g454854/U$2 ( \10831 , \8313 , RIfc9dbf8_6817);
and \g454854/U$3 ( \10832 , RIdeb1a40_485, \8323 );
nor \g454854/U$1 ( \10833 , \10831 , \10832 );
not \g450068/U$3 ( \10834 , \10833 );
not \g450068/U$4 ( \10835 , \8347 );
and \g450068/U$2 ( \10836 , \10834 , \10835 );
and \g450068/U$5 ( \10837 , \8351 , RIdec5540_709);
nor \g450068/U$1 ( \10838 , \10836 , \10837 );
and \g452428/U$2 ( \10839 , \8378 , RIdeb7440_549);
and \g452428/U$3 ( \10840 , RIfc9d7c0_6814, \8417 );
nor \g452428/U$1 ( \10841 , \10839 , \10840 );
nand \g447752/U$1 ( \10842 , \10827 , \10830 , \10838 , \10841 );
nor \g446136/U$1 ( \10843 , \10822 , \10823 , \10842 );
and \g452423/U$2 ( \10844 , \8335 , RIde9d568_357);
and \g452423/U$3 ( \10845 , RIfcb8610_7120, \8340 );
nor \g452423/U$1 ( \10846 , \10844 , \10845 );
and \g452422/U$2 ( \10847 , \8326 , RIdeaa768_421);
and \g452422/U$3 ( \10848 , RIdebfb40_645, \8404 );
nor \g452422/U$1 ( \10849 , \10847 , \10848 );
and \g445246/U$2 ( \10850 , \10843 , \10846 , \10849 );
nor \g445246/U$1 ( \10851 , \10850 , \8589 );
or \g444398/U$1 ( \10852 , \10731 , \10792 , \10821 , \10851 );
and \g446126/U$2 ( \10853 , RIe15ce40_2434, \8409 );
and \g446126/U$3 ( \10854 , RIe154740_2338, \8378 );
and \g449042/U$2 ( \10855 , RIee37528_5088, \8373 );
and \g449042/U$3 ( \10856 , \8383 , RIe162840_2498);
and \g449042/U$4 ( \10857 , RIe151a40_2306, \8488 );
nor \g449042/U$1 ( \10858 , \10855 , \10856 , \10857 );
and \g452389/U$2 ( \10859 , \8335 , RIe146640_2178);
and \g452389/U$3 ( \10860 , RIfcc6170_7276, \8340 );
nor \g452389/U$1 ( \10861 , \10859 , \10860 );
and \g452387/U$2 ( \10862 , \8404 , RIe15fb40_2466);
and \g452387/U$3 ( \10863 , RIe165540_2530, \8351 );
nor \g452387/U$1 ( \10864 , \10862 , \10863 );
and \g454302/U$2 ( \10865 , \8313 , RIe149340_2210);
and \g454302/U$3 ( \10866 , RIe14c040_2242, \8323 );
nor \g454302/U$1 ( \10867 , \10865 , \10866 );
not \g454301/U$1 ( \10868 , \10867 );
and \g450057/U$2 ( \10869 , \10868 , \8316 );
and \g450057/U$3 ( \10870 , RIfcd35c8_7427, \8359 );
nor \g450057/U$1 ( \10871 , \10869 , \10870 );
nand \g448197/U$1 ( \10872 , \10858 , \10861 , \10864 , \10871 );
nor \g446126/U$1 ( \10873 , \10853 , \10854 , \10872 );
and \g452382/U$2 ( \10874 , \8356 , RIe14ed40_2274);
and \g452382/U$3 ( \10875 , RIfcb5be0_7090, \8417 );
nor \g452382/U$1 ( \10876 , \10874 , \10875 );
and \g452381/U$2 ( \10877 , \8531 , RIfc53a80_5974);
and \g452381/U$3 ( \10878 , RIe157440_2370, \8414 );
nor \g452381/U$1 ( \10879 , \10877 , \10878 );
and \g445238/U$2 ( \10880 , \10873 , \10876 , \10879 );
nor \g445238/U$1 ( \10881 , \10880 , \8368 );
and \g446130/U$2 ( \10882 , RIdf3ee18_2092, \8409 );
and \g446130/U$3 ( \10883 , RIdf3a7c8_2042, \8378 );
and \g449047/U$2 ( \10884 , RIfcb4f38_7081, \8373 );
and \g449047/U$3 ( \10885 , \8330 , RIee33310_5041);
and \g449047/U$4 ( \10886 , RIfcd27b8_7417, \8488 );
nor \g449047/U$1 ( \10887 , \10884 , \10885 , \10886 );
and \g452402/U$2 ( \10888 , \8335 , RIdf2f260_1913);
and \g452402/U$3 ( \10889 , RIdf35908_1986, \8340 );
nor \g452402/U$1 ( \10890 , \10888 , \10889 );
and \g452398/U$2 ( \10891 , \8404 , RIfc47f78_5841);
and \g452398/U$3 ( \10892 , RIfc7f130_6468, \8351 );
nor \g452398/U$1 ( \10893 , \10891 , \10892 );
and \g454292/U$2 ( \10894 , \8313 , RIfebe9f8_8289);
and \g454292/U$3 ( \10895 , RIdf33478_1960, \8323 );
nor \g454292/U$1 ( \10896 , \10894 , \10895 );
not \g454291/U$1 ( \10897 , \10896 );
and \g450061/U$2 ( \10898 , \10897 , \8316 );
and \g450061/U$3 ( \10899 , RIfc7fc70_6476, \8359 );
nor \g450061/U$1 ( \10900 , \10898 , \10899 );
nand \g448198/U$1 ( \10901 , \10887 , \10890 , \10893 , \10900 );
nor \g446130/U$1 ( \10902 , \10882 , \10883 , \10901 );
and \g452397/U$2 ( \10903 , \8356 , RIfcc6b48_7283);
and \g452397/U$3 ( \10904 , RIe140f10_2116, \8417 );
nor \g452397/U$1 ( \10905 , \10903 , \10904 );
and \g452396/U$2 ( \10906 , \8531 , RIfca1000_6854);
and \g452396/U$3 ( \10907 , RIdf3cc58_2068, \8414 );
nor \g452396/U$1 ( \10908 , \10906 , \10907 );
and \g445242/U$2 ( \10909 , \10902 , \10905 , \10908 );
nor \g445242/U$1 ( \10910 , \10909 , \8422 );
or \g444244/U$1 ( \10911 , \10852 , \10881 , \10910 );
_DC \g26e2/U$1 ( \10912 , \10911 , \8654 );
and \g447177/U$2 ( \10913 , \10044 , RIfe7dc28_7775);
and \g447177/U$3 ( \10914 , RIee38770_5101, \10046 );
nor \g447177/U$1 ( \10915 , \10913 , \10914 );
and \g446438/U$2 ( \10916 , RIee1cde0_4787, \8351 );
and \g446438/U$3 ( \10917 , RIee1bd00_4775, \8383 );
and \g449447/U$2 ( \10918 , RIfe7dac0_7774, \8414 );
and \g449447/U$3 ( \10919 , \8409 , RIde8d8c0_280);
and \g449447/U$4 ( \10920 , RIfe7dd90_7776, \8326 );
nor \g449447/U$1 ( \10921 , \10918 , \10919 , \10920 );
and \g453875/U$2 ( \10922 , \8356 , RIfc768c8_6371);
and \g453875/U$3 ( \10923 , RIee1a518_4758, \8359 );
nor \g453875/U$1 ( \10924 , \10922 , \10923 );
and \g455053/U$2 ( \10925 , \8313 , RIee19b40_4751);
and \g455053/U$3 ( \10926 , RIee19e10_4753, \8323 );
nor \g455053/U$1 ( \10927 , \10925 , \10926 );
not \g450466/U$3 ( \10928 , \10927 );
not \g450466/U$4 ( \10929 , \8347 );
and \g450466/U$2 ( \10930 , \10928 , \10929 );
and \g450466/U$5 ( \10931 , \8340 , RIfcd05f8_7393);
nor \g450466/U$1 ( \10932 , \10930 , \10931 );
and \g453870/U$2 ( \10933 , \8378 , RIfe7d958_7773);
and \g453870/U$3 ( \10934 , RIde91088_297, \8417 );
nor \g453870/U$1 ( \10935 , \10933 , \10934 );
nand \g447972/U$1 ( \10936 , \10921 , \10924 , \10932 , \10935 );
nor \g446438/U$1 ( \10937 , \10916 , \10917 , \10936 );
not \g444822/U$3 ( \10938 , \10937 );
not \g444822/U$4 ( \10939 , \8558 );
and \g444822/U$2 ( \10940 , \10938 , \10939 );
and \g446448/U$2 ( \10941 , RIdeb9fd8_580, \8414 );
and \g446448/U$3 ( \10942 , RIdeaebd8_452, \8356 );
and \g449457/U$2 ( \10943 , RIdea3b20_388, \8319 );
and \g449457/U$3 ( \10944 , \8324 , RIdeaa420_420);
and \g449457/U$4 ( \10945 , RIdebccd8_612, \8409 );
nor \g449457/U$1 ( \10946 , \10943 , \10944 , \10945 );
and \g453916/U$2 ( \10947 , \8335 , RIde9d220_356);
and \g453916/U$3 ( \10948 , RIee1da88_4796, \8340 );
nor \g453916/U$1 ( \10949 , \10947 , \10948 );
and \g453911/U$2 ( \10950 , \8404 , RIdebf9d8_644);
and \g453911/U$3 ( \10951 , RIdec53d8_708, \8351 );
nor \g453911/U$1 ( \10952 , \10950 , \10951 );
and \g455046/U$2 ( \10953 , \8313 , RIee20080_4823);
and \g455046/U$3 ( \10954 , RIdec26d8_676, \8323 );
nor \g455046/U$1 ( \10955 , \10953 , \10954 );
not \g450476/U$3 ( \10956 , \10955 );
not \g450476/U$4 ( \10957 , \8328 );
and \g450476/U$2 ( \10958 , \10956 , \10957 );
and \g450476/U$5 ( \10959 , \8417 , RIee1f3d8_4814);
nor \g450476/U$1 ( \10960 , \10958 , \10959 );
nand \g447978/U$1 ( \10961 , \10946 , \10949 , \10952 , \10960 );
nor \g446448/U$1 ( \10962 , \10941 , \10942 , \10961 );
and \g453901/U$2 ( \10963 , \8378 , RIdeb72d8_548);
and \g453901/U$3 ( \10964 , RIee1ee38_4810, \8359 );
nor \g453901/U$1 ( \10965 , \10963 , \10964 );
and \g453898/U$2 ( \10966 , \8531 , RIee1e898_4806);
and \g453898/U$3 ( \10967 , RIdeb18d8_484, \8488 );
nor \g453898/U$1 ( \10968 , \10966 , \10967 );
and \g445460/U$2 ( \10969 , \10962 , \10965 , \10968 );
nor \g445460/U$1 ( \10970 , \10969 , \8589 );
nor \g444822/U$1 ( \10971 , \10940 , \10970 );
and \g447184/U$2 ( \10972 , \10039 , RIfcd8a28_7487);
and \g447184/U$3 ( \10973 , RIee1b490_4769, \10041 );
nor \g447184/U$1 ( \10974 , \10972 , \10973 );
nand \g444439/U$1 ( \10975 , \10915 , \10971 , \10974 );
and \g453968/U$2 ( \10976 , \8378 , RIdf034a8_1414);
and \g453968/U$3 ( \10977 , RIdefada8_1318, \8488 );
nor \g453968/U$1 ( \10978 , \10976 , \10977 );
and \g446462/U$2 ( \10979 , RIdf061a8_1446, \8414 );
and \g446462/U$3 ( \10980 , RIdef80a8_1286, \8523 );
and \g449476/U$2 ( \10981 , RIdf08ea8_1478, \8409 );
and \g449476/U$3 ( \10982 , \8373 , RIdf115a8_1574);
and \g449476/U$4 ( \10983 , RIdf142a8_1606, \8383 );
nor \g449476/U$1 ( \10984 , \10981 , \10982 , \10983 );
and \g453985/U$2 ( \10985 , \8335 , RIdee9fa8_1126);
and \g453985/U$3 ( \10986 , RIdef26a8_1222, \8340 );
nor \g453985/U$1 ( \10987 , \10985 , \10986 );
and \g453979/U$2 ( \10988 , \8404 , RIdf0e8a8_1542);
and \g453979/U$3 ( \10989 , RIdf16fa8_1638, \8351 );
nor \g453979/U$1 ( \10990 , \10988 , \10989 );
and \g455005/U$2 ( \10991 , \8313 , RIdeecca8_1158);
and \g455005/U$3 ( \10992 , RIdeef9a8_1190, \8323 );
nor \g455005/U$1 ( \10993 , \10991 , \10992 );
not \g455004/U$1 ( \10994 , \10993 );
and \g450497/U$2 ( \10995 , \10994 , \8316 );
and \g450497/U$3 ( \10996 , RIdf0bba8_1510, \8417 );
nor \g450497/U$1 ( \10997 , \10995 , \10996 );
nand \g448246/U$1 ( \10998 , \10984 , \10987 , \10990 , \10997 );
nor \g446462/U$1 ( \10999 , \10979 , \10980 , \10998 );
and \g453967/U$2 ( \11000 , \8356 , RIdef53a8_1254);
and \g453967/U$3 ( \11001 , RIdefdaa8_1350, \8359 );
nor \g453967/U$1 ( \11002 , \11000 , \11001 );
nand \g445694/U$1 ( \11003 , \10978 , \10999 , \11002 );
and \g444808/U$2 ( \11004 , \11003 , \8478 );
and \g449466/U$2 ( \11005 , RIfebe188_8283, \8409 );
and \g449466/U$3 ( \11006 , \8373 , RIfebe020_8282);
and \g449466/U$4 ( \11007 , RIee249a0_4875, \8330 );
nor \g449466/U$1 ( \11008 , \11005 , \11006 , \11007 );
and \g453945/U$2 ( \11009 , \8335 , RIded2dd0_863);
and \g453945/U$3 ( \11010 , RIded98b0_939, \8340 );
nor \g453945/U$1 ( \11011 , \11009 , \11010 );
and \g453944/U$2 ( \11012 , \8404 , RIee23488_4860);
and \g453944/U$3 ( \11013 , RIee25648_4884, \8351 );
nor \g453944/U$1 ( \11014 , \11012 , \11013 );
and \g454361/U$2 ( \11015 , \8313 , RIded5530_891);
and \g454361/U$3 ( \11016 , RIded72b8_912, \8323 );
nor \g454361/U$1 ( \11017 , \11015 , \11016 );
not \g454360/U$1 ( \11018 , \11017 );
and \g450485/U$2 ( \11019 , \11018 , \8316 );
and \g450485/U$3 ( \11020 , RIfebe2f0_8284, \8417 );
nor \g450485/U$1 ( \11021 , \11019 , \11020 );
nand \g448245/U$1 ( \11022 , \11008 , \11011 , \11014 , \11021 );
and \g444808/U$3 ( \11023 , \8482 , \11022 );
nor \g444808/U$1 ( \11024 , \11004 , \11023 );
and \g447198/U$2 ( \11025 , \8521 , RIfc618b0_6132);
and \g447198/U$3 ( \11026 , RIfc787b8_6393, \8525 );
nor \g447198/U$1 ( \11027 , \11025 , \11026 );
and \g447197/U$2 ( \11028 , \10290 , RIfc7aae0_6418);
and \g447197/U$3 ( \11029 , RIfcbf7f8_7201, \10293 );
nor \g447197/U$1 ( \11030 , \11028 , \11029 );
and \g447199/U$2 ( \11031 , \8974 , RIfe7e060_7778);
and \g447199/U$3 ( \11032 , RIfe7e1c8_7779, \8976 );
nor \g447199/U$1 ( \11033 , \11031 , \11032 );
nand \g444543/U$1 ( \11034 , \11024 , \11027 , \11030 , \11033 );
and \g446423/U$2 ( \11035 , RIee373c0_5087, \8373 );
and \g446423/U$3 ( \11036 , RIe1626d8_2497, \8330 );
and \g449425/U$2 ( \11037 , RIe1572d8_2369, \8414 );
and \g449425/U$3 ( \11038 , \8409 , RIe15ccd8_2433);
and \g449425/U$4 ( \11039 , RIe14bed8_2241, \8324 );
nor \g449425/U$1 ( \11040 , \11037 , \11038 , \11039 );
and \g453807/U$2 ( \11041 , \8356 , RIe14ebd8_2273);
and \g453807/U$3 ( \11042 , RIfe7def8_7777, \8359 );
nor \g453807/U$1 ( \11043 , \11041 , \11042 );
and \g455061/U$2 ( \11044 , \8313 , RIfebdeb8_8281);
and \g455061/U$3 ( \11045 , RIe1518d8_2305, \8323 );
nor \g455061/U$1 ( \11046 , \11044 , \11045 );
not \g450447/U$3 ( \11047 , \11046 );
not \g450447/U$4 ( \11048 , \8347 );
and \g450447/U$2 ( \11049 , \11047 , \11048 );
and \g450447/U$5 ( \11050 , \8340 , RIfc649e8_6167);
nor \g450447/U$1 ( \11051 , \11049 , \11050 );
and \g453802/U$2 ( \11052 , \8378 , RIe1545d8_2337);
and \g453802/U$3 ( \11053 , RIee362e0_5075, \8417 );
nor \g453802/U$1 ( \11054 , \11052 , \11053 );
nand \g447961/U$1 ( \11055 , \11040 , \11043 , \11051 , \11054 );
nor \g446423/U$1 ( \11056 , \11035 , \11036 , \11055 );
and \g453788/U$2 ( \11057 , \8335 , RIe1464d8_2177);
and \g453788/U$3 ( \11058 , RIe1653d8_2529, \8351 );
nor \g453788/U$1 ( \11059 , \11057 , \11058 );
and \g453794/U$2 ( \11060 , \8317 , RIe1491d8_2209);
and \g453794/U$3 ( \11061 , RIe15f9d8_2465, \8404 );
nor \g453794/U$1 ( \11062 , \11060 , \11061 );
and \g445444/U$2 ( \11063 , \11056 , \11059 , \11062 );
nor \g445444/U$1 ( \11064 , \11063 , \8368 );
and \g446430/U$2 ( \11065 , RIfebdbe8_8279, \8412 );
and \g446430/U$3 ( \11066 , RIee2d7a8_4976, \8356 );
and \g449435/U$2 ( \11067 , RIdf312b8_1936, \8319 );
and \g449435/U$3 ( \11068 , \8324 , RIdf33310_1959);
and \g449435/U$4 ( \11069 , RIfe7d520_7770, \8409 );
nor \g449435/U$1 ( \11070 , \11067 , \11068 , \11069 );
and \g453837/U$2 ( \11071 , \8335 , RIdf2f0f8_1912);
and \g453837/U$3 ( \11072 , RIdf357a0_1985, \8340 );
nor \g453837/U$1 ( \11073 , \11071 , \11072 );
and \g453833/U$2 ( \11074 , \8404 , RIfceb9e8_7703);
and \g453833/U$3 ( \11075 , RIfe7d7f0_7772, \8351 );
nor \g453833/U$1 ( \11076 , \11074 , \11075 );
and \g454534/U$2 ( \11077 , \8313 , RIee32230_5029);
and \g454534/U$3 ( \11078 , RIfe7d688_7771, \8323 );
nor \g454534/U$1 ( \11079 , \11077 , \11078 );
not \g450455/U$3 ( \11080 , \11079 );
not \g450455/U$4 ( \11081 , \8328 );
and \g450455/U$2 ( \11082 , \11080 , \11081 );
and \g450455/U$5 ( \11083 , \8417 , RIfebdd50_8280);
nor \g450455/U$1 ( \11084 , \11082 , \11083 );
nand \g447965/U$1 ( \11085 , \11070 , \11073 , \11076 , \11084 );
nor \g446430/U$1 ( \11086 , \11065 , \11066 , \11085 );
and \g453822/U$2 ( \11087 , \8378 , RIfe7d3b8_7769);
and \g453822/U$3 ( \11088 , RIfc734c0_6334, \8359 );
nor \g453822/U$1 ( \11089 , \11087 , \11088 );
and \g453820/U$2 ( \11090 , \8523 , RIfccfab8_7385);
and \g453820/U$3 ( \11091 , RIee2f968_5000, \8488 );
nor \g453820/U$1 ( \11092 , \11090 , \11091 );
and \g445450/U$2 ( \11093 , \11086 , \11089 , \11092 );
nor \g445450/U$1 ( \11094 , \11093 , \8422 );
or \g444304/U$1 ( \11095 , \10975 , \11034 , \11064 , \11094 );
and \g446409/U$2 ( \11096 , RIfe7ce18_7765, \8417 );
and \g446409/U$3 ( \11097 , RIfe7d0e8_7767, \8335 );
and \g449407/U$2 ( \11098 , RIfe7d250_7768, \8326 );
and \g449407/U$3 ( \11099 , \8373 , RIee28e88_4924);
and \g449407/U$4 ( \11100 , RIee2a238_4938, \8383 );
nor \g449407/U$1 ( \11101 , \11098 , \11099 , \11100 );
and \g455112/U$2 ( \11102 , \8313 , RIee26890_4897);
and \g455112/U$3 ( \11103 , RIee26e30_4901, \8323 );
nor \g455112/U$1 ( \11104 , \11102 , \11103 );
not \g450427/U$3 ( \11105 , \11104 );
not \g450427/U$4 ( \11106 , \8347 );
and \g450427/U$2 ( \11107 , \11105 , \11106 );
and \g450427/U$5 ( \11108 , \8340 , RIee262f0_4893);
nor \g450427/U$1 ( \11109 , \11107 , \11108 );
and \g453731/U$2 ( \11110 , \8404 , RIee27c40_4911);
and \g453731/U$3 ( \11111 , RIee2bcf0_4957, \8351 );
nor \g453731/U$1 ( \11112 , \11110 , \11111 );
and \g453740/U$2 ( \11113 , \8356 , RIfcaa0d8_6957);
and \g453740/U$3 ( \11114 , RIee27268_4904, \8359 );
nor \g453740/U$1 ( \11115 , \11113 , \11114 );
nand \g447950/U$1 ( \11116 , \11101 , \11109 , \11112 , \11115 );
nor \g446409/U$1 ( \11117 , \11096 , \11097 , \11116 );
and \g453721/U$2 ( \11118 , \8317 , RIee26020_4891);
and \g453721/U$3 ( \11119 , RIfe7cb48_7763, \8378 );
nor \g453721/U$1 ( \11120 , \11118 , \11119 );
and \g453716/U$2 ( \11121 , \8414 , RIfe7cf80_7766);
and \g453716/U$3 ( \11122 , RIfe7ccb0_7764, \8409 );
nor \g453716/U$1 ( \11123 , \11121 , \11122 );
and \g445435/U$2 ( \11124 , \11117 , \11120 , \11123 );
nor \g445435/U$1 ( \11125 , \11124 , \8621 );
and \g446415/U$2 ( \11126 , RIe16e1e0_2630, \8414 );
and \g446415/U$3 ( \11127 , RIdf1d0b0_1707, \8356 );
and \g449417/U$2 ( \11128 , RIdedc010_967, \8319 );
and \g449417/U$3 ( \11129 , \8324 , RIdee72a8_1094);
and \g449417/U$4 ( \11130 , RIde96920_324, \8407 );
nor \g449417/U$1 ( \11131 , \11128 , \11129 , \11130 );
and \g453767/U$2 ( \11132 , \8335 , RIde7c868_197);
and \g453767/U$3 ( \11133 , RIdf007a8_1382, \8340 );
nor \g453767/U$1 ( \11134 , \11132 , \11133 );
and \g453762/U$2 ( \11135 , \8404 , RIdec80d8_740);
and \g453762/U$3 ( \11136 , RIded07d8_836, \8351 );
nor \g453762/U$1 ( \11137 , \11135 , \11136 );
and \g454319/U$2 ( \11138 , \8313 , RIdecadd8_772);
and \g454319/U$3 ( \11139 , RIdecdad8_804, \8323 );
nor \g454319/U$1 ( \11140 , \11138 , \11139 );
not \g450437/U$3 ( \11141 , \11140 );
not \g450437/U$4 ( \11142 , \8328 );
and \g450437/U$2 ( \11143 , \11141 , \11142 );
and \g450437/U$5 ( \11144 , \8417 , RIdeb45d8_516);
nor \g450437/U$1 ( \11145 , \11143 , \11144 );
nand \g447956/U$1 ( \11146 , \11131 , \11134 , \11137 , \11145 );
nor \g446415/U$1 ( \11147 , \11126 , \11127 , \11146 );
and \g453755/U$2 ( \11148 , \8378 , RIe159fd8_2401);
and \g453755/U$3 ( \11149 , RIe1437d8_2145, \8359 );
nor \g453755/U$1 ( \11150 , \11148 , \11149 );
and \g453751/U$2 ( \11151 , \8523 , RIdf2c830_1883);
and \g453751/U$3 ( \11152 , RIdf381d0_2015, \8486 );
nor \g453751/U$1 ( \11153 , \11151 , \11152 );
and \g445440/U$2 ( \11154 , \11147 , \11150 , \11153 );
nor \g445440/U$1 ( \11155 , \11154 , \8651 );
or \g444174/U$1 ( \11156 , \11095 , \11125 , \11155 );
_DC \g2767/U$1 ( \11157 , \11156 , \8654 );
and \g450915/U$2 ( \11158 , \8531 , RIdf22c18_1772);
and \g450915/U$3 ( \11159 , RIfe7f6e0_7794, \8414 );
nor \g450915/U$1 ( \11160 , \11158 , \11159 );
and \g445780/U$2 ( \11161 , RIdf27f10_1831, \8409 );
and \g445780/U$3 ( \11162 , RIdf246d0_1791, \8378 );
and \g448602/U$2 ( \11163 , RIee28d20_4923, \8373 );
and \g448602/U$3 ( \11164 , \8330 , RIee2a0d0_4937);
and \g448602/U$4 ( \11165 , RIfc63638_6153, \8486 );
nor \g448602/U$1 ( \11166 , \11163 , \11164 , \11165 );
and \g450932/U$2 ( \11167 , \8335 , RIdf19168_1662);
and \g450932/U$3 ( \11168 , RIdf21700_1757, \8340 );
nor \g450932/U$1 ( \11169 , \11167 , \11168 );
and \g450925/U$2 ( \11170 , \8404 , RIfe7f578_7793);
and \g450925/U$3 ( \11171 , RIee2bb88_4956, \8351 );
nor \g450925/U$1 ( \11172 , \11170 , \11171 );
and \g454503/U$2 ( \11173 , \8313 , RIfeaa958_8257);
and \g454503/U$3 ( \11174 , RIdf1f810_1735, \8323 );
nor \g454503/U$1 ( \11175 , \11173 , \11174 );
not \g454502/U$1 ( \11176 , \11175 );
and \g449627/U$2 ( \11177 , \11176 , \8316 );
and \g449627/U$3 ( \11178 , RIfcce9d8_7373, \8359 );
nor \g449627/U$1 ( \11179 , \11177 , \11178 );
nand \g448145/U$1 ( \11180 , \11166 , \11169 , \11172 , \11179 );
nor \g445780/U$1 ( \11181 , \11161 , \11162 , \11180 );
and \g450920/U$2 ( \11182 , \8356 , RIfc62990_6144);
and \g450920/U$3 ( \11183 , RIdf2a238_1856, \8417 );
nor \g450920/U$1 ( \11184 , \11182 , \11183 );
nand \g445525/U$1 ( \11185 , \11160 , \11181 , \11184 );
and \g444839/U$2 ( \11186 , \11185 , \8752 );
and \g448591/U$2 ( \11187 , RIdecac70_771, \8371 );
and \g448591/U$3 ( \11188 , \8383 , RIdecd970_803);
and \g448591/U$4 ( \11189 , RIdf38068_2014, \8488 );
nor \g448591/U$1 ( \11190 , \11187 , \11188 , \11189 );
and \g450900/U$2 ( \11191 , \8335 , RIde7c520_196);
and \g450900/U$3 ( \11192 , RIdf00640_1381, \8340 );
nor \g450900/U$1 ( \11193 , \11191 , \11192 );
and \g450895/U$2 ( \11194 , \8404 , RIdec7f70_739);
and \g450895/U$3 ( \11195 , RIded0670_835, \8351 );
nor \g450895/U$1 ( \11196 , \11194 , \11195 );
and \g454607/U$2 ( \11197 , \8313 , RIdedbea8_966);
and \g454607/U$3 ( \11198 , RIdee7140_1093, \8323 );
nor \g454607/U$1 ( \11199 , \11197 , \11198 );
not \g454606/U$1 ( \11200 , \11199 );
and \g449617/U$2 ( \11201 , \11200 , \8316 );
and \g449617/U$3 ( \11202 , RIe143670_2144, \8359 );
nor \g449617/U$1 ( \11203 , \11201 , \11202 );
nand \g448144/U$1 ( \11204 , \11190 , \11193 , \11196 , \11203 );
and \g444839/U$3 ( \11205 , \9010 , \11204 );
nor \g444839/U$1 ( \11206 , \11186 , \11205 );
and \g446574/U$2 ( \11207 , \9031 , RIe159e70_2400);
and \g446574/U$3 ( \11208 , RIe16e078_2629, \9033 );
nor \g446574/U$1 ( \11209 , \11207 , \11208 );
and \g446575/U$2 ( \11210 , \9036 , RIde965d8_323);
and \g446575/U$3 ( \11211 , RIdeb4470_515, \9038 );
nor \g446575/U$1 ( \11212 , \11210 , \11211 );
nor \g448386/U$1 ( \11213 , \8651 , \8520 );
and \g446576/U$2 ( \11214 , \11213 , RIdf1cf48_1706);
nor \g448385/U$1 ( \11215 , \8651 , \8524 );
and \g446576/U$3 ( \11216 , RIdf2c6c8_1882, \11215 );
nor \g446576/U$1 ( \11217 , \11214 , \11216 );
nand \g444557/U$1 ( \11218 , \11206 , \11209 , \11212 , \11217 );
and \g450847/U$2 ( \11219 , \8324 , RIdeef840_1189);
and \g450847/U$3 ( \11220 , RIdf0e740_1541, \8404 );
nor \g450847/U$1 ( \11221 , \11219 , \11220 );
and \g445765/U$2 ( \11222 , RIdf11440_1573, \8371 );
and \g445765/U$3 ( \11223 , RIdeecb40_1157, \8319 );
and \g448582/U$2 ( \11224 , RIdf06040_1445, \8412 );
and \g448582/U$3 ( \11225 , \8409 , RIdf08d40_1477);
and \g448582/U$4 ( \11226 , RIdf14140_1605, \8383 );
nor \g448582/U$1 ( \11227 , \11224 , \11225 , \11226 );
and \g450864/U$2 ( \11228 , \8356 , RIdef5240_1253);
and \g450864/U$3 ( \11229 , RIdefd940_1349, \8359 );
nor \g450864/U$1 ( \11230 , \11228 , \11229 );
and \g454635/U$2 ( \11231 , \8313 , RIdef7f40_1285);
and \g454635/U$3 ( \11232 , RIdefac40_1317, \8323 );
nor \g454635/U$1 ( \11233 , \11231 , \11232 );
not \g449606/U$3 ( \11234 , \11233 );
not \g449606/U$4 ( \11235 , \8347 );
and \g449606/U$2 ( \11236 , \11234 , \11235 );
and \g449606/U$5 ( \11237 , \8351 , RIdf16e40_1637);
nor \g449606/U$1 ( \11238 , \11236 , \11237 );
and \g450858/U$2 ( \11239 , \8378 , RIdf03340_1413);
and \g450858/U$3 ( \11240 , RIdf0ba40_1509, \8417 );
nor \g450858/U$1 ( \11241 , \11239 , \11240 );
nand \g447492/U$1 ( \11242 , \11227 , \11230 , \11238 , \11241 );
nor \g445765/U$1 ( \11243 , \11222 , \11223 , \11242 );
and \g450852/U$2 ( \11244 , \8335 , RIdee9e40_1125);
and \g450852/U$3 ( \11245 , RIdef2540_1221, \8340 );
nor \g450852/U$1 ( \11246 , \11244 , \11245 );
nand \g445520/U$1 ( \11247 , \11221 , \11243 , \11246 );
and \g444754/U$2 ( \11248 , \11247 , \8478 );
and \g448572/U$2 ( \11249 , RIfc4cb68_5895, \8373 );
and \g448572/U$3 ( \11250 , \8383 , RIee24838_4874);
and \g448572/U$4 ( \11251 , RIee223a8_4848, \8486 );
nor \g448572/U$1 ( \11252 , \11249 , \11250 , \11251 );
and \g450828/U$2 ( \11253 , \8335 , RIded2c68_862);
and \g450828/U$3 ( \11254 , RIded9748_938, \8340 );
nor \g450828/U$1 ( \11255 , \11253 , \11254 );
and \g450823/U$2 ( \11256 , \8404 , RIee23320_4859);
and \g450823/U$3 ( \11257 , RIfcb7800_7110, \8351 );
nor \g450823/U$1 ( \11258 , \11256 , \11257 );
and \g455237/U$2 ( \11259 , \8313 , RIded53c8_890);
and \g455237/U$3 ( \11260 , RIfe804f0_7804, \8323 );
nor \g455237/U$1 ( \11261 , \11259 , \11260 );
not \g455236/U$1 ( \11262 , \11261 );
and \g449597/U$2 ( \11263 , \11262 , \8316 );
and \g449597/U$3 ( \11264 , RIfc98900_6758, \8359 );
nor \g449597/U$1 ( \11265 , \11263 , \11264 );
nand \g448140/U$1 ( \11266 , \11252 , \11255 , \11258 , \11265 );
and \g444754/U$3 ( \11267 , \8482 , \11266 );
nor \g444754/U$1 ( \11268 , \11248 , \11267 );
and \g446553/U$2 ( \11269 , \8964 , RIdee2c58_1044);
and \g446553/U$3 ( \11270 , RIfe80388_7803, \8966 );
nor \g446553/U$1 ( \11271 , \11269 , \11270 );
and \g446554/U$2 ( \11272 , \8521 , RIee212c8_4836);
and \g446554/U$3 ( \11273 , RIfcc8600_7302, \8525 );
nor \g446554/U$1 ( \11274 , \11272 , \11273 );
and \g446560/U$2 ( \11275 , \8974 , RIdedea40_997);
and \g446560/U$3 ( \11276 , RIfe80220_7802, \8976 );
nor \g446560/U$1 ( \11277 , \11275 , \11276 );
nand \g444453/U$1 ( \11278 , \11268 , \11271 , \11274 , \11277 );
and \g445744/U$2 ( \11279 , RIee36178_5074, \8417 );
and \g445744/U$3 ( \11280 , RIe14ea70_2272, \8356 );
and \g448551/U$2 ( \11281 , RIee37258_5086, \8371 );
and \g448551/U$3 ( \11282 , \8330 , RIe162570_2496);
and \g448551/U$4 ( \11283 , RIe151770_2304, \8488 );
nor \g448551/U$1 ( \11284 , \11281 , \11282 , \11283 );
and \g450765/U$2 ( \11285 , \8335 , RIe146370_2176);
and \g450765/U$3 ( \11286 , RIfce1290_7584, \8340 );
nor \g450765/U$1 ( \11287 , \11285 , \11286 );
and \g450760/U$2 ( \11288 , \8404 , RIe15f870_2464);
and \g450760/U$3 ( \11289 , RIe165270_2528, \8351 );
nor \g450760/U$1 ( \11290 , \11288 , \11289 );
and \g454242/U$2 ( \11291 , \8313 , RIe149070_2208);
and \g454242/U$3 ( \11292 , RIe14bd70_2240, \8323 );
nor \g454242/U$1 ( \11293 , \11291 , \11292 );
not \g454241/U$1 ( \11294 , \11293 );
and \g449577/U$2 ( \11295 , \11294 , \8316 );
and \g449577/U$3 ( \11296 , RIfc86fc0_6558, \8359 );
nor \g449577/U$1 ( \11297 , \11295 , \11296 );
nand \g448136/U$1 ( \11298 , \11284 , \11287 , \11290 , \11297 );
nor \g445744/U$1 ( \11299 , \11279 , \11280 , \11298 );
and \g450747/U$2 ( \11300 , \8378 , RIe154470_2336);
and \g450747/U$3 ( \11301 , RIfc4eff8_5921, \8523 );
nor \g450747/U$1 ( \11302 , \11300 , \11301 );
and \g450746/U$2 ( \11303 , \8414 , RIe157170_2368);
and \g450746/U$3 ( \11304 , RIe15cb70_2432, \8407 );
nor \g450746/U$1 ( \11305 , \11303 , \11304 );
and \g444956/U$2 ( \11306 , \11299 , \11302 , \11305 );
nor \g444956/U$1 ( \11307 , \11306 , \8368 );
and \g445751/U$2 ( \11308 , RIfe800b8_7801, \8417 );
and \g445751/U$3 ( \11309 , RIee2d640_4975, \8356 );
and \g448562/U$2 ( \11310 , RIdf31150_1935, \8319 );
and \g448562/U$3 ( \11311 , \8326 , RIdf331a8_1958);
and \g448562/U$4 ( \11312 , RIee2f800_4999, \8488 );
nor \g448562/U$1 ( \11313 , \11310 , \11311 , \11312 );
and \g450795/U$2 ( \11314 , \8335 , RIdf2ef90_1911);
and \g450795/U$3 ( \11315 , RIdf35638_1984, \8340 );
nor \g450795/U$1 ( \11316 , \11314 , \11315 );
and \g450791/U$2 ( \11317 , \8404 , RIee31150_5017);
and \g450791/U$3 ( \11318 , RIee34558_5054, \8351 );
nor \g450791/U$1 ( \11319 , \11317 , \11318 );
and \g454409/U$2 ( \11320 , \8313 , RIee320c8_5028);
and \g454409/U$3 ( \11321 , RIee331a8_5040, \8323 );
nor \g454409/U$1 ( \11322 , \11320 , \11321 );
not \g449587/U$3 ( \11323 , \11322 );
not \g449587/U$4 ( \11324 , \8328 );
and \g449587/U$2 ( \11325 , \11323 , \11324 );
and \g449587/U$5 ( \11326 , \8359 , RIfcc8330_7300);
nor \g449587/U$1 ( \11327 , \11325 , \11326 );
nand \g447485/U$1 ( \11328 , \11313 , \11316 , \11319 , \11327 );
nor \g445751/U$1 ( \11329 , \11308 , \11309 , \11328 );
and \g450783/U$2 ( \11330 , \8378 , RIfe7fde8_7799);
and \g450783/U$3 ( \11331 , RIfca0d30_6852, \8531 );
nor \g450783/U$1 ( \11332 , \11330 , \11331 );
and \g450780/U$2 ( \11333 , \8414 , RIdf3caf0_2067);
and \g450780/U$3 ( \11334 , RIfe7ff50_7800, \8409 );
nor \g450780/U$1 ( \11335 , \11333 , \11334 );
and \g444963/U$2 ( \11336 , \11329 , \11332 , \11335 );
nor \g444963/U$1 ( \11337 , \11336 , \8422 );
or \g444358/U$1 ( \11338 , \11218 , \11278 , \11307 , \11337 );
and \g445731/U$2 ( \11339 , RIfcaf808_7019, \8340 );
and \g445731/U$3 ( \11340 , RIdebf870_643, \8404 );
and \g448534/U$2 ( \11341 , RIfca5d58_6909, \8531 );
and \g448534/U$3 ( \11342 , \8486 , RIdeb1770_483);
and \g448534/U$4 ( \11343 , RIdec2570_675, \8383 );
nor \g448534/U$1 ( \11344 , \11341 , \11342 , \11343 );
and \g450702/U$2 ( \11345 , \8356 , RIdeaea70_451);
and \g450702/U$3 ( \11346 , RIfe7fc80_7798, \8359 );
nor \g450702/U$1 ( \11347 , \11345 , \11346 );
and \g454218/U$2 ( \11348 , \8313 , RIdeb9e70_579);
and \g454218/U$3 ( \11349 , RIdebcb70_611, \8323 );
nor \g454218/U$1 ( \11350 , \11348 , \11349 );
not \g449556/U$3 ( \11351 , \11350 );
not \g449556/U$4 ( \11352 , \8376 );
and \g449556/U$2 ( \11353 , \11351 , \11352 );
and \g449556/U$5 ( \11354 , \8351 , RIdec5270_707);
nor \g449556/U$1 ( \11355 , \11353 , \11354 );
and \g450697/U$2 ( \11356 , \8378 , RIdeb7170_547);
and \g450697/U$3 ( \11357 , RIfe7f848_7795, \8417 );
nor \g450697/U$1 ( \11358 , \11356 , \11357 );
nand \g447474/U$1 ( \11359 , \11344 , \11347 , \11355 , \11358 );
nor \g445731/U$1 ( \11360 , \11339 , \11340 , \11359 );
and \g450687/U$2 ( \11361 , \8335 , RIde9ced8_355);
and \g450687/U$3 ( \11362 , RIee1ff18_4822, \8371 );
nor \g450687/U$1 ( \11363 , \11361 , \11362 );
and \g450690/U$2 ( \11364 , \8319 , RIdea37d8_387);
and \g450690/U$3 ( \11365 , RIdeaa0d8_419, \8326 );
nor \g450690/U$1 ( \11366 , \11364 , \11365 );
and \g444950/U$2 ( \11367 , \11360 , \11363 , \11366 );
nor \g444950/U$1 ( \11368 , \11367 , \8589 );
and \g445738/U$2 ( \11369 , RIfcb0a50_7032, \8373 );
and \g445738/U$3 ( \11370 , RIe167ca0_2558, \8335 );
and \g448542/U$2 ( \11371 , RIfc82100_6502, \8523 );
and \g448542/U$3 ( \11372 , \8488 , RIfc52f40_5966);
and \g448542/U$4 ( \11373 , RIfcce438_7369, \8383 );
nor \g448542/U$1 ( \11374 , \11371 , \11372 , \11373 );
and \g450728/U$2 ( \11375 , \8356 , RIfca7108_6923);
and \g450728/U$3 ( \11376 , RIde81728_221, \8359 );
nor \g450728/U$1 ( \11377 , \11375 , \11376 );
and \g454900/U$2 ( \11378 , \8313 , RIde89720_260);
and \g454900/U$3 ( \11379 , RIfe7f9b0_7796, \8323 );
nor \g454900/U$1 ( \11380 , \11378 , \11379 );
not \g449566/U$3 ( \11381 , \11380 );
not \g449566/U$4 ( \11382 , \8376 );
and \g449566/U$2 ( \11383 , \11381 , \11382 );
and \g449566/U$5 ( \11384 , \8351 , RIfcdc3d0_7528);
nor \g449566/U$1 ( \11385 , \11383 , \11384 );
and \g450723/U$2 ( \11386 , \8378 , RIde85580_240);
and \g450723/U$3 ( \11387 , RIde90d40_296, \8417 );
nor \g450723/U$1 ( \11388 , \11386 , \11387 );
nand \g447478/U$1 ( \11389 , \11374 , \11377 , \11385 , \11388 );
nor \g445738/U$1 ( \11390 , \11369 , \11370 , \11389 );
and \g450719/U$2 ( \11391 , \8340 , RIfe7fb18_7797);
and \g450719/U$3 ( \11392 , RIfc75680_6358, \8404 );
nor \g450719/U$1 ( \11393 , \11391 , \11392 );
and \g450720/U$2 ( \11394 , \8319 , RIe169a28_2579);
and \g450720/U$3 ( \11395 , RIe16b648_2599, \8326 );
nor \g450720/U$1 ( \11396 , \11394 , \11395 );
and \g444955/U$2 ( \11397 , \11390 , \11393 , \11396 );
nor \g444955/U$1 ( \11398 , \11397 , \8558 );
or \g444266/U$1 ( \11399 , \11338 , \11368 , \11398 );
_DC \g27ec/U$1 ( \11400 , \11399 , \8654 );
and \g448730/U$2 ( \11401 , RIee34dc8_5060, \8531 );
and \g448730/U$3 ( \11402 , \8488 , RIe1514a0_2302);
and \g448730/U$4 ( \11403 , RIe1622a0_2494, \8330 );
nor \g448730/U$1 ( \11404 , \11401 , \11402 , \11403 );
and \g451363/U$2 ( \11405 , \8335 , RIe1460a0_2174);
and \g451363/U$3 ( \11406 , RIfc861b0_6548, \8340 );
nor \g451363/U$1 ( \11407 , \11405 , \11406 );
and \g454678/U$2 ( \11408 , \8313 , RIe148da0_2206);
and \g454678/U$3 ( \11409 , RIe14baa0_2238, \8323 );
nor \g454678/U$1 ( \11410 , \11408 , \11409 );
not \g454677/U$1 ( \11411 , \11410 );
and \g449757/U$2 ( \11412 , \11411 , \8316 );
and \g449757/U$3 ( \11413 , RIe164fa0_2526, \8351 );
nor \g449757/U$1 ( \11414 , \11412 , \11413 );
and \g451358/U$2 ( \11415 , \8356 , RIe14e7a0_2270);
and \g451358/U$3 ( \11416 , RIfe85c20_7866, \8359 );
nor \g451358/U$1 ( \11417 , \11415 , \11416 );
nand \g448156/U$1 ( \11418 , \11404 , \11407 , \11414 , \11417 );
and \g444763/U$2 ( \11419 , \11418 , \8369 );
and \g445891/U$2 ( \11420 , RIee2d4d8_4974, \8356 );
and \g445891/U$3 ( \11421 , RIdf35368_1982, \8340 );
and \g448748/U$2 ( \11422 , RIdf3c820_2065, \8414 );
and \g448748/U$3 ( \11423 , \8409 , RIdf3eb48_2090);
and \g448748/U$4 ( \11424 , RIee2f698_4998, \8488 );
nor \g448748/U$1 ( \11425 , \11422 , \11423 , \11424 );
and \g454401/U$2 ( \11426 , \8313 , RIfe857e8_7863);
and \g454401/U$3 ( \11427 , RIfe85518_7861, \8323 );
nor \g454401/U$1 ( \11428 , \11426 , \11427 );
not \g449776/U$3 ( \11429 , \11428 );
not \g449776/U$4 ( \11430 , \8328 );
and \g449776/U$2 ( \11431 , \11429 , \11430 );
and \g449776/U$5 ( \11432 , \8359 , RIfc9d4f0_6812);
nor \g449776/U$1 ( \11433 , \11431 , \11432 );
and \g451429/U$2 ( \11434 , \8404 , RIfe85680_7862);
and \g451429/U$3 ( \11435 , RIee343f0_5053, \8351 );
nor \g451429/U$1 ( \11436 , \11434 , \11435 );
and \g451438/U$2 ( \11437 , \8378 , RIdf3a660_2041);
and \g451438/U$3 ( \11438 , RIe140c40_2114, \8417 );
nor \g451438/U$1 ( \11439 , \11437 , \11438 );
nand \g447590/U$1 ( \11440 , \11425 , \11433 , \11436 , \11439 );
nor \g445891/U$1 ( \11441 , \11420 , \11421 , \11440 );
and \g451406/U$2 ( \11442 , \8335 , RIfe85ab8_7865);
and \g451406/U$3 ( \11443 , RIfc52298_5957, \8531 );
nor \g451406/U$1 ( \11444 , \11442 , \11443 );
and \g451400/U$2 ( \11445 , \8319 , RIdf30e80_1933);
and \g451400/U$3 ( \11446 , RIdf32ed8_1956, \8326 );
nor \g451400/U$1 ( \11447 , \11445 , \11446 );
and \g445066/U$2 ( \11448 , \11441 , \11444 , \11447 );
nor \g445066/U$1 ( \11449 , \11448 , \8422 );
nor \g444763/U$1 ( \11450 , \11419 , \11449 );
and \g446662/U$2 ( \11451 , \8426 , RIe15f5a0_2462);
and \g446662/U$3 ( \11452 , RIfe85950_7864, \8428 );
nor \g446662/U$1 ( \11453 , \11451 , \11452 );
and \g446661/U$2 ( \11454 , \8431 , RIe15c8a0_2430);
and \g446661/U$3 ( \11455 , RIee36010_5073, \8434 );
nor \g446661/U$1 ( \11456 , \11454 , \11455 );
and \g446664/U$2 ( \11457 , \8438 , RIe1541a0_2334);
and \g446664/U$3 ( \11458 , RIe156ea0_2366, \8440 );
nor \g446664/U$1 ( \11459 , \11457 , \11458 );
nand \g444469/U$1 ( \11460 , \11450 , \11453 , \11456 , \11459 );
and \g451536/U$2 ( \11461 , \8324 , RIdee6e70_1091);
and \g451536/U$3 ( \11462 , RIdf1cc78_1704, \8356 );
nor \g451536/U$1 ( \11463 , \11461 , \11462 );
and \g445922/U$2 ( \11464 , RIdf2c3f8_1880, \8523 );
and \g445922/U$3 ( \11465 , RIdedbbd8_964, \8319 );
and \g448788/U$2 ( \11466 , RIe16dda8_2627, \8412 );
and \g448788/U$3 ( \11467 , \8409 , RIde95f48_321);
and \g448788/U$4 ( \11468 , RIdf37d98_2012, \8488 );
nor \g448788/U$1 ( \11469 , \11466 , \11467 , \11468 );
and \g454680/U$2 ( \11470 , \8313 , RIdeca9a0_769);
and \g454680/U$3 ( \11471 , RIdecd6a0_801, \8323 );
nor \g454680/U$1 ( \11472 , \11470 , \11471 );
not \g449812/U$3 ( \11473 , \11472 );
not \g449812/U$4 ( \11474 , \8328 );
and \g449812/U$2 ( \11475 , \11473 , \11474 );
and \g449812/U$5 ( \11476 , \8359 , RIe1433a0_2142);
nor \g449812/U$1 ( \11477 , \11475 , \11476 );
and \g451560/U$2 ( \11478 , \8404 , RIdec7ca0_737);
and \g451560/U$3 ( \11479 , RIded03a0_833, \8351 );
nor \g451560/U$1 ( \11480 , \11478 , \11479 );
and \g451561/U$2 ( \11481 , \8378 , RIe159ba0_2398);
and \g451561/U$3 ( \11482 , RIdeb41a0_513, \8417 );
nor \g451561/U$1 ( \11483 , \11481 , \11482 );
nand \g447612/U$1 ( \11484 , \11469 , \11477 , \11480 , \11483 );
nor \g445922/U$1 ( \11485 , \11464 , \11465 , \11484 );
and \g451540/U$2 ( \11486 , \8335 , RIde7be90_194);
and \g451540/U$3 ( \11487 , RIdf00370_1379, \8340 );
nor \g451540/U$1 ( \11488 , \11486 , \11487 );
nand \g445556/U$1 ( \11489 , \11463 , \11485 , \11488 );
and \g444875/U$2 ( \11490 , \11489 , \9010 );
and \g448770/U$2 ( \11491 , RIfcd32f8_7425, \8531 );
and \g448770/U$3 ( \11492 , \8488 , RIee26b60_4899);
and \g448770/U$4 ( \11493 , RIee29f68_4936, \8330 );
nor \g448770/U$1 ( \11494 , \11491 , \11492 , \11493 );
and \g451496/U$2 ( \11495 , \8335 , RIfe84b40_7854);
and \g451496/U$3 ( \11496 , RIfc9e300_6822, \8340 );
nor \g451496/U$1 ( \11497 , \11495 , \11496 );
and \g454562/U$2 ( \11498 , \8313 , RIee25eb8_4890);
and \g454562/U$3 ( \11499 , RIdf1f540_1733, \8323 );
nor \g454562/U$1 ( \11500 , \11498 , \11499 );
not \g454561/U$1 ( \11501 , \11500 );
and \g449795/U$2 ( \11502 , \11501 , \8316 );
and \g449795/U$3 ( \11503 , RIee2b8b8_4954, \8351 );
nor \g449795/U$1 ( \11504 , \11502 , \11503 );
and \g451491/U$2 ( \11505 , \8356 , RIee265c0_4895);
and \g451491/U$3 ( \11506 , RIee27100_4903, \8359 );
nor \g451491/U$1 ( \11507 , \11505 , \11506 );
nand \g448162/U$1 ( \11508 , \11494 , \11497 , \11504 , \11507 );
and \g444875/U$3 ( \11509 , \8752 , \11508 );
nor \g444875/U$1 ( \11510 , \11490 , \11509 );
nor \g448424/U$1 ( \11511 , \8621 , \8425 );
and \g446695/U$2 ( \11512 , \11511 , RIee27970_4909);
nor \g448418/U$1 ( \11513 , \8621 , \8372 );
and \g446695/U$3 ( \11514 , RIee28bb8_4922, \11513 );
nor \g446695/U$1 ( \11515 , \11512 , \11514 );
nor \g448423/U$1 ( \11516 , \8621 , \8408 );
and \g446689/U$2 ( \11517 , \11516 , RIfe84e10_7856);
nor \g448411/U$1 ( \11518 , \8621 , \8433 );
and \g446689/U$3 ( \11519 , RIdf2a0d0_1855, \11518 );
nor \g446689/U$1 ( \11520 , \11517 , \11519 );
nor \g448443/U$1 ( \11521 , \8621 , \8437 );
and \g446698/U$2 ( \11522 , \11521 , RIfe84ca8_7855);
nor \g448442/U$1 ( \11523 , \8621 , \8413 );
and \g446698/U$3 ( \11524 , RIdf262f0_1811, \11523 );
nor \g446698/U$1 ( \11525 , \11522 , \11524 );
nand \g444578/U$1 ( \11526 , \11510 , \11515 , \11520 , \11525 );
and \g445841/U$2 ( \11527 , RIee1fdb0_4821, \8373 );
and \g445841/U$3 ( \11528 , RIdeb6ea0_545, \8378 );
and \g448683/U$2 ( \11529 , RIdea3148_385, \8319 );
and \g448683/U$3 ( \11530 , \8326 , RIdea9a48_417);
and \g448683/U$4 ( \11531 , RIdec22a0_673, \8383 );
nor \g448683/U$1 ( \11532 , \11529 , \11530 , \11531 );
and \g451218/U$2 ( \11533 , \8335 , RIde9c848_353);
and \g451218/U$3 ( \11534 , RIee1d920_4795, \8340 );
nor \g451218/U$1 ( \11535 , \11533 , \11534 );
and \g454568/U$2 ( \11536 , \8313 , RIee1e730_4805);
and \g454568/U$3 ( \11537 , RIdeb14a0_481, \8323 );
nor \g454568/U$1 ( \11538 , \11536 , \11537 );
not \g449708/U$3 ( \11539 , \11538 );
not \g449708/U$4 ( \11540 , \8347 );
and \g449708/U$2 ( \11541 , \11539 , \11540 );
and \g449708/U$5 ( \11542 , \8351 , RIdec4fa0_705);
nor \g449708/U$1 ( \11543 , \11541 , \11542 );
and \g451208/U$2 ( \11544 , \8356 , RIdeae7a0_449);
and \g451208/U$3 ( \11545 , RIee1ecd0_4809, \8359 );
nor \g451208/U$1 ( \11546 , \11544 , \11545 );
nand \g447558/U$1 ( \11547 , \11532 , \11535 , \11543 , \11546 );
nor \g445841/U$1 ( \11548 , \11527 , \11528 , \11547 );
and \g451193/U$2 ( \11549 , \8404 , RIdebf5a0_641);
and \g451193/U$3 ( \11550 , RIdebc8a0_609, \8409 );
nor \g451193/U$1 ( \11551 , \11549 , \11550 );
and \g451188/U$2 ( \11552 , \8414 , RIdeb9ba0_577);
and \g451188/U$3 ( \11553 , RIee1f270_4813, \8417 );
nor \g451188/U$1 ( \11554 , \11552 , \11553 );
and \g445030/U$2 ( \11555 , \11548 , \11551 , \11554 );
nor \g445030/U$1 ( \11556 , \11555 , \8589 );
and \g445858/U$2 ( \11557 , RIee199d8_4750, \8531 );
and \g445858/U$3 ( \11558 , RIe167b38_2557, \8335 );
and \g448703/U$2 ( \11559 , RIee1b1c0_4767, \8373 );
and \g448703/U$3 ( \11560 , \8383 , RIee1ba30_4773);
and \g448703/U$4 ( \11561 , RIfe853b0_7860, \8486 );
nor \g448703/U$1 ( \11562 , \11559 , \11560 , \11561 );
and \g454453/U$2 ( \11563 , \8313 , RIfea9cb0_8248);
and \g454453/U$3 ( \11564 , RIde8d230_278, \8323 );
nor \g454453/U$1 ( \11565 , \11563 , \11564 );
not \g449730/U$3 ( \11566 , \11565 );
not \g449730/U$4 ( \11567 , \8376 );
and \g449730/U$2 ( \11568 , \11566 , \11567 );
and \g449730/U$5 ( \11569 , \8359 , RIee1a3b0_4757);
nor \g449730/U$1 ( \11570 , \11568 , \11569 );
and \g451284/U$2 ( \11571 , \8404 , RIfec04b0_8308);
and \g451284/U$3 ( \11572 , RIee1cb10_4785, \8351 );
nor \g451284/U$1 ( \11573 , \11571 , \11572 );
and \g451293/U$2 ( \11574 , \8378 , RIfe84f78_7857);
and \g451293/U$3 ( \11575 , RIfe850e0_7858, \8417 );
nor \g451293/U$1 ( \11576 , \11574 , \11575 );
nand \g447566/U$1 ( \11577 , \11562 , \11570 , \11573 , \11576 );
nor \g445858/U$1 ( \11578 , \11557 , \11558 , \11577 );
and \g451258/U$2 ( \11579 , \8356 , RIfe85248_7859);
and \g451258/U$3 ( \11580 , RIee39148_5108, \8340 );
nor \g451258/U$1 ( \11581 , \11579 , \11580 );
and \g451268/U$2 ( \11582 , \8319 , RIee38608_5100);
and \g451268/U$3 ( \11583 , RIe16b378_2597, \8326 );
nor \g451268/U$1 ( \11584 , \11582 , \11583 );
and \g445045/U$2 ( \11585 , \11578 , \11581 , \11584 );
nor \g445045/U$1 ( \11586 , \11585 , \8558 );
or \g444387/U$1 ( \11587 , \11460 , \11526 , \11556 , \11586 );
and \g445813/U$2 ( \11588 , RIfc88eb0_6580, \8523 );
and \g445813/U$3 ( \11589 , RIded50f8_888, \8319 );
and \g448645/U$2 ( \11590 , RIee23cf8_4866, \8371 );
and \g448645/U$3 ( \11591 , \8383 , RIfcb54d8_7085);
and \g448645/U$4 ( \11592 , RIfcd43d8_7437, \8488 );
nor \g448645/U$1 ( \11593 , \11590 , \11591 , \11592 );
and \g454367/U$2 ( \11594 , \8313 , RIfec01e0_8306);
and \g454367/U$3 ( \11595 , RIdee2988_1042, \8323 );
nor \g454367/U$1 ( \11596 , \11594 , \11595 );
not \g449668/U$3 ( \11597 , \11596 );
not \g449668/U$4 ( \11598 , \8376 );
and \g449668/U$2 ( \11599 , \11597 , \11598 );
and \g449668/U$5 ( \11600 , \8359 , RIfcd7ee8_7479);
nor \g449668/U$1 ( \11601 , \11599 , \11600 );
and \g451078/U$2 ( \11602 , \8404 , RIfc54e30_5988);
and \g451078/U$3 ( \11603 , RIfec0348_8307, \8351 );
nor \g451078/U$1 ( \11604 , \11602 , \11603 );
and \g451084/U$2 ( \11605 , \8378 , RIdede770_995);
and \g451084/U$3 ( \11606 , RIfec0078_8305, \8417 );
nor \g451084/U$1 ( \11607 , \11605 , \11606 );
nand \g447531/U$1 ( \11608 , \11593 , \11601 , \11604 , \11607 );
nor \g445813/U$1 ( \11609 , \11588 , \11589 , \11608 );
and \g451062/U$2 ( \11610 , \8335 , RIfeab330_8264);
and \g451062/U$3 ( \11611 , RIded9478_936, \8340 );
nor \g451062/U$1 ( \11612 , \11610 , \11611 );
and \g451059/U$2 ( \11613 , \8324 , RIded6fe8_910);
and \g451059/U$3 ( \11614 , RIfc9e5d0_6824, \8356 );
nor \g451059/U$1 ( \11615 , \11613 , \11614 );
and \g445007/U$2 ( \11616 , \11609 , \11612 , \11615 );
nor \g445007/U$1 ( \11617 , \11616 , \8481 );
and \g445828/U$2 ( \11618 , RIdef7c70_1283, \8523 );
and \g445828/U$3 ( \11619 , RIdeec870_1155, \8319 );
and \g448663/U$2 ( \11620 , RIdf05d70_1443, \8412 );
and \g448663/U$3 ( \11621 , \8409 , RIdf08a70_1475);
and \g448663/U$4 ( \11622 , RIdefa970_1315, \8488 );
nor \g448663/U$1 ( \11623 , \11620 , \11621 , \11622 );
and \g454867/U$2 ( \11624 , \8313 , RIdf11170_1571);
and \g454867/U$3 ( \11625 , RIdf13e70_1603, \8323 );
nor \g454867/U$1 ( \11626 , \11624 , \11625 );
not \g449687/U$3 ( \11627 , \11626 );
not \g449687/U$4 ( \11628 , \8328 );
and \g449687/U$2 ( \11629 , \11627 , \11628 );
and \g449687/U$5 ( \11630 , \8359 , RIdefd670_1347);
nor \g449687/U$1 ( \11631 , \11629 , \11630 );
and \g451137/U$2 ( \11632 , \8404 , RIdf0e470_1539);
and \g451137/U$3 ( \11633 , RIdf16b70_1635, \8351 );
nor \g451137/U$1 ( \11634 , \11632 , \11633 );
and \g451148/U$2 ( \11635 , \8378 , RIdf03070_1411);
and \g451148/U$3 ( \11636 , RIdf0b770_1507, \8417 );
nor \g451148/U$1 ( \11637 , \11635 , \11636 );
nand \g447546/U$1 ( \11638 , \11623 , \11631 , \11634 , \11637 );
nor \g445828/U$1 ( \11639 , \11618 , \11619 , \11638 );
and \g451122/U$2 ( \11640 , \8335 , RIdee9b70_1123);
and \g451122/U$3 ( \11641 , RIdef2270_1219, \8340 );
nor \g451122/U$1 ( \11642 , \11640 , \11641 );
and \g451114/U$2 ( \11643 , \8326 , RIdeef570_1187);
and \g451114/U$3 ( \11644 , RIdef4f70_1251, \8356 );
nor \g451114/U$1 ( \11645 , \11643 , \11644 );
and \g445016/U$2 ( \11646 , \11639 , \11642 , \11645 );
nor \g445016/U$1 ( \11647 , \11646 , \8477 );
or \g444194/U$1 ( \11648 , \11587 , \11617 , \11647 );
_DC \g2871/U$1 ( \11649 , \11648 , \8654 );
and \g452285/U$2 ( \11650 , \8326 , RIe16b210_2596);
and \g452285/U$3 ( \11651 , RIfce4530_7620, \8356 );
nor \g452285/U$1 ( \11652 , \11650 , \11651 );
and \g446109/U$2 ( \11653 , RIfcd2d58_7421, \8531 );
and \g446109/U$3 ( \11654 , RIe1698c0_2578, \8317 );
and \g449022/U$2 ( \11655 , RIfe86d00_7878, \8414 );
and \g449022/U$3 ( \11656 , \8409 , RIde8cee8_277);
and \g449022/U$4 ( \11657 , RIfc8b8e0_6610, \8488 );
nor \g449022/U$1 ( \11658 , \11655 , \11656 , \11657 );
and \g454791/U$2 ( \11659 , \8313 , RIfc80918_6485);
and \g454791/U$3 ( \11660 , RIee1b8c8_4772, \8323 );
nor \g454791/U$1 ( \11661 , \11659 , \11660 );
not \g450034/U$3 ( \11662 , \11661 );
not \g450034/U$4 ( \11663 , \8328 );
and \g450034/U$2 ( \11664 , \11662 , \11663 );
and \g450034/U$5 ( \11665 , \8359 , RIde81098_219);
nor \g450034/U$1 ( \11666 , \11664 , \11665 );
and \g452297/U$2 ( \11667 , \8404 , RIfcdad50_7512);
and \g452297/U$3 ( \11668 , RIee1c9a8_4784, \8351 );
nor \g452297/U$1 ( \11669 , \11667 , \11668 );
and \g452303/U$2 ( \11670 , \8378 , RIfec0d20_8314);
and \g452303/U$3 ( \11671 , RIfe86e68_7879, \8417 );
nor \g452303/U$1 ( \11672 , \11670 , \11671 );
nand \g447736/U$1 ( \11673 , \11658 , \11666 , \11669 , \11672 );
nor \g446109/U$1 ( \11674 , \11653 , \11654 , \11673 );
and \g452290/U$2 ( \11675 , \8335 , RIe1679d0_2556);
and \g452290/U$3 ( \11676 , RIfc8ba48_6611, \8340 );
nor \g452290/U$1 ( \11677 , \11675 , \11676 );
nand \g445600/U$1 ( \11678 , \11652 , \11674 , \11677 );
and \g444745/U$2 ( \11679 , \11678 , \9700 );
and \g449010/U$2 ( \11680 , RIfcd9b08_7499, \8531 );
and \g449010/U$3 ( \11681 , \8488 , RIdeb1338_480);
and \g449010/U$4 ( \11682 , RIdec2138_672, \8383 );
nor \g449010/U$1 ( \11683 , \11680 , \11681 , \11682 );
and \g452268/U$2 ( \11684 , \8335 , RIde9c500_352);
and \g452268/U$3 ( \11685 , RIfc8b610_6608, \8340 );
nor \g452268/U$1 ( \11686 , \11684 , \11685 );
and \g454778/U$2 ( \11687 , \8313 , RIdea2e00_384);
and \g454778/U$3 ( \11688 , RIdea9700_416, \8323 );
nor \g454778/U$1 ( \11689 , \11687 , \11688 );
not \g454777/U$1 ( \11690 , \11689 );
and \g450022/U$2 ( \11691 , \11690 , \8316 );
and \g450022/U$3 ( \11692 , RIdec4e38_704, \8351 );
nor \g450022/U$1 ( \11693 , \11691 , \11692 );
and \g452263/U$2 ( \11694 , \8356 , RIdeae638_448);
and \g452263/U$3 ( \11695 , RIfc48ef0_5852, \8359 );
nor \g452263/U$1 ( \11696 , \11694 , \11695 );
nand \g448189/U$1 ( \11697 , \11683 , \11686 , \11693 , \11696 );
and \g444745/U$3 ( \11698 , \9702 , \11697 );
nor \g444745/U$1 ( \11699 , \11679 , \11698 );
nor \g448348/U$1 ( \11700 , \8589 , \8408 );
and \g446871/U$2 ( \11701 , \11700 , RIdebc738_608);
nor \g448347/U$1 ( \11702 , \8589 , \8433 );
and \g446871/U$3 ( \11703 , RIfc49490_5856, \11702 );
nor \g446871/U$1 ( \11704 , \11701 , \11703 );
and \g446873/U$2 ( \11705 , \9724 , RIdebf438_640);
and \g446873/U$3 ( \11706 , RIee1fc48_4820, \9726 );
nor \g446873/U$1 ( \11707 , \11705 , \11706 );
and \g446872/U$2 ( \11708 , \9170 , RIdeb6d38_544);
and \g446872/U$3 ( \11709 , RIdeb9a38_576, \9172 );
nor \g446872/U$1 ( \11710 , \11708 , \11709 );
nand \g444496/U$1 ( \11711 , \11699 , \11704 , \11707 , \11710 );
and \g452360/U$2 ( \11712 , \8378 , RIe159a38_2397);
and \g452360/U$3 ( \11713 , RIdf37c30_2011, \8488 );
nor \g452360/U$1 ( \11714 , \11712 , \11713 );
and \g446125/U$2 ( \11715 , RIe16dc40_2626, \8414 );
and \g446125/U$3 ( \11716 , RIdf2c290_1879, \8531 );
and \g449039/U$2 ( \11717 , RIde95c00_320, \8409 );
and \g449039/U$3 ( \11718 , \8373 , RIdeca838_768);
and \g449039/U$4 ( \11719 , RIdecd538_800, \8383 );
nor \g449039/U$1 ( \11720 , \11717 , \11718 , \11719 );
and \g452374/U$2 ( \11721 , \8335 , RIde7bb48_193);
and \g452374/U$3 ( \11722 , RIdf00208_1378, \8340 );
nor \g452374/U$1 ( \11723 , \11721 , \11722 );
and \g452369/U$2 ( \11724 , \8404 , RIdec7b38_736);
and \g452369/U$3 ( \11725 , RIded0238_832, \8351 );
nor \g452369/U$1 ( \11726 , \11724 , \11725 );
and \g454826/U$2 ( \11727 , \8313 , RIdedba70_963);
and \g454826/U$3 ( \11728 , RIdee6d08_1090, \8323 );
nor \g454826/U$1 ( \11729 , \11727 , \11728 );
not \g454825/U$1 ( \11730 , \11729 );
and \g450053/U$2 ( \11731 , \11730 , \8316 );
and \g450053/U$3 ( \11732 , RIdeb4038_512, \8417 );
nor \g450053/U$1 ( \11733 , \11731 , \11732 );
nand \g448194/U$1 ( \11734 , \11720 , \11723 , \11726 , \11733 );
nor \g446125/U$1 ( \11735 , \11715 , \11716 , \11734 );
and \g452358/U$2 ( \11736 , \8356 , RIdf1cb10_1703);
and \g452358/U$3 ( \11737 , RIe143238_2141, \8359 );
nor \g452358/U$1 ( \11738 , \11736 , \11737 );
nand \g445604/U$1 ( \11739 , \11714 , \11735 , \11738 );
and \g444878/U$2 ( \11740 , \11739 , \9010 );
and \g449032/U$2 ( \11741 , RIdf26188_1810, \8412 );
and \g449032/U$3 ( \11742 , \8409 , RIdf27da8_1830);
and \g449032/U$4 ( \11743 , RIdf1f3d8_1732, \8326 );
nor \g449032/U$1 ( \11744 , \11741 , \11742 , \11743 );
and \g452340/U$2 ( \11745 , \8356 , RIfc475a0_5834);
and \g452340/U$3 ( \11746 , RIfc8cb28_6623, \8359 );
nor \g452340/U$1 ( \11747 , \11745 , \11746 );
and \g454811/U$2 ( \11748 , \8313 , RIdf22948_1770);
and \g454811/U$3 ( \11749 , RIfcdb188_7515, \8323 );
nor \g454811/U$1 ( \11750 , \11748 , \11749 );
not \g450044/U$3 ( \11751 , \11750 );
not \g450044/U$4 ( \11752 , \8347 );
and \g450044/U$2 ( \11753 , \11751 , \11752 );
and \g450044/U$5 ( \11754 , \8340 , RIdf21430_1755);
nor \g450044/U$1 ( \11755 , \11753 , \11754 );
and \g452335/U$2 ( \11756 , \8378 , RIdf24568_1790);
and \g452335/U$3 ( \11757 , RIdf29f68_1854, \8417 );
nor \g452335/U$1 ( \11758 , \11756 , \11757 );
nand \g447740/U$1 ( \11759 , \11744 , \11747 , \11755 , \11758 );
and \g444878/U$3 ( \11760 , \8752 , \11759 );
nor \g444878/U$1 ( \11761 , \11740 , \11760 );
nor \g448426/U$1 ( \11762 , \8621 , \8508 );
and \g446890/U$2 ( \11763 , \11762 , RIfe868c8_7875);
nor \g448425/U$1 ( \11764 , \8621 , \8318 );
and \g446890/U$3 ( \11765 , RIfec0bb8_8313, \11764 );
nor \g446890/U$1 ( \11766 , \11763 , \11765 );
nor \g448420/U$1 ( \11767 , \8621 , \8382 );
and \g446889/U$2 ( \11768 , \11767 , RIfc8c858_6621);
nor \g448412/U$1 ( \11769 , \8621 , \9295 );
and \g446889/U$3 ( \11770 , RIfcd2a88_7419, \11769 );
nor \g446889/U$1 ( \11771 , \11768 , \11770 );
and \g446891/U$2 ( \11772 , \11511 , RIfcd6430_7460);
and \g446891/U$3 ( \11773 , RIfc47ca8_5839, \11513 );
nor \g446891/U$1 ( \11774 , \11772 , \11773 );
nand \g444613/U$1 ( \11775 , \11761 , \11766 , \11771 , \11774 );
and \g446084/U$2 ( \11776 , RIfc48518_5845, \8531 );
and \g446084/U$3 ( \11777 , RIe148c38_2205, \8319 );
and \g448990/U$2 ( \11778 , RIee370f0_5085, \8373 );
and \g448990/U$3 ( \11779 , \8330 , RIe162138_2493);
and \g448990/U$4 ( \11780 , RIe151338_2301, \8488 );
nor \g448990/U$1 ( \11781 , \11778 , \11779 , \11780 );
and \g454406/U$2 ( \11782 , \8313 , RIe156d38_2365);
and \g454406/U$3 ( \11783 , RIe15c738_2429, \8323 );
nor \g454406/U$1 ( \11784 , \11782 , \11783 );
not \g450002/U$3 ( \11785 , \11784 );
not \g450002/U$4 ( \11786 , \8376 );
and \g450002/U$2 ( \11787 , \11785 , \11786 );
and \g450002/U$5 ( \11788 , \8359 , RIfc3f260_5744);
nor \g450002/U$1 ( \11789 , \11787 , \11788 );
and \g452193/U$2 ( \11790 , \8404 , RIe15f438_2461);
and \g452193/U$3 ( \11791 , RIe164e38_2525, \8351 );
nor \g452193/U$1 ( \11792 , \11790 , \11791 );
and \g452197/U$2 ( \11793 , \8378 , RIe154038_2333);
and \g452197/U$3 ( \11794 , RIfc999e0_6770, \8417 );
nor \g452197/U$1 ( \11795 , \11793 , \11794 );
nand \g447720/U$1 ( \11796 , \11781 , \11789 , \11792 , \11795 );
nor \g446084/U$1 ( \11797 , \11776 , \11777 , \11796 );
and \g452179/U$2 ( \11798 , \8335 , RIe145f38_2173);
and \g452179/U$3 ( \11799 , RIfc99e18_6773, \8340 );
nor \g452179/U$1 ( \11800 , \11798 , \11799 );
and \g452178/U$2 ( \11801 , \8326 , RIe14b938_2237);
and \g452178/U$3 ( \11802 , RIe14e638_2269, \8356 );
nor \g452178/U$1 ( \11803 , \11801 , \11802 );
and \g445211/U$2 ( \11804 , \11797 , \11800 , \11803 );
nor \g445211/U$1 ( \11805 , \11804 , \8368 );
and \g446092/U$2 ( \11806 , RIee2d370_4973, \8356 );
and \g446092/U$3 ( \11807 , RIfcc3470_7244, \8359 );
and \g449000/U$2 ( \11808 , RIfec0ff0_8316, \8326 );
and \g449000/U$3 ( \11809 , \8373 , RIee31f60_5027);
and \g449000/U$4 ( \11810 , RIee33040_5039, \8383 );
nor \g449000/U$1 ( \11811 , \11808 , \11809 , \11810 );
and \g454762/U$2 ( \11812 , \8313 , RIfe86a30_7876);
and \g454762/U$3 ( \11813 , RIdf3e9e0_2089, \8323 );
nor \g454762/U$1 ( \11814 , \11812 , \11813 );
not \g450011/U$3 ( \11815 , \11814 );
not \g450011/U$4 ( \11816 , \8376 );
and \g450011/U$2 ( \11817 , \11815 , \11816 );
and \g450011/U$5 ( \11818 , \8340 , RIdf35200_1981);
nor \g450011/U$1 ( \11819 , \11817 , \11818 );
and \g452229/U$2 ( \11820 , \8404 , RIfcd99a0_7498);
and \g452229/U$3 ( \11821 , RIee34288_5052, \8351 );
nor \g452229/U$1 ( \11822 , \11820 , \11821 );
and \g452230/U$2 ( \11823 , \8378 , RIdf3a4f8_2040);
and \g452230/U$3 ( \11824 , RIfe86b98_7877, \8417 );
nor \g452230/U$1 ( \11825 , \11823 , \11824 );
nand \g447726/U$1 ( \11826 , \11811 , \11819 , \11822 , \11825 );
nor \g446092/U$1 ( \11827 , \11806 , \11807 , \11826 );
and \g452218/U$2 ( \11828 , \8335 , RIfec0e88_8315);
and \g452218/U$3 ( \11829 , RIee2f530_4997, \8488 );
nor \g452218/U$1 ( \11830 , \11828 , \11829 );
and \g452213/U$2 ( \11831 , \8317 , RIdf30d18_1932);
and \g452213/U$3 ( \11832 , RIfc7fdd8_6477, \8531 );
nor \g452213/U$1 ( \11833 , \11831 , \11832 );
and \g445221/U$2 ( \11834 , \11827 , \11830 , \11833 );
nor \g445221/U$1 ( \11835 , \11834 , \8422 );
or \g444369/U$1 ( \11836 , \11711 , \11775 , \11805 , \11835 );
and \g446055/U$2 ( \11837 , RIfcc3038_7241, \8531 );
and \g446055/U$3 ( \11838 , RIded4f90_887, \8319 );
and \g448959/U$2 ( \11839 , RIee23b90_4865, \8373 );
and \g448959/U$3 ( \11840 , \8383 , RIee246d0_4873);
and \g448959/U$4 ( \11841 , RIfc98a68_6759, \8488 );
nor \g448959/U$1 ( \11842 , \11839 , \11840 , \11841 );
and \g455132/U$2 ( \11843 , \8313 , RIdee0930_1019);
and \g455132/U$3 ( \11844 , RIdee2820_1041, \8323 );
nor \g455132/U$1 ( \11845 , \11843 , \11844 );
not \g449974/U$3 ( \11846 , \11845 );
not \g449974/U$4 ( \11847 , \8376 );
and \g449974/U$2 ( \11848 , \11846 , \11847 );
and \g449974/U$5 ( \11849 , \8359 , RIfc55da8_5999);
nor \g449974/U$1 ( \11850 , \11848 , \11849 );
and \g452081/U$2 ( \11851 , \8404 , RIee231b8_4858);
and \g452081/U$3 ( \11852 , RIee254e0_4883, \8351 );
nor \g452081/U$1 ( \11853 , \11851 , \11852 );
and \g452086/U$2 ( \11854 , \8378 , RIdede608_994);
and \g452086/U$3 ( \11855 , RIfe86fd0_7880, \8417 );
nor \g452086/U$1 ( \11856 , \11854 , \11855 );
nand \g447702/U$1 ( \11857 , \11842 , \11850 , \11853 , \11856 );
nor \g446055/U$1 ( \11858 , \11837 , \11838 , \11857 );
and \g452067/U$2 ( \11859 , \8335 , RIded2b00_861);
and \g452067/U$3 ( \11860 , RIded9310_935, \8340 );
nor \g452067/U$1 ( \11861 , \11859 , \11860 );
and \g452059/U$2 ( \11862 , \8326 , RIded6e80_909);
and \g452059/U$3 ( \11863 , RIfc464c0_5822, \8356 );
nor \g452059/U$1 ( \11864 , \11862 , \11863 );
and \g445188/U$2 ( \11865 , \11858 , \11861 , \11864 );
nor \g445188/U$1 ( \11866 , \11865 , \8481 );
and \g446071/U$2 ( \11867 , RIdf16a08_1634, \8351 );
and \g446071/U$3 ( \11868 , RIdee9a08_1122, \8335 );
and \g448977/U$2 ( \11869 , RIdf05c08_1442, \8414 );
and \g448977/U$3 ( \11870 , \8409 , RIdf08908_1474);
and \g448977/U$4 ( \11871 , RIdeef408_1186, \8326 );
nor \g448977/U$1 ( \11872 , \11869 , \11870 , \11871 );
and \g452144/U$2 ( \11873 , \8356 , RIdef4e08_1250);
and \g452144/U$3 ( \11874 , RIdefd508_1346, \8359 );
nor \g452144/U$1 ( \11875 , \11873 , \11874 );
and \g454603/U$2 ( \11876 , \8313 , RIdef7b08_1282);
and \g454603/U$3 ( \11877 , RIdefa808_1314, \8323 );
nor \g454603/U$1 ( \11878 , \11876 , \11877 );
not \g449990/U$3 ( \11879 , \11878 );
not \g449990/U$4 ( \11880 , \8347 );
and \g449990/U$2 ( \11881 , \11879 , \11880 );
and \g449990/U$5 ( \11882 , \8340 , RIdef2108_1218);
nor \g449990/U$1 ( \11883 , \11881 , \11882 );
and \g452063/U$2 ( \11884 , \8378 , RIdf02f08_1410);
and \g452063/U$3 ( \11885 , RIdf0b608_1506, \8417 );
nor \g452063/U$1 ( \11886 , \11884 , \11885 );
nand \g447712/U$1 ( \11887 , \11872 , \11875 , \11883 , \11886 );
nor \g446071/U$1 ( \11888 , \11867 , \11868 , \11887 );
and \g452122/U$2 ( \11889 , \8317 , RIdeec708_1154);
and \g452122/U$3 ( \11890 , RIdf0e308_1538, \8404 );
nor \g452122/U$1 ( \11891 , \11889 , \11890 );
and \g453854/U$2 ( \11892 , \8373 , RIdf11008_1570);
and \g453854/U$3 ( \11893 , RIdf13d08_1602, \8383 );
nor \g453854/U$1 ( \11894 , \11892 , \11893 );
and \g445202/U$2 ( \11895 , \11888 , \11891 , \11894 );
nor \g445202/U$1 ( \11896 , \11895 , \8477 );
or \g444200/U$1 ( \11897 , \11836 , \11866 , \11896 );
_DC \g28f6/U$1 ( \11898 , \11897 , \8654 );
and \g451964/U$2 ( \11899 , \8404 , RIfcecac8_7715);
and \g451964/U$3 ( \11900 , RIdee26b8_1040, \8409 );
nor \g451964/U$1 ( \11901 , \11899 , \11900 );
and \g446029/U$2 ( \11902 , RIfc931d0_6696, \8371 );
and \g446029/U$3 ( \11903 , RIdede4a0_993, \8378 );
and \g448953/U$2 ( \11904 , RIfc792f8_6401, \8531 );
and \g448953/U$3 ( \11905 , \8486 , RIfcbf528_7199);
and \g448953/U$4 ( \11906 , RIfc5b640_6062, \8383 );
nor \g448953/U$1 ( \11907 , \11904 , \11905 , \11906 );
and \g452003/U$2 ( \11908 , \8335 , RIded2998_860);
and \g452003/U$3 ( \11909 , RIded91a8_934, \8340 );
nor \g452003/U$1 ( \11910 , \11908 , \11909 );
and \g454523/U$2 ( \11911 , \8313 , RIded4e28_886);
and \g454523/U$3 ( \11912 , RIded6d18_908, \8323 );
nor \g454523/U$1 ( \11913 , \11911 , \11912 );
not \g454522/U$1 ( \11914 , \11913 );
and \g449957/U$2 ( \11915 , \11914 , \8316 );
and \g449957/U$3 ( \11916 , RIfc5b7a8_6063, \8351 );
nor \g449957/U$1 ( \11917 , \11915 , \11916 );
and \g451997/U$2 ( \11918 , \8356 , RIfc93068_6695);
and \g451997/U$3 ( \11919 , RIfcbf0f0_7196, \8359 );
nor \g451997/U$1 ( \11920 , \11918 , \11919 );
nand \g448183/U$1 ( \11921 , \11907 , \11910 , \11917 , \11920 );
nor \g446029/U$1 ( \11922 , \11902 , \11903 , \11921 );
and \g451913/U$2 ( \11923 , \8412 , RIdee07c8_1018);
and \g451913/U$3 ( \11924 , RIdee4710_1063, \8417 );
nor \g451913/U$1 ( \11925 , \11923 , \11924 );
nand \g445576/U$1 ( \11926 , \11901 , \11922 , \11925 );
and \g444827/U$2 ( \11927 , \11926 , \8482 );
and \g448878/U$2 ( \11928 , RIdf10ea0_1569, \8373 );
and \g448878/U$3 ( \11929 , \8383 , RIdf13ba0_1601);
and \g448878/U$4 ( \11930 , RIdefa6a0_1313, \8488 );
nor \g448878/U$1 ( \11931 , \11928 , \11929 , \11930 );
and \g454583/U$2 ( \11932 , \8313 , RIdf05aa0_1441);
and \g454583/U$3 ( \11933 , RIdf087a0_1473, \8323 );
nor \g454583/U$1 ( \11934 , \11932 , \11933 );
not \g449893/U$3 ( \11935 , \11934 );
not \g449893/U$4 ( \11936 , \8376 );
and \g449893/U$2 ( \11937 , \11935 , \11936 );
and \g449893/U$5 ( \11938 , \8359 , RIdefd3a0_1345);
nor \g449893/U$1 ( \11939 , \11937 , \11938 );
and \g453258/U$2 ( \11940 , \8404 , RIdf0e1a0_1537);
and \g453258/U$3 ( \11941 , RIdf168a0_1633, \8351 );
nor \g453258/U$1 ( \11942 , \11940 , \11941 );
and \g451813/U$2 ( \11943 , \8378 , RIdf02da0_1409);
and \g451813/U$3 ( \11944 , RIdf0b4a0_1505, \8417 );
nor \g451813/U$1 ( \11945 , \11943 , \11944 );
nand \g447640/U$1 ( \11946 , \11931 , \11939 , \11942 , \11945 );
and \g444827/U$3 ( \11947 , \8478 , \11946 );
nor \g444827/U$1 ( \11948 , \11927 , \11947 );
and \g446732/U$2 ( \11949 , \8775 , RIdef4ca0_1249);
and \g446732/U$3 ( \11950 , RIdef79a0_1281, \8777 );
nor \g446732/U$1 ( \11951 , \11949 , \11950 );
and \g446740/U$2 ( \11952 , \8780 , RIdeef2a0_1185);
and \g446740/U$3 ( \11953 , RIdef1fa0_1217, \8782 );
nor \g446740/U$1 ( \11954 , \11952 , \11953 );
and \g446753/U$2 ( \11955 , \8785 , RIdee98a0_1121);
and \g446753/U$3 ( \11956 , RIdeec5a0_1153, \8787 );
nor \g446753/U$1 ( \11957 , \11955 , \11956 );
nand \g444572/U$1 ( \11958 , \11948 , \11951 , \11954 , \11957 );
and \g451396/U$2 ( \11959 , \8319 , RIfc43220_5786);
and \g451396/U$3 ( \11960 , RIfea9e18_8249, \8326 );
nor \g451396/U$1 ( \11961 , \11959 , \11960 );
and \g445904/U$2 ( \11962 , RIee195a0_4747, \8356 );
and \g445904/U$3 ( \11963 , RIfcbe718_7189, \8340 );
and \g448791/U$2 ( \11964 , RIfe82f20_7834, \8414 );
and \g448791/U$3 ( \11965 , \8409 , RIde8cba0_276);
and \g448791/U$4 ( \11966 , RIfe831f0_7836, \8488 );
nor \g448791/U$1 ( \11967 , \11964 , \11965 , \11966 );
and \g454967/U$2 ( \11968 , \8313 , RIfe83088_7835);
and \g454967/U$3 ( \11969 , RIfc7af18_6421, \8323 );
nor \g454967/U$1 ( \11970 , \11968 , \11969 );
not \g449806/U$3 ( \11971 , \11970 );
not \g449806/U$4 ( \11972 , \8328 );
and \g449806/U$2 ( \11973 , \11971 , \11972 );
and \g449806/U$5 ( \11974 , \8359 , RIee1a248_4756);
nor \g449806/U$1 ( \11975 , \11973 , \11974 );
and \g451483/U$2 ( \11976 , \8404 , RIee1a950_4761);
and \g451483/U$3 ( \11977 , RIfc90ea8_6671, \8351 );
nor \g451483/U$1 ( \11978 , \11976 , \11977 );
and \g451518/U$2 ( \11979 , \8378 , RIfe82db8_7833);
and \g451518/U$3 ( \11980 , RIde906b0_294, \8417 );
nor \g451518/U$1 ( \11981 , \11979 , \11980 );
nand \g447599/U$1 ( \11982 , \11967 , \11975 , \11978 , \11981 );
nor \g445904/U$1 ( \11983 , \11962 , \11963 , \11982 );
and \g451431/U$2 ( \11984 , \8335 , RIe167868_2555);
and \g451431/U$3 ( \11985 , RIfcc2390_7232, \8523 );
nor \g451431/U$1 ( \11986 , \11984 , \11985 );
nand \g445549/U$1 ( \11987 , \11961 , \11983 , \11986 );
and \g444744/U$2 ( \11988 , \11987 , \9700 );
and \g448716/U$2 ( \11989 , RIee1e5c8_4804, \8531 );
and \g448716/U$3 ( \11990 , \8488 , RIdeb11d0_479);
and \g448716/U$4 ( \11991 , RIdec1fd0_671, \8383 );
nor \g448716/U$1 ( \11992 , \11989 , \11990 , \11991 );
and \g451255/U$2 ( \11993 , \8335 , RIde9c1b8_351);
and \g451255/U$3 ( \11994 , RIfc437c0_5790, \8340 );
nor \g451255/U$1 ( \11995 , \11993 , \11994 );
and \g455384/U$2 ( \11996 , \8313 , RIdea2ab8_383);
and \g455384/U$3 ( \11997 , RIdea93b8_415, \8323 );
nor \g455384/U$1 ( \11998 , \11996 , \11997 );
not \g455383/U$1 ( \11999 , \11998 );
and \g449722/U$2 ( \12000 , \11999 , \8316 );
and \g449722/U$3 ( \12001 , RIdec4cd0_703, \8351 );
nor \g449722/U$1 ( \12002 , \12000 , \12001 );
and \g451234/U$2 ( \12003 , \8356 , RIdeae4d0_447);
and \g451234/U$3 ( \12004 , RIfe83358_7837, \8359 );
nor \g451234/U$1 ( \12005 , \12003 , \12004 );
nand \g448151/U$1 ( \12006 , \11992 , \11995 , \12002 , \12005 );
and \g444744/U$3 ( \12007 , \9702 , \12006 );
nor \g444744/U$1 ( \12008 , \11988 , \12007 );
and \g446610/U$2 ( \12009 , \11700 , RIdebc5d0_607);
and \g446610/U$3 ( \12010 , RIfc7b1e8_6423, \11702 );
nor \g446610/U$1 ( \12011 , \12009 , \12010 );
and \g446627/U$2 ( \12012 , \9724 , RIdebf2d0_639);
and \g446627/U$3 ( \12013 , RIfc7b4b8_6425, \9726 );
nor \g446627/U$1 ( \12014 , \12012 , \12013 );
and \g446618/U$2 ( \12015 , \9170 , RIdeb6bd0_543);
and \g446618/U$3 ( \12016 , RIdeb98d0_575, \9172 );
nor \g446618/U$1 ( \12017 , \12015 , \12016 );
nand \g444459/U$1 ( \12018 , \12008 , \12011 , \12014 , \12017 );
and \g445730/U$2 ( \12019 , RIee36f88_5084, \8373 );
and \g445730/U$3 ( \12020 , RIe156bd0_2364, \8412 );
and \g448553/U$2 ( \12021 , RIfebfda8_8303, \8523 );
and \g448553/U$3 ( \12022 , \8486 , RIe1511d0_2300);
and \g448553/U$4 ( \12023 , RIe161fd0_2492, \8330 );
nor \g448553/U$1 ( \12024 , \12021 , \12022 , \12023 );
and \g450705/U$2 ( \12025 , \8335 , RIe145dd0_2172);
and \g450705/U$3 ( \12026 , RIfebfc40_8302, \8340 );
nor \g450705/U$1 ( \12027 , \12025 , \12026 );
and \g454765/U$2 ( \12028 , \8313 , RIe148ad0_2204);
and \g454765/U$3 ( \12029 , RIe14b7d0_2236, \8323 );
nor \g454765/U$1 ( \12030 , \12028 , \12029 );
not \g454764/U$1 ( \12031 , \12030 );
and \g449563/U$2 ( \12032 , \12031 , \8316 );
and \g449563/U$3 ( \12033 , RIe164cd0_2524, \8351 );
nor \g449563/U$1 ( \12034 , \12032 , \12033 );
and \g450682/U$2 ( \12035 , \8356 , RIe14e4d0_2268);
and \g450682/U$3 ( \12036 , RIfe83628_7839, \8359 );
nor \g450682/U$1 ( \12037 , \12035 , \12036 );
nand \g448135/U$1 ( \12038 , \12024 , \12027 , \12034 , \12037 );
nor \g445730/U$1 ( \12039 , \12019 , \12020 , \12038 );
and \g450582/U$2 ( \12040 , \8404 , RIe15f2d0_2460);
and \g450582/U$3 ( \12041 , RIee35ea8_5072, \8417 );
nor \g450582/U$1 ( \12042 , \12040 , \12041 );
and \g450608/U$2 ( \12043 , \8378 , RIe153ed0_2332);
and \g450608/U$3 ( \12044 , RIe15c5d0_2428, \8409 );
nor \g450608/U$1 ( \12045 , \12043 , \12044 );
and \g444929/U$2 ( \12046 , \12039 , \12042 , \12045 );
nor \g444929/U$1 ( \12047 , \12046 , \8368 );
and \g445786/U$2 ( \12048 , RIfc96a10_6736, \8356 );
and \g445786/U$3 ( \12049 , RIdf35098_1980, \8340 );
and \g448624/U$2 ( \12050 , RIee31df8_5026, \8373 );
and \g448624/U$3 ( \12051 , \8383 , RIee32ed8_5038);
and \g448624/U$4 ( \12052 , RIfc91e20_6682, \8488 );
nor \g448624/U$1 ( \12053 , \12050 , \12051 , \12052 );
and \g454336/U$2 ( \12054 , \8313 , RIfe834c0_7838);
and \g454336/U$3 ( \12055 , RIdf3e878_2088, \8323 );
nor \g454336/U$1 ( \12056 , \12054 , \12055 );
not \g449642/U$3 ( \12057 , \12056 );
not \g449642/U$4 ( \12058 , \8376 );
and \g449642/U$2 ( \12059 , \12057 , \12058 );
and \g449642/U$5 ( \12060 , \8359 , RIfc5a6c8_6051);
nor \g449642/U$1 ( \12061 , \12059 , \12060 );
and \g450939/U$2 ( \12062 , \8404 , RIfcc1f58_7229);
and \g450939/U$3 ( \12063 , RIee34120_5051, \8351 );
nor \g450939/U$1 ( \12064 , \12062 , \12063 );
and \g450967/U$2 ( \12065 , \8378 , RIdf3a390_2039);
and \g450967/U$3 ( \12066 , RIe140ad8_2113, \8417 );
nor \g450967/U$1 ( \12067 , \12065 , \12066 );
nand \g447511/U$1 ( \12068 , \12053 , \12061 , \12064 , \12067 );
nor \g445786/U$1 ( \12069 , \12048 , \12049 , \12068 );
and \g450869/U$2 ( \12070 , \8335 , RIfeab768_8267);
and \g450869/U$3 ( \12071 , RIee2e888_4988, \8523 );
nor \g450869/U$1 ( \12072 , \12070 , \12071 );
and \g450838/U$2 ( \12073 , \8319 , RIdf30bb0_1931);
and \g450838/U$3 ( \12074 , RIfeab600_8266, \8324 );
nor \g450838/U$1 ( \12075 , \12073 , \12074 );
and \g444971/U$2 ( \12076 , \12069 , \12072 , \12075 );
nor \g444971/U$1 ( \12077 , \12076 , \8422 );
or \g444360/U$1 ( \12078 , \11958 , \12018 , \12047 , \12077 );
and \g446392/U$2 ( \12079 , RIfcbe9e8_7191, \8351 );
and \g446392/U$3 ( \12080 , RIfc92258_6685, \8404 );
and \g449438/U$2 ( \12081 , RIfc79730_6404, \8317 );
and \g449438/U$3 ( \12082 , \8326 , RIdf1f270_1731);
and \g449438/U$4 ( \12083 , RIfc5add0_6056, \8488 );
nor \g449438/U$1 ( \12084 , \12081 , \12082 , \12083 );
and \g455409/U$2 ( \12085 , \8313 , RIdf26020_1809);
and \g455409/U$3 ( \12086 , RIfea95a8_8243, \8323 );
nor \g455409/U$1 ( \12087 , \12085 , \12086 );
not \g450436/U$3 ( \12088 , \12087 );
not \g450436/U$4 ( \12089 , \8376 );
and \g450436/U$2 ( \12090 , \12088 , \12089 );
and \g450436/U$5 ( \12091 , \8359 , RIfc79a00_6406);
nor \g450436/U$1 ( \12092 , \12090 , \12091 );
and \g453760/U$2 ( \12093 , \8335 , RIdf19000_1661);
and \g453760/U$3 ( \12094 , RIfce3018_7605, \8340 );
nor \g453760/U$1 ( \12095 , \12093 , \12094 );
and \g453711/U$2 ( \12096 , \8378 , RIdf24400_1789);
and \g453711/U$3 ( \12097 , RIfea7118_8217, \8417 );
nor \g453711/U$1 ( \12098 , \12096 , \12097 );
nand \g447948/U$1 ( \12099 , \12084 , \12092 , \12095 , \12098 );
nor \g446392/U$1 ( \12100 , \12079 , \12080 , \12099 );
and \g453640/U$2 ( \12101 , \8356 , RIfc92690_6688);
and \g453640/U$3 ( \12102 , RIfc79fa0_6410, \8383 );
nor \g453640/U$1 ( \12103 , \12101 , \12102 );
and \g453620/U$2 ( \12104 , \8531 , RIfce5d18_7637);
and \g453620/U$3 ( \12105 , RIfc96740_6734, \8373 );
nor \g453620/U$1 ( \12106 , \12104 , \12105 );
and \g445419/U$2 ( \12107 , \12100 , \12103 , \12106 );
nor \g445419/U$1 ( \12108 , \12107 , \8621 );
and \g446452/U$2 ( \12109 , RIdf2c128_1878, \8531 );
and \g446452/U$3 ( \12110 , RIdedb908_962, \8319 );
and \g449502/U$2 ( \12111 , RIdeca6d0_767, \8373 );
and \g449502/U$3 ( \12112 , \8330 , RIdecd3d0_799);
and \g449502/U$4 ( \12113 , RIdf37ac8_2010, \8488 );
nor \g449502/U$1 ( \12114 , \12111 , \12112 , \12113 );
and \g454871/U$2 ( \12115 , \8313 , RIe16dad8_2625);
and \g454871/U$3 ( \12116 , RIde958b8_319, \8323 );
nor \g454871/U$1 ( \12117 , \12115 , \12116 );
not \g450514/U$3 ( \12118 , \12117 );
not \g450514/U$4 ( \12119 , \8376 );
and \g450514/U$2 ( \12120 , \12118 , \12119 );
and \g450514/U$5 ( \12121 , \8359 , RIe1430d0_2140);
nor \g450514/U$1 ( \12122 , \12120 , \12121 );
and \g453994/U$2 ( \12123 , \8404 , RIdec79d0_735);
and \g453994/U$3 ( \12124 , RIded00d0_831, \8351 );
nor \g453994/U$1 ( \12125 , \12123 , \12124 );
and \g454033/U$2 ( \12126 , \8378 , RIe1598d0_2396);
and \g454033/U$3 ( \12127 , RIdeb3ed0_511, \8417 );
nor \g454033/U$1 ( \12128 , \12126 , \12127 );
nand \g447985/U$1 ( \12129 , \12114 , \12122 , \12125 , \12128 );
nor \g446452/U$1 ( \12130 , \12109 , \12110 , \12129 );
and \g453910/U$2 ( \12131 , \8335 , RIde7b800_192);
and \g453910/U$3 ( \12132 , RIdf000a0_1377, \8340 );
nor \g453910/U$1 ( \12133 , \12131 , \12132 );
and \g453882/U$2 ( \12134 , \8326 , RIdee6ba0_1089);
and \g453882/U$3 ( \12135 , RIdf1c9a8_1702, \8356 );
nor \g453882/U$1 ( \12136 , \12134 , \12135 );
and \g445449/U$2 ( \12137 , \12130 , \12133 , \12136 );
nor \g445449/U$1 ( \12138 , \12137 , \8651 );
or \g444187/U$1 ( \12139 , \12078 , \12108 , \12138 );
_DC \g297b/U$1 ( \12140 , \12139 , \8654 );
and \g446663/U$2 ( \12141 , \11213 , RIdf1c840_1701);
and \g446663/U$3 ( \12142 , RIdf2bfc0_1877, \11215 );
nor \g446663/U$1 ( \12143 , \12141 , \12142 );
and \g445888/U$2 ( \12144 , RIdf37960_2009, \8488 );
and \g445888/U$3 ( \12145 , RIe142f68_2139, \8359 );
and \g448755/U$2 ( \12146 , RIde95570_318, \8409 );
and \g448755/U$3 ( \12147 , \8373 , RIdeca568_766);
and \g448755/U$4 ( \12148 , RIdecd268_798, \8383 );
nor \g448755/U$1 ( \12149 , \12146 , \12147 , \12148 );
and \g451437/U$2 ( \12150 , \8335 , RIde7b4b8_191);
and \g451437/U$3 ( \12151 , RIdefff38_1376, \8340 );
nor \g451437/U$1 ( \12152 , \12150 , \12151 );
and \g451420/U$2 ( \12153 , \8404 , RIdec7868_734);
and \g451420/U$3 ( \12154 , RIdecff68_830, \8351 );
nor \g451420/U$1 ( \12155 , \12153 , \12154 );
and \g454847/U$2 ( \12156 , \8313 , RIdedb7a0_961);
and \g454847/U$3 ( \12157 , RIdee6a38_1088, \8323 );
nor \g454847/U$1 ( \12158 , \12156 , \12157 );
not \g454846/U$1 ( \12159 , \12158 );
and \g449778/U$2 ( \12160 , \12159 , \8316 );
and \g449778/U$3 ( \12161 , RIdeb3d68_510, \8417 );
nor \g449778/U$1 ( \12162 , \12160 , \12161 );
nand \g448159/U$1 ( \12163 , \12149 , \12152 , \12155 , \12162 );
nor \g445888/U$1 ( \12164 , \12144 , \12145 , \12163 );
not \g444847/U$3 ( \12165 , \12164 );
not \g444847/U$4 ( \12166 , \8651 );
and \g444847/U$2 ( \12167 , \12165 , \12166 );
and \g445916/U$2 ( \12168 , RIfcb08e8_7031, \8351 );
and \g445916/U$3 ( \12169 , RIdf18e98_1660, \8335 );
and \g448792/U$2 ( \12170 , RIfeaa520_8254, \8326 );
and \g448792/U$3 ( \12171 , \8531 , RIdf227e0_1769);
and \g448792/U$4 ( \12172 , RIfcee850_7736, \8488 );
nor \g448792/U$1 ( \12173 , \12170 , \12171 , \12172 );
and \g450660/U$2 ( \12174 , \8356 , RIfc5efe8_6103);
and \g450660/U$3 ( \12175 , RIfc5ed18_6101, \8359 );
nor \g450660/U$1 ( \12176 , \12174 , \12175 );
and \g454588/U$2 ( \12177 , \8313 , RIdf25eb8_1808);
and \g454588/U$3 ( \12178 , RIdf27c40_1829, \8323 );
nor \g454588/U$1 ( \12179 , \12177 , \12178 );
not \g449813/U$3 ( \12180 , \12179 );
not \g449813/U$4 ( \12181 , \8376 );
and \g449813/U$2 ( \12182 , \12180 , \12181 );
and \g449813/U$5 ( \12183 , \8340 , RIdf212c8_1754);
nor \g449813/U$1 ( \12184 , \12182 , \12183 );
and \g451547/U$2 ( \12185 , \8378 , RIdf24298_1788);
and \g451547/U$3 ( \12186 , RIdf29e00_1853, \8417 );
nor \g451547/U$1 ( \12187 , \12185 , \12186 );
nand \g447611/U$1 ( \12188 , \12173 , \12176 , \12184 , \12187 );
nor \g445916/U$1 ( \12189 , \12168 , \12169 , \12188 );
and \g451514/U$2 ( \12190 , \8319 , RIdf1ad88_1682);
and \g451514/U$3 ( \12191 , RIfcdef68_7559, \8404 );
nor \g451514/U$1 ( \12192 , \12190 , \12191 );
and \g451501/U$2 ( \12193 , \8373 , RIfc95ed0_6728);
and \g451501/U$3 ( \12194 , RIfcee418_7733, \8383 );
nor \g451501/U$1 ( \12195 , \12193 , \12194 );
and \g445079/U$2 ( \12196 , \12189 , \12192 , \12195 );
nor \g445079/U$1 ( \12197 , \12196 , \8621 );
nor \g444847/U$1 ( \12198 , \12167 , \12197 );
and \g446676/U$2 ( \12199 , \9031 , RIe159768_2395);
and \g446676/U$3 ( \12200 , RIe16d970_2624, \9033 );
nor \g446676/U$1 ( \12201 , \12199 , \12200 );
nand \g444421/U$1 ( \12202 , \12143 , \12198 , \12201 );
and \g448833/U$2 ( \12203 , RIe169758_2577, \8319 );
and \g448833/U$3 ( \12204 , \8324 , RIe16b0a8_2595);
and \g448833/U$4 ( \12205 , RIde8c858_275, \8409 );
nor \g448833/U$1 ( \12206 , \12203 , \12204 , \12205 );
and \g451359/U$2 ( \12207 , \8335 , RIe167700_2554);
and \g451359/U$3 ( \12208 , RIfcedfe0_7730, \8340 );
nor \g451359/U$1 ( \12209 , \12207 , \12208 );
and \g451677/U$2 ( \12210 , \8404 , RIfcec0f0_7708);
and \g451677/U$3 ( \12211 , RIfced4a0_7722, \8351 );
nor \g451677/U$1 ( \12212 , \12210 , \12211 );
and \g454657/U$2 ( \12213 , \8313 , RIfc95930_6724);
and \g454657/U$3 ( \12214 , RIfcc1418_7221, \8323 );
nor \g454657/U$1 ( \12215 , \12213 , \12214 );
not \g449851/U$3 ( \12216 , \12215 );
not \g449851/U$4 ( \12217 , \8328 );
and \g449851/U$2 ( \12218 , \12216 , \12217 );
and \g449851/U$5 ( \12219 , \8417 , RIde90368_293);
nor \g449851/U$1 ( \12220 , \12218 , \12219 );
nand \g447631/U$1 ( \12221 , \12206 , \12209 , \12212 , \12220 );
and \g444681/U$2 ( \12222 , \12221 , \9700 );
and \g445976/U$2 ( \12223 , RIdec4b68_702, \8351 );
and \g445976/U$3 ( \12224 , RIde9be70_350, \8335 );
and \g448868/U$2 ( \12225 , RIdea9070_414, \8326 );
and \g448868/U$3 ( \12226 , \8523 , RIfcc12b0_7220);
and \g448868/U$4 ( \12227 , RIdeb1068_478, \8486 );
nor \g448868/U$1 ( \12228 , \12225 , \12226 , \12227 );
and \g451805/U$2 ( \12229 , \8356 , RIdeae368_446);
and \g451805/U$3 ( \12230 , RIfc75ef0_6364, \8359 );
nor \g451805/U$1 ( \12231 , \12229 , \12230 );
and \g455052/U$2 ( \12232 , \8313 , RIdeb9768_574);
and \g455052/U$3 ( \12233 , RIdebc468_606, \8323 );
nor \g455052/U$1 ( \12234 , \12232 , \12233 );
not \g449886/U$3 ( \12235 , \12234 );
not \g449886/U$4 ( \12236 , \8376 );
and \g449886/U$2 ( \12237 , \12235 , \12236 );
and \g449886/U$5 ( \12238 , \8340 , RIfc5e340_6094);
nor \g449886/U$1 ( \12239 , \12237 , \12238 );
and \g451793/U$2 ( \12240 , \8378 , RIdeb6a68_542);
and \g451793/U$3 ( \12241 , RIfce6df8_7649, \8417 );
nor \g451793/U$1 ( \12242 , \12240 , \12241 );
nand \g447650/U$1 ( \12243 , \12228 , \12231 , \12239 , \12242 );
nor \g445976/U$1 ( \12244 , \12223 , \12224 , \12243 );
and \g451767/U$2 ( \12245 , \8319 , RIdea2770_382);
and \g451767/U$3 ( \12246 , RIdebf168_638, \8404 );
nor \g451767/U$1 ( \12247 , \12245 , \12246 );
and \g451752/U$2 ( \12248 , \8373 , RIfc5df08_6091);
and \g451752/U$3 ( \12249 , RIdec1e68_670, \8330 );
nor \g451752/U$1 ( \12250 , \12248 , \12249 );
and \g445132/U$2 ( \12251 , \12244 , \12247 , \12250 );
nor \g445132/U$1 ( \12252 , \12251 , \8589 );
nor \g444681/U$1 ( \12253 , \12222 , \12252 );
nor \g448255/U$1 ( \12254 , \8558 , \8437 );
and \g446727/U$2 ( \12255 , \12254 , RIde84ef0_238);
nor \g448287/U$1 ( \12256 , \8558 , \8413 );
and \g446727/U$3 ( \12257 , RIde893d8_259, \12256 );
nor \g446727/U$1 ( \12258 , \12255 , \12257 );
nor \g448286/U$1 ( \12259 , \8558 , \8487 );
and \g446724/U$2 ( \12260 , \12259 , RIfc95a98_6725);
nor \g448285/U$1 ( \12261 , \8558 , \10292 );
and \g446724/U$3 ( \12262 , RIde80d50_218, \12261 );
nor \g446724/U$1 ( \12263 , \12260 , \12262 );
nor \g448256/U$1 ( \12264 , \8558 , \8520 );
and \g446738/U$2 ( \12265 , \12264 , RIfced1d0_7720);
nor \g448295/U$1 ( \12266 , \8558 , \8524 );
and \g446738/U$3 ( \12267 , RIfced068_7719, \12266 );
nor \g446738/U$1 ( \12268 , \12265 , \12267 );
nand \g444476/U$1 ( \12269 , \12253 , \12258 , \12263 , \12268 );
and \g445822/U$2 ( \12270 , RIfccfef0_7388, \8351 );
and \g445822/U$3 ( \12271 , RIfcafda8_7023, \8404 );
and \g448668/U$2 ( \12272 , RIdf3c6b8_2064, \8414 );
and \g448668/U$3 ( \12273 , \8409 , RIdf3e710_2087);
and \g448668/U$4 ( \12274 , RIfebf100_8294, \8326 );
nor \g448668/U$1 ( \12275 , \12272 , \12273 , \12274 );
and \g451144/U$2 ( \12276 , \8356 , RIee2d208_4972);
and \g451144/U$3 ( \12277 , RIfc5fc90_6112, \8359 );
nor \g451144/U$1 ( \12278 , \12276 , \12277 );
and \g454801/U$2 ( \12279 , \8313 , RIfc742d0_6344);
and \g454801/U$3 ( \12280 , RIee2f3c8_4996, \8323 );
nor \g454801/U$1 ( \12281 , \12279 , \12280 );
not \g449689/U$3 ( \12282 , \12281 );
not \g449689/U$4 ( \12283 , \8347 );
and \g449689/U$2 ( \12284 , \12282 , \12283 );
and \g449689/U$5 ( \12285 , \8340 , RIdf34f30_1979);
nor \g449689/U$1 ( \12286 , \12284 , \12285 );
and \g451129/U$2 ( \12287 , \8378 , RIdf3a228_2038);
and \g451129/U$3 ( \12288 , RIe140970_2112, \8417 );
nor \g451129/U$1 ( \12289 , \12287 , \12288 );
nand \g447542/U$1 ( \12290 , \12275 , \12278 , \12286 , \12289 );
nor \g445822/U$1 ( \12291 , \12270 , \12271 , \12290 );
and \g451101/U$2 ( \12292 , \8335 , RIdf2ecc0_1909);
and \g451101/U$3 ( \12293 , RIfca57b8_6905, \8383 );
nor \g451101/U$1 ( \12294 , \12292 , \12293 );
and \g451085/U$2 ( \12295 , \8319 , RIdf30a48_1930);
and \g451085/U$3 ( \12296 , RIfc600c8_6115, \8373 );
nor \g451085/U$1 ( \12297 , \12295 , \12296 );
and \g445013/U$2 ( \12298 , \12291 , \12294 , \12297 );
nor \g445013/U$1 ( \12299 , \12298 , \8422 );
and \g445853/U$2 ( \12300 , RIe153d68_2331, \8378 );
and \g445853/U$3 ( \12301 , RIfe82818_7829, \8359 );
and \g448708/U$2 ( \12302 , RIe148968_2203, \8319 );
and \g448708/U$3 ( \12303 , \8324 , RIe14b668_2235);
and \g448708/U$4 ( \12304 , RIe15c468_2427, \8407 );
nor \g448708/U$1 ( \12305 , \12302 , \12303 , \12304 );
and \g451280/U$2 ( \12306 , \8335 , RIe145c68_2171);
and \g451280/U$3 ( \12307 , RIfc5f9c0_6110, \8340 );
nor \g451280/U$1 ( \12308 , \12306 , \12307 );
and \g451274/U$2 ( \12309 , \8404 , RIe15f168_2459);
and \g451274/U$3 ( \12310 , RIe164b68_2523, \8351 );
nor \g451274/U$1 ( \12311 , \12309 , \12310 );
and \g454373/U$2 ( \12312 , \8313 , RIee36e20_5083);
and \g454373/U$3 ( \12313 , RIe161e68_2491, \8323 );
nor \g454373/U$1 ( \12314 , \12312 , \12313 );
not \g449731/U$3 ( \12315 , \12314 );
not \g449731/U$4 ( \12316 , \8328 );
and \g449731/U$2 ( \12317 , \12315 , \12316 );
and \g449731/U$5 ( \12318 , \8417 , RIfc426e0_5778);
nor \g449731/U$1 ( \12319 , \12317 , \12318 );
nand \g447564/U$1 ( \12320 , \12305 , \12308 , \12311 , \12319 );
nor \g445853/U$1 ( \12321 , \12300 , \12301 , \12320 );
and \g451230/U$2 ( \12322 , \8356 , RIe14e368_2267);
and \g451230/U$3 ( \12323 , RIe156a68_2363, \8414 );
nor \g451230/U$1 ( \12324 , \12322 , \12323 );
and \g451216/U$2 ( \12325 , \8531 , RIee34c60_5059);
and \g451216/U$3 ( \12326 , RIe151068_2299, \8488 );
nor \g451216/U$1 ( \12327 , \12325 , \12326 );
and \g445034/U$2 ( \12328 , \12321 , \12324 , \12327 );
nor \g445034/U$1 ( \12329 , \12328 , \8368 );
or \g444302/U$1 ( \12330 , \12202 , \12269 , \12299 , \12329 );
and \g445767/U$2 ( \12331 , RIdee0660_1017, \8414 );
and \g445767/U$3 ( \12332 , RIfc73a60_6338, \8356 );
and \g448599/U$2 ( \12333 , RIdee2550_1039, \8409 );
and \g448599/U$3 ( \12334 , \8371 , RIfc60aa0_6122);
and \g448599/U$4 ( \12335 , RIfccfd88_7387, \8383 );
nor \g448599/U$1 ( \12336 , \12333 , \12334 , \12335 );
and \g450891/U$2 ( \12337 , \8335 , RIded2830_859);
and \g450891/U$3 ( \12338 , RIfe82980_7830, \8340 );
nor \g450891/U$1 ( \12339 , \12337 , \12338 );
and \g450879/U$2 ( \12340 , \8404 , RIfca5ec0_6910);
and \g450879/U$3 ( \12341 , RIfcc96e0_7314, \8351 );
nor \g450879/U$1 ( \12342 , \12340 , \12341 );
and \g454156/U$2 ( \12343 , \8313 , RIded4cc0_885);
and \g454156/U$3 ( \12344 , RIded6bb0_907, \8323 );
nor \g454156/U$1 ( \12345 , \12343 , \12344 );
not \g454155/U$1 ( \12346 , \12345 );
and \g449620/U$2 ( \12347 , \12346 , \8316 );
and \g449620/U$3 ( \12348 , RIdee45a8_1062, \8417 );
nor \g449620/U$1 ( \12349 , \12347 , \12348 );
nand \g448143/U$1 ( \12350 , \12336 , \12339 , \12342 , \12349 );
nor \g445767/U$1 ( \12351 , \12331 , \12332 , \12350 );
and \g450846/U$2 ( \12352 , \8378 , RIfe826b0_7828);
and \g450846/U$3 ( \12353 , RIfcdeb30_7556, \8359 );
nor \g450846/U$1 ( \12354 , \12352 , \12353 );
and \g450832/U$2 ( \12355 , \8523 , RIfca5bf0_6908);
and \g450832/U$3 ( \12356 , RIfc73bc8_6339, \8488 );
nor \g450832/U$1 ( \12357 , \12355 , \12356 );
and \g444973/U$2 ( \12358 , \12351 , \12354 , \12357 );
nor \g444973/U$1 ( \12359 , \12358 , \8481 );
and \g445795/U$2 ( \12360 , RIdf02c38_1408, \8378 );
and \g445795/U$3 ( \12361 , RIdefd238_1344, \8359 );
and \g448636/U$2 ( \12362 , RIdeec438_1152, \8319 );
and \g448636/U$3 ( \12363 , \8324 , RIdeef138_1184);
and \g448636/U$4 ( \12364 , RIdf08638_1472, \8409 );
nor \g448636/U$1 ( \12365 , \12362 , \12363 , \12364 );
and \g451015/U$2 ( \12366 , \8335 , RIdee9738_1120);
and \g451015/U$3 ( \12367 , RIdef1e38_1216, \8340 );
nor \g451015/U$1 ( \12368 , \12366 , \12367 );
and \g451005/U$2 ( \12369 , \8404 , RIdf0e038_1536);
and \g451005/U$3 ( \12370 , RIdf16738_1632, \8351 );
nor \g451005/U$1 ( \12371 , \12369 , \12370 );
and \g454433/U$2 ( \12372 , \8313 , RIdf10d38_1568);
and \g454433/U$3 ( \12373 , RIdf13a38_1600, \8323 );
nor \g454433/U$1 ( \12374 , \12372 , \12373 );
not \g449653/U$3 ( \12375 , \12374 );
not \g449653/U$4 ( \12376 , \8328 );
and \g449653/U$2 ( \12377 , \12375 , \12376 );
and \g449653/U$5 ( \12378 , \8417 , RIdf0b338_1504);
nor \g449653/U$1 ( \12379 , \12377 , \12378 );
nand \g447521/U$1 ( \12380 , \12365 , \12368 , \12371 , \12379 );
nor \g445795/U$1 ( \12381 , \12360 , \12361 , \12380 );
and \g450976/U$2 ( \12382 , \8356 , RIdef4b38_1248);
and \g450976/U$3 ( \12383 , RIdf05938_1440, \8414 );
nor \g450976/U$1 ( \12384 , \12382 , \12383 );
and \g450971/U$2 ( \12385 , \8531 , RIdef7838_1280);
and \g450971/U$3 ( \12386 , RIdefa538_1312, \8488 );
nor \g450971/U$1 ( \12387 , \12385 , \12386 );
and \g444994/U$2 ( \12388 , \12381 , \12384 , \12387 );
nor \g444994/U$1 ( \12389 , \12388 , \8477 );
or \g444177/U$1 ( \12390 , \12330 , \12359 , \12389 );
_DC \g2a00/U$1 ( \12391 , \12390 , \8654 );
and \g448888/U$2 ( \12392 , RIfc65c30_6180, \8319 );
and \g448888/U$3 ( \12393 , \8324 , RIe16af40_2594);
and \g448888/U$4 ( \12394 , RIde8c510_274, \8409 );
nor \g448888/U$1 ( \12395 , \12392 , \12393 , \12394 );
and \g451888/U$2 ( \12396 , \8335 , RIe167598_2553);
and \g451888/U$3 ( \12397 , RIfc51488_5947, \8340 );
nor \g451888/U$1 ( \12398 , \12396 , \12397 );
and \g453300/U$2 ( \12399 , \8404 , RIfe8b8f0_7932);
and \g453300/U$3 ( \12400 , RIfc6fc80_6294, \8351 );
nor \g453300/U$1 ( \12401 , \12399 , \12400 );
and \g454570/U$2 ( \12402 , \8313 , RIfca8080_6934);
and \g454570/U$3 ( \12403 , RIee1b760_4771, \8323 );
nor \g454570/U$1 ( \12404 , \12402 , \12403 );
not \g449910/U$3 ( \12405 , \12404 );
not \g449910/U$4 ( \12406 , \8328 );
and \g449910/U$2 ( \12407 , \12405 , \12406 );
and \g449910/U$5 ( \12408 , \8417 , RIde90020_292);
nor \g449910/U$1 ( \12409 , \12407 , \12408 );
nand \g447663/U$1 ( \12410 , \12395 , \12398 , \12401 , \12409 );
and \g444683/U$2 ( \12411 , \12410 , \9700 );
and \g446008/U$2 ( \12412 , RIdec4a00_701, \8351 );
and \g446008/U$3 ( \12413 , RIde9bb28_349, \8335 );
and \g448890/U$2 ( \12414 , RIdea8d28_413, \8324 );
and \g448890/U$3 ( \12415 , \8523 , RIfc657f8_6177);
and \g448890/U$4 ( \12416 , RIdeb0f00_477, \8488 );
nor \g448890/U$1 ( \12417 , \12414 , \12415 , \12416 );
and \g451893/U$2 ( \12418 , \8356 , RIdeae200_445);
and \g451893/U$3 ( \12419 , RIfc6f9b0_6292, \8359 );
nor \g451893/U$1 ( \12420 , \12418 , \12419 );
and \g454731/U$2 ( \12421 , \8313 , RIdeb9600_573);
and \g454731/U$3 ( \12422 , RIdebc300_605, \8323 );
nor \g454731/U$1 ( \12423 , \12421 , \12422 );
not \g449912/U$3 ( \12424 , \12423 );
not \g449912/U$4 ( \12425 , \8376 );
and \g449912/U$2 ( \12426 , \12424 , \12425 );
and \g449912/U$5 ( \12427 , \8340 , RIfce69c0_7646);
nor \g449912/U$1 ( \12428 , \12426 , \12427 );
and \g451892/U$2 ( \12429 , \8378 , RIdeb6900_541);
and \g451892/U$3 ( \12430 , RIfc64cb8_6169, \8417 );
nor \g451892/U$1 ( \12431 , \12429 , \12430 );
nand \g447664/U$1 ( \12432 , \12417 , \12420 , \12428 , \12431 );
nor \g446008/U$1 ( \12433 , \12412 , \12413 , \12432 );
and \g451890/U$2 ( \12434 , \8319 , RIdea2428_381);
and \g451890/U$3 ( \12435 , RIdebf000_637, \8404 );
nor \g451890/U$1 ( \12436 , \12434 , \12435 );
and \g453223/U$2 ( \12437 , \8371 , RIfcad7b0_6996);
and \g453223/U$3 ( \12438 , RIdec1d00_669, \8383 );
nor \g453223/U$1 ( \12439 , \12437 , \12438 );
and \g445157/U$2 ( \12440 , \12433 , \12436 , \12439 );
nor \g445157/U$1 ( \12441 , \12440 , \8589 );
nor \g444683/U$1 ( \12442 , \12411 , \12441 );
and \g446794/U$2 ( \12443 , \12254 , RIde84ba8_237);
and \g446794/U$3 ( \12444 , RIde89090_258, \12256 );
nor \g446794/U$1 ( \12445 , \12443 , \12444 );
and \g446792/U$2 ( \12446 , \12259 , RIfcad210_6992);
and \g446792/U$3 ( \12447 , RIfc65ac8_6179, \12261 );
nor \g446792/U$1 ( \12448 , \12446 , \12447 );
and \g446795/U$2 ( \12449 , \12264 , RIfcce2d0_7368);
and \g446795/U$3 ( \12450 , RIfcce168_7367, \12266 );
nor \g446795/U$1 ( \12451 , \12449 , \12450 );
nand \g444483/U$1 ( \12452 , \12442 , \12445 , \12448 , \12451 );
and \g448892/U$2 ( \12453 , RIe15c300_2426, \8409 );
and \g448892/U$3 ( \12454 , \8373 , RIfc66e78_6193);
and \g448892/U$4 ( \12455 , RIe161d00_2490, \8383 );
nor \g448892/U$1 ( \12456 , \12453 , \12454 , \12455 );
and \g451898/U$2 ( \12457 , \8335 , RIe145b00_2170);
and \g451898/U$3 ( \12458 , RIfc6e1c8_6275, \8340 );
nor \g451898/U$1 ( \12459 , \12457 , \12458 );
and \g451897/U$2 ( \12460 , \8404 , RIe15f000_2458);
and \g451897/U$3 ( \12461 , RIe164a00_2522, \8351 );
nor \g451897/U$1 ( \12462 , \12460 , \12461 );
and \g454567/U$2 ( \12463 , \8313 , RIe148800_2202);
and \g454567/U$3 ( \12464 , RIe14b500_2234, \8323 );
nor \g454567/U$1 ( \12465 , \12463 , \12464 );
not \g454566/U$1 ( \12466 , \12465 );
and \g449914/U$2 ( \12467 , \12466 , \8316 );
and \g449914/U$3 ( \12468 , RIfc6e498_6277, \8417 );
nor \g449914/U$1 ( \12469 , \12467 , \12468 );
nand \g448181/U$1 ( \12470 , \12456 , \12459 , \12462 , \12469 );
and \g444769/U$2 ( \12471 , \12470 , \8369 );
and \g446010/U$2 ( \12472 , RIee33fb8_5050, \8351 );
and \g446010/U$3 ( \12473 , RIee30fe8_5016, \8404 );
and \g448893/U$2 ( \12474 , RIdf3c550_2063, \8414 );
and \g448893/U$3 ( \12475 , \8409 , RIdf3e5a8_2086);
and \g448893/U$4 ( \12476 , RIdf32d70_1955, \8324 );
nor \g448893/U$1 ( \12477 , \12474 , \12475 , \12476 );
and \g451904/U$2 ( \12478 , \8356 , RIfc6e600_6278);
and \g451904/U$3 ( \12479 , RIfc6e060_6274, \8359 );
nor \g451904/U$1 ( \12480 , \12478 , \12479 );
and \g455372/U$2 ( \12481 , \8313 , RIfc56078_6001);
and \g455372/U$3 ( \12482 , RIfcac6d0_6984, \8323 );
nor \g455372/U$1 ( \12483 , \12481 , \12482 );
not \g449916/U$3 ( \12484 , \12483 );
not \g449916/U$4 ( \12485 , \8347 );
and \g449916/U$2 ( \12486 , \12484 , \12485 );
and \g449916/U$5 ( \12487 , \8340 , RIdf34dc8_1978);
nor \g449916/U$1 ( \12488 , \12486 , \12487 );
and \g451902/U$2 ( \12489 , \8378 , RIfea8798_8233);
and \g451902/U$3 ( \12490 , RIfea8630_8232, \8417 );
nor \g451902/U$1 ( \12491 , \12489 , \12490 );
nand \g447665/U$1 ( \12492 , \12477 , \12480 , \12488 , \12491 );
nor \g446010/U$1 ( \12493 , \12472 , \12473 , \12492 );
and \g452845/U$2 ( \12494 , \8335 , RIdf2eb58_1908);
and \g452845/U$3 ( \12495 , RIee32d70_5037, \8383 );
nor \g452845/U$1 ( \12496 , \12494 , \12495 );
and \g451899/U$2 ( \12497 , \8319 , RIfea84c8_8231);
and \g451899/U$3 ( \12498 , RIee31c90_5025, \8371 );
nor \g451899/U$1 ( \12499 , \12497 , \12498 );
and \g445159/U$2 ( \12500 , \12493 , \12496 , \12499 );
nor \g445159/U$1 ( \12501 , \12500 , \8422 );
nor \g444769/U$1 ( \12502 , \12471 , \12501 );
and \g446797/U$2 ( \12503 , \8438 , RIe153c00_2330);
and \g446797/U$3 ( \12504 , RIe156900_2362, \8440 );
nor \g446797/U$1 ( \12505 , \12503 , \12504 );
nor \g448401/U$1 ( \12506 , \8368 , \8487 );
and \g446798/U$2 ( \12507 , \12506 , RIe150f00_2298);
nor \g448321/U$1 ( \12508 , \8368 , \10292 );
and \g446798/U$3 ( \12509 , RIfc6e330_6276, \12508 );
nor \g446798/U$1 ( \12510 , \12507 , \12509 );
and \g446799/U$2 ( \12511 , \8717 , RIe14e200_2266);
and \g446799/U$3 ( \12512 , RIfccda60_7362, \8719 );
nor \g446799/U$1 ( \12513 , \12511 , \12512 );
nand \g444484/U$1 ( \12514 , \12502 , \12505 , \12510 , \12513 );
and \g446005/U$2 ( \12515 , RIdf057d0_1439, \8414 );
and \g446005/U$3 ( \12516 , RIdef49d0_1247, \8356 );
and \g448884/U$2 ( \12517 , RIdf084d0_1471, \8407 );
and \g448884/U$3 ( \12518 , \8373 , RIdf10bd0_1567);
and \g448884/U$4 ( \12519 , RIdf138d0_1599, \8383 );
nor \g448884/U$1 ( \12520 , \12517 , \12518 , \12519 );
and \g451879/U$2 ( \12521 , \8335 , RIdee95d0_1119);
and \g451879/U$3 ( \12522 , RIdef1cd0_1215, \8340 );
nor \g451879/U$1 ( \12523 , \12521 , \12522 );
and \g453636/U$2 ( \12524 , \8404 , RIdf0ded0_1535);
and \g453636/U$3 ( \12525 , RIdf165d0_1631, \8351 );
nor \g453636/U$1 ( \12526 , \12524 , \12525 );
and \g454832/U$2 ( \12527 , \8313 , RIdeec2d0_1151);
and \g454832/U$3 ( \12528 , RIdeeefd0_1183, \8323 );
nor \g454832/U$1 ( \12529 , \12527 , \12528 );
not \g454831/U$1 ( \12530 , \12529 );
and \g449907/U$2 ( \12531 , \12530 , \8316 );
and \g449907/U$3 ( \12532 , RIdf0b1d0_1503, \8417 );
nor \g449907/U$1 ( \12533 , \12531 , \12532 );
nand \g448179/U$1 ( \12534 , \12520 , \12523 , \12526 , \12533 );
nor \g446005/U$1 ( \12535 , \12515 , \12516 , \12534 );
and \g451878/U$2 ( \12536 , \8378 , RIdf02ad0_1407);
and \g451878/U$3 ( \12537 , RIdefd0d0_1343, \8359 );
nor \g451878/U$1 ( \12538 , \12536 , \12537 );
and \g453723/U$2 ( \12539 , \8523 , RIdef76d0_1279);
and \g453723/U$3 ( \12540 , RIdefa3d0_1311, \8488 );
nor \g453723/U$1 ( \12541 , \12539 , \12540 );
and \g445154/U$2 ( \12542 , \12535 , \12538 , \12541 );
nor \g445154/U$1 ( \12543 , \12542 , \8477 );
and \g446006/U$2 ( \12544 , RIfc6efd8_6285, \8373 );
and \g446006/U$3 ( \12545 , RIfc6ee70_6284, \8330 );
and \g448886/U$2 ( \12546 , RIfeaaef8_8261, \8324 );
and \g448886/U$3 ( \12547 , \8531 , RIfc66a40_6190);
and \g448886/U$4 ( \12548 , RIfccde98_7365, \8488 );
nor \g448886/U$1 ( \12549 , \12546 , \12547 , \12548 );
and \g451886/U$2 ( \12550 , \8356 , RIfc668d8_6189);
and \g451886/U$3 ( \12551 , RIfc66608_6187, \8359 );
nor \g451886/U$1 ( \12552 , \12550 , \12551 );
and \g455092/U$2 ( \12553 , \8313 , RIdf25d50_1807);
and \g455092/U$3 ( \12554 , RIdf27ad8_1828, \8323 );
nor \g455092/U$1 ( \12555 , \12553 , \12554 );
not \g449909/U$3 ( \12556 , \12555 );
not \g449909/U$4 ( \12557 , \8376 );
and \g449909/U$2 ( \12558 , \12556 , \12557 );
and \g449909/U$5 ( \12559 , \8340 , RIfcacf40_6990);
nor \g449909/U$1 ( \12560 , \12558 , \12559 );
and \g451887/U$2 ( \12561 , \8378 , RIdf24130_1787);
and \g451887/U$3 ( \12562 , RIfe8b788_7931, \8417 );
nor \g451887/U$1 ( \12563 , \12561 , \12562 );
nand \g447662/U$1 ( \12564 , \12549 , \12552 , \12560 , \12563 );
nor \g446006/U$1 ( \12565 , \12544 , \12545 , \12564 );
and \g451884/U$2 ( \12566 , \8335 , RIdf18d30_1659);
and \g451884/U$3 ( \12567 , RIee2b750_4953, \8351 );
nor \g451884/U$1 ( \12568 , \12566 , \12567 );
and \g451885/U$2 ( \12569 , \8319 , RIfc6e8d0_6280);
and \g451885/U$3 ( \12570 , RIee27808_4908, \8404 );
nor \g451885/U$1 ( \12571 , \12569 , \12570 );
and \g445155/U$2 ( \12572 , \12565 , \12568 , \12571 );
nor \g445155/U$1 ( \12573 , \12572 , \8621 );
or \g444377/U$1 ( \12574 , \12452 , \12514 , \12543 , \12573 );
and \g446001/U$2 ( \12575 , RIfccb300_7334, \8373 );
and \g446001/U$3 ( \12576 , RIfc67c88_6203, \8383 );
and \g448882/U$2 ( \12577 , RIdee04f8_1016, \8414 );
and \g448882/U$3 ( \12578 , \8409 , RIfea8360_8230);
and \g448882/U$4 ( \12579 , RIded6a48_906, \8326 );
nor \g448882/U$1 ( \12580 , \12577 , \12578 , \12579 );
and \g451868/U$2 ( \12581 , \8356 , RIfc67df0_6204);
and \g451868/U$3 ( \12582 , RIfc6def8_6273, \8359 );
nor \g451868/U$1 ( \12583 , \12581 , \12582 );
and \g454548/U$2 ( \12584 , \8313 , RIfc67b20_6202);
and \g454548/U$3 ( \12585 , RIfcac130_6980, \8323 );
nor \g454548/U$1 ( \12586 , \12584 , \12585 );
not \g449903/U$3 ( \12587 , \12586 );
not \g449903/U$4 ( \12588 , \8347 );
and \g449903/U$2 ( \12589 , \12587 , \12588 );
and \g449903/U$5 ( \12590 , \8340 , RIded9040_933);
nor \g449903/U$1 ( \12591 , \12589 , \12590 );
and \g453986/U$2 ( \12592 , \8378 , RIdede338_992);
and \g453986/U$3 ( \12593 , RIfea81f8_8229, \8417 );
nor \g453986/U$1 ( \12594 , \12592 , \12593 );
nand \g447660/U$1 ( \12595 , \12580 , \12583 , \12591 , \12594 );
nor \g446001/U$1 ( \12596 , \12575 , \12576 , \12595 );
and \g451866/U$2 ( \12597 , \8335 , RIded26c8_858);
and \g451866/U$3 ( \12598 , RIfc6dc28_6271, \8351 );
nor \g451866/U$1 ( \12599 , \12597 , \12598 );
and \g451867/U$2 ( \12600 , \8319 , RIded4b58_884);
and \g451867/U$3 ( \12601 , RIfccd4c0_7358, \8404 );
nor \g451867/U$1 ( \12602 , \12600 , \12601 );
and \g445151/U$2 ( \12603 , \12596 , \12599 , \12602 );
nor \g445151/U$1 ( \12604 , \12603 , \8481 );
and \g446002/U$2 ( \12605 , RIe159600_2394, \8378 );
and \g446002/U$3 ( \12606 , RIe142e00_2138, \8359 );
and \g448883/U$2 ( \12607 , RIdedb638_960, \8319 );
and \g448883/U$3 ( \12608 , \8324 , RIdee68d0_1087);
and \g448883/U$4 ( \12609 , RIde95228_317, \8409 );
nor \g448883/U$1 ( \12610 , \12607 , \12608 , \12609 );
and \g451876/U$2 ( \12611 , \8335 , RIde7b170_190);
and \g451876/U$3 ( \12612 , RIdeffdd0_1375, \8340 );
nor \g451876/U$1 ( \12613 , \12611 , \12612 );
and \g451875/U$2 ( \12614 , \8404 , RIdec7700_733);
and \g451875/U$3 ( \12615 , RIdecfe00_829, \8351 );
nor \g451875/U$1 ( \12616 , \12614 , \12615 );
and \g454681/U$2 ( \12617 , \8313 , RIdeca400_765);
and \g454681/U$3 ( \12618 , RIdecd100_797, \8323 );
nor \g454681/U$1 ( \12619 , \12617 , \12618 );
not \g449905/U$3 ( \12620 , \12619 );
not \g449905/U$4 ( \12621 , \8328 );
and \g449905/U$2 ( \12622 , \12620 , \12621 );
and \g449905/U$5 ( \12623 , \8417 , RIdeb3c00_509);
nor \g449905/U$1 ( \12624 , \12622 , \12623 );
nand \g447661/U$1 ( \12625 , \12610 , \12613 , \12616 , \12624 );
nor \g446002/U$1 ( \12626 , \12605 , \12606 , \12625 );
and \g451873/U$2 ( \12627 , \8356 , RIdf1c6d8_1700);
and \g451873/U$3 ( \12628 , RIe16d808_2623, \8412 );
nor \g451873/U$1 ( \12629 , \12627 , \12628 );
and \g451872/U$2 ( \12630 , \8531 , RIdf2be58_1876);
and \g451872/U$3 ( \12631 , RIdf377f8_2008, \8488 );
nor \g451872/U$1 ( \12632 , \12630 , \12631 );
and \g445153/U$2 ( \12633 , \12626 , \12629 , \12632 );
nor \g445153/U$1 ( \12634 , \12633 , \8651 );
or \g444170/U$1 ( \12635 , \12574 , \12604 , \12634 );
_DC \g2a85/U$1 ( \12636 , \12635 , \8654 );
and \g448920/U$2 ( \12637 , RIe1695f0_2576, \8317 );
and \g448920/U$3 ( \12638 , \8326 , RIe16add8_2593);
and \g448920/U$4 ( \12639 , RIfe8aae0_7922, \8409 );
nor \g448920/U$1 ( \12640 , \12637 , \12638 , \12639 );
and \g451977/U$2 ( \12641 , \8335 , RIe167430_2552);
and \g451977/U$3 ( \12642 , RIee38fe0_5107, \8340 );
nor \g451977/U$1 ( \12643 , \12641 , \12642 );
and \g451520/U$2 ( \12644 , \8404 , RIfcaa240_6958);
and \g451520/U$3 ( \12645 , RIfcab320_6970, \8351 );
nor \g451520/U$1 ( \12646 , \12644 , \12645 );
and \g454427/U$2 ( \12647 , \8313 , RIfc6f6e0_6290);
and \g454427/U$3 ( \12648 , RIfca8350_6936, \8323 );
nor \g454427/U$1 ( \12649 , \12647 , \12648 );
not \g449935/U$3 ( \12650 , \12649 );
not \g449935/U$4 ( \12651 , \8328 );
and \g449935/U$2 ( \12652 , \12650 , \12651 );
and \g449935/U$5 ( \12653 , \8417 , RIde8fcd8_291);
nor \g449935/U$1 ( \12654 , \12652 , \12653 );
nand \g447680/U$1 ( \12655 , \12640 , \12643 , \12646 , \12654 );
and \g444684/U$2 ( \12656 , \12655 , \9700 );
and \g446033/U$2 ( \12657 , RIdec4898_700, \8351 );
and \g446033/U$3 ( \12658 , RIdebee98_636, \8404 );
and \g448922/U$2 ( \12659 , RIdea89e0_412, \8326 );
and \g448922/U$3 ( \12660 , \8523 , RIfcad648_6995);
and \g448922/U$4 ( \12661 , RIdeb0d98_476, \8486 );
nor \g448922/U$1 ( \12662 , \12659 , \12660 , \12661 );
and \g451986/U$2 ( \12663 , \8356 , RIdeae098_444);
and \g451986/U$3 ( \12664 , RIfc40d18_5763, \8359 );
nor \g451986/U$1 ( \12665 , \12663 , \12664 );
and \g455007/U$2 ( \12666 , \8313 , RIdeb9498_572);
and \g455007/U$3 ( \12667 , RIdebc198_604, \8323 );
nor \g455007/U$1 ( \12668 , \12666 , \12667 );
not \g449939/U$3 ( \12669 , \12668 );
not \g449939/U$4 ( \12670 , \8376 );
and \g449939/U$2 ( \12671 , \12669 , \12670 );
and \g449939/U$5 ( \12672 , \8340 , RIfcaa510_6960);
nor \g449939/U$1 ( \12673 , \12671 , \12672 );
and \g451985/U$2 ( \12674 , \8378 , RIdeb6798_540);
and \g451985/U$3 ( \12675 , RIfce6b28_7647, \8417 );
nor \g451985/U$1 ( \12676 , \12674 , \12675 );
nand \g447682/U$1 ( \12677 , \12662 , \12665 , \12673 , \12676 );
nor \g446033/U$1 ( \12678 , \12657 , \12658 , \12677 );
and \g451983/U$2 ( \12679 , \8335 , RIde9b7e0_348);
and \g451983/U$3 ( \12680 , RIdec1b98_668, \8383 );
nor \g451983/U$1 ( \12681 , \12679 , \12680 );
and \g451982/U$2 ( \12682 , \8319 , RIdea20e0_380);
and \g451982/U$3 ( \12683 , RIfc661d0_6184, \8371 );
nor \g451982/U$1 ( \12684 , \12682 , \12683 );
and \g445175/U$2 ( \12685 , \12678 , \12681 , \12684 );
nor \g445175/U$1 ( \12686 , \12685 , \8589 );
nor \g444684/U$1 ( \12687 , \12656 , \12686 );
and \g446815/U$2 ( \12688 , \12254 , RIde84860_236);
and \g446815/U$3 ( \12689 , RIde88d48_257, \12256 );
nor \g446815/U$1 ( \12690 , \12688 , \12689 );
and \g446814/U$2 ( \12691 , \12259 , RIfc64718_6165);
and \g446814/U$3 ( \12692 , RIde80a08_217, \12261 );
nor \g446814/U$1 ( \12693 , \12691 , \12692 );
and \g446816/U$2 ( \12694 , \12264 , RIfcadeb8_7001);
and \g446816/U$3 ( \12695 , RIfcae020_7002, \12266 );
nor \g446816/U$1 ( \12696 , \12694 , \12695 );
nand \g444486/U$1 ( \12697 , \12687 , \12690 , \12693 , \12696 );
and \g451996/U$2 ( \12698 , \8523 , RIfcab050_6968);
and \g451996/U$3 ( \12699 , RIe150d98_2297, \8488 );
nor \g451996/U$1 ( \12700 , \12698 , \12699 );
and \g446036/U$2 ( \12701 , RIe153a98_2329, \8378 );
and \g446036/U$3 ( \12702 , RIfc3f0f8_5743, \8359 );
and \g448927/U$2 ( \12703 , RIe15c198_2425, \8409 );
and \g448927/U$3 ( \12704 , \8373 , RIfe8a3d8_7917);
and \g448927/U$4 ( \12705 , RIe161b98_2489, \8383 );
nor \g448927/U$1 ( \12706 , \12703 , \12704 , \12705 );
and \g452000/U$2 ( \12707 , \8335 , RIe145998_2169);
and \g452000/U$3 ( \12708 , RIfcca658_7325, \8340 );
nor \g452000/U$1 ( \12709 , \12707 , \12708 );
and \g451042/U$2 ( \12710 , \8404 , RIe15ee98_2457);
and \g451042/U$3 ( \12711 , RIe164898_2521, \8351 );
nor \g451042/U$1 ( \12712 , \12710 , \12711 );
and \g454394/U$2 ( \12713 , \8313 , RIe148698_2201);
and \g454394/U$3 ( \12714 , RIe14b398_2233, \8323 );
nor \g454394/U$1 ( \12715 , \12713 , \12714 );
not \g454393/U$1 ( \12716 , \12715 );
and \g449943/U$2 ( \12717 , \12716 , \8316 );
and \g449943/U$3 ( \12718 , RIfe8a270_7916, \8417 );
nor \g449943/U$1 ( \12719 , \12717 , \12718 );
nand \g448184/U$1 ( \12720 , \12706 , \12709 , \12712 , \12719 );
nor \g446036/U$1 ( \12721 , \12701 , \12702 , \12720 );
and \g452351/U$2 ( \12722 , \8356 , RIe14e098_2265);
and \g452351/U$3 ( \12723 , RIe156798_2361, \8414 );
nor \g452351/U$1 ( \12724 , \12722 , \12723 );
nand \g445583/U$1 ( \12725 , \12700 , \12721 , \12724 );
and \g444852/U$2 ( \12726 , \12725 , \8369 );
and \g448924/U$2 ( \12727 , RIdf3c3e8_2062, \8414 );
and \g448924/U$3 ( \12728 , \8409 , RIfe8a540_7918);
and \g448924/U$4 ( \12729 , RIdf32c08_1954, \8324 );
nor \g448924/U$1 ( \12730 , \12727 , \12728 , \12729 );
and \g451992/U$2 ( \12731 , \8356 , RIee2d0a0_4971);
and \g451992/U$3 ( \12732 , RIfc6b1f8_6241, \8359 );
nor \g451992/U$1 ( \12733 , \12731 , \12732 );
and \g454475/U$2 ( \12734 , \8313 , RIfc70d60_6306);
and \g454475/U$3 ( \12735 , RIee2f260_4995, \8323 );
nor \g454475/U$1 ( \12736 , \12734 , \12735 );
not \g449940/U$3 ( \12737 , \12736 );
not \g449940/U$4 ( \12738 , \8347 );
and \g449940/U$2 ( \12739 , \12737 , \12738 );
and \g449940/U$5 ( \12740 , \8340 , RIfe8a978_7921);
nor \g449940/U$1 ( \12741 , \12739 , \12740 );
and \g451991/U$2 ( \12742 , \8378 , RIdf3a0c0_2037);
and \g451991/U$3 ( \12743 , RIe140808_2111, \8417 );
nor \g451991/U$1 ( \12744 , \12742 , \12743 );
nand \g447683/U$1 ( \12745 , \12730 , \12733 , \12741 , \12744 );
and \g444852/U$3 ( \12746 , \9266 , \12745 );
nor \g444852/U$1 ( \12747 , \12726 , \12746 );
and \g446818/U$2 ( \12748 , \9288 , RIee30e80_5015);
and \g446818/U$3 ( \12749 , RIee31b28_5024, \9290 );
nor \g446818/U$1 ( \12750 , \12748 , \12749 );
and \g446817/U$2 ( \12751 , \9293 , RIfe8a6a8_7919);
and \g446817/U$3 ( \12752 , RIfe8a810_7920, \9296 );
nor \g446817/U$1 ( \12753 , \12751 , \12752 );
and \g446819/U$2 ( \12754 , \9299 , RIdf2e9f0_1907);
and \g446819/U$3 ( \12755 , RIdf308e0_1929, \9301 );
nor \g446819/U$1 ( \12756 , \12754 , \12755 );
nand \g444603/U$1 ( \12757 , \12747 , \12750 , \12753 , \12756 );
and \g446027/U$2 ( \12758 , RIdf23fc8_1786, \8378 );
and \g446027/U$3 ( \12759 , RIfc6aaf0_6236, \8359 );
and \g448916/U$2 ( \12760 , RIdf27970_1827, \8409 );
and \g448916/U$3 ( \12761 , \8373 , RIee28a50_4921);
and \g448916/U$4 ( \12762 , RIee29e00_4935, \8383 );
nor \g448916/U$1 ( \12763 , \12760 , \12761 , \12762 );
and \g451965/U$2 ( \12764 , \8335 , RIfeaa7f0_8256);
and \g451965/U$3 ( \12765 , RIdf21160_1753, \8340 );
nor \g451965/U$1 ( \12766 , \12764 , \12765 );
and \g450990/U$2 ( \12767 , \8404 , RIee276a0_4907);
and \g450990/U$3 ( \12768 , RIee2b5e8_4952, \8351 );
nor \g450990/U$1 ( \12769 , \12767 , \12768 );
and \g454308/U$2 ( \12770 , \8313 , RIdf1ac20_1681);
and \g454308/U$3 ( \12771 , RIdf1f108_1730, \8323 );
nor \g454308/U$1 ( \12772 , \12770 , \12771 );
not \g454307/U$1 ( \12773 , \12772 );
and \g449933/U$2 ( \12774 , \12773 , \8316 );
and \g449933/U$3 ( \12775 , RIdf29c98_1852, \8417 );
nor \g449933/U$1 ( \12776 , \12774 , \12775 );
nand \g448182/U$1 ( \12777 , \12763 , \12766 , \12769 , \12776 );
nor \g446027/U$1 ( \12778 , \12758 , \12759 , \12777 );
and \g451962/U$2 ( \12779 , \8356 , RIfcdd4b0_7540);
and \g451962/U$3 ( \12780 , RIdf25be8_1806, \8414 );
nor \g451962/U$1 ( \12781 , \12779 , \12780 );
and \g451961/U$2 ( \12782 , \8531 , RIdf22678_1768);
and \g451961/U$3 ( \12783 , RIfc6ac58_6237, \8488 );
nor \g451961/U$1 ( \12784 , \12782 , \12783 );
and \g445172/U$2 ( \12785 , \12778 , \12781 , \12784 );
nor \g445172/U$1 ( \12786 , \12785 , \8621 );
and \g446030/U$2 ( \12787 , RIdecfc98_828, \8351 );
and \g446030/U$3 ( \12788 , RIde7ae28_189, \8335 );
and \g448919/U$2 ( \12789 , RIe16d6a0_2622, \8414 );
and \g448919/U$3 ( \12790 , \8409 , RIde94ee0_316);
and \g448919/U$4 ( \12791 , RIdee6768_1086, \8326 );
nor \g448919/U$1 ( \12792 , \12789 , \12790 , \12791 );
and \g451971/U$2 ( \12793 , \8356 , RIdf1c570_1699);
and \g451971/U$3 ( \12794 , RIe142c98_2137, \8359 );
nor \g451971/U$1 ( \12795 , \12793 , \12794 );
and \g454195/U$2 ( \12796 , \8313 , RIdf2bcf0_1875);
and \g454195/U$3 ( \12797 , RIdf37690_2007, \8323 );
nor \g454195/U$1 ( \12798 , \12796 , \12797 );
not \g449555/U$3 ( \12799 , \12798 );
not \g449555/U$4 ( \12800 , \8347 );
and \g449555/U$2 ( \12801 , \12799 , \12800 );
and \g449555/U$5 ( \12802 , \8340 , RIdeffc68_1374);
nor \g449555/U$1 ( \12803 , \12801 , \12802 );
and \g451970/U$2 ( \12804 , \8378 , RIe159498_2393);
and \g451970/U$3 ( \12805 , RIdeb3a98_508, \8417 );
nor \g451970/U$1 ( \12806 , \12804 , \12805 );
nand \g447679/U$1 ( \12807 , \12792 , \12795 , \12803 , \12806 );
nor \g446030/U$1 ( \12808 , \12787 , \12788 , \12807 );
and \g451969/U$2 ( \12809 , \8319 , RIdedb4d0_959);
and \g451969/U$3 ( \12810 , RIdec7598_732, \8404 );
nor \g451969/U$1 ( \12811 , \12809 , \12810 );
and \g451968/U$2 ( \12812 , \8373 , RIdeca298_764);
and \g451968/U$3 ( \12813 , RIdeccf98_796, \8383 );
nor \g451968/U$1 ( \12814 , \12812 , \12813 );
and \g445173/U$2 ( \12815 , \12808 , \12811 , \12814 );
nor \g445173/U$1 ( \12816 , \12815 , \8651 );
or \g444333/U$1 ( \12817 , \12697 , \12757 , \12786 , \12816 );
and \g446023/U$2 ( \12818 , RIdf10a68_1566, \8373 );
and \g446023/U$3 ( \12819 , RIdf13768_1598, \8330 );
and \g448911/U$2 ( \12820 , RIdf05668_1438, \8414 );
and \g448911/U$3 ( \12821 , \8409 , RIdf08368_1470);
and \g448911/U$4 ( \12822 , RIdeeee68_1182, \8326 );
nor \g448911/U$1 ( \12823 , \12820 , \12821 , \12822 );
and \g451949/U$2 ( \12824 , \8356 , RIdef4868_1246);
and \g451949/U$3 ( \12825 , RIdefcf68_1342, \8359 );
nor \g451949/U$1 ( \12826 , \12824 , \12825 );
and \g454510/U$2 ( \12827 , \8313 , RIdef7568_1278);
and \g454510/U$3 ( \12828 , RIdefa268_1310, \8323 );
nor \g454510/U$1 ( \12829 , \12827 , \12828 );
not \g449930/U$3 ( \12830 , \12829 );
not \g449930/U$4 ( \12831 , \8347 );
and \g449930/U$2 ( \12832 , \12830 , \12831 );
and \g449930/U$5 ( \12833 , \8340 , RIdef1b68_1214);
nor \g449930/U$1 ( \12834 , \12832 , \12833 );
and \g451446/U$2 ( \12835 , \8378 , RIdf02968_1406);
and \g451446/U$3 ( \12836 , RIdf0b068_1502, \8417 );
nor \g451446/U$1 ( \12837 , \12835 , \12836 );
nand \g447674/U$1 ( \12838 , \12823 , \12826 , \12834 , \12837 );
nor \g446023/U$1 ( \12839 , \12818 , \12819 , \12838 );
and \g451527/U$2 ( \12840 , \8335 , RIdee9468_1118);
and \g451527/U$3 ( \12841 , RIdf16468_1630, \8351 );
nor \g451527/U$1 ( \12842 , \12840 , \12841 );
and \g451947/U$2 ( \12843 , \8319 , RIdeec168_1150);
and \g451947/U$3 ( \12844 , RIdf0dd68_1534, \8404 );
nor \g451947/U$1 ( \12845 , \12843 , \12844 );
and \g445167/U$2 ( \12846 , \12839 , \12842 , \12845 );
nor \g445167/U$1 ( \12847 , \12846 , \8477 );
and \g446026/U$2 ( \12848 , RIfe8ac48_7923, \8414 );
and \g446026/U$3 ( \12849 , RIee20ff8_4834, \8356 );
and \g448914/U$2 ( \12850 , RIded49f0_883, \8317 );
and \g448914/U$3 ( \12851 , \8326 , RIfe8af18_7925);
and \g448914/U$4 ( \12852 , RIdee23e8_1038, \8407 );
nor \g448914/U$1 ( \12853 , \12850 , \12851 , \12852 );
and \g451958/U$2 ( \12854 , \8335 , RIfe8b080_7926);
and \g451958/U$3 ( \12855 , RIded8ed8_932, \8340 );
nor \g451958/U$1 ( \12856 , \12854 , \12855 );
and \g451957/U$2 ( \12857 , \8404 , RIee23050_4857);
and \g451957/U$3 ( \12858 , RIee25378_4882, \8351 );
nor \g451957/U$1 ( \12859 , \12857 , \12858 );
and \g454565/U$2 ( \12860 , \8313 , RIee23a28_4864);
and \g454565/U$3 ( \12861 , RIee24568_4872, \8323 );
nor \g454565/U$1 ( \12862 , \12860 , \12861 );
not \g449692/U$3 ( \12863 , \12862 );
not \g449692/U$4 ( \12864 , \8328 );
and \g449692/U$2 ( \12865 , \12863 , \12864 );
and \g449692/U$5 ( \12866 , \8417 , RIfe8adb0_7924);
nor \g449692/U$1 ( \12867 , \12865 , \12866 );
nand \g447676/U$1 ( \12868 , \12853 , \12856 , \12859 , \12867 );
nor \g446026/U$1 ( \12869 , \12848 , \12849 , \12868 );
and \g451956/U$2 ( \12870 , \8378 , RIdede1d0_991);
and \g451956/U$3 ( \12871 , RIfca5650_6904, \8359 );
nor \g451956/U$1 ( \12872 , \12870 , \12871 );
and \g451955/U$2 ( \12873 , \8523 , RIfceeb20_7738);
and \g451955/U$3 ( \12874 , RIee220d8_4846, \8488 );
nor \g451955/U$1 ( \12875 , \12873 , \12874 );
and \g445169/U$2 ( \12876 , \12869 , \12872 , \12875 );
nor \g445169/U$1 ( \12877 , \12876 , \8481 );
or \g444199/U$1 ( \12878 , \12817 , \12847 , \12877 );
_DC \g2b0a/U$1 ( \12879 , \12878 , \8654 );
and \g451462/U$2 ( \12880 , \8371 , RIdf10900_1565);
and \g451462/U$3 ( \12881 , RIdf13600_1597, \8383 );
nor \g451462/U$1 ( \12882 , \12880 , \12881 );
and \g445903/U$2 ( \12883 , RIdf16300_1629, \8351 );
and \g445903/U$3 ( \12884 , RIdee9300_1117, \8335 );
and \g448754/U$2 ( \12885 , RIdeeed00_1181, \8326 );
and \g448754/U$3 ( \12886 , \8531 , RIdef7400_1277);
and \g448754/U$4 ( \12887 , RIdefa100_1309, \8488 );
nor \g448754/U$1 ( \12888 , \12885 , \12886 , \12887 );
and \g451466/U$2 ( \12889 , \8356 , RIdef4700_1245);
and \g451466/U$3 ( \12890 , RIdefce00_1341, \8359 );
nor \g451466/U$1 ( \12891 , \12889 , \12890 );
and \g454533/U$2 ( \12892 , \8313 , RIdf05500_1437);
and \g454533/U$3 ( \12893 , RIdf08200_1469, \8323 );
nor \g454533/U$1 ( \12894 , \12892 , \12893 );
not \g449783/U$3 ( \12895 , \12894 );
not \g449783/U$4 ( \12896 , \8376 );
and \g449783/U$2 ( \12897 , \12895 , \12896 );
and \g449783/U$5 ( \12898 , \8340 , RIdef1a00_1213);
nor \g449783/U$1 ( \12899 , \12897 , \12898 );
and \g451465/U$2 ( \12900 , \8378 , RIdf02800_1405);
and \g451465/U$3 ( \12901 , RIdf0af00_1501, \8417 );
nor \g451465/U$1 ( \12902 , \12900 , \12901 );
nand \g447596/U$1 ( \12903 , \12888 , \12891 , \12899 , \12902 );
nor \g445903/U$1 ( \12904 , \12883 , \12884 , \12903 );
and \g451464/U$2 ( \12905 , \8319 , RIdeec000_1149);
and \g451464/U$3 ( \12906 , RIdf0dc00_1533, \8404 );
nor \g451464/U$1 ( \12907 , \12905 , \12906 );
nand \g445552/U$1 ( \12908 , \12882 , \12904 , \12907 );
and \g444765/U$2 ( \12909 , \12908 , \8478 );
and \g448750/U$2 ( \12910 , RIdf25a80_1805, \8414 );
and \g448750/U$3 ( \12911 , \8407 , RIdf27808_1826);
and \g448750/U$4 ( \12912 , RIdf1efa0_1729, \8326 );
nor \g448750/U$1 ( \12913 , \12910 , \12911 , \12912 );
and \g451459/U$2 ( \12914 , \8356 , RIfc54cc8_5987);
and \g451459/U$3 ( \12915 , RIfc55100_5990, \8359 );
nor \g451459/U$1 ( \12916 , \12914 , \12915 );
and \g454261/U$2 ( \12917 , \8313 , RIfc54f98_5989);
and \g454261/U$3 ( \12918 , RIfcd9f40_7502, \8323 );
nor \g454261/U$1 ( \12919 , \12917 , \12918 );
not \g449781/U$3 ( \12920 , \12919 );
not \g449781/U$4 ( \12921 , \8347 );
and \g449781/U$2 ( \12922 , \12920 , \12921 );
and \g449781/U$5 ( \12923 , \8340 , RIfc4b218_5877);
nor \g449781/U$1 ( \12924 , \12922 , \12923 );
and \g451457/U$2 ( \12925 , \8378 , RIdf23e60_1785);
and \g451457/U$3 ( \12926 , RIdf29b30_1851, \8417 );
nor \g451457/U$1 ( \12927 , \12925 , \12926 );
nand \g447595/U$1 ( \12928 , \12913 , \12916 , \12924 , \12927 );
and \g444765/U$3 ( \12929 , \8752 , \12928 );
nor \g444765/U$1 ( \12930 , \12909 , \12929 );
and \g446687/U$2 ( \12931 , \11762 , RIdf18bc8_1658);
and \g446687/U$3 ( \12932 , RIfcc69e0_7282, \11764 );
nor \g446687/U$1 ( \12933 , \12931 , \12932 );
and \g446686/U$2 ( \12934 , \11767 , RIfec23a0_8330);
and \g446686/U$3 ( \12935 , RIee2b480_4951, \11769 );
nor \g446686/U$1 ( \12936 , \12934 , \12935 );
and \g446688/U$2 ( \12937 , \11511 , RIfec2238_8329);
and \g446688/U$3 ( \12938 , RIee288e8_4920, \11513 );
nor \g446688/U$1 ( \12939 , \12937 , \12938 );
nand \g444472/U$1 ( \12940 , \12930 , \12933 , \12936 , \12939 );
and \g451474/U$2 ( \12941 , \8317 , RIe148530_2200);
and \g451474/U$3 ( \12942 , RIe15ed30_2456, \8404 );
nor \g451474/U$1 ( \12943 , \12941 , \12942 );
and \g445907/U$2 ( \12944 , RIee36cb8_5082, \8373 );
and \g445907/U$3 ( \12945 , RIe161a30_2488, \8330 );
and \g448759/U$2 ( \12946 , RIe14b230_2232, \8324 );
and \g448759/U$3 ( \12947 , \8531 , RIfc8af08_6603);
and \g448759/U$4 ( \12948 , RIe150c30_2296, \8488 );
nor \g448759/U$1 ( \12949 , \12946 , \12947 , \12948 );
and \g451477/U$2 ( \12950 , \8356 , RIe14df30_2264);
and \g451477/U$3 ( \12951 , RIfcc7688_7291, \8359 );
nor \g451477/U$1 ( \12952 , \12950 , \12951 );
and \g455228/U$2 ( \12953 , \8313 , RIe156630_2360);
and \g455228/U$3 ( \12954 , RIe15c030_2424, \8323 );
nor \g455228/U$1 ( \12955 , \12953 , \12954 );
not \g449787/U$3 ( \12956 , \12955 );
not \g449787/U$4 ( \12957 , \8376 );
and \g449787/U$2 ( \12958 , \12956 , \12957 );
and \g449787/U$5 ( \12959 , \8340 , RIfc9a250_6776);
nor \g449787/U$1 ( \12960 , \12958 , \12959 );
and \g451476/U$2 ( \12961 , \8378 , RIe153930_2328);
and \g451476/U$3 ( \12962 , RIfcc7250_7288, \8417 );
nor \g451476/U$1 ( \12963 , \12961 , \12962 );
nand \g447600/U$1 ( \12964 , \12949 , \12952 , \12960 , \12963 );
nor \g445907/U$1 ( \12965 , \12944 , \12945 , \12964 );
and \g451472/U$2 ( \12966 , \8335 , RIe145830_2168);
and \g451472/U$3 ( \12967 , RIe164730_2520, \8351 );
nor \g451472/U$1 ( \12968 , \12966 , \12967 );
nand \g445553/U$1 ( \12969 , \12943 , \12965 , \12968 );
and \g444850/U$2 ( \12970 , \12969 , \8369 );
and \g448757/U$2 ( \12971 , RIfec2940_8334, \8324 );
and \g448757/U$3 ( \12972 , \8531 , RIfcdb458_7517);
and \g448757/U$4 ( \12973 , RIee2f0f8_4994, \8488 );
nor \g448757/U$1 ( \12974 , \12971 , \12972 , \12973 );
and \g451471/U$2 ( \12975 , \8356 , RIee2cf38_4970);
and \g451471/U$3 ( \12976 , RIfc9a958_6781, \8359 );
nor \g451471/U$1 ( \12977 , \12975 , \12976 );
and \g454538/U$2 ( \12978 , \8313 , RIdf3c280_2061);
and \g454538/U$3 ( \12979 , RIdf3e440_2085, \8323 );
nor \g454538/U$1 ( \12980 , \12978 , \12979 );
not \g449786/U$3 ( \12981 , \12980 );
not \g449786/U$4 ( \12982 , \8376 );
and \g449786/U$2 ( \12983 , \12981 , \12982 );
and \g449786/U$5 ( \12984 , \8340 , RIdf34c60_1977);
nor \g449786/U$1 ( \12985 , \12983 , \12984 );
and \g453735/U$2 ( \12986 , \8378 , RIdf39f58_2036);
and \g453735/U$3 ( \12987 , RIe1406a0_2110, \8417 );
nor \g453735/U$1 ( \12988 , \12986 , \12987 );
nand \g447598/U$1 ( \12989 , \12974 , \12977 , \12985 , \12988 );
and \g444850/U$3 ( \12990 , \9266 , \12989 );
nor \g444850/U$1 ( \12991 , \12970 , \12990 );
and \g446693/U$2 ( \12992 , \9288 , RIfcec960_7714);
and \g446693/U$3 ( \12993 , RIfca1ca8_6863, \9290 );
nor \g446693/U$1 ( \12994 , \12992 , \12993 );
and \g446692/U$2 ( \12995 , \9293 , RIfc56bb8_6009);
and \g446692/U$3 ( \12996 , RIfc9aac0_6782, \9296 );
nor \g446692/U$1 ( \12997 , \12995 , \12996 );
and \g446694/U$2 ( \12998 , \9299 , RIdf2e888_1906);
and \g446694/U$3 ( \12999 , RIdf30778_1928, \9301 );
nor \g446694/U$1 ( \13000 , \12998 , \12999 );
nand \g444579/U$1 ( \13001 , \12991 , \12994 , \12997 , \13000 );
and \g445898/U$2 ( \13002 , RIdee0390_1015, \8414 );
and \g445898/U$3 ( \13003 , RIfca0790_6848, \8531 );
and \g448745/U$2 ( \13004 , RIdee2280_1037, \8407 );
and \g448745/U$3 ( \13005 , \8373 , RIfcc46b8_7257);
and \g448745/U$4 ( \13006 , RIfc9e8a0_6826, \8330 );
nor \g448745/U$1 ( \13007 , \13004 , \13005 , \13006 );
and \g451444/U$2 ( \13008 , \8335 , RIded2560_857);
and \g451444/U$3 ( \13009 , RIded8d70_931, \8340 );
nor \g451444/U$1 ( \13010 , \13008 , \13009 );
and \g453085/U$2 ( \13011 , \8404 , RIfcd4108_7435);
and \g453085/U$3 ( \13012 , RIfce4ad0_7624, \8351 );
nor \g453085/U$1 ( \13013 , \13011 , \13012 );
and \g455284/U$2 ( \13014 , \8313 , RIded4888_882);
and \g455284/U$3 ( \13015 , RIded68e0_905, \8323 );
nor \g455284/U$1 ( \13016 , \13014 , \13015 );
not \g455283/U$1 ( \13017 , \13016 );
and \g449775/U$2 ( \13018 , \13017 , \8316 );
and \g449775/U$3 ( \13019 , RIdee4440_1061, \8417 );
nor \g449775/U$1 ( \13020 , \13018 , \13019 );
nand \g448160/U$1 ( \13021 , \13007 , \13010 , \13013 , \13020 );
nor \g445898/U$1 ( \13022 , \13002 , \13003 , \13021 );
and \g451439/U$2 ( \13023 , \8356 , RIfc50ee8_5943);
and \g451439/U$3 ( \13024 , RIfcda0a8_7503, \8359 );
nor \g451439/U$1 ( \13025 , \13023 , \13024 );
and \g451441/U$2 ( \13026 , \8378 , RIdede068_990);
and \g451441/U$3 ( \13027 , RIfce54a8_7631, \8488 );
nor \g451441/U$1 ( \13028 , \13026 , \13027 );
and \g445074/U$2 ( \13029 , \13022 , \13025 , \13028 );
nor \g445074/U$1 ( \13030 , \13029 , \8481 );
and \g445901/U$2 ( \13031 , RIe16d538_2621, \8414 );
and \g445901/U$3 ( \13032 , RIdf2bb88_1874, \8531 );
and \g448747/U$2 ( \13033 , RIdedb368_958, \8319 );
and \g448747/U$3 ( \13034 , \8326 , RIdee6600_1085);
and \g448747/U$4 ( \13035 , RIde94b98_315, \8409 );
nor \g448747/U$1 ( \13036 , \13033 , \13034 , \13035 );
and \g451452/U$2 ( \13037 , \8335 , RIde7aae0_188);
and \g451452/U$3 ( \13038 , RIdeffb00_1373, \8340 );
nor \g451452/U$1 ( \13039 , \13037 , \13038 );
and \g452164/U$2 ( \13040 , \8404 , RIdec7430_731);
and \g452164/U$3 ( \13041 , RIdecfb30_827, \8351 );
nor \g452164/U$1 ( \13042 , \13040 , \13041 );
and \g454707/U$2 ( \13043 , \8313 , RIdeca130_763);
and \g454707/U$3 ( \13044 , RIdecce30_795, \8323 );
nor \g454707/U$1 ( \13045 , \13043 , \13044 );
not \g449777/U$3 ( \13046 , \13045 );
not \g449777/U$4 ( \13047 , \8328 );
and \g449777/U$2 ( \13048 , \13046 , \13047 );
and \g449777/U$5 ( \13049 , \8417 , RIdeb3930_507);
nor \g449777/U$1 ( \13050 , \13048 , \13049 );
nand \g447593/U$1 ( \13051 , \13036 , \13039 , \13042 , \13050 );
nor \g445901/U$1 ( \13052 , \13031 , \13032 , \13051 );
and \g451447/U$2 ( \13053 , \8356 , RIdf1c408_1698);
and \g451447/U$3 ( \13054 , RIe142b30_2136, \8359 );
nor \g451447/U$1 ( \13055 , \13053 , \13054 );
and \g451449/U$2 ( \13056 , \8378 , RIe159330_2392);
and \g451449/U$3 ( \13057 , RIdf37528_2006, \8488 );
nor \g451449/U$1 ( \13058 , \13056 , \13057 );
and \g445076/U$2 ( \13059 , \13052 , \13055 , \13058 );
nor \g445076/U$1 ( \13060 , \13059 , \8651 );
or \g444322/U$1 ( \13061 , \12940 , \13001 , \13030 , \13060 );
and \g445894/U$2 ( \13062 , RIfce3f90_7616, \8371 );
and \g445894/U$3 ( \13063 , RIdec1a30_667, \8330 );
and \g448740/U$2 ( \13064 , RIdea8698_411, \8326 );
and \g448740/U$3 ( \13065 , \8531 , RIfc5a998_6053);
and \g448740/U$4 ( \13066 , RIdeb0c30_475, \8488 );
nor \g448740/U$1 ( \13067 , \13064 , \13065 , \13066 );
and \g451424/U$2 ( \13068 , \8356 , RIdeadf30_443);
and \g451424/U$3 ( \13069 , RIfc8c588_6619, \8359 );
nor \g451424/U$1 ( \13070 , \13068 , \13069 );
and \g454804/U$2 ( \13071 , \8313 , RIdeb9330_571);
and \g454804/U$3 ( \13072 , RIdebc030_603, \8323 );
nor \g454804/U$1 ( \13073 , \13071 , \13072 );
not \g449770/U$3 ( \13074 , \13073 );
not \g449770/U$4 ( \13075 , \8376 );
and \g449770/U$2 ( \13076 , \13074 , \13075 );
and \g449770/U$5 ( \13077 , \8340 , RIfc99b48_6771);
nor \g449770/U$1 ( \13078 , \13076 , \13077 );
and \g451422/U$2 ( \13079 , \8378 , RIdeb6630_539);
and \g451422/U$3 ( \13080 , RIfcc3308_7243, \8417 );
nor \g451422/U$1 ( \13081 , \13079 , \13080 );
nand \g447589/U$1 ( \13082 , \13067 , \13070 , \13078 , \13081 );
nor \g445894/U$1 ( \13083 , \13062 , \13063 , \13082 );
and \g451417/U$2 ( \13084 , \8335 , RIde9b498_347);
and \g451417/U$3 ( \13085 , RIdec4730_699, \8351 );
nor \g451417/U$1 ( \13086 , \13084 , \13085 );
and \g451418/U$2 ( \13087 , \8319 , RIdea1d98_379);
and \g451418/U$3 ( \13088 , RIdebed30_635, \8404 );
nor \g451418/U$1 ( \13089 , \13087 , \13088 );
and \g445069/U$2 ( \13090 , \13083 , \13086 , \13089 );
nor \g445069/U$1 ( \13091 , \13090 , \8589 );
and \g445896/U$2 ( \13092 , RIde88a00_256, \8414 );
and \g445896/U$3 ( \13093 , RIfca3058_6877, \8356 );
and \g448742/U$2 ( \13094 , RIfca3328_6879, \8319 );
and \g448742/U$3 ( \13095 , \8326 , RIfec27d8_8333);
and \g448742/U$4 ( \13096 , RIfec2508_8331, \8409 );
nor \g448742/U$1 ( \13097 , \13094 , \13095 , \13096 );
and \g451433/U$2 ( \13098 , \8335 , RIe1672c8_2551);
and \g451433/U$3 ( \13099 , RIee38e78_5106, \8340 );
nor \g451433/U$1 ( \13100 , \13098 , \13099 );
and \g451432/U$2 ( \13101 , \8404 , RIfca3fd0_6888);
and \g451432/U$3 ( \13102 , RIfc78bf0_6396, \8351 );
nor \g451432/U$1 ( \13103 , \13101 , \13102 );
and \g454988/U$2 ( \13104 , \8313 , RIfca12d0_6856);
and \g454988/U$3 ( \13105 , RIfcbc558_7165, \8323 );
nor \g454988/U$1 ( \13106 , \13104 , \13105 );
not \g449773/U$3 ( \13107 , \13106 );
not \g449773/U$4 ( \13108 , \8328 );
and \g449773/U$2 ( \13109 , \13107 , \13108 );
and \g449773/U$5 ( \13110 , \8417 , RIfec2670_8332);
nor \g449773/U$1 ( \13111 , \13109 , \13110 );
nand \g447591/U$1 ( \13112 , \13097 , \13100 , \13103 , \13111 );
nor \g445896/U$1 ( \13113 , \13092 , \13093 , \13112 );
and \g451430/U$2 ( \13114 , \8378 , RIde84518_235);
and \g451430/U$3 ( \13115 , RIfcc35d8_7245, \8359 );
nor \g451430/U$1 ( \13116 , \13114 , \13115 );
and \g450696/U$2 ( \13117 , \8531 , RIfc5a290_6048);
and \g450696/U$3 ( \13118 , RIfcb57a8_7087, \8488 );
nor \g450696/U$1 ( \13119 , \13117 , \13118 );
and \g445071/U$2 ( \13120 , \13113 , \13116 , \13119 );
nor \g445071/U$1 ( \13121 , \13120 , \8558 );
or \g444271/U$1 ( \13122 , \13061 , \13091 , \13121 );
_DC \g2b8f/U$1 ( \13123 , \13122 , \8654 );
and \g451583/U$2 ( \13124 , \8324 , RIe16ac70_2592);
and \g451583/U$3 ( \13125 , RIfcb8778_7121, \8404 );
nor \g451583/U$1 ( \13126 , \13124 , \13125 );
and \g445931/U$2 ( \13127 , RIfce13f8_7585, \8371 );
and \g445931/U$3 ( \13128 , RIfc850d0_6536, \8319 );
and \g448790/U$2 ( \13129 , RIfce1128_7583, \8531 );
and \g448790/U$3 ( \13130 , \8486 , RIfcb8070_7116);
and \g448790/U$4 ( \13131 , RIfc9c9b0_6804, \8330 );
nor \g448790/U$1 ( \13132 , \13129 , \13130 , \13131 );
and \g451588/U$2 ( \13133 , \8356 , RIfc9c140_6798);
and \g451588/U$3 ( \13134 , RIde806c0_216, \8359 );
nor \g451588/U$1 ( \13135 , \13133 , \13134 );
and \g454596/U$2 ( \13136 , \8313 , RIde886b8_255);
and \g454596/U$3 ( \13137 , RIfe8d3a8_7951, \8323 );
nor \g454596/U$1 ( \13138 , \13136 , \13137 );
not \g449819/U$3 ( \13139 , \13138 );
not \g449819/U$4 ( \13140 , \8376 );
and \g449819/U$2 ( \13141 , \13139 , \13140 );
and \g449819/U$5 ( \13142 , \8351 , RIfc85ee0_6546);
nor \g449819/U$1 ( \13143 , \13141 , \13142 );
and \g450638/U$2 ( \13144 , \8378 , RIde841d0_234);
and \g450638/U$3 ( \13145 , RIfe8d510_7952, \8417 );
nor \g450638/U$1 ( \13146 , \13144 , \13145 );
nand \g447620/U$1 ( \13147 , \13132 , \13135 , \13143 , \13146 );
nor \g445931/U$1 ( \13148 , \13127 , \13128 , \13147 );
and \g451585/U$2 ( \13149 , \8335 , RIe167160_2550);
and \g451585/U$3 ( \13150 , RIee38d10_5105, \8340 );
nor \g451585/U$1 ( \13151 , \13149 , \13150 );
nand \g445560/U$1 ( \13152 , \13126 , \13148 , \13151 );
and \g444694/U$2 ( \13153 , \13152 , \9700 );
and \g448787/U$2 ( \13154 , RIdeb91c8_570, \8412 );
and \g448787/U$3 ( \13155 , \8407 , RIdebbec8_602);
and \g448787/U$4 ( \13156 , RIdec18c8_666, \8383 );
nor \g448787/U$1 ( \13157 , \13154 , \13155 , \13156 );
and \g451580/U$2 ( \13158 , \8356 , RIdeaddc8_442);
and \g451580/U$3 ( \13159 , RIfc85d78_6545, \8359 );
nor \g451580/U$1 ( \13160 , \13158 , \13159 );
and \g455115/U$2 ( \13161 , \8313 , RIfc85aa8_6543);
and \g455115/U$3 ( \13162 , RIdeb0ac8_474, \8323 );
nor \g455115/U$1 ( \13163 , \13161 , \13162 );
not \g449817/U$3 ( \13164 , \13163 );
not \g449817/U$4 ( \13165 , \8347 );
and \g449817/U$2 ( \13166 , \13164 , \13165 );
and \g449817/U$5 ( \13167 , \8351 , RIdec45c8_698);
nor \g449817/U$1 ( \13168 , \13166 , \13167 );
and \g451579/U$2 ( \13169 , \8378 , RIdeb64c8_538);
and \g451579/U$3 ( \13170 , RIfcb8bb0_7124, \8417 );
nor \g451579/U$1 ( \13171 , \13169 , \13170 );
nand \g447618/U$1 ( \13172 , \13157 , \13160 , \13168 , \13171 );
and \g444694/U$3 ( \13173 , \9702 , \13172 );
nor \g444694/U$1 ( \13174 , \13153 , \13173 );
and \g446720/U$2 ( \13175 , \9724 , RIdebebc8_634);
and \g446720/U$3 ( \13176 , RIfce85e0_7666, \9726 );
nor \g446720/U$1 ( \13177 , \13175 , \13176 );
and \g446719/U$2 ( \13178 , \9729 , RIde9b150_346);
and \g446719/U$3 ( \13179 , RIdea1a50_378, \9731 );
nor \g446719/U$1 ( \13180 , \13178 , \13179 );
and \g446718/U$2 ( \13181 , \9734 , RIdea8350_410);
and \g446718/U$3 ( \13182 , RIfc4d3d8_5901, \9736 );
nor \g446718/U$1 ( \13183 , \13181 , \13182 );
nand \g444475/U$1 ( \13184 , \13174 , \13177 , \13180 , \13183 );
and \g451599/U$2 ( \13185 , \8531 , RIfcb6cc0_7102);
and \g451599/U$3 ( \13186 , RIfe8cb38_7945, \8414 );
nor \g451599/U$1 ( \13187 , \13185 , \13186 );
and \g445934/U$2 ( \13188 , RIdee2118_1036, \8409 );
and \g445934/U$3 ( \13189 , RIdeddf00_989, \8378 );
and \g448796/U$2 ( \13190 , RIded4720_881, \8317 );
and \g448796/U$3 ( \13191 , \8326 , RIded6778_904);
and \g448796/U$4 ( \13192 , RIee21f70_4845, \8488 );
nor \g448796/U$1 ( \13193 , \13190 , \13191 , \13192 );
and \g451603/U$2 ( \13194 , \8335 , RIded23f8_856);
and \g451603/U$3 ( \13195 , RIded8c08_930, \8340 );
nor \g451603/U$1 ( \13196 , \13194 , \13195 );
and \g451602/U$2 ( \13197 , \8404 , RIee22ee8_4856);
and \g451602/U$3 ( \13198 , RIee25210_4881, \8351 );
nor \g451602/U$1 ( \13199 , \13197 , \13198 );
and \g455088/U$2 ( \13200 , \8313 , RIee238c0_4863);
and \g455088/U$3 ( \13201 , RIee24400_4871, \8323 );
nor \g455088/U$1 ( \13202 , \13200 , \13201 );
not \g449823/U$3 ( \13203 , \13202 );
not \g449823/U$4 ( \13204 , \8328 );
and \g449823/U$2 ( \13205 , \13203 , \13204 );
and \g449823/U$5 ( \13206 , \8359 , RIfcc5a68_7271);
nor \g449823/U$1 ( \13207 , \13205 , \13206 );
nand \g447623/U$1 ( \13208 , \13193 , \13196 , \13199 , \13207 );
nor \g445934/U$1 ( \13209 , \13188 , \13189 , \13208 );
and \g451600/U$2 ( \13210 , \8356 , RIee20e90_4833);
and \g451600/U$3 ( \13211 , RIfe8cca0_7946, \8417 );
nor \g451600/U$1 ( \13212 , \13210 , \13211 );
nand \g445561/U$1 ( \13213 , \13187 , \13209 , \13212 );
and \g444910/U$2 ( \13214 , \13213 , \8482 );
and \g448793/U$2 ( \13215 , RIe16d3d0_2620, \8414 );
and \g448793/U$3 ( \13216 , \8409 , RIde94850_314);
and \g448793/U$4 ( \13217 , RIdecccc8_794, \8330 );
nor \g448793/U$1 ( \13218 , \13215 , \13216 , \13217 );
and \g451594/U$2 ( \13219 , \8356 , RIdf1c2a0_1697);
and \g451594/U$3 ( \13220 , RIe1429c8_2135, \8359 );
nor \g451594/U$1 ( \13221 , \13219 , \13220 );
and \g455376/U$2 ( \13222 , \8313 , RIdf2ba20_1873);
and \g455376/U$3 ( \13223 , RIdf373c0_2005, \8323 );
nor \g455376/U$1 ( \13224 , \13222 , \13223 );
not \g449820/U$3 ( \13225 , \13224 );
not \g449820/U$4 ( \13226 , \8347 );
and \g449820/U$2 ( \13227 , \13225 , \13226 );
and \g449820/U$5 ( \13228 , \8351 , RIdecf9c8_826);
nor \g449820/U$1 ( \13229 , \13227 , \13228 );
and \g451592/U$2 ( \13230 , \8378 , RIe1591c8_2391);
and \g451592/U$3 ( \13231 , RIdeb37c8_506, \8417 );
nor \g451592/U$1 ( \13232 , \13230 , \13231 );
nand \g447621/U$1 ( \13233 , \13218 , \13221 , \13229 , \13232 );
and \g444910/U$3 ( \13234 , \9010 , \13233 );
nor \g444910/U$1 ( \13235 , \13214 , \13234 );
and \g446721/U$2 ( \13236 , \9041 , RIdec72c8_730);
and \g446721/U$3 ( \13237 , RIdec9fc8_762, \9043 );
nor \g446721/U$1 ( \13238 , \13236 , \13237 );
nor \g448382/U$1 ( \13239 , \8651 , \8325 );
and \g446722/U$2 ( \13240 , \13239 , RIdee6498_1084);
nor \g448316/U$1 ( \13241 , \8651 , \8516 );
and \g446722/U$3 ( \13242 , RIdeff998_1372, \13241 );
nor \g446722/U$1 ( \13243 , \13240 , \13242 );
nor \g448384/U$1 ( \13244 , \8651 , \8508 );
and \g446723/U$2 ( \13245 , \13244 , RIde7a798_187);
nor \g448383/U$1 ( \13246 , \8651 , \8318 );
and \g446723/U$3 ( \13247 , RIdedb200_957, \13246 );
nor \g446723/U$1 ( \13248 , \13245 , \13247 );
nand \g444585/U$1 ( \13249 , \13235 , \13238 , \13243 , \13248 );
and \g445927/U$2 ( \13250 , RIdf276a0_1825, \8409 );
and \g445927/U$3 ( \13251 , RIdf23cf8_1784, \8378 );
and \g448782/U$2 ( \13252 , RIee28780_4919, \8373 );
and \g448782/U$3 ( \13253 , \8383 , RIee29c98_4934);
and \g448782/U$4 ( \13254 , RIfcb73c8_7107, \8488 );
nor \g448782/U$1 ( \13255 , \13252 , \13253 , \13254 );
and \g451568/U$2 ( \13256 , \8335 , RIdf18a60_1657);
and \g451568/U$3 ( \13257 , RIfc83d20_6522, \8340 );
nor \g451568/U$1 ( \13258 , \13256 , \13257 );
and \g451566/U$2 ( \13259 , \8404 , RIee27538_4906);
and \g451566/U$3 ( \13260 , RIee2b318_4950, \8351 );
nor \g451566/U$1 ( \13261 , \13259 , \13260 );
and \g454414/U$2 ( \13262 , \8313 , RIfc51b90_5952);
and \g454414/U$3 ( \13263 , RIdf1ee38_1728, \8323 );
nor \g454414/U$1 ( \13264 , \13262 , \13263 );
not \g454413/U$1 ( \13265 , \13264 );
and \g449810/U$2 ( \13266 , \13265 , \8316 );
and \g449810/U$3 ( \13267 , RIfc83ff0_6524, \8359 );
nor \g449810/U$1 ( \13268 , \13266 , \13267 );
nand \g448167/U$1 ( \13269 , \13255 , \13258 , \13261 , \13268 );
nor \g445927/U$1 ( \13270 , \13250 , \13251 , \13269 );
and \g451565/U$2 ( \13271 , \8356 , RIfcdaa80_7510);
and \g451565/U$3 ( \13272 , RIdf299c8_1850, \8417 );
nor \g451565/U$1 ( \13273 , \13271 , \13272 );
and \g451563/U$2 ( \13274 , \8531 , RIfc51320_5946);
and \g451563/U$3 ( \13275 , RIdf25918_1804, \8412 );
nor \g451563/U$1 ( \13276 , \13274 , \13275 );
and \g445096/U$2 ( \13277 , \13270 , \13273 , \13276 );
nor \g445096/U$1 ( \13278 , \13277 , \8621 );
and \g445928/U$2 ( \13279 , RIdf05398_1436, \8414 );
and \g445928/U$3 ( \13280 , RIdeebe98_1148, \8319 );
and \g448784/U$2 ( \13281 , RIdf08098_1468, \8409 );
and \g448784/U$3 ( \13282 , \8531 , RIdef7298_1276);
and \g448784/U$4 ( \13283 , RIdef9f98_1308, \8488 );
nor \g448784/U$1 ( \13284 , \13281 , \13282 , \13283 );
and \g455140/U$2 ( \13285 , \8313 , RIdf10798_1564);
and \g455140/U$3 ( \13286 , RIdf13498_1596, \8323 );
nor \g455140/U$1 ( \13287 , \13285 , \13286 );
not \g449814/U$3 ( \13288 , \13287 );
not \g449814/U$4 ( \13289 , \8328 );
and \g449814/U$2 ( \13290 , \13288 , \13289 );
and \g449814/U$5 ( \13291 , \8417 , RIdf0ad98_1500);
nor \g449814/U$1 ( \13292 , \13290 , \13291 );
and \g453980/U$2 ( \13293 , \8404 , RIdf0da98_1532);
and \g453980/U$3 ( \13294 , RIdf16198_1628, \8351 );
nor \g453980/U$1 ( \13295 , \13293 , \13294 );
and \g451574/U$2 ( \13296 , \8356 , RIdef4598_1244);
and \g451574/U$3 ( \13297 , RIdefcc98_1340, \8359 );
nor \g451574/U$1 ( \13298 , \13296 , \13297 );
nand \g447616/U$1 ( \13299 , \13284 , \13292 , \13295 , \13298 );
nor \g445928/U$1 ( \13300 , \13279 , \13280 , \13299 );
and \g451573/U$2 ( \13301 , \8335 , RIdee9198_1116);
and \g451573/U$3 ( \13302 , RIdef1898_1212, \8340 );
nor \g451573/U$1 ( \13303 , \13301 , \13302 );
and \g451572/U$2 ( \13304 , \8326 , RIdeeeb98_1180);
and \g451572/U$3 ( \13305 , RIdf02698_1404, \8378 );
nor \g451572/U$1 ( \13306 , \13304 , \13305 );
and \g445097/U$2 ( \13307 , \13300 , \13303 , \13306 );
nor \g445097/U$1 ( \13308 , \13307 , \8477 );
or \g444376/U$1 ( \13309 , \13184 , \13249 , \13278 , \13308 );
and \g445923/U$2 ( \13310 , RIee35d40_5071, \8417 );
and \g445923/U$3 ( \13311 , RIe14ddc8_2263, \8356 );
and \g448778/U$2 ( \13312 , RIee36b50_5081, \8373 );
and \g448778/U$3 ( \13313 , \8330 , RIe1618c8_2487);
and \g448778/U$4 ( \13314 , RIe150ac8_2295, \8488 );
nor \g448778/U$1 ( \13315 , \13312 , \13313 , \13314 );
and \g451554/U$2 ( \13316 , \8335 , RIe1456c8_2167);
and \g451554/U$3 ( \13317 , RIfce0fc0_7582, \8340 );
nor \g451554/U$1 ( \13318 , \13316 , \13317 );
and \g451553/U$2 ( \13319 , \8404 , RIe15ebc8_2455);
and \g451553/U$3 ( \13320 , RIe1645c8_2519, \8351 );
nor \g451553/U$1 ( \13321 , \13319 , \13320 );
and \g454417/U$2 ( \13322 , \8313 , RIe1483c8_2199);
and \g454417/U$3 ( \13323 , RIe14b0c8_2231, \8323 );
nor \g454417/U$1 ( \13324 , \13322 , \13323 );
not \g454416/U$1 ( \13325 , \13324 );
and \g449578/U$2 ( \13326 , \13325 , \8316 );
and \g449578/U$3 ( \13327 , RIfc3ef90_5742, \8359 );
nor \g449578/U$1 ( \13328 , \13326 , \13327 );
nand \g448165/U$1 ( \13329 , \13315 , \13318 , \13321 , \13328 );
nor \g445923/U$1 ( \13330 , \13310 , \13311 , \13329 );
and \g451550/U$2 ( \13331 , \8378 , RIe1537c8_2327);
and \g451550/U$3 ( \13332 , RIfe8d7e0_7954, \8531 );
nor \g451550/U$1 ( \13333 , \13331 , \13332 );
and \g451548/U$2 ( \13334 , \8412 , RIe1564c8_2359);
and \g451548/U$3 ( \13335 , RIe15bec8_2423, \8409 );
nor \g451548/U$1 ( \13336 , \13334 , \13335 );
and \g445092/U$2 ( \13337 , \13330 , \13333 , \13336 );
nor \g445092/U$1 ( \13338 , \13337 , \8368 );
and \g445925/U$2 ( \13339 , RIfe8ce08_7947, \8409 );
and \g445925/U$3 ( \13340 , RIfe8d0d8_7949, \8378 );
and \g448780/U$2 ( \13341 , RIdf30610_1927, \8319 );
and \g448780/U$3 ( \13342 , \8326 , RIfe8d678_7953);
and \g448780/U$4 ( \13343 , RIee2ef90_4993, \8488 );
nor \g448780/U$1 ( \13344 , \13341 , \13342 , \13343 );
and \g450619/U$2 ( \13345 , \8335 , RIdf2e720_1905);
and \g450619/U$3 ( \13346 , RIdf34af8_1976, \8340 );
nor \g450619/U$1 ( \13347 , \13345 , \13346 );
and \g450666/U$2 ( \13348 , \8404 , RIee30d18_5014);
and \g450666/U$3 ( \13349 , RIee33e50_5049, \8351 );
nor \g450666/U$1 ( \13350 , \13348 , \13349 );
and \g454682/U$2 ( \13351 , \8313 , RIee319c0_5023);
and \g454682/U$3 ( \13352 , RIee32c08_5036, \8323 );
nor \g454682/U$1 ( \13353 , \13351 , \13352 );
not \g449809/U$3 ( \13354 , \13353 );
not \g449809/U$4 ( \13355 , \8328 );
and \g449809/U$2 ( \13356 , \13354 , \13355 );
and \g449809/U$5 ( \13357 , \8359 , RIfce9dc8_7683);
nor \g449809/U$1 ( \13358 , \13356 , \13357 );
nand \g447615/U$1 ( \13359 , \13344 , \13347 , \13350 , \13358 );
nor \g445925/U$1 ( \13360 , \13339 , \13340 , \13359 );
and \g451558/U$2 ( \13361 , \8356 , RIee2cdd0_4969);
and \g451558/U$3 ( \13362 , RIfe8cf70_7948, \8417 );
nor \g451558/U$1 ( \13363 , \13361 , \13362 );
and \g450788/U$2 ( \13364 , \8531 , RIfce51d8_7629);
and \g450788/U$3 ( \13365 , RIfe8d240_7950, \8414 );
nor \g450788/U$1 ( \13366 , \13364 , \13365 );
and \g445093/U$2 ( \13367 , \13360 , \13363 , \13366 );
nor \g445093/U$1 ( \13368 , \13367 , \8422 );
or \g444241/U$1 ( \13369 , \13309 , \13338 , \13368 );
_DC \g2c14/U$1 ( \13370 , \13369 , \8654 );
and \g450983/U$2 ( \13371 , \8356 , RIe14dc60_2262);
and \g450983/U$3 ( \13372 , RIe15bd60_2422, \8409 );
nor \g450983/U$1 ( \13373 , \13371 , \13372 );
and \g445793/U$2 ( \13374 , RIe156360_2358, \8414 );
and \g445793/U$3 ( \13375 , RIfe94158_8029, \8417 );
and \g448614/U$2 ( \13376 , RIfe942c0_8030, \8373 );
and \g448614/U$3 ( \13377 , \8383 , RIe161760_2486);
and \g448614/U$4 ( \13378 , RIe150960_2294, \8488 );
nor \g448614/U$1 ( \13379 , \13376 , \13377 , \13378 );
and \g450987/U$2 ( \13380 , \8335 , RIe145560_2166);
and \g450987/U$3 ( \13381 , RIfc5c2e8_6071, \8340 );
nor \g450987/U$1 ( \13382 , \13380 , \13381 );
and \g450985/U$2 ( \13383 , \8404 , RIe15ea60_2454);
and \g450985/U$3 ( \13384 , RIe164460_2518, \8351 );
nor \g450985/U$1 ( \13385 , \13383 , \13384 );
and \g454520/U$2 ( \13386 , \8313 , RIe148260_2198);
and \g454520/U$3 ( \13387 , RIe14af60_2230, \8323 );
nor \g454520/U$1 ( \13388 , \13386 , \13387 );
not \g454519/U$1 ( \13389 , \13388 );
and \g449640/U$2 ( \13390 , \13389 , \8316 );
and \g449640/U$3 ( \13391 , RIfe94428_8031, \8359 );
nor \g449640/U$1 ( \13392 , \13390 , \13391 );
nand \g448147/U$1 ( \13393 , \13379 , \13382 , \13385 , \13392 );
nor \g445793/U$1 ( \13394 , \13374 , \13375 , \13393 );
and \g450982/U$2 ( \13395 , \8378 , RIe153660_2326);
and \g450982/U$3 ( \13396 , RIfe94590_8032, \8531 );
nor \g450982/U$1 ( \13397 , \13395 , \13396 );
nand \g445530/U$1 ( \13398 , \13373 , \13394 , \13397 );
and \g444849/U$2 ( \13399 , \13398 , \8369 );
and \g448613/U$2 ( \13400 , RIfcc88d0_7304, \8531 );
and \g448613/U$3 ( \13401 , \8486 , RIee2ee28_4992);
and \g448613/U$4 ( \13402 , RIee32aa0_5035, \8330 );
nor \g448613/U$1 ( \13403 , \13400 , \13401 , \13402 );
and \g450981/U$2 ( \13404 , \8356 , RIee2cc68_4968);
and \g450981/U$3 ( \13405 , RIfcdd780_7542, \8359 );
nor \g450981/U$1 ( \13406 , \13404 , \13405 );
and \g454372/U$2 ( \13407 , \8313 , RIdf3c118_2060);
and \g454372/U$3 ( \13408 , RIdf3e2d8_2084, \8323 );
nor \g454372/U$1 ( \13409 , \13407 , \13408 );
not \g449639/U$3 ( \13410 , \13409 );
not \g449639/U$4 ( \13411 , \8376 );
and \g449639/U$2 ( \13412 , \13410 , \13411 );
and \g449639/U$5 ( \13413 , \8351 , RIee33ce8_5048);
nor \g449639/U$1 ( \13414 , \13412 , \13413 );
and \g450980/U$2 ( \13415 , \8378 , RIdf39df0_2035);
and \g450980/U$3 ( \13416 , RIe140538_2109, \8417 );
nor \g450980/U$1 ( \13417 , \13415 , \13416 );
nand \g447518/U$1 ( \13418 , \13403 , \13406 , \13414 , \13417 );
and \g444849/U$3 ( \13419 , \9266 , \13418 );
nor \g444849/U$1 ( \13420 , \13399 , \13419 );
and \g446592/U$2 ( \13421 , \9288 , RIfc5d530_6084);
and \g446592/U$3 ( \13422 , RIee31858_5022, \9290 );
nor \g446592/U$1 ( \13423 , \13421 , \13422 );
nor \g448419/U$1 ( \13424 , \8422 , \8325 );
and \g446593/U$2 ( \13425 , \13424 , RIdf32aa0_1953);
nor \g448427/U$1 ( \13426 , \8422 , \8516 );
and \g446593/U$3 ( \13427 , RIdf34990_1975, \13426 );
nor \g446593/U$1 ( \13428 , \13425 , \13427 );
and \g446594/U$2 ( \13429 , \9299 , RIdf2e5b8_1904);
and \g446594/U$3 ( \13430 , RIdf304a8_1926, \9301 );
nor \g446594/U$1 ( \13431 , \13429 , \13430 );
nand \g444563/U$1 ( \13432 , \13420 , \13423 , \13428 , \13431 );
and \g450972/U$2 ( \13433 , \8317 , RIdedb098_956);
and \g450972/U$3 ( \13434 , RIdee6330_1083, \8326 );
nor \g450972/U$1 ( \13435 , \13433 , \13434 );
and \g445791/U$2 ( \13436 , RIdec9e60_761, \8373 );
and \g445791/U$3 ( \13437 , RIde7a450_186, \8335 );
and \g448610/U$2 ( \13438 , RIe16d268_2619, \8414 );
and \g448610/U$3 ( \13439 , \8409 , RIde94508_313);
and \g448610/U$4 ( \13440 , RIdeccb60_793, \8383 );
nor \g448610/U$1 ( \13441 , \13438 , \13439 , \13440 );
and \g450975/U$2 ( \13442 , \8356 , RIdf1c138_1696);
and \g450975/U$3 ( \13443 , RIe142860_2134, \8359 );
nor \g450975/U$1 ( \13444 , \13442 , \13443 );
and \g454912/U$2 ( \13445 , \8313 , RIdf2b8b8_1872);
and \g454912/U$3 ( \13446 , RIdf37258_2004, \8323 );
nor \g454912/U$1 ( \13447 , \13445 , \13446 );
not \g449637/U$3 ( \13448 , \13447 );
not \g449637/U$4 ( \13449 , \8347 );
and \g449637/U$2 ( \13450 , \13448 , \13449 );
and \g449637/U$5 ( \13451 , \8351 , RIdecf860_825);
nor \g449637/U$1 ( \13452 , \13450 , \13451 );
and \g450973/U$2 ( \13453 , \8378 , RIe159060_2390);
and \g450973/U$3 ( \13454 , RIdeb3660_505, \8417 );
nor \g450973/U$1 ( \13455 , \13453 , \13454 );
nand \g447517/U$1 ( \13456 , \13441 , \13444 , \13452 , \13455 );
nor \g445791/U$1 ( \13457 , \13436 , \13437 , \13456 );
and \g450970/U$2 ( \13458 , \8340 , RIdeff830_1371);
and \g450970/U$3 ( \13459 , RIdec7160_729, \8404 );
nor \g450970/U$1 ( \13460 , \13458 , \13459 );
nand \g445528/U$1 ( \13461 , \13435 , \13457 , \13460 );
and \g444872/U$2 ( \13462 , \13461 , \9010 );
and \g448609/U$2 ( \13463 , RIfcb2940_7054, \8373 );
and \g448609/U$3 ( \13464 , \8383 , RIfe946f8_8033);
and \g448609/U$4 ( \13465 , RIee269f8_4898, \8488 );
nor \g448609/U$1 ( \13466 , \13463 , \13464 , \13465 );
and \g450966/U$2 ( \13467 , \8335 , RIfea9170_8240);
and \g450966/U$3 ( \13468 , RIee26188_4892, \8340 );
nor \g450966/U$1 ( \13469 , \13467 , \13468 );
and \g450965/U$2 ( \13470 , \8404 , RIee273d0_4905);
and \g450965/U$3 ( \13471 , RIee2b1b0_4949, \8351 );
nor \g450965/U$1 ( \13472 , \13470 , \13471 );
and \g454317/U$2 ( \13473 , \8313 , RIee25d50_4889);
and \g454317/U$3 ( \13474 , RIfe94c98_8037, \8323 );
nor \g454317/U$1 ( \13475 , \13473 , \13474 );
not \g454316/U$1 ( \13476 , \13475 );
and \g449636/U$2 ( \13477 , \13476 , \8316 );
and \g449636/U$3 ( \13478 , RIee26f98_4902, \8359 );
nor \g449636/U$1 ( \13479 , \13477 , \13478 );
nand \g448146/U$1 ( \13480 , \13466 , \13469 , \13472 , \13479 );
and \g444872/U$3 ( \13481 , \8752 , \13480 );
nor \g444872/U$1 ( \13482 , \13462 , \13481 );
and \g446589/U$2 ( \13483 , \11516 , RIdf27538_1824);
and \g446589/U$3 ( \13484 , RIfe949c8_8035, \11518 );
nor \g446589/U$1 ( \13485 , \13483 , \13484 );
nor \g448441/U$1 ( \13486 , \8621 , \8520 );
and \g446590/U$2 ( \13487 , \13486 , RIee26458_4894);
nor \g448440/U$1 ( \13488 , \8621 , \8524 );
and \g446590/U$3 ( \13489 , RIee26728_4896, \13488 );
nor \g446590/U$1 ( \13490 , \13487 , \13489 );
and \g446591/U$2 ( \13491 , \11521 , RIfe94860_8034);
and \g446591/U$3 ( \13492 , RIfe94b30_8036, \11523 );
nor \g446591/U$1 ( \13493 , \13491 , \13492 );
nand \g444562/U$1 ( \13494 , \13482 , \13485 , \13490 , \13493 );
and \g445787/U$2 ( \13495 , RIee1fae0_4819, \8371 );
and \g445787/U$3 ( \13496 , RIdea1708_377, \8319 );
and \g448605/U$2 ( \13497 , RIee1e460_4803, \8531 );
and \g448605/U$3 ( \13498 , \8488 , RIdeb0960_473);
and \g448605/U$4 ( \13499 , RIdec1760_665, \8383 );
nor \g448605/U$1 ( \13500 , \13497 , \13498 , \13499 );
and \g450951/U$2 ( \13501 , \8356 , RIdeadc60_441);
and \g450951/U$3 ( \13502 , RIee1eb68_4808, \8359 );
nor \g450951/U$1 ( \13503 , \13501 , \13502 );
and \g454312/U$2 ( \13504 , \8313 , RIdeb9060_569);
and \g454312/U$3 ( \13505 , RIdebbd60_601, \8323 );
nor \g454312/U$1 ( \13506 , \13504 , \13505 );
not \g449631/U$3 ( \13507 , \13506 );
not \g449631/U$4 ( \13508 , \8376 );
and \g449631/U$2 ( \13509 , \13507 , \13508 );
and \g449631/U$5 ( \13510 , \8351 , RIdec4460_697);
nor \g449631/U$1 ( \13511 , \13509 , \13510 );
and \g450950/U$2 ( \13512 , \8378 , RIdeb6360_537);
and \g450950/U$3 ( \13513 , RIee1f108_4812, \8417 );
nor \g450950/U$1 ( \13514 , \13512 , \13513 );
nand \g447510/U$1 ( \13515 , \13500 , \13503 , \13511 , \13514 );
nor \g445787/U$1 ( \13516 , \13495 , \13496 , \13515 );
and \g450948/U$2 ( \13517 , \8335 , RIde9ae08_345);
and \g450948/U$3 ( \13518 , RIee1d7b8_4794, \8340 );
nor \g450948/U$1 ( \13519 , \13517 , \13518 );
and \g450947/U$2 ( \13520 , \8324 , RIdea8008_409);
and \g450947/U$3 ( \13521 , RIdebea60_633, \8404 );
nor \g450947/U$1 ( \13522 , \13520 , \13521 );
and \g444993/U$2 ( \13523 , \13516 , \13519 , \13522 );
nor \g444993/U$1 ( \13524 , \13523 , \8589 );
and \g445789/U$2 ( \13525 , RIfe95670_8044, \8371 );
and \g445789/U$3 ( \13526 , RIfea9440_8242, \8335 );
and \g448606/U$2 ( \13527 , RIfe95940_8046, \8414 );
and \g448606/U$3 ( \13528 , \8409 , RIfe95238_8041);
and \g448606/U$4 ( \13529 , RIfe95508_8043, \8383 );
nor \g448606/U$1 ( \13530 , \13527 , \13528 , \13529 );
and \g450960/U$2 ( \13531 , \8356 , RIee19438_4746);
and \g450960/U$3 ( \13532 , RIee1a0e0_4755, \8359 );
nor \g450960/U$1 ( \13533 , \13531 , \13532 );
and \g454464/U$2 ( \13534 , \8313 , RIee19870_4749);
and \g454464/U$3 ( \13535 , RIee19ca8_4752, \8323 );
nor \g454464/U$1 ( \13536 , \13534 , \13535 );
not \g449632/U$3 ( \13537 , \13536 );
not \g449632/U$4 ( \13538 , \8347 );
and \g449632/U$2 ( \13539 , \13537 , \13538 );
and \g449632/U$5 ( \13540 , \8351 , RIfe957d8_8045);
nor \g449632/U$1 ( \13541 , \13539 , \13540 );
and \g450957/U$2 ( \13542 , \8378 , RIfe953a0_8042);
and \g450957/U$3 ( \13543 , RIfe95aa8_8047, \8417 );
nor \g450957/U$1 ( \13544 , \13542 , \13543 );
nand \g447514/U$1 ( \13545 , \13530 , \13533 , \13541 , \13544 );
nor \g445789/U$1 ( \13546 , \13525 , \13526 , \13545 );
and \g450953/U$2 ( \13547 , \8340 , RIee38ba8_5104);
and \g450953/U$3 ( \13548 , RIee1a7e8_4760, \8404 );
nor \g450953/U$1 ( \13549 , \13547 , \13548 );
and \g450954/U$2 ( \13550 , \8319 , RIee384a0_5099);
and \g450954/U$3 ( \13551 , RIfe95c10_8048, \8324 );
nor \g450954/U$1 ( \13552 , \13550 , \13551 );
and \g444995/U$2 ( \13553 , \13546 , \13549 , \13552 );
nor \g444995/U$1 ( \13554 , \13553 , \8558 );
or \g444384/U$1 ( \13555 , \13432 , \13494 , \13524 , \13554 );
and \g445785/U$2 ( \13556 , RIdf10630_1563, \8371 );
and \g445785/U$3 ( \13557 , RIdeebd30_1147, \8317 );
and \g448603/U$2 ( \13558 , RIdef7130_1275, \8531 );
and \g448603/U$3 ( \13559 , \8486 , RIdef9e30_1307);
and \g448603/U$4 ( \13560 , RIdf13330_1595, \8383 );
nor \g448603/U$1 ( \13561 , \13558 , \13559 , \13560 );
and \g450944/U$2 ( \13562 , \8356 , RIdef4430_1243);
and \g450944/U$3 ( \13563 , RIdefcb30_1339, \8359 );
nor \g450944/U$1 ( \13564 , \13562 , \13563 );
and \g454463/U$2 ( \13565 , \8313 , RIdf05230_1435);
and \g454463/U$3 ( \13566 , RIdf07f30_1467, \8323 );
nor \g454463/U$1 ( \13567 , \13565 , \13566 );
not \g449629/U$3 ( \13568 , \13567 );
not \g449629/U$4 ( \13569 , \8376 );
and \g449629/U$2 ( \13570 , \13568 , \13569 );
and \g449629/U$5 ( \13571 , \8351 , RIdf16030_1627);
nor \g449629/U$1 ( \13572 , \13570 , \13571 );
and \g450942/U$2 ( \13573 , \8378 , RIdf02530_1403);
and \g450942/U$3 ( \13574 , RIdf0ac30_1499, \8417 );
nor \g450942/U$1 ( \13575 , \13573 , \13574 );
nand \g447509/U$1 ( \13576 , \13561 , \13564 , \13572 , \13575 );
nor \g445785/U$1 ( \13577 , \13556 , \13557 , \13576 );
and \g450941/U$2 ( \13578 , \8335 , RIdee9030_1115);
and \g450941/U$3 ( \13579 , RIdef1730_1211, \8340 );
nor \g450941/U$1 ( \13580 , \13578 , \13579 );
and \g450940/U$2 ( \13581 , \8324 , RIdeeea30_1179);
and \g450940/U$3 ( \13582 , RIdf0d930_1531, \8404 );
nor \g450940/U$1 ( \13583 , \13581 , \13582 );
and \g444990/U$2 ( \13584 , \13577 , \13580 , \13583 );
nor \g444990/U$1 ( \13585 , \13584 , \8477 );
and \g445783/U$2 ( \13586 , RIee23758_4862, \8373 );
and \g445783/U$3 ( \13587 , RIfe95d78_8049, \8319 );
and \g448601/U$2 ( \13588 , RIfe94e00_8038, \8414 );
and \g448601/U$3 ( \13589 , \8409 , RIfe94f68_8039);
and \g448601/U$4 ( \13590 , RIee24298_4870, \8330 );
nor \g448601/U$1 ( \13591 , \13588 , \13589 , \13590 );
and \g450936/U$2 ( \13592 , \8356 , RIfc5dad0_6088);
and \g450936/U$3 ( \13593 , RIee22ab0_4853, \8359 );
nor \g450936/U$1 ( \13594 , \13592 , \13593 );
and \g454424/U$2 ( \13595 , \8313 , RIfca46d8_6893);
and \g454424/U$3 ( \13596 , RIee21e08_4844, \8323 );
nor \g454424/U$1 ( \13597 , \13595 , \13596 );
not \g449628/U$3 ( \13598 , \13597 );
not \g449628/U$4 ( \13599 , \8347 );
and \g449628/U$2 ( \13600 , \13598 , \13599 );
and \g449628/U$5 ( \13601 , \8351 , RIee250a8_4880);
nor \g449628/U$1 ( \13602 , \13600 , \13601 );
and \g450935/U$2 ( \13603 , \8378 , RIdeddd98_988);
and \g450935/U$3 ( \13604 , RIfe950d0_8040, \8417 );
nor \g450935/U$1 ( \13605 , \13603 , \13604 );
nand \g447507/U$1 ( \13606 , \13591 , \13594 , \13602 , \13605 );
nor \g445783/U$1 ( \13607 , \13586 , \13587 , \13606 );
and \g450934/U$2 ( \13608 , \8335 , RIfe95ee0_8050);
and \g450934/U$3 ( \13609 , RIfeaa250_8252, \8340 );
nor \g450934/U$1 ( \13610 , \13608 , \13609 );
and \g450933/U$2 ( \13611 , \8326 , RIfe96048_8051);
and \g450933/U$3 ( \13612 , RIee22d80_4855, \8404 );
nor \g450933/U$1 ( \13613 , \13611 , \13612 );
and \g444989/U$2 ( \13614 , \13607 , \13610 , \13613 );
nor \g444989/U$1 ( \13615 , \13614 , \8481 );
or \g444196/U$1 ( \13616 , \13555 , \13585 , \13615 );
_DC \g2c99/U$1 ( \13617 , \13616 , \8654 );
and \g446609/U$2 ( \13618 , \8969 , RIee22c18_4854);
and \g446609/U$3 ( \13619 , RIee235f0_4861, \8971 );
nor \g446609/U$1 ( \13620 , \13618 , \13619 );
and \g445817/U$2 ( \13621 , RIee24f40_4879, \8351 );
and \g445817/U$3 ( \13622 , RIee24130_4869, \8383 );
and \g448641/U$2 ( \13623 , RIfe93ff0_8028, \8326 );
and \g448641/U$3 ( \13624 , \8523 , RIfc68390_6208);
and \g448641/U$4 ( \13625 , RIee21ca0_4843, \8488 );
nor \g448641/U$1 ( \13626 , \13623 , \13624 , \13625 );
and \g451088/U$2 ( \13627 , \8356 , RIee20d28_4832);
and \g451088/U$3 ( \13628 , RIfc684f8_6209, \8359 );
nor \g451088/U$1 ( \13629 , \13627 , \13628 );
and \g454366/U$2 ( \13630 , \8313 , RIdee0228_1014);
and \g454366/U$3 ( \13631 , RIdee1fb0_1035, \8323 );
nor \g454366/U$1 ( \13632 , \13630 , \13631 );
not \g449666/U$3 ( \13633 , \13632 );
not \g449666/U$4 ( \13634 , \8376 );
and \g449666/U$2 ( \13635 , \13633 , \13634 );
and \g449666/U$5 ( \13636 , \8340 , RIded8aa0_929);
nor \g449666/U$1 ( \13637 , \13635 , \13636 );
and \g451087/U$2 ( \13638 , \8378 , RIdeddc30_987);
and \g451087/U$3 ( \13639 , RIfe93d20_8026, \8417 );
nor \g451087/U$1 ( \13640 , \13638 , \13639 );
nand \g447534/U$1 ( \13641 , \13626 , \13629 , \13637 , \13640 );
nor \g445817/U$1 ( \13642 , \13621 , \13622 , \13641 );
not \g444813/U$3 ( \13643 , \13642 );
not \g444813/U$4 ( \13644 , \8481 );
and \g444813/U$2 ( \13645 , \13643 , \13644 );
and \g445819/U$2 ( \13646 , RIdf15ec8_1626, \8351 );
and \g445819/U$3 ( \13647 , RIdf0d7c8_1530, \8404 );
and \g448643/U$2 ( \13648 , RIdeee8c8_1178, \8326 );
and \g448643/U$3 ( \13649 , \8531 , RIdef6fc8_1274);
and \g448643/U$4 ( \13650 , RIdef9cc8_1306, \8488 );
nor \g448643/U$1 ( \13651 , \13648 , \13649 , \13650 );
and \g451097/U$2 ( \13652 , \8356 , RIdef42c8_1242);
and \g451097/U$3 ( \13653 , RIdefc9c8_1338, \8359 );
nor \g451097/U$1 ( \13654 , \13652 , \13653 );
and \g455206/U$2 ( \13655 , \8313 , RIdf050c8_1434);
and \g455206/U$3 ( \13656 , RIdf07dc8_1466, \8323 );
nor \g455206/U$1 ( \13657 , \13655 , \13656 );
not \g449669/U$3 ( \13658 , \13657 );
not \g449669/U$4 ( \13659 , \8376 );
and \g449669/U$2 ( \13660 , \13658 , \13659 );
and \g449669/U$5 ( \13661 , \8340 , RIdef15c8_1210);
nor \g449669/U$1 ( \13662 , \13660 , \13661 );
and \g451095/U$2 ( \13663 , \8378 , RIdf023c8_1402);
and \g451095/U$3 ( \13664 , RIdf0aac8_1498, \8417 );
nor \g451095/U$1 ( \13665 , \13663 , \13664 );
nand \g447536/U$1 ( \13666 , \13651 , \13654 , \13662 , \13665 );
nor \g445819/U$1 ( \13667 , \13646 , \13647 , \13666 );
and \g451093/U$2 ( \13668 , \8335 , RIdee8ec8_1114);
and \g451093/U$3 ( \13669 , RIdf131c8_1594, \8383 );
nor \g451093/U$1 ( \13670 , \13668 , \13669 );
and \g451092/U$2 ( \13671 , \8319 , RIdeebbc8_1146);
and \g451092/U$3 ( \13672 , RIdf104c8_1562, \8373 );
nor \g451092/U$1 ( \13673 , \13671 , \13672 );
and \g445015/U$2 ( \13674 , \13667 , \13670 , \13673 );
nor \g445015/U$1 ( \13675 , \13674 , \8477 );
nor \g444813/U$1 ( \13676 , \13645 , \13675 );
and \g446608/U$2 ( \13677 , \8509 , RIfe93e88_8027);
and \g446608/U$3 ( \13678 , RIded45b8_880, \8511 );
nor \g446608/U$1 ( \13679 , \13677 , \13678 );
nand \g444420/U$1 ( \13680 , \13620 , \13676 , \13679 );
and \g448646/U$2 ( \13681 , RIe1561f8_2357, \8414 );
and \g448646/U$3 ( \13682 , \8409 , RIe15bbf8_2421);
and \g448646/U$4 ( \13683 , RIe14adf8_2229, \8324 );
nor \g448646/U$1 ( \13684 , \13681 , \13682 , \13683 );
and \g451100/U$2 ( \13685 , \8356 , RIe14daf8_2261);
and \g451100/U$3 ( \13686 , RIfc3ee28_5741, \8359 );
nor \g451100/U$1 ( \13687 , \13685 , \13686 );
and \g455269/U$2 ( \13688 , \8313 , RIfce6c90_7648);
and \g455269/U$3 ( \13689 , RIe1507f8_2293, \8323 );
nor \g455269/U$1 ( \13690 , \13688 , \13689 );
not \g449671/U$3 ( \13691 , \13690 );
not \g449671/U$4 ( \13692 , \8347 );
and \g449671/U$2 ( \13693 , \13691 , \13692 );
and \g449671/U$5 ( \13694 , \8340 , RIfcca7c0_7326);
nor \g449671/U$1 ( \13695 , \13693 , \13694 );
and \g451099/U$2 ( \13696 , \8378 , RIe1534f8_2325);
and \g451099/U$3 ( \13697 , RIee35bd8_5070, \8417 );
nor \g451099/U$1 ( \13698 , \13696 , \13697 );
nand \g447537/U$1 ( \13699 , \13684 , \13687 , \13695 , \13698 );
and \g444757/U$2 ( \13700 , \13699 , \8369 );
and \g445820/U$2 ( \13701 , RIdf3bfb0_2059, \8412 );
and \g445820/U$3 ( \13702 , RIee2cb00_4967, \8356 );
and \g448647/U$2 ( \13703 , RIdf30340_1925, \8317 );
and \g448647/U$3 ( \13704 , \8326 , RIdf32938_1952);
and \g448647/U$4 ( \13705 , RIfe93618_8021, \8409 );
nor \g448647/U$1 ( \13706 , \13703 , \13704 , \13705 );
and \g451106/U$2 ( \13707 , \8335 , RIdf2e450_1903);
and \g451106/U$3 ( \13708 , RIfe93bb8_8025, \8340 );
nor \g451106/U$1 ( \13709 , \13707 , \13708 );
and \g451105/U$2 ( \13710 , \8404 , RIee30bb0_5013);
and \g451105/U$3 ( \13711 , RIee33b80_5047, \8351 );
nor \g451105/U$1 ( \13712 , \13710 , \13711 );
and \g454371/U$2 ( \13713 , \8313 , RIee316f0_5021);
and \g454371/U$3 ( \13714 , RIee32938_5034, \8323 );
nor \g454371/U$1 ( \13715 , \13713 , \13714 );
not \g449672/U$3 ( \13716 , \13715 );
not \g449672/U$4 ( \13717 , \8328 );
and \g449672/U$2 ( \13718 , \13716 , \13717 );
and \g449672/U$5 ( \13719 , \8417 , RIe1403d0_2108);
nor \g449672/U$1 ( \13720 , \13718 , \13719 );
nand \g447538/U$1 ( \13721 , \13706 , \13709 , \13712 , \13720 );
nor \g445820/U$1 ( \13722 , \13701 , \13702 , \13721 );
and \g451104/U$2 ( \13723 , \8378 , RIfe934b0_8020);
and \g451104/U$3 ( \13724 , RIfcd0d00_7398, \8359 );
nor \g451104/U$1 ( \13725 , \13723 , \13724 );
and \g451103/U$2 ( \13726 , \8531 , RIee2e720_4987);
and \g451103/U$3 ( \13727 , RIee2ecc0_4991, \8488 );
nor \g451103/U$1 ( \13728 , \13726 , \13727 );
and \g445017/U$2 ( \13729 , \13722 , \13725 , \13728 );
nor \g445017/U$1 ( \13730 , \13729 , \8422 );
nor \g444757/U$1 ( \13731 , \13700 , \13730 );
and \g446612/U$2 ( \13732 , \8426 , RIe15e8f8_2453);
and \g446612/U$3 ( \13733 , RIee369e8_5080, \8428 );
nor \g446612/U$1 ( \13734 , \13732 , \13733 );
nor \g448396/U$1 ( \13735 , \8368 , \8382 );
and \g446611/U$2 ( \13736 , \13735 , RIe1615f8_2485);
nor \g448320/U$1 ( \13737 , \8368 , \9295 );
and \g446611/U$3 ( \13738 , RIe1642f8_2517, \13737 );
nor \g446611/U$1 ( \13739 , \13736 , \13738 );
and \g446613/U$2 ( \13740 , \8707 , RIe1453f8_2165);
and \g446613/U$3 ( \13741 , RIe1480f8_2197, \8709 );
nor \g446613/U$1 ( \13742 , \13740 , \13741 );
nand \g444460/U$1 ( \13743 , \13731 , \13734 , \13739 , \13742 );
and \g445812/U$2 ( \13744 , RIdeb8ef8_568, \8412 );
and \g445812/U$3 ( \13745 , RIdeadaf8_440, \8356 );
and \g448637/U$2 ( \13746 , RIdebbbf8_600, \8409 );
and \g448637/U$3 ( \13747 , \8371 , RIfcc6cb0_7284);
and \g448637/U$4 ( \13748 , RIdec15f8_664, \8383 );
nor \g448637/U$1 ( \13749 , \13746 , \13747 , \13748 );
and \g451074/U$2 ( \13750 , \8335 , RIde9aac0_344);
and \g451074/U$3 ( \13751 , RIfc5d3c8_6083, \8340 );
nor \g451074/U$1 ( \13752 , \13750 , \13751 );
and \g451073/U$2 ( \13753 , \8404 , RIdebe8f8_632);
and \g451073/U$3 ( \13754 , RIdec42f8_696, \8351 );
nor \g451073/U$1 ( \13755 , \13753 , \13754 );
and \g454359/U$2 ( \13756 , \8313 , RIdea13c0_376);
and \g454359/U$3 ( \13757 , RIdea7cc0_408, \8323 );
nor \g454359/U$1 ( \13758 , \13756 , \13757 );
not \g454358/U$1 ( \13759 , \13758 );
and \g449663/U$2 ( \13760 , \13759 , \8316 );
and \g449663/U$3 ( \13761 , RIfe93780_8022, \8417 );
nor \g449663/U$1 ( \13762 , \13760 , \13761 );
nand \g448150/U$1 ( \13763 , \13749 , \13752 , \13755 , \13762 );
nor \g445812/U$1 ( \13764 , \13744 , \13745 , \13763 );
and \g451072/U$2 ( \13765 , \8378 , RIdeb61f8_536);
and \g451072/U$3 ( \13766 , RIee1ea00_4807, \8359 );
nor \g451072/U$1 ( \13767 , \13765 , \13766 );
and \g451071/U$2 ( \13768 , \8531 , RIee1e2f8_4802);
and \g451071/U$3 ( \13769 , RIdeb07f8_472, \8488 );
nor \g451071/U$1 ( \13770 , \13768 , \13769 );
and \g445011/U$2 ( \13771 , \13764 , \13767 , \13770 );
nor \g445011/U$1 ( \13772 , \13771 , \8589 );
and \g445815/U$2 ( \13773 , RIfc58238_6025, \8351 );
and \g445815/U$3 ( \13774 , RIfc59750_6040, \8404 );
and \g448638/U$2 ( \13775 , RIe16ab08_2591, \8326 );
and \g448638/U$3 ( \13776 , \8531 , RIfc90a70_6668);
and \g448638/U$4 ( \13777 , RIfc976b8_6745, \8488 );
nor \g448638/U$1 ( \13778 , \13775 , \13776 , \13777 );
and \g451081/U$2 ( \13779 , \8356 , RIfc60500_6118);
and \g451081/U$3 ( \13780 , RIfc5f420_6106, \8359 );
nor \g451081/U$1 ( \13781 , \13779 , \13780 );
and \g454151/U$2 ( \13782 , \8313 , RIde88370_254);
and \g454151/U$3 ( \13783 , RIfe938e8_8023, \8323 );
nor \g454151/U$1 ( \13784 , \13782 , \13783 );
not \g449664/U$3 ( \13785 , \13784 );
not \g449664/U$4 ( \13786 , \8376 );
and \g449664/U$2 ( \13787 , \13785 , \13786 );
and \g449664/U$5 ( \13788 , \8340 , RIee38a40_5103);
nor \g449664/U$1 ( \13789 , \13787 , \13788 );
and \g451079/U$2 ( \13790 , \8378 , RIde83e88_233);
and \g451079/U$3 ( \13791 , RIfe93a50_8024, \8417 );
nor \g451079/U$1 ( \13792 , \13790 , \13791 );
nand \g447533/U$1 ( \13793 , \13778 , \13781 , \13789 , \13792 );
nor \g445815/U$1 ( \13794 , \13773 , \13774 , \13793 );
and \g451077/U$2 ( \13795 , \8335 , RIe166ff8_2549);
and \g451077/U$3 ( \13796 , RIfcc3b78_7249, \8330 );
nor \g451077/U$1 ( \13797 , \13795 , \13796 );
and \g451076/U$2 ( \13798 , \8319 , RIe169488_2575);
and \g451076/U$3 ( \13799 , RIfc7d0d8_6445, \8373 );
nor \g451076/U$1 ( \13800 , \13798 , \13799 );
and \g445012/U$2 ( \13801 , \13794 , \13797 , \13800 );
nor \g445012/U$1 ( \13802 , \13801 , \8558 );
or \g444308/U$1 ( \13803 , \13680 , \13743 , \13772 , \13802 );
and \g445809/U$2 ( \13804 , RIfe93348_8019, \8414 );
and \g445809/U$3 ( \13805 , RIdf22510_1767, \8531 );
and \g448632/U$2 ( \13806 , RIfe931e0_8018, \8409 );
and \g448632/U$3 ( \13807 , \8373 , RIfc67148_6195);
and \g448632/U$4 ( \13808 , RIee29b30_4933, \8383 );
nor \g448632/U$1 ( \13809 , \13806 , \13807 , \13808 );
and \g451061/U$2 ( \13810 , \8335 , RIfea7c58_8225);
and \g451061/U$3 ( \13811 , RIdf20ff8_1752, \8340 );
nor \g451061/U$1 ( \13812 , \13810 , \13811 );
and \g451060/U$2 ( \13813 , \8404 , RIfc6fb18_6293);
and \g451060/U$3 ( \13814 , RIee2b048_4948, \8351 );
nor \g451060/U$1 ( \13815 , \13813 , \13814 );
and \g454353/U$2 ( \13816 , \8313 , RIdf1aab8_1680);
and \g454353/U$3 ( \13817 , RIdf1ecd0_1727, \8323 );
nor \g454353/U$1 ( \13818 , \13816 , \13817 );
not \g454352/U$1 ( \13819 , \13818 );
and \g449660/U$2 ( \13820 , \13819 , \8316 );
and \g449660/U$3 ( \13821 , RIdf29860_1849, \8417 );
nor \g449660/U$1 ( \13822 , \13820 , \13821 );
nand \g448149/U$1 ( \13823 , \13809 , \13812 , \13815 , \13822 );
nor \g445809/U$1 ( \13824 , \13804 , \13805 , \13823 );
and \g451056/U$2 ( \13825 , \8356 , RIfcea7a0_7690);
and \g451056/U$3 ( \13826 , RIfc672b0_6196, \8359 );
nor \g451056/U$1 ( \13827 , \13825 , \13826 );
and \g451057/U$2 ( \13828 , \8378 , RIfe93078_8017);
and \g451057/U$3 ( \13829 , RIfca8788_6939, \8488 );
nor \g451057/U$1 ( \13830 , \13828 , \13829 );
and \g445008/U$2 ( \13831 , \13824 , \13827 , \13830 );
nor \g445008/U$1 ( \13832 , \13831 , \8621 );
and \g445811/U$2 ( \13833 , RIdec9cf8_760, \8371 );
and \g445811/U$3 ( \13834 , RIdecc9f8_792, \8383 );
and \g448634/U$2 ( \13835 , RIdee61c8_1082, \8326 );
and \g448634/U$3 ( \13836 , \8531 , RIdf2b750_1871);
and \g448634/U$4 ( \13837 , RIdf370f0_2003, \8488 );
nor \g448634/U$1 ( \13838 , \13835 , \13836 , \13837 );
and \g451069/U$2 ( \13839 , \8356 , RIdf1bfd0_1695);
and \g451069/U$3 ( \13840 , RIe1426f8_2133, \8359 );
nor \g451069/U$1 ( \13841 , \13839 , \13840 );
and \g454191/U$2 ( \13842 , \8313 , RIe16d100_2618);
and \g454191/U$3 ( \13843 , RIde941c0_312, \8323 );
nor \g454191/U$1 ( \13844 , \13842 , \13843 );
not \g449661/U$3 ( \13845 , \13844 );
not \g449661/U$4 ( \13846 , \8376 );
and \g449661/U$2 ( \13847 , \13845 , \13846 );
and \g449661/U$5 ( \13848 , \8340 , RIdeff6c8_1370);
nor \g449661/U$1 ( \13849 , \13847 , \13848 );
and \g451067/U$2 ( \13850 , \8378 , RIe158ef8_2389);
and \g451067/U$3 ( \13851 , RIdeb34f8_504, \8417 );
nor \g451067/U$1 ( \13852 , \13850 , \13851 );
nand \g447530/U$1 ( \13853 , \13838 , \13841 , \13849 , \13852 );
nor \g445811/U$1 ( \13854 , \13833 , \13834 , \13853 );
and \g451065/U$2 ( \13855 , \8335 , RIde7a108_185);
and \g451065/U$3 ( \13856 , RIdecf6f8_824, \8351 );
nor \g451065/U$1 ( \13857 , \13855 , \13856 );
and \g451066/U$2 ( \13858 , \8317 , RIdedaf30_955);
and \g451066/U$3 ( \13859 , RIdec6ff8_728, \8404 );
nor \g451066/U$1 ( \13860 , \13858 , \13859 );
and \g445010/U$2 ( \13861 , \13854 , \13857 , \13860 );
nor \g445010/U$1 ( \13862 , \13861 , \8651 );
or \g444184/U$1 ( \13863 , \13803 , \13832 , \13862 );
_DC \g2d1e/U$1 ( \13864 , \13863 , \8654 );
and \g447221/U$2 ( \13865 , \8785 , RIdeeb8f8_1144);
and \g447221/U$3 ( \13866 , RIdeee5f8_1176, \8787 );
nor \g447221/U$1 ( \13867 , \13865 , \13866 );
and \g446485/U$2 ( \13868 , RIdf188f8_1656, \8351 );
and \g446485/U$3 ( \13869 , RIdf15bf8_1624, \8383 );
and \g449496/U$2 ( \13870 , RIdf07af8_1464, \8414 );
and \g449496/U$3 ( \13871 , \8409 , RIdf0a7f8_1496);
and \g449496/U$4 ( \13872 , RIdef12f8_1208, \8326 );
nor \g449496/U$1 ( \13873 , \13870 , \13871 , \13872 );
and \g454070/U$2 ( \13874 , \8356 , RIdef6cf8_1272);
and \g454070/U$3 ( \13875 , RIdeff3f8_1368, \8359 );
nor \g454070/U$1 ( \13876 , \13874 , \13875 );
and \g455221/U$2 ( \13877 , \8313 , RIdef99f8_1304);
and \g455221/U$3 ( \13878 , RIdefc6f8_1336, \8323 );
nor \g455221/U$1 ( \13879 , \13877 , \13878 );
not \g450519/U$3 ( \13880 , \13879 );
not \g450519/U$4 ( \13881 , \8347 );
and \g450519/U$2 ( \13882 , \13880 , \13881 );
and \g450519/U$5 ( \13883 , \8340 , RIdef3ff8_1240);
nor \g450519/U$1 ( \13884 , \13882 , \13883 );
and \g454069/U$2 ( \13885 , \8378 , RIdf04df8_1432);
and \g454069/U$3 ( \13886 , RIdf0d4f8_1528, \8417 );
nor \g454069/U$1 ( \13887 , \13885 , \13886 );
nand \g447996/U$1 ( \13888 , \13873 , \13876 , \13884 , \13887 );
nor \g446485/U$1 ( \13889 , \13868 , \13869 , \13888 );
not \g444927/U$3 ( \13890 , \13889 );
not \g444927/U$4 ( \13891 , \8477 );
and \g444927/U$2 ( \13892 , \13890 , \13891 );
and \g446487/U$2 ( \13893 , RIfc4ff70_5932, \8373 );
and \g446487/U$3 ( \13894 , RIee24dd8_4878, \8383 );
and \g449499/U$2 ( \13895 , RIfe915c0_7998, \8412 );
and \g449499/U$3 ( \13896 , \8409 , RIdee4170_1059);
and \g449499/U$4 ( \13897 , RIfe91728_7999, \8326 );
nor \g449499/U$1 ( \13898 , \13895 , \13896 , \13897 );
and \g454078/U$2 ( \13899 , \8356 , RIee219d0_4841);
and \g454078/U$3 ( \13900 , RIfcd4810_7440, \8359 );
nor \g454078/U$1 ( \13901 , \13899 , \13900 );
and \g455404/U$2 ( \13902 , \8313 , RIfce1560_7586);
and \g455404/U$3 ( \13903 , RIee22948_4852, \8323 );
nor \g455404/U$1 ( \13904 , \13902 , \13903 );
not \g450521/U$3 ( \13905 , \13904 );
not \g450521/U$4 ( \13906 , \8347 );
and \g450521/U$2 ( \13907 , \13905 , \13906 );
and \g450521/U$5 ( \13908 , \8340 , RIdedac60_953);
nor \g450521/U$1 ( \13909 , \13907 , \13908 );
and \g454076/U$2 ( \13910 , \8378 , RIdedff58_1012);
and \g454076/U$3 ( \13911 , RIdee5ef8_1080, \8417 );
nor \g454076/U$1 ( \13912 , \13910 , \13911 );
nand \g447997/U$1 ( \13913 , \13898 , \13901 , \13909 , \13912 );
nor \g446487/U$1 ( \13914 , \13893 , \13894 , \13913 );
and \g454072/U$2 ( \13915 , \8335 , RIfe91890_8000);
and \g454072/U$3 ( \13916 , RIfc857d8_6541, \8351 );
nor \g454072/U$1 ( \13917 , \13915 , \13916 );
and \g454074/U$2 ( \13918 , \8319 , RIded64a8_902);
and \g454074/U$3 ( \13919 , RIfc50240_5934, \8404 );
nor \g454074/U$1 ( \13920 , \13918 , \13919 );
and \g445493/U$2 ( \13921 , \13914 , \13917 , \13920 );
nor \g445493/U$1 ( \13922 , \13921 , \8481 );
nor \g444927/U$1 ( \13923 , \13892 , \13922 );
and \g447222/U$2 ( \13924 , \9480 , RIdf101f8_1560);
and \g447222/U$3 ( \13925 , RIdf12ef8_1592, \9482 );
nor \g447222/U$1 ( \13926 , \13924 , \13925 );
nand \g444442/U$1 ( \13927 , \13867 , \13923 , \13926 );
and \g454091/U$2 ( \13928 , \8523 , RIfc9ea08_6827);
and \g454091/U$3 ( \13929 , RIdeb3228_502, \8486 );
nor \g454091/U$1 ( \13930 , \13928 , \13929 );
and \g446492/U$2 ( \13931 , RIdebb928_598, \8414 );
and \g446492/U$3 ( \13932 , RIdeb0528_470, \8356 );
and \g449504/U$2 ( \13933 , RIdebe628_630, \8407 );
and \g449504/U$3 ( \13934 , \8373 , RIee20bc0_4831);
and \g449504/U$4 ( \13935 , RIdec4028_694, \8383 );
nor \g449504/U$1 ( \13936 , \13933 , \13934 , \13935 );
and \g454098/U$2 ( \13937 , \8335 , RIdea0d30_374);
and \g454098/U$3 ( \13938 , RIee1e028_4800, \8340 );
nor \g454098/U$1 ( \13939 , \13937 , \13938 );
and \g454096/U$2 ( \13940 , \8404 , RIdec1328_662);
and \g454096/U$3 ( \13941 , RIdec6d28_726, \8351 );
nor \g454096/U$1 ( \13942 , \13940 , \13941 );
and \g455243/U$2 ( \13943 , \8313 , RIdea7630_406);
and \g455243/U$3 ( \13944 , RIdead828_438, \8323 );
nor \g455243/U$1 ( \13945 , \13943 , \13944 );
not \g455242/U$1 ( \13946 , \13945 );
and \g450526/U$2 ( \13947 , \13946 , \8316 );
and \g450526/U$3 ( \13948 , RIfcbaed8_7149, \8417 );
nor \g450526/U$1 ( \13949 , \13947 , \13948 );
nand \g448253/U$1 ( \13950 , \13936 , \13939 , \13942 , \13949 );
nor \g446492/U$1 ( \13951 , \13931 , \13932 , \13950 );
and \g454092/U$2 ( \13952 , \8378 , RIdeb8c28_566);
and \g454092/U$3 ( \13953 , RIfc412b8_5767, \8359 );
nor \g454092/U$1 ( \13954 , \13952 , \13953 );
nand \g445699/U$1 ( \13955 , \13930 , \13951 , \13954 );
and \g444731/U$2 ( \13956 , \13955 , \9702 );
and \g449501/U$2 ( \13957 , RIfe91458_7997, \8407 );
and \g449501/U$3 ( \13958 , \8373 , RIfcba668_7143);
and \g449501/U$4 ( \13959 , RIfc55538_5993, \8330 );
nor \g449501/U$1 ( \13960 , \13957 , \13958 , \13959 );
and \g454086/U$2 ( \13961 , \8335 , RIe169320_2574);
and \g454086/U$3 ( \13962 , RIee39418_5110, \8340 );
nor \g454086/U$1 ( \13963 , \13961 , \13962 );
and \g454084/U$2 ( \13964 , \8404 , RIfc4af48_5875);
and \g454084/U$3 ( \13965 , RIfcbac08_7147, \8351 );
nor \g454084/U$1 ( \13966 , \13964 , \13965 );
and \g455076/U$2 ( \13967 , \8313 , RIfc884d8_6573);
and \g455076/U$3 ( \13968 , RIe16ce30_2616, \8323 );
nor \g455076/U$1 ( \13969 , \13967 , \13968 );
not \g455075/U$1 ( \13970 , \13969 );
and \g450523/U$2 ( \13971 , \13970 , \8316 );
and \g450523/U$3 ( \13972 , RIfe912f0_7996, \8417 );
nor \g450523/U$1 ( \13973 , \13971 , \13972 );
nand \g448251/U$1 ( \13974 , \13960 , \13963 , \13966 , \13973 );
and \g444731/U$3 ( \13975 , \9700 , \13974 );
nor \g444731/U$1 ( \13976 , \13956 , \13975 );
and \g447226/U$2 ( \13977 , \12254 , RIde87ce0_252);
and \g447226/U$3 ( \13978 , RIde8be80_272, \12256 );
nor \g447226/U$1 ( \13979 , \13977 , \13978 );
and \g447225/U$2 ( \13980 , \12259 , RIfc88640_6574);
and \g447225/U$3 ( \13981 , RIfc85238_6537, \12261 );
nor \g447225/U$1 ( \13982 , \13980 , \13981 );
and \g447227/U$2 ( \13983 , \12264 , RIfcd5788_7451);
and \g447227/U$3 ( \13984 , RIfcda210_7504, \12266 );
nor \g447227/U$1 ( \13985 , \13983 , \13984 );
nand \g444548/U$1 ( \13986 , \13976 , \13979 , \13982 , \13985 );
and \g446480/U$2 ( \13987 , RIe158c28_2387, \8414 );
and \g446480/U$3 ( \13988 , RIe150528_2291, \8356 );
and \g449492/U$2 ( \13989 , RIe15e628_2451, \8407 );
and \g449492/U$3 ( \13990 , \8373 , RIfe90918_7989);
and \g449492/U$4 ( \13991 , RIe164028_2515, \8383 );
nor \g449492/U$1 ( \13992 , \13989 , \13990 , \13991 );
and \g454055/U$2 ( \13993 , \8335 , RIe147e28_2195);
and \g454055/U$3 ( \13994 , RIfcda378_7505, \8340 );
nor \g454055/U$1 ( \13995 , \13993 , \13994 );
and \g454054/U$2 ( \13996 , \8404 , RIe161328_2483);
and \g454054/U$3 ( \13997 , RIe166d28_2547, \8351 );
nor \g454054/U$1 ( \13998 , \13996 , \13997 );
and \g455258/U$2 ( \13999 , \8313 , RIe14ab28_2227);
and \g455258/U$3 ( \14000 , RIe14d828_2259, \8323 );
nor \g455258/U$1 ( \14001 , \13999 , \14000 );
not \g455257/U$1 ( \14002 , \14001 );
and \g450513/U$2 ( \14003 , \14002 , \8316 );
and \g450513/U$3 ( \14004 , RIee36880_5079, \8417 );
nor \g450513/U$1 ( \14005 , \14003 , \14004 );
nand \g448250/U$1 ( \14006 , \13992 , \13995 , \13998 , \14005 );
nor \g446480/U$1 ( \14007 , \13987 , \13988 , \14006 );
and \g454051/U$2 ( \14008 , \8378 , RIe155f28_2355);
and \g454051/U$3 ( \14009 , RIfe91188_7995, \8359 );
nor \g454051/U$1 ( \14010 , \14008 , \14009 );
and \g454050/U$2 ( \14011 , \8531 , RIfe91020_7994);
and \g454050/U$3 ( \14012 , RIe153228_2323, \8488 );
nor \g454050/U$1 ( \14013 , \14011 , \14012 );
and \g445488/U$2 ( \14014 , \14007 , \14010 , \14013 );
nor \g445488/U$1 ( \14015 , \14014 , \8368 );
and \g446482/U$2 ( \14016 , RIfcb99c0_7134, \8373 );
and \g446482/U$3 ( \14017 , RIfe90d50_7992, \8383 );
and \g449495/U$2 ( \14018 , RIdf346c0_1973, \8326 );
and \g449495/U$3 ( \14019 , \8531 , RIfc87dd0_6568);
and \g449495/U$4 ( \14020 , RIee30778_5010, \8488 );
nor \g449495/U$1 ( \14021 , \14018 , \14019 , \14020 );
and \g454064/U$2 ( \14022 , \8356 , RIee2e5b8_4986);
and \g454064/U$3 ( \14023 , RIfcec690_7712, \8359 );
nor \g454064/U$1 ( \14024 , \14022 , \14023 );
and \g455401/U$2 ( \14025 , \8313 , RIdf3e008_2082);
and \g455401/U$3 ( \14026 , RIfe90a80_7990, \8323 );
nor \g455401/U$1 ( \14027 , \14025 , \14026 );
not \g450518/U$3 ( \14028 , \14027 );
not \g450518/U$4 ( \14029 , \8376 );
and \g450518/U$2 ( \14030 , \14028 , \14029 );
and \g450518/U$5 ( \14031 , \8340 , RIdf36e20_2001);
nor \g450518/U$1 ( \14032 , \14030 , \14031 );
and \g454063/U$2 ( \14033 , \8378 , RIdf3bce0_2057);
and \g454063/U$3 ( \14034 , RIfe90be8_7991, \8417 );
nor \g454063/U$1 ( \14035 , \14033 , \14034 );
nand \g447995/U$1 ( \14036 , \14021 , \14024 , \14032 , \14035 );
nor \g446482/U$1 ( \14037 , \14016 , \14017 , \14036 );
and \g454059/U$2 ( \14038 , \8335 , RIdf30070_1923);
and \g454059/U$3 ( \14039 , RIfe90eb8_7993, \8351 );
nor \g454059/U$1 ( \14040 , \14038 , \14039 );
and \g454062/U$2 ( \14041 , \8319 , RIdf32668_1950);
and \g454062/U$3 ( \14042 , RIfc9c2a8_6799, \8404 );
nor \g454062/U$1 ( \14043 , \14041 , \14042 );
and \g445490/U$2 ( \14044 , \14037 , \14040 , \14043 );
nor \g445490/U$1 ( \14045 , \14044 , \8422 );
or \g444305/U$1 ( \14046 , \13927 , \13986 , \14015 , \14045 );
and \g446477/U$2 ( \14047 , RIfe904e0_7986, \8414 );
and \g446477/U$3 ( \14048 , RIfcb92b8_7129, \8531 );
and \g449489/U$2 ( \14049 , RIfe907b0_7988, \8407 );
and \g449489/U$3 ( \14050 , \8373 , RIee299c8_4932);
and \g449489/U$4 ( \14051 , RIee2aee0_4947, \8383 );
nor \g449489/U$1 ( \14052 , \14049 , \14050 , \14051 );
and \g454037/U$2 ( \14053 , \8335 , RIdf1a950_1679);
and \g454037/U$3 ( \14054 , RIfc86a20_6554, \8340 );
nor \g454037/U$1 ( \14055 , \14053 , \14054 );
and \g454036/U$2 ( \14056 , \8404 , RIee28618_4918);
and \g454036/U$3 ( \14057 , RIee2c998_4966, \8351 );
nor \g454036/U$1 ( \14058 , \14056 , \14057 );
and \g454954/U$2 ( \14059 , \8313 , RIfcb8fe8_7127);
and \g454954/U$3 ( \14060 , RIdf20e90_1751, \8323 );
nor \g454954/U$1 ( \14061 , \14059 , \14060 );
not \g454953/U$1 ( \14062 , \14061 );
and \g450510/U$2 ( \14063 , \14062 , \8316 );
and \g450510/U$3 ( \14064 , RIfe90378_7985, \8417 );
nor \g450510/U$1 ( \14065 , \14063 , \14064 );
nand \g448249/U$1 ( \14066 , \14052 , \14055 , \14058 , \14065 );
nor \g446477/U$1 ( \14067 , \14047 , \14048 , \14066 );
and \g454031/U$2 ( \14068 , \8356 , RIfc4ee90_5920);
and \g454031/U$3 ( \14069 , RIfc9d928_6815, \8359 );
nor \g454031/U$1 ( \14070 , \14068 , \14069 );
and \g454032/U$2 ( \14071 , \8378 , RIfe90648_7987);
and \g454032/U$3 ( \14072 , RIfc86048_6547, \8488 );
nor \g454032/U$1 ( \14073 , \14071 , \14072 );
and \g445483/U$2 ( \14074 , \14067 , \14070 , \14073 );
nor \g445483/U$1 ( \14075 , \14074 , \8621 );
and \g446479/U$2 ( \14076 , RIdecc728_790, \8371 );
and \g446479/U$3 ( \14077 , RIdecf428_822, \8383 );
and \g449490/U$2 ( \14078 , RIe16fb30_2648, \8414 );
and \g449490/U$3 ( \14079 , \8409 , RIde9a430_342);
and \g449490/U$4 ( \14080 , RIdee8bf8_1112, \8326 );
nor \g449490/U$1 ( \14081 , \14078 , \14079 , \14080 );
and \g454046/U$2 ( \14082 , \8356 , RIdf1ea00_1725);
and \g454046/U$3 ( \14083 , RIe145128_2163, \8359 );
nor \g454046/U$1 ( \14084 , \14082 , \14083 );
and \g455300/U$2 ( \14085 , \8313 , RIdf2e180_1901);
and \g455300/U$3 ( \14086 , RIdf39b20_2033, \8323 );
nor \g455300/U$1 ( \14087 , \14085 , \14086 );
not \g450511/U$3 ( \14088 , \14087 );
not \g450511/U$4 ( \14089 , \8347 );
and \g450511/U$2 ( \14090 , \14088 , \14089 );
and \g450511/U$5 ( \14091 , \8340 , RIdf020f8_1400);
nor \g450511/U$1 ( \14092 , \14090 , \14091 );
and \g454045/U$2 ( \14093 , \8378 , RIe15b928_2419);
and \g454045/U$3 ( \14094 , RIdeb5f28_534, \8417 );
nor \g454045/U$1 ( \14095 , \14093 , \14094 );
nand \g447993/U$1 ( \14096 , \14081 , \14084 , \14092 , \14095 );
nor \g446479/U$1 ( \14097 , \14076 , \14077 , \14096 );
and \g454039/U$2 ( \14098 , \8335 , RIde80378_215);
and \g454039/U$3 ( \14099 , RIded2128_854, \8351 );
nor \g454039/U$1 ( \14100 , \14098 , \14099 );
and \g454041/U$2 ( \14101 , \8319 , RIdedd960_985);
and \g454041/U$3 ( \14102 , RIdec9a28_758, \8404 );
nor \g454041/U$1 ( \14103 , \14101 , \14102 );
and \g445487/U$2 ( \14104 , \14097 , \14100 , \14103 );
nor \g445487/U$1 ( \14105 , \14104 , \8651 );
or \g444175/U$1 ( \14106 , \14046 , \14075 , \14105 );
_DC \g2da3/U$1 ( \14107 , \14106 , \8654 );
and \g446518/U$2 ( \14108 , \10230 , RIee2e450_4985);
and \g446518/U$3 ( \14109 , RIfcbe010_7184, \10232 );
nor \g446518/U$1 ( \14110 , \14108 , \14109 );
and \g445713/U$2 ( \14111 , RIe142428_2131, \8417 );
and \g445713/U$3 ( \14112 , RIe140100_2106, \8409 );
and \g448510/U$2 ( \14113 , RIee327d0_5033, \8373 );
and \g448510/U$3 ( \14114 , \8383 , RIee33a18_5046);
and \g448510/U$4 ( \14115 , RIee30610_5009, \8486 );
nor \g448510/U$1 ( \14116 , \14113 , \14114 , \14115 );
and \g450611/U$2 ( \14117 , \8335 , RIfec2d78_8337);
and \g450611/U$3 ( \14118 , RIfec2ee0_8338, \8340 );
nor \g450611/U$1 ( \14119 , \14117 , \14118 );
and \g450609/U$2 ( \14120 , \8404 , RIfcbcf30_7172);
and \g450609/U$3 ( \14121 , RIee34af8_5058, \8351 );
nor \g450609/U$1 ( \14122 , \14120 , \14121 );
and \g454176/U$2 ( \14123 , \8313 , RIfec2c10_8336);
and \g454176/U$3 ( \14124 , RIfec3048_8339, \8323 );
nor \g454176/U$1 ( \14125 , \14123 , \14124 );
not \g454175/U$1 ( \14126 , \14125 );
and \g449531/U$2 ( \14127 , \14126 , \8316 );
and \g449531/U$3 ( \14128 , RIfc731f0_6332, \8359 );
nor \g449531/U$1 ( \14129 , \14127 , \14128 );
nand \g448131/U$1 ( \14130 , \14116 , \14119 , \14122 , \14129 );
nor \g445713/U$1 ( \14131 , \14111 , \14112 , \14130 );
not \g444867/U$3 ( \14132 , \14131 );
not \g444867/U$4 ( \14133 , \8422 );
and \g444867/U$2 ( \14134 , \14132 , \14133 );
and \g445716/U$2 ( \14135 , RIe158ac0_2386, \8414 );
and \g445716/U$3 ( \14136 , RIfc54b60_5986, \8417 );
and \g448512/U$2 ( \14137 , RIee38338_5098, \8373 );
and \g448512/U$3 ( \14138 , \8383 , RIe163ec0_2514);
and \g448512/U$4 ( \14139 , RIe1530c0_2322, \8486 );
nor \g448512/U$1 ( \14140 , \14137 , \14138 , \14139 );
and \g450621/U$2 ( \14141 , \8335 , RIe147cc0_2194);
and \g450621/U$3 ( \14142 , RIfc9fdb8_6841, \8340 );
nor \g450621/U$1 ( \14143 , \14141 , \14142 );
and \g450620/U$2 ( \14144 , \8404 , RIe1611c0_2482);
and \g450620/U$3 ( \14145 , RIe166bc0_2546, \8351 );
nor \g450620/U$1 ( \14146 , \14144 , \14145 );
and \g454182/U$2 ( \14147 , \8313 , RIe14a9c0_2226);
and \g454182/U$3 ( \14148 , RIe14d6c0_2258, \8323 );
nor \g454182/U$1 ( \14149 , \14147 , \14148 );
not \g454181/U$1 ( \14150 , \14149 );
and \g449533/U$2 ( \14151 , \14150 , \8316 );
and \g449533/U$3 ( \14152 , RIee35a70_5069, \8359 );
nor \g449533/U$1 ( \14153 , \14151 , \14152 );
nand \g448132/U$1 ( \14154 , \14140 , \14143 , \14146 , \14153 );
nor \g445716/U$1 ( \14155 , \14135 , \14136 , \14154 );
and \g450617/U$2 ( \14156 , \8378 , RIe155dc0_2354);
and \g450617/U$3 ( \14157 , RIee357a0_5067, \8531 );
nor \g450617/U$1 ( \14158 , \14156 , \14157 );
and \g450618/U$2 ( \14159 , \8356 , RIe1503c0_2290);
and \g450618/U$3 ( \14160 , RIe15e4c0_2450, \8409 );
nor \g450618/U$1 ( \14161 , \14159 , \14160 );
and \g444939/U$2 ( \14162 , \14155 , \14158 , \14161 );
nor \g444939/U$1 ( \14163 , \14162 , \8368 );
nor \g444867/U$1 ( \14164 , \14134 , \14163 );
nor \g448407/U$1 ( \14165 , \8422 , \8437 );
and \g446519/U$2 ( \14166 , \14165 , RIdf3bb78_2056);
nor \g448438/U$1 ( \14167 , \8422 , \8413 );
and \g446519/U$3 ( \14168 , RIfea7280_8218, \14167 );
nor \g446519/U$1 ( \14169 , \14166 , \14168 );
nand \g444416/U$1 ( \14170 , \14110 , \14164 , \14169 );
and \g450633/U$2 ( \14171 , \8317 , RIdeee490_1175);
and \g450633/U$3 ( \14172 , RIdef1190_1207, \8326 );
nor \g450633/U$1 ( \14173 , \14171 , \14172 );
and \g445718/U$2 ( \14174 , RIdf12d90_1591, \8373 );
and \g445718/U$3 ( \14175 , RIdeeb790_1143, \8335 );
and \g448514/U$2 ( \14176 , RIdef9890_1303, \8531 );
and \g448514/U$3 ( \14177 , \8488 , RIdefc590_1335);
and \g448514/U$4 ( \14178 , RIdf15a90_1623, \8330 );
nor \g448514/U$1 ( \14179 , \14176 , \14177 , \14178 );
and \g450636/U$2 ( \14180 , \8356 , RIdef6b90_1271);
and \g450636/U$3 ( \14181 , RIdeff290_1367, \8359 );
nor \g450636/U$1 ( \14182 , \14180 , \14181 );
and \g454192/U$2 ( \14183 , \8313 , RIdf07990_1463);
and \g454192/U$3 ( \14184 , RIdf0a690_1495, \8323 );
nor \g454192/U$1 ( \14185 , \14183 , \14184 );
not \g449538/U$3 ( \14186 , \14185 );
not \g449538/U$4 ( \14187 , \8376 );
and \g449538/U$2 ( \14188 , \14186 , \14187 );
and \g449538/U$5 ( \14189 , \8351 , RIdf18790_1655);
nor \g449538/U$1 ( \14190 , \14188 , \14189 );
and \g450635/U$2 ( \14191 , \8378 , RIdf04c90_1431);
and \g450635/U$3 ( \14192 , RIdf0d390_1527, \8417 );
nor \g450635/U$1 ( \14193 , \14191 , \14192 );
nand \g447469/U$1 ( \14194 , \14179 , \14182 , \14190 , \14193 );
nor \g445718/U$1 ( \14195 , \14174 , \14175 , \14194 );
and \g450632/U$2 ( \14196 , \8340 , RIdef3e90_1239);
and \g450632/U$3 ( \14197 , RIdf10090_1559, \8404 );
nor \g450632/U$1 ( \14198 , \14196 , \14197 );
nand \g445510/U$1 ( \14199 , \14173 , \14195 , \14198 );
and \g444752/U$2 ( \14200 , \14199 , \8478 );
and \g448513/U$2 ( \14201 , RIfe8f568_7975, \8317 );
and \g448513/U$3 ( \14202 , \8324 , RIded87d0_927);
and \g448513/U$4 ( \14203 , RIfc534e0_5970, \8488 );
nor \g448513/U$1 ( \14204 , \14201 , \14202 , \14203 );
and \g450628/U$2 ( \14205 , \8335 , RIded42e8_878);
and \g450628/U$3 ( \14206 , RIfe8f6d0_7976, \8340 );
nor \g450628/U$1 ( \14207 , \14205 , \14206 );
and \g450627/U$2 ( \14208 , \8404 , RIfccf680_7382);
and \g450627/U$3 ( \14209 , RIee25be8_4888, \8351 );
nor \g450627/U$1 ( \14210 , \14208 , \14209 );
and \g454187/U$2 ( \14211 , \8313 , RIee23fc8_4868);
and \g454187/U$3 ( \14212 , RIfc6af28_6239, \8323 );
nor \g454187/U$1 ( \14213 , \14211 , \14212 );
not \g449534/U$3 ( \14214 , \14213 );
not \g449534/U$4 ( \14215 , \8328 );
and \g449534/U$2 ( \14216 , \14214 , \14215 );
and \g449534/U$5 ( \14217 , \8359 , RIfc6b090_6240);
nor \g449534/U$1 ( \14218 , \14216 , \14217 );
nand \g447468/U$1 ( \14219 , \14204 , \14207 , \14210 , \14218 );
and \g444752/U$3 ( \14220 , \8482 , \14219 );
nor \g444752/U$1 ( \14221 , \14200 , \14220 );
and \g446523/U$2 ( \14222 , \8964 , RIdee4008_1058);
and \g446523/U$3 ( \14223 , RIdee5d90_1079, \8966 );
nor \g446523/U$1 ( \14224 , \14222 , \14223 );
and \g446524/U$2 ( \14225 , \8521 , RIfc66770_6188);
and \g446524/U$3 ( \14226 , RIfca5920_6906, \8525 );
nor \g446524/U$1 ( \14227 , \14225 , \14226 );
and \g446525/U$2 ( \14228 , \8974 , RIdedfdf0_1011);
and \g446525/U$3 ( \14229 , RIdee1ce0_1033, \8976 );
nor \g446525/U$1 ( \14230 , \14228 , \14229 );
nand \g444446/U$1 ( \14231 , \14221 , \14224 , \14227 , \14230 );
and \g445711/U$2 ( \14232 , RIee29860_4931, \8373 );
and \g445711/U$3 ( \14233 , RIdf1a7e8_1678, \8335 );
and \g448506/U$2 ( \14234 , RIdf23a28_1782, \8531 );
and \g448506/U$3 ( \14235 , \8488 , RIfc53648_5971);
and \g448506/U$4 ( \14236 , RIfcb4830_7076, \8383 );
nor \g448506/U$1 ( \14237 , \14234 , \14235 , \14236 );
and \g450598/U$2 ( \14238 , \8356 , RIfc823d0_6504);
and \g450598/U$3 ( \14239 , RIfcc9de8_7319, \8359 );
nor \g450598/U$1 ( \14240 , \14238 , \14239 );
and \g454169/U$2 ( \14241 , \8313 , RIdf27268_1822);
and \g454169/U$3 ( \14242 , RIdf29590_1847, \8323 );
nor \g454169/U$1 ( \14243 , \14241 , \14242 );
not \g449527/U$3 ( \14244 , \14243 );
not \g449527/U$4 ( \14245 , \8376 );
and \g449527/U$2 ( \14246 , \14244 , \14245 );
and \g449527/U$5 ( \14247 , \8351 , RIfcb46c8_7075);
nor \g449527/U$1 ( \14248 , \14246 , \14247 );
and \g450597/U$2 ( \14249 , \8378 , RIdf25648_1802);
and \g450597/U$3 ( \14250 , RIdf2b480_1869, \8417 );
nor \g450597/U$1 ( \14251 , \14249 , \14250 );
nand \g447462/U$1 ( \14252 , \14237 , \14240 , \14248 , \14251 );
nor \g445711/U$1 ( \14253 , \14232 , \14233 , \14252 );
and \g450592/U$2 ( \14254 , \8340 , RIdf223a8_1766);
and \g450592/U$3 ( \14255 , RIfcb88e0_7122, \8404 );
nor \g450592/U$1 ( \14256 , \14254 , \14255 );
and \g450594/U$2 ( \14257 , \8319 , RIdf1bd00_1693);
and \g450594/U$3 ( \14258 , RIdf20d28_1750, \8324 );
nor \g450594/U$1 ( \14259 , \14257 , \14258 );
and \g444936/U$2 ( \14260 , \14253 , \14256 , \14259 );
nor \g444936/U$1 ( \14261 , \14260 , \8621 );
and \g445712/U$2 ( \14262 , RIde9a0e8_341, \8407 );
and \g445712/U$3 ( \14263 , RIe15b7c0_2418, \8378 );
and \g448508/U$2 ( \14264 , RIdedd7f8_984, \8319 );
and \g448508/U$3 ( \14265 , \8326 , RIdee8a90_1111);
and \g448508/U$4 ( \14266 , RIdf399b8_2032, \8488 );
nor \g448508/U$1 ( \14267 , \14264 , \14265 , \14266 );
and \g450605/U$2 ( \14268 , \8335 , RIde80030_214);
and \g450605/U$3 ( \14269 , RIdf01f90_1399, \8340 );
nor \g450605/U$1 ( \14270 , \14268 , \14269 );
and \g450603/U$2 ( \14271 , \8404 , RIdec98c0_757);
and \g450603/U$3 ( \14272 , RIded1fc0_853, \8351 );
nor \g450603/U$1 ( \14273 , \14271 , \14272 );
and \g454172/U$2 ( \14274 , \8313 , RIdecc5c0_789);
and \g454172/U$3 ( \14275 , RIdecf2c0_821, \8323 );
nor \g454172/U$1 ( \14276 , \14274 , \14275 );
not \g449529/U$3 ( \14277 , \14276 );
not \g449529/U$4 ( \14278 , \8328 );
and \g449529/U$2 ( \14279 , \14277 , \14278 );
and \g449529/U$5 ( \14280 , \8359 , RIe144fc0_2162);
nor \g449529/U$1 ( \14281 , \14279 , \14280 );
nand \g447463/U$1 ( \14282 , \14267 , \14270 , \14273 , \14281 );
nor \g445712/U$1 ( \14283 , \14262 , \14263 , \14282 );
and \g450602/U$2 ( \14284 , \8356 , RIdf1e898_1724);
and \g450602/U$3 ( \14285 , RIdeb5dc0_533, \8417 );
nor \g450602/U$1 ( \14286 , \14284 , \14285 );
and \g450601/U$2 ( \14287 , \8531 , RIdf2e018_1900);
and \g450601/U$3 ( \14288 , RIe16f9c8_2647, \8412 );
nor \g450601/U$1 ( \14289 , \14287 , \14288 );
and \g444938/U$2 ( \14290 , \14283 , \14286 , \14289 );
nor \g444938/U$1 ( \14291 , \14290 , \8651 );
or \g444290/U$1 ( \14292 , \14170 , \14231 , \14261 , \14291 );
and \g445706/U$2 ( \14293 , RIfc5d800_6086, \8371 );
and \g445706/U$3 ( \14294 , RIe1691b8_2573, \8335 );
and \g448500/U$2 ( \14295 , RIfea73e8_8219, \8412 );
and \g448500/U$3 ( \14296 , \8409 , RIfea7820_8222);
and \g448500/U$4 ( \14297 , RIfcd16d8_7405, \8383 );
nor \g448500/U$1 ( \14298 , \14295 , \14296 , \14297 );
and \g450578/U$2 ( \14299 , \8356 , RIfc7a108_6411);
and \g450578/U$3 ( \14300 , RIde837f8_231, \8359 );
nor \g450578/U$1 ( \14301 , \14299 , \14300 );
and \g454158/U$2 ( \14302 , \8313 , RIfcc7ef8_7297);
and \g454158/U$3 ( \14303 , RIfc7bd28_6431, \8323 );
nor \g454158/U$1 ( \14304 , \14302 , \14303 );
not \g449523/U$3 ( \14305 , \14304 );
not \g449523/U$4 ( \14306 , \8347 );
and \g449523/U$2 ( \14307 , \14305 , \14306 );
and \g449523/U$5 ( \14308 , \8351 , RIfcb2508_7051);
nor \g449523/U$1 ( \14309 , \14307 , \14308 );
and \g450577/U$2 ( \14310 , \8378 , RIde87998_251);
and \g450577/U$3 ( \14311 , RIde93b30_310, \8417 );
nor \g450577/U$1 ( \14312 , \14310 , \14311 );
nand \g447458/U$1 ( \14313 , \14298 , \14301 , \14309 , \14312 );
nor \g445706/U$1 ( \14314 , \14293 , \14294 , \14313 );
and \g450575/U$2 ( \14315 , \8340 , RIfc7a6a8_6415);
and \g450575/U$3 ( \14316 , RIfc63d40_6158, \8404 );
nor \g450575/U$1 ( \14317 , \14315 , \14316 );
and \g450576/U$2 ( \14318 , \8319 , RIe16a838_2589);
and \g450576/U$3 ( \14319 , RIe16ccc8_2615, \8326 );
nor \g450576/U$1 ( \14320 , \14318 , \14319 );
and \g444933/U$2 ( \14321 , \14314 , \14317 , \14320 );
nor \g444933/U$1 ( \14322 , \14321 , \8558 );
and \g445708/U$2 ( \14323 , RIee1f978_4818, \8417 );
and \g445708/U$3 ( \14324 , RIdeb03c0_469, \8356 );
and \g448504/U$2 ( \14325 , RIdea72e8_405, \8317 );
and \g448504/U$3 ( \14326 , \8326 , RIdead6c0_437);
and \g448504/U$4 ( \14327 , RIdeb30c0_501, \8486 );
nor \g448504/U$1 ( \14328 , \14325 , \14326 , \14327 );
and \g450588/U$2 ( \14329 , \8335 , RIdea09e8_373);
and \g450588/U$3 ( \14330 , RIfc5e4a8_6095, \8340 );
nor \g450588/U$1 ( \14331 , \14329 , \14330 );
and \g450587/U$2 ( \14332 , \8404 , RIdec11c0_661);
and \g450587/U$3 ( \14333 , RIdec6bc0_725, \8351 );
nor \g450587/U$1 ( \14334 , \14332 , \14333 );
and \g454664/U$2 ( \14335 , \8313 , RIee20a58_4830);
and \g454664/U$3 ( \14336 , RIdec3ec0_693, \8323 );
nor \g454664/U$1 ( \14337 , \14335 , \14336 );
not \g449525/U$3 ( \14338 , \14337 );
not \g449525/U$4 ( \14339 , \8328 );
and \g449525/U$2 ( \14340 , \14338 , \14339 );
and \g449525/U$5 ( \14341 , \8359 , RIee1efa0_4811);
nor \g449525/U$1 ( \14342 , \14340 , \14341 );
nand \g447460/U$1 ( \14343 , \14328 , \14331 , \14334 , \14342 );
nor \g445708/U$1 ( \14344 , \14323 , \14324 , \14343 );
and \g450585/U$2 ( \14345 , \8378 , RIdeb8ac0_565);
and \g450585/U$3 ( \14346 , RIfcb04b0_7028, \8531 );
nor \g450585/U$1 ( \14347 , \14345 , \14346 );
and \g450584/U$2 ( \14348 , \8414 , RIdebb7c0_597);
and \g450584/U$3 ( \14349 , RIdebe4c0_629, \8409 );
nor \g450584/U$1 ( \14350 , \14348 , \14349 );
and \g444934/U$2 ( \14351 , \14344 , \14347 , \14350 );
nor \g444934/U$1 ( \14352 , \14351 , \8589 );
or \g444232/U$1 ( \14353 , \14292 , \14322 , \14352 );
_DC \g2e28/U$1 ( \14354 , \14353 , \8654 );
and \g449373/U$2 ( \14355 , RIe14a858_2225, \8319 );
and \g449373/U$3 ( \14356 , \8326 , RIe14d558_2257);
and \g449373/U$4 ( \14357 , RIe15e358_2449, \8407 );
nor \g449373/U$1 ( \14358 , \14355 , \14356 , \14357 );
and \g453619/U$2 ( \14359 , \8335 , RIe147b58_2193);
and \g453619/U$3 ( \14360 , RIfcb9b28_7135, \8340 );
nor \g453619/U$1 ( \14361 , \14359 , \14360 );
and \g453617/U$2 ( \14362 , \8404 , RIe161058_2481);
and \g453617/U$3 ( \14363 , RIe166a58_2545, \8351 );
nor \g453617/U$1 ( \14364 , \14362 , \14363 );
and \g455150/U$2 ( \14365 , \8313 , RIfec3cf0_8348);
and \g455150/U$3 ( \14366 , RIe163d58_2513, \8323 );
nor \g455150/U$1 ( \14367 , \14365 , \14366 );
not \g450395/U$3 ( \14368 , \14367 );
not \g450395/U$4 ( \14369 , \8328 );
and \g450395/U$2 ( \14370 , \14368 , \14369 );
and \g450395/U$5 ( \14371 , \8417 , RIfcd54b8_7449);
nor \g450395/U$1 ( \14372 , \14370 , \14371 );
nand \g447931/U$1 ( \14373 , \14358 , \14361 , \14364 , \14372 );
and \g444802/U$2 ( \14374 , \14373 , \8369 );
and \g446386/U$2 ( \14375 , RIfc9a0e8_6775, \8373 );
and \g446386/U$3 ( \14376 , RIfc553d0_5992, \8383 );
and \g449377/U$2 ( \14377 , RIfec3fc0_8350, \8326 );
and \g449377/U$3 ( \14378 , \8531 , RIfcc51f8_7265);
and \g449377/U$4 ( \14379 , RIee304a8_5008, \8486 );
nor \g449377/U$1 ( \14380 , \14377 , \14378 , \14379 );
and \g453624/U$2 ( \14381 , \8356 , RIee2e2e8_4984);
and \g453624/U$3 ( \14382 , RIfc87128_6559, \8359 );
nor \g453624/U$1 ( \14383 , \14381 , \14382 );
and \g455146/U$2 ( \14384 , \8313 , RIdf3dea0_2081);
and \g455146/U$3 ( \14385 , RIe13ff98_2105, \8323 );
nor \g455146/U$1 ( \14386 , \14384 , \14385 );
not \g450397/U$3 ( \14387 , \14386 );
not \g450397/U$4 ( \14388 , \8376 );
and \g450397/U$2 ( \14389 , \14387 , \14388 );
and \g450397/U$5 ( \14390 , \8340 , RIdf36cb8_2000);
nor \g450397/U$1 ( \14391 , \14389 , \14390 );
and \g453623/U$2 ( \14392 , \8378 , RIdf3ba10_2055);
and \g453623/U$3 ( \14393 , RIe1422c0_2130, \8417 );
nor \g453623/U$1 ( \14394 , \14392 , \14393 );
nand \g447932/U$1 ( \14395 , \14380 , \14383 , \14391 , \14394 );
nor \g446386/U$1 ( \14396 , \14375 , \14376 , \14395 );
and \g453621/U$2 ( \14397 , \8335 , RIfec3e58_8349);
and \g453621/U$3 ( \14398 , RIfcdb2f0_7516, \8351 );
nor \g453621/U$1 ( \14399 , \14397 , \14398 );
and \g453622/U$2 ( \14400 , \8319 , RIdf32500_1949);
and \g453622/U$3 ( \14401 , RIfcbd908_7179, \8404 );
nor \g453622/U$1 ( \14402 , \14400 , \14401 );
and \g445421/U$2 ( \14403 , \14396 , \14399 , \14402 );
nor \g445421/U$1 ( \14404 , \14403 , \8422 );
nor \g444802/U$1 ( \14405 , \14374 , \14404 );
and \g447136/U$2 ( \14406 , \8438 , RIe155c58_2353);
and \g447136/U$3 ( \14407 , RIe158958_2385, \8440 );
nor \g447136/U$1 ( \14408 , \14406 , \14407 );
and \g447135/U$2 ( \14409 , \12506 , RIe152f58_2321);
and \g447135/U$3 ( \14410 , RIfe9ba48_8115, \12508 );
nor \g447135/U$1 ( \14411 , \14409 , \14410 );
and \g447137/U$2 ( \14412 , \8717 , RIe150258_2289);
and \g447137/U$3 ( \14413 , RIfec4128_8351, \8719 );
nor \g447137/U$1 ( \14414 , \14412 , \14413 );
nand \g444534/U$1 ( \14415 , \14405 , \14408 , \14411 , \14414 );
and \g453607/U$2 ( \14416 , \8319 , RIdeee328_1174);
and \g453607/U$3 ( \14417 , RIdf0ff28_1558, \8404 );
nor \g453607/U$1 ( \14418 , \14416 , \14417 );
and \g446383/U$2 ( \14419 , RIdf12c28_1590, \8373 );
and \g446383/U$3 ( \14420 , RIdf15928_1622, \8383 );
and \g449372/U$2 ( \14421 , RIdf07828_1462, \8414 );
and \g449372/U$3 ( \14422 , \8407 , RIdf0a528_1494);
and \g449372/U$4 ( \14423 , RIdef1028_1206, \8326 );
nor \g449372/U$1 ( \14424 , \14421 , \14422 , \14423 );
and \g453610/U$2 ( \14425 , \8356 , RIdef6a28_1270);
and \g453610/U$3 ( \14426 , RIdeff128_1366, \8359 );
nor \g453610/U$1 ( \14427 , \14425 , \14426 );
and \g454266/U$2 ( \14428 , \8313 , RIdef9728_1302);
and \g454266/U$3 ( \14429 , RIdefc428_1334, \8323 );
nor \g454266/U$1 ( \14430 , \14428 , \14429 );
not \g450392/U$3 ( \14431 , \14430 );
not \g450392/U$4 ( \14432 , \8347 );
and \g450392/U$2 ( \14433 , \14431 , \14432 );
and \g450392/U$5 ( \14434 , \8340 , RIdef3d28_1238);
nor \g450392/U$1 ( \14435 , \14433 , \14434 );
and \g453608/U$2 ( \14436 , \8378 , RIdf04b28_1430);
and \g453608/U$3 ( \14437 , RIdf0d228_1526, \8417 );
nor \g453608/U$1 ( \14438 , \14436 , \14437 );
nand \g447928/U$1 ( \14439 , \14424 , \14427 , \14435 , \14438 );
nor \g446383/U$1 ( \14440 , \14419 , \14420 , \14439 );
and \g453605/U$2 ( \14441 , \8335 , RIdeeb628_1142);
and \g453605/U$3 ( \14442 , RIdf18628_1654, \8351 );
nor \g453605/U$1 ( \14443 , \14441 , \14442 );
nand \g445676/U$1 ( \14444 , \14418 , \14440 , \14443 );
and \g444801/U$2 ( \14445 , \14444 , \8478 );
and \g449370/U$2 ( \14446 , RIfeaa3b8_8253, \8324 );
and \g449370/U$3 ( \14447 , \8531 , RIdf238c0_1781);
and \g449370/U$4 ( \14448 , RIfc86b88_6555, \8488 );
nor \g449370/U$1 ( \14449 , \14446 , \14447 , \14448 );
and \g453600/U$2 ( \14450 , \8356 , RIfc75ab8_6361);
and \g453600/U$3 ( \14451 , RIfcb7c38_7113, \8359 );
nor \g453600/U$1 ( \14452 , \14450 , \14451 );
and \g454326/U$2 ( \14453 , \8313 , RIfe9b778_8113);
and \g454326/U$3 ( \14454 , RIfe9b610_8112, \8323 );
nor \g454326/U$1 ( \14455 , \14453 , \14454 );
not \g450390/U$3 ( \14456 , \14455 );
not \g450390/U$4 ( \14457 , \8376 );
and \g450390/U$2 ( \14458 , \14456 , \14457 );
and \g450390/U$5 ( \14459 , \8340 , RIdf22240_1765);
nor \g450390/U$1 ( \14460 , \14458 , \14459 );
and \g453599/U$2 ( \14461 , \8378 , RIfe9b4a8_8111);
and \g453599/U$3 ( \14462 , RIfe9b8e0_8114, \8417 );
nor \g453599/U$1 ( \14463 , \14461 , \14462 );
nand \g447927/U$1 ( \14464 , \14449 , \14452 , \14460 , \14463 );
and \g444801/U$3 ( \14465 , \8752 , \14464 );
nor \g444801/U$1 ( \14466 , \14445 , \14465 );
and \g447133/U$2 ( \14467 , \11762 , RIdf1a680_1677);
and \g447133/U$3 ( \14468 , RIdf1bb98_1692, \11764 );
nor \g447133/U$1 ( \14469 , \14467 , \14468 );
and \g447132/U$2 ( \14470 , \11767 , RIee2ad78_4946);
and \g447132/U$3 ( \14471 , RIee2c830_4965, \11769 );
nor \g447132/U$1 ( \14472 , \14470 , \14471 );
and \g447134/U$2 ( \14473 , \11511 , RIee284b0_4917);
and \g447134/U$3 ( \14474 , RIee296f8_4930, \11513 );
nor \g447134/U$1 ( \14475 , \14473 , \14474 );
nand \g444533/U$1 ( \14476 , \14466 , \14469 , \14472 , \14475 );
and \g446378/U$2 ( \14477 , RIdeb8958_564, \8378 );
and \g446378/U$3 ( \14478 , RIfcb96f0_7132, \8359 );
and \g449366/U$2 ( \14479 , RIdebe358_628, \8407 );
and \g449366/U$3 ( \14480 , \8371 , RIfc723e0_6322);
and \g449366/U$4 ( \14481 , RIdec3d58_692, \8383 );
nor \g449366/U$1 ( \14482 , \14479 , \14480 , \14481 );
and \g453585/U$2 ( \14483 , \8335 , RIdea06a0_372);
and \g453585/U$3 ( \14484 , RIfc9b498_6789, \8340 );
nor \g453585/U$1 ( \14485 , \14483 , \14484 );
and \g453583/U$2 ( \14486 , \8404 , RIdec1058_660);
and \g453583/U$3 ( \14487 , RIdec6a58_724, \8351 );
nor \g453583/U$1 ( \14488 , \14486 , \14487 );
and \g454462/U$2 ( \14489 , \8313 , RIdea6fa0_404);
and \g454462/U$3 ( \14490 , RIdead558_436, \8323 );
nor \g454462/U$1 ( \14491 , \14489 , \14490 );
not \g454461/U$1 ( \14492 , \14491 );
and \g450386/U$2 ( \14493 , \14492 , \8316 );
and \g450386/U$3 ( \14494 , RIfc59fc0_6046, \8417 );
nor \g450386/U$1 ( \14495 , \14493 , \14494 );
nand \g448233/U$1 ( \14496 , \14482 , \14485 , \14488 , \14495 );
nor \g446378/U$1 ( \14497 , \14477 , \14478 , \14496 );
and \g453578/U$2 ( \14498 , \8356 , RIdeb0258_468);
and \g453578/U$3 ( \14499 , RIdebb658_596, \8414 );
nor \g453578/U$1 ( \14500 , \14498 , \14499 );
and \g453577/U$2 ( \14501 , \8531 , RIfce1c68_7591);
and \g453577/U$3 ( \14502 , RIdeb2f58_500, \8488 );
nor \g453577/U$1 ( \14503 , \14501 , \14502 );
and \g445415/U$2 ( \14504 , \14497 , \14500 , \14503 );
nor \g445415/U$1 ( \14505 , \14504 , \8589 );
and \g446380/U$2 ( \14506 , RIde87650_250, \8378 );
and \g446380/U$3 ( \14507 , RIde834b0_230, \8359 );
and \g449368/U$2 ( \14508 , RIe16a6d0_2588, \8319 );
and \g449368/U$3 ( \14509 , \8326 , RIe16cb60_2614);
and \g449368/U$4 ( \14510 , RIde8f990_290, \8407 );
nor \g449368/U$1 ( \14511 , \14508 , \14509 , \14510 );
and \g453592/U$2 ( \14512 , \8335 , RIe169050_2572);
and \g453592/U$3 ( \14513 , RIee392b0_5109, \8340 );
nor \g453592/U$1 ( \14514 , \14512 , \14513 );
and \g453590/U$2 ( \14515 , \8404 , RIfcd3e38_7433);
and \g453590/U$3 ( \14516 , RIfc81458_6493, \8351 );
nor \g453590/U$1 ( \14517 , \14515 , \14516 );
and \g455161/U$2 ( \14518 , \8313 , RIfc4e620_5914);
and \g455161/U$3 ( \14519 , RIfc83780_6518, \8323 );
nor \g455161/U$1 ( \14520 , \14518 , \14519 );
not \g450388/U$3 ( \14521 , \14520 );
not \g450388/U$4 ( \14522 , \8328 );
and \g450388/U$2 ( \14523 , \14521 , \14522 );
and \g450388/U$5 ( \14524 , \8417 , RIde937e8_309);
nor \g450388/U$1 ( \14525 , \14523 , \14524 );
nand \g447926/U$1 ( \14526 , \14511 , \14514 , \14517 , \14525 );
nor \g446380/U$1 ( \14527 , \14506 , \14507 , \14526 );
and \g453587/U$2 ( \14528 , \8356 , RIfc6c710_6256);
and \g453587/U$3 ( \14529 , RIde8bb38_271, \8414 );
nor \g453587/U$1 ( \14530 , \14528 , \14529 );
and \g453586/U$2 ( \14531 , \8531 , RIfc65960_6178);
and \g453586/U$3 ( \14532 , RIfc42c80_5782, \8488 );
nor \g453586/U$1 ( \14533 , \14531 , \14532 );
and \g445416/U$2 ( \14534 , \14527 , \14530 , \14533 );
nor \g445416/U$1 ( \14535 , \14534 , \8558 );
or \g444410/U$1 ( \14536 , \14415 , \14476 , \14505 , \14535 );
and \g446375/U$2 ( \14537 , RIdeb5c58_532, \8417 );
and \g446375/U$3 ( \14538 , RIdec9758_756, \8404 );
and \g449360/U$2 ( \14539 , RIdf2deb0_1899, \8531 );
and \g449360/U$3 ( \14540 , \8488 , RIdf39850_2031);
and \g449360/U$4 ( \14541 , RIdecf158_820, \8383 );
nor \g449360/U$1 ( \14542 , \14539 , \14540 , \14541 );
and \g453567/U$2 ( \14543 , \8335 , RIde7fce8_213);
and \g453567/U$3 ( \14544 , RIdf01e28_1398, \8340 );
nor \g453567/U$1 ( \14545 , \14543 , \14544 );
and \g454633/U$2 ( \14546 , \8313 , RIdedd690_983);
and \g454633/U$3 ( \14547 , RIdee8928_1110, \8323 );
nor \g454633/U$1 ( \14548 , \14546 , \14547 );
not \g454632/U$1 ( \14549 , \14548 );
and \g450380/U$2 ( \14550 , \14549 , \8316 );
and \g450380/U$3 ( \14551 , RIded1e58_852, \8351 );
nor \g450380/U$1 ( \14552 , \14550 , \14551 );
and \g453566/U$2 ( \14553 , \8356 , RIdf1e730_1723);
and \g453566/U$3 ( \14554 , RIe144e58_2161, \8359 );
nor \g453566/U$1 ( \14555 , \14553 , \14554 );
nand \g448232/U$1 ( \14556 , \14542 , \14545 , \14552 , \14555 );
nor \g446375/U$1 ( \14557 , \14537 , \14538 , \14556 );
and \g453563/U$2 ( \14558 , \8378 , RIe15b658_2417);
and \g453563/U$3 ( \14559 , RIdecc458_788, \8373 );
nor \g453563/U$1 ( \14560 , \14558 , \14559 );
and \g453562/U$2 ( \14561 , \8414 , RIe16f860_2646);
and \g453562/U$3 ( \14562 , RIde99da0_340, \8409 );
nor \g453562/U$1 ( \14563 , \14561 , \14562 );
and \g445410/U$2 ( \14564 , \14557 , \14560 , \14563 );
nor \g445410/U$1 ( \14565 , \14564 , \8651 );
and \g446376/U$2 ( \14566 , RIdee1b78_1032, \8414 );
and \g446376/U$3 ( \14567 , RIee21868_4840, \8356 );
and \g449363/U$2 ( \14568 , RIded6340_901, \8319 );
and \g449363/U$3 ( \14569 , \8324 , RIded8668_926);
and \g449363/U$4 ( \14570 , RIdee3ea0_1057, \8409 );
nor \g449363/U$1 ( \14571 , \14568 , \14569 , \14570 );
and \g453574/U$2 ( \14572 , \8335 , RIded4180_877);
and \g453574/U$3 ( \14573 , RIdedaaf8_952, \8340 );
nor \g453574/U$1 ( \14574 , \14572 , \14573 );
and \g453573/U$2 ( \14575 , \8404 , RIfccc110_7344);
and \g453573/U$3 ( \14576 , RIee25a80_4887, \8351 );
nor \g453573/U$1 ( \14577 , \14575 , \14576 );
and \g454535/U$2 ( \14578 , \8313 , RIfcddd20_7546);
and \g454535/U$3 ( \14579 , RIee24c70_4877, \8323 );
nor \g454535/U$1 ( \14580 , \14578 , \14579 );
not \g450385/U$3 ( \14581 , \14580 );
not \g450385/U$4 ( \14582 , \8328 );
and \g450385/U$2 ( \14583 , \14581 , \14582 );
and \g450385/U$5 ( \14584 , \8417 , RIdee5c28_1078);
nor \g450385/U$1 ( \14585 , \14583 , \14584 );
nand \g447923/U$1 ( \14586 , \14571 , \14574 , \14577 , \14585 );
nor \g446376/U$1 ( \14587 , \14566 , \14567 , \14586 );
and \g453572/U$2 ( \14588 , \8378 , RIdedfc88_1010);
and \g453572/U$3 ( \14589 , RIfc6a6b8_6233, \8359 );
nor \g453572/U$1 ( \14590 , \14588 , \14589 );
and \g453571/U$2 ( \14591 , \8531 , RIfc88be0_6578);
and \g453571/U$3 ( \14592 , RIee227e0_4851, \8486 );
nor \g453571/U$1 ( \14593 , \14591 , \14592 );
and \g445411/U$2 ( \14594 , \14587 , \14590 , \14593 );
nor \g445411/U$1 ( \14595 , \14594 , \8481 );
or \g444173/U$1 ( \14596 , \14536 , \14565 , \14595 );
_DC \g2ead/U$1 ( \14597 , \14596 , \8654 );
and \g453739/U$2 ( \14598 , \8414 , RIde8b7f0_270);
and \g453739/U$3 ( \14599 , RIfe9b1d8_8109, \8407 );
nor \g453739/U$1 ( \14600 , \14598 , \14599 );
and \g446412/U$2 ( \14601 , RIde934a0_308, \8417 );
and \g446412/U$3 ( \14602 , RIee1b058_4766, \8404 );
and \g449408/U$2 ( \14603 , RIfcb27d8_7053, \8319 );
and \g449408/U$3 ( \14604 , \8326 , RIe16c9f8_2613);
and \g449408/U$4 ( \14605 , RIee1c6d8_4782, \8383 );
nor \g449408/U$1 ( \14606 , \14603 , \14604 , \14605 );
and \g453744/U$2 ( \14607 , \8335 , RIe168ee8_2571);
and \g453744/U$3 ( \14608 , RIfc511b8_5945, \8340 );
nor \g453744/U$1 ( \14609 , \14607 , \14608 );
and \g454595/U$2 ( \14610 , \8313 , RIfcd3a00_7430);
and \g454595/U$3 ( \14611 , RIfcb2238_7049, \8323 );
nor \g454595/U$1 ( \14612 , \14610 , \14611 );
not \g450428/U$3 ( \14613 , \14612 );
not \g450428/U$4 ( \14614 , \8347 );
and \g450428/U$2 ( \14615 , \14613 , \14614 );
and \g450428/U$5 ( \14616 , \8351 , RIfce5070_7628);
nor \g450428/U$1 ( \14617 , \14615 , \14616 );
and \g453742/U$2 ( \14618 , \8356 , RIfcdb020_7514);
and \g453742/U$3 ( \14619 , RIfc6b798_6245, \8359 );
nor \g453742/U$1 ( \14620 , \14618 , \14619 );
nand \g447952/U$1 ( \14621 , \14606 , \14609 , \14617 , \14620 );
nor \g446412/U$1 ( \14622 , \14601 , \14602 , \14621 );
and \g453741/U$2 ( \14623 , \8378 , RIfe9b340_8110);
and \g453741/U$3 ( \14624 , RIfce70c8_7651, \8373 );
nor \g453741/U$1 ( \14625 , \14623 , \14624 );
nand \g445682/U$1 ( \14626 , \14600 , \14622 , \14625 );
and \g444747/U$2 ( \14627 , \14626 , \9700 );
and \g449406/U$2 ( \14628 , RIfcc6710_7280, \8523 );
and \g449406/U$3 ( \14629 , \8486 , RIdeb2df0_499);
and \g449406/U$4 ( \14630 , RIdec3bf0_691, \8330 );
nor \g449406/U$1 ( \14631 , \14628 , \14629 , \14630 );
and \g453738/U$2 ( \14632 , \8335 , RIdea0358_371);
and \g453738/U$3 ( \14633 , RIfc5ff60_6114, \8340 );
nor \g453738/U$1 ( \14634 , \14632 , \14633 );
and \g454629/U$2 ( \14635 , \8313 , RIdea6c58_403);
and \g454629/U$3 ( \14636 , RIdead3f0_435, \8323 );
nor \g454629/U$1 ( \14637 , \14635 , \14636 );
not \g454628/U$1 ( \14638 , \14637 );
and \g450426/U$2 ( \14639 , \14638 , \8316 );
and \g450426/U$3 ( \14640 , RIdec68f0_723, \8351 );
nor \g450426/U$1 ( \14641 , \14639 , \14640 );
and \g453737/U$2 ( \14642 , \8356 , RIdeb00f0_467);
and \g453737/U$3 ( \14643 , RIfc9b8d0_6792, \8359 );
nor \g453737/U$1 ( \14644 , \14642 , \14643 );
nand \g448236/U$1 ( \14645 , \14631 , \14634 , \14641 , \14644 );
and \g444747/U$3 ( \14646 , \9702 , \14645 );
nor \g444747/U$1 ( \14647 , \14627 , \14646 );
and \g447158/U$2 ( \14648 , \11700 , RIdebe1f0_627);
and \g447158/U$3 ( \14649 , RIfc7ce08_6443, \11702 );
nor \g447158/U$1 ( \14650 , \14648 , \14649 );
and \g447160/U$2 ( \14651 , \9724 , RIdec0ef0_659);
and \g447160/U$3 ( \14652 , RIee208f0_4829, \9726 );
nor \g447160/U$1 ( \14653 , \14651 , \14652 );
and \g447159/U$2 ( \14654 , \9170 , RIdeb87f0_563);
and \g447159/U$3 ( \14655 , RIdebb4f0_595, \9172 );
nor \g447159/U$1 ( \14656 , \14654 , \14655 );
nand \g444539/U$1 ( \14657 , \14647 , \14650 , \14653 , \14656 );
and \g453756/U$2 ( \14658 , \8414 , RIdf076c0_1461);
and \g453756/U$3 ( \14659 , RIdf0a3c0_1493, \8409 );
nor \g453756/U$1 ( \14660 , \14658 , \14659 );
and \g446414/U$2 ( \14661 , RIdf0d0c0_1525, \8417 );
and \g446414/U$3 ( \14662 , RIdf0fdc0_1557, \8404 );
and \g449412/U$2 ( \14663 , RIdeee1c0_1173, \8317 );
and \g449412/U$3 ( \14664 , \8324 , RIdef0ec0_1205);
and \g449412/U$4 ( \14665 , RIdf157c0_1621, \8383 );
nor \g449412/U$1 ( \14666 , \14663 , \14664 , \14665 );
and \g453759/U$2 ( \14667 , \8335 , RIdeeb4c0_1141);
and \g453759/U$3 ( \14668 , RIdef3bc0_1237, \8340 );
nor \g453759/U$1 ( \14669 , \14667 , \14668 );
and \g455106/U$2 ( \14670 , \8313 , RIdef95c0_1301);
and \g455106/U$3 ( \14671 , RIdefc2c0_1333, \8323 );
nor \g455106/U$1 ( \14672 , \14670 , \14671 );
not \g450433/U$3 ( \14673 , \14672 );
not \g450433/U$4 ( \14674 , \8347 );
and \g450433/U$2 ( \14675 , \14673 , \14674 );
and \g450433/U$5 ( \14676 , \8351 , RIdf184c0_1653);
nor \g450433/U$1 ( \14677 , \14675 , \14676 );
and \g453758/U$2 ( \14678 , \8356 , RIdef68c0_1269);
and \g453758/U$3 ( \14679 , RIdefefc0_1365, \8359 );
nor \g453758/U$1 ( \14680 , \14678 , \14679 );
nand \g447954/U$1 ( \14681 , \14666 , \14669 , \14677 , \14680 );
nor \g446414/U$1 ( \14682 , \14661 , \14662 , \14681 );
and \g453757/U$2 ( \14683 , \8378 , RIdf049c0_1429);
and \g453757/U$3 ( \14684 , RIdf12ac0_1589, \8373 );
nor \g453757/U$1 ( \14685 , \14683 , \14684 );
nand \g445684/U$1 ( \14686 , \14660 , \14682 , \14685 );
and \g444806/U$2 ( \14687 , \14686 , \8478 );
and \g449410/U$2 ( \14688 , RIfcb5640_7086, \8531 );
and \g449410/U$3 ( \14689 , \8488 , RIfca4408_6891);
and \g449410/U$4 ( \14690 , RIfc6b900_6246, \8383 );
nor \g449410/U$1 ( \14691 , \14688 , \14689 , \14690 );
and \g453750/U$2 ( \14692 , \8335 , RIded4018_876);
and \g453750/U$3 ( \14693 , RIdeda990_951, \8340 );
nor \g453750/U$1 ( \14694 , \14692 , \14693 );
and \g454512/U$2 ( \14695 , \8313 , RIded61d8_900);
and \g454512/U$3 ( \14696 , RIded8500_925, \8323 );
nor \g454512/U$1 ( \14697 , \14695 , \14696 );
not \g454511/U$1 ( \14698 , \14697 );
and \g450431/U$2 ( \14699 , \14698 , \8316 );
and \g450431/U$3 ( \14700 , RIfc69b78_6225, \8351 );
nor \g450431/U$1 ( \14701 , \14699 , \14700 );
and \g453748/U$2 ( \14702 , \8356 , RIee21700_4839);
and \g453748/U$3 ( \14703 , RIfc7ff40_6478, \8359 );
nor \g453748/U$1 ( \14704 , \14702 , \14703 );
nand \g448237/U$1 ( \14705 , \14691 , \14694 , \14701 , \14704 );
and \g444806/U$3 ( \14706 , \8482 , \14705 );
nor \g444806/U$1 ( \14707 , \14687 , \14706 );
and \g447164/U$2 ( \14708 , \8964 , RIdee3d38_1056);
and \g447164/U$3 ( \14709 , RIdee5ac0_1077, \8966 );
nor \g447164/U$1 ( \14710 , \14708 , \14709 );
and \g447165/U$2 ( \14711 , \8969 , RIfced770_7724);
and \g447165/U$3 ( \14712 , RIfc4d270_5900, \8971 );
nor \g447165/U$1 ( \14713 , \14711 , \14712 );
and \g447166/U$2 ( \14714 , \8974 , RIdedfb20_1009);
and \g447166/U$3 ( \14715 , RIdee1a10_1031, \8976 );
nor \g447166/U$1 ( \14716 , \14714 , \14715 );
nand \g444540/U$1 ( \14717 , \14707 , \14710 , \14713 , \14716 );
and \g446405/U$2 ( \14718 , RIfc691a0_6218, \8356 );
and \g446405/U$3 ( \14719 , RIfcaad80_6966, \8340 );
and \g449402/U$2 ( \14720 , RIdf27100_1821, \8414 );
and \g449402/U$3 ( \14721 , \8409 , RIdf29428_1846);
and \g449402/U$4 ( \14722 , RIfcdcda8_7535, \8486 );
nor \g449402/U$1 ( \14723 , \14720 , \14721 , \14722 );
and \g454488/U$2 ( \14724 , \8313 , RIfc5c018_6069);
and \g454488/U$3 ( \14725 , RIfca1b40_6862, \8323 );
nor \g454488/U$1 ( \14726 , \14724 , \14725 );
not \g450422/U$3 ( \14727 , \14726 );
not \g450422/U$4 ( \14728 , \8328 );
and \g450422/U$2 ( \14729 , \14727 , \14728 );
and \g450422/U$5 ( \14730 , \8359 , RIfc5e1d8_6093);
nor \g450422/U$1 ( \14731 , \14729 , \14730 );
and \g453713/U$2 ( \14732 , \8404 , RIfe9ada0_8106);
and \g453713/U$3 ( \14733 , RIfcb1860_7042, \8351 );
nor \g453713/U$1 ( \14734 , \14732 , \14733 );
and \g453715/U$2 ( \14735 , \8378 , RIfe9af08_8107);
and \g453715/U$3 ( \14736 , RIdf2b318_1868, \8417 );
nor \g453715/U$1 ( \14737 , \14735 , \14736 );
nand \g447947/U$1 ( \14738 , \14723 , \14731 , \14734 , \14737 );
nor \g446405/U$1 ( \14739 , \14718 , \14719 , \14738 );
and \g453710/U$2 ( \14740 , \8335 , RIdf1a518_1676);
and \g453710/U$3 ( \14741 , RIfcac400_6982, \8531 );
nor \g453710/U$1 ( \14742 , \14740 , \14741 );
and \g453709/U$2 ( \14743 , \8319 , RIfc61b80_6134);
and \g453709/U$3 ( \14744 , RIdf20bc0_1749, \8326 );
nor \g453709/U$1 ( \14745 , \14743 , \14744 );
and \g445434/U$2 ( \14746 , \14739 , \14742 , \14745 );
nor \g445434/U$1 ( \14747 , \14746 , \8621 );
and \g446407/U$2 ( \14748 , RIdeb5af0_531, \8417 );
and \g446407/U$3 ( \14749 , RIdec95f0_755, \8404 );
and \g449404/U$2 ( \14750 , RIdedd528_982, \8319 );
and \g449404/U$3 ( \14751 , \8326 , RIdee87c0_1109);
and \g449404/U$4 ( \14752 , RIdeceff0_819, \8383 );
nor \g449404/U$1 ( \14753 , \14750 , \14751 , \14752 );
and \g453725/U$2 ( \14754 , \8335 , RIde7f9a0_212);
and \g453725/U$3 ( \14755 , RIdf01cc0_1397, \8340 );
nor \g453725/U$1 ( \14756 , \14754 , \14755 );
and \g455116/U$2 ( \14757 , \8313 , RIdf2dd48_1898);
and \g455116/U$3 ( \14758 , RIdf396e8_2030, \8323 );
nor \g455116/U$1 ( \14759 , \14757 , \14758 );
not \g450424/U$3 ( \14760 , \14759 );
not \g450424/U$4 ( \14761 , \8347 );
and \g450424/U$2 ( \14762 , \14760 , \14761 );
and \g450424/U$5 ( \14763 , \8351 , RIded1cf0_851);
nor \g450424/U$1 ( \14764 , \14762 , \14763 );
and \g453724/U$2 ( \14765 , \8356 , RIdf1e5c8_1722);
and \g453724/U$3 ( \14766 , RIe144cf0_2160, \8359 );
nor \g453724/U$1 ( \14767 , \14765 , \14766 );
nand \g447949/U$1 ( \14768 , \14753 , \14756 , \14764 , \14767 );
nor \g446407/U$1 ( \14769 , \14748 , \14749 , \14768 );
and \g453722/U$2 ( \14770 , \8378 , RIe15b4f0_2416);
and \g453722/U$3 ( \14771 , RIdecc2f0_787, \8373 );
nor \g453722/U$1 ( \14772 , \14770 , \14771 );
and \g453719/U$2 ( \14773 , \8414 , RIe16f6f8_2645);
and \g453719/U$3 ( \14774 , RIde99a58_339, \8407 );
nor \g453719/U$1 ( \14775 , \14773 , \14774 );
and \g445437/U$2 ( \14776 , \14769 , \14772 , \14775 );
nor \g445437/U$1 ( \14777 , \14776 , \8651 );
or \g444334/U$1 ( \14778 , \14657 , \14717 , \14747 , \14777 );
and \g446402/U$2 ( \14779 , RIee2e180_4983, \8356 );
and \g446402/U$3 ( \14780 , RIdf36b50_1999, \8340 );
and \g449397/U$2 ( \14781 , RIfc54890_5984, \8373 );
and \g449397/U$3 ( \14782 , \8383 , RIfc92f00_6694);
and \g449397/U$4 ( \14783 , RIee30340_5007, \8488 );
nor \g449397/U$1 ( \14784 , \14781 , \14782 , \14783 );
and \g455362/U$2 ( \14785 , \8313 , RIdf3dd38_2080);
and \g455362/U$3 ( \14786 , RIe13fe30_2104, \8323 );
nor \g455362/U$1 ( \14787 , \14785 , \14786 );
not \g450417/U$3 ( \14788 , \14787 );
not \g450417/U$4 ( \14789 , \8376 );
and \g450417/U$2 ( \14790 , \14788 , \14789 );
and \g450417/U$5 ( \14791 , \8359 , RIfc57590_6016);
nor \g450417/U$1 ( \14792 , \14790 , \14791 );
and \g453695/U$2 ( \14793 , \8404 , RIfcdcc40_7534);
and \g453695/U$3 ( \14794 , RIfcea098_7685, \8351 );
nor \g453695/U$1 ( \14795 , \14793 , \14794 );
and \g453696/U$2 ( \14796 , \8378 , RIdf3b8a8_2054);
and \g453696/U$3 ( \14797 , RIe142158_2129, \8417 );
nor \g453696/U$1 ( \14798 , \14796 , \14797 );
nand \g447943/U$1 ( \14799 , \14784 , \14792 , \14795 , \14798 );
nor \g446402/U$1 ( \14800 , \14779 , \14780 , \14799 );
and \g453693/U$2 ( \14801 , \8335 , RIfe9b070_8108);
and \g453693/U$3 ( \14802 , RIfcd0490_7392, \8531 );
nor \g453693/U$1 ( \14803 , \14801 , \14802 );
and \g453691/U$2 ( \14804 , \8317 , RIdf32398_1948);
and \g453691/U$3 ( \14805 , RIdf34558_1972, \8326 );
nor \g453691/U$1 ( \14806 , \14804 , \14805 );
and \g445430/U$2 ( \14807 , \14800 , \14803 , \14806 );
nor \g445430/U$1 ( \14808 , \14807 , \8422 );
and \g446404/U$2 ( \14809 , RIfcd5080_7446, \8531 );
and \g446404/U$3 ( \14810 , RIe14a6f0_2224, \8319 );
and \g449399/U$2 ( \14811 , RIe1587f0_2384, \8414 );
and \g449399/U$3 ( \14812 , \8409 , RIe15e1f0_2448);
and \g449399/U$4 ( \14813 , RIe152df0_2320, \8488 );
nor \g449399/U$1 ( \14814 , \14811 , \14812 , \14813 );
and \g455365/U$2 ( \14815 , \8313 , RIee381d0_5097);
and \g455365/U$3 ( \14816 , RIe163bf0_2512, \8323 );
nor \g455365/U$1 ( \14817 , \14815 , \14816 );
not \g450420/U$3 ( \14818 , \14817 );
not \g450420/U$4 ( \14819 , \8328 );
and \g450420/U$2 ( \14820 , \14818 , \14819 );
and \g450420/U$5 ( \14821 , \8359 , RIfc3f968_5749);
nor \g450420/U$1 ( \14822 , \14820 , \14821 );
and \g453705/U$2 ( \14823 , \8404 , RIe160ef0_2480);
and \g453705/U$3 ( \14824 , RIe1668f0_2544, \8351 );
nor \g453705/U$1 ( \14825 , \14823 , \14824 );
and \g453708/U$2 ( \14826 , \8378 , RIe155af0_2352);
and \g453708/U$3 ( \14827 , RIfcdfaa8_7567, \8417 );
nor \g453708/U$1 ( \14828 , \14826 , \14827 );
nand \g447945/U$1 ( \14829 , \14814 , \14822 , \14825 , \14828 );
nor \g446404/U$1 ( \14830 , \14809 , \14810 , \14829 );
and \g453703/U$2 ( \14831 , \8335 , RIe1479f0_2192);
and \g453703/U$3 ( \14832 , RIfc84b30_6532, \8340 );
nor \g453703/U$1 ( \14833 , \14831 , \14832 );
and \g453702/U$2 ( \14834 , \8326 , RIe14d3f0_2256);
and \g453702/U$3 ( \14835 , RIe1500f0_2288, \8356 );
nor \g453702/U$1 ( \14836 , \14834 , \14835 );
and \g445431/U$2 ( \14837 , \14830 , \14833 , \14836 );
nor \g445431/U$1 ( \14838 , \14837 , \8368 );
or \g444250/U$1 ( \14839 , \14778 , \14808 , \14838 );
_DC \g2f32/U$1 ( \14840 , \14839 , \8654 );
and \g447041/U$2 ( \14841 , \11521 , RIfe999f0_8092);
and \g447041/U$3 ( \14842 , RIfe99b58_8093, \11523 );
nor \g447041/U$1 ( \14843 , \14841 , \14842 );
and \g446272/U$2 ( \14844 , RIfc4a9a8_5871, \8488 );
and \g446272/U$3 ( \14845 , RIfc9ac28_6783, \8359 );
and \g449231/U$2 ( \14846 , RIdf1ba30_1691, \8319 );
and \g449231/U$3 ( \14847 , \8326 , RIdf20a58_1748);
and \g449231/U$4 ( \14848 , RIdf292c0_1845, \8409 );
nor \g449231/U$1 ( \14849 , \14846 , \14847 , \14848 );
and \g453080/U$2 ( \14850 , \8335 , RIfe99cc0_8094);
and \g453080/U$3 ( \14851 , RIdf220d8_1764, \8340 );
nor \g453080/U$1 ( \14852 , \14850 , \14851 );
and \g453079/U$2 ( \14853 , \8404 , RIfcbad70_7148);
and \g453079/U$3 ( \14854 , RIfc83078_6513, \8351 );
nor \g453079/U$1 ( \14855 , \14853 , \14854 );
and \g455208/U$2 ( \14856 , \8313 , RIfc9ad90_6784);
and \g455208/U$3 ( \14857 , RIfcb6e28_7103, \8323 );
nor \g455208/U$1 ( \14858 , \14856 , \14857 );
not \g450247/U$3 ( \14859 , \14858 );
not \g450247/U$4 ( \14860 , \8328 );
and \g450247/U$2 ( \14861 , \14859 , \14860 );
and \g450247/U$5 ( \14862 , \8417 , RIdf2b1b0_1867);
nor \g450247/U$1 ( \14863 , \14861 , \14862 );
nand \g447849/U$1 ( \14864 , \14849 , \14852 , \14855 , \14863 );
nor \g446272/U$1 ( \14865 , \14844 , \14845 , \14864 );
not \g444819/U$3 ( \14866 , \14865 );
not \g444819/U$4 ( \14867 , \8621 );
and \g444819/U$2 ( \14868 , \14866 , \14867 );
and \g446274/U$2 ( \14869 , RIdf07558_1460, \8412 );
and \g446274/U$3 ( \14870 , RIdef6758_1268, \8356 );
and \g449233/U$2 ( \14871 , RIdf0a258_1492, \8409 );
and \g449233/U$3 ( \14872 , \8373 , RIdf12958_1588);
and \g449233/U$4 ( \14873 , RIdf15658_1620, \8383 );
nor \g449233/U$1 ( \14874 , \14871 , \14872 , \14873 );
and \g453091/U$2 ( \14875 , \8335 , RIdeeb358_1140);
and \g453091/U$3 ( \14876 , RIdef3a58_1236, \8340 );
nor \g453091/U$1 ( \14877 , \14875 , \14876 );
and \g453090/U$2 ( \14878 , \8404 , RIdf0fc58_1556);
and \g453090/U$3 ( \14879 , RIdf18358_1652, \8351 );
nor \g453090/U$1 ( \14880 , \14878 , \14879 );
and \g455216/U$2 ( \14881 , \8313 , RIdeee058_1172);
and \g455216/U$3 ( \14882 , RIdef0d58_1204, \8323 );
nor \g455216/U$1 ( \14883 , \14881 , \14882 );
not \g455215/U$1 ( \14884 , \14883 );
and \g450248/U$2 ( \14885 , \14884 , \8316 );
and \g450248/U$3 ( \14886 , RIdf0cf58_1524, \8417 );
nor \g450248/U$1 ( \14887 , \14885 , \14886 );
nand \g448213/U$1 ( \14888 , \14874 , \14877 , \14880 , \14887 );
nor \g446274/U$1 ( \14889 , \14869 , \14870 , \14888 );
and \g453087/U$2 ( \14890 , \8378 , RIdf04858_1428);
and \g453087/U$3 ( \14891 , RIdefee58_1364, \8359 );
nor \g453087/U$1 ( \14892 , \14890 , \14891 );
and \g453086/U$2 ( \14893 , \8531 , RIdef9458_1300);
and \g453086/U$3 ( \14894 , RIdefc158_1332, \8488 );
nor \g453086/U$1 ( \14895 , \14893 , \14894 );
and \g445347/U$2 ( \14896 , \14889 , \14892 , \14895 );
nor \g445347/U$1 ( \14897 , \14896 , \8477 );
nor \g444819/U$1 ( \14898 , \14868 , \14897 );
and \g447040/U$2 ( \14899 , \13486 , RIfc82da8_6511);
and \g447040/U$3 ( \14900 , RIdf23758_1780, \13488 );
nor \g447040/U$1 ( \14901 , \14899 , \14900 );
nand \g444430/U$1 ( \14902 , \14843 , \14898 , \14901 );
and \g453104/U$2 ( \14903 , \8531 , RIfc9f3e0_6834);
and \g453104/U$3 ( \14904 , RIfc89b58_6589, \8486 );
nor \g453104/U$1 ( \14905 , \14903 , \14904 );
and \g446277/U$2 ( \14906 , RIfe99f90_8096, \8414 );
and \g446277/U$3 ( \14907 , RIfc82538_6505, \8356 );
and \g449238/U$2 ( \14908 , RIdee3bd0_1055, \8409 );
and \g449238/U$3 ( \14909 , \8373 , RIfc52568_5959);
and \g449238/U$4 ( \14910 , RIee24b08_4876, \8383 );
nor \g449238/U$1 ( \14911 , \14908 , \14909 , \14910 );
and \g453109/U$2 ( \14912 , \8335 , RIded3eb0_875);
and \g453109/U$3 ( \14913 , RIdeda828_950, \8340 );
nor \g453109/U$1 ( \14914 , \14912 , \14913 );
and \g453108/U$2 ( \14915 , \8404 , RIfc826a0_6506);
and \g453108/U$3 ( \14916 , RIee25918_4886, \8351 );
nor \g453108/U$1 ( \14917 , \14915 , \14916 );
and \g454515/U$2 ( \14918 , \8313 , RIfeabe70_8272);
and \g454515/U$3 ( \14919 , RIded8398_924, \8323 );
nor \g454515/U$1 ( \14920 , \14918 , \14919 );
not \g454514/U$1 ( \14921 , \14920 );
and \g450254/U$2 ( \14922 , \14921 , \8316 );
and \g450254/U$3 ( \14923 , RIdee5958_1076, \8417 );
nor \g450254/U$1 ( \14924 , \14922 , \14923 );
nand \g448216/U$1 ( \14925 , \14911 , \14914 , \14917 , \14924 );
nor \g446277/U$1 ( \14926 , \14906 , \14907 , \14925 );
and \g453106/U$2 ( \14927 , \8378 , RIdedf9b8_1008);
and \g453106/U$3 ( \14928 , RIfce4800_7622, \8359 );
nor \g453106/U$1 ( \14929 , \14927 , \14928 );
nand \g445645/U$1 ( \14930 , \14905 , \14926 , \14929 );
and \g444921/U$2 ( \14931 , \14930 , \8482 );
and \g449236/U$2 ( \14932 , RIdee8658_1108, \8326 );
and \g449236/U$3 ( \14933 , \8531 , RIdf2dbe0_1897);
and \g449236/U$4 ( \14934 , RIdf39580_2029, \8488 );
nor \g449236/U$1 ( \14935 , \14932 , \14933 , \14934 );
and \g453101/U$2 ( \14936 , \8356 , RIdf1e460_1721);
and \g453101/U$3 ( \14937 , RIe144b88_2159, \8359 );
nor \g453101/U$1 ( \14938 , \14936 , \14937 );
and \g455222/U$2 ( \14939 , \8313 , RIe16f590_2644);
and \g455222/U$3 ( \14940 , RIde99710_338, \8323 );
nor \g455222/U$1 ( \14941 , \14939 , \14940 );
not \g450251/U$3 ( \14942 , \14941 );
not \g450251/U$4 ( \14943 , \8376 );
and \g450251/U$2 ( \14944 , \14942 , \14943 );
and \g450251/U$5 ( \14945 , \8340 , RIdf01b58_1396);
nor \g450251/U$1 ( \14946 , \14944 , \14945 );
and \g453099/U$2 ( \14947 , \8378 , RIe15b388_2415);
and \g453099/U$3 ( \14948 , RIdeb5988_530, \8417 );
nor \g453099/U$1 ( \14949 , \14947 , \14948 );
nand \g447850/U$1 ( \14950 , \14935 , \14938 , \14946 , \14949 );
and \g444921/U$3 ( \14951 , \9010 , \14950 );
nor \g444921/U$1 ( \14952 , \14931 , \14951 );
and \g447046/U$2 ( \14953 , \9041 , RIdec9488_754);
and \g447046/U$3 ( \14954 , RIdecc188_786, \9043 );
nor \g447046/U$1 ( \14955 , \14953 , \14954 );
nor \g448375/U$1 ( \14956 , \8651 , \8382 );
and \g447045/U$2 ( \14957 , \14956 , RIdecee88_818);
nor \g448317/U$1 ( \14958 , \8651 , \9295 );
and \g447045/U$3 ( \14959 , RIded1b88_850, \14958 );
nor \g447045/U$1 ( \14960 , \14957 , \14959 );
and \g447048/U$2 ( \14961 , \13244 , RIde7f658_211);
and \g447048/U$3 ( \14962 , RIdedd3c0_981, \13246 );
nor \g447048/U$1 ( \14963 , \14961 , \14962 );
nand \g444640/U$1 ( \14964 , \14952 , \14955 , \14960 , \14963 );
and \g446268/U$2 ( \14965 , RIfc831e0_6514, \8373 );
and \g446268/U$3 ( \14966 , RIee338b0_5045, \8383 );
and \g449226/U$2 ( \14967 , RIdf343f0_1971, \8326 );
and \g449226/U$3 ( \14968 , \8531 , RIfcba938_7145);
and \g449226/U$4 ( \14969 , RIee301d8_5006, \8488 );
nor \g449226/U$1 ( \14970 , \14967 , \14968 , \14969 );
and \g453063/U$2 ( \14971 , \8356 , RIee2e018_4982);
and \g453063/U$3 ( \14972 , RIfcb6f90_7104, \8359 );
nor \g453063/U$1 ( \14973 , \14971 , \14972 );
and \g454407/U$2 ( \14974 , \8313 , RIdf3dbd0_2079);
and \g454407/U$3 ( \14975 , RIe13fcc8_2103, \8323 );
nor \g454407/U$1 ( \14976 , \14974 , \14975 );
not \g450241/U$3 ( \14977 , \14976 );
not \g450241/U$4 ( \14978 , \8376 );
and \g450241/U$2 ( \14979 , \14977 , \14978 );
and \g450241/U$5 ( \14980 , \8340 , RIdf369e8_1998);
nor \g450241/U$1 ( \14981 , \14979 , \14980 );
and \g453062/U$2 ( \14982 , \8378 , RIdf3b740_2053);
and \g453062/U$3 ( \14983 , RIe141ff0_2128, \8417 );
nor \g453062/U$1 ( \14984 , \14982 , \14983 );
nand \g447844/U$1 ( \14985 , \14970 , \14973 , \14981 , \14984 );
nor \g446268/U$1 ( \14986 , \14965 , \14966 , \14985 );
and \g453055/U$2 ( \14987 , \8335 , RIfe99e28_8095);
and \g453055/U$3 ( \14988 , RIee34990_5057, \8351 );
nor \g453055/U$1 ( \14989 , \14987 , \14988 );
and \g453058/U$2 ( \14990 , \8319 , RIdf32230_1947);
and \g453058/U$3 ( \14991 , RIfcd3b68_7431, \8404 );
nor \g453058/U$1 ( \14992 , \14990 , \14991 );
and \g445343/U$2 ( \14993 , \14986 , \14989 , \14992 );
nor \g445343/U$1 ( \14994 , \14993 , \8422 );
and \g446270/U$2 ( \14995 , RIe158688_2383, \8414 );
and \g446270/U$3 ( \14996 , RIe14ff88_2287, \8356 );
and \g449228/U$2 ( \14997 , RIe14a588_2223, \8319 );
and \g449228/U$3 ( \14998 , \8326 , RIe14d288_2255);
and \g449228/U$4 ( \14999 , RIe15e088_2447, \8409 );
nor \g449228/U$1 ( \15000 , \14997 , \14998 , \14999 );
and \g453071/U$2 ( \15001 , \8335 , RIe147888_2191);
and \g453071/U$3 ( \15002 , RIfc51cf8_5953, \8340 );
nor \g453071/U$1 ( \15003 , \15001 , \15002 );
and \g453070/U$2 ( \15004 , \8404 , RIe160d88_2479);
and \g453070/U$3 ( \15005 , RIe166788_2543, \8351 );
nor \g453070/U$1 ( \15006 , \15004 , \15005 );
and \g454743/U$2 ( \15007 , \8313 , RIfc83618_6517);
and \g454743/U$3 ( \15008 , RIe163a88_2511, \8323 );
nor \g454743/U$1 ( \15009 , \15007 , \15008 );
not \g450244/U$3 ( \15010 , \15009 );
not \g450244/U$4 ( \15011 , \8328 );
and \g450244/U$2 ( \15012 , \15010 , \15011 );
and \g450244/U$5 ( \15013 , \8417 , RIee36718_5078);
nor \g450244/U$1 ( \15014 , \15012 , \15013 );
nand \g447847/U$1 ( \15015 , \15000 , \15003 , \15006 , \15014 );
nor \g446270/U$1 ( \15016 , \14995 , \14996 , \15015 );
and \g453068/U$2 ( \15017 , \8378 , RIe155988_2351);
and \g453068/U$3 ( \15018 , RIfc3f800_5748, \8359 );
nor \g453068/U$1 ( \15019 , \15017 , \15018 );
and \g453066/U$2 ( \15020 , \8531 , RIfc895b8_6585);
and \g453066/U$3 ( \15021 , RIe152c88_2319, \8488 );
nor \g453066/U$1 ( \15022 , \15020 , \15021 );
and \g445345/U$2 ( \15023 , \15016 , \15019 , \15022 );
nor \g445345/U$1 ( \15024 , \15023 , \8368 );
or \g444303/U$1 ( \15025 , \14902 , \14964 , \14994 , \15024 );
and \g446263/U$2 ( \15026 , RIee1b5f8_4770, \8373 );
and \g446263/U$3 ( \15027 , RIee1c570_4781, \8383 );
and \g449222/U$2 ( \15028 , RIfe99720_8090, \8414 );
and \g449222/U$3 ( \15029 , \8409 , RIfe99450_8088);
and \g449222/U$4 ( \15030 , RIe16c890_2612, \8326 );
nor \g449222/U$1 ( \15031 , \15028 , \15029 , \15030 );
and \g453044/U$2 ( \15032 , \8356 , RIfc89450_6584);
and \g453044/U$3 ( \15033 , RIde83168_229, \8359 );
nor \g453044/U$1 ( \15034 , \15032 , \15033 );
and \g455189/U$2 ( \15035 , \8313 , RIfcd5a58_7453);
and \g455189/U$3 ( \15036 , RIfcc43e8_7255, \8323 );
nor \g455189/U$1 ( \15037 , \15035 , \15036 );
not \g450237/U$3 ( \15038 , \15037 );
not \g450237/U$4 ( \15039 , \8347 );
and \g450237/U$2 ( \15040 , \15038 , \15039 );
and \g450237/U$5 ( \15041 , \8340 , RIfcc5798_7269);
nor \g450237/U$1 ( \15042 , \15040 , \15041 );
and \g453043/U$2 ( \15043 , \8378 , RIfe995b8_8089);
and \g453043/U$3 ( \15044 , RIfe99888_8091, \8417 );
nor \g453043/U$1 ( \15045 , \15043 , \15044 );
nand \g447841/U$1 ( \15046 , \15031 , \15034 , \15042 , \15045 );
nor \g446263/U$1 ( \15047 , \15026 , \15027 , \15046 );
and \g453036/U$2 ( \15048 , \8335 , RIe168d80_2570);
and \g453036/U$3 ( \15049 , RIee1d650_4793, \8351 );
nor \g453036/U$1 ( \15050 , \15048 , \15049 );
and \g453039/U$2 ( \15051 , \8319 , RIe16a568_2587);
and \g453039/U$3 ( \15052 , RIee1aef0_4765, \8404 );
nor \g453039/U$1 ( \15053 , \15051 , \15052 );
and \g445337/U$2 ( \15054 , \15047 , \15050 , \15053 );
nor \g445337/U$1 ( \15055 , \15054 , \8558 );
and \g446265/U$2 ( \15056 , RIdebb388_594, \8414 );
and \g446265/U$3 ( \15057 , RIfce1f38_7593, \8531 );
and \g449224/U$2 ( \15058 , RIdea6910_402, \8319 );
and \g449224/U$3 ( \15059 , \8326 , RIdead210_434);
and \g449224/U$4 ( \15060 , RIdebe088_626, \8409 );
nor \g449224/U$1 ( \15061 , \15058 , \15059 , \15060 );
and \g453051/U$2 ( \15062 , \8335 , RIdea0010_370);
and \g453051/U$3 ( \15063 , RIfc892e8_6583, \8340 );
nor \g453051/U$1 ( \15064 , \15062 , \15063 );
and \g453050/U$2 ( \15065 , \8404 , RIdec0d88_658);
and \g453050/U$3 ( \15066 , RIdec6788_722, \8351 );
nor \g453050/U$1 ( \15067 , \15065 , \15066 );
and \g454378/U$2 ( \15068 , \8313 , RIee20788_4828);
and \g454378/U$3 ( \15069 , RIdec3a88_690, \8323 );
nor \g454378/U$1 ( \15070 , \15068 , \15069 );
not \g450239/U$3 ( \15071 , \15070 );
not \g450239/U$4 ( \15072 , \8328 );
and \g450239/U$2 ( \15073 , \15071 , \15072 );
and \g450239/U$5 ( \15074 , \8417 , RIee1f810_4817);
nor \g450239/U$1 ( \15075 , \15073 , \15074 );
nand \g447843/U$1 ( \15076 , \15061 , \15064 , \15067 , \15075 );
nor \g446265/U$1 ( \15077 , \15056 , \15057 , \15076 );
and \g453047/U$2 ( \15078 , \8356 , RIdeaff88_466);
and \g453047/U$3 ( \15079 , RIfc9b1c8_6787, \8359 );
nor \g453047/U$1 ( \15080 , \15078 , \15079 );
and \g453048/U$2 ( \15081 , \8378 , RIdeb8688_562);
and \g453048/U$3 ( \15082 , RIdeb2c88_498, \8488 );
nor \g453048/U$1 ( \15083 , \15081 , \15082 );
and \g445340/U$2 ( \15084 , \15077 , \15080 , \15083 );
nor \g445340/U$1 ( \15085 , \15084 , \8589 );
or \g444247/U$1 ( \15086 , \15025 , \15055 , \15085 );
_DC \g2fb7/U$1 ( \15087 , \15086 , \8654 );
and \g453270/U$2 ( \15088 , \8326 , RIdee84f0_1107);
and \g453270/U$3 ( \15089 , RIdec9320_753, \8404 );
nor \g453270/U$1 ( \15090 , \15088 , \15089 );
and \g446311/U$2 ( \15091 , RIdecc020_785, \8371 );
and \g446311/U$3 ( \15092 , RIdedd258_980, \8317 );
and \g449283/U$2 ( \15093 , RIdf2da78_1896, \8531 );
and \g449283/U$3 ( \15094 , \8486 , RIdf39418_2028);
and \g449283/U$4 ( \15095 , RIdeced20_817, \8383 );
nor \g449283/U$1 ( \15096 , \15093 , \15094 , \15095 );
and \g453275/U$2 ( \15097 , \8356 , RIdf1e2f8_1720);
and \g453275/U$3 ( \15098 , RIe144a20_2158, \8359 );
nor \g453275/U$1 ( \15099 , \15097 , \15098 );
and \g455270/U$2 ( \15100 , \8313 , RIe16f428_2643);
and \g455270/U$3 ( \15101 , RIde993c8_337, \8323 );
nor \g455270/U$1 ( \15102 , \15100 , \15101 );
not \g450299/U$3 ( \15103 , \15102 );
not \g450299/U$4 ( \15104 , \8376 );
and \g450299/U$2 ( \15105 , \15103 , \15104 );
and \g450299/U$5 ( \15106 , \8351 , RIded1a20_849);
nor \g450299/U$1 ( \15107 , \15105 , \15106 );
and \g453273/U$2 ( \15108 , \8378 , RIe15b220_2414);
and \g453273/U$3 ( \15109 , RIdeb5820_529, \8417 );
nor \g453273/U$1 ( \15110 , \15108 , \15109 );
nand \g447876/U$1 ( \15111 , \15096 , \15099 , \15107 , \15110 );
nor \g446311/U$1 ( \15112 , \15091 , \15092 , \15111 );
and \g453271/U$2 ( \15113 , \8335 , RIde7f310_210);
and \g453271/U$3 ( \15114 , RIdf019f0_1395, \8340 );
nor \g453271/U$1 ( \15115 , \15113 , \15114 );
nand \g445655/U$1 ( \15116 , \15090 , \15112 , \15115 );
and \g444884/U$2 ( \15117 , \15116 , \9010 );
and \g449281/U$2 ( \15118 , RIdf1b8c8_1690, \8319 );
and \g449281/U$3 ( \15119 , \8326 , RIdf208f0_1747);
and \g449281/U$4 ( \15120 , RIfc48950_5848, \8488 );
nor \g449281/U$1 ( \15121 , \15118 , \15119 , \15120 );
and \g453267/U$2 ( \15122 , \8335 , RIdf1a3b0_1675);
and \g453267/U$3 ( \15123 , RIdf21f70_1763, \8340 );
nor \g453267/U$1 ( \15124 , \15122 , \15123 );
and \g453266/U$2 ( \15125 , \8404 , RIfc80210_6480);
and \g453266/U$3 ( \15126 , RIfcc3740_7246, \8351 );
nor \g453266/U$1 ( \15127 , \15125 , \15126 );
and \g454457/U$2 ( \15128 , \8313 , RIfce05e8_7575);
and \g454457/U$3 ( \15129 , RIfc48ab8_5849, \8323 );
nor \g454457/U$1 ( \15130 , \15128 , \15129 );
not \g450298/U$3 ( \15131 , \15130 );
not \g450298/U$4 ( \15132 , \8328 );
and \g450298/U$2 ( \15133 , \15131 , \15132 );
and \g450298/U$5 ( \15134 , \8359 , RIfc8bbb0_6612);
nor \g450298/U$1 ( \15135 , \15133 , \15134 );
nand \g447875/U$1 ( \15136 , \15121 , \15124 , \15127 , \15135 );
and \g444884/U$3 ( \15137 , \8752 , \15136 );
nor \g444884/U$1 ( \15138 , \15117 , \15137 );
and \g447081/U$2 ( \15139 , \11516 , RIdf29158_1844);
and \g447081/U$3 ( \15140 , RIdf2b048_1866, \11518 );
nor \g447081/U$1 ( \15141 , \15139 , \15140 );
and \g447082/U$2 ( \15142 , \13486 , RIfc8bd18_6613);
and \g447082/U$3 ( \15143 , RIdf235f0_1779, \13488 );
nor \g447082/U$1 ( \15144 , \15142 , \15143 );
and \g447084/U$2 ( \15145 , \11521 , RIdf254e0_1801);
and \g447084/U$3 ( \15146 , RIdf26f98_1820, \11523 );
nor \g447084/U$1 ( \15147 , \15145 , \15146 );
nand \g444648/U$1 ( \15148 , \15138 , \15141 , \15144 , \15147 );
and \g453283/U$2 ( \15149 , \8531 , RIfce43c8_7619);
and \g453283/U$3 ( \15150 , RIdee18a8_1030, \8414 );
nor \g453283/U$1 ( \15151 , \15149 , \15150 );
and \g446313/U$2 ( \15152 , RIdee3a68_1054, \8409 );
and \g446313/U$3 ( \15153 , RIdedf850_1007, \8378 );
and \g449287/U$2 ( \15154 , RIfc99710_6768, \8373 );
and \g449287/U$3 ( \15155 , \8383 , RIfcd9838_7497);
and \g449287/U$4 ( \15156 , RIfcb5370_7084, \8488 );
nor \g449287/U$1 ( \15157 , \15154 , \15155 , \15156 );
and \g453287/U$2 ( \15158 , \8335 , RIded3d48_874);
and \g453287/U$3 ( \15159 , RIdeda6c0_949, \8340 );
nor \g453287/U$1 ( \15160 , \15158 , \15159 );
and \g453286/U$2 ( \15161 , \8404 , RIfca1168_6855);
and \g453286/U$3 ( \15162 , RIfcbc120_7162, \8351 );
nor \g453286/U$1 ( \15163 , \15161 , \15162 );
and \g455308/U$2 ( \15164 , \8313 , RIded6070_899);
and \g455308/U$3 ( \15165 , RIded8230_923, \8323 );
nor \g455308/U$1 ( \15166 , \15164 , \15165 );
not \g455307/U$1 ( \15167 , \15166 );
and \g450303/U$2 ( \15168 , \15167 , \8316 );
and \g450303/U$3 ( \15169 , RIfc549f8_5985, \8359 );
nor \g450303/U$1 ( \15170 , \15168 , \15169 );
nand \g448224/U$1 ( \15171 , \15157 , \15160 , \15163 , \15170 );
nor \g446313/U$1 ( \15172 , \15152 , \15153 , \15171 );
and \g453284/U$2 ( \15173 , \8356 , RIfce0480_7574);
and \g453284/U$3 ( \15174 , RIdee57f0_1075, \8417 );
nor \g453284/U$1 ( \15175 , \15173 , \15174 );
nand \g445656/U$1 ( \15176 , \15151 , \15172 , \15175 );
and \g444829/U$2 ( \15177 , \15176 , \8482 );
and \g449285/U$2 ( \15178 , RIdef92f0_1299, \8531 );
and \g449285/U$3 ( \15179 , \8486 , RIdefbff0_1331);
and \g449285/U$4 ( \15180 , RIdf154f0_1619, \8383 );
nor \g449285/U$1 ( \15181 , \15178 , \15179 , \15180 );
and \g453280/U$2 ( \15182 , \8356 , RIdef65f0_1267);
and \g453280/U$3 ( \15183 , RIdefecf0_1363, \8359 );
nor \g453280/U$1 ( \15184 , \15182 , \15183 );
and \g455306/U$2 ( \15185 , \8313 , RIdf073f0_1459);
and \g455306/U$3 ( \15186 , RIdf0a0f0_1491, \8323 );
nor \g455306/U$1 ( \15187 , \15185 , \15186 );
not \g450302/U$3 ( \15188 , \15187 );
not \g450302/U$4 ( \15189 , \8376 );
and \g450302/U$2 ( \15190 , \15188 , \15189 );
and \g450302/U$5 ( \15191 , \8351 , RIdf181f0_1651);
nor \g450302/U$1 ( \15192 , \15190 , \15191 );
and \g453279/U$2 ( \15193 , \8378 , RIdf046f0_1427);
and \g453279/U$3 ( \15194 , RIdf0cdf0_1523, \8417 );
nor \g453279/U$1 ( \15195 , \15193 , \15194 );
nand \g447877/U$1 ( \15196 , \15181 , \15184 , \15192 , \15195 );
and \g444829/U$3 ( \15197 , \8478 , \15196 );
nor \g444829/U$1 ( \15198 , \15177 , \15197 );
and \g447086/U$2 ( \15199 , \8780 , RIdef0bf0_1203);
and \g447086/U$3 ( \15200 , RIdef38f0_1235, \8782 );
nor \g447086/U$1 ( \15201 , \15199 , \15200 );
and \g447085/U$2 ( \15202 , \9480 , RIdf0faf0_1555);
and \g447085/U$3 ( \15203 , RIdf127f0_1587, \9482 );
nor \g447085/U$1 ( \15204 , \15202 , \15203 );
and \g447087/U$2 ( \15205 , \8785 , RIdeeb1f0_1139);
and \g447087/U$3 ( \15206 , RIdeedef0_1171, \8787 );
nor \g447087/U$1 ( \15207 , \15205 , \15206 );
nand \g444649/U$1 ( \15208 , \15198 , \15201 , \15204 , \15207 );
and \g446306/U$2 ( \15209 , RIdebdf20_625, \8409 );
and \g446306/U$3 ( \15210 , RIdeb8520_561, \8378 );
and \g449276/U$2 ( \15211 , RIfc49328_5855, \8373 );
and \g449276/U$3 ( \15212 , \8383 , RIdec3920_689);
and \g449276/U$4 ( \15213 , RIdeb2b20_497, \8488 );
nor \g449276/U$1 ( \15214 , \15211 , \15212 , \15213 );
and \g453253/U$2 ( \15215 , \8335 , RIde9fcc8_369);
and \g453253/U$3 ( \15216 , RIfc491c0_5854, \8340 );
nor \g453253/U$1 ( \15217 , \15215 , \15216 );
and \g453252/U$2 ( \15218 , \8404 , RIdec0c20_657);
and \g453252/U$3 ( \15219 , RIdec6620_721, \8351 );
nor \g453252/U$1 ( \15220 , \15218 , \15219 );
and \g455302/U$2 ( \15221 , \8313 , RIdea65c8_401);
and \g455302/U$3 ( \15222 , RIdeacec8_433, \8323 );
nor \g455302/U$1 ( \15223 , \15221 , \15222 );
not \g455301/U$1 ( \15224 , \15223 );
and \g450294/U$2 ( \15225 , \15224 , \8316 );
and \g450294/U$3 ( \15226 , RIfc80648_6483, \8359 );
nor \g450294/U$1 ( \15227 , \15225 , \15226 );
nand \g448223/U$1 ( \15228 , \15214 , \15217 , \15220 , \15227 );
nor \g446306/U$1 ( \15229 , \15209 , \15210 , \15228 );
and \g453250/U$2 ( \15230 , \8356 , RIdeafe20_465);
and \g453250/U$3 ( \15231 , RIfc80eb8_6489, \8417 );
nor \g453250/U$1 ( \15232 , \15230 , \15231 );
and \g453249/U$2 ( \15233 , \8531 , RIfc8b340_6606);
and \g453249/U$3 ( \15234 , RIdebb220_593, \8414 );
nor \g453249/U$1 ( \15235 , \15233 , \15234 );
and \g445368/U$2 ( \15236 , \15229 , \15232 , \15235 );
nor \g445368/U$1 ( \15237 , \15236 , \8589 );
and \g446309/U$2 ( \15238 , RIfce4698_7621, \8371 );
and \g446309/U$3 ( \15239 , RIe16a400_2586, \8319 );
and \g449278/U$2 ( \15240 , RIfc48d88_5851, \8531 );
and \g449278/U$3 ( \15241 , \8488 , RIfcbba18_7157);
and \g449278/U$4 ( \15242 , RIfe98208_8075, \8383 );
nor \g449278/U$1 ( \15243 , \15240 , \15241 , \15242 );
and \g453261/U$2 ( \15244 , \8356 , RIfc99f80_6774);
and \g453261/U$3 ( \15245 , RIde82e20_228, \8359 );
nor \g453261/U$1 ( \15246 , \15244 , \15245 );
and \g454472/U$2 ( \15247 , \8313 , RIde8b4a8_269);
and \g454472/U$3 ( \15248 , RIde8f648_289, \8323 );
nor \g454472/U$1 ( \15249 , \15247 , \15248 );
not \g450295/U$3 ( \15250 , \15249 );
not \g450295/U$4 ( \15251 , \8376 );
and \g450295/U$2 ( \15252 , \15250 , \15251 );
and \g450295/U$5 ( \15253 , \8351 , RIfcd9c70_7500);
nor \g450295/U$1 ( \15254 , \15252 , \15253 );
and \g453260/U$2 ( \15255 , \8378 , RIde87308_249);
and \g453260/U$3 ( \15256 , RIde93158_307, \8417 );
nor \g453260/U$1 ( \15257 , \15255 , \15256 );
nand \g447871/U$1 ( \15258 , \15243 , \15246 , \15254 , \15257 );
nor \g446309/U$1 ( \15259 , \15238 , \15239 , \15258 );
and \g453257/U$2 ( \15260 , \8335 , RIe168c18_2569);
and \g453257/U$3 ( \15261 , RIfc8b4a8_6607, \8340 );
nor \g453257/U$1 ( \15262 , \15260 , \15261 );
and \g453256/U$2 ( \15263 , \8326 , RIe16c728_2611);
and \g453256/U$3 ( \15264 , RIfe980a0_8074, \8404 );
nor \g453256/U$1 ( \15265 , \15263 , \15264 );
and \g445369/U$2 ( \15266 , \15259 , \15262 , \15265 );
nor \g445369/U$1 ( \15267 , \15266 , \8558 );
or \g444407/U$1 ( \15268 , \15148 , \15208 , \15237 , \15267 );
and \g446304/U$2 ( \15269 , RIfc48248_5843, \8417 );
and \g446304/U$3 ( \15270 , RIe14fe20_2286, \8356 );
and \g449272/U$2 ( \15271 , RIe14a420_2222, \8317 );
and \g449272/U$3 ( \15272 , \8326 , RIe14d120_2254);
and \g449272/U$4 ( \15273 , RIe152b20_2318, \8486 );
nor \g449272/U$1 ( \15274 , \15271 , \15272 , \15273 );
and \g453240/U$2 ( \15275 , \8335 , RIe147720_2190);
and \g453240/U$3 ( \15276 , RIfca0e98_6853, \8340 );
nor \g453240/U$1 ( \15277 , \15275 , \15276 );
and \g453239/U$2 ( \15278 , \8404 , RIe160c20_2478);
and \g453239/U$3 ( \15279 , RIe166620_2542, \8351 );
nor \g453239/U$1 ( \15280 , \15278 , \15279 );
and \g454530/U$2 ( \15281 , \8313 , RIee38068_5096);
and \g454530/U$3 ( \15282 , RIe163920_2510, \8323 );
nor \g454530/U$1 ( \15283 , \15281 , \15282 );
not \g450289/U$3 ( \15284 , \15283 );
not \g450289/U$4 ( \15285 , \8328 );
and \g450289/U$2 ( \15286 , \15284 , \15285 );
and \g450289/U$5 ( \15287 , \8359 , RIfcbbe50_7160);
nor \g450289/U$1 ( \15288 , \15286 , \15287 );
nand \g447869/U$1 ( \15289 , \15274 , \15277 , \15280 , \15288 );
nor \g446304/U$1 ( \15290 , \15269 , \15270 , \15289 );
and \g453238/U$2 ( \15291 , \8378 , RIe155820_2350);
and \g453238/U$3 ( \15292 , RIfc47e10_5840, \8531 );
nor \g453238/U$1 ( \15293 , \15291 , \15292 );
and \g453237/U$2 ( \15294 , \8414 , RIe158520_2382);
and \g453237/U$3 ( \15295 , RIe15df20_2446, \8409 );
nor \g453237/U$1 ( \15296 , \15294 , \15295 );
and \g445365/U$2 ( \15297 , \15290 , \15293 , \15296 );
nor \g445365/U$1 ( \15298 , \15297 , \8368 );
and \g446305/U$2 ( \15299 , RIe13fb60_2102, \8409 );
and \g446305/U$3 ( \15300 , RIdf3b5d8_2052, \8378 );
and \g449274/U$2 ( \15301 , RIdf320c8_1946, \8319 );
and \g449274/U$3 ( \15302 , \8326 , RIdf34288_1970);
and \g449274/U$4 ( \15303 , RIee30070_5005, \8486 );
nor \g449274/U$1 ( \15304 , \15301 , \15302 , \15303 );
and \g453246/U$2 ( \15305 , \8335 , RIfe97dd0_8072);
and \g453246/U$3 ( \15306 , RIdf36880_1997, \8340 );
nor \g453246/U$1 ( \15307 , \15305 , \15306 );
and \g453245/U$2 ( \15308 , \8404 , RIfc99878_6769);
and \g453245/U$3 ( \15309 , RIfc8be80_6614, \8351 );
nor \g453245/U$1 ( \15310 , \15308 , \15309 );
and \g455275/U$2 ( \15311 , \8313 , RIfc480e0_5842);
and \g455275/U$3 ( \15312 , RIfc7fb08_6475, \8323 );
nor \g455275/U$1 ( \15313 , \15311 , \15312 );
not \g450291/U$3 ( \15314 , \15313 );
not \g450291/U$4 ( \15315 , \8328 );
and \g450291/U$2 ( \15316 , \15314 , \15315 );
and \g450291/U$5 ( \15317 , \8359 , RIfe97f38_8073);
nor \g450291/U$1 ( \15318 , \15316 , \15317 );
nand \g447870/U$1 ( \15319 , \15304 , \15307 , \15310 , \15318 );
nor \g446305/U$1 ( \15320 , \15299 , \15300 , \15319 );
and \g453244/U$2 ( \15321 , \8356 , RIee2deb0_4981);
and \g453244/U$3 ( \15322 , RIe141e88_2127, \8417 );
nor \g453244/U$1 ( \15323 , \15321 , \15322 );
and \g453243/U$2 ( \15324 , \8531 , RIee2eb58_4990);
and \g453243/U$3 ( \15325 , RIdf3da68_2078, \8414 );
nor \g453243/U$1 ( \15326 , \15324 , \15325 );
and \g445366/U$2 ( \15327 , \15320 , \15323 , \15326 );
nor \g445366/U$1 ( \15328 , \15327 , \8422 );
or \g444248/U$1 ( \15329 , \15268 , \15298 , \15328 );
_DC \g303c/U$1 ( \15330 , \15329 , \8654 );
and \g453152/U$2 ( \15331 , \8404 , RIe160ab8_2477);
and \g453152/U$3 ( \15332 , RIe15ddb8_2445, \8409 );
nor \g453152/U$1 ( \15333 , \15331 , \15332 );
and \g446287/U$2 ( \15334 , RIee37f00_5095, \8371 );
and \g446287/U$3 ( \15335 , RIe1556b8_2349, \8378 );
and \g449250/U$2 ( \15336 , RIe14a2b8_2221, \8317 );
and \g449250/U$3 ( \15337 , \8326 , RIe14cfb8_2253);
and \g449250/U$4 ( \15338 , RIe1637b8_2509, \8383 );
nor \g449250/U$1 ( \15339 , \15336 , \15337 , \15338 );
and \g453154/U$2 ( \15340 , \8335 , RIe1475b8_2189);
and \g453154/U$3 ( \15341 , RIfcbd368_7175, \8340 );
nor \g453154/U$1 ( \15342 , \15340 , \15341 );
and \g455264/U$2 ( \15343 , \8313 , RIfe9f990_8160);
and \g455264/U$3 ( \15344 , RIe1529b8_2317, \8323 );
nor \g455264/U$1 ( \15345 , \15343 , \15344 );
not \g450266/U$3 ( \15346 , \15345 );
not \g450266/U$4 ( \15347 , \8347 );
and \g450266/U$2 ( \15348 , \15346 , \15347 );
and \g450266/U$5 ( \15349 , \8351 , RIe1664b8_2541);
nor \g450266/U$1 ( \15350 , \15348 , \15349 );
and \g453153/U$2 ( \15351 , \8356 , RIe14fcb8_2285);
and \g453153/U$3 ( \15352 , RIfe9f828_8159, \8359 );
nor \g453153/U$1 ( \15353 , \15351 , \15352 );
nand \g447857/U$1 ( \15354 , \15339 , \15342 , \15350 , \15353 );
nor \g446287/U$1 ( \15355 , \15334 , \15335 , \15354 );
and \g453151/U$2 ( \15356 , \8414 , RIe1583b8_2381);
and \g453151/U$3 ( \15357 , RIfc8ea18_6645, \8417 );
nor \g453151/U$1 ( \15358 , \15356 , \15357 );
nand \g445647/U$1 ( \15359 , \15333 , \15355 , \15358 );
and \g444854/U$2 ( \15360 , \15359 , \8369 );
and \g449248/U$2 ( \15361 , RIfc98360_6754, \8373 );
and \g449248/U$3 ( \15362 , \8383 , RIfc45278_5809);
and \g449248/U$4 ( \15363 , RIee2ff08_5004, \8488 );
nor \g449248/U$1 ( \15364 , \15361 , \15362 , \15363 );
and \g454683/U$2 ( \15365 , \8313 , RIdf3d900_2077);
and \g454683/U$3 ( \15366 , RIe13f9f8_2101, \8323 );
nor \g454683/U$1 ( \15367 , \15365 , \15366 );
not \g450263/U$3 ( \15368 , \15367 );
not \g450263/U$4 ( \15369 , \8376 );
and \g450263/U$2 ( \15370 , \15368 , \15369 );
and \g450263/U$5 ( \15371 , \8359 , RIfcd6ca0_7466);
nor \g450263/U$1 ( \15372 , \15370 , \15371 );
and \g453145/U$2 ( \15373 , \8404 , RIfca2248_6867);
and \g453145/U$3 ( \15374 , RIfc8ee50_6648, \8351 );
nor \g453145/U$1 ( \15375 , \15373 , \15374 );
and \g453146/U$2 ( \15376 , \8378 , RIdf3b470_2051);
and \g453146/U$3 ( \15377 , RIe141d20_2126, \8417 );
nor \g453146/U$1 ( \15378 , \15376 , \15377 );
nand \g447855/U$1 ( \15379 , \15364 , \15372 , \15375 , \15378 );
and \g444854/U$3 ( \15380 , \9266 , \15379 );
nor \g444854/U$1 ( \15381 , \15360 , \15380 );
and \g447052/U$2 ( \15382 , \10230 , RIee2dd48_4980);
and \g447052/U$3 ( \15383 , RIfc8ece8_6647, \10232 );
nor \g447052/U$1 ( \15384 , \15382 , \15383 );
and \g447053/U$2 ( \15385 , \13424 , RIdf34120_1969);
and \g447053/U$3 ( \15386 , RIdf36718_1996, \13426 );
nor \g447053/U$1 ( \15387 , \15385 , \15386 );
and \g447054/U$2 ( \15388 , \9299 , RIfe9f6c0_8158);
and \g447054/U$3 ( \15389 , RIdf31f60_1945, \9301 );
nor \g447054/U$1 ( \15390 , \15388 , \15389 );
nand \g444642/U$1 ( \15391 , \15381 , \15384 , \15387 , \15390 );
and \g453160/U$2 ( \15392 , \8326 , RIdf20788_1746);
and \g453160/U$3 ( \15393 , RIfc7d678_6449, \8404 );
nor \g453160/U$1 ( \15394 , \15392 , \15393 );
and \g446290/U$2 ( \15395 , RIfc8e1a8_6639, \8371 );
and \g446290/U$3 ( \15396 , RIdf1b760_1689, \8319 );
and \g449253/U$2 ( \15397 , RIdf26e30_1819, \8414 );
and \g449253/U$3 ( \15398 , \8409 , RIdf28ff0_1843);
and \g449253/U$4 ( \15399 , RIfc45db8_5817, \8383 );
nor \g449253/U$1 ( \15400 , \15397 , \15398 , \15399 );
and \g453163/U$2 ( \15401 , \8356 , RIfcc2c00_7238);
and \g453163/U$3 ( \15402 , RIfcb43f8_7073, \8359 );
nor \g453163/U$1 ( \15403 , \15401 , \15402 );
and \g455271/U$2 ( \15404 , \8313 , RIdf23488_1778);
and \g455271/U$3 ( \15405 , RIfc8e748_6643, \8323 );
nor \g455271/U$1 ( \15406 , \15404 , \15405 );
not \g450269/U$3 ( \15407 , \15406 );
not \g450269/U$4 ( \15408 , \8347 );
and \g450269/U$2 ( \15409 , \15407 , \15408 );
and \g450269/U$5 ( \15410 , \8351 , RIfcb4560_7074);
nor \g450269/U$1 ( \15411 , \15409 , \15410 );
and \g453162/U$2 ( \15412 , \8378 , RIdf25378_1800);
and \g453162/U$3 ( \15413 , RIdf2aee0_1865, \8417 );
nor \g453162/U$1 ( \15414 , \15412 , \15413 );
nand \g447859/U$1 ( \15415 , \15400 , \15403 , \15411 , \15414 );
nor \g446290/U$1 ( \15416 , \15395 , \15396 , \15415 );
and \g453161/U$2 ( \15417 , \8335 , RIdf1a248_1674);
and \g453161/U$3 ( \15418 , RIdf21e08_1762, \8340 );
nor \g453161/U$1 ( \15419 , \15417 , \15418 );
nand \g445648/U$1 ( \15420 , \15394 , \15416 , \15419 );
and \g444728/U$2 ( \15421 , \15420 , \8752 );
and \g449252/U$2 ( \15422 , RIdef9188_1298, \8531 );
and \g449252/U$3 ( \15423 , \8488 , RIdefbe88_1330);
and \g449252/U$4 ( \15424 , RIdf15388_1618, \8383 );
nor \g449252/U$1 ( \15425 , \15422 , \15423 , \15424 );
and \g453157/U$2 ( \15426 , \8356 , RIdef6488_1266);
and \g453157/U$3 ( \15427 , RIdefeb88_1362, \8359 );
nor \g453157/U$1 ( \15428 , \15426 , \15427 );
and \g454600/U$2 ( \15429 , \8313 , RIdf07288_1458);
and \g454600/U$3 ( \15430 , RIdf09f88_1490, \8323 );
nor \g454600/U$1 ( \15431 , \15429 , \15430 );
not \g450267/U$3 ( \15432 , \15431 );
not \g450267/U$4 ( \15433 , \8376 );
and \g450267/U$2 ( \15434 , \15432 , \15433 );
and \g450267/U$5 ( \15435 , \8351 , RIdf18088_1650);
nor \g450267/U$1 ( \15436 , \15434 , \15435 );
and \g453156/U$2 ( \15437 , \8378 , RIdf04588_1426);
and \g453156/U$3 ( \15438 , RIdf0cc88_1522, \8417 );
nor \g453156/U$1 ( \15439 , \15437 , \15438 );
nand \g447858/U$1 ( \15440 , \15425 , \15428 , \15436 , \15439 );
and \g444728/U$3 ( \15441 , \8478 , \15440 );
nor \g444728/U$1 ( \15442 , \15421 , \15441 );
and \g447056/U$2 ( \15443 , \8780 , RIdef0a88_1202);
and \g447056/U$3 ( \15444 , RIdef3788_1234, \8782 );
nor \g447056/U$1 ( \15445 , \15443 , \15444 );
and \g447055/U$2 ( \15446 , \9480 , RIdf0f988_1554);
and \g447055/U$3 ( \15447 , RIdf12688_1586, \9482 );
nor \g447055/U$1 ( \15448 , \15446 , \15447 );
and \g447057/U$2 ( \15449 , \8785 , RIdeeb088_1138);
and \g447057/U$3 ( \15450 , RIdeedd88_1170, \8787 );
nor \g447057/U$1 ( \15451 , \15449 , \15450 );
nand \g444643/U$1 ( \15452 , \15442 , \15445 , \15448 , \15451 );
and \g446282/U$2 ( \15453 , RIfc98090_6752, \8531 );
and \g446282/U$3 ( \15454 , RIfe9fdc8_8163, \8319 );
and \g449243/U$2 ( \15455 , RIfc57860_6018, \8373 );
and \g449243/U$3 ( \15456 , \8383 , RIfc44e40_5806);
and \g449243/U$4 ( \15457 , RIee22678_4850, \8488 );
nor \g449243/U$1 ( \15458 , \15455 , \15456 , \15457 );
and \g455245/U$2 ( \15459 , \8313 , RIdee1740_1029);
and \g455245/U$3 ( \15460 , RIdee3900_1053, \8323 );
nor \g455245/U$1 ( \15461 , \15459 , \15460 );
not \g450260/U$3 ( \15462 , \15461 );
not \g450260/U$4 ( \15463 , \8376 );
and \g450260/U$2 ( \15464 , \15462 , \15463 );
and \g450260/U$5 ( \15465 , \8359 , RIfcbd4d0_7176);
nor \g450260/U$1 ( \15466 , \15464 , \15465 );
and \g453133/U$2 ( \15467 , \8404 , RIfca23b0_6868);
and \g453133/U$3 ( \15468 , RIfc8efb8_6649, \8351 );
nor \g453133/U$1 ( \15469 , \15467 , \15468 );
and \g453134/U$2 ( \15470 , \8378 , RIdedf6e8_1006);
and \g453134/U$3 ( \15471 , RIfe9faf8_8161, \8417 );
nor \g453134/U$1 ( \15472 , \15470 , \15471 );
nand \g447853/U$1 ( \15473 , \15458 , \15466 , \15469 , \15472 );
nor \g446282/U$1 ( \15474 , \15453 , \15454 , \15473 );
and \g453130/U$2 ( \15475 , \8335 , RIded3be0_873);
and \g453130/U$3 ( \15476 , RIfe9fc60_8162, \8340 );
nor \g453130/U$1 ( \15477 , \15475 , \15476 );
and \g453129/U$2 ( \15478 , \8326 , RIded80c8_922);
and \g453129/U$3 ( \15479 , RIee21598_4838, \8356 );
nor \g453129/U$1 ( \15480 , \15478 , \15479 );
and \g445352/U$2 ( \15481 , \15474 , \15477 , \15480 );
nor \g445352/U$1 ( \15482 , \15481 , \8481 );
and \g446284/U$2 ( \15483 , RIdecbeb8_784, \8371 );
and \g446284/U$3 ( \15484 , RIde7efc8_209, \8335 );
and \g449245/U$2 ( \15485 , RIdf2d910_1895, \8531 );
and \g449245/U$3 ( \15486 , \8488 , RIdf392b0_2027);
and \g449245/U$4 ( \15487 , RIdecebb8_816, \8383 );
nor \g449245/U$1 ( \15488 , \15485 , \15486 , \15487 );
and \g453141/U$2 ( \15489 , \8356 , RIdf1e190_1719);
and \g453141/U$3 ( \15490 , RIe1448b8_2157, \8359 );
nor \g453141/U$1 ( \15491 , \15489 , \15490 );
and \g455250/U$2 ( \15492 , \8313 , RIe16f2c0_2642);
and \g455250/U$3 ( \15493 , RIde99080_336, \8323 );
nor \g455250/U$1 ( \15494 , \15492 , \15493 );
not \g450262/U$3 ( \15495 , \15494 );
not \g450262/U$4 ( \15496 , \8376 );
and \g450262/U$2 ( \15497 , \15495 , \15496 );
and \g450262/U$5 ( \15498 , \8351 , RIded18b8_848);
nor \g450262/U$1 ( \15499 , \15497 , \15498 );
and \g453139/U$2 ( \15500 , \8378 , RIe15b0b8_2413);
and \g453139/U$3 ( \15501 , RIdeb56b8_528, \8417 );
nor \g453139/U$1 ( \15502 , \15500 , \15501 );
nand \g447854/U$1 ( \15503 , \15488 , \15491 , \15499 , \15502 );
nor \g446284/U$1 ( \15504 , \15483 , \15484 , \15503 );
and \g453136/U$2 ( \15505 , \8340 , RIdf01888_1394);
and \g453136/U$3 ( \15506 , RIdec91b8_752, \8404 );
nor \g453136/U$1 ( \15507 , \15505 , \15506 );
and \g453138/U$2 ( \15508 , \8317 , RIdedd0f0_979);
and \g453138/U$3 ( \15509 , RIdee8388_1106, \8326 );
nor \g453138/U$1 ( \15510 , \15508 , \15509 );
and \g445354/U$2 ( \15511 , \15504 , \15507 , \15510 );
nor \g445354/U$1 ( \15512 , \15511 , \8651 );
or \g444327/U$1 ( \15513 , \15391 , \15452 , \15482 , \15512 );
and \g446279/U$2 ( \15514 , RIfc8daa0_6634, \8373 );
and \g446279/U$3 ( \15515 , RIdebb0b8_592, \8414 );
and \g449239/U$2 ( \15516 , RIfcbd098_7173, \8523 );
and \g449239/U$3 ( \15517 , \8488 , RIdeb29b8_496);
and \g449239/U$4 ( \15518 , RIdec37b8_688, \8383 );
nor \g449239/U$1 ( \15519 , \15516 , \15517 , \15518 );
and \g453118/U$2 ( \15520 , \8335 , RIde9f980_368);
and \g453118/U$3 ( \15521 , RIfc8dc08_6635, \8340 );
nor \g453118/U$1 ( \15522 , \15520 , \15521 );
and \g455233/U$2 ( \15523 , \8313 , RIdea6280_400);
and \g455233/U$3 ( \15524 , RIdeacb80_432, \8323 );
nor \g455233/U$1 ( \15525 , \15523 , \15524 );
not \g455232/U$1 ( \15526 , \15525 );
and \g450255/U$2 ( \15527 , \15526 , \8316 );
and \g450255/U$3 ( \15528 , RIdec64b8_720, \8351 );
nor \g450255/U$1 ( \15529 , \15527 , \15528 );
and \g453116/U$2 ( \15530 , \8356 , RIdeafcb8_464);
and \g453116/U$3 ( \15531 , RIfc98798_6757, \8359 );
nor \g453116/U$1 ( \15532 , \15530 , \15531 );
nand \g448217/U$1 ( \15533 , \15519 , \15522 , \15529 , \15532 );
nor \g446279/U$1 ( \15534 , \15514 , \15515 , \15533 );
and \g453113/U$2 ( \15535 , \8404 , RIdec0ab8_656);
and \g453113/U$3 ( \15536 , RIfc56348_6003, \8417 );
nor \g453113/U$1 ( \15537 , \15535 , \15536 );
and \g453114/U$2 ( \15538 , \8378 , RIdeb83b8_560);
and \g453114/U$3 ( \15539 , RIdebddb8_624, \8409 );
nor \g453114/U$1 ( \15540 , \15538 , \15539 );
and \g445350/U$2 ( \15541 , \15534 , \15537 , \15540 );
nor \g445350/U$1 ( \15542 , \15541 , \8589 );
and \g446280/U$2 ( \15543 , RIfc7dd80_6454, \8373 );
and \g446280/U$3 ( \15544 , RIde86fc0_248, \8378 );
and \g449241/U$2 ( \15545 , RIfcd96d0_7496, \8531 );
and \g449241/U$3 ( \15546 , \8488 , RIfc8e040_6638);
and \g449241/U$4 ( \15547 , RIfc8ded8_6637, \8383 );
nor \g449241/U$1 ( \15548 , \15545 , \15546 , \15547 );
and \g453126/U$2 ( \15549 , \8335 , RIe168ab0_2568);
and \g453126/U$3 ( \15550 , RIfcbd200_7174, \8340 );
nor \g453126/U$1 ( \15551 , \15549 , \15550 );
and \g454537/U$2 ( \15552 , \8313 , RIe16a298_2585);
and \g454537/U$3 ( \15553 , RIe16c5c0_2610, \8323 );
nor \g454537/U$1 ( \15554 , \15552 , \15553 );
not \g454536/U$1 ( \15555 , \15554 );
and \g450258/U$2 ( \15556 , \15555 , \8316 );
and \g450258/U$3 ( \15557 , RIfcd6868_7463, \8351 );
nor \g450258/U$1 ( \15558 , \15556 , \15557 );
and \g453125/U$2 ( \15559 , \8356 , RIfca1e10_6864);
and \g453125/U$3 ( \15560 , RIde82ad8_227, \8359 );
nor \g453125/U$1 ( \15561 , \15559 , \15560 );
nand \g448218/U$1 ( \15562 , \15548 , \15551 , \15558 , \15561 );
nor \g446280/U$1 ( \15563 , \15543 , \15544 , \15562 );
and \g453124/U$2 ( \15564 , \8404 , RIfc56618_6005);
and \g453124/U$3 ( \15565 , RIde8f300_288, \8409 );
nor \g453124/U$1 ( \15566 , \15564 , \15565 );
and \g453122/U$2 ( \15567 , \8412 , RIde8b160_268);
and \g453122/U$3 ( \15568 , RIde92e10_306, \8417 );
nor \g453122/U$1 ( \15569 , \15567 , \15568 );
and \g445351/U$2 ( \15570 , \15563 , \15566 , \15569 );
nor \g445351/U$1 ( \15571 , \15570 , \8558 );
or \g444282/U$1 ( \15572 , \15513 , \15542 , \15571 );
_DC \g30c1/U$1 ( \15573 , \15572 , \8654 );
and \g448655/U$2 ( \15574 , RIe157f80_2378, \8414 );
and \g448655/U$3 ( \15575 , \8407 , RIe15d980_2442);
and \g448655/U$4 ( \15576 , RIe152580_2314, \8486 );
nor \g448655/U$1 ( \15577 , \15574 , \15575 , \15576 );
and \g454392/U$2 ( \15578 , \8313 , RIee37ac8_5092);
and \g454392/U$3 ( \15579 , RIe163380_2506, \8323 );
nor \g454392/U$1 ( \15580 , \15578 , \15579 );
not \g449680/U$3 ( \15581 , \15580 );
not \g449680/U$4 ( \15582 , \8328 );
and \g449680/U$2 ( \15583 , \15581 , \15582 );
and \g449680/U$5 ( \15584 , \8359 , RIfc3f530_5746);
nor \g449680/U$1 ( \15585 , \15583 , \15584 );
and \g451136/U$2 ( \15586 , \8404 , RIe160680_2474);
and \g451136/U$3 ( \15587 , RIe166080_2538, \8351 );
nor \g451136/U$1 ( \15588 , \15586 , \15587 );
and \g451138/U$2 ( \15589 , \8378 , RIe155280_2346);
and \g451138/U$3 ( \15590 , RIfcd1c78_7409, \8417 );
nor \g451138/U$1 ( \15591 , \15589 , \15590 );
nand \g447547/U$1 ( \15592 , \15577 , \15585 , \15588 , \15591 );
and \g444758/U$2 ( \15593 , \15592 , \8369 );
and \g445830/U$2 ( \15594 , RIfc5a560_6050, \8373 );
and \g445830/U$3 ( \15595 , RIdf3d4c8_2074, \8414 );
and \g448657/U$2 ( \15596 , RIdf31c90_1943, \8317 );
and \g448657/U$3 ( \15597 , \8326 , RIdf33e50_1967);
and \g448657/U$4 ( \15598 , RIfc7a270_6412, \8330 );
nor \g448657/U$1 ( \15599 , \15596 , \15597 , \15598 );
and \g451146/U$2 ( \15600 , \8335 , RIdf2fda0_1921);
and \g451146/U$3 ( \15601 , RIdf362e0_1993, \8340 );
nor \g451146/U$1 ( \15602 , \15600 , \15601 );
and \g455361/U$2 ( \15603 , \8313 , RIfc91cb8_6681);
and \g455361/U$3 ( \15604 , RIee2fc38_5002, \8323 );
nor \g455361/U$1 ( \15605 , \15603 , \15604 );
not \g449682/U$3 ( \15606 , \15605 );
not \g449682/U$4 ( \15607 , \8347 );
and \g449682/U$2 ( \15608 , \15606 , \15607 );
and \g449682/U$5 ( \15609 , \8351 , RIfc42b18_5781);
nor \g449682/U$1 ( \15610 , \15608 , \15609 );
and \g451145/U$2 ( \15611 , \8356 , RIee2d910_4977);
and \g451145/U$3 ( \15612 , RIfce5bb0_7636, \8359 );
nor \g451145/U$1 ( \15613 , \15611 , \15612 );
nand \g447549/U$1 ( \15614 , \15599 , \15602 , \15610 , \15613 );
nor \g445830/U$1 ( \15615 , \15594 , \15595 , \15614 );
and \g451142/U$2 ( \15616 , \8404 , RIfc96b78_6737);
and \g451142/U$3 ( \15617 , RIfea6fb0_8216, \8417 );
nor \g451142/U$1 ( \15618 , \15616 , \15617 );
and \g451143/U$2 ( \15619 , \8378 , RIdf3b038_2048);
and \g451143/U$3 ( \15620 , RIe13f5c0_2098, \8409 );
nor \g451143/U$1 ( \15621 , \15619 , \15620 );
and \g445023/U$2 ( \15622 , \15615 , \15618 , \15621 );
nor \g445023/U$1 ( \15623 , \15622 , \8422 );
nor \g444758/U$1 ( \15624 , \15593 , \15623 );
and \g446621/U$2 ( \15625 , \8707 , RIe147180_2186);
and \g446621/U$3 ( \15626 , RIe149e80_2218, \8709 );
nor \g446621/U$1 ( \15627 , \15625 , \15626 );
and \g446620/U$2 ( \15628 , \8712 , RIe14cb80_2250);
and \g446620/U$3 ( \15629 , RIfc7a3d8_6413, \8714 );
nor \g446620/U$1 ( \15630 , \15628 , \15629 );
and \g446622/U$2 ( \15631 , \8717 , RIe14f880_2282);
and \g446622/U$3 ( \15632 , RIee35368_5064, \8719 );
nor \g446622/U$1 ( \15633 , \15631 , \15632 );
nand \g444461/U$1 ( \15634 , \15624 , \15627 , \15630 , \15633 );
and \g451156/U$2 ( \15635 , \8414 , RIe16ee88_2639);
and \g451156/U$3 ( \15636 , RIde986a8_333, \8409 );
nor \g451156/U$1 ( \15637 , \15635 , \15636 );
and \g445831/U$2 ( \15638 , RIdeb5280_525, \8417 );
and \g445831/U$3 ( \15639 , RIdec8d80_749, \8404 );
and \g448661/U$2 ( \15640 , RIdedccb8_976, \8317 );
and \g448661/U$3 ( \15641 , \8326 , RIdee7f50_1103);
and \g448661/U$4 ( \15642 , RIdece780_813, \8383 );
nor \g448661/U$1 ( \15643 , \15640 , \15641 , \15642 );
and \g451159/U$2 ( \15644 , \8335 , RIde7e5f0_206);
and \g451159/U$3 ( \15645 , RIdf01450_1391, \8340 );
nor \g451159/U$1 ( \15646 , \15644 , \15645 );
and \g454395/U$2 ( \15647 , \8313 , RIdf2d4d8_1892);
and \g454395/U$3 ( \15648 , RIdf38e78_2024, \8323 );
nor \g454395/U$1 ( \15649 , \15647 , \15648 );
not \g449688/U$3 ( \15650 , \15649 );
not \g449688/U$4 ( \15651 , \8347 );
and \g449688/U$2 ( \15652 , \15650 , \15651 );
and \g449688/U$5 ( \15653 , \8351 , RIded1480_845);
nor \g449688/U$1 ( \15654 , \15652 , \15653 );
and \g451158/U$2 ( \15655 , \8356 , RIdf1dd58_1716);
and \g451158/U$3 ( \15656 , RIe144480_2154, \8359 );
nor \g451158/U$1 ( \15657 , \15655 , \15656 );
nand \g447552/U$1 ( \15658 , \15643 , \15646 , \15654 , \15657 );
nor \g445831/U$1 ( \15659 , \15638 , \15639 , \15658 );
and \g451157/U$2 ( \15660 , \8378 , RIe15ac80_2410);
and \g451157/U$3 ( \15661 , RIdecba80_781, \8371 );
nor \g451157/U$1 ( \15662 , \15660 , \15661 );
nand \g445535/U$1 ( \15663 , \15637 , \15659 , \15662 );
and \g444874/U$2 ( \15664 , \15663 , \9010 );
and \g448658/U$2 ( \15665 , RIfc7a978_6417, \8319 );
and \g448658/U$3 ( \15666 , \8326 , RIdf20350_1743);
and \g448658/U$4 ( \15667 , RIfc59e58_6045, \8383 );
nor \g448658/U$1 ( \15668 , \15665 , \15666 , \15667 );
and \g451153/U$2 ( \15669 , \8335 , RIdf19e10_1671);
and \g451153/U$3 ( \15670 , RIfc430b8_5785, \8340 );
nor \g451153/U$1 ( \15671 , \15669 , \15670 );
and \g454913/U$2 ( \15672 , \8313 , RIfc919e8_6679);
and \g454913/U$3 ( \15673 , RIfcb3318_7061, \8323 );
nor \g454913/U$1 ( \15674 , \15672 , \15673 );
not \g449683/U$3 ( \15675 , \15674 );
not \g449683/U$4 ( \15676 , \8347 );
and \g449683/U$2 ( \15677 , \15675 , \15676 );
and \g449683/U$5 ( \15678 , \8351 , RIfc43658_5789);
nor \g449683/U$1 ( \15679 , \15677 , \15678 );
and \g451152/U$2 ( \15680 , \8356 , RIfc91880_6678);
and \g451152/U$3 ( \15681 , RIfc91718_6677, \8359 );
nor \g451152/U$1 ( \15682 , \15680 , \15681 );
nand \g447551/U$1 ( \15683 , \15668 , \15671 , \15679 , \15682 );
and \g444874/U$3 ( \15684 , \8752 , \15683 );
nor \g444874/U$1 ( \15685 , \15664 , \15684 );
and \g446625/U$2 ( \15686 , \11511 , RIfc7ac48_6419);
and \g446625/U$3 ( \15687 , RIfc96fb0_6740, \11513 );
nor \g446625/U$1 ( \15688 , \15686 , \15687 );
and \g446624/U$2 ( \15689 , \11516 , RIdf28bb8_1840);
and \g446624/U$3 ( \15690 , RIfea0368_8167, \11518 );
nor \g446624/U$1 ( \15691 , \15689 , \15690 );
and \g446626/U$2 ( \15692 , \11521 , RIdf25210_1799);
and \g446626/U$3 ( \15693 , RIdf26cc8_1818, \11523 );
nor \g446626/U$1 ( \15694 , \15692 , \15693 );
nand \g444568/U$1 ( \15695 , \15685 , \15688 , \15691 , \15694 );
and \g445826/U$2 ( \15696 , RIdef6050_1263, \8356 );
and \g445826/U$3 ( \15697 , RIdef3350_1231, \8340 );
and \g448652/U$2 ( \15698 , RIdf12250_1583, \8373 );
and \g448652/U$3 ( \15699 , \8383 , RIdf14f50_1615);
and \g448652/U$4 ( \15700 , RIdefba50_1327, \8488 );
nor \g448652/U$1 ( \15701 , \15698 , \15699 , \15700 );
and \g454383/U$2 ( \15702 , \8313 , RIdf06e50_1455);
and \g454383/U$3 ( \15703 , RIdf09b50_1487, \8323 );
nor \g454383/U$1 ( \15704 , \15702 , \15703 );
not \g449677/U$3 ( \15705 , \15704 );
not \g449677/U$4 ( \15706 , \8376 );
and \g449677/U$2 ( \15707 , \15705 , \15706 );
and \g449677/U$5 ( \15708 , \8359 , RIdefe750_1359);
nor \g449677/U$1 ( \15709 , \15707 , \15708 );
and \g451126/U$2 ( \15710 , \8404 , RIdf0f550_1551);
and \g451126/U$3 ( \15711 , RIdf17c50_1647, \8351 );
nor \g451126/U$1 ( \15712 , \15710 , \15711 );
and \g451128/U$2 ( \15713 , \8378 , RIdf04150_1423);
and \g451128/U$3 ( \15714 , RIdf0c850_1519, \8417 );
nor \g451128/U$1 ( \15715 , \15713 , \15714 );
nand \g447544/U$1 ( \15716 , \15701 , \15709 , \15712 , \15715 );
nor \g445826/U$1 ( \15717 , \15696 , \15697 , \15716 );
and \g451124/U$2 ( \15718 , \8335 , RIdeeac50_1135);
and \g451124/U$3 ( \15719 , RIdef8d50_1295, \8531 );
nor \g451124/U$1 ( \15720 , \15718 , \15719 );
and \g451123/U$2 ( \15721 , \8319 , RIdeed950_1167);
and \g451123/U$3 ( \15722 , RIdef0650_1199, \8324 );
nor \g451123/U$1 ( \15723 , \15721 , \15722 );
and \g445020/U$2 ( \15724 , \15717 , \15720 , \15723 );
nor \g445020/U$1 ( \15725 , \15724 , \8477 );
and \g445827/U$2 ( \15726 , RIfc5a830_6052, \8356 );
and \g445827/U$3 ( \15727 , RIdeda3f0_947, \8340 );
and \g448654/U$2 ( \15728 , RIdee1308_1026, \8412 );
and \g448654/U$3 ( \15729 , \8409 , RIdee3630_1051);
and \g448654/U$4 ( \15730 , RIfcd85f0_7484, \8488 );
nor \g448654/U$1 ( \15731 , \15728 , \15729 , \15730 );
and \g455038/U$2 ( \15732 , \8313 , RIfc91f88_6683);
and \g455038/U$3 ( \15733 , RIfc968a8_6735, \8323 );
nor \g455038/U$1 ( \15734 , \15732 , \15733 );
not \g449679/U$3 ( \15735 , \15734 );
not \g449679/U$4 ( \15736 , \8328 );
and \g449679/U$2 ( \15737 , \15735 , \15736 );
and \g449679/U$5 ( \15738 , \8359 , RIfcc7d90_7296);
nor \g449679/U$1 ( \15739 , \15737 , \15738 );
and \g451132/U$2 ( \15740 , \8404 , RIfcdfc10_7568);
and \g451132/U$3 ( \15741 , RIfcd1b10_7408, \8351 );
nor \g451132/U$1 ( \15742 , \15740 , \15741 );
and \g451133/U$2 ( \15743 , \8378 , RIdedf2b0_1003);
and \g451133/U$3 ( \15744 , RIfea99e0_8246, \8417 );
nor \g451133/U$1 ( \15745 , \15743 , \15744 );
nand \g447545/U$1 ( \15746 , \15731 , \15739 , \15742 , \15745 );
nor \g445827/U$1 ( \15747 , \15726 , \15727 , \15746 );
and \g451131/U$2 ( \15748 , \8335 , RIded37a8_870);
and \g451131/U$3 ( \15749 , RIfce3888_7611, \8531 );
nor \g451131/U$1 ( \15750 , \15748 , \15749 );
and \g451130/U$2 ( \15751 , \8319 , RIded5f08_898);
and \g451130/U$3 ( \15752 , RIfea9878_8245, \8326 );
nor \g451130/U$1 ( \15753 , \15751 , \15752 );
and \g445021/U$2 ( \15754 , \15747 , \15750 , \15753 );
nor \g445021/U$1 ( \15755 , \15754 , \8481 );
or \g444335/U$1 ( \15756 , \15634 , \15695 , \15725 , \15755 );
and \g445823/U$2 ( \15757 , RIfcd70d8_7469, \8417 );
and \g445823/U$3 ( \15758 , RIdec0680_653, \8404 );
and \g448649/U$2 ( \15759 , RIdea58a8_397, \8319 );
and \g448649/U$3 ( \15760 , \8326 , RIdeac1a8_429);
and \g448649/U$4 ( \15761 , RIdec3380_685, \8383 );
nor \g448649/U$1 ( \15762 , \15759 , \15760 , \15761 );
and \g451115/U$2 ( \15763 , \8335 , RIde9efa8_365);
and \g451115/U$3 ( \15764 , RIfc43928_5791, \8340 );
nor \g451115/U$1 ( \15765 , \15763 , \15764 );
and \g454377/U$2 ( \15766 , \8313 , RIfcb3480_7062);
and \g454377/U$3 ( \15767 , RIdeb2580_493, \8323 );
nor \g454377/U$1 ( \15768 , \15766 , \15767 );
not \g449674/U$3 ( \15769 , \15768 );
not \g449674/U$4 ( \15770 , \8347 );
and \g449674/U$2 ( \15771 , \15769 , \15770 );
and \g449674/U$5 ( \15772 , \8351 , RIdec6080_717);
nor \g449674/U$1 ( \15773 , \15771 , \15772 );
and \g451113/U$2 ( \15774 , \8356 , RIdeaf880_461);
and \g451113/U$3 ( \15775 , RIfcbe448_7187, \8359 );
nor \g451113/U$1 ( \15776 , \15774 , \15775 );
nand \g447540/U$1 ( \15777 , \15762 , \15765 , \15773 , \15776 );
nor \g445823/U$1 ( \15778 , \15757 , \15758 , \15777 );
and \g451111/U$2 ( \15779 , \8378 , RIdeb7f80_557);
and \g451111/U$3 ( \15780 , RIee204b8_4826, \8371 );
nor \g451111/U$1 ( \15781 , \15779 , \15780 );
and \g451110/U$2 ( \15782 , \8414 , RIdebac80_589);
and \g451110/U$3 ( \15783 , RIdebd980_621, \8409 );
nor \g451110/U$1 ( \15784 , \15782 , \15783 );
and \g445018/U$2 ( \15785 , \15778 , \15781 , \15784 );
nor \g445018/U$1 ( \15786 , \15785 , \8589 );
and \g445824/U$2 ( \15787 , RIfcd1de0_7410, \8523 );
and \g445824/U$3 ( \15788 , RIfc97118_6741, \8317 );
and \g448650/U$2 ( \15789 , RIfcc77f0_7292, \8371 );
and \g448650/U$3 ( \15790 , \8330 , RIee1c408_4780);
and \g448650/U$4 ( \15791 , RIfc59a20_6042, \8488 );
nor \g448650/U$1 ( \15792 , \15789 , \15790 , \15791 );
and \g455159/U$2 ( \15793 , \8313 , RIde8aad0_266);
and \g455159/U$3 ( \15794 , RIde8ec70_286, \8323 );
nor \g455159/U$1 ( \15795 , \15793 , \15794 );
not \g449676/U$3 ( \15796 , \15795 );
not \g449676/U$4 ( \15797 , \8376 );
and \g449676/U$2 ( \15798 , \15796 , \15797 );
and \g449676/U$5 ( \15799 , \8359 , RIfca31c0_6878);
nor \g449676/U$1 ( \15800 , \15798 , \15799 );
and \g451119/U$2 ( \15801 , \8404 , RIfea04d0_8168);
and \g451119/U$3 ( \15802 , RIfcd88c0_7486, \8351 );
nor \g451119/U$1 ( \15803 , \15801 , \15802 );
and \g451121/U$2 ( \15804 , \8378 , RIde86930_246);
and \g451121/U$3 ( \15805 , RIde92438_303, \8417 );
nor \g451121/U$1 ( \15806 , \15804 , \15805 );
nand \g447541/U$1 ( \15807 , \15792 , \15800 , \15803 , \15806 );
nor \g445824/U$1 ( \15808 , \15787 , \15788 , \15807 );
and \g451118/U$2 ( \15809 , \8335 , RIe168948_2567);
and \g451118/U$3 ( \15810 , RIfc97280_6742, \8340 );
nor \g451118/U$1 ( \15811 , \15809 , \15810 );
and \g451116/U$2 ( \15812 , \8326 , RIe16c188_2607);
and \g451116/U$3 ( \15813 , RIfc91448_6675, \8356 );
nor \g451116/U$1 ( \15814 , \15812 , \15813 );
and \g445019/U$2 ( \15815 , \15808 , \15811 , \15814 );
nor \g445019/U$1 ( \15816 , \15815 , \8558 );
or \g444268/U$1 ( \15817 , \15756 , \15786 , \15816 );
_DC \g3146/U$1 ( \15818 , \15817 , \8654 );
and \g448935/U$2 ( \15819 , RIfea8ea0_8238, \8414 );
and \g448935/U$3 ( \15820 , \8409 , RIde8d578_279);
and \g448935/U$4 ( \15821 , RIfc938d8_6701, \8486 );
nor \g448935/U$1 ( \15822 , \15819 , \15820 , \15821 );
and \g454980/U$2 ( \15823 , \8313 , RIee1b328_4768);
and \g454980/U$3 ( \15824 , RIee1bb98_4774, \8323 );
nor \g454980/U$1 ( \15825 , \15823 , \15824 );
not \g449949/U$3 ( \15826 , \15825 );
not \g449949/U$4 ( \15827 , \8328 );
and \g449949/U$2 ( \15828 , \15826 , \15827 );
and \g449949/U$5 ( \15829 , \8359 , RIde813e0_220);
nor \g449949/U$1 ( \15830 , \15828 , \15829 );
and \g452023/U$2 ( \15831 , \8404 , RIee1aab8_4762);
and \g452023/U$3 ( \15832 , RIee1cc78_4786, \8351 );
nor \g452023/U$1 ( \15833 , \15831 , \15832 );
and \g452024/U$2 ( \15834 , \8378 , RIde85238_239);
and \g452024/U$3 ( \15835 , RIde909f8_295, \8417 );
nor \g452024/U$1 ( \15836 , \15834 , \15835 );
nand \g447693/U$1 ( \15837 , \15822 , \15830 , \15833 , \15836 );
and \g444685/U$2 ( \15838 , \15837 , \9700 );
and \g446044/U$2 ( \15839 , RIfc78218_6389, \8523 );
and \g446044/U$3 ( \15840 , RIde9cb90_354, \8335 );
and \g448904/U$2 ( \15841 , RIdeb9d08_578, \8414 );
and \g448904/U$3 ( \15842 , \8409 , RIdebca08_610);
and \g448904/U$4 ( \15843 , RIdeb1608_482, \8488 );
nor \g448904/U$1 ( \15844 , \15841 , \15842 , \15843 );
and \g454379/U$2 ( \15845 , \8313 , RIfc93608_6699);
and \g454379/U$3 ( \15846 , RIdec2408_674, \8323 );
nor \g454379/U$1 ( \15847 , \15845 , \15846 );
not \g449951/U$3 ( \15848 , \15847 );
not \g449951/U$4 ( \15849 , \8328 );
and \g449951/U$2 ( \15850 , \15848 , \15849 );
and \g449951/U$5 ( \15851 , \8359 , RIfcdf7d8_7565);
nor \g449951/U$1 ( \15852 , \15850 , \15851 );
and \g452403/U$2 ( \15853 , \8404 , RIdebf708_642);
and \g452403/U$3 ( \15854 , RIdec5108_706, \8351 );
nor \g452403/U$1 ( \15855 , \15853 , \15854 );
and \g452029/U$2 ( \15856 , \8378 , RIdeb7008_546);
and \g452029/U$3 ( \15857 , RIfc934a0_6698, \8417 );
nor \g452029/U$1 ( \15858 , \15856 , \15857 );
nand \g447694/U$1 ( \15859 , \15844 , \15852 , \15855 , \15858 );
nor \g446044/U$1 ( \15860 , \15839 , \15840 , \15859 );
and \g452025/U$2 ( \15861 , \8356 , RIdeae908_450);
and \g452025/U$3 ( \15862 , RIfcc8498_7301, \8340 );
nor \g452025/U$1 ( \15863 , \15861 , \15862 );
and \g452026/U$2 ( \15864 , \8319 , RIdea3490_386);
and \g452026/U$3 ( \15865 , RIdea9d90_418, \8326 );
nor \g452026/U$1 ( \15866 , \15864 , \15865 );
and \g445184/U$2 ( \15867 , \15860 , \15863 , \15866 );
nor \g445184/U$1 ( \15868 , \15867 , \8589 );
nor \g444685/U$1 ( \15869 , \15838 , \15868 );
and \g446827/U$2 ( \15870 , \10044 , RIfea9f80_8250);
and \g446827/U$3 ( \15871 , RIfea8d38_8237, \10046 );
nor \g446827/U$1 ( \15872 , \15870 , \15871 );
and \g446826/U$2 ( \15873 , \10034 , RIe16b4e0_2598);
and \g446826/U$3 ( \15874 , RIfce8ce8_7671, \10036 );
nor \g446826/U$1 ( \15875 , \15873 , \15874 );
and \g446828/U$2 ( \15876 , \12264 , RIfcbfd98_7205);
and \g446828/U$3 ( \15877 , RIfce5e80_7638, \12266 );
nor \g446828/U$1 ( \15878 , \15876 , \15877 );
nand \g444490/U$1 ( \15879 , \15869 , \15872 , \15875 , \15878 );
and \g452033/U$2 ( \15880 , \8317 , RIdeec9d8_1156);
and \g452033/U$3 ( \15881 , RIdeef6d8_1188, \8326 );
nor \g452033/U$1 ( \15882 , \15880 , \15881 );
and \g446046/U$2 ( \15883 , RIdef7dd8_1284, \8523 );
and \g446046/U$3 ( \15884 , RIdee9cd8_1124, \8335 );
and \g448940/U$2 ( \15885 , RIdf112d8_1572, \8373 );
and \g448940/U$3 ( \15886 , \8383 , RIdf13fd8_1604);
and \g448940/U$4 ( \15887 , RIdefaad8_1316, \8486 );
nor \g448940/U$1 ( \15888 , \15885 , \15886 , \15887 );
and \g454663/U$2 ( \15889 , \8313 , RIdf05ed8_1444);
and \g454663/U$3 ( \15890 , RIdf08bd8_1476, \8323 );
nor \g454663/U$1 ( \15891 , \15889 , \15890 );
not \g449953/U$3 ( \15892 , \15891 );
not \g449953/U$4 ( \15893 , \8376 );
and \g449953/U$2 ( \15894 , \15892 , \15893 );
and \g449953/U$5 ( \15895 , \8359 , RIdefd7d8_1348);
nor \g449953/U$1 ( \15896 , \15894 , \15895 );
and \g452035/U$2 ( \15897 , \8404 , RIdf0e5d8_1540);
and \g452035/U$3 ( \15898 , RIdf16cd8_1636, \8351 );
nor \g452035/U$1 ( \15899 , \15897 , \15898 );
and \g452036/U$2 ( \15900 , \8378 , RIdf031d8_1412);
and \g452036/U$3 ( \15901 , RIdf0b8d8_1508, \8417 );
nor \g452036/U$1 ( \15902 , \15900 , \15901 );
nand \g447697/U$1 ( \15903 , \15888 , \15896 , \15899 , \15902 );
nor \g446046/U$1 ( \15904 , \15883 , \15884 , \15903 );
and \g452034/U$2 ( \15905 , \8356 , RIdef50d8_1252);
and \g452034/U$3 ( \15906 , RIdef23d8_1220, \8340 );
nor \g452034/U$1 ( \15907 , \15905 , \15906 );
nand \g445585/U$1 ( \15908 , \15882 , \15904 , \15907 );
and \g444773/U$2 ( \15909 , \15908 , \8478 );
and \g448938/U$2 ( \15910 , RIfcc8768_7303, \8531 );
and \g448938/U$3 ( \15911 , \8488 , RIee22240_4847);
and \g448938/U$4 ( \15912 , RIfcde6f8_7553, \8383 );
nor \g448938/U$1 ( \15913 , \15910 , \15911 , \15912 );
and \g452065/U$2 ( \15914 , \8335 , RIfea76b8_8221);
and \g452065/U$3 ( \15915 , RIded95e0_937, \8340 );
nor \g452065/U$1 ( \15916 , \15914 , \15915 );
and \g454429/U$2 ( \15917 , \8313 , RIded5260_889);
and \g454429/U$3 ( \15918 , RIded7150_911, \8323 );
nor \g454429/U$1 ( \15919 , \15917 , \15918 );
not \g454428/U$1 ( \15920 , \15919 );
and \g449952/U$2 ( \15921 , \15920 , \8316 );
and \g449952/U$3 ( \15922 , RIfc942b0_6708, \8351 );
nor \g449952/U$1 ( \15923 , \15921 , \15922 );
and \g451941/U$2 ( \15924 , \8356 , RIee21160_4835);
and \g451941/U$3 ( \15925 , RIfc5c9f0_6076, \8359 );
nor \g451941/U$1 ( \15926 , \15924 , \15925 );
nand \g448185/U$1 ( \15927 , \15913 , \15916 , \15923 , \15926 );
and \g444773/U$3 ( \15928 , \8482 , \15927 );
nor \g444773/U$1 ( \15929 , \15909 , \15928 );
and \g446831/U$2 ( \15930 , \8964 , RIdee2af0_1043);
and \g446831/U$3 ( \15931 , RIdee4878_1064, \8966 );
nor \g446831/U$1 ( \15932 , \15930 , \15931 );
and \g446832/U$2 ( \15933 , \8969 , RIfcde860_7554);
and \g446832/U$3 ( \15934 , RIfcd1138_7401, \8971 );
nor \g446832/U$1 ( \15935 , \15933 , \15934 );
and \g446833/U$2 ( \15936 , \8974 , RIdede8d8_996);
and \g446833/U$3 ( \15937 , RIdee0a98_1020, \8976 );
nor \g446833/U$1 ( \15938 , \15936 , \15937 );
nand \g444491/U$1 ( \15939 , \15929 , \15932 , \15935 , \15938 );
and \g446040/U$2 ( \15940 , RIfc93fe0_6706, \8356 );
and \g446040/U$3 ( \15941 , RIdf354d0_1983, \8340 );
and \g448932/U$2 ( \15942 , RIfc93e78_6705, \8373 );
and \g448932/U$3 ( \15943 , \8383 , RIfcb19c8_7043);
and \g448932/U$4 ( \15944 , RIfcdbf98_7525, \8486 );
nor \g448932/U$1 ( \15945 , \15942 , \15943 , \15944 );
and \g454516/U$2 ( \15946 , \8313 , RIdf3c988_2066);
and \g454516/U$3 ( \15947 , RIdf3ecb0_2091, \8323 );
nor \g454516/U$1 ( \15948 , \15946 , \15947 );
not \g449946/U$3 ( \15949 , \15948 );
not \g449946/U$4 ( \15950 , \8376 );
and \g449946/U$2 ( \15951 , \15949 , \15950 );
and \g449946/U$5 ( \15952 , \8359 , RIfce8478_7665);
nor \g449946/U$1 ( \15953 , \15951 , \15952 );
and \g452014/U$2 ( \15954 , \8404 , RIfce7938_7657);
and \g452014/U$3 ( \15955 , RIfceb718_7701, \8351 );
nor \g452014/U$1 ( \15956 , \15954 , \15955 );
and \g453770/U$2 ( \15957 , \8378 , RIfe9daa0_8138);
and \g453770/U$3 ( \15958 , RIe140da8_2115, \8417 );
nor \g453770/U$1 ( \15959 , \15957 , \15958 );
nand \g447689/U$1 ( \15960 , \15945 , \15953 , \15956 , \15959 );
nor \g446040/U$1 ( \15961 , \15940 , \15941 , \15960 );
and \g452012/U$2 ( \15962 , \8335 , RIdf2ee28_1910);
and \g452012/U$3 ( \15963 , RIfc776d8_6381, \8523 );
nor \g452012/U$1 ( \15964 , \15962 , \15963 );
and \g452011/U$2 ( \15965 , \8319 , RIdf30fe8_1934);
and \g452011/U$3 ( \15966 , RIdf33040_1957, \8326 );
nor \g452011/U$1 ( \15967 , \15965 , \15966 );
and \g445180/U$2 ( \15968 , \15961 , \15964 , \15967 );
nor \g445180/U$1 ( \15969 , \15968 , \8422 );
and \g446042/U$2 ( \15970 , RIfcd6160_7458, \8531 );
and \g446042/U$3 ( \15971 , RIe146208_2175, \8335 );
and \g448933/U$2 ( \15972 , RIe157008_2367, \8414 );
and \g448933/U$3 ( \15973 , \8409 , RIe15ca08_2431);
and \g448933/U$4 ( \15974 , RIe151608_2303, \8488 );
nor \g448933/U$1 ( \15975 , \15972 , \15973 , \15974 );
and \g454471/U$2 ( \15976 , \8313 , RIfc779a8_6383);
and \g454471/U$3 ( \15977 , RIe162408_2495, \8323 );
nor \g454471/U$1 ( \15978 , \15976 , \15977 );
not \g449947/U$3 ( \15979 , \15978 );
not \g449947/U$4 ( \15980 , \8328 );
and \g449947/U$2 ( \15981 , \15979 , \15980 );
and \g449947/U$5 ( \15982 , \8359 , RIfea7550_8220);
nor \g449947/U$1 ( \15983 , \15981 , \15982 );
and \g452020/U$2 ( \15984 , \8404 , RIe15f708_2463);
and \g452020/U$3 ( \15985 , RIe165108_2527, \8351 );
nor \g452020/U$1 ( \15986 , \15984 , \15985 );
and \g452021/U$2 ( \15987 , \8378 , RIe154308_2335);
and \g452021/U$3 ( \15988 , RIfe9dc08_8139, \8417 );
nor \g452021/U$1 ( \15989 , \15987 , \15988 );
nand \g447691/U$1 ( \15990 , \15975 , \15983 , \15986 , \15989 );
nor \g446042/U$1 ( \15991 , \15970 , \15971 , \15990 );
and \g452016/U$2 ( \15992 , \8356 , RIe14e908_2271);
and \g452016/U$3 ( \15993 , RIfcd1408_7403, \8340 );
nor \g452016/U$1 ( \15994 , \15992 , \15993 );
and \g452017/U$2 ( \15995 , \8319 , RIe148f08_2207);
and \g452017/U$3 ( \15996 , RIe14bc08_2239, \8326 );
nor \g452017/U$1 ( \15997 , \15995 , \15996 );
and \g445182/U$2 ( \15998 , \15991 , \15994 , \15997 );
nor \g445182/U$1 ( \15999 , \15998 , \8368 );
or \g444367/U$1 ( \16000 , \15879 , \15939 , \15969 , \15999 );
and \g446038/U$2 ( \16001 , RIdf22ab0_1771, \8531 );
and \g446038/U$3 ( \16002 , RIdf1aef0_1683, \8319 );
and \g448929/U$2 ( \16003 , RIdf26458_1812, \8414 );
and \g448929/U$3 ( \16004 , \8409 , RIfea8bd0_8236);
and \g448929/U$4 ( \16005 , RIee26cc8_4900, \8488 );
nor \g448929/U$1 ( \16006 , \16003 , \16004 , \16005 );
and \g454698/U$2 ( \16007 , \8313 , RIfc77de0_6386);
and \g454698/U$3 ( \16008 , RIfc93ba8_6703, \8323 );
nor \g454698/U$1 ( \16009 , \16007 , \16008 );
not \g449684/U$3 ( \16010 , \16009 );
not \g449684/U$4 ( \16011 , \8328 );
and \g449684/U$2 ( \16012 , \16010 , \16011 );
and \g449684/U$5 ( \16013 , \8359 , RIfcb1c98_7045);
nor \g449684/U$1 ( \16014 , \16012 , \16013 );
and \g452004/U$2 ( \16015 , \8404 , RIee27ad8_4910);
and \g452004/U$3 ( \16016 , RIee2ba20_4955, \8351 );
nor \g452004/U$1 ( \16017 , \16015 , \16016 );
and \g452005/U$2 ( \16018 , \8378 , RIfe9d7d0_8136);
and \g452005/U$3 ( \16019 , RIfe9d668_8135, \8417 );
nor \g452005/U$1 ( \16020 , \16018 , \16019 );
nand \g447686/U$1 ( \16021 , \16006 , \16014 , \16017 , \16020 );
nor \g446038/U$1 ( \16022 , \16001 , \16002 , \16021 );
and \g452002/U$2 ( \16023 , \8335 , RIfe9d938_8137);
and \g452002/U$3 ( \16024 , RIdf21598_1756, \8340 );
nor \g452002/U$1 ( \16025 , \16023 , \16024 );
and \g452001/U$2 ( \16026 , \8326 , RIdf1f6a8_1734);
and \g452001/U$3 ( \16027 , RIfcc0068_7207, \8356 );
nor \g452001/U$1 ( \16028 , \16026 , \16027 );
and \g445178/U$2 ( \16029 , \16022 , \16025 , \16028 );
nor \g445178/U$1 ( \16030 , \16029 , \8621 );
and \g446039/U$2 ( \16031 , RIdf2c560_1881, \8523 );
and \g446039/U$3 ( \16032 , RIde7c1d8_195, \8335 );
and \g448930/U$2 ( \16033 , RIe16df10_2628, \8414 );
and \g448930/U$3 ( \16034 , \8407 , RIde96290_322);
and \g448930/U$4 ( \16035 , RIdf37f00_2013, \8488 );
nor \g448930/U$1 ( \16036 , \16033 , \16034 , \16035 );
and \g454582/U$2 ( \16037 , \8313 , RIdecab08_770);
and \g454582/U$3 ( \16038 , RIdecd808_802, \8323 );
nor \g454582/U$1 ( \16039 , \16037 , \16038 );
not \g449945/U$3 ( \16040 , \16039 );
not \g449945/U$4 ( \16041 , \8328 );
and \g449945/U$2 ( \16042 , \16040 , \16041 );
and \g449945/U$5 ( \16043 , \8359 , RIe143508_2143);
nor \g449945/U$1 ( \16044 , \16042 , \16043 );
and \g453096/U$2 ( \16045 , \8404 , RIdec7e08_738);
and \g453096/U$3 ( \16046 , RIded0508_834, \8351 );
nor \g453096/U$1 ( \16047 , \16045 , \16046 );
and \g452010/U$2 ( \16048 , \8378 , RIe159d08_2399);
and \g452010/U$3 ( \16049 , RIdeb4308_514, \8417 );
nor \g452010/U$1 ( \16050 , \16048 , \16049 );
nand \g447688/U$1 ( \16051 , \16036 , \16044 , \16047 , \16050 );
nor \g446039/U$1 ( \16052 , \16031 , \16032 , \16051 );
and \g452569/U$2 ( \16053 , \8356 , RIdf1cde0_1705);
and \g452569/U$3 ( \16054 , RIdf004d8_1380, \8340 );
nor \g452569/U$1 ( \16055 , \16053 , \16054 );
and \g452008/U$2 ( \16056 , \8319 , RIdedbd40_965);
and \g452008/U$3 ( \16057 , RIdee6fd8_1092, \8326 );
nor \g452008/U$1 ( \16058 , \16056 , \16057 );
and \g445179/U$2 ( \16059 , \16052 , \16055 , \16058 );
nor \g445179/U$1 ( \16060 , \16059 , \8651 );
or \g444190/U$1 ( \16061 , \16000 , \16030 , \16060 );
_DC \g31cb/U$1 ( \16062 , \16061 , \8654 );
and \g450871/U$2 ( \16063 , \8319 , RIfcc8fd8_7309);
and \g450871/U$3 ( \16064 , RIe16a9a0_2590, \8324 );
nor \g450871/U$1 ( \16065 , \16063 , \16064 );
and \g445771/U$2 ( \16066 , RIfc75d88_6363, \8531 );
and \g445771/U$3 ( \16067 , RIe166e90_2548, \8335 );
and \g448593/U$2 ( \16068 , RIde88028_253, \8414 );
and \g448593/U$3 ( \16069 , \8407 , RIde8c1c8_273);
and \g448593/U$4 ( \16070 , RIfca4b10_6896, \8486 );
nor \g448593/U$1 ( \16071 , \16068 , \16069 , \16070 );
and \g454859/U$2 ( \16072 , \8313 , RIfcc8e70_7308);
and \g454859/U$3 ( \16073 , RIfc957c8_6723, \8323 );
nor \g454859/U$1 ( \16074 , \16072 , \16073 );
not \g449616/U$3 ( \16075 , \16074 );
not \g449616/U$4 ( \16076 , \8328 );
and \g449616/U$2 ( \16077 , \16075 , \16076 );
and \g449616/U$5 ( \16078 , \8359 , RIfcb0bb8_7033);
nor \g449616/U$1 ( \16079 , \16077 , \16078 );
and \g450885/U$2 ( \16080 , \8404 , RIfc5e610_6096);
and \g450885/U$3 ( \16081 , RIee1c840_4783, \8351 );
nor \g450885/U$1 ( \16082 , \16080 , \16081 );
and \g450892/U$2 ( \16083 , \8378 , RIde83b40_232);
and \g450892/U$3 ( \16084 , RIfe9e8b0_8148, \8417 );
nor \g450892/U$1 ( \16085 , \16083 , \16084 );
nand \g447495/U$1 ( \16086 , \16071 , \16079 , \16082 , \16085 );
nor \g445771/U$1 ( \16087 , \16066 , \16067 , \16086 );
and \g450866/U$2 ( \16088 , \8356 , RIfca4c78_6897);
and \g450866/U$3 ( \16089 , RIfc95390_6720, \8340 );
nor \g450866/U$1 ( \16090 , \16088 , \16089 );
nand \g445521/U$1 ( \16091 , \16065 , \16087 , \16090 );
and \g444743/U$2 ( \16092 , \16091 , \9700 );
and \g448576/U$2 ( \16093 , RIee1e190_4801, \8531 );
and \g448576/U$3 ( \16094 , \8488 , RIdeb0690_471);
and \g448576/U$4 ( \16095 , RIdec1490_663, \8383 );
nor \g448576/U$1 ( \16096 , \16093 , \16094 , \16095 );
and \g450826/U$2 ( \16097 , \8335 , RIde9a778_343);
and \g450826/U$3 ( \16098 , RIfcdf0d0_7560, \8340 );
nor \g450826/U$1 ( \16099 , \16097 , \16098 );
and \g454797/U$2 ( \16100 , \8313 , RIdea1078_375);
and \g454797/U$3 ( \16101 , RIdea7978_407, \8323 );
nor \g454797/U$1 ( \16102 , \16100 , \16101 );
not \g454796/U$1 ( \16103 , \16102 );
and \g449598/U$2 ( \16104 , \16103 , \8316 );
and \g449598/U$3 ( \16105 , RIdec4190_695, \8351 );
nor \g449598/U$1 ( \16106 , \16104 , \16105 );
and \g450820/U$2 ( \16107 , \8356 , RIdead990_439);
and \g450820/U$3 ( \16108 , RIfcebb50_7704, \8359 );
nor \g450820/U$1 ( \16109 , \16107 , \16108 );
nand \g448139/U$1 ( \16110 , \16096 , \16099 , \16106 , \16109 );
and \g444743/U$3 ( \16111 , \9702 , \16110 );
nor \g444743/U$1 ( \16112 , \16092 , \16111 );
and \g446550/U$2 ( \16113 , \11700 , RIdebba90_599);
and \g446550/U$3 ( \16114 , RIfc954f8_6721, \11702 );
nor \g446550/U$1 ( \16115 , \16113 , \16114 );
and \g446552/U$2 ( \16116 , \9724 , RIdebe790_631);
and \g446552/U$3 ( \16117 , RIfceaa70_7692, \9726 );
nor \g446552/U$1 ( \16118 , \16116 , \16117 );
and \g446551/U$2 ( \16119 , \9170 , RIdeb6090_535);
and \g446551/U$3 ( \16120 , RIdeb8d90_567, \9172 );
nor \g446551/U$1 ( \16121 , \16119 , \16120 );
nand \g444451/U$1 ( \16122 , \16112 , \16115 , \16118 , \16121 );
and \g450993/U$2 ( \16123 , \8326 , RIdf1eb68_1726);
and \g450993/U$3 ( \16124 , RIfc75518_6357, \8356 );
nor \g450993/U$1 ( \16125 , \16123 , \16124 );
and \g445798/U$2 ( \16126 , RIfe9eb80_8150, \8523 );
and \g445798/U$3 ( \16127 , RIfe9ece8_8151, \8319 );
and \g448629/U$2 ( \16128 , RIdf257b0_1803, \8414 );
and \g448629/U$3 ( \16129 , \8407 , RIdf273d0_1823);
and \g448629/U$4 ( \16130 , RIfceda40_7726, \8488 );
nor \g448629/U$1 ( \16131 , \16128 , \16129 , \16130 );
and \g455096/U$2 ( \16132 , \8313 , RIfc757e8_6359);
and \g455096/U$3 ( \16133 , RIfcd0328_7391, \8323 );
nor \g455096/U$1 ( \16134 , \16132 , \16133 );
not \g449652/U$3 ( \16135 , \16134 );
not \g449652/U$4 ( \16136 , \8328 );
and \g449652/U$2 ( \16137 , \16135 , \16136 );
and \g449652/U$5 ( \16138 , \8359 , RIfc95d68_6727);
nor \g449652/U$1 ( \16139 , \16137 , \16138 );
and \g451018/U$2 ( \16140 , \8404 , RIfcee6e8_7735);
and \g451018/U$3 ( \16141 , RIfc5e778_6097, \8351 );
nor \g451018/U$1 ( \16142 , \16140 , \16141 );
and \g451026/U$2 ( \16143 , \8378 , RIdf23b90_1783);
and \g451026/U$3 ( \16144 , RIdf296f8_1848, \8417 );
nor \g451026/U$1 ( \16145 , \16143 , \16144 );
nand \g447523/U$1 ( \16146 , \16131 , \16139 , \16142 , \16145 );
nor \g445798/U$1 ( \16147 , \16126 , \16127 , \16146 );
and \g450998/U$2 ( \16148 , \8335 , RIfe9ea18_8149);
and \g450998/U$3 ( \16149 , RIfcd01c0_7390, \8340 );
nor \g450998/U$1 ( \16150 , \16148 , \16149 );
nand \g445529/U$1 ( \16151 , \16125 , \16147 , \16150 );
and \g444840/U$2 ( \16152 , \16151 , \8752 );
and \g448612/U$2 ( \16153 , RIdec9b90_759, \8373 );
and \g448612/U$3 ( \16154 , \8383 , RIdecc890_791);
and \g448612/U$4 ( \16155 , RIdf36f88_2002, \8486 );
nor \g448612/U$1 ( \16156 , \16153 , \16154 , \16155 );
and \g454934/U$2 ( \16157 , \8313 , RIe16cf98_2617);
and \g454934/U$3 ( \16158 , RIde93e78_311, \8323 );
nor \g454934/U$1 ( \16159 , \16157 , \16158 );
not \g449634/U$3 ( \16160 , \16159 );
not \g449634/U$4 ( \16161 , \8376 );
and \g449634/U$2 ( \16162 , \16160 , \16161 );
and \g449634/U$5 ( \16163 , \8359 , RIe142590_2132);
nor \g449634/U$1 ( \16164 , \16162 , \16163 );
and \g450956/U$2 ( \16165 , \8404 , RIdec6e90_727);
and \g450956/U$3 ( \16166 , RIdecf590_823, \8351 );
nor \g450956/U$1 ( \16167 , \16165 , \16166 );
and \g450964/U$2 ( \16168 , \8378 , RIe158d90_2388);
and \g450964/U$3 ( \16169 , RIdeb3390_503, \8417 );
nor \g450964/U$1 ( \16170 , \16168 , \16169 );
nand \g447512/U$1 ( \16171 , \16156 , \16164 , \16167 , \16170 );
and \g444840/U$3 ( \16172 , \9010 , \16171 );
nor \g444840/U$1 ( \16173 , \16152 , \16172 );
and \g446583/U$2 ( \16174 , \11213 , RIdf1be68_1694);
and \g446583/U$3 ( \16175 , RIdf2b5e8_1870, \11215 );
nor \g446583/U$1 ( \16176 , \16174 , \16175 );
and \g446584/U$2 ( \16177 , \13239 , RIdee6060_1081);
and \g446584/U$3 ( \16178 , RIdeff560_1369, \13241 );
nor \g446584/U$1 ( \16179 , \16177 , \16178 );
and \g446585/U$2 ( \16180 , \13244 , RIde79dc0_184);
and \g446585/U$3 ( \16181 , RIdedadc8_954, \13246 );
nor \g446585/U$1 ( \16182 , \16180 , \16181 );
nand \g444559/U$1 ( \16183 , \16173 , \16176 , \16179 , \16182 );
and \g445728/U$2 ( \16184 , RIfe9e748_8147, \8373 );
and \g445728/U$3 ( \16185 , RIe153390_2324, \8378 );
and \g448536/U$2 ( \16186 , RIe147f90_2196, \8319 );
and \g448536/U$3 ( \16187 , \8326 , RIe14ac90_2228);
and \g448536/U$4 ( \16188 , RIe161490_2484, \8330 );
nor \g448536/U$1 ( \16189 , \16186 , \16187 , \16188 );
and \g450700/U$2 ( \16190 , \8335 , RIe145290_2164);
and \g450700/U$3 ( \16191 , RIfca6730_6916, \8340 );
nor \g450700/U$1 ( \16192 , \16190 , \16191 );
and \g454219/U$2 ( \16193 , \8313 , RIfce8b80_7670);
and \g454219/U$3 ( \16194 , RIe150690_2292, \8323 );
nor \g454219/U$1 ( \16195 , \16193 , \16194 );
not \g449558/U$3 ( \16196 , \16195 );
not \g449558/U$4 ( \16197 , \8347 );
and \g449558/U$2 ( \16198 , \16196 , \16197 );
and \g449558/U$5 ( \16199 , \8351 , RIe164190_2516);
nor \g449558/U$1 ( \16200 , \16198 , \16199 );
and \g450693/U$2 ( \16201 , \8356 , RIe14d990_2260);
and \g450693/U$3 ( \16202 , RIfc3ecc0_5740, \8359 );
nor \g450693/U$1 ( \16203 , \16201 , \16202 );
nand \g447473/U$1 ( \16204 , \16189 , \16192 , \16200 , \16203 );
nor \g445728/U$1 ( \16205 , \16184 , \16185 , \16204 );
and \g450677/U$2 ( \16206 , \8404 , RIe15e790_2452);
and \g450677/U$3 ( \16207 , RIe15ba90_2420, \8407 );
nor \g450677/U$1 ( \16208 , \16206 , \16207 );
and \g450669/U$2 ( \16209 , \8414 , RIe156090_2356);
and \g450669/U$3 ( \16210 , RIfc74f78_6353, \8417 );
nor \g450669/U$1 ( \16211 , \16209 , \16210 );
and \g444947/U$2 ( \16212 , \16205 , \16208 , \16211 );
nor \g444947/U$1 ( \16213 , \16212 , \8368 );
and \g445740/U$2 ( \16214 , RIe140268_2107, \8417 );
and \g445740/U$3 ( \16215 , RIfc74b40_6350, \8404 );
and \g448554/U$2 ( \16216 , RIdf301d8_1924, \8317 );
and \g448554/U$3 ( \16217 , \8326 , RIdf327d0_1951);
and \g448554/U$4 ( \16218 , RIfc5f2b8_6105, \8330 );
nor \g448554/U$1 ( \16219 , \16216 , \16217 , \16218 );
and \g450759/U$2 ( \16220 , \8335 , RIdf2e2e8_1902);
and \g450759/U$3 ( \16221 , RIdf34828_1974, \8340 );
nor \g450759/U$1 ( \16222 , \16220 , \16221 );
and \g454244/U$2 ( \16223 , \8313 , RIfc965d8_6733);
and \g454244/U$3 ( \16224 , RIfcc1850_7224, \8323 );
nor \g454244/U$1 ( \16225 , \16223 , \16224 );
not \g449575/U$3 ( \16226 , \16225 );
not \g449575/U$4 ( \16227 , \8347 );
and \g449575/U$2 ( \16228 , \16226 , \16227 );
and \g449575/U$5 ( \16229 , \8351 , RIfcee2b0_7732);
nor \g449575/U$1 ( \16230 , \16228 , \16229 );
and \g450751/U$2 ( \16231 , \8356 , RIfc96038_6729);
and \g450751/U$3 ( \16232 , RIfcc1c88_7227, \8359 );
nor \g450751/U$1 ( \16233 , \16231 , \16232 );
nand \g447484/U$1 ( \16234 , \16219 , \16222 , \16230 , \16233 );
nor \g445740/U$1 ( \16235 , \16214 , \16215 , \16234 );
and \g450733/U$2 ( \16236 , \8378 , RIdf39c88_2034);
and \g450733/U$3 ( \16237 , RIfc753b0_6356, \8371 );
nor \g450733/U$1 ( \16238 , \16236 , \16237 );
and \g450732/U$2 ( \16239 , \8412 , RIdf3be48_2058);
and \g450732/U$3 ( \16240 , RIdf3e170_2083, \8409 );
nor \g450732/U$1 ( \16241 , \16239 , \16240 );
and \g444965/U$2 ( \16242 , \16235 , \16238 , \16241 );
nor \g444965/U$1 ( \16243 , \16242 , \8422 );
or \g444357/U$1 ( \16244 , \16122 , \16183 , \16213 , \16243 );
and \g445701/U$2 ( \16245 , RIdef4160_1241, \8356 );
and \g445701/U$3 ( \16246 , RIdefc860_1337, \8359 );
and \g448501/U$2 ( \16247 , RIdeee760_1177, \8326 );
and \g448501/U$3 ( \16248 , \8371 , RIdf10360_1561);
and \g448501/U$4 ( \16249 , RIdf13060_1593, \8383 );
nor \g448501/U$1 ( \16250 , \16247 , \16248 , \16249 );
and \g454557/U$2 ( \16251 , \8313 , RIdf04f60_1433);
and \g454557/U$3 ( \16252 , RIdf07c60_1465, \8323 );
nor \g454557/U$1 ( \16253 , \16251 , \16252 );
not \g449520/U$3 ( \16254 , \16253 );
not \g449520/U$4 ( \16255 , \8376 );
and \g449520/U$2 ( \16256 , \16254 , \16255 );
and \g449520/U$5 ( \16257 , \8340 , RIdef1460_1209);
nor \g449520/U$1 ( \16258 , \16256 , \16257 );
and \g450558/U$2 ( \16259 , \8404 , RIdf0d660_1529);
and \g450558/U$3 ( \16260 , RIdf15d60_1625, \8351 );
nor \g450558/U$1 ( \16261 , \16259 , \16260 );
and \g450565/U$2 ( \16262 , \8378 , RIdf02260_1401);
and \g450565/U$3 ( \16263 , RIdf0a960_1497, \8417 );
nor \g450565/U$1 ( \16264 , \16262 , \16263 );
nand \g447454/U$1 ( \16265 , \16250 , \16258 , \16261 , \16264 );
nor \g445701/U$1 ( \16266 , \16245 , \16246 , \16265 );
and \g450545/U$2 ( \16267 , \8335 , RIdee8d60_1113);
and \g450545/U$3 ( \16268 , RIdef9b60_1305, \8488 );
nor \g450545/U$1 ( \16269 , \16267 , \16268 );
and \g454123/U$2 ( \16270 , \8319 , RIdeeba60_1145);
and \g454123/U$3 ( \16271 , RIdef6e60_1273, \8531 );
nor \g454123/U$1 ( \16272 , \16270 , \16271 );
and \g445500/U$2 ( \16273 , \16266 , \16269 , \16272 );
nor \g445500/U$1 ( \16274 , \16273 , \8477 );
and \g445714/U$2 ( \16275 , RIfc5ee80_6102, \8371 );
and \g445714/U$3 ( \16276 , RIdee00c0_1013, \8414 );
and \g448518/U$2 ( \16277 , RIded4450_879, \8317 );
and \g448518/U$3 ( \16278 , \8326 , RIded6610_903);
and \g448518/U$4 ( \16279 , RIfc96308_6731, \8383 );
nor \g448518/U$1 ( \16280 , \16277 , \16278 , \16279 );
and \g450625/U$2 ( \16281 , \8335 , RIded2290_855);
and \g450625/U$3 ( \16282 , RIded8938_928, \8340 );
nor \g450625/U$1 ( \16283 , \16281 , \16282 );
and \g454422/U$2 ( \16284 , \8313 , RIfc74ca8_6351);
and \g454422/U$3 ( \16285 , RIfc75248_6355, \8323 );
nor \g454422/U$1 ( \16286 , \16284 , \16285 );
not \g449536/U$3 ( \16287 , \16286 );
not \g449536/U$4 ( \16288 , \8347 );
and \g449536/U$2 ( \16289 , \16287 , \16288 );
and \g449536/U$5 ( \16290 , \8351 , RIfc961a0_6730);
nor \g449536/U$1 ( \16291 , \16289 , \16290 );
and \g450622/U$2 ( \16292 , \8356 , RIfcb0618_7029);
and \g450622/U$3 ( \16293 , RIfc96470_6732, \8359 );
nor \g450622/U$1 ( \16294 , \16292 , \16293 );
nand \g447467/U$1 ( \16295 , \16280 , \16283 , \16291 , \16294 );
nor \g445714/U$1 ( \16296 , \16275 , \16276 , \16295 );
and \g450599/U$2 ( \16297 , \8404 , RIfce6150_7640);
and \g450599/U$3 ( \16298 , RIdee42d8_1060, \8417 );
nor \g450599/U$1 ( \16299 , \16297 , \16298 );
and \g450604/U$2 ( \16300 , \8378 , RIdeddac8_986);
and \g450604/U$3 ( \16301 , RIdee1e48_1034, \8409 );
nor \g450604/U$1 ( \16302 , \16300 , \16301 );
and \g444937/U$2 ( \16303 , \16296 , \16299 , \16302 );
nor \g444937/U$1 ( \16304 , \16303 , \8481 );
or \g444202/U$1 ( \16305 , \16244 , \16274 , \16304 );
_DC \g3250/U$1 ( \16306 , \16305 , \8654 );
not \g455683/U$2 ( \16307 , RIbc62550_11);
nand \g455683/U$1 ( \16308 , \16307 , RIbc625c8_12);
not \g455724/U$1 ( \16309 , RIbc62460_9);
not \g455726/U$1 ( \16310 , RIbc624d8_10);
or \g455703/U$1 ( \16311 , \16309 , \16310 );
nor \g455604/U$1 ( \16312 , \16308 , \16311 );
buf \g455594/U$1 ( \16313 , \16312 );
and \g452532/U$2 ( \16314 , \16313 , RIfcb6180_7094);
not \g455718/U$2 ( \16315 , RIbc62550_11);
nor \g455718/U$1 ( \16316 , \16315 , RIbc625c8_12);
buf \g455717/U$1 ( \16317 , \16316 );
not \g455701/U$1 ( \16318 , \16311 );
and \g455593/U$1 ( \16319 , \16317 , \16318 );
not \drc_bufs455844/U$1 ( \16320 , \16319 );
not \drc_bufs455843/U$1 ( \16321 , \16320 );
and \g452532/U$3 ( \16322 , RIe224940_4706, \16321 );
nor \g452532/U$1 ( \16323 , \16314 , \16322 );
and \g455706/U$1 ( \16324 , RIbc625c8_12, RIbc62550_11);
buf \g455704/U$1 ( \16325 , \16324 );
and \g455537/U$1 ( \16326 , \16325 , \16318 );
not \drc_bufs455870/U$1 ( \16327 , \16326 );
not \drc_bufs455868/U$1 ( \16328 , \16327 );
and \g446159/U$2 ( \16329 , RIfc44cd8_5805, \16328 );
or \g455711/U$1 ( \16330 , \16309 , RIbc624d8_10);
nor \g455689/U$1 ( \16331 , RIbc625c8_12, RIbc62550_11);
not \g455688/U$1 ( \16332 , \16331 );
nor \g455519/U$1 ( \16333 , \16330 , \16332 );
buf \g455510/U$1 ( \16334 , \16333 );
and \g446159/U$3 ( \16335 , RIe216840_4546, \16334 );
and \g455699/U$1 ( \16336 , \16310 , \16309 );
and \g455576/U$1 ( \16337 , \16317 , \16336 );
and \g449083/U$2 ( \16338 , RIe20e140_4450, \16337 );
and \g455572/U$1 ( \16339 , \16325 , \16336 );
not \drc_bufs455766/U$1 ( \16340 , \16339 );
not \drc_bufs455764/U$1 ( \16341 , \16340 );
and \g449083/U$3 ( \16342 , \16341 , RIfcab1b8_6969);
not \g455709/U$1 ( \16343 , \16330 );
and \g455648/U$1 ( \16344 , \16317 , \16343 );
and \g449083/U$4 ( \16345 , RIe21ef40_4642, \16344 );
nor \g449083/U$1 ( \16346 , \16338 , \16342 , \16345 );
and \g454186/U$2 ( \16347 , \16317 , RIe213b40_4514);
and \g454186/U$3 ( \16348 , RIfc4dc48_5907, \16325 );
nor \g454186/U$1 ( \16349 , \16347 , \16348 );
not \g450097/U$3 ( \16350 , \16349 );
or \g455708/U$1 ( \16351 , \16310 , RIbc62460_9);
not \g450097/U$4 ( \16352 , \16351 );
and \g450097/U$2 ( \16353 , \16350 , \16352 );
and \g455615/U$1 ( \16354 , \16343 , \16325 );
not \drc_bufs455805/U$1 ( \16355 , \16354 );
not \drc_bufs455804/U$1 ( \16356 , \16355 );
and \g450097/U$5 ( \16357 , \16356 , RIfc55ad8_5997);
nor \g450097/U$1 ( \16358 , \16353 , \16357 );
not \g455698/U$1 ( \16359 , \16336 );
nor \g455498/U$1 ( \16360 , \16359 , \16332 );
buf \g455497/U$1 ( \16361 , \16360 );
and \g452536/U$2 ( \16362 , \16361 , RIe208740_4386);
nor \g455586/U$1 ( \16363 , \16359 , \16308 );
buf \g455585/U$1 ( \16364 , \16363 );
and \g452536/U$3 ( \16365 , RIe20b440_4418, \16364 );
nor \g452536/U$1 ( \16366 , \16362 , \16365 );
nor \g455509/U$1 ( \16367 , \16351 , \16332 );
buf \g455508/U$1 ( \16368 , \16367 );
and \g452535/U$2 ( \16369 , \16368 , RIe210e40_4482);
nor \g455626/U$1 ( \16370 , \16351 , \16308 );
buf \g455625/U$1 ( \16371 , \16370 );
and \g452535/U$3 ( \16372 , RIfcdcf10_7536, \16371 );
nor \g452535/U$1 ( \16373 , \16369 , \16372 );
nand \g447770/U$1 ( \16374 , \16346 , \16358 , \16366 , \16373 );
nor \g446159/U$1 ( \16375 , \16329 , \16335 , \16374 );
nor \g455530/U$1 ( \16376 , \16332 , \16311 );
buf \g455520/U$1 ( \16377 , \16376 );
and \g452533/U$2 ( \16378 , \16377 , RIe221c40_4674);
nor \g455679/U$1 ( \16379 , \16330 , \16308 );
buf \g455678/U$1 ( \16380 , \16379 );
and \g452533/U$3 ( \16381 , RIe219540_4578, \16380 );
nor \g452533/U$1 ( \16382 , \16378 , \16381 );
nand \g445614/U$1 ( \16383 , \16323 , \16375 , \16382 );
or \g455680/U$1 ( \16384 , RIbc62208_4, RIbc62190_3, RIbc62280_5, RIbc62118_2);
not \g454132/U$2 ( \16385 , \16384 );
nand \g454132/U$1 ( \16386 , \16385 , RIbc622f8_6);
not \g450540/U$2 ( \16387 , \16386 );
nand \g450540/U$1 ( \16388 , \16387 , RIbc623e8_8);
or \g448480/U$1 ( \16389 , \16388 , RIbc62370_7);
not \g448479/U$1 ( \16390 , \16389 );
and \g444859/U$2 ( \16391 , \16383 , \16390 );
or \g450541/U$1 ( \16392 , \16386 , RIbc623e8_8);
or \g448458/U$1 ( \16393 , \16392 , RIbc62370_7);
not \g448457/U$1 ( \16394 , \16393 );
and \g449081/U$2 ( \16395 , RIf164828_5603, \16344 );
and \g449081/U$3 ( \16396 , \16354 , RIfcd2ec0_7422);
not \drc_bufs455753/U$1 ( \16397 , \16337 );
not \drc_bufs455751/U$1 ( \16398 , \16397 );
and \g449081/U$4 ( \16399 , RIfc4f160_5922, \16398 );
nor \g449081/U$1 ( \16400 , \16395 , \16396 , \16399 );
and \g454893/U$2 ( \16401 , \16317 , RIfc64178_6161);
and \g454893/U$3 ( \16402 , RIfce3720_7610, \16325 );
nor \g454893/U$1 ( \16403 , \16401 , \16402 );
not \g450095/U$3 ( \16404 , \16403 );
not \g450095/U$4 ( \16405 , \16311 );
and \g450095/U$2 ( \16406 , \16404 , \16405 );
and \g450095/U$5 ( \16407 , \16341 , RIfc59318_6037);
nor \g450095/U$1 ( \16408 , \16406 , \16407 );
and \g452525/U$2 ( \16409 , \16377 , RIe201558_4305);
and \g452525/U$3 ( \16410 , RIe203178_4325, \16313 );
nor \g452525/U$1 ( \16411 , \16409 , \16410 );
and \g452527/U$2 ( \16412 , \16334 , RIf162398_5577);
and \g452527/U$3 ( \16413 , RIfc7f838_6473, \16380 );
nor \g452527/U$1 ( \16414 , \16412 , \16413 );
nand \g447358/U$1 ( \16415 , \16400 , \16408 , \16411 , \16414 );
and \g444859/U$3 ( \16416 , \16394 , \16415 );
nor \g444859/U$1 ( \16417 , \16391 , \16416 );
not \g455491/U$1 ( \16418 , \16360 );
nor \g448413/U$1 ( \16419 , \16393 , \16418 );
and \g446934/U$2 ( \16420 , \16419 , RIfcebf88_7707);
not \g455579/U$1 ( \16421 , \16363 );
nor \g448421/U$1 ( \16422 , \16393 , \16421 );
and \g446934/U$3 ( \16423 , RIf15ac10_5492, \16422 );
nor \g446934/U$1 ( \16424 , \16420 , \16423 );
not \g455924/U$2 ( \16425 , \16317 );
nor \g455924/U$1 ( \16426 , \16425 , \16351 );
buf \g455635/U$1 ( \16427 , \16426 );
not \g455629/U$1 ( \16428 , \16427 );
nor \g448429/U$1 ( \16429 , \16393 , \16428 );
and \g446932/U$2 ( \16430 , \16429 , RIfca8bc0_6942);
not \g455923/U$2 ( \16431 , \16325 );
nor \g455923/U$1 ( \16432 , \16431 , \16351 );
not \drc_bufs455831/U$1 ( \16433 , \16432 );
nor \g448428/U$1 ( \16434 , \16393 , \16433 );
and \g446932/U$3 ( \16435 , RIfcc9c80_7318, \16434 );
nor \g446932/U$1 ( \16436 , \16430 , \16435 );
not \g455500/U$1 ( \16437 , \16367 );
nor \g448414/U$1 ( \16438 , \16393 , \16437 );
and \g446933/U$2 ( \16439 , \16438 , RIfea2c30_8196);
not \g455617/U$1 ( \16440 , \16370 );
nor \g448430/U$1 ( \16441 , \16393 , \16440 );
and \g446933/U$3 ( \16442 , RIfea2ac8_8195, \16441 );
nor \g446933/U$1 ( \16443 , \16439 , \16442 );
nand \g444621/U$1 ( \16444 , \16417 , \16424 , \16436 , \16443 );
and \g452518/U$2 ( \16445 , \16371 , RIe1b31c8_3415);
and \g452518/U$3 ( \16446 , RIfc50d80_5942, \16427 );
nor \g452518/U$1 ( \16447 , \16445 , \16446 );
not \drc_bufs455829/U$1 ( \16448 , \16433 );
and \g446155/U$2 ( \16449 , RIfc9bfd8_6797, \16448 );
and \g446155/U$3 ( \16450 , RIe1ab8d8_3329, \16361 );
and \g449080/U$2 ( \16451 , RIfc6bd38_6249, \16321 );
and \g449080/U$3 ( \16452 , \16328 , RIfc63908_6155);
and \g449080/U$4 ( \16453 , RIfc9d658_6813, \16337 );
nor \g449080/U$1 ( \16454 , \16451 , \16452 , \16453 );
and \g454891/U$2 ( \16455 , \16317 , RIfc92ac8_6691);
and \g454891/U$3 ( \16456 , RIfc66fe0_6194, \16325 );
nor \g454891/U$1 ( \16457 , \16455 , \16456 );
not \g450094/U$3 ( \16458 , \16457 );
not \g450094/U$4 ( \16459 , \16330 );
and \g450094/U$2 ( \16460 , \16458 , \16459 );
and \g450094/U$5 ( \16461 , \16341 , RIfc4df18_5909);
nor \g450094/U$1 ( \16462 , \16460 , \16461 );
and \g452520/U$2 ( \16463 , \16377 , RIe1b7f20_3470);
and \g452520/U$3 ( \16464 , RIe1ba0e0_3494, \16313 );
nor \g452520/U$1 ( \16465 , \16463 , \16464 );
and \g452521/U$2 ( \16466 , \16334 , RIfea2f00_8198);
and \g452521/U$3 ( \16467 , RIe1b5d60_3446, \16380 );
nor \g452521/U$1 ( \16468 , \16466 , \16467 );
nand \g447357/U$1 ( \16469 , \16454 , \16462 , \16465 , \16468 );
nor \g446155/U$1 ( \16470 , \16449 , \16450 , \16469 );
and \g452519/U$2 ( \16471 , \16364 , RIe1ad0c0_3346);
and \g452519/U$3 ( \16472 , RIe1b1878_3397, \16368 );
nor \g452519/U$1 ( \16473 , \16471 , \16472 );
nand \g445613/U$1 ( \16474 , \16447 , \16470 , \16473 );
nor \g454134/U$1 ( \16475 , \16384 , RIbc622f8_6);
nand \g450544/U$1 ( \16476 , RIbc623e8_8, \16475 );
nor \g448462/U$1 ( \16477 , \16476 , RIbc62370_7);
and \g444917/U$2 ( \16478 , \16474 , \16477 );
not \g455727/U$1 ( \16479 , RIbc62370_7);
or \g448472/U$1 ( \16480 , \16476 , \16479 );
not \g448471/U$1 ( \16481 , \16480 );
and \g449076/U$2 ( \16482 , RIfc434f0_5788, \16398 );
and \g449076/U$3 ( \16483 , \16341 , RIfc64010_6160);
not \drc_bufs455792/U$1 ( \16484 , \16344 );
not \drc_bufs455790/U$1 ( \16485 , \16484 );
and \g449076/U$4 ( \16486 , RIf155a80_5434, \16485 );
nor \g449076/U$1 ( \16487 , \16482 , \16483 , \16486 );
and \g454206/U$2 ( \16488 , \16317 , RIfcccae8_7351);
and \g454206/U$3 ( \16489 , RIfccdbc8_7363, \16325 );
nor \g454206/U$1 ( \16490 , \16488 , \16489 );
not \g450091/U$3 ( \16491 , \16490 );
not \g450091/U$4 ( \16492 , \16351 );
and \g450091/U$2 ( \16493 , \16491 , \16492 );
and \g450091/U$5 ( \16494 , \16356 , RIf1565c0_5442);
nor \g450091/U$1 ( \16495 , \16493 , \16494 );
and \g452515/U$2 ( \16496 , \16361 , RIe1eee08_4095);
and \g452515/U$3 ( \16497 , RIfc4c028_5887, \16364 );
nor \g452515/U$1 ( \16498 , \16496 , \16497 );
and \g452513/U$2 ( \16499 , \16368 , RIfec6018_8373);
and \g452513/U$3 ( \16500 , RIfca6cd0_6920, \16371 );
nor \g452513/U$1 ( \16501 , \16499 , \16500 );
nand \g447768/U$1 ( \16502 , \16487 , \16495 , \16498 , \16501 );
and \g444917/U$3 ( \16503 , \16481 , \16502 );
nor \g444917/U$1 ( \16504 , \16478 , \16503 );
nor \g448444/U$1 ( \16505 , \16480 , \16320 );
and \g446928/U$2 ( \16506 , \16505 , RIfca1870_6860);
nor \g448422/U$1 ( \16507 , \16480 , \16327 );
and \g446928/U$3 ( \16508 , RIfcbb040_7150, \16507 );
nor \g446928/U$1 ( \16509 , \16506 , \16508 );
not \g455513/U$1 ( \16510 , \16334 );
nor \g448450/U$1 ( \16511 , \16480 , \16510 );
and \g446931/U$2 ( \16512 , \16511 , RIe1f6428_4179);
not \g455677/U$1 ( \16513 , \16380 );
nor \g448449/U$1 ( \16514 , \16480 , \16513 );
and \g446931/U$3 ( \16515 , RIfc45c50_5816, \16514 );
nor \g446931/U$1 ( \16516 , \16512 , \16515 );
not \g455522/U$1 ( \16517 , \16376 );
nor \g448448/U$1 ( \16518 , \16480 , \16517 );
and \g446929/U$2 ( \16519 , \16518 , RIe1faeb0_4232);
not \g455596/U$1 ( \16520 , \16312 );
nor \g448445/U$1 ( \16521 , \16480 , \16520 );
and \g446929/U$3 ( \16522 , RIfc93d10_6704, \16521 );
nor \g446929/U$1 ( \16523 , \16519 , \16522 );
nand \g444620/U$1 ( \16524 , \16504 , \16509 , \16516 , \16523 );
and \g446152/U$2 ( \16525 , RIe1e12a8_3939, \16354 );
and \g446152/U$3 ( \16526 , RIe1caaa8_3683, \16368 );
and \g449071/U$2 ( \16527 , RIe1e99a8_4035, \16321 );
and \g449071/U$3 ( \16528 , \16328 , RIe1ec6a8_4067);
and \g449071/U$4 ( \16529 , RIe1d04a8_3747, \16427 );
nor \g449071/U$1 ( \16530 , \16527 , \16528 , \16529 );
and \g452504/U$2 ( \16531 , \16361 , RIe1bf6a8_3555);
and \g452504/U$3 ( \16532 , RIe1c23a8_3587, \16364 );
nor \g452504/U$1 ( \16533 , \16531 , \16532 );
and \g452502/U$2 ( \16534 , \16377 , RIe1e3fa8_3971);
and \g452502/U$3 ( \16535 , RIe1e6ca8_4003, \16313 );
nor \g452502/U$1 ( \16536 , \16534 , \16535 );
and \g454878/U$2 ( \16537 , \16317 , RIe1c50a8_3619);
and \g454878/U$3 ( \16538 , RIe1c7da8_3651, \16325 );
nor \g454878/U$1 ( \16539 , \16537 , \16538 );
not \g454877/U$1 ( \16540 , \16539 );
and \g450087/U$2 ( \16541 , \16540 , \16336 );
and \g450087/U$3 ( \16542 , RIe1d31a8_3779, \16432 );
nor \g450087/U$1 ( \16543 , \16541 , \16542 );
nand \g448074/U$1 ( \16544 , \16530 , \16533 , \16536 , \16543 );
nor \g446152/U$1 ( \16545 , \16525 , \16526 , \16544 );
and \g452500/U$2 ( \16546 , \16334 , RIe1d8ba8_3843);
and \g452500/U$3 ( \16547 , RIe1cd7a8_3715, \16371 );
nor \g452500/U$1 ( \16548 , \16546 , \16547 );
and \g452499/U$2 ( \16549 , \16380 , RIe1db8a8_3875);
and \g452499/U$3 ( \16550 , RIe1de5a8_3907, \16485 );
nor \g452499/U$1 ( \16551 , \16549 , \16550 );
and \g445258/U$2 ( \16552 , \16545 , \16548 , \16551 );
not \g450539/U$2 ( \16553 , RIbc623e8_8);
nand \g450539/U$1 ( \16554 , \16553 , \16475 );
or \g448478/U$1 ( \16555 , \16554 , \16479 );
nor \g445258/U$1 ( \16556 , \16552 , \16555 );
and \g446153/U$2 ( \16557 , RIe1ffaa0_4286, \16427 );
and \g446153/U$3 ( \16558 , RIe1f19a0_4126, \16368 );
and \g449074/U$2 ( \16559 , RIe179ce8_2763, \16485 );
and \g449074/U$3 ( \16560 , \16354 , RIe18d7e8_2987);
and \g449074/U$4 ( \16561 , RIe1bc9a8_3523, \16398 );
nor \g449074/U$1 ( \16562 , \16559 , \16560 , \16561 );
and \g454881/U$2 ( \16563 , \16317 , RIe1a6ce8_3275);
and \g454881/U$3 ( \16564 , RIe1a99e8_3307, \16325 );
nor \g454881/U$1 ( \16565 , \16563 , \16564 );
not \g450090/U$3 ( \16566 , \16565 );
not \g450090/U$4 ( \16567 , \16311 );
and \g450090/U$2 ( \16568 , \16566 , \16567 );
and \g450090/U$5 ( \16569 , \16341 , RIe1d5ea8_3811);
nor \g450090/U$1 ( \16570 , \16568 , \16569 );
and \g452508/U$2 ( \16571 , \16377 , RIe1a12e8_3211);
and \g452508/U$3 ( \16572 , RIe1a3fe8_3243, \16313 );
nor \g452508/U$1 ( \16573 , \16571 , \16572 );
and \g452509/U$2 ( \16574 , \16334 , RIe21c240_4610);
and \g452509/U$3 ( \16575 , RIe227640_4738, \16380 );
nor \g452509/U$1 ( \16576 , \16574 , \16575 );
nand \g447356/U$1 ( \16577 , \16562 , \16570 , \16573 , \16576 );
nor \g446153/U$1 ( \16578 , \16557 , \16558 , \16577 );
and \g452507/U$2 ( \16579 , \16361 , RIe171e58_2673);
and \g452507/U$3 ( \16580 , RIe205a40_4354, \16432 );
nor \g452507/U$1 ( \16581 , \16579 , \16580 );
and \g452506/U$2 ( \16582 , \16364 , RIe1af820_3374);
and \g452506/U$3 ( \16583 , RIe1f8e58_4209, \16371 );
nor \g452506/U$1 ( \16584 , \16582 , \16583 );
and \g445260/U$2 ( \16585 , \16578 , \16581 , \16584 );
or \g448486/U$1 ( \16586 , \16554 , RIbc62370_7);
nor \g445260/U$1 ( \16587 , \16585 , \16586 );
or \g444355/U$1 ( \16588 , \16444 , \16524 , \16556 , \16587 );
and \g446149/U$2 ( \16589 , RIe19e5e8_3179, \16326 );
and \g446149/U$3 ( \16590 , RIe1904e8_3019, \16334 );
and \g449068/U$2 ( \16591 , RIe1823e8_2859, \16337 );
and \g449068/U$3 ( \16592 , \16341 , RIfc8e310_6640);
and \g449068/U$4 ( \16593 , RIe195ee8_3083, \16485 );
nor \g449068/U$1 ( \16594 , \16591 , \16592 , \16593 );
and \g454225/U$2 ( \16595 , \16317 , RIe187de8_2923);
and \g454225/U$3 ( \16596 , RIe18aae8_2955, \16325 );
nor \g454225/U$1 ( \16597 , \16595 , \16596 );
not \g450082/U$3 ( \16598 , \16597 );
not \g450082/U$4 ( \16599 , \16351 );
and \g450082/U$2 ( \16600 , \16598 , \16599 );
and \g450082/U$5 ( \16601 , \16356 , RIfc846f8_6529);
nor \g450082/U$1 ( \16602 , \16600 , \16601 );
and \g452487/U$2 ( \16603 , \16361 , RIe17c9e8_2795);
and \g452487/U$3 ( \16604 , RIe17f6e8_2827, \16364 );
nor \g452487/U$1 ( \16605 , \16603 , \16604 );
and \g452486/U$2 ( \16606 , \16368 , RIe1850e8_2891);
and \g452486/U$3 ( \16607 , RIfce2be0_7602, \16371 );
nor \g452486/U$1 ( \16608 , \16606 , \16607 );
nand \g447764/U$1 ( \16609 , \16594 , \16602 , \16605 , \16608 );
nor \g446149/U$1 ( \16610 , \16589 , \16590 , \16609 );
and \g452483/U$2 ( \16611 , \16377 , RIe198be8_3115);
and \g452483/U$3 ( \16612 , RIe1931e8_3051, \16380 );
nor \g452483/U$1 ( \16613 , \16611 , \16612 );
and \g452482/U$2 ( \16614 , \16313 , RIfca84b8_6937);
and \g452482/U$3 ( \16615 , RIe19b8e8_3147, \16319 );
nor \g452482/U$1 ( \16616 , \16614 , \16615 );
and \g445255/U$2 ( \16617 , \16610 , \16613 , \16616 );
or \g448484/U$1 ( \16618 , \16388 , \16479 );
nor \g445255/U$1 ( \16619 , \16617 , \16618 );
and \g446150/U$2 ( \16620 , RIfc642e0_6162, \16448 );
and \g446150/U$3 ( \16621 , RIfccaec8_7331, \16361 );
and \g449070/U$2 ( \16622 , RIfccc278_7345, \16321 );
and \g449070/U$3 ( \16623 , \16326 , RIfcd1570_7404);
and \g449070/U$4 ( \16624 , RIfc5c720_6074, \16398 );
nor \g449070/U$1 ( \16625 , \16622 , \16623 , \16624 );
and \g454875/U$2 ( \16626 , \16317 , RIfc60398_6117);
and \g454875/U$3 ( \16627 , RIfcc1b20_7226, \16325 );
nor \g454875/U$1 ( \16628 , \16626 , \16627 );
not \g450085/U$3 ( \16629 , \16628 );
not \g450085/U$4 ( \16630 , \16330 );
and \g450085/U$2 ( \16631 , \16629 , \16630 );
and \g450085/U$5 ( \16632 , \16341 , RIfca9598_6949);
nor \g450085/U$1 ( \16633 , \16631 , \16632 );
and \g452493/U$2 ( \16634 , \16377 , RIfea2d98_8197);
and \g452493/U$3 ( \16635 , RIf1404c8_5191, \16313 );
nor \g452493/U$1 ( \16636 , \16634 , \16635 );
and \g452494/U$2 ( \16637 , \16334 , RIee3da68_5160);
and \g452494/U$3 ( \16638 , RIee3e5a8_5168, \16380 );
nor \g452494/U$1 ( \16639 , \16637 , \16638 );
nand \g447354/U$1 ( \16640 , \16625 , \16633 , \16636 , \16639 );
nor \g446150/U$1 ( \16641 , \16620 , \16621 , \16640 );
and \g452492/U$2 ( \16642 , \16364 , RIfc6bea0_6250);
and \g452492/U$3 ( \16643 , RIfec6180_8374, \16368 );
nor \g452492/U$1 ( \16644 , \16642 , \16643 );
and \g452491/U$2 ( \16645 , \16371 , RIee3a228_5120);
and \g452491/U$3 ( \16646 , RIfca7f18_6933, \16427 );
nor \g452491/U$1 ( \16647 , \16645 , \16646 );
and \g445256/U$2 ( \16648 , \16641 , \16644 , \16647 );
or \g448460/U$1 ( \16649 , \16392 , \16479 );
nor \g445256/U$1 ( \16650 , \16648 , \16649 );
or \g444276/U$1 ( \16651 , \16588 , \16619 , \16650 );
buf \g455926/U$1 ( \16652 , \16384 );
_DC \g3362/U$1 ( \16653 , \16651 , \16652 );
and \g452643/U$2 ( \16654 , \16361 , RIe2085d8_4385);
and \g452643/U$3 ( \16655 , RIe2139d8_4513, \16427 );
nor \g452643/U$1 ( \16656 , \16654 , \16655 );
and \g446182/U$2 ( \16657 , RIfc40070_5754, \16432 );
and \g446182/U$3 ( \16658 , RIf169850_5660, \16371 );
and \g449114/U$2 ( \16659 , RIe2247d8_4705, \16321 );
and \g449114/U$3 ( \16660 , \16328 , RIfc40bb0_5762);
and \g449114/U$4 ( \16661 , RIe20dfd8_4449, \16337 );
nor \g449114/U$1 ( \16662 , \16659 , \16660 , \16661 );
and \g454952/U$2 ( \16663 , \16317 , RIe21edd8_4641);
and \g454952/U$3 ( \16664 , RIfcd7d80_7478, \16325 );
nor \g454952/U$1 ( \16665 , \16663 , \16664 );
not \g450129/U$3 ( \16666 , \16665 );
not \g450129/U$4 ( \16667 , \16330 );
and \g450129/U$2 ( \16668 , \16666 , \16667 );
and \g450129/U$5 ( \16669 , \16341 , RIfcc1580_7222);
nor \g450129/U$1 ( \16670 , \16668 , \16669 );
and \g452645/U$2 ( \16671 , \16377 , RIe221ad8_4673);
and \g452645/U$3 ( \16672 , RIfc77138_6377, \16313 );
nor \g452645/U$1 ( \16673 , \16671 , \16672 );
and \g452646/U$2 ( \16674 , \16334 , RIe2166d8_4545);
and \g452646/U$3 ( \16675 , RIe2193d8_4577, \16380 );
nor \g452646/U$1 ( \16676 , \16674 , \16675 );
nand \g447365/U$1 ( \16677 , \16662 , \16670 , \16673 , \16676 );
nor \g446182/U$1 ( \16678 , \16657 , \16658 , \16677 );
and \g452640/U$2 ( \16679 , \16364 , RIe20b2d8_4417);
and \g452640/U$3 ( \16680 , RIe210cd8_4481, \16368 );
nor \g452640/U$1 ( \16681 , \16679 , \16680 );
nand \g445619/U$1 ( \16682 , \16656 , \16678 , \16681 );
and \g444860/U$2 ( \16683 , \16682 , \16390 );
and \g449111/U$2 ( \16684 , RIfc49b98_5861, \16337 );
and \g449111/U$3 ( \16685 , \16341 , RIfc72110_6320);
and \g449111/U$4 ( \16686 , RIfc60668_6119, \16485 );
nor \g449111/U$1 ( \16687 , \16684 , \16685 , \16686 );
and \g454946/U$2 ( \16688 , \16317 , RIf15eb58_5537);
and \g454946/U$3 ( \16689 , RIf160a48_5559, \16325 );
nor \g454946/U$1 ( \16690 , \16688 , \16689 );
not \g450126/U$3 ( \16691 , \16690 );
not \g450126/U$4 ( \16692 , \16351 );
and \g450126/U$2 ( \16693 , \16691 , \16692 );
and \g450126/U$5 ( \16694 , \16356 , RIfc60230_6116);
nor \g450126/U$1 ( \16695 , \16693 , \16694 );
and \g452637/U$2 ( \16696 , \16361 , RIfc71738_6313);
and \g452637/U$3 ( \16697 , RIfcca0b8_7321, \16364 );
nor \g452637/U$1 ( \16698 , \16696 , \16697 );
and \g452636/U$2 ( \16699 , \16368 , RIfea19e8_8183);
and \g452636/U$3 ( \16700 , RIfea1880_8182, \16371 );
nor \g452636/U$1 ( \16701 , \16699 , \16700 );
nand \g447785/U$1 ( \16702 , \16687 , \16695 , \16698 , \16701 );
and \g444860/U$3 ( \16703 , \16394 , \16702 );
nor \g444860/U$1 ( \16704 , \16683 , \16703 );
nor \g448415/U$1 ( \16705 , \16393 , \16510 );
and \g446952/U$2 ( \16706 , \16705 , RIfc45818_5813);
nor \g448433/U$1 ( \16707 , \16393 , \16513 );
and \g446952/U$3 ( \16708 , RIfcaf970_7020, \16707 );
nor \g446952/U$1 ( \16709 , \16706 , \16708 );
nor \g448432/U$1 ( \16710 , \16393 , \16320 );
and \g446951/U$2 ( \16711 , \16710 , RIfc749d8_6349);
nor \g448431/U$1 ( \16712 , \16393 , \16327 );
and \g446951/U$3 ( \16713 , RIfcd0058_7389, \16712 );
nor \g446951/U$1 ( \16714 , \16711 , \16713 );
nor \g448416/U$1 ( \16715 , \16393 , \16517 );
and \g446953/U$2 ( \16716 , \16715 , RIe2013f0_4304);
nor \g448434/U$1 ( \16717 , \16393 , \16520 );
and \g446953/U$3 ( \16718 , RIe203010_4324, \16717 );
nor \g446953/U$1 ( \16719 , \16716 , \16718 );
nand \g444625/U$1 ( \16720 , \16704 , \16709 , \16714 , \16719 );
and \g452660/U$2 ( \16721 , \16361 , RIe1bf540_3554);
and \g452660/U$3 ( \16722 , RIe1d0340_3746, \16427 );
nor \g452660/U$1 ( \16723 , \16721 , \16722 );
and \g446186/U$2 ( \16724 , RIe1d3040_3778, \16432 );
and \g446186/U$3 ( \16725 , RIe1cd640_3714, \16371 );
and \g449119/U$2 ( \16726 , RIe1e9840_4034, \16321 );
and \g449119/U$3 ( \16727 , \16326 , RIe1ec540_4066);
and \g449119/U$4 ( \16728 , RIe1c4f40_3618, \16337 );
nor \g449119/U$1 ( \16729 , \16726 , \16727 , \16728 );
and \g455373/U$2 ( \16730 , \16317 , RIe1de440_3906);
and \g455373/U$3 ( \16731 , RIe1e1140_3938, \16325 );
nor \g455373/U$1 ( \16732 , \16730 , \16731 );
not \g450133/U$3 ( \16733 , \16732 );
not \g450133/U$4 ( \16734 , \16330 );
and \g450133/U$2 ( \16735 , \16733 , \16734 );
and \g450133/U$5 ( \16736 , \16341 , RIe1c7c40_3650);
nor \g450133/U$1 ( \16737 , \16735 , \16736 );
and \g452662/U$2 ( \16738 , \16377 , RIe1e3e40_3970);
and \g452662/U$3 ( \16739 , RIe1e6b40_4002, \16313 );
nor \g452662/U$1 ( \16740 , \16738 , \16739 );
and \g452663/U$2 ( \16741 , \16334 , RIe1d8a40_3842);
and \g452663/U$3 ( \16742 , RIe1db740_3874, \16380 );
nor \g452663/U$1 ( \16743 , \16741 , \16742 );
nand \g447369/U$1 ( \16744 , \16729 , \16737 , \16740 , \16743 );
nor \g446186/U$1 ( \16745 , \16724 , \16725 , \16744 );
and \g452659/U$2 ( \16746 , \16364 , RIe1c2240_3586);
and \g452659/U$3 ( \16747 , RIe1ca940_3682, \16368 );
nor \g452659/U$1 ( \16748 , \16746 , \16747 );
nand \g445620/U$1 ( \16749 , \16723 , \16745 , \16748 );
not \g448477/U$1 ( \16750 , \16555 );
and \g444783/U$2 ( \16751 , \16749 , \16750 );
not \g448485/U$1 ( \16752 , \16586 );
and \g449116/U$2 ( \16753 , RIe179b80_2762, \16344 );
and \g449116/U$3 ( \16754 , \16356 , RIe18d680_2986);
and \g449116/U$4 ( \16755 , RIe1bc840_3522, \16398 );
nor \g449116/U$1 ( \16756 , \16753 , \16754 , \16755 );
and \g454956/U$2 ( \16757 , \16317 , RIe1a6b80_3274);
and \g454956/U$3 ( \16758 , RIe1a9880_3306, \16325 );
nor \g454956/U$1 ( \16759 , \16757 , \16758 );
not \g450130/U$3 ( \16760 , \16759 );
not \g450130/U$4 ( \16761 , \16311 );
and \g450130/U$2 ( \16762 , \16760 , \16761 );
and \g450130/U$5 ( \16763 , \16341 , RIe1d5d40_3810);
nor \g450130/U$1 ( \16764 , \16762 , \16763 );
and \g452653/U$2 ( \16765 , \16377 , RIe1a1180_3210);
and \g452653/U$3 ( \16766 , RIe1a3e80_3242, \16313 );
nor \g452653/U$1 ( \16767 , \16765 , \16766 );
and \g452655/U$2 ( \16768 , \16334 , RIe21c0d8_4609);
and \g452655/U$3 ( \16769 , RIe2274d8_4737, \16380 );
nor \g452655/U$1 ( \16770 , \16768 , \16769 );
nand \g447367/U$1 ( \16771 , \16756 , \16764 , \16767 , \16770 );
and \g444783/U$3 ( \16772 , \16752 , \16771 );
nor \g444783/U$1 ( \16773 , \16751 , \16772 );
nor \g448363/U$1 ( \16774 , \16586 , \16418 );
and \g446956/U$2 ( \16775 , \16774 , RIe171cf0_2672);
nor \g448362/U$1 ( \16776 , \16586 , \16421 );
and \g446956/U$3 ( \16777 , RIe1af6b8_3373, \16776 );
nor \g446956/U$1 ( \16778 , \16775 , \16777 );
nor \g448361/U$1 ( \16779 , \16586 , \16437 );
and \g446955/U$2 ( \16780 , \16779 , RIe1f1838_4125);
nor \g448360/U$1 ( \16781 , \16586 , \16440 );
and \g446955/U$3 ( \16782 , RIe1f8cf0_4208, \16781 );
nor \g446955/U$1 ( \16783 , \16780 , \16782 );
nor \g448359/U$1 ( \16784 , \16586 , \16428 );
and \g446954/U$2 ( \16785 , \16784 , RIe1ff938_4285);
nor \g448344/U$1 ( \16786 , \16586 , \16433 );
and \g446954/U$3 ( \16787 , RIe2058d8_4353, \16786 );
nor \g446954/U$1 ( \16788 , \16785 , \16787 );
nand \g444508/U$1 ( \16789 , \16773 , \16778 , \16783 , \16788 );
and \g446176/U$2 ( \16790 , RIe19e480_3178, \16326 );
and \g446176/U$3 ( \16791 , RIe190380_3018, \16334 );
and \g449106/U$2 ( \16792 , RIe187c80_2922, \16427 );
and \g449106/U$3 ( \16793 , \16448 , RIe18a980_2954);
and \g449106/U$4 ( \16794 , RIe195d80_3082, \16485 );
nor \g449106/U$1 ( \16795 , \16792 , \16793 , \16794 );
and \g454938/U$2 ( \16796 , \16317 , RIe182280_2858);
and \g454938/U$3 ( \16797 , RIfc615e0_6130, \16325 );
nor \g454938/U$1 ( \16798 , \16796 , \16797 );
not \g454937/U$1 ( \16799 , \16798 );
and \g450122/U$2 ( \16800 , \16799 , \16336 );
and \g450122/U$3 ( \16801 , RIfcc1148_7219, \16356 );
nor \g450122/U$1 ( \16802 , \16800 , \16801 );
and \g452619/U$2 ( \16803 , \16361 , RIe17c880_2794);
and \g452619/U$3 ( \16804 , RIe17f580_2826, \16364 );
nor \g452619/U$1 ( \16805 , \16803 , \16804 );
and \g452617/U$2 ( \16806 , \16368 , RIe184f80_2890);
and \g452617/U$3 ( \16807 , RIfcb2ee0_7058, \16371 );
nor \g452617/U$1 ( \16808 , \16806 , \16807 );
nand \g448082/U$1 ( \16809 , \16795 , \16802 , \16805 , \16808 );
nor \g446176/U$1 ( \16810 , \16790 , \16791 , \16809 );
and \g452615/U$2 ( \16811 , \16377 , RIe198a80_3114);
and \g452615/U$3 ( \16812 , RIe193080_3050, \16380 );
nor \g452615/U$1 ( \16813 , \16811 , \16812 );
and \g452614/U$2 ( \16814 , \16313 , RIfccc980_7350);
and \g452614/U$3 ( \16815 , RIe19b780_3146, \16321 );
nor \g452614/U$1 ( \16816 , \16814 , \16815 );
and \g445276/U$2 ( \16817 , \16810 , \16813 , \16816 );
nor \g445276/U$1 ( \16818 , \16817 , \16618 );
and \g446179/U$2 ( \16819 , RIfea1f88_8187, \16432 );
and \g446179/U$3 ( \16820 , RIfea1cb8_8185, \16371 );
and \g449108/U$2 ( \16821 , RIfc6adc0_6238, \16344 );
and \g449108/U$3 ( \16822 , \16356 , RIfcad0a8_6991);
and \g449108/U$4 ( \16823 , RIfc6a820_6234, \16337 );
nor \g449108/U$1 ( \16824 , \16821 , \16822 , \16823 );
and \g454944/U$2 ( \16825 , \16317 , RIfc4c898_5893);
and \g454944/U$3 ( \16826 , RIfc69038_6217, \16325 );
nor \g454944/U$1 ( \16827 , \16825 , \16826 );
not \g450123/U$3 ( \16828 , \16827 );
not \g450123/U$4 ( \16829 , \16311 );
and \g450123/U$2 ( \16830 , \16828 , \16829 );
and \g450123/U$5 ( \16831 , \16341 , RIfc60d70_6124);
nor \g450123/U$1 ( \16832 , \16830 , \16831 );
and \g452626/U$2 ( \16833 , \16377 , RIe1764a8_2723);
and \g452626/U$3 ( \16834 , RIfc6f2a8_6287, \16313 );
nor \g452626/U$1 ( \16835 , \16833 , \16834 );
and \g452628/U$2 ( \16836 , \16334 , RIfea1b50_8184);
and \g452628/U$3 ( \16837 , RIfc70388_6299, \16380 );
nor \g452628/U$1 ( \16838 , \16836 , \16837 );
nand \g447362/U$1 ( \16839 , \16824 , \16832 , \16835 , \16838 );
nor \g446179/U$1 ( \16840 , \16819 , \16820 , \16839 );
and \g452621/U$2 ( \16841 , \16364 , RIfea1e20_8186);
and \g452621/U$3 ( \16842 , RIe174450_2700, \16368 );
nor \g452621/U$1 ( \16843 , \16841 , \16842 );
and \g452623/U$2 ( \16844 , \16361 , RIf16d798_5705);
and \g452623/U$3 ( \16845 , RIfc56e88_6011, \16427 );
nor \g452623/U$1 ( \16846 , \16844 , \16845 );
and \g445279/U$2 ( \16847 , \16840 , \16843 , \16846 );
nor \g445279/U$1 ( \16848 , \16847 , \16649 );
or \g444403/U$1 ( \16849 , \16720 , \16789 , \16818 , \16848 );
and \g446173/U$2 ( \16850 , RIfcada80_6998, \16448 );
and \g446173/U$3 ( \16851 , RIe1eeca0_4094, \16361 );
and \g449101/U$2 ( \16852 , RIfc71030_6308, \16321 );
and \g449101/U$3 ( \16853 , \16328 , RIfc4ca00_5894);
and \g449101/U$4 ( \16854 , RIfcad378_6993, \16398 );
nor \g449101/U$1 ( \16855 , \16852 , \16853 , \16854 );
and \g454928/U$2 ( \16856 , \16317 , RIfc63a70_6156);
and \g454928/U$3 ( \16857 , RIfc70bf8_6305, \16325 );
nor \g454928/U$1 ( \16858 , \16856 , \16857 );
not \g450116/U$3 ( \16859 , \16858 );
not \g450116/U$4 ( \16860 , \16330 );
and \g450116/U$2 ( \16861 , \16859 , \16860 );
and \g450116/U$5 ( \16862 , \16339 , RIfcde158_7549);
nor \g450116/U$1 ( \16863 , \16861 , \16862 );
and \g452602/U$2 ( \16864 , \16377 , RIe1fad48_4231);
and \g452602/U$3 ( \16865 , RIfcde428_7551, \16313 );
nor \g452602/U$1 ( \16866 , \16864 , \16865 );
and \g452603/U$2 ( \16867 , \16334 , RIe1f62c0_4178);
and \g452603/U$3 ( \16868 , RIfca7db0_6932, \16380 );
nor \g452603/U$1 ( \16869 , \16867 , \16868 );
nand \g447361/U$1 ( \16870 , \16855 , \16863 , \16866 , \16869 );
nor \g446173/U$1 ( \16871 , \16850 , \16851 , \16870 );
and \g452600/U$2 ( \16872 , \16364 , RIfc65f00_6182);
and \g452600/U$3 ( \16873 , RIe1f3f98_4153, \16368 );
nor \g452600/U$1 ( \16874 , \16872 , \16873 );
and \g452599/U$2 ( \16875 , \16371 , RIfc6f578_6289);
and \g452599/U$3 ( \16876 , RIfc6fde8_6295, \16427 );
nor \g452599/U$1 ( \16877 , \16875 , \16876 );
and \g445272/U$2 ( \16878 , \16871 , \16874 , \16877 );
nor \g445272/U$1 ( \16879 , \16878 , \16480 );
and \g446174/U$2 ( \16880 , RIfc69308_6219, \16328 );
and \g446174/U$3 ( \16881 , RIe1b4578_3429, \16334 );
and \g449104/U$2 ( \16882 , RIfcb9c90_7136, \16398 );
and \g449104/U$3 ( \16883 , \16341 , RIfc9f818_6837);
and \g449104/U$4 ( \16884 , RIfc69740_6222, \16344 );
nor \g449104/U$1 ( \16885 , \16882 , \16883 , \16884 );
and \g454932/U$2 ( \16886 , \16317 , RIf148088_5279);
and \g454932/U$3 ( \16887 , RIfccf950_7384, \16325 );
nor \g454932/U$1 ( \16888 , \16886 , \16887 );
not \g450120/U$3 ( \16889 , \16888 );
not \g450120/U$4 ( \16890 , \16351 );
and \g450120/U$2 ( \16891 , \16889 , \16890 );
and \g450120/U$5 ( \16892 , \16354 , RIfccd628_7359);
nor \g450120/U$1 ( \16893 , \16891 , \16892 );
and \g452610/U$2 ( \16894 , \16361 , RIe1ab770_3328);
and \g452610/U$3 ( \16895 , RIe1acf58_3345, \16364 );
nor \g452610/U$1 ( \16896 , \16894 , \16895 );
and \g452609/U$2 ( \16897 , \16368 , RIe1b1710_3396);
and \g452609/U$3 ( \16898 , RIe1b3060_3414, \16371 );
nor \g452609/U$1 ( \16899 , \16897 , \16898 );
nand \g447783/U$1 ( \16900 , \16885 , \16893 , \16896 , \16899 );
nor \g446174/U$1 ( \16901 , \16880 , \16881 , \16900 );
and \g452608/U$2 ( \16902 , \16377 , RIe1b7db8_3469);
and \g452608/U$3 ( \16903 , RIe1b5bf8_3445, \16380 );
nor \g452608/U$1 ( \16904 , \16902 , \16903 );
and \g452607/U$2 ( \16905 , \16313 , RIe1b9f78_3493);
and \g452607/U$3 ( \16906 , RIfccba08_7339, \16321 );
nor \g452607/U$1 ( \16907 , \16905 , \16906 );
and \g445273/U$2 ( \16908 , \16901 , \16904 , \16907 );
not \g448461/U$1 ( \16909 , \16477 );
nor \g445273/U$1 ( \16910 , \16908 , \16909 );
or \g444178/U$1 ( \16911 , \16849 , \16879 , \16910 );
_DC \g33e7/U$1 ( \16912 , \16911 , \16652 );
and \g446763/U$2 ( \16913 , \16419 , RIfc7c430_6436);
and \g446763/U$3 ( \16914 , RIf15aaa8_5491, \16422 );
nor \g446763/U$1 ( \16915 , \16913 , \16914 );
and \g445979/U$2 ( \16916 , RIfc77f48_6387, \16341 );
and \g445979/U$3 ( \16917 , RIfc41fd8_5773, \16337 );
and \g448851/U$2 ( \16918 , RIfc59cf0_6044, \16319 );
and \g448851/U$3 ( \16919 , \16485 , RIfcd19a8_7407);
and \g448851/U$4 ( \16920 , RIfc79cd0_6408, \16356 );
nor \g448851/U$1 ( \16921 , \16918 , \16919 , \16920 );
and \g453097/U$2 ( \16922 , \16368 , RIfea46e8_8215);
and \g453097/U$3 ( \16923 , RIfea4580_8214, \16371 );
nor \g453097/U$1 ( \16924 , \16922 , \16923 );
and \g454188/U$2 ( \16925 , \16317 , RIf15e888_5535);
and \g454188/U$3 ( \16926 , RIf160778_5557, \16325 );
nor \g454188/U$1 ( \16927 , \16925 , \16926 );
not \g449874/U$3 ( \16928 , \16927 );
not \g449874/U$4 ( \16929 , \16351 );
and \g449874/U$2 ( \16930 , \16928 , \16929 );
and \g449874/U$5 ( \16931 , \16326 , RIfc7b080_6422);
nor \g449874/U$1 ( \16932 , \16930 , \16931 );
and \g451779/U$2 ( \16933 , \16334 , RIf162230_5576);
and \g451779/U$3 ( \16934 , RIfcc81c8_7299, \16380 );
nor \g451779/U$1 ( \16935 , \16933 , \16934 );
nand \g447648/U$1 ( \16936 , \16921 , \16924 , \16932 , \16935 );
nor \g445979/U$1 ( \16937 , \16916 , \16917 , \16936 );
not \g444815/U$3 ( \16938 , \16937 );
not \g444815/U$4 ( \16939 , \16393 );
and \g444815/U$2 ( \16940 , \16938 , \16939 );
and \g445981/U$2 ( \16941 , RIfc87290_6560, \16356 );
and \g445981/U$3 ( \16942 , RIe184cb0_2888, \16368 );
and \g448857/U$2 ( \16943 , RIe1879b0_2920, \16427 );
and \g448857/U$3 ( \16944 , \16398 , RIe181fb0_2856);
and \g448857/U$4 ( \16945 , RIfc83a50_6520, \16341 );
nor \g448857/U$1 ( \16946 , \16943 , \16944 , \16945 );
and \g451795/U$2 ( \16947 , \16361 , RIe17c5b0_2792);
and \g451795/U$3 ( \16948 , RIe17f2b0_2824, \16364 );
nor \g451795/U$1 ( \16949 , \16947 , \16948 );
and \g452648/U$2 ( \16950 , \16377 , RIe1987b0_3112);
and \g452648/U$3 ( \16951 , RIfc9cf50_6808, \16313 );
nor \g452648/U$1 ( \16952 , \16950 , \16951 );
and \g454869/U$2 ( \16953 , \16317 , RIe19b4b0_3144);
and \g454869/U$3 ( \16954 , RIe19e1b0_3176, \16325 );
nor \g454869/U$1 ( \16955 , \16953 , \16954 );
not \g450098/U$3 ( \16956 , \16955 );
not \g450098/U$4 ( \16957 , \16311 );
and \g450098/U$2 ( \16958 , \16956 , \16957 );
and \g450098/U$5 ( \16959 , \16448 , RIe18a6b0_2952);
nor \g450098/U$1 ( \16960 , \16958 , \16959 );
nand \g447649/U$1 ( \16961 , \16946 , \16949 , \16952 , \16960 );
nor \g445981/U$1 ( \16962 , \16941 , \16942 , \16961 );
and \g451788/U$2 ( \16963 , \16334 , RIe1900b0_3016);
and \g451788/U$3 ( \16964 , RIfc842c0_6526, \16371 );
nor \g451788/U$1 ( \16965 , \16963 , \16964 );
and \g452827/U$2 ( \16966 , \16380 , RIe192db0_3048);
and \g452827/U$3 ( \16967 , RIe195ab0_3080, \16485 );
nor \g452827/U$1 ( \16968 , \16966 , \16967 );
and \g445137/U$2 ( \16969 , \16962 , \16965 , \16968 );
nor \g445137/U$1 ( \16970 , \16969 , \16618 );
nor \g444815/U$1 ( \16971 , \16940 , \16970 );
and \g446764/U$2 ( \16972 , \16715 , RIfea4418_8213);
and \g446764/U$3 ( \16973 , RIfea9b48_8247, \16717 );
nor \g446764/U$1 ( \16974 , \16972 , \16973 );
nand \g444424/U$1 ( \16975 , \16915 , \16971 , \16974 );
and \g451817/U$2 ( \16976 , \16380 , RIe1b5928_3443);
and \g451817/U$3 ( \16977 , RIfca6190_6912, \16485 );
nor \g451817/U$1 ( \16978 , \16976 , \16977 );
and \g445988/U$2 ( \16979 , RIfcc20c0_7230, \16354 );
and \g445988/U$3 ( \16980 , RIe1b1440_3394, \16368 );
and \g448864/U$2 ( \16981 , RIfcc5090_7264, \16427 );
and \g448864/U$3 ( \16982 , \16337 , RIfcb9588_7131);
and \g448864/U$4 ( \16983 , RIfcd5350_7448, \16341 );
nor \g448864/U$1 ( \16984 , \16981 , \16982 , \16983 );
and \g451822/U$2 ( \16985 , \16361 , RIe1ab4a0_3326);
and \g451822/U$3 ( \16986 , RIe1acc88_3343, \16364 );
nor \g451822/U$1 ( \16987 , \16985 , \16986 );
and \g451821/U$2 ( \16988 , \16377 , RIe1b7ae8_3467);
and \g451821/U$3 ( \16989 , RIe1b9ca8_3491, \16313 );
nor \g451821/U$1 ( \16990 , \16988 , \16989 );
and \g454753/U$2 ( \16991 , \16317 , RIfcbef88_7195);
and \g454753/U$3 ( \16992 , RIfc784e8_6391, \16325 );
nor \g454753/U$1 ( \16993 , \16991 , \16992 );
not \g449888/U$3 ( \16994 , \16993 );
not \g449888/U$4 ( \16995 , \16311 );
and \g449888/U$2 ( \16996 , \16994 , \16995 );
and \g449888/U$5 ( \16997 , \16432 , RIfcb81d8_7117);
nor \g449888/U$1 ( \16998 , \16996 , \16997 );
nand \g447653/U$1 ( \16999 , \16984 , \16987 , \16990 , \16998 );
nor \g445988/U$1 ( \17000 , \16979 , \16980 , \16999 );
and \g451819/U$2 ( \17001 , \16334 , RIe1b4410_3428);
and \g451819/U$3 ( \17002 , RIe1b2d90_3412, \16371 );
nor \g451819/U$1 ( \17003 , \17001 , \17002 );
nand \g445573/U$1 ( \17004 , \16978 , \17000 , \17003 );
and \g444913/U$2 ( \17005 , \17004 , \16477 );
and \g448859/U$2 ( \17006 , RIe1a68b0_3272, \16321 );
and \g448859/U$3 ( \17007 , \16328 , RIe1a95b0_3304);
and \g448859/U$4 ( \17008 , RIe1798b0_2760, \16485 );
nor \g448859/U$1 ( \17009 , \17006 , \17007 , \17008 );
and \g454709/U$2 ( \17010 , \16317 , RIe1ff668_4283);
and \g454709/U$3 ( \17011 , RIe205608_4351, \16325 );
nor \g454709/U$1 ( \17012 , \17010 , \17011 );
not \g449966/U$3 ( \17013 , \17012 );
not \g449966/U$4 ( \17014 , \16351 );
and \g449966/U$2 ( \17015 , \17013 , \17014 );
and \g449966/U$5 ( \17016 , \16356 , RIe18d3b0_2984);
nor \g449966/U$1 ( \17017 , \17015 , \17016 );
and \g451925/U$2 ( \17018 , \16377 , RIe1a0eb0_3208);
and \g451925/U$3 ( \17019 , RIe1a3bb0_3240, \16313 );
nor \g451925/U$1 ( \17020 , \17018 , \17019 );
and \g451812/U$2 ( \17021 , \16368 , RIe1f1568_4123);
and \g451812/U$3 ( \17022 , RIe1f8a20_4206, \16371 );
nor \g451812/U$1 ( \17023 , \17021 , \17022 );
nand \g447651/U$1 ( \17024 , \17009 , \17017 , \17020 , \17023 );
and \g444913/U$3 ( \17025 , \16752 , \17024 );
nor \g444913/U$1 ( \17026 , \17005 , \17025 );
nor \g448346/U$1 ( \17027 , \16586 , \16397 );
and \g446769/U$2 ( \17028 , \17027 , RIe1bc570_3520);
nor \g448371/U$1 ( \17029 , \16586 , \16513 );
and \g446769/U$3 ( \17030 , RIe227208_4735, \17029 );
nor \g446769/U$1 ( \17031 , \17028 , \17030 );
nor \g448372/U$1 ( \17032 , \16586 , \16510 );
and \g446768/U$2 ( \17033 , \17032 , RIe21be08_4607);
nor \g448345/U$1 ( \17034 , \16586 , \16340 );
and \g446768/U$3 ( \17035 , RIe1d5a70_3808, \17034 );
nor \g446768/U$1 ( \17036 , \17033 , \17035 );
and \g446770/U$2 ( \17037 , \16774 , RIe171a20_2670);
and \g446770/U$3 ( \17038 , RIe1af3e8_3371, \16776 );
nor \g446770/U$1 ( \17039 , \17037 , \17038 );
nand \g444594/U$1 ( \17040 , \17026 , \17031 , \17036 , \17039 );
and \g445969/U$2 ( \17041 , RIe177420_2734, \16313 );
and \g445969/U$3 ( \17042 , RIfc472d0_5832, \16361 );
and \g448841/U$2 ( \17043 , RIfc9e030_6820, \16319 );
and \g448841/U$3 ( \17044 , \16344 , RIfcc4820_7258);
and \g448841/U$4 ( \17045 , RIfc4f700_5926, \16356 );
nor \g448841/U$1 ( \17046 , \17043 , \17044 , \17045 );
and \g451747/U$2 ( \17047 , \16368 , RIe174180_2698);
and \g451747/U$3 ( \17048 , RIfc812f0_6492, \16371 );
nor \g451747/U$1 ( \17049 , \17047 , \17048 );
and \g455034/U$2 ( \17050 , \16317 , RIee3b308_5132);
and \g455034/U$3 ( \17051 , RIee3c6b8_5146, \16325 );
nor \g455034/U$1 ( \17052 , \17050 , \17051 );
not \g449865/U$3 ( \17053 , \17052 );
not \g449865/U$4 ( \17054 , \16351 );
and \g449865/U$2 ( \17055 , \17053 , \17054 );
and \g449865/U$5 ( \17056 , \16328 , RIfc9d0b8_6809);
nor \g449865/U$1 ( \17057 , \17055 , \17056 );
and \g451745/U$2 ( \17058 , \16334 , RIfce8040_7662);
and \g451745/U$3 ( \17059 , RIfc4fb38_5929, \16380 );
nor \g451745/U$1 ( \17060 , \17058 , \17059 );
nand \g447638/U$1 ( \17061 , \17046 , \17049 , \17057 , \17060 );
nor \g445969/U$1 ( \17062 , \17041 , \17042 , \17061 );
and \g451742/U$2 ( \17063 , \16364 , RIfc46a60_5826);
and \g451742/U$3 ( \17064 , RIfcd3028_7423, \16341 );
nor \g451742/U$1 ( \17065 , \17063 , \17064 );
and \g451739/U$2 ( \17066 , \16398 , RIfc7f400_6470);
and \g451739/U$3 ( \17067 , RIe176340_2722, \16377 );
nor \g451739/U$1 ( \17068 , \17066 , \17067 );
and \g445124/U$2 ( \17069 , \17062 , \17065 , \17068 );
nor \g445124/U$1 ( \17070 , \17069 , \16649 );
and \g445973/U$2 ( \17071 , RIfc97c58_6749, \16356 );
and \g445973/U$3 ( \17072 , RIe210a08_4479, \16368 );
and \g448846/U$2 ( \17073 , RIe213708_4511, \16427 );
and \g448846/U$3 ( \17074 , \16398 , RIe20dd08_4447);
and \g448846/U$4 ( \17075 , RIfca4570_6892, \16339 );
nor \g448846/U$1 ( \17076 , \17073 , \17074 , \17075 );
and \g451770/U$2 ( \17077 , \16361 , RIe208308_4383);
and \g451770/U$3 ( \17078 , RIe20b008_4415, \16364 );
nor \g451770/U$1 ( \17079 , \17077 , \17078 );
and \g453632/U$2 ( \17080 , \16377 , RIe221808_4671);
and \g453632/U$3 ( \17081 , RIfc7d3a8_6447, \16313 );
nor \g453632/U$1 ( \17082 , \17080 , \17081 );
and \g455167/U$2 ( \17083 , \16317 , RIe224508_4703);
and \g455167/U$3 ( \17084 , RIf16cc58_5697, \16325 );
nor \g455167/U$1 ( \17085 , \17083 , \17084 );
not \g449870/U$3 ( \17086 , \17085 );
not \g449870/U$4 ( \17087 , \16311 );
and \g449870/U$2 ( \17088 , \17086 , \17087 );
and \g449870/U$5 ( \17089 , \16448 , RIfcdbe30_7524);
nor \g449870/U$1 ( \17090 , \17088 , \17089 );
nand \g447644/U$1 ( \17091 , \17076 , \17079 , \17082 , \17090 );
nor \g445973/U$1 ( \17092 , \17071 , \17072 , \17091 );
and \g451759/U$2 ( \17093 , \16334 , RIe216408_4543);
and \g451759/U$3 ( \17094 , RIf169580_5658, \16371 );
nor \g451759/U$1 ( \17095 , \17093 , \17094 );
and \g451757/U$2 ( \17096 , \16380 , RIe219108_4575);
and \g451757/U$3 ( \17097 , RIe21eb08_4639, \16485 );
nor \g451757/U$1 ( \17098 , \17096 , \17097 );
and \g445128/U$2 ( \17099 , \17092 , \17095 , \17098 );
nor \g445128/U$1 ( \17100 , \17099 , \16389 );
or \g444298/U$1 ( \17101 , \16975 , \17040 , \17070 , \17100 );
and \g445961/U$2 ( \17102 , RIfc4a840_5870, \16354 );
and \g445961/U$3 ( \17103 , RIe1f5ff0_4176, \16334 );
and \g448829/U$2 ( \17104 , RIf157f10_5460, \16321 );
and \g448829/U$3 ( \17105 , \16328 , RIf159158_5473);
and \g448829/U$4 ( \17106 , RIf151f70_5392, \16427 );
nor \g448829/U$1 ( \17107 , \17104 , \17105 , \17106 );
and \g451714/U$2 ( \17108 , \16361 , RIe1ee9d0_4092);
and \g451714/U$3 ( \17109 , RIfca9ca0_6954, \16364 );
nor \g451714/U$1 ( \17110 , \17108 , \17109 );
and \g451710/U$2 ( \17111 , \16377 , RIe1faa78_4229);
and \g451710/U$3 ( \17112 , RIfcae890_7008, \16313 );
nor \g451710/U$1 ( \17113 , \17111 , \17112 );
and \g454845/U$2 ( \17114 , \16317 , RIfc6d250_6264);
and \g454845/U$3 ( \17115 , RIfc68ed0_6216, \16325 );
nor \g454845/U$1 ( \17116 , \17114 , \17115 );
not \g454844/U$1 ( \17117 , \17116 );
and \g449857/U$2 ( \17118 , \17117 , \16336 );
and \g449857/U$3 ( \17119 , RIf153758_5409, \16448 );
nor \g449857/U$1 ( \17120 , \17118 , \17119 );
nand \g448051/U$1 ( \17121 , \17107 , \17110 , \17113 , \17120 );
nor \g445961/U$1 ( \17122 , \17102 , \17103 , \17121 );
and \g451703/U$2 ( \17123 , \16371 , RIfccb468_7335);
and \g451703/U$3 ( \17124 , RIfce0e58_7581, \16380 );
nor \g451703/U$1 ( \17125 , \17123 , \17124 );
and \g451706/U$2 ( \17126 , \16368 , RIe1f3cc8_4151);
and \g451706/U$3 ( \17127 , RIfc4ed28_5919, \16344 );
nor \g451706/U$1 ( \17128 , \17126 , \17127 );
and \g445116/U$2 ( \17129 , \17122 , \17125 , \17128 );
nor \g445116/U$1 ( \17130 , \17129 , \16480 );
and \g445965/U$2 ( \17131 , RIe1c7970_3648, \16341 );
and \g445965/U$3 ( \17132 , RIe1e3b70_3968, \16377 );
and \g448836/U$2 ( \17133 , RIe1d0070_3744, \16427 );
and \g448836/U$3 ( \17134 , \16448 , RIe1d2d70_3776);
and \g448836/U$4 ( \17135 , RIe1e9570_4032, \16321 );
nor \g448836/U$1 ( \17136 , \17133 , \17134 , \17135 );
and \g451731/U$2 ( \17137 , \16368 , RIe1ca670_3680);
and \g451731/U$3 ( \17138 , RIe1cd370_3712, \16371 );
nor \g451731/U$1 ( \17139 , \17137 , \17138 );
and \g454142/U$2 ( \17140 , \16317 , RIe1de170_3904);
and \g454142/U$3 ( \17141 , RIe1e0e70_3936, \16325 );
nor \g454142/U$1 ( \17142 , \17140 , \17141 );
not \g449860/U$3 ( \17143 , \17142 );
not \g449860/U$4 ( \17144 , \16330 );
and \g449860/U$2 ( \17145 , \17143 , \17144 );
and \g449860/U$5 ( \17146 , \16328 , RIe1ec270_4064);
nor \g449860/U$1 ( \17147 , \17145 , \17146 );
and \g451728/U$2 ( \17148 , \16334 , RIe1d8770_3840);
and \g451728/U$3 ( \17149 , RIe1db470_3872, \16380 );
nor \g451728/U$1 ( \17150 , \17148 , \17149 );
nand \g447635/U$1 ( \17151 , \17136 , \17139 , \17147 , \17150 );
nor \g445965/U$1 ( \17152 , \17131 , \17132 , \17151 );
and \g451723/U$2 ( \17153 , \16361 , RIe1bf270_3552);
and \g451723/U$3 ( \17154 , RIe1e6870_4000, \16313 );
nor \g451723/U$1 ( \17155 , \17153 , \17154 );
and \g452407/U$2 ( \17156 , \16364 , RIe1c1f70_3584);
and \g452407/U$3 ( \17157 , RIe1c4c70_3616, \16337 );
nor \g452407/U$1 ( \17158 , \17156 , \17157 );
and \g445121/U$2 ( \17159 , \17152 , \17155 , \17158 );
nor \g445121/U$1 ( \17160 , \17159 , \16555 );
or \g444183/U$1 ( \17161 , \17101 , \17130 , \17160 );
_DC \g346c/U$1 ( \17162 , \17161 , \16652 );
and \g452156/U$2 ( \17163 , \16377 , RIe2216a0_4670);
and \g452156/U$3 ( \17164 , RIe218fa0_4574, \16380 );
nor \g452156/U$1 ( \17165 , \17163 , \17164 );
and \g446079/U$2 ( \17166 , RIe2243a0_4702, \16321 );
and \g446079/U$3 ( \17167 , RIfca0358_6845, \16313 );
and \g448979/U$2 ( \17168 , RIe20dba0_4446, \16398 );
and \g448979/U$3 ( \17169 , \16339 , RIfc8bfe8_6615);
and \g448979/U$4 ( \17170 , RIe21e9a0_4638, \16344 );
nor \g448979/U$1 ( \17171 , \17168 , \17169 , \17170 );
and \g454431/U$2 ( \17172 , \16317 , RIe2135a0_4510);
and \g454431/U$3 ( \17173 , RIfc456b0_5812, \16325 );
nor \g454431/U$1 ( \17174 , \17172 , \17173 );
not \g449570/U$3 ( \17175 , \17174 );
not \g449570/U$4 ( \17176 , \16351 );
and \g449570/U$2 ( \17177 , \17175 , \17176 );
and \g449570/U$5 ( \17178 , \16356 , RIfc9a688_6779);
nor \g449570/U$1 ( \17179 , \17177 , \17178 );
and \g452165/U$2 ( \17180 , \16361 , RIe2081a0_4382);
and \g452165/U$3 ( \17181 , RIe20aea0_4414, \16364 );
nor \g452165/U$1 ( \17182 , \17180 , \17181 );
and \g453698/U$2 ( \17183 , \16368 , RIe2108a0_4478);
and \g453698/U$3 ( \17184 , RIf169418_5657, \16371 );
nor \g453698/U$1 ( \17185 , \17183 , \17184 );
nand \g447718/U$1 ( \17186 , \17171 , \17179 , \17182 , \17185 );
nor \g446079/U$1 ( \17187 , \17166 , \17167 , \17186 );
and \g452154/U$2 ( \17188 , \16334 , RIe2162a0_4542);
and \g452154/U$3 ( \17189 , RIfc48c20_5850, \16328 );
nor \g452154/U$1 ( \17190 , \17188 , \17189 );
nand \g445593/U$1 ( \17191 , \17165 , \17187 , \17190 );
and \g444857/U$2 ( \17192 , \17191 , \16390 );
and \g448973/U$2 ( \17193 , RIfc487e8_5847, \16485 );
and \g448973/U$3 ( \17194 , \16356 , RIfce2910_7600);
and \g448973/U$4 ( \17195 , RIfcbdbd8_7181, \16398 );
nor \g448973/U$1 ( \17196 , \17193 , \17194 , \17195 );
and \g454143/U$2 ( \17197 , \16317 , RIfc7f568_6471);
and \g454143/U$3 ( \17198 , RIfc8c9c0_6622, \16325 );
nor \g454143/U$1 ( \17199 , \17197 , \17198 );
not \g449988/U$3 ( \17200 , \17199 );
not \g449988/U$4 ( \17201 , \16311 );
and \g449988/U$2 ( \17202 , \17200 , \17201 );
and \g449988/U$5 ( \17203 , \16341 , RIfc580d0_6024);
nor \g449988/U$1 ( \17204 , \17202 , \17203 );
and \g452147/U$2 ( \17205 , \16377 , RIe201120_4302);
and \g452147/U$3 ( \17206 , RIe202d40_4322, \16313 );
nor \g452147/U$1 ( \17207 , \17205 , \17206 );
and \g452148/U$2 ( \17208 , \16334 , RIfc992d8_6765);
and \g452148/U$3 ( \17209 , RIfc46d30_5828, \16380 );
nor \g452148/U$1 ( \17210 , \17208 , \17209 );
nand \g447242/U$1 ( \17211 , \17196 , \17204 , \17207 , \17210 );
and \g444857/U$3 ( \17212 , \16394 , \17211 );
nor \g444857/U$1 ( \17213 , \17192 , \17212 );
and \g446849/U$2 ( \17214 , \16419 , RIfce01b0_7572);
and \g446849/U$3 ( \17215 , RIfc8dd70_6636, \16422 );
nor \g446849/U$1 ( \17216 , \17214 , \17215 );
and \g446848/U$2 ( \17217 , \16429 , RIfc44a08_5803);
and \g446848/U$3 ( \17218 , RIfca2680_6870, \16434 );
nor \g446848/U$1 ( \17219 , \17217 , \17218 );
and \g446850/U$2 ( \17220 , \16438 , RIe1fbf90_4244);
and \g446850/U$3 ( \17221 , RIe1fd1d8_4257, \16441 );
nor \g446850/U$1 ( \17222 , \17220 , \17221 );
nand \g444606/U$1 ( \17223 , \17213 , \17216 , \17219 , \17222 );
and \g452126/U$2 ( \17224 , \16377 , RIfec5910_8368);
and \g452126/U$3 ( \17225 , RIe1b57c0_3442, \16380 );
nor \g452126/U$1 ( \17226 , \17224 , \17225 );
and \g446073/U$2 ( \17227 , RIfc78d58_6397, \16321 );
and \g446073/U$3 ( \17228 , RIe1b9b40_3490, \16313 );
and \g448970/U$2 ( \17229 , RIfec5a78_8369, \16427 );
and \g448970/U$3 ( \17230 , \16432 , RIf1492d0_5292);
and \g448970/U$4 ( \17231 , RIfcd51e8_7447, \16344 );
nor \g448970/U$1 ( \17232 , \17229 , \17230 , \17231 );
and \g454750/U$2 ( \17233 , \16317 , RIf146a08_5263);
and \g454750/U$3 ( \17234 , RIfec5640_8366, \16325 );
nor \g454750/U$1 ( \17235 , \17233 , \17234 );
not \g454749/U$1 ( \17236 , \17235 );
and \g449983/U$2 ( \17237 , \17236 , \16336 );
and \g449983/U$3 ( \17238 , RIfc78a88_6395, \16356 );
nor \g449983/U$1 ( \17239 , \17237 , \17238 );
and \g452134/U$2 ( \17240 , \16361 , RIfea1178_8177);
and \g452134/U$3 ( \17241 , RIfec57a8_8367, \16364 );
nor \g452134/U$1 ( \17242 , \17240 , \17241 );
and \g452132/U$2 ( \17243 , \16368 , RIe1b12d8_3393);
and \g452132/U$3 ( \17244 , RIe1b2c28_3411, \16371 );
nor \g452132/U$1 ( \17245 , \17243 , \17244 );
nand \g448065/U$1 ( \17246 , \17232 , \17239 , \17242 , \17245 );
nor \g446073/U$1 ( \17247 , \17227 , \17228 , \17246 );
and \g452125/U$2 ( \17248 , \16334 , RIfea1010_8176);
and \g452125/U$3 ( \17249 , RIf14cf48_5335, \16326 );
nor \g452125/U$1 ( \17250 , \17248 , \17249 );
nand \g445591/U$1 ( \17251 , \17226 , \17247 , \17250 );
and \g444915/U$2 ( \17252 , \17251 , \16477 );
and \g449311/U$2 ( \17253 , RIfc90368_6663, \16321 );
and \g449311/U$3 ( \17254 , \16328 , RIfc7bbc0_6430);
and \g449311/U$4 ( \17255 , RIfcdb728_7519, \16398 );
nor \g449311/U$1 ( \17256 , \17253 , \17254 , \17255 );
and \g454665/U$2 ( \17257 , \16317 , RIfc43ec8_5795);
and \g454665/U$3 ( \17258 , RIfcd8b90_7488, \16325 );
nor \g454665/U$1 ( \17259 , \17257 , \17258 );
not \g449979/U$3 ( \17260 , \17259 );
not \g449979/U$4 ( \17261 , \16330 );
and \g449979/U$2 ( \17262 , \17260 , \17261 );
and \g449979/U$5 ( \17263 , \16339 , RIfc91010_6672);
nor \g449979/U$1 ( \17264 , \17262 , \17263 );
and \g452117/U$2 ( \17265 , \16377 , RIe1fa910_4228);
and \g452117/U$3 ( \17266 , RIfc7b8f0_6428, \16313 );
nor \g452117/U$1 ( \17267 , \17265 , \17266 );
and \g452120/U$2 ( \17268 , \16334 , RIe1f5e88_4175);
and \g452120/U$3 ( \17269 , RIfc7b788_6427, \16380 );
nor \g452120/U$1 ( \17270 , \17268 , \17269 );
nand \g447333/U$1 ( \17271 , \17256 , \17264 , \17267 , \17270 );
and \g444915/U$3 ( \17272 , \16481 , \17271 );
nor \g444915/U$1 ( \17273 , \17252 , \17272 );
nor \g448451/U$1 ( \17274 , \16480 , \16428 );
and \g446839/U$2 ( \17275 , \17274 , RIfc90d40_6670);
nor \g448446/U$1 ( \17276 , \16480 , \16433 );
and \g446839/U$3 ( \17277 , RIfc7b350_6424, \17276 );
nor \g446839/U$1 ( \17278 , \17275 , \17277 );
nor \g448455/U$1 ( \17279 , \16480 , \16437 );
and \g446844/U$2 ( \17280 , \17279 , RIe1f3b60_4150);
nor \g448454/U$1 ( \17281 , \16480 , \16440 );
and \g446844/U$3 ( \17282 , RIfca3490_6880, \17281 );
nor \g446844/U$1 ( \17283 , \17280 , \17282 );
nor \g448453/U$1 ( \17284 , \16480 , \16418 );
and \g446843/U$2 ( \17285 , \17284 , RIe1ee868_4091);
nor \g448452/U$1 ( \17286 , \16480 , \16421 );
and \g446843/U$3 ( \17287 , RIfcd8758_7485, \17286 );
nor \g446843/U$1 ( \17288 , \17285 , \17287 );
nand \g444604/U$1 ( \17289 , \17273 , \17278 , \17283 , \17288 );
and \g446059/U$2 ( \17290 , RIee3c550_5145, \16432 );
and \g446059/U$3 ( \17291 , RIee3a0c0_5119, \16371 );
and \g448957/U$2 ( \17292 , RIfc995a8_6767, \16319 );
and \g448957/U$3 ( \17293 , \16328 , RIfcb5d48_7091);
and \g448957/U$4 ( \17294 , RIfcbc288_7163, \16337 );
nor \g448957/U$1 ( \17295 , \17292 , \17293 , \17294 );
and \g454467/U$2 ( \17296 , \16317 , RIfcd2bf0_7420);
and \g454467/U$3 ( \17297 , RIfc54188_5979, \16325 );
nor \g454467/U$1 ( \17298 , \17296 , \17297 );
not \g449973/U$3 ( \17299 , \17298 );
not \g449973/U$4 ( \17300 , \16330 );
and \g449973/U$2 ( \17301 , \17299 , \17300 );
and \g449973/U$5 ( \17302 , \16339 , RIfc46628_5823);
nor \g449973/U$1 ( \17303 , \17301 , \17302 );
and \g452168/U$2 ( \17304 , \16377 , RIe1761d8_2721);
and \g452168/U$3 ( \17305 , RIfc9a3b8_6777, \16313 );
nor \g452168/U$1 ( \17306 , \17304 , \17305 );
and \g452091/U$2 ( \17307 , \16334 , RIfc7dee8_6455);
and \g452091/U$3 ( \17308 , RIfc8b778_6609, \16380 );
nor \g452091/U$1 ( \17309 , \17307 , \17308 );
nand \g447331/U$1 ( \17310 , \17295 , \17303 , \17306 , \17309 );
nor \g446059/U$1 ( \17311 , \17290 , \17291 , \17310 );
and \g453209/U$2 ( \17312 , \16364 , RIf16e710_5716);
and \g453209/U$3 ( \17313 , RIfeaba38_8269, \16368 );
nor \g453209/U$1 ( \17314 , \17312 , \17313 );
and \g452085/U$2 ( \17315 , \16361 , RIfc8fdc8_6659);
and \g452085/U$3 ( \17316 , RIfc8c420_6618, \16427 );
nor \g452085/U$1 ( \17317 , \17315 , \17316 );
and \g445194/U$2 ( \17318 , \17311 , \17314 , \17317 );
nor \g445194/U$1 ( \17319 , \17318 , \16649 );
and \g446063/U$2 ( \17320 , RIe187848_2919, \16427 );
and \g446063/U$3 ( \17321 , RIe184b48_2887, \16368 );
and \g448962/U$2 ( \17322 , RIe195948_3079, \16344 );
and \g448962/U$3 ( \17323 , \16354 , RIfc7efc8_6467);
and \g448962/U$4 ( \17324 , RIe181e48_2855, \16398 );
nor \g448962/U$1 ( \17325 , \17322 , \17323 , \17324 );
and \g455114/U$2 ( \17326 , \16317 , RIe19b348_3143);
and \g455114/U$3 ( \17327 , RIe19e048_3175, \16325 );
nor \g455114/U$1 ( \17328 , \17326 , \17327 );
not \g449976/U$3 ( \17329 , \17328 );
not \g449976/U$4 ( \17330 , \16311 );
and \g449976/U$2 ( \17331 , \17329 , \17330 );
and \g449976/U$5 ( \17332 , \16341 , RIfc98d38_6761);
nor \g449976/U$1 ( \17333 , \17331 , \17332 );
and \g452103/U$2 ( \17334 , \16377 , RIe198648_3111);
and \g452103/U$3 ( \17335 , RIfcc3ce0_7250, \16313 );
nor \g452103/U$1 ( \17336 , \17334 , \17335 );
and \g452106/U$2 ( \17337 , \16334 , RIe18ff48_3015);
and \g452106/U$3 ( \17338 , RIe192c48_3047, \16380 );
nor \g452106/U$1 ( \17339 , \17337 , \17338 );
nand \g447332/U$1 ( \17340 , \17325 , \17333 , \17336 , \17339 );
nor \g446063/U$1 ( \17341 , \17320 , \17321 , \17340 );
and \g452099/U$2 ( \17342 , \16361 , RIe17c448_2791);
and \g452099/U$3 ( \17343 , RIe18a548_2951, \16448 );
nor \g452099/U$1 ( \17344 , \17342 , \17343 );
and \g452097/U$2 ( \17345 , \16364 , RIe17f148_2823);
and \g452097/U$3 ( \17346 , RIfc46790_5824, \16371 );
nor \g452097/U$1 ( \17347 , \17345 , \17346 );
and \g445195/U$2 ( \17348 , \17341 , \17344 , \17347 );
nor \g445195/U$1 ( \17349 , \17348 , \16618 );
or \g444394/U$1 ( \17350 , \17223 , \17289 , \17319 , \17349 );
and \g446052/U$2 ( \17351 , RIe1e9408_4031, \16321 );
and \g446052/U$3 ( \17352 , RIe1e6708_3999, \16313 );
and \g448948/U$2 ( \17353 , RIe1c4b08_3615, \16398 );
and \g448948/U$3 ( \17354 , \16341 , RIe1c7808_3647);
and \g448948/U$4 ( \17355 , RIe1de008_3903, \16485 );
nor \g448948/U$1 ( \17356 , \17353 , \17354 , \17355 );
and \g454713/U$2 ( \17357 , \16317 , RIe1cff08_3743);
and \g454713/U$3 ( \17358 , RIe1d2c08_3775, \16325 );
nor \g454713/U$1 ( \17359 , \17357 , \17358 );
not \g449965/U$3 ( \17360 , \17359 );
not \g449965/U$4 ( \17361 , \16351 );
and \g449965/U$2 ( \17362 , \17360 , \17361 );
and \g449965/U$5 ( \17363 , \16356 , RIe1e0d08_3935);
nor \g449965/U$1 ( \17364 , \17362 , \17363 );
and \g452061/U$2 ( \17365 , \16361 , RIe1bf108_3551);
and \g452061/U$3 ( \17366 , RIe1c1e08_3583, \16364 );
nor \g452061/U$1 ( \17367 , \17365 , \17366 );
and \g452057/U$2 ( \17368 , \16368 , RIe1ca508_3679);
and \g452057/U$3 ( \17369 , RIe1cd208_3711, \16371 );
nor \g452057/U$1 ( \17370 , \17368 , \17369 );
nand \g447700/U$1 ( \17371 , \17356 , \17364 , \17367 , \17370 );
nor \g446052/U$1 ( \17372 , \17351 , \17352 , \17371 );
and \g452054/U$2 ( \17373 , \16377 , RIe1e3a08_3967);
and \g452054/U$3 ( \17374 , RIe1db308_3871, \16380 );
nor \g452054/U$1 ( \17375 , \17373 , \17374 );
and \g452157/U$2 ( \17376 , \16334 , RIe1d8608_3839);
and \g452157/U$3 ( \17377 , RIe1ec108_4063, \16326 );
nor \g452157/U$1 ( \17378 , \17376 , \17377 );
and \g445189/U$2 ( \17379 , \17372 , \17375 , \17378 );
nor \g445189/U$1 ( \17380 , \17379 , \16555 );
and \g446056/U$2 ( \17381 , RIe1ff500_4282, \16427 );
and \g446056/U$3 ( \17382 , RIe1f1400_4122, \16368 );
and \g448952/U$2 ( \17383 , RIe179748_2759, \16485 );
and \g448952/U$3 ( \17384 , \16356 , RIe18d248_2983);
and \g448952/U$4 ( \17385 , RIe1bc408_3519, \16337 );
nor \g448952/U$1 ( \17386 , \17383 , \17384 , \17385 );
and \g454998/U$2 ( \17387 , \16317 , RIe1a6748_3271);
and \g454998/U$3 ( \17388 , RIe1a9448_3303, \16325 );
nor \g454998/U$1 ( \17389 , \17387 , \17388 );
not \g449969/U$3 ( \17390 , \17389 );
not \g449969/U$4 ( \17391 , \16311 );
and \g449969/U$2 ( \17392 , \17390 , \17391 );
and \g449969/U$5 ( \17393 , \16341 , RIe1d5908_3807);
nor \g449969/U$1 ( \17394 , \17392 , \17393 );
and \g452076/U$2 ( \17395 , \16377 , RIe1a0d48_3207);
and \g452076/U$3 ( \17396 , RIe1a3a48_3239, \16313 );
nor \g452076/U$1 ( \17397 , \17395 , \17396 );
and \g452079/U$2 ( \17398 , \16334 , RIe21bca0_4606);
and \g452079/U$3 ( \17399 , RIe2270a0_4734, \16380 );
nor \g452079/U$1 ( \17400 , \17398 , \17399 );
nand \g447328/U$1 ( \17401 , \17386 , \17394 , \17397 , \17400 );
nor \g446056/U$1 ( \17402 , \17381 , \17382 , \17401 );
and \g452072/U$2 ( \17403 , \16361 , RIe1718b8_2669);
and \g452072/U$3 ( \17404 , RIe2054a0_4350, \16432 );
nor \g452072/U$1 ( \17405 , \17403 , \17404 );
and \g452071/U$2 ( \17406 , \16364 , RIe1af280_3370);
and \g452071/U$3 ( \17407 , RIe1f88b8_4205, \16371 );
nor \g452071/U$1 ( \17408 , \17406 , \17407 );
and \g445191/U$2 ( \17409 , \17402 , \17405 , \17408 );
nor \g445191/U$1 ( \17410 , \17409 , \16586 );
or \g444225/U$1 ( \17411 , \17350 , \17380 , \17410 );
_DC \g34f1/U$1 ( \17412 , \17411 , \16652 );
and \g450835/U$2 ( \17413 , \16313 , RIfc7e050_6456);
and \g450835/U$3 ( \17414 , RIfc5dda0_6090, \16321 );
nor \g450835/U$1 ( \17415 , \17413 , \17414 );
and \g445762/U$2 ( \17416 , RIfc5e070_6092, \16328 );
and \g445762/U$3 ( \17417 , RIe1f5d20_4174, \16334 );
and \g448574/U$2 ( \17418 , RIfc8cdf8_6625, \16427 );
and \g448574/U$3 ( \17419 , \16432 , RIfca4138_6889);
and \g448574/U$4 ( \17420 , RIfcd9568_7495, \16485 );
nor \g448574/U$1 ( \17421 , \17418 , \17419 , \17420 );
and \g454495/U$2 ( \17422 , \16317 , RIfcbc3f0_7164);
and \g454495/U$3 ( \17423 , RIfc99440_6766, \16325 );
nor \g454495/U$1 ( \17424 , \17422 , \17423 );
not \g454494/U$1 ( \17425 , \17424 );
and \g449601/U$2 ( \17426 , \17425 , \16336 );
and \g449601/U$3 ( \17427 , RIfc5d968_6087, \16356 );
nor \g449601/U$1 ( \17428 , \17426 , \17427 );
and \g450845/U$2 ( \17429 , \16361 , RIe1ee700_4090);
and \g450845/U$3 ( \17430 , RIfc5a128_6047, \16364 );
nor \g450845/U$1 ( \17431 , \17429 , \17430 );
and \g450844/U$2 ( \17432 , \16368 , RIe1f39f8_4149);
and \g450844/U$3 ( \17433 , RIfcc7c28_7295, \16371 );
nor \g450844/U$1 ( \17434 , \17432 , \17433 );
nand \g448013/U$1 ( \17435 , \17421 , \17428 , \17431 , \17434 );
nor \g445762/U$1 ( \17436 , \17416 , \17417 , \17435 );
and \g450839/U$2 ( \17437 , \16377 , RIe1fa7a8_4227);
and \g450839/U$3 ( \17438 , RIfc8d668_6631, \16380 );
nor \g450839/U$1 ( \17439 , \17437 , \17438 );
nand \g445519/U$1 ( \17440 , \17415 , \17436 , \17439 );
and \g444831/U$2 ( \17441 , \17440 , \16481 );
and \g448569/U$2 ( \17442 , RIf14bb98_5321, \16321 );
and \g448569/U$3 ( \17443 , \16328 , RIf14cde0_5334);
and \g448569/U$4 ( \17444 , RIf1468a0_5262, \16398 );
nor \g448569/U$1 ( \17445 , \17442 , \17443 , \17444 );
and \g455057/U$2 ( \17446 , \16317 , RIfc9e738_6825);
and \g455057/U$3 ( \17447 , RIfc4c460_5890, \16325 );
nor \g455057/U$1 ( \17448 , \17446 , \17447 );
not \g449595/U$3 ( \17449 , \17448 );
not \g449595/U$4 ( \17450 , \16330 );
and \g449595/U$2 ( \17451 , \17449 , \17450 );
and \g449595/U$5 ( \17452 , \16339 , RIf1473e0_5270);
nor \g449595/U$1 ( \17453 , \17451 , \17452 );
and \g452687/U$2 ( \17454 , \16377 , RIe1b7980_3466);
and \g452687/U$3 ( \17455 , RIe1b99d8_3489, \16313 );
nor \g452687/U$1 ( \17456 , \17454 , \17455 );
and \g450829/U$2 ( \17457 , \16334 , RIfec54d8_8365);
and \g450829/U$3 ( \17458 , RIe1b5658_3441, \16380 );
nor \g450829/U$1 ( \17459 , \17457 , \17458 );
nand \g447254/U$1 ( \17460 , \17445 , \17453 , \17456 , \17459 );
and \g444831/U$3 ( \17461 , \16477 , \17460 );
nor \g444831/U$1 ( \17462 , \17441 , \17461 );
nor \g448282/U$1 ( \17463 , \16909 , \16418 );
and \g446559/U$2 ( \17464 , \17463 , RIe1ab338_3325);
nor \g448281/U$1 ( \17465 , \16909 , \16428 );
and \g446559/U$3 ( \17466 , RIf147f20_5278, \17465 );
nor \g446559/U$1 ( \17467 , \17464 , \17466 );
nor \g448280/U$1 ( \17468 , \16909 , \16421 );
and \g446558/U$2 ( \17469 , \17468 , RIe1acb20_3342);
nor \g448278/U$1 ( \17470 , \16909 , \16433 );
and \g446558/U$3 ( \17471 , RIf149168_5291, \17470 );
nor \g446558/U$1 ( \17472 , \17469 , \17471 );
nor \g448284/U$1 ( \17473 , \16909 , \16437 );
and \g446561/U$2 ( \17474 , \17473 , RIe1b1170_3392);
nor \g448283/U$1 ( \17475 , \16909 , \16440 );
and \g446561/U$3 ( \17476 , RIe1b2ac0_3410, \17475 );
nor \g446561/U$1 ( \17477 , \17474 , \17476 );
nand \g444556/U$1 ( \17478 , \17462 , \17467 , \17472 , \17477 );
and \g450872/U$2 ( \17479 , \16364 , RIe1c1ca0_3582);
and \g450872/U$3 ( \17480 , RIe1cd0a0_3710, \16371 );
nor \g450872/U$1 ( \17481 , \17479 , \17480 );
and \g445770/U$2 ( \17482 , RIe1cfda0_3742, \16427 );
and \g445770/U$3 ( \17483 , RIe1ca3a0_3678, \16368 );
and \g448585/U$2 ( \17484 , RIe1e92a0_4030, \16321 );
and \g448585/U$3 ( \17485 , \16328 , RIe1ebfa0_4062);
and \g448585/U$4 ( \17486 , RIe1c49a0_3614, \16398 );
nor \g448585/U$1 ( \17487 , \17484 , \17485 , \17486 );
and \g454290/U$2 ( \17488 , \16317 , RIe1ddea0_3902);
and \g454290/U$3 ( \17489 , RIe1e0ba0_3934, \16325 );
nor \g454290/U$1 ( \17490 , \17488 , \17489 );
not \g449611/U$3 ( \17491 , \17490 );
not \g449611/U$4 ( \17492 , \16330 );
and \g449611/U$2 ( \17493 , \17491 , \17492 );
and \g449611/U$5 ( \17494 , \16341 , RIe1c76a0_3646);
nor \g449611/U$1 ( \17495 , \17493 , \17494 );
and \g450876/U$2 ( \17496 , \16377 , RIe1e38a0_3966);
and \g450876/U$3 ( \17497 , RIe1e65a0_3998, \16313 );
nor \g450876/U$1 ( \17498 , \17496 , \17497 );
and \g450903/U$2 ( \17499 , \16334 , RIe1d84a0_3838);
and \g450903/U$3 ( \17500 , RIe1db1a0_3870, \16380 );
nor \g450903/U$1 ( \17501 , \17499 , \17500 );
nand \g447257/U$1 ( \17502 , \17487 , \17495 , \17498 , \17501 );
nor \g445770/U$1 ( \17503 , \17482 , \17483 , \17502 );
and \g450875/U$2 ( \17504 , \16361 , RIe1befa0_3550);
and \g450875/U$3 ( \17505 , RIe1d2aa0_3774, \16448 );
nor \g450875/U$1 ( \17506 , \17504 , \17505 );
nand \g445522/U$1 ( \17507 , \17481 , \17503 , \17506 );
and \g444755/U$2 ( \17508 , \17507 , \16750 );
and \g448579/U$2 ( \17509 , RIe1795e0_2758, \16485 );
and \g448579/U$3 ( \17510 , \16356 , RIe18d0e0_2982);
and \g448579/U$4 ( \17511 , RIe1bc2a0_3518, \16398 );
nor \g448579/U$1 ( \17512 , \17509 , \17510 , \17511 );
and \g454473/U$2 ( \17513 , \16317 , RIe1a65e0_3270);
and \g454473/U$3 ( \17514 , RIe1a92e0_3302, \16325 );
nor \g454473/U$1 ( \17515 , \17513 , \17514 );
not \g449605/U$3 ( \17516 , \17515 );
not \g449605/U$4 ( \17517 , \16311 );
and \g449605/U$2 ( \17518 , \17516 , \17517 );
and \g449605/U$5 ( \17519 , \16339 , RIe1d57a0_3806);
nor \g449605/U$1 ( \17520 , \17518 , \17519 );
and \g450861/U$2 ( \17521 , \16377 , RIe1a0be0_3206);
and \g450861/U$3 ( \17522 , RIe1a38e0_3238, \16313 );
nor \g450861/U$1 ( \17523 , \17521 , \17522 );
and \g450865/U$2 ( \17524 , \16334 , RIe21bb38_4605);
and \g450865/U$3 ( \17525 , RIe226f38_4733, \16380 );
nor \g450865/U$1 ( \17526 , \17524 , \17525 );
nand \g447256/U$1 ( \17527 , \17512 , \17520 , \17523 , \17526 );
and \g444755/U$3 ( \17528 , \16752 , \17527 );
nor \g444755/U$1 ( \17529 , \17508 , \17528 );
and \g446567/U$2 ( \17530 , \16774 , RIe171750_2668);
and \g446567/U$3 ( \17531 , RIe1af118_3369, \16776 );
nor \g446567/U$1 ( \17532 , \17530 , \17531 );
and \g446566/U$2 ( \17533 , \16779 , RIe1f1298_4121);
and \g446566/U$3 ( \17534 , RIe1f8750_4204, \16781 );
nor \g446566/U$1 ( \17535 , \17533 , \17534 );
and \g446565/U$2 ( \17536 , \16784 , RIe1ff398_4281);
and \g446565/U$3 ( \17537 , RIe205338_4349, \16786 );
nor \g446565/U$1 ( \17538 , \17536 , \17537 );
nand \g444455/U$1 ( \17539 , \17529 , \17532 , \17535 , \17538 );
and \g445752/U$2 ( \17540 , RIe19b1e0_3142, \16321 );
and \g445752/U$3 ( \17541 , RIfc67580_6198, \16313 );
and \g448560/U$2 ( \17542 , RIe1876e0_2918, \16427 );
and \g448560/U$3 ( \17543 , \16432 , RIe18a3e0_2950);
and \g448560/U$4 ( \17544 , RIe1957e0_3078, \16485 );
nor \g448560/U$1 ( \17545 , \17542 , \17543 , \17544 );
and \g454443/U$2 ( \17546 , \16317 , RIe181ce0_2854);
and \g454443/U$3 ( \17547 , RIfcaa7e0_6962, \16325 );
nor \g454443/U$1 ( \17548 , \17546 , \17547 );
not \g454442/U$1 ( \17549 , \17548 );
and \g449586/U$2 ( \17550 , \17549 , \16336 );
and \g449586/U$3 ( \17551 , RIfccb030_7332, \16356 );
nor \g449586/U$1 ( \17552 , \17550 , \17551 );
and \g450796/U$2 ( \17553 , \16361 , RIe17c2e0_2790);
and \g450796/U$3 ( \17554 , RIe17efe0_2822, \16364 );
nor \g450796/U$1 ( \17555 , \17553 , \17554 );
and \g450794/U$2 ( \17556 , \16368 , RIe1849e0_2886);
and \g450794/U$3 ( \17557 , RIfc6a550_6232, \16371 );
nor \g450794/U$1 ( \17558 , \17556 , \17557 );
nand \g448012/U$1 ( \17559 , \17545 , \17552 , \17555 , \17558 );
nor \g445752/U$1 ( \17560 , \17540 , \17541 , \17559 );
and \g450787/U$2 ( \17561 , \16377 , RIe1984e0_3110);
and \g450787/U$3 ( \17562 , RIe192ae0_3046, \16380 );
nor \g450787/U$1 ( \17563 , \17561 , \17562 );
and \g450786/U$2 ( \17564 , \16334 , RIe18fde0_3014);
and \g450786/U$3 ( \17565 , RIe19dee0_3174, \16328 );
nor \g450786/U$1 ( \17566 , \17564 , \17565 );
and \g444966/U$2 ( \17567 , \17560 , \17563 , \17566 );
nor \g444966/U$1 ( \17568 , \17567 , \16618 );
and \g445756/U$2 ( \17569 , RIfca9430_6948, \16427 );
and \g445756/U$3 ( \17570 , RIe174018_2697, \16368 );
and \g448565/U$2 ( \17571 , RIfc607d0_6120, \16485 );
and \g448565/U$3 ( \17572 , \16354 , RIfcca928_7327);
and \g448565/U$4 ( \17573 , RIfc650f0_6172, \16398 );
nor \g448565/U$1 ( \17574 , \17571 , \17572 , \17573 );
and \g454258/U$2 ( \17575 , \16317 , RIfc65690_6176);
and \g454258/U$3 ( \17576 , RIfc65d98_6181, \16325 );
nor \g454258/U$1 ( \17577 , \17575 , \17576 );
not \g449591/U$3 ( \17578 , \17577 );
not \g449591/U$4 ( \17579 , \16311 );
and \g449591/U$2 ( \17580 , \17578 , \17579 );
and \g449591/U$5 ( \17581 , \16339 , RIfcecf00_7718);
nor \g449591/U$1 ( \17582 , \17580 , \17581 );
and \g450812/U$2 ( \17583 , \16377 , RIfea0638_8169);
and \g450812/U$3 ( \17584 , RIe1772b8_2733, \16313 );
nor \g450812/U$1 ( \17585 , \17583 , \17584 );
and \g450813/U$2 ( \17586 , \16334 , RIee3d798_5158);
and \g450813/U$3 ( \17587 , RIfc65258_6173, \16380 );
nor \g450813/U$1 ( \17588 , \17586 , \17587 );
nand \g447253/U$1 ( \17589 , \17574 , \17582 , \17585 , \17588 );
nor \g445756/U$1 ( \17590 , \17569 , \17570 , \17589 );
and \g450806/U$2 ( \17591 , \16361 , RIfc43a90_5792);
and \g450806/U$3 ( \17592 , RIee3c3e8_5144, \16448 );
nor \g450806/U$1 ( \17593 , \17591 , \17592 );
and \g450805/U$2 ( \17594 , \16364 , RIf16e5a8_5715);
and \g450805/U$3 ( \17595 , RIee39f58_5118, \16371 );
nor \g450805/U$1 ( \17596 , \17594 , \17595 );
and \g444967/U$2 ( \17597 , \17590 , \17593 , \17596 );
nor \g444967/U$1 ( \17598 , \17597 , \16649 );
or \g444383/U$1 ( \17599 , \17478 , \17539 , \17568 , \17598 );
and \g445745/U$2 ( \17600 , RIfc65528_6175, \16328 );
and \g445745/U$3 ( \17601 , RIe221538_4669, \16377 );
and \g448549/U$2 ( \17602 , RIe20da38_4445, \16398 );
and \g448549/U$3 ( \17603 , \16339 , RIfc60c08_6123);
and \g448549/U$4 ( \17604 , RIe21e838_4637, \16485 );
nor \g448549/U$1 ( \17605 , \17602 , \17603 , \17604 );
and \g454719/U$2 ( \17606 , \16317 , RIe213438_4509);
and \g454719/U$3 ( \17607 , RIfc3fda0_5752, \16325 );
nor \g454719/U$1 ( \17608 , \17606 , \17607 );
not \g449573/U$3 ( \17609 , \17608 );
not \g449573/U$4 ( \17610 , \16351 );
and \g449573/U$2 ( \17611 , \17609 , \17610 );
and \g449573/U$5 ( \17612 , \16356 , RIfc6b4c8_6243);
nor \g449573/U$1 ( \17613 , \17611 , \17612 );
and \g450762/U$2 ( \17614 , \16361 , RIe208038_4381);
and \g450762/U$3 ( \17615 , RIe20ad38_4413, \16364 );
nor \g450762/U$1 ( \17616 , \17614 , \17615 );
and \g450761/U$2 ( \17617 , \16368 , RIe210738_4477);
and \g450761/U$3 ( \17618 , RIfc61310_6128, \16371 );
nor \g450761/U$1 ( \17619 , \17617 , \17618 );
nand \g447483/U$1 ( \17620 , \17605 , \17613 , \17616 , \17619 );
nor \g445745/U$1 ( \17621 , \17600 , \17601 , \17620 );
and \g450754/U$2 ( \17622 , \16334 , RIe216138_4541);
and \g450754/U$3 ( \17623 , RIfca9f70_6956, \16313 );
nor \g450754/U$1 ( \17624 , \17622 , \17623 );
and \g450753/U$2 ( \17625 , \16380 , RIe218e38_4573);
and \g450753/U$3 ( \17626 , RIe224238_4701, \16321 );
nor \g450753/U$1 ( \17627 , \17625 , \17626 );
and \g444957/U$2 ( \17628 , \17621 , \17624 , \17627 );
nor \g444957/U$1 ( \17629 , \17628 , \16389 );
and \g445749/U$2 ( \17630 , RIfc73358_6333, \16427 );
and \g445749/U$3 ( \17631 , RIe1fbe28_4243, \16368 );
and \g448555/U$2 ( \17632 , RIfccbcd8_7341, \16319 );
and \g448555/U$3 ( \17633 , \16326 , RIfc66ba8_6191);
and \g448555/U$4 ( \17634 , RIfc44468_5799, \16398 );
nor \g448555/U$1 ( \17635 , \17632 , \17633 , \17634 );
and \g454637/U$2 ( \17636 , \16317 , RIfccbe40_7342);
and \g454637/U$3 ( \17637 , RIfcadbe8_6999, \16325 );
nor \g454637/U$1 ( \17638 , \17636 , \17637 );
not \g449582/U$3 ( \17639 , \17638 );
not \g449582/U$4 ( \17640 , \16330 );
and \g449582/U$2 ( \17641 , \17639 , \17640 );
and \g449582/U$5 ( \17642 , \16339 , RIfcc2660_7234);
nor \g449582/U$1 ( \17643 , \17641 , \17642 );
and \g450776/U$2 ( \17644 , \16377 , RIe200fb8_4301);
and \g450776/U$3 ( \17645 , RIe202bd8_4321, \16313 );
nor \g450776/U$1 ( \17646 , \17644 , \17645 );
and \g450777/U$2 ( \17647 , \16334 , RIfc6a3e8_6231);
and \g450777/U$3 ( \17648 , RIfca7540_6926, \16380 );
nor \g450777/U$1 ( \17649 , \17647 , \17648 );
nand \g447251/U$1 ( \17650 , \17635 , \17643 , \17646 , \17649 );
nor \g445749/U$1 ( \17651 , \17630 , \17631 , \17650 );
and \g450772/U$2 ( \17652 , \16361 , RIfca7270_6924);
and \g450772/U$3 ( \17653 , RIfca6898_6917, \16448 );
nor \g450772/U$1 ( \17654 , \17652 , \17653 );
and \g451988/U$2 ( \17655 , \16364 , RIf15a940_5490);
and \g451988/U$3 ( \17656 , RIe1fd070_4256, \16371 );
nor \g451988/U$1 ( \17657 , \17655 , \17656 );
and \g444960/U$2 ( \17658 , \17651 , \17654 , \17657 );
nor \g444960/U$1 ( \17659 , \17658 , \16393 );
or \g444205/U$1 ( \17660 , \17599 , \17629 , \17659 );
_DC \g3576/U$1 ( \17661 , \17660 , \16652 );
and \g446605/U$2 ( \17662 , \17284 , RIe1ee598_4089);
and \g446605/U$3 ( \17663 , RIfc73e98_6341, \17286 );
nor \g446605/U$1 ( \17664 , \17662 , \17663 );
and \g445814/U$2 ( \17665 , RIf14fc48_5367, \16341 );
and \g445814/U$3 ( \17666 , RIfc72c50_6328, \16398 );
and \g448640/U$2 ( \17667 , RIfc6ba68_6247, \16321 );
and \g448640/U$3 ( \17668 , \16485 , RIfc53918_5973);
and \g448640/U$4 ( \17669 , RIfcce000_7366, \16356 );
nor \g448640/U$1 ( \17670 , \17667 , \17668 , \17669 );
and \g453679/U$2 ( \17671 , \16368 , RIe1f3890_4148);
and \g453679/U$3 ( \17672 , RIfc72db8_6329, \16371 );
nor \g453679/U$1 ( \17673 , \17671 , \17672 );
and \g454363/U$2 ( \17674 , \16317 , RIf151e08_5391);
and \g454363/U$3 ( \17675 , RIf1535f0_5408, \16325 );
nor \g454363/U$1 ( \17676 , \17674 , \17675 );
not \g449665/U$3 ( \17677 , \17676 );
not \g449665/U$4 ( \17678 , \16351 );
and \g449665/U$2 ( \17679 , \17677 , \17678 );
and \g449665/U$5 ( \17680 , \16328 , RIfcce5a0_7370);
nor \g449665/U$1 ( \17681 , \17679 , \17680 );
and \g451080/U$2 ( \17682 , \16334 , RIe1f5bb8_4173);
and \g451080/U$3 ( \17683 , RIfcce708_7371, \16380 );
nor \g451080/U$1 ( \17684 , \17682 , \17683 );
nand \g447532/U$1 ( \17685 , \17670 , \17673 , \17681 , \17684 );
nor \g445814/U$1 ( \17686 , \17665 , \17666 , \17685 );
not \g444812/U$3 ( \17687 , \17686 );
not \g444812/U$4 ( \17688 , \16480 );
and \g444812/U$2 ( \17689 , \17687 , \17688 );
and \g445818/U$2 ( \17690 , RIe1e0a38_3933, \16356 );
and \g445818/U$3 ( \17691 , RIe1ca238_3677, \16368 );
and \g448644/U$2 ( \17692 , RIe1cfc38_3741, \16427 );
and \g448644/U$3 ( \17693 , \16398 , RIe1c4838_3613);
and \g448644/U$4 ( \17694 , RIe1c7538_3645, \16341 );
nor \g448644/U$1 ( \17695 , \17692 , \17693 , \17694 );
and \g453450/U$2 ( \17696 , \16361 , RIe1bee38_3549);
and \g453450/U$3 ( \17697 , RIe1c1b38_3581, \16364 );
nor \g453450/U$1 ( \17698 , \17696 , \17697 );
and \g451096/U$2 ( \17699 , \16377 , RIe1e3738_3965);
and \g451096/U$3 ( \17700 , RIe1e6438_3997, \16313 );
nor \g451096/U$1 ( \17701 , \17699 , \17700 );
and \g454370/U$2 ( \17702 , \16317 , RIe1e9138_4029);
and \g454370/U$3 ( \17703 , RIe1ebe38_4061, \16325 );
nor \g454370/U$1 ( \17704 , \17702 , \17703 );
not \g449670/U$3 ( \17705 , \17704 );
not \g449670/U$4 ( \17706 , \16311 );
and \g449670/U$2 ( \17707 , \17705 , \17706 );
and \g449670/U$5 ( \17708 , \16448 , RIe1d2938_3773);
nor \g449670/U$1 ( \17709 , \17707 , \17708 );
nand \g447535/U$1 ( \17710 , \17695 , \17698 , \17701 , \17709 );
nor \g445818/U$1 ( \17711 , \17690 , \17691 , \17710 );
and \g451091/U$2 ( \17712 , \16334 , RIe1d8338_3837);
and \g451091/U$3 ( \17713 , RIe1ccf38_3709, \16371 );
nor \g451091/U$1 ( \17714 , \17712 , \17713 );
and \g451089/U$2 ( \17715 , \16380 , RIe1db038_3869);
and \g451089/U$3 ( \17716 , RIe1ddd38_3901, \16485 );
nor \g451089/U$1 ( \17717 , \17715 , \17716 );
and \g445014/U$2 ( \17718 , \17711 , \17714 , \17717 );
nor \g445014/U$1 ( \17719 , \17718 , \16555 );
nor \g444812/U$1 ( \17720 , \17689 , \17719 );
and \g446606/U$2 ( \17721 , \16518 , RIe1fa640_4226);
and \g446606/U$3 ( \17722 , RIfc6f410_6288, \16521 );
nor \g446606/U$1 ( \17723 , \17721 , \17722 );
nand \g444419/U$1 ( \17724 , \17664 , \17720 , \17723 );
and \g451120/U$2 ( \17725 , \16364 , RIe1ac9b8_3341);
and \g451120/U$3 ( \17726 , RIfc82ad8_6509, \16337 );
nor \g451120/U$1 ( \17727 , \17725 , \17726 );
and \g445825/U$2 ( \17728 , RIfcc5900_7270, \16341 );
and \g445825/U$3 ( \17729 , RIe1b7818_3465, \16377 );
and \g448653/U$2 ( \17730 , RIfcb84a8_7119, \16321 );
and \g448653/U$3 ( \17731 , \16485 , RIfc9e198_6821);
and \g448653/U$4 ( \17732 , RIfc85940_6542, \16354 );
nor \g448653/U$1 ( \17733 , \17730 , \17731 , \17732 );
and \g451127/U$2 ( \17734 , \16368 , RIe1b1008_3391);
and \g451127/U$3 ( \17735 , RIfe884e8_7895, \16371 );
nor \g451127/U$1 ( \17736 , \17734 , \17735 );
and \g455085/U$2 ( \17737 , \16317 , RIfc838e8_6519);
and \g455085/U$3 ( \17738 , RIfc518c0_5950, \16325 );
nor \g455085/U$1 ( \17739 , \17737 , \17738 );
not \g449678/U$3 ( \17740 , \17739 );
not \g449678/U$4 ( \17741 , \16351 );
and \g449678/U$2 ( \17742 , \17740 , \17741 );
and \g449678/U$5 ( \17743 , \16326 , RIfcb8a48_7123);
nor \g449678/U$1 ( \17744 , \17742 , \17743 );
and \g451125/U$2 ( \17745 , \16334 , RIe1b42a8_3427);
and \g451125/U$3 ( \17746 , RIfeac140_8274, \16380 );
nor \g451125/U$1 ( \17747 , \17745 , \17746 );
nand \g447543/U$1 ( \17748 , \17733 , \17736 , \17744 , \17747 );
nor \g445825/U$1 ( \17749 , \17728 , \17729 , \17748 );
and \g451117/U$2 ( \17750 , \16361 , RIfe88650_7896);
and \g451117/U$3 ( \17751 , RIe1b9870_3488, \16313 );
nor \g451117/U$1 ( \17752 , \17750 , \17751 );
nand \g445534/U$1 ( \17753 , \17727 , \17749 , \17752 );
and \g444907/U$2 ( \17754 , \17753 , \16477 );
and \g448648/U$2 ( \17755 , RIe1ff230_4280, \16427 );
and \g448648/U$3 ( \17756 , \16432 , RIe2051d0_4348);
and \g448648/U$4 ( \17757 , RIe1a6478_3269, \16319 );
nor \g448648/U$1 ( \17758 , \17755 , \17756 , \17757 );
and \g451108/U$2 ( \17759 , \16368 , RIe1f1130_4120);
and \g451108/U$3 ( \17760 , RIe1f85e8_4203, \16371 );
nor \g451108/U$1 ( \17761 , \17759 , \17760 );
and \g455253/U$2 ( \17762 , \16317 , RIe179478_2757);
and \g455253/U$3 ( \17763 , RIe18cf78_2981, \16325 );
nor \g455253/U$1 ( \17764 , \17762 , \17763 );
not \g449673/U$3 ( \17765 , \17764 );
not \g449673/U$4 ( \17766 , \16330 );
and \g449673/U$2 ( \17767 , \17765 , \17766 );
and \g449673/U$5 ( \17768 , \16328 , RIe1a9178_3301);
nor \g449673/U$1 ( \17769 , \17767 , \17768 );
and \g451107/U$2 ( \17770 , \16334 , RIe21b9d0_4604);
and \g451107/U$3 ( \17771 , RIe226dd0_4732, \16380 );
nor \g451107/U$1 ( \17772 , \17770 , \17771 );
nand \g447539/U$1 ( \17773 , \17758 , \17761 , \17769 , \17772 );
and \g444907/U$3 ( \17774 , \16752 , \17773 );
nor \g444907/U$1 ( \17775 , \17754 , \17774 );
and \g446615/U$2 ( \17776 , \17027 , RIe1bc138_3517);
and \g446615/U$3 ( \17777 , RIe1d5638_3805, \17034 );
nor \g446615/U$1 ( \17778 , \17776 , \17777 );
nor \g448373/U$1 ( \17779 , \16586 , \16517 );
and \g446614/U$2 ( \17780 , \17779 , RIe1a0a78_3205);
nor \g448343/U$1 ( \17781 , \16586 , \16520 );
and \g446614/U$3 ( \17782 , RIe1a3778_3237, \17781 );
nor \g446614/U$1 ( \17783 , \17780 , \17782 );
and \g446616/U$2 ( \17784 , \16774 , RIe1715e8_2667);
and \g446616/U$3 ( \17785 , RIe1aefb0_3368, \16776 );
nor \g446616/U$1 ( \17786 , \17784 , \17785 );
nand \g444566/U$1 ( \17787 , \17775 , \17778 , \17783 , \17786 );
and \g445807/U$2 ( \17788 , RIfc87c68_6567, \16356 );
and \g445807/U$3 ( \17789 , RIe173eb0_2696, \16368 );
and \g448631/U$2 ( \17790 , RIfc9bd08_6795, \16321 );
and \g448631/U$3 ( \17791 , \16328 , RIfc9be70_6796);
and \g448631/U$4 ( \17792 , RIfc876c8_6563, \16427 );
nor \g448631/U$1 ( \17793 , \17790 , \17791 , \17792 );
and \g451053/U$2 ( \17794 , \16361 , RIfc9d388_6811);
and \g451053/U$3 ( \17795 , RIfc4e350_5912, \16364 );
nor \g451053/U$1 ( \17796 , \17794 , \17795 );
and \g451051/U$2 ( \17797 , \16377 , RIe176070_2720);
and \g451051/U$3 ( \17798 , RIfc4ccd0_5896, \16313 );
nor \g451051/U$1 ( \17799 , \17797 , \17798 );
and \g454349/U$2 ( \17800 , \16317 , RIfc4e080_5910);
and \g454349/U$3 ( \17801 , RIfcb9420_7130, \16325 );
nor \g454349/U$1 ( \17802 , \17800 , \17801 );
not \g454348/U$1 ( \17803 , \17802 );
and \g449658/U$2 ( \17804 , \17803 , \16336 );
and \g449658/U$3 ( \17805 , RIfc4f598_5925, \16448 );
nor \g449658/U$1 ( \17806 , \17804 , \17805 );
nand \g448019/U$1 ( \17807 , \17793 , \17796 , \17799 , \17806 );
nor \g445807/U$1 ( \17808 , \17788 , \17789 , \17807 );
and \g451045/U$2 ( \17809 , \16334 , RIfc4fca0_5930);
and \g451045/U$3 ( \17810 , RIfc4dae0_5906, \16371 );
nor \g451045/U$1 ( \17811 , \17809 , \17810 );
and \g451044/U$2 ( \17812 , \16380 , RIfcc4c58_7261);
and \g451044/U$3 ( \17813 , RIfc87b00_6566, \16485 );
nor \g451044/U$1 ( \17814 , \17812 , \17813 );
and \g445006/U$2 ( \17815 , \17808 , \17811 , \17814 );
nor \g445006/U$1 ( \17816 , \17815 , \16649 );
and \g445810/U$2 ( \17817 , RIfc9ba38_6793, \16356 );
and \g445810/U$3 ( \17818 , RIe2105d0_4476, \16368 );
and \g448635/U$2 ( \17819 , RIe2240d0_4700, \16321 );
and \g448635/U$3 ( \17820 , \16328 , RIfc40a48_5761);
and \g448635/U$4 ( \17821 , RIe2132d0_4508, \16427 );
nor \g448635/U$1 ( \17822 , \17819 , \17820 , \17821 );
and \g451070/U$2 ( \17823 , \16361 , RIe207ed0_4380);
and \g451070/U$3 ( \17824 , RIe20abd0_4412, \16364 );
nor \g451070/U$1 ( \17825 , \17823 , \17824 );
and \g451068/U$2 ( \17826 , \16377 , RIe2213d0_4668);
and \g451068/U$3 ( \17827 , RIfc85508_6539, \16313 );
nor \g451068/U$1 ( \17828 , \17826 , \17827 );
and \g454451/U$2 ( \17829 , \16317 , RIe20d8d0_4444);
and \g454451/U$3 ( \17830 , RIfc97988_6747, \16325 );
nor \g454451/U$1 ( \17831 , \17829 , \17830 );
not \g454450/U$1 ( \17832 , \17831 );
and \g449662/U$2 ( \17833 , \17832 , \16336 );
and \g449662/U$3 ( \17834 , RIfc52c70_5964, \16432 );
nor \g449662/U$1 ( \17835 , \17833 , \17834 );
nand \g448021/U$1 ( \17836 , \17822 , \17825 , \17828 , \17835 );
nor \g445810/U$1 ( \17837 , \17817 , \17818 , \17836 );
and \g451064/U$2 ( \17838 , \16334 , RIe215fd0_4540);
and \g451064/U$3 ( \17839 , RIfca3760_6882, \16371 );
nor \g451064/U$1 ( \17840 , \17838 , \17839 );
and \g451063/U$2 ( \17841 , \16380 , RIe218cd0_4572);
and \g451063/U$3 ( \17842 , RIe21e6d0_4636, \16485 );
nor \g451063/U$1 ( \17843 , \17841 , \17842 );
and \g445009/U$2 ( \17844 , \17837 , \17840 , \17843 );
nor \g445009/U$1 ( \17845 , \17844 , \16389 );
or \g444297/U$1 ( \17846 , \17724 , \17787 , \17816 , \17845 );
and \g445801/U$2 ( \17847 , RIf142d90_5220, \16339 );
and \g445801/U$3 ( \17848 , RIe198378_3109, \16377 );
and \g448622/U$2 ( \17849 , RIe19b078_3141, \16321 );
and \g448622/U$3 ( \17850 , \16485 , RIe195678_3077);
and \g448622/U$4 ( \17851 , RIfca35f8_6881, \16356 );
nor \g448622/U$1 ( \17852 , \17849 , \17850 , \17851 );
and \g451025/U$2 ( \17853 , \16368 , RIe184878_2885);
and \g451025/U$3 ( \17854 , RIfcba230_7140, \16371 );
nor \g451025/U$1 ( \17855 , \17853 , \17854 );
and \g454338/U$2 ( \17856 , \16317 , RIe187578_2917);
and \g454338/U$3 ( \17857 , RIe18a278_2949, \16325 );
nor \g454338/U$1 ( \17858 , \17856 , \17857 );
not \g449649/U$3 ( \17859 , \17858 );
not \g449649/U$4 ( \17860 , \16351 );
and \g449649/U$2 ( \17861 , \17859 , \17860 );
and \g449649/U$5 ( \17862 , \16328 , RIe19dd78_3173);
nor \g449649/U$1 ( \17863 , \17861 , \17862 );
and \g451022/U$2 ( \17864 , \16334 , RIe18fc78_3013);
and \g451022/U$3 ( \17865 , RIe192978_3045, \16380 );
nor \g451022/U$1 ( \17866 , \17864 , \17865 );
nand \g447524/U$1 ( \17867 , \17852 , \17855 , \17863 , \17866 );
nor \g445801/U$1 ( \17868 , \17847 , \17848 , \17867 );
and \g451013/U$2 ( \17869 , \16361 , RIe17c178_2789);
and \g451013/U$3 ( \17870 , RIfca1438_6857, \16313 );
nor \g451013/U$1 ( \17871 , \17869 , \17870 );
and \g451016/U$2 ( \17872 , \16364 , RIe17ee78_2821);
and \g451016/U$3 ( \17873 , RIe181b78_2853, \16398 );
nor \g451016/U$1 ( \17874 , \17872 , \17873 );
and \g445001/U$2 ( \17875 , \17868 , \17871 , \17874 );
nor \g445001/U$1 ( \17876 , \17875 , \16618 );
and \g445804/U$2 ( \17877 , RIfc6c008_6251, \16341 );
and \g445804/U$3 ( \17878 , RIe200e50_4300, \16377 );
and \g448627/U$2 ( \17879 , RIfcddbb8_7545, \16319 );
and \g448627/U$3 ( \17880 , \16344 , RIfcaf100_7014);
and \g448627/U$4 ( \17881 , RIfc73d30_6340, \16356 );
nor \g448627/U$1 ( \17882 , \17879 , \17880 , \17881 );
and \g451036/U$2 ( \17883 , \16368 , RIe1fbcc0_4242);
and \g451036/U$3 ( \17884 , RIe1fcf08_4255, \16371 );
nor \g451036/U$1 ( \17885 , \17883 , \17884 );
and \g454888/U$2 ( \17886 , \16317 , RIfca8620_6938);
and \g454888/U$3 ( \17887 , RIfcdda50_7544, \16325 );
nor \g454888/U$1 ( \17888 , \17886 , \17887 );
not \g449655/U$3 ( \17889 , \17888 );
not \g449655/U$4 ( \17890 , \16351 );
and \g449655/U$2 ( \17891 , \17889 , \17890 );
and \g449655/U$5 ( \17892 , \16328 , RIfceb5b0_7700);
nor \g449655/U$1 ( \17893 , \17891 , \17892 );
and \g451034/U$2 ( \17894 , \16334 , RIfcdcad8_7533);
and \g451034/U$3 ( \17895 , RIfc71468_6311, \16380 );
nor \g451034/U$1 ( \17896 , \17894 , \17895 );
nand \g447527/U$1 ( \17897 , \17882 , \17885 , \17893 , \17896 );
nor \g445804/U$1 ( \17898 , \17877 , \17878 , \17897 );
and \g451029/U$2 ( \17899 , \16361 , RIfca92c8_6947);
and \g451029/U$3 ( \17900 , RIe202a70_4320, \16313 );
nor \g451029/U$1 ( \17901 , \17899 , \17900 );
and \g451030/U$2 ( \17902 , \16364 , RIfca9700_6950);
and \g451030/U$3 ( \17903 , RIfcdd1e0_7538, \16398 );
nor \g451030/U$1 ( \17904 , \17902 , \17903 );
and \g445004/U$2 ( \17905 , \17898 , \17901 , \17904 );
nor \g445004/U$1 ( \17906 , \17905 , \16393 );
or \g444207/U$1 ( \17907 , \17846 , \17876 , \17906 );
_DC \g35fb/U$1 ( \17908 , \17907 , \16652 );
and \g453386/U$2 ( \17909 , \16377 , RIe198210_3108);
and \g453386/U$3 ( \17910 , RIe192810_3044, \16380 );
nor \g453386/U$1 ( \17911 , \17909 , \17910 );
and \g446336/U$2 ( \17912 , RIe19af10_3140, \16321 );
and \g446336/U$3 ( \17913 , RIfec1590_8320, \16313 );
and \g449315/U$2 ( \17914 , RIe181a10_2852, \16337 );
and \g449315/U$3 ( \17915 , \16341 , RIfc88370_6572);
and \g449315/U$4 ( \17916 , RIe195510_3076, \16344 );
nor \g449315/U$1 ( \17917 , \17914 , \17915 , \17916 );
and \g454213/U$2 ( \17918 , \16317 , RIe187410_2916);
and \g454213/U$3 ( \17919 , RIe18a110_2948, \16325 );
nor \g454213/U$1 ( \17920 , \17918 , \17919 );
not \g450332/U$3 ( \17921 , \17920 );
not \g450332/U$4 ( \17922 , \16351 );
and \g450332/U$2 ( \17923 , \17921 , \17922 );
and \g450332/U$5 ( \17924 , \16356 , RIfec1428_8319);
nor \g450332/U$1 ( \17925 , \17923 , \17924 );
and \g453394/U$2 ( \17926 , \16361 , RIe17c010_2788);
and \g453394/U$3 ( \17927 , RIe17ed10_2820, \16364 );
nor \g453394/U$1 ( \17928 , \17926 , \17927 );
and \g453392/U$2 ( \17929 , \16368 , RIe184710_2884);
and \g453392/U$3 ( \17930 , RIfec12c0_8318, \16371 );
nor \g453392/U$1 ( \17931 , \17929 , \17930 );
nand \g447891/U$1 ( \17932 , \17917 , \17925 , \17928 , \17931 );
nor \g446336/U$1 ( \17933 , \17912 , \17913 , \17932 );
and \g453385/U$2 ( \17934 , \16334 , RIe18fb10_3012);
and \g453385/U$3 ( \17935 , RIe19dc10_3172, \16328 );
nor \g453385/U$1 ( \17936 , \17934 , \17935 );
nand \g445662/U$1 ( \17937 , \17911 , \17933 , \17936 );
not \g448483/U$1 ( \17938 , \16618 );
and \g444798/U$2 ( \17939 , \17937 , \17938 );
and \g449310/U$2 ( \17940 , RIf15e720_5534, \16427 );
and \g449310/U$3 ( \17941 , \16448 , RIf160610_5556);
and \g449310/U$4 ( \17942 , RIfc50ab0_5940, \16485 );
nor \g449310/U$1 ( \17943 , \17940 , \17941 , \17942 );
and \g455323/U$2 ( \17944 , \16317 , RIfc86480_6550);
and \g455323/U$3 ( \17945 , RIfce7668_7655, \16325 );
nor \g455323/U$1 ( \17946 , \17944 , \17945 );
not \g455322/U$1 ( \17947 , \17946 );
and \g450328/U$2 ( \17948 , \17947 , \16336 );
and \g450328/U$3 ( \17949 , RIfc58c10_6032, \16354 );
nor \g450328/U$1 ( \17950 , \17948 , \17949 );
and \g453378/U$2 ( \17951 , \16361 , RIfcb01e0_7026);
and \g453378/U$3 ( \17952 , RIfcd2218_7413, \16364 );
nor \g453378/U$1 ( \17953 , \17951 , \17952 );
and \g453375/U$2 ( \17954 , \16368 , RIfe87f48_7891);
and \g453375/U$3 ( \17955 , RIfe87c78_7889, \16371 );
nor \g453375/U$1 ( \17956 , \17954 , \17955 );
nand \g448108/U$1 ( \17957 , \17943 , \17950 , \17953 , \17956 );
and \g444798/U$3 ( \17958 , \16394 , \17957 );
nor \g444798/U$1 ( \17959 , \17939 , \17958 );
and \g447098/U$2 ( \17960 , \16705 , RIfccd1f0_7356);
and \g447098/U$3 ( \17961 , RIfccd790_7360, \16707 );
nor \g447098/U$1 ( \17962 , \17960 , \17961 );
and \g447097/U$2 ( \17963 , \16710 , RIf1662e0_5622);
and \g447097/U$3 ( \17964 , RIfca6460_6914, \16712 );
nor \g447097/U$1 ( \17965 , \17963 , \17964 );
and \g447099/U$2 ( \17966 , \16715 , RIfe87b10_7888);
and \g447099/U$3 ( \17967 , RIe202908_4319, \16717 );
nor \g447099/U$1 ( \17968 , \17966 , \17967 );
nand \g444528/U$1 ( \17969 , \17959 , \17962 , \17965 , \17968 );
and \g453349/U$2 ( \17970 , \16380 , RIfc4ea58_5917);
and \g453349/U$3 ( \17971 , RIfc5f858_6109, \16321 );
nor \g453349/U$1 ( \17972 , \17970 , \17971 );
and \g446329/U$2 ( \17973 , RIfc6ccb0_6260, \16328 );
and \g446329/U$3 ( \17974 , RIe175f08_2719, \16377 );
and \g449303/U$2 ( \17975 , RIfc5ac68_6055, \16427 );
and \g449303/U$3 ( \17976 , \16448 , RIfca3b98_6885);
and \g449303/U$4 ( \17977 , RIfcc6008_7275, \16485 );
nor \g449303/U$1 ( \17978 , \17975 , \17976 , \17977 );
and \g455235/U$2 ( \17979 , \16317 , RIf16f688_5727);
and \g455235/U$3 ( \17980 , RIfc9b330_6788, \16325 );
nor \g455235/U$1 ( \17981 , \17979 , \17980 );
not \g455234/U$1 ( \17982 , \17981 );
and \g450320/U$2 ( \17983 , \17982 , \16336 );
and \g450320/U$3 ( \17984 , RIfc81020_6490, \16354 );
nor \g450320/U$1 ( \17985 , \17983 , \17984 );
and \g453359/U$2 ( \17986 , \16361 , RIfc5f588_6107);
and \g453359/U$3 ( \17987 , RIfc42410_5776, \16364 );
nor \g453359/U$1 ( \17988 , \17986 , \17987 );
and \g453357/U$2 ( \17989 , \16368 , RIe173d48_2695);
and \g453357/U$3 ( \17990 , RIfc984c8_6755, \16371 );
nor \g453357/U$1 ( \17991 , \17989 , \17990 );
nand \g448107/U$1 ( \17992 , \17978 , \17985 , \17988 , \17991 );
nor \g446329/U$1 ( \17993 , \17973 , \17974 , \17992 );
and \g453353/U$2 ( \17994 , \16334 , RIfc42140_5774);
and \g453353/U$3 ( \17995 , RIfca88f0_6940, \16313 );
nor \g453353/U$1 ( \17996 , \17994 , \17995 );
nand \g445660/U$1 ( \17997 , \17972 , \17993 , \17996 );
not \g448459/U$1 ( \17998 , \16649 );
and \g444797/U$2 ( \17999 , \17997 , \17998 );
and \g449300/U$2 ( \18000 , RIe213168_4507, \16427 );
and \g449300/U$3 ( \18001 , \16448 , RIfe87de0_7890);
and \g449300/U$4 ( \18002 , RIe21e568_4635, \16344 );
nor \g449300/U$1 ( \18003 , \18000 , \18001 , \18002 );
and \g455241/U$2 ( \18004 , \16317 , RIe20d768_4443);
and \g455241/U$3 ( \18005 , RIfcdf670_7564, \16325 );
nor \g455241/U$1 ( \18006 , \18004 , \18005 );
not \g455240/U$1 ( \18007 , \18006 );
and \g450317/U$2 ( \18008 , \18007 , \16336 );
and \g450317/U$3 ( \18009 , RIfc86cf0_6556, \16356 );
nor \g450317/U$1 ( \18010 , \18008 , \18009 );
and \g453340/U$2 ( \18011 , \16361 , RIe207d68_4379);
and \g453340/U$3 ( \18012 , RIe20aa68_4411, \16364 );
nor \g453340/U$1 ( \18013 , \18011 , \18012 );
and \g453339/U$2 ( \18014 , \16368 , RIe210468_4475);
and \g453339/U$3 ( \18015 , RIf1692b0_5656, \16371 );
nor \g453339/U$1 ( \18016 , \18014 , \18015 );
nand \g448105/U$1 ( \18017 , \18003 , \18010 , \18013 , \18016 );
and \g444797/U$3 ( \18018 , \16390 , \18017 );
nor \g444797/U$1 ( \18019 , \17999 , \18018 );
nor \g448331/U$1 ( \18020 , \16389 , \16320 );
and \g447091/U$2 ( \18021 , \18020 , RIe223f68_4699);
nor \g448330/U$1 ( \18022 , \16389 , \16327 );
and \g447091/U$3 ( \18023 , RIfe880b0_7892, \18022 );
nor \g447091/U$1 ( \18024 , \18021 , \18023 );
nor \g448333/U$1 ( \18025 , \16389 , \16517 );
and \g447092/U$2 ( \18026 , \18025 , RIe221268_4667);
nor \g448332/U$1 ( \18027 , \16389 , \16520 );
and \g447092/U$3 ( \18028 , RIf16bfb0_5688, \18027 );
nor \g447092/U$1 ( \18029 , \18026 , \18028 );
nor \g448335/U$1 ( \18030 , \16389 , \16510 );
and \g447093/U$2 ( \18031 , \18030 , RIe215e68_4539);
nor \g448334/U$1 ( \18032 , \16389 , \16513 );
and \g447093/U$3 ( \18033 , RIe218b68_4571, \18032 );
nor \g447093/U$1 ( \18034 , \18031 , \18033 );
nand \g444526/U$1 ( \18035 , \18019 , \18024 , \18029 , \18034 );
and \g446318/U$2 ( \18036 , RIfce0b88_7579, \16328 );
and \g446318/U$3 ( \18037 , RIe1b76b0_3464, \16377 );
and \g449292/U$2 ( \18038 , RIfce9af8_7681, \16427 );
and \g449292/U$3 ( \18039 , \16432 , RIfc89f90_6592);
and \g449292/U$4 ( \18040 , RIfc8a260_6594, \16337 );
nor \g449292/U$1 ( \18041 , \18038 , \18039 , \18040 );
and \g453308/U$2 ( \18042 , \16368 , RIe1b0ea0_3390);
and \g453308/U$3 ( \18043 , RIe1b2958_3409, \16371 );
nor \g453308/U$1 ( \18044 , \18042 , \18043 );
and \g455256/U$2 ( \18045 , \16317 , RIfcb69f0_7100);
and \g455256/U$3 ( \18046 , RIfcd5bc0_7454, \16325 );
nor \g455256/U$1 ( \18047 , \18045 , \18046 );
not \g450308/U$3 ( \18048 , \18047 );
not \g450308/U$4 ( \18049 , \16330 );
and \g450308/U$2 ( \18050 , \18048 , \18049 );
and \g450308/U$5 ( \18051 , \16341 , RIfc4a138_5865);
nor \g450308/U$1 ( \18052 , \18050 , \18051 );
and \g453307/U$2 ( \18053 , \16334 , RIe1b4140_3426);
and \g453307/U$3 ( \18054 , RIe1b54f0_3440, \16380 );
nor \g453307/U$1 ( \18055 , \18053 , \18054 );
nand \g447409/U$1 ( \18056 , \18041 , \18044 , \18052 , \18055 );
nor \g446318/U$1 ( \18057 , \18036 , \18037 , \18056 );
and \g453304/U$2 ( \18058 , \16361 , RIe1ab1d0_3324);
and \g453304/U$3 ( \18059 , RIe1b9708_3487, \16313 );
nor \g453304/U$1 ( \18060 , \18058 , \18059 );
and \g453301/U$2 ( \18061 , \16364 , RIe1ac850_3340);
and \g453301/U$3 ( \18062 , RIfc82808_6507, \16319 );
nor \g453301/U$1 ( \18063 , \18061 , \18062 );
and \g445375/U$2 ( \18064 , \18057 , \18060 , \18063 );
nor \g445375/U$1 ( \18065 , \18064 , \16909 );
and \g446321/U$2 ( \18066 , RIe1ff0c8_4279, \16427 );
and \g446321/U$3 ( \18067 , RIe1f0fc8_4119, \16368 );
and \g449296/U$2 ( \18068 , RIe1a6310_3268, \16321 );
and \g449296/U$3 ( \18069 , \16326 , RIe1a9010_3300);
and \g449296/U$4 ( \18070 , RIe1bbfd0_3516, \16398 );
nor \g449296/U$1 ( \18071 , \18068 , \18069 , \18070 );
and \g455247/U$2 ( \18072 , \16317 , RIe179310_2756);
and \g455247/U$3 ( \18073 , RIe18ce10_2980, \16325 );
nor \g455247/U$1 ( \18074 , \18072 , \18073 );
not \g450312/U$3 ( \18075 , \18074 );
not \g450312/U$4 ( \18076 , \16330 );
and \g450312/U$2 ( \18077 , \18075 , \18076 );
and \g450312/U$5 ( \18078 , \16339 , RIe1d54d0_3804);
nor \g450312/U$1 ( \18079 , \18077 , \18078 );
and \g453326/U$2 ( \18080 , \16377 , RIe1a0910_3204);
and \g453326/U$3 ( \18081 , RIe1a3610_3236, \16313 );
nor \g453326/U$1 ( \18082 , \18080 , \18081 );
and \g453328/U$2 ( \18083 , \16334 , RIe21b868_4603);
and \g453328/U$3 ( \18084 , RIe226c68_4731, \16380 );
nor \g453328/U$1 ( \18085 , \18083 , \18084 );
nand \g447411/U$1 ( \18086 , \18071 , \18079 , \18082 , \18085 );
nor \g446321/U$1 ( \18087 , \18066 , \18067 , \18086 );
and \g453323/U$2 ( \18088 , \16361 , RIe171480_2666);
and \g453323/U$3 ( \18089 , RIe205068_4347, \16432 );
nor \g453323/U$1 ( \18090 , \18088 , \18089 );
and \g453319/U$2 ( \18091 , \16364 , RIe1aee48_3367);
and \g453319/U$3 ( \18092 , RIe1f8480_4202, \16371 );
nor \g453319/U$1 ( \18093 , \18091 , \18092 );
and \g445380/U$2 ( \18094 , \18087 , \18090 , \18093 );
nor \g445380/U$1 ( \18095 , \18094 , \16586 );
or \g444320/U$1 ( \18096 , \17969 , \18035 , \18065 , \18095 );
and \g446310/U$2 ( \18097 , RIfc84158_6525, \16319 );
and \g446310/U$3 ( \18098 , RIfc4b920_5882, \16313 );
and \g449286/U$2 ( \18099 , RIf151ca0_5390, \16427 );
and \g449286/U$3 ( \18100 , \16448 , RIf153488_5407);
and \g449286/U$4 ( \18101 , RIfcb7530_7108, \16344 );
nor \g449286/U$1 ( \18102 , \18099 , \18100 , \18101 );
and \g454435/U$2 ( \18103 , \16317 , RIfcbaaa0_7146);
and \g454435/U$3 ( \18104 , RIfc9aef8_6785, \16325 );
nor \g454435/U$1 ( \18105 , \18103 , \18104 );
not \g454434/U$1 ( \18106 , \18105 );
and \g450300/U$2 ( \18107 , \18106 , \16336 );
and \g450300/U$3 ( \18108 , RIfc4ba88_5883, \16354 );
nor \g450300/U$1 ( \18109 , \18107 , \18108 );
and \g453277/U$2 ( \18110 , \16361 , RIe1ee430_4088);
and \g453277/U$3 ( \18111 , RIfc52130_5956, \16364 );
nor \g453277/U$1 ( \18112 , \18110 , \18111 );
and \g453276/U$2 ( \18113 , \16368 , RIe1f3728_4147);
and \g453276/U$3 ( \18114 , RIfc51e60_5954, \16371 );
nor \g453276/U$1 ( \18115 , \18113 , \18114 );
nand \g448101/U$1 ( \18116 , \18102 , \18109 , \18112 , \18115 );
nor \g446310/U$1 ( \18117 , \18097 , \18098 , \18116 );
and \g453272/U$2 ( \18118 , \16377 , RIe1fa4d8_4225);
and \g453272/U$3 ( \18119 , RIfcd58f0_7452, \16380 );
nor \g453272/U$1 ( \18120 , \18118 , \18119 );
and \g453269/U$2 ( \18121 , \16334 , RIe1f5a50_4172);
and \g453269/U$3 ( \18122 , RIfc47b40_5838, \16328 );
nor \g453269/U$1 ( \18123 , \18121 , \18122 );
and \g445370/U$2 ( \18124 , \18117 , \18120 , \18123 );
nor \g445370/U$1 ( \18125 , \18124 , \16480 );
and \g446314/U$2 ( \18126 , RIe1e62d0_3996, \16313 );
and \g446314/U$3 ( \18127 , RIe1c19d0_3580, \16364 );
and \g449288/U$2 ( \18128 , RIe1cfad0_3740, \16427 );
and \g449288/U$3 ( \18129 , \16448 , RIe1d27d0_3772);
and \g449288/U$4 ( \18130 , RIe1e8fd0_4028, \16319 );
nor \g449288/U$1 ( \18131 , \18128 , \18129 , \18130 );
and \g453290/U$2 ( \18132 , \16368 , RIe1ca0d0_3676);
and \g453290/U$3 ( \18133 , RIe1ccdd0_3708, \16371 );
nor \g453290/U$1 ( \18134 , \18132 , \18133 );
and \g455309/U$2 ( \18135 , \16317 , RIe1ddbd0_3900);
and \g455309/U$3 ( \18136 , RIe1e08d0_3932, \16325 );
nor \g455309/U$1 ( \18137 , \18135 , \18136 );
not \g450304/U$3 ( \18138 , \18137 );
not \g450304/U$4 ( \18139 , \16330 );
and \g450304/U$2 ( \18140 , \18138 , \18139 );
and \g450304/U$5 ( \18141 , \16328 , RIe1ebcd0_4060);
nor \g450304/U$1 ( \18142 , \18140 , \18141 );
and \g453289/U$2 ( \18143 , \16334 , RIe1d81d0_3836);
and \g453289/U$3 ( \18144 , RIe1daed0_3868, \16380 );
nor \g453289/U$1 ( \18145 , \18143 , \18144 );
nand \g447879/U$1 ( \18146 , \18131 , \18134 , \18142 , \18145 );
nor \g446314/U$1 ( \18147 , \18126 , \18127 , \18146 );
and \g453282/U$2 ( \18148 , \16341 , RIe1c73d0_3644);
and \g453282/U$3 ( \18149 , RIe1e35d0_3964, \16377 );
nor \g453282/U$1 ( \18150 , \18148 , \18149 );
and \g453285/U$2 ( \18151 , \16361 , RIe1becd0_3548);
and \g453285/U$3 ( \18152 , RIe1c46d0_3612, \16398 );
nor \g453285/U$1 ( \18153 , \18151 , \18152 );
and \g445373/U$2 ( \18154 , \18147 , \18150 , \18153 );
nor \g445373/U$1 ( \18155 , \18154 , \16555 );
or \g444263/U$1 ( \18156 , \18096 , \18125 , \18155 );
_DC \g3680/U$1 ( \18157 , \18156 , \16652 );
and \g453641/U$2 ( \18158 , \16364 , RIfc93338_6697);
and \g453641/U$3 ( \18159 , RIfe872a0_7882, \16371 );
nor \g453641/U$1 ( \18160 , \18158 , \18159 );
and \g446390/U$2 ( \18161 , RIf15e5b8_5533, \16427 );
and \g446390/U$3 ( \18162 , RIfe87138_7881, \16368 );
and \g449384/U$2 ( \18163 , RIfcdf940_7566, \16485 );
and \g449384/U$3 ( \18164 , \16356 , RIfcb2670_7052);
and \g449384/U$4 ( \18165 , RIfec1158_8317, \16398 );
nor \g449384/U$1 ( \18166 , \18163 , \18164 , \18165 );
and \g455354/U$2 ( \18167 , \16317 , RIfcd73a8_7471);
and \g455354/U$3 ( \18168 , RIfc5af38_6057, \16325 );
nor \g455354/U$1 ( \18169 , \18167 , \18168 );
not \g450403/U$3 ( \18170 , \18169 );
not \g450403/U$4 ( \18171 , \16311 );
and \g450403/U$2 ( \18172 , \18170 , \18171 );
and \g450403/U$5 ( \18173 , \16341 , RIfc78920_6394);
nor \g450403/U$1 ( \18174 , \18172 , \18173 );
and \g453646/U$2 ( \18175 , \16377 , RIe200ce8_4299);
and \g453646/U$3 ( \18176 , RIe2027a0_4318, \16313 );
nor \g453646/U$1 ( \18177 , \18175 , \18176 );
and \g453651/U$2 ( \18178 , \16334 , RIfcbf3c0_7198);
and \g453651/U$3 ( \18179 , RIfc5b208_6059, \16380 );
nor \g453651/U$1 ( \18180 , \18178 , \18179 );
nand \g447420/U$1 ( \18181 , \18166 , \18174 , \18177 , \18180 );
nor \g446390/U$1 ( \18182 , \18161 , \18162 , \18181 );
and \g453642/U$2 ( \18183 , \16361 , RIfcea368_7687);
and \g453642/U$3 ( \18184 , RIf1604a8_5555, \16448 );
nor \g453642/U$1 ( \18185 , \18183 , \18184 );
nand \g445677/U$1 ( \18186 , \18160 , \18182 , \18185 );
and \g444803/U$2 ( \18187 , \18186 , \16394 );
and \g449380/U$2 ( \18188 , RIe213000_4506, \16427 );
and \g449380/U$3 ( \18189 , \16448 , RIfc79e38_6409);
and \g449380/U$4 ( \18190 , RIe21e400_4634, \16485 );
nor \g449380/U$1 ( \18191 , \18188 , \18189 , \18190 );
and \g455145/U$2 ( \18192 , \16317 , RIe20d600_4442);
and \g455145/U$3 ( \18193 , RIf168068_5643, \16325 );
nor \g455145/U$1 ( \18194 , \18192 , \18193 );
not \g455144/U$1 ( \18195 , \18194 );
and \g450399/U$2 ( \18196 , \18195 , \16336 );
and \g450399/U$3 ( \18197 , RIfc920f0_6684, \16356 );
nor \g450399/U$1 ( \18198 , \18196 , \18197 );
and \g453630/U$2 ( \18199 , \16361 , RIe207c00_4378);
and \g453630/U$3 ( \18200 , RIe20a900_4410, \16364 );
nor \g453630/U$1 ( \18201 , \18199 , \18200 );
and \g453627/U$2 ( \18202 , \16368 , RIe210300_4474);
and \g453627/U$3 ( \18203 , RIfcbee20_7194, \16371 );
nor \g453627/U$1 ( \18204 , \18202 , \18203 );
nand \g448115/U$1 ( \18205 , \18191 , \18198 , \18201 , \18204 );
and \g444803/U$3 ( \18206 , \16390 , \18205 );
nor \g444803/U$1 ( \18207 , \18187 , \18206 );
and \g447139/U$2 ( \18208 , \18020 , RIe223e00_4698);
and \g447139/U$3 ( \18209 , RIfea9710_8244, \18022 );
nor \g447139/U$1 ( \18210 , \18208 , \18209 );
and \g447140/U$2 ( \18211 , \18025 , RIe221100_4666);
and \g447140/U$3 ( \18212 , RIfcd8488_7483, \18027 );
nor \g447140/U$1 ( \18213 , \18211 , \18212 );
and \g447141/U$2 ( \18214 , \18030 , RIe215d00_4538);
and \g447141/U$3 ( \18215 , RIe218a00_4570, \18032 );
nor \g447141/U$1 ( \18216 , \18214 , \18215 );
nand \g444535/U$1 ( \18217 , \18207 , \18210 , \18213 , \18216 );
and \g453671/U$2 ( \18218 , \16377 , RIe1fa370_4224);
and \g453671/U$3 ( \18219 , RIfcbf960_7202, \16380 );
nor \g453671/U$1 ( \18220 , \18218 , \18219 );
and \g446397/U$2 ( \18221 , RIfc5bbe0_6066, \16319 );
and \g446397/U$3 ( \18222 , RIfcede78_7729, \16313 );
and \g449394/U$2 ( \18223 , RIfce1b00_7590, \16398 );
and \g449394/U$3 ( \18224 , \16339 , RIfcb1f68_7047);
and \g449394/U$4 ( \18225 , RIfce1dd0_7592, \16485 );
nor \g449394/U$1 ( \18226 , \18223 , \18224 , \18225 );
and \g455188/U$2 ( \18227 , \16317 , RIfc78380_6390);
and \g455188/U$3 ( \18228 , RIfcbfc30_7204, \16325 );
nor \g455188/U$1 ( \18229 , \18227 , \18228 );
not \g450413/U$3 ( \18230 , \18229 );
not \g450413/U$4 ( \18231 , \16351 );
and \g450413/U$2 ( \18232 , \18230 , \18231 );
and \g450413/U$5 ( \18233 , \16356 , RIfcd4c48_7443);
nor \g450413/U$1 ( \18234 , \18232 , \18233 );
and \g453676/U$2 ( \18235 , \16361 , RIe1ee2c8_4087);
and \g453676/U$3 ( \18236 , RIfc93a40_6702, \16364 );
nor \g453676/U$1 ( \18237 , \18235 , \18236 );
and \g453674/U$2 ( \18238 , \16368 , RIe1f35c0_4146);
and \g453674/U$3 ( \18239 , RIfc93770_6700, \16371 );
nor \g453674/U$1 ( \18240 , \18238 , \18239 );
nand \g447940/U$1 ( \18241 , \18226 , \18234 , \18237 , \18240 );
nor \g446397/U$1 ( \18242 , \18221 , \18222 , \18241 );
and \g453670/U$2 ( \18243 , \16334 , RIe1f58e8_4171);
and \g453670/U$3 ( \18244 , RIfcb23a0_7050, \16328 );
nor \g453670/U$1 ( \18245 , \18243 , \18244 );
nand \g445679/U$1 ( \18246 , \18220 , \18242 , \18245 );
and \g444836/U$2 ( \18247 , \18246 , \16481 );
and \g449388/U$2 ( \18248 , RIfcd7c18_7477, \16427 );
and \g449388/U$3 ( \18249 , \16448 , RIfc94850_6712);
and \g449388/U$4 ( \18250 , RIfceabd8_7693, \16485 );
nor \g449388/U$1 ( \18251 , \18248 , \18249 , \18250 );
and \g455358/U$2 ( \18252 , \16317 , RIfce2640_7598);
and \g455358/U$3 ( \18253 , RIfc76a30_6372, \16325 );
nor \g455358/U$1 ( \18254 , \18252 , \18253 );
not \g455357/U$1 ( \18255 , \18254 );
and \g450409/U$2 ( \18256 , \18255 , \16336 );
and \g450409/U$3 ( \18257 , RIfcd12a0_7402, \16354 );
nor \g450409/U$1 ( \18258 , \18256 , \18257 );
and \g453664/U$2 ( \18259 , \16361 , RIe1ab068_3323);
and \g453664/U$3 ( \18260 , RIe1ac6e8_3339, \16364 );
nor \g453664/U$1 ( \18261 , \18259 , \18260 );
and \g453661/U$2 ( \18262 , \16368 , RIe1b0d38_3389);
and \g453661/U$3 ( \18263 , RIe1b27f0_3408, \16371 );
nor \g453661/U$1 ( \18264 , \18262 , \18263 );
nand \g448116/U$1 ( \18265 , \18251 , \18258 , \18261 , \18264 );
and \g444836/U$3 ( \18266 , \16477 , \18265 );
nor \g444836/U$1 ( \18267 , \18247 , \18266 );
nor \g448276/U$1 ( \18268 , \16909 , \16320 );
and \g447147/U$2 ( \18269 , \18268 , RIfc94148_6707);
nor \g448272/U$1 ( \18270 , \16909 , \16327 );
and \g447147/U$3 ( \18271 , RIfcdec98_7557, \18270 );
nor \g447147/U$1 ( \18272 , \18269 , \18271 );
nor \g448292/U$1 ( \18273 , \16909 , \16517 );
and \g447148/U$2 ( \18274 , \18273 , RIe1b7548_3463);
nor \g448277/U$1 ( \18275 , \16909 , \16520 );
and \g447148/U$3 ( \18276 , RIe1b95a0_3486, \18275 );
nor \g447148/U$1 ( \18277 , \18274 , \18276 );
nor \g448294/U$1 ( \18278 , \16909 , \16510 );
and \g447150/U$2 ( \18279 , \18278 , RIe1b3fd8_3425);
nor \g448293/U$1 ( \18280 , \16909 , \16513 );
and \g447150/U$3 ( \18281 , RIe1b5388_3439, \18280 );
nor \g447150/U$1 ( \18282 , \18279 , \18281 );
nand \g444657/U$1 ( \18283 , \18267 , \18272 , \18277 , \18282 );
and \g446381/U$2 ( \18284 , RIfc915b0_6676, \16328 );
and \g446381/U$3 ( \18285 , RIfc96e48_6739, \16334 );
and \g449371/U$2 ( \18286 , RIfc96ce0_6738, \16427 );
and \g449371/U$3 ( \18287 , \16448 , RIfc7a810_6416);
and \g449371/U$4 ( \18288 , RIfcc7958_7293, \16344 );
nor \g449371/U$1 ( \18289 , \18286 , \18287 , \18288 );
and \g454314/U$2 ( \18290 , \16317 , RIfc7a540_6414);
and \g454314/U$3 ( \18291 , RIfce39f0_7612, \16325 );
nor \g454314/U$1 ( \18292 , \18290 , \18291 );
not \g454313/U$1 ( \18293 , \18292 );
and \g450391/U$2 ( \18294 , \18293 , \16336 );
and \g450391/U$3 ( \18295 , RIfceb448_7699, \16356 );
nor \g450391/U$1 ( \18296 , \18294 , \18295 );
and \g453601/U$2 ( \18297 , \16361 , RIfc429b0_5780);
and \g453601/U$3 ( \18298 , RIfc91b50_6680, \16364 );
nor \g453601/U$1 ( \18299 , \18297 , \18298 );
and \g453598/U$2 ( \18300 , \16368 , RIe173be0_2694);
and \g453598/U$3 ( \18301 , RIfcc7ac0_7294, \16371 );
nor \g453598/U$1 ( \18302 , \18300 , \18301 );
nand \g448114/U$1 ( \18303 , \18289 , \18296 , \18299 , \18302 );
nor \g446381/U$1 ( \18304 , \18284 , \18285 , \18303 );
and \g453595/U$2 ( \18305 , \16377 , RIe175da0_2718);
and \g453595/U$3 ( \18306 , RIfc42de8_5783, \16380 );
nor \g453595/U$1 ( \18307 , \18305 , \18306 );
and \g453593/U$2 ( \18308 , \16313 , RIfce3b58_7613);
and \g453593/U$3 ( \18309 , RIfcbe5b0_7188, \16319 );
nor \g453593/U$1 ( \18310 , \18308 , \18309 );
and \g445417/U$2 ( \18311 , \18304 , \18307 , \18310 );
nor \g445417/U$1 ( \18312 , \18311 , \16649 );
and \g446385/U$2 ( \18313 , RIe19daa8_3171, \16328 );
and \g446385/U$3 ( \18314 , RIe18f9a8_3011, \16334 );
and \g449375/U$2 ( \18315 , RIe1818a8_2851, \16398 );
and \g449375/U$3 ( \18316 , \16341 , RIfc912e0_6674);
and \g449375/U$4 ( \18317 , RIe1953a8_3075, \16485 );
nor \g449375/U$1 ( \18318 , \18315 , \18316 , \18317 );
and \g455148/U$2 ( \18319 , \16317 , RIe1872a8_2915);
and \g455148/U$3 ( \18320 , RIe189fa8_2947, \16325 );
nor \g455148/U$1 ( \18321 , \18319 , \18320 );
not \g450396/U$3 ( \18322 , \18321 );
not \g450396/U$4 ( \18323 , \16351 );
and \g450396/U$2 ( \18324 , \18322 , \18323 );
and \g450396/U$5 ( \18325 , \16354 , RIf1449b0_5240);
nor \g450396/U$1 ( \18326 , \18324 , \18325 );
and \g453618/U$2 ( \18327 , \16361 , RIe17bea8_2787);
and \g453618/U$3 ( \18328 , RIe17eba8_2819, \16364 );
nor \g453618/U$1 ( \18329 , \18327 , \18328 );
and \g453616/U$2 ( \18330 , \16368 , RIe1845a8_2883);
and \g453616/U$3 ( \18331 , RIf143ba0_5230, \16371 );
nor \g453616/U$1 ( \18332 , \18330 , \18331 );
nand \g447930/U$1 ( \18333 , \18318 , \18326 , \18329 , \18332 );
nor \g446385/U$1 ( \18334 , \18313 , \18314 , \18333 );
and \g453613/U$2 ( \18335 , \16377 , RIe1980a8_3107);
and \g453613/U$3 ( \18336 , RIe1926a8_3043, \16380 );
nor \g453613/U$1 ( \18337 , \18335 , \18336 );
and \g453611/U$2 ( \18338 , \16313 , RIf1457c0_5250);
and \g453611/U$3 ( \18339 , RIe19ada8_3139, \16321 );
nor \g453611/U$1 ( \18340 , \18338 , \18339 );
and \g445420/U$2 ( \18341 , \18334 , \18337 , \18340 );
nor \g445420/U$1 ( \18342 , \18341 , \16618 );
or \g444409/U$1 ( \18343 , \18217 , \18283 , \18312 , \18342 );
and \g446374/U$2 ( \18344 , RIe1d2668_3771, \16432 );
and \g446374/U$3 ( \18345 , RIe1ccc68_3707, \16371 );
and \g449361/U$2 ( \18346 , RIe1e8e68_4027, \16321 );
and \g449361/U$3 ( \18347 , \16328 , RIe1ebb68_4059);
and \g449361/U$4 ( \18348 , RIe1c4568_3611, \16398 );
nor \g449361/U$1 ( \18349 , \18346 , \18347 , \18348 );
and \g454577/U$2 ( \18350 , \16317 , RIe1dda68_3899);
and \g454577/U$3 ( \18351 , RIe1e0768_3931, \16325 );
nor \g454577/U$1 ( \18352 , \18350 , \18351 );
not \g450381/U$3 ( \18353 , \18352 );
not \g450381/U$4 ( \18354 , \16330 );
and \g450381/U$2 ( \18355 , \18353 , \18354 );
and \g450381/U$5 ( \18356 , \16341 , RIe1c7268_3643);
nor \g450381/U$1 ( \18357 , \18355 , \18356 );
and \g453565/U$2 ( \18358 , \16377 , RIe1e3468_3963);
and \g453565/U$3 ( \18359 , RIe1e6168_3995, \16313 );
nor \g453565/U$1 ( \18360 , \18358 , \18359 );
and \g453568/U$2 ( \18361 , \16334 , RIe1d8068_3835);
and \g453568/U$3 ( \18362 , RIe1dad68_3867, \16380 );
nor \g453568/U$1 ( \18363 , \18361 , \18362 );
nand \g447417/U$1 ( \18364 , \18349 , \18357 , \18360 , \18363 );
nor \g446374/U$1 ( \18365 , \18344 , \18345 , \18364 );
and \g453556/U$2 ( \18366 , \16364 , RIe1c1868_3579);
and \g453556/U$3 ( \18367 , RIe1c9f68_3675, \16368 );
nor \g453556/U$1 ( \18368 , \18366 , \18367 );
and \g453559/U$2 ( \18369 , \16361 , RIe1beb68_3547);
and \g453559/U$3 ( \18370 , RIe1cf968_3739, \16427 );
nor \g453559/U$1 ( \18371 , \18369 , \18370 );
and \g445409/U$2 ( \18372 , \18365 , \18368 , \18371 );
nor \g445409/U$1 ( \18373 , \18372 , \16555 );
and \g446377/U$2 ( \18374 , RIe1fef60_4278, \16427 );
and \g446377/U$3 ( \18375 , RIe1f0e60_4118, \16368 );
and \g449367/U$2 ( \18376 , RIe1a61a8_3267, \16319 );
and \g449367/U$3 ( \18377 , \16326 , RIe1a8ea8_3299);
and \g449367/U$4 ( \18378 , RIe1bbe68_3515, \16398 );
nor \g449367/U$1 ( \18379 , \18376 , \18377 , \18378 );
and \g455165/U$2 ( \18380 , \16317 , RIe1791a8_2755);
and \g455165/U$3 ( \18381 , RIe18cca8_2979, \16325 );
nor \g455165/U$1 ( \18382 , \18380 , \18381 );
not \g450387/U$3 ( \18383 , \18382 );
not \g450387/U$4 ( \18384 , \16330 );
and \g450387/U$2 ( \18385 , \18383 , \18384 );
and \g450387/U$5 ( \18386 , \16341 , RIe1d5368_3803);
nor \g450387/U$1 ( \18387 , \18385 , \18386 );
and \g453581/U$2 ( \18388 , \16377 , RIe1a07a8_3203);
and \g453581/U$3 ( \18389 , RIe1a34a8_3235, \16313 );
nor \g453581/U$1 ( \18390 , \18388 , \18389 );
and \g453584/U$2 ( \18391 , \16334 , RIe21b700_4602);
and \g453584/U$3 ( \18392 , RIe226b00_4730, \16380 );
nor \g453584/U$1 ( \18393 , \18391 , \18392 );
nand \g447418/U$1 ( \18394 , \18379 , \18387 , \18390 , \18393 );
nor \g446377/U$1 ( \18395 , \18374 , \18375 , \18394 );
and \g453576/U$2 ( \18396 , \16361 , RIe171318_2665);
and \g453576/U$3 ( \18397 , RIe204f00_4346, \16432 );
nor \g453576/U$1 ( \18398 , \18396 , \18397 );
and \g453575/U$2 ( \18399 , \16364 , RIe1aece0_3366);
and \g453575/U$3 ( \18400 , RIe1f8318_4201, \16371 );
nor \g453575/U$1 ( \18401 , \18399 , \18400 );
and \g445412/U$2 ( \18402 , \18395 , \18398 , \18401 );
nor \g445412/U$1 ( \18403 , \18402 , \16586 );
or \g444229/U$1 ( \18404 , \18343 , \18373 , \18403 );
_DC \g3705/U$1 ( \18405 , \18404 , \16652 );
and \g449024/U$2 ( \18406 , RIe195240_3074, \16485 );
and \g449024/U$3 ( \18407 , \16354 , RIf144848_5239);
and \g449024/U$4 ( \18408 , RIe181740_2850, \16398 );
nor \g449024/U$1 ( \18409 , \18406 , \18407 , \18408 );
and \g454800/U$2 ( \18410 , \16317 , RIe19ac40_3138);
and \g454800/U$3 ( \18411 , RIe19d940_3170, \16325 );
nor \g454800/U$1 ( \18412 , \18410 , \18411 );
not \g450038/U$3 ( \18413 , \18412 );
not \g450038/U$4 ( \18414 , \16311 );
and \g450038/U$2 ( \18415 , \18413 , \18414 );
and \g450038/U$5 ( \18416 , \16341 , RIfc6f140_6286);
nor \g450038/U$1 ( \18417 , \18415 , \18416 );
and \g452318/U$2 ( \18418 , \16377 , RIe197f40_3106);
and \g452318/U$3 ( \18419 , RIfc64880_6166, \16313 );
nor \g452318/U$1 ( \18420 , \18418 , \18419 );
and \g452321/U$2 ( \18421 , \16334 , RIe18f840_3010);
and \g452321/U$3 ( \18422 , RIe192540_3042, \16380 );
nor \g452321/U$1 ( \18423 , \18421 , \18422 );
nand \g447347/U$1 ( \18424 , \18409 , \18417 , \18420 , \18423 );
and \g444708/U$2 ( \18425 , \18424 , \17938 );
and \g446116/U$2 ( \18426 , RIfcacb08_6987, \16326 );
and \g446116/U$3 ( \18427 , RIfc67418_6197, \16334 );
and \g449029/U$2 ( \18428 , RIf15ba20_5502, \16398 );
and \g449029/U$3 ( \18429 , \16341 , RIfc6dac0_6270);
and \g449029/U$4 ( \18430 , RIfccad60_7330, \16485 );
nor \g449029/U$1 ( \18431 , \18428 , \18429 , \18430 );
and \g454324/U$2 ( \18432 , \16317 , RIf15e450_5532);
and \g454324/U$3 ( \18433 , RIf160340_5554, \16325 );
nor \g454324/U$1 ( \18434 , \18432 , \18433 );
not \g450042/U$3 ( \18435 , \18434 );
not \g450042/U$4 ( \18436 , \16351 );
and \g450042/U$2 ( \18437 , \18435 , \18436 );
and \g450042/U$5 ( \18438 , \16356 , RIfca8a58_6941);
nor \g450042/U$1 ( \18439 , \18437 , \18438 );
and \g452336/U$2 ( \18440 , \16361 , RIfc6d7f0_6268);
and \g452336/U$3 ( \18441 , RIfc6d958_6269, \16364 );
nor \g452336/U$1 ( \18442 , \18440 , \18441 );
and \g452334/U$2 ( \18443 , \16368 , RIfe81300_7814);
and \g452334/U$3 ( \18444 , RIfe81a08_7819, \16371 );
nor \g452334/U$1 ( \18445 , \18443 , \18444 );
nand \g447741/U$1 ( \18446 , \18431 , \18439 , \18442 , \18445 );
nor \g446116/U$1 ( \18447 , \18426 , \18427 , \18446 );
and \g452329/U$2 ( \18448 , \16377 , RIfe818a0_7818);
and \g452329/U$3 ( \18449 , RIfcac838_6985, \16380 );
nor \g452329/U$1 ( \18450 , \18448 , \18449 );
and \g452328/U$2 ( \18451 , \16313 , RIfea8900_8234);
and \g452328/U$3 ( \18452 , RIfcac9a0_6986, \16319 );
nor \g452328/U$1 ( \18453 , \18451 , \18452 );
and \g445232/U$2 ( \18454 , \18447 , \18450 , \18453 );
nor \g445232/U$1 ( \18455 , \18454 , \16393 );
nor \g444708/U$1 ( \18456 , \18425 , \18455 );
nor \g448390/U$1 ( \18457 , \16618 , \16428 );
and \g446886/U$2 ( \18458 , \18457 , RIe187140_2914);
nor \g448389/U$1 ( \18459 , \16618 , \16433 );
and \g446886/U$3 ( \18460 , RIe189e40_2946, \18459 );
nor \g446886/U$1 ( \18461 , \18458 , \18460 );
nor \g448327/U$1 ( \18462 , \16618 , \16437 );
and \g446887/U$2 ( \18463 , \18462 , RIe184440_2882);
nor \g448391/U$1 ( \18464 , \16618 , \16440 );
and \g446887/U$3 ( \18465 , RIf143a38_5229, \18464 );
nor \g446887/U$1 ( \18466 , \18463 , \18465 );
nor \g448326/U$1 ( \18467 , \16618 , \16418 );
and \g446888/U$2 ( \18468 , \18467 , RIe17bd40_2786);
nor \g448377/U$1 ( \18469 , \16618 , \16421 );
and \g446888/U$3 ( \18470 , RIe17ea40_2818, \18469 );
nor \g446888/U$1 ( \18471 , \18468 , \18470 );
nand \g444499/U$1 ( \18472 , \18456 , \18461 , \18466 , \18471 );
and \g452365/U$2 ( \18473 , \16313 , RIfc66d10_6192);
and \g452365/U$3 ( \18474 , RIe223c98_4697, \16321 );
nor \g452365/U$1 ( \18475 , \18473 , \18474 );
and \g446122/U$2 ( \18476 , RIfe81468_7815, \16328 );
and \g446122/U$3 ( \18477 , RIe215b98_4537, \16334 );
and \g449038/U$2 ( \18478 , RIe212e98_4505, \16427 );
and \g449038/U$3 ( \18479 , \16448 , RIfc3fc38_5751);
and \g449038/U$4 ( \18480 , RIe21e298_4633, \16485 );
nor \g449038/U$1 ( \18481 , \18478 , \18479 , \18480 );
and \g454824/U$2 ( \18482 , \16317 , RIe20d498_4441);
and \g454824/U$3 ( \18483 , RIf167f00_5642, \16325 );
nor \g454824/U$1 ( \18484 , \18482 , \18483 );
not \g454823/U$1 ( \18485 , \18484 );
and \g450051/U$2 ( \18486 , \18485 , \16336 );
and \g450051/U$3 ( \18487 , RIf16b038_5677, \16356 );
nor \g450051/U$1 ( \18488 , \18486 , \18487 );
and \g452373/U$2 ( \18489 , \16361 , RIe207a98_4377);
and \g452373/U$3 ( \18490 , RIe20a798_4409, \16364 );
nor \g452373/U$1 ( \18491 , \18489 , \18490 );
and \g452370/U$2 ( \18492 , \16368 , RIe210198_4473);
and \g452370/U$3 ( \18493 , RIfc67850_6200, \16371 );
nor \g452370/U$1 ( \18494 , \18492 , \18493 );
nand \g448072/U$1 ( \18495 , \18481 , \18488 , \18491 , \18494 );
nor \g446122/U$1 ( \18496 , \18476 , \18477 , \18495 );
and \g452366/U$2 ( \18497 , \16377 , RIe220f98_4665);
and \g452366/U$3 ( \18498 , RIe218898_4569, \16380 );
nor \g452366/U$1 ( \18499 , \18497 , \18498 );
nand \g445607/U$1 ( \18500 , \18475 , \18496 , \18499 );
and \g444741/U$2 ( \18501 , \18500 , \16390 );
and \g449035/U$2 ( \18502 , RIf13f3e8_5179, \16344 );
and \g449035/U$3 ( \18503 , \16356 , RIfccabf8_7329);
and \g449035/U$4 ( \18504 , RIfc6eba0_6282, \16398 );
nor \g449035/U$1 ( \18505 , \18502 , \18503 , \18504 );
and \g454816/U$2 ( \18506 , \16317 , RIf141008_5199);
and \g454816/U$3 ( \18507 , RIfc64f88_6171, \16325 );
nor \g454816/U$1 ( \18508 , \18506 , \18507 );
not \g450047/U$3 ( \18509 , \18508 );
not \g450047/U$4 ( \18510 , \16311 );
and \g450047/U$2 ( \18511 , \18509 , \18510 );
and \g450047/U$5 ( \18512 , \16341 , RIfc66338_6185);
nor \g450047/U$1 ( \18513 , \18511 , \18512 );
and \g452354/U$2 ( \18514 , \16377 , RIfe81738_7817);
and \g452354/U$3 ( \18515 , RIe177150_2732, \16313 );
nor \g452354/U$1 ( \18516 , \18514 , \18515 );
and \g452355/U$2 ( \18517 , \16334 , RIee3d630_5157);
and \g452355/U$3 ( \18518 , RIfca81e8_6935, \16380 );
nor \g452355/U$1 ( \18519 , \18517 , \18518 );
nand \g447348/U$1 ( \18520 , \18505 , \18513 , \18516 , \18519 );
and \g444741/U$3 ( \18521 , \17998 , \18520 );
nor \g444741/U$1 ( \18522 , \18501 , \18521 );
nor \g448263/U$1 ( \18523 , \16649 , \16437 );
and \g446896/U$2 ( \18524 , \18523 , RIe173a78_2693);
nor \g448270/U$1 ( \18525 , \16649 , \16433 );
and \g446896/U$3 ( \18526 , RIfc66068_6183, \18525 );
nor \g446896/U$1 ( \18527 , \18524 , \18526 );
nor \g448269/U$1 ( \18528 , \16649 , \16440 );
and \g446895/U$2 ( \18529 , \18528 , RIfcdde88_7547);
nor \g448268/U$1 ( \18530 , \16649 , \16428 );
and \g446895/U$3 ( \18531 , RIfc6ed08_6283, \18530 );
nor \g446895/U$1 ( \18532 , \18529 , \18531 );
nor \g448262/U$1 ( \18533 , \16649 , \16418 );
and \g446897/U$2 ( \18534 , \18533 , RIfcacdd8_6989);
nor \g448266/U$1 ( \18535 , \16649 , \16421 );
and \g446897/U$3 ( \18536 , RIfc664a0_6186, \18535 );
nor \g446897/U$1 ( \18537 , \18534 , \18536 );
nand \g444615/U$1 ( \18538 , \18522 , \18527 , \18532 , \18537 );
and \g446106/U$2 ( \18539 , RIfc6cf80_6262, \16319 );
and \g446106/U$3 ( \18540 , RIfc6d3b8_6265, \16313 );
and \g449013/U$2 ( \18541 , RIfc68d68_6215, \16427 );
and \g449013/U$3 ( \18542 , \16432 , RIfc6c5a8_6255);
and \g449013/U$4 ( \18543 , RIfcabe60_6978, \16485 );
nor \g449013/U$1 ( \18544 , \18541 , \18542 , \18543 );
and \g454785/U$2 ( \18545 , \16317 , RIfccb8a0_7338);
and \g454785/U$3 ( \18546 , RIfc68a98_6213, \16325 );
nor \g454785/U$1 ( \18547 , \18545 , \18546 );
not \g454784/U$1 ( \18548 , \18547 );
and \g450027/U$2 ( \18549 , \18548 , \16336 );
and \g450027/U$3 ( \18550 , RIfc6d520_6266, \16356 );
nor \g450027/U$1 ( \18551 , \18549 , \18550 );
and \g452286/U$2 ( \18552 , \16361 , RIe1ee160_4086);
and \g452286/U$3 ( \18553 , RIfca9b38_6953, \16364 );
nor \g452286/U$1 ( \18554 , \18552 , \18553 );
and \g452282/U$2 ( \18555 , \16368 , RIe1f3458_4145);
and \g452282/U$3 ( \18556 , RIfc68c00_6214, \16371 );
nor \g452282/U$1 ( \18557 , \18555 , \18556 );
nand \g448069/U$1 ( \18558 , \18544 , \18551 , \18554 , \18557 );
nor \g446106/U$1 ( \18559 , \18539 , \18540 , \18558 );
and \g452279/U$2 ( \18560 , \16377 , RIfe815d0_7816);
and \g452279/U$3 ( \18561 , RIfc6d0e8_6263, \16380 );
nor \g452279/U$1 ( \18562 , \18560 , \18561 );
and \g452275/U$2 ( \18563 , \16334 , RIe1f5780_4170);
and \g452275/U$3 ( \18564 , RIfc587d8_6029, \16328 );
nor \g452275/U$1 ( \18565 , \18563 , \18564 );
and \g445226/U$2 ( \18566 , \18559 , \18562 , \18565 );
nor \g445226/U$1 ( \18567 , \18566 , \16480 );
and \g446110/U$2 ( \18568 , RIe1cf800_3738, \16427 );
and \g446110/U$3 ( \18569 , RIe1c9e00_3674, \16368 );
and \g449019/U$2 ( \18570 , RIe1dd900_3898, \16485 );
and \g449019/U$3 ( \18571 , \16354 , RIe1e0600_3930);
and \g449019/U$4 ( \18572 , RIe1c4400_3610, \16337 );
nor \g449019/U$1 ( \18573 , \18570 , \18571 , \18572 );
and \g454790/U$2 ( \18574 , \16317 , RIe1e8d00_4026);
and \g454790/U$3 ( \18575 , RIe1eba00_4058, \16325 );
nor \g454790/U$1 ( \18576 , \18574 , \18575 );
not \g450032/U$3 ( \18577 , \18576 );
not \g450032/U$4 ( \18578 , \16311 );
and \g450032/U$2 ( \18579 , \18577 , \18578 );
and \g450032/U$5 ( \18580 , \16341 , RIe1c7100_3642);
nor \g450032/U$1 ( \18581 , \18579 , \18580 );
and \g452301/U$2 ( \18582 , \16377 , RIe1e3300_3962);
and \g452301/U$3 ( \18583 , RIe1e6000_3994, \16313 );
nor \g452301/U$1 ( \18584 , \18582 , \18583 );
and \g452305/U$2 ( \18585 , \16334 , RIe1d7f00_3834);
and \g452305/U$3 ( \18586 , RIe1dac00_3866, \16380 );
nor \g452305/U$1 ( \18587 , \18585 , \18586 );
nand \g447344/U$1 ( \18588 , \18573 , \18581 , \18584 , \18587 );
nor \g446110/U$1 ( \18589 , \18568 , \18569 , \18588 );
and \g452296/U$2 ( \18590 , \16361 , RIe1bea00_3546);
and \g452296/U$3 ( \18591 , RIe1d2500_3770, \16448 );
nor \g452296/U$1 ( \18592 , \18590 , \18591 );
and \g452295/U$2 ( \18593 , \16364 , RIe1c1700_3578);
and \g452295/U$3 ( \18594 , RIe1ccb00_3706, \16371 );
nor \g452295/U$1 ( \18595 , \18593 , \18594 );
and \g445230/U$2 ( \18596 , \18589 , \18592 , \18595 );
nor \g445230/U$1 ( \18597 , \18596 , \16555 );
or \g444380/U$1 ( \18598 , \18472 , \18538 , \18567 , \18597 );
and \g446098/U$2 ( \18599 , RIfc6bbd0_6248, \16326 );
and \g446098/U$3 ( \18600 , RIe1b73e0_3462, \16377 );
and \g449003/U$2 ( \18601 , RIfcab488_6971, \16427 );
and \g449003/U$3 ( \18602 , \16448 , RIfc6c9e0_6258);
and \g449003/U$4 ( \18603 , RIfccbb70_7340, \16485 );
nor \g449003/U$1 ( \18604 , \18601 , \18602 , \18603 );
and \g454771/U$2 ( \18605 , \16317 , RIfcabfc8_6979);
and \g454771/U$3 ( \18606 , RIfc6ce18_6261, \16325 );
nor \g454771/U$1 ( \18607 , \18605 , \18606 );
not \g454770/U$1 ( \18608 , \18607 );
and \g450017/U$2 ( \18609 , \18608 , \16336 );
and \g450017/U$3 ( \18610 , RIfcab5f0_6972, \16356 );
nor \g450017/U$1 ( \18611 , \18609 , \18610 );
and \g452250/U$2 ( \18612 , \16361 , RIe1aaf00_3322);
and \g452250/U$3 ( \18613 , RIe1ac580_3338, \16364 );
nor \g452250/U$1 ( \18614 , \18612 , \18613 );
and \g452249/U$2 ( \18615 , \16368 , RIe1b0bd0_3388);
and \g452249/U$3 ( \18616 , RIfea7dc0_8226, \16371 );
nor \g452249/U$1 ( \18617 , \18615 , \18616 );
nand \g448067/U$1 ( \18618 , \18604 , \18611 , \18614 , \18617 );
nor \g446098/U$1 ( \18619 , \18599 , \18600 , \18618 );
and \g452246/U$2 ( \18620 , \16334 , RIe1b3e70_3424);
and \g452246/U$3 ( \18621 , RIe1b9438_3485, \16313 );
nor \g452246/U$1 ( \18622 , \18620 , \18621 );
and \g452243/U$2 ( \18623 , \16380 , RIe1b5220_3438);
and \g452243/U$3 ( \18624 , RIfcdd348_7539, \16319 );
nor \g452243/U$1 ( \18625 , \18623 , \18624 );
and \g445219/U$2 ( \18626 , \18619 , \18622 , \18625 );
nor \g445219/U$1 ( \18627 , \18626 , \16909 );
and \g446101/U$2 ( \18628 , RIe1a8d40_3298, \16328 );
and \g446101/U$3 ( \18629 , RIe21b598_4601, \16334 );
and \g449008/U$2 ( \18630 , RIe1bbd00_3514, \16398 );
and \g449008/U$3 ( \18631 , \16341 , RIe1d5200_3802);
and \g449008/U$4 ( \18632 , RIe179040_2754, \16485 );
nor \g449008/U$1 ( \18633 , \18630 , \18631 , \18632 );
and \g454362/U$2 ( \18634 , \16317 , RIe1fedf8_4277);
and \g454362/U$3 ( \18635 , RIe204d98_4345, \16325 );
nor \g454362/U$1 ( \18636 , \18634 , \18635 );
not \g450020/U$3 ( \18637 , \18636 );
not \g450020/U$4 ( \18638 , \16351 );
and \g450020/U$2 ( \18639 , \18637 , \18638 );
and \g450020/U$5 ( \18640 , \16356 , RIe18cb40_2978);
nor \g450020/U$1 ( \18641 , \18639 , \18640 );
and \g452267/U$2 ( \18642 , \16361 , RIe1711b0_2664);
and \g452267/U$3 ( \18643 , RIe1aeb78_3365, \16364 );
nor \g452267/U$1 ( \18644 , \18642 , \18643 );
and \g452264/U$2 ( \18645 , \16368 , RIe1f0cf8_4117);
and \g452264/U$3 ( \18646 , RIe1f81b0_4200, \16371 );
nor \g452264/U$1 ( \18647 , \18645 , \18646 );
nand \g447734/U$1 ( \18648 , \18633 , \18641 , \18644 , \18647 );
nor \g446101/U$1 ( \18649 , \18628 , \18629 , \18648 );
and \g452260/U$2 ( \18650 , \16377 , RIe1a0640_3202);
and \g452260/U$3 ( \18651 , RIe226998_4729, \16380 );
nor \g452260/U$1 ( \18652 , \18650 , \18651 );
and \g452259/U$2 ( \18653 , \16313 , RIe1a3340_3234);
and \g452259/U$3 ( \18654 , RIe1a6040_3266, \16321 );
nor \g452259/U$1 ( \18655 , \18653 , \18654 );
and \g445223/U$2 ( \18656 , \18649 , \18652 , \18655 );
nor \g445223/U$1 ( \18657 , \18656 , \16586 );
or \g444167/U$1 ( \18658 , \18598 , \18627 , \18657 );
_DC \g378a/U$1 ( \18659 , \18658 , \16652 );
and \g452598/U$2 ( \18660 , \16368 , RIe210030_4472);
and \g452598/U$3 ( \18661 , RIe21e130_4632, \16485 );
nor \g452598/U$1 ( \18662 , \18660 , \18661 );
and \g446172/U$2 ( \18663 , RIfcecc30_7716, \16356 );
and \g446172/U$3 ( \18664 , RIe215a30_4536, \16334 );
and \g449102/U$2 ( \18665 , RIe212d30_4504, \16427 );
and \g449102/U$3 ( \18666 , \16398 , RIe20d330_4440);
and \g449102/U$4 ( \18667 , RIfc545c0_5982, \16339 );
nor \g449102/U$1 ( \18668 , \18665 , \18666 , \18667 );
and \g452605/U$2 ( \18669 , \16361 , RIe207930_4376);
and \g452605/U$3 ( \18670 , RIe20a630_4408, \16364 );
nor \g452605/U$1 ( \18671 , \18669 , \18670 );
and \g452604/U$2 ( \18672 , \16377 , RIe220e30_4664);
and \g452604/U$3 ( \18673 , RIfc82970_6508, \16313 );
nor \g452604/U$1 ( \18674 , \18672 , \18673 );
and \g454931/U$2 ( \18675 , \16317 , RIe223b30_4696);
and \g454931/U$3 ( \18676 , RIfc408e0_5760, \16325 );
nor \g454931/U$1 ( \18677 , \18675 , \18676 );
not \g450117/U$3 ( \18678 , \18677 );
not \g450117/U$4 ( \18679 , \16311 );
and \g450117/U$2 ( \18680 , \18678 , \18679 );
and \g450117/U$5 ( \18681 , \16448 , RIfc3fad0_5750);
nor \g450117/U$1 ( \18682 , \18680 , \18681 );
nand \g447782/U$1 ( \18683 , \18668 , \18671 , \18674 , \18682 );
nor \g446172/U$1 ( \18684 , \18663 , \18664 , \18683 );
and \g452597/U$2 ( \18685 , \16371 , RIf169148_5655);
and \g452597/U$3 ( \18686 , RIe218730_4568, \16380 );
nor \g452597/U$1 ( \18687 , \18685 , \18686 );
nand \g445618/U$1 ( \18688 , \18662 , \18684 , \18687 );
and \g444742/U$2 ( \18689 , \18688 , \16390 );
and \g449098/U$2 ( \18690 , RIfc59480_6038, \16321 );
and \g449098/U$3 ( \18691 , \16344 , RIfc59b88_6043);
and \g449098/U$4 ( \18692 , RIfcdb890_7520, \16356 );
nor \g449098/U$1 ( \18693 , \18690 , \18691 , \18692 );
and \g452589/U$2 ( \18694 , \16368 , RIe173910_2692);
and \g452589/U$3 ( \18695 , RIfc58aa8_6031, \16371 );
nor \g452589/U$1 ( \18696 , \18694 , \18695 );
and \g454981/U$2 ( \18697 , \16317 , RIfc57158_6013);
and \g454981/U$3 ( \18698 , RIfc57c98_6021, \16325 );
nor \g454981/U$1 ( \18699 , \18697 , \18698 );
not \g450113/U$3 ( \18700 , \18699 );
not \g450113/U$4 ( \18701 , \16351 );
and \g450113/U$2 ( \18702 , \18700 , \18701 );
and \g450113/U$5 ( \18703 , \16328 , RIfcbb748_7155);
nor \g450113/U$1 ( \18704 , \18702 , \18703 );
and \g452587/U$2 ( \18705 , \16334 , RIfcb5eb0_7092);
and \g452587/U$3 ( \18706 , RIfc8ada0_6602, \16380 );
nor \g452587/U$1 ( \18707 , \18705 , \18706 );
nand \g447780/U$1 ( \18708 , \18693 , \18696 , \18704 , \18707 );
and \g444742/U$3 ( \18709 , \17998 , \18708 );
nor \g444742/U$1 ( \18710 , \18689 , \18709 );
nor \g448264/U$1 ( \18711 , \16649 , \16517 );
and \g446945/U$2 ( \18712 , \18711 , RIe175c38_2717);
nor \g448271/U$1 ( \18713 , \16649 , \16520 );
and \g446945/U$3 ( \18714 , RIfcbbce8_7159, \18713 );
nor \g446945/U$1 ( \18715 , \18712 , \18714 );
nor \g448265/U$1 ( \18716 , \16649 , \16397 );
and \g446950/U$2 ( \18717 , \18716 , RIfc8a968_6599);
nor \g448267/U$1 ( \18718 , \16649 , \16340 );
and \g446950/U$3 ( \18719 , RIfcc62d8_7277, \18718 );
nor \g446950/U$1 ( \18720 , \18717 , \18719 );
and \g446948/U$2 ( \18721 , \18533 , RIfc56d20_6010);
and \g446948/U$3 ( \18722 , RIfc57428_6015, \18535 );
nor \g446948/U$1 ( \18723 , \18721 , \18722 );
nand \g444623/U$1 ( \18724 , \18710 , \18715 , \18720 , \18723 );
and \g449090/U$2 ( \18725 , RIe186fd8_2913, \16427 );
and \g449090/U$3 ( \18726 , \16448 , RIe189cd8_2945);
and \g449090/U$4 ( \18727 , RIe19aad8_3137, \16321 );
nor \g449090/U$1 ( \18728 , \18725 , \18726 , \18727 );
and \g452562/U$2 ( \18729 , \16368 , RIe1842d8_2881);
and \g452562/U$3 ( \18730 , RIf1438d0_5228, \16371 );
nor \g452562/U$1 ( \18731 , \18729 , \18730 );
and \g454904/U$2 ( \18732 , \16317 , RIe1950d8_3073);
and \g454904/U$3 ( \18733 , RIfc5c5b8_6073, \16325 );
nor \g454904/U$1 ( \18734 , \18732 , \18733 );
not \g450105/U$3 ( \18735 , \18734 );
not \g450105/U$4 ( \18736 , \16330 );
and \g450105/U$2 ( \18737 , \18735 , \18736 );
and \g450105/U$5 ( \18738 , \16326 , RIe19d7d8_3169);
nor \g450105/U$1 ( \18739 , \18737 , \18738 );
and \g452560/U$2 ( \18740 , \16334 , RIe18f6d8_3009);
and \g452560/U$3 ( \18741 , RIe1923d8_3041, \16380 );
nor \g452560/U$1 ( \18742 , \18740 , \18741 );
nand \g447773/U$1 ( \18743 , \18728 , \18731 , \18739 , \18742 );
and \g444709/U$2 ( \18744 , \18743 , \17938 );
and \g446168/U$2 ( \18745 , RIe202638_4317, \16313 );
and \g446168/U$3 ( \18746 , RIfc537b0_5972, \16364 );
and \g449094/U$2 ( \18747 , RIfcba0c8_7139, \16427 );
and \g449094/U$3 ( \18748 , \16432 , RIfcd4270_7436);
and \g449094/U$4 ( \18749 , RIfc4bec0_5886, \16321 );
nor \g449094/U$1 ( \18750 , \18747 , \18748 , \18749 );
and \g452575/U$2 ( \18751 , \16368 , RIe1fbb58_4241);
and \g452575/U$3 ( \18752 , RIe1fcda0_4254, \16371 );
nor \g452575/U$1 ( \18753 , \18751 , \18752 );
and \g454150/U$2 ( \18754 , \16317 , RIfc4c190_5888);
and \g454150/U$3 ( \18755 , RIfc88910_6576, \16325 );
nor \g454150/U$1 ( \18756 , \18754 , \18755 );
not \g450109/U$3 ( \18757 , \18756 );
not \g450109/U$4 ( \18758 , \16330 );
and \g450109/U$2 ( \18759 , \18757 , \18758 );
and \g450109/U$5 ( \18760 , \16326 , RIfc88d48_6579);
nor \g450109/U$1 ( \18761 , \18759 , \18760 );
and \g452573/U$2 ( \18762 , \16334 , RIfcba398_7141);
and \g452573/U$3 ( \18763 , RIfc4c2f8_5889, \16380 );
nor \g452573/U$1 ( \18764 , \18762 , \18763 );
nand \g447776/U$1 ( \18765 , \18750 , \18753 , \18761 , \18764 );
nor \g446168/U$1 ( \18766 , \18745 , \18746 , \18765 );
and \g452567/U$2 ( \18767 , \16341 , RIfc53d50_5976);
and \g452567/U$3 ( \18768 , RIe200b80_4298, \16377 );
nor \g452567/U$1 ( \18769 , \18767 , \18768 );
and \g452568/U$2 ( \18770 , \16361 , RIfc4c5c8_5891);
and \g452568/U$3 ( \18771 , RIfc9b768_6791, \16337 );
nor \g452568/U$1 ( \18772 , \18770 , \18771 );
and \g445270/U$2 ( \18773 , \18766 , \18769 , \18772 );
nor \g445270/U$1 ( \18774 , \18773 , \16393 );
nor \g444709/U$1 ( \18775 , \18744 , \18774 );
nor \g448329/U$1 ( \18776 , \16618 , \16517 );
and \g446936/U$2 ( \18777 , \18776 , RIe197dd8_3105);
nor \g448379/U$1 ( \18778 , \16618 , \16520 );
and \g446936/U$3 ( \18779 , RIfcc2d68_7239, \18778 );
nor \g446936/U$1 ( \18780 , \18777 , \18779 );
nor \g448376/U$1 ( \18781 , \16618 , \16397 );
and \g446937/U$2 ( \18782 , \18781 , RIe1815d8_2849);
nor \g448378/U$1 ( \18783 , \16618 , \16340 );
and \g446937/U$3 ( \18784 , RIfc5b370_6060, \18783 );
nor \g446937/U$1 ( \18785 , \18782 , \18784 );
and \g446938/U$2 ( \18786 , \18467 , RIe17bbd8_2785);
and \g446938/U$3 ( \18787 , RIe17e8d8_2817, \18469 );
nor \g446938/U$1 ( \18788 , \18786 , \18787 );
nand \g444506/U$1 ( \18789 , \18775 , \18780 , \18785 , \18788 );
and \g446156/U$2 ( \18790 , RIf14a7e8_5307, \16356 );
and \g446156/U$3 ( \18791 , RIfe807c0_7806, \16334 );
and \g449082/U$2 ( \18792 , RIf14ba30_5320, \16321 );
and \g449082/U$3 ( \18793 , \16328 , RIf14cc78_5333);
and \g449082/U$4 ( \18794 , RIfce4f08_7627, \16427 );
nor \g449082/U$1 ( \18795 , \18792 , \18793 , \18794 );
and \g452528/U$2 ( \18796 , \16361 , RIfebe728_8287);
and \g452528/U$3 ( \18797 , RIfe80928_7807, \16364 );
nor \g452528/U$1 ( \18798 , \18796 , \18797 );
and \g452526/U$2 ( \18799 , \16377 , RIe1b7278_3461);
and \g452526/U$3 ( \18800 , RIe1b92d0_3484, \16313 );
nor \g452526/U$1 ( \18801 , \18799 , \18800 );
and \g454895/U$2 ( \18802 , \16317 , RIfc87560_6562);
and \g454895/U$3 ( \18803 , RIfc9cde8_6807, \16325 );
nor \g454895/U$1 ( \18804 , \18802 , \18803 );
not \g454894/U$1 ( \18805 , \18804 );
and \g450096/U$2 ( \18806 , \18805 , \16336 );
and \g450096/U$3 ( \18807 , RIfc50510_5936, \16448 );
nor \g450096/U$1 ( \18808 , \18806 , \18807 );
nand \g448075/U$1 ( \18809 , \18795 , \18798 , \18801 , \18808 );
nor \g446156/U$1 ( \18810 , \18790 , \18791 , \18809 );
and \g452523/U$2 ( \18811 , \16371 , RIfe80a90_7808);
and \g452523/U$3 ( \18812 , RIfebe5c0_8286, \16380 );
nor \g452523/U$1 ( \18813 , \18811 , \18812 );
and \g452524/U$2 ( \18814 , \16368 , RIfebe890_8288);
and \g452524/U$3 ( \18815 , RIf149ca8_5299, \16485 );
nor \g452524/U$1 ( \18816 , \18814 , \18815 );
and \g445262/U$2 ( \18817 , \18810 , \18813 , \18816 );
nor \g445262/U$1 ( \18818 , \18817 , \16909 );
and \g446162/U$2 ( \18819 , RIe18c9d8_2977, \16356 );
and \g446162/U$3 ( \18820 , RIe1f0b90_4116, \16368 );
and \g449085/U$2 ( \18821 , RIe1a5ed8_3265, \16321 );
and \g449085/U$3 ( \18822 , \16328 , RIe1a8bd8_3297);
and \g449085/U$4 ( \18823 , RIe1fec90_4276, \16427 );
nor \g449085/U$1 ( \18824 , \18821 , \18822 , \18823 );
and \g452548/U$2 ( \18825 , \16361 , RIe171048_2663);
and \g452548/U$3 ( \18826 , RIe1aea10_3364, \16364 );
nor \g452548/U$1 ( \18827 , \18825 , \18826 );
and \g452545/U$2 ( \18828 , \16377 , RIe1a04d8_3201);
and \g452545/U$3 ( \18829 , RIe1a31d8_3233, \16313 );
nor \g452545/U$1 ( \18830 , \18828 , \18829 );
and \g454180/U$2 ( \18831 , \16317 , RIe1bbb98_3513);
and \g454180/U$3 ( \18832 , RIe1d5098_3801, \16325 );
nor \g454180/U$1 ( \18833 , \18831 , \18832 );
not \g454179/U$1 ( \18834 , \18833 );
and \g450100/U$2 ( \18835 , \18834 , \16336 );
and \g450100/U$3 ( \18836 , RIe204c30_4344, \16448 );
nor \g450100/U$1 ( \18837 , \18835 , \18836 );
nand \g448078/U$1 ( \18838 , \18824 , \18827 , \18830 , \18837 );
nor \g446162/U$1 ( \18839 , \18819 , \18820 , \18838 );
and \g452539/U$2 ( \18840 , \16334 , RIe21b430_4600);
and \g452539/U$3 ( \18841 , RIe1f8048_4199, \16371 );
nor \g452539/U$1 ( \18842 , \18840 , \18841 );
and \g452538/U$2 ( \18843 , \16380 , RIe226830_4728);
and \g452538/U$3 ( \18844 , RIe178ed8_2753, \16485 );
nor \g452538/U$1 ( \18845 , \18843 , \18844 );
and \g445263/U$2 ( \18846 , \18839 , \18842 , \18845 );
nor \g445263/U$1 ( \18847 , \18846 , \16586 );
or \g444318/U$1 ( \18848 , \18724 , \18789 , \18818 , \18847 );
and \g446151/U$2 ( \18849 , RIe1c6f98_3641, \16341 );
and \g446151/U$3 ( \18850 , RIe1e3198_3961, \16377 );
and \g449073/U$2 ( \18851 , RIe1cf698_3737, \16427 );
and \g449073/U$3 ( \18852 , \16432 , RIe1d2398_3769);
and \g449073/U$4 ( \18853 , RIe1e8b98_4025, \16321 );
nor \g449073/U$1 ( \18854 , \18851 , \18852 , \18853 );
and \g452505/U$2 ( \18855 , \16368 , RIe1c9c98_3673);
and \g452505/U$3 ( \18856 , RIe1cc998_3705, \16371 );
nor \g452505/U$1 ( \18857 , \18855 , \18856 );
and \g454880/U$2 ( \18858 , \16317 , RIe1dd798_3897);
and \g454880/U$3 ( \18859 , RIe1e0498_3929, \16325 );
nor \g454880/U$1 ( \18860 , \18858 , \18859 );
not \g450088/U$3 ( \18861 , \18860 );
not \g450088/U$4 ( \18862 , \16330 );
and \g450088/U$2 ( \18863 , \18861 , \18862 );
and \g450088/U$5 ( \18864 , \16328 , RIe1eb898_4057);
nor \g450088/U$1 ( \18865 , \18863 , \18864 );
and \g452503/U$2 ( \18866 , \16334 , RIe1d7d98_3833);
and \g452503/U$3 ( \18867 , RIe1daa98_3865, \16380 );
nor \g452503/U$1 ( \18868 , \18866 , \18867 );
nand \g447765/U$1 ( \18869 , \18854 , \18857 , \18865 , \18868 );
nor \g446151/U$1 ( \18870 , \18849 , \18850 , \18869 );
and \g452495/U$2 ( \18871 , \16361 , RIe1be898_3545);
and \g452495/U$3 ( \18872 , RIe1e5e98_3993, \16313 );
nor \g452495/U$1 ( \18873 , \18871 , \18872 );
and \g452497/U$2 ( \18874 , \16364 , RIe1c1598_3577);
and \g452497/U$3 ( \18875 , RIe1c4298_3609, \16398 );
nor \g452497/U$1 ( \18876 , \18874 , \18875 );
and \g445257/U$2 ( \18877 , \18870 , \18873 , \18876 );
nor \g445257/U$1 ( \18878 , \18877 , \16555 );
and \g446154/U$2 ( \18879 , RIfc849c8_6531, \16356 );
and \g446154/U$3 ( \18880 , RIfebe458_8285, \16368 );
and \g449078/U$2 ( \18881 , RIfcc4988_7259, \16427 );
and \g449078/U$3 ( \18882 , \16398 , RIfcb7f08_7115);
and \g449078/U$4 ( \18883 , RIfc87f38_6569, \16341 );
nor \g449078/U$1 ( \18884 , \18881 , \18882 , \18883 );
and \g452516/U$2 ( \18885 , \16361 , RIfe80658_7805);
and \g452516/U$3 ( \18886 , RIf14e190_5348, \16364 );
nor \g452516/U$1 ( \18887 , \18885 , \18886 );
and \g452512/U$2 ( \18888 , \16377 , RIe1fa208_4223);
and \g452512/U$3 ( \18889 , RIfcb9f60_7138, \16313 );
nor \g452512/U$1 ( \18890 , \18888 , \18889 );
and \g454889/U$2 ( \18891 , \16317 , RIf157da8_5459);
and \g454889/U$3 ( \18892 , RIfc9e468_6823, \16325 );
nor \g454889/U$1 ( \18893 , \18891 , \18892 );
not \g450092/U$3 ( \18894 , \18893 );
not \g450092/U$4 ( \18895 , \16311 );
and \g450092/U$2 ( \18896 , \18894 , \18895 );
and \g450092/U$5 ( \18897 , \16448 , RIf153320_5406);
nor \g450092/U$1 ( \18898 , \18896 , \18897 );
nand \g447766/U$1 ( \18899 , \18884 , \18887 , \18890 , \18898 );
nor \g446154/U$1 ( \18900 , \18879 , \18880 , \18899 );
and \g452511/U$2 ( \18901 , \16334 , RIe1f5618_4169);
and \g452511/U$3 ( \18902 , RIf150d28_5379, \16371 );
nor \g452511/U$1 ( \18903 , \18901 , \18902 );
and \g452510/U$2 ( \18904 , \16380 , RIfc9f6b0_6836);
and \g452510/U$3 ( \18905 , RIfc529a0_5962, \16485 );
nor \g452510/U$1 ( \18906 , \18904 , \18905 );
and \g445259/U$2 ( \18907 , \18900 , \18903 , \18906 );
nor \g445259/U$1 ( \18908 , \18907 , \16480 );
or \g444261/U$1 ( \18909 , \18848 , \18878 , \18908 );
_DC \g380f/U$1 ( \18910 , \18909 , \16652 );
and \g450583/U$2 ( \18911 , \16313 , RIf140360_5190);
and \g450583/U$3 ( \18912 , RIf140ea0_5198, \16321 );
nor \g450583/U$1 ( \18913 , \18911 , \18912 );
and \g445709/U$2 ( \18914 , RIf1423b8_5213, \16326 );
and \g445709/U$3 ( \18915 , RIee3d4c8_5156, \16334 );
and \g448507/U$2 ( \18916 , RIfe7af28_7743, \16427 );
and \g448507/U$3 ( \18917 , \16432 , RIfe7b090_7744);
and \g448507/U$4 ( \18918 , RIf13f280_5178, \16485 );
nor \g448507/U$1 ( \18919 , \18916 , \18917 , \18918 );
and \g454614/U$2 ( \18920 , \16317 , RIfe7ac58_7741);
and \g454614/U$3 ( \18921 , RIfe7adc0_7742, \16325 );
nor \g454614/U$1 ( \18922 , \18920 , \18921 );
not \g454613/U$1 ( \18923 , \18922 );
and \g449528/U$2 ( \18924 , \18923 , \16336 );
and \g449528/U$3 ( \18925 , RIf13fc58_5185, \16356 );
nor \g449528/U$1 ( \18926 , \18924 , \18925 );
and \g450600/U$2 ( \18927 , \16361 , RIfcb20d0_7048);
and \g450600/U$3 ( \18928 , RIf16e440_5714, \16364 );
nor \g450600/U$1 ( \18929 , \18927 , \18928 );
and \g450596/U$2 ( \18930 , \16368 , RIe1737a8_2691);
and \g450596/U$3 ( \18931 , RIee39df0_5117, \16371 );
nor \g450596/U$1 ( \18932 , \18930 , \18931 );
nand \g448005/U$1 ( \18933 , \18919 , \18926 , \18929 , \18932 );
nor \g445709/U$1 ( \18934 , \18914 , \18915 , \18933 );
and \g450586/U$2 ( \18935 , \16377 , RIfe7b798_7749);
and \g450586/U$3 ( \18936 , RIfc79460_6402, \16380 );
nor \g450586/U$1 ( \18937 , \18935 , \18936 );
nand \g445508/U$1 ( \18938 , \18913 , \18934 , \18937 );
and \g444749/U$2 ( \18939 , \18938 , \17998 );
and \g448499/U$2 ( \18940 , RIe186e70_2912, \16427 );
and \g448499/U$3 ( \18941 , \16448 , RIe189b70_2944);
and \g448499/U$4 ( \18942 , RIe194f70_3072, \16344 );
nor \g448499/U$1 ( \18943 , \18940 , \18941 , \18942 );
and \g454525/U$2 ( \18944 , \16317 , RIe181470_2848);
and \g454525/U$3 ( \18945 , RIfe7b1f8_7745, \16325 );
nor \g454525/U$1 ( \18946 , \18944 , \18945 );
not \g454524/U$1 ( \18947 , \18946 );
and \g449519/U$2 ( \18948 , \18947 , \16336 );
and \g449519/U$3 ( \18949 , RIfe7b4c8_7747, \16356 );
nor \g449519/U$1 ( \18950 , \18948 , \18949 );
and \g450566/U$2 ( \18951 , \16361 , RIe17ba70_2784);
and \g450566/U$3 ( \18952 , RIe17e770_2816, \16364 );
nor \g450566/U$1 ( \18953 , \18951 , \18952 );
and \g450563/U$2 ( \18954 , \16368 , RIe184170_2880);
and \g450563/U$3 ( \18955 , RIfe7b360_7746, \16371 );
nor \g450563/U$1 ( \18956 , \18954 , \18955 );
nand \g448004/U$1 ( \18957 , \18943 , \18950 , \18953 , \18956 );
and \g444749/U$3 ( \18958 , \17938 , \18957 );
nor \g444749/U$1 ( \18959 , \18939 , \18958 );
nor \g448328/U$1 ( \18960 , \16618 , \16510 );
and \g446505/U$2 ( \18961 , \18960 , RIe18f570_3008);
nor \g448394/U$1 ( \18962 , \16618 , \16513 );
and \g446505/U$3 ( \18963 , RIe192270_3040, \18962 );
nor \g446505/U$1 ( \18964 , \18961 , \18963 );
nor \g448392/U$1 ( \18965 , \16618 , \16320 );
and \g446503/U$2 ( \18966 , \18965 , RIe19a970_3136);
nor \g448393/U$1 ( \18967 , \16618 , \16327 );
and \g446503/U$3 ( \18968 , RIe19d670_3168, \18967 );
nor \g446503/U$1 ( \18969 , \18966 , \18968 );
and \g446506/U$2 ( \18970 , \18776 , RIe197c70_3104);
and \g446506/U$3 ( \18971 , RIfe7b630_7748, \18778 );
nor \g446506/U$1 ( \18972 , \18970 , \18971 );
nand \g444444/U$1 ( \18973 , \18959 , \18964 , \18969 , \18972 );
and \g450648/U$2 ( \18974 , \16371 , RIf150bc0_5378);
and \g450648/U$3 ( \18975 , RIf151b38_5389, \16427 );
nor \g450648/U$1 ( \18976 , \18974 , \18975 );
and \g445723/U$2 ( \18977 , RIfe7c008_7755, \16448 );
and \g445723/U$3 ( \18978 , RIe1edff8_4085, \16361 );
and \g448526/U$2 ( \18979 , RIf157c40_5458, \16319 );
and \g448526/U$3 ( \18980 , \16328 , RIf158ff0_5472);
and \g448526/U$4 ( \18981 , RIf14ee38_5357, \16398 );
nor \g448526/U$1 ( \18982 , \18979 , \18980 , \18981 );
and \g454278/U$2 ( \18983 , \16317 , RIf155918_5433);
and \g454278/U$3 ( \18984 , RIf156458_5441, \16325 );
nor \g454278/U$1 ( \18985 , \18983 , \18984 );
not \g449546/U$3 ( \18986 , \18985 );
not \g449546/U$4 ( \18987 , \16330 );
and \g449546/U$2 ( \18988 , \18986 , \18987 );
and \g449546/U$5 ( \18989 , \16341 , RIf14fae0_5366);
nor \g449546/U$1 ( \18990 , \18988 , \18989 );
and \g450661/U$2 ( \18991 , \16377 , RIfe7c170_7756);
and \g450661/U$3 ( \18992 , RIf156f98_5449, \16313 );
nor \g450661/U$1 ( \18993 , \18991 , \18992 );
and \g450664/U$2 ( \18994 , \16334 , RIe1f54b0_4168);
and \g450664/U$3 ( \18995 , RIf1549a0_5422, \16380 );
nor \g450664/U$1 ( \18996 , \18994 , \18995 );
nand \g447238/U$1 ( \18997 , \18982 , \18990 , \18993 , \18996 );
nor \g445723/U$1 ( \18998 , \18977 , \18978 , \18997 );
and \g450651/U$2 ( \18999 , \16364 , RIf14e028_5347);
and \g450651/U$3 ( \19000 , RIe1f32f0_4144, \16368 );
nor \g450651/U$1 ( \19001 , \18999 , \19000 );
nand \g445511/U$1 ( \19002 , \18976 , \18998 , \19001 );
and \g444830/U$2 ( \19003 , \19002 , \16481 );
and \g448516/U$2 ( \19004 , RIf147db8_5277, \16427 );
and \g448516/U$3 ( \19005 , \16448 , RIf149000_5290);
and \g448516/U$4 ( \19006 , RIfe7c2d8_7757, \16485 );
nor \g448516/U$1 ( \19007 , \19004 , \19005 , \19006 );
and \g454437/U$2 ( \19008 , \16317 , RIf146738_5261);
and \g454437/U$3 ( \19009 , RIfe7c5a8_7759, \16325 );
nor \g454437/U$1 ( \19010 , \19008 , \19009 );
not \g454436/U$1 ( \19011 , \19010 );
and \g449537/U$2 ( \19012 , \19011 , \16336 );
and \g449537/U$3 ( \19013 , RIf14a680_5306, \16356 );
nor \g449537/U$1 ( \19014 , \19012 , \19013 );
and \g450631/U$2 ( \19015 , \16361 , RIe1aad98_3321);
and \g450631/U$3 ( \19016 , RIfe7c710_7760, \16364 );
nor \g450631/U$1 ( \19017 , \19015 , \19016 );
and \g450626/U$2 ( \19018 , \16368 , RIfebd918_8277);
and \g450626/U$3 ( \19019 , RIe1b2688_3407, \16371 );
nor \g450626/U$1 ( \19020 , \19018 , \19019 );
nand \g448006/U$1 ( \19021 , \19007 , \19014 , \19017 , \19020 );
and \g444830/U$3 ( \19022 , \16477 , \19021 );
nor \g444830/U$1 ( \19023 , \19003 , \19022 );
and \g446520/U$2 ( \19024 , \18268 , RIf14b8c8_5319);
and \g446520/U$3 ( \19025 , RIf14cb10_5332, \18270 );
nor \g446520/U$1 ( \19026 , \19024 , \19025 );
and \g446521/U$2 ( \19027 , \18273 , RIfe7c878_7761);
and \g446521/U$3 ( \19028 , RIfebda80_8278, \18275 );
nor \g446521/U$1 ( \19029 , \19027 , \19028 );
and \g446522/U$2 ( \19030 , \18278 , RIfe7c440_7758);
and \g446522/U$3 ( \19031 , RIfe7c9e0_7762, \18280 );
nor \g446522/U$1 ( \19032 , \19030 , \19031 );
nand \g444551/U$1 ( \19033 , \19023 , \19026 , \19029 , \19032 );
and \g446488/U$2 ( \19034 , RIe2239c8_4695, \16321 );
and \g446488/U$3 ( \19035 , RIf16be48_5687, \16313 );
and \g449505/U$2 ( \19036 , RIe20d1c8_4439, \16398 );
and \g449505/U$3 ( \19037 , \16341 , RIfe7b900_7750);
and \g449505/U$4 ( \19038 , RIe21dfc8_4631, \16344 );
nor \g449505/U$1 ( \19039 , \19036 , \19037 , \19038 );
and \g455020/U$2 ( \19040 , \16317 , RIe212bc8_4503);
and \g455020/U$3 ( \19041 , RIfebd7b0_8276, \16325 );
nor \g455020/U$1 ( \19042 , \19040 , \19041 );
not \g450524/U$3 ( \19043 , \19042 );
not \g450524/U$4 ( \19044 , \16351 );
and \g450524/U$2 ( \19045 , \19043 , \19044 );
and \g450524/U$5 ( \19046 , \16356 , RIf16aed0_5676);
nor \g450524/U$1 ( \19047 , \19045 , \19046 );
and \g454088/U$2 ( \19048 , \16361 , RIe2077c8_4375);
and \g454088/U$3 ( \19049 , RIe20a4c8_4407, \16364 );
nor \g454088/U$1 ( \19050 , \19048 , \19049 );
and \g454085/U$2 ( \19051 , \16368 , RIe20fec8_4471);
and \g454085/U$3 ( \19052 , RIfebd648_8275, \16371 );
nor \g454085/U$1 ( \19053 , \19051 , \19052 );
nand \g447999/U$1 ( \19054 , \19039 , \19047 , \19050 , \19053 );
nor \g446488/U$1 ( \19055 , \19034 , \19035 , \19054 );
and \g454075/U$2 ( \19056 , \16377 , RIe220cc8_4663);
and \g454075/U$3 ( \19057 , RIe2185c8_4567, \16380 );
nor \g454075/U$1 ( \19058 , \19056 , \19057 );
and \g454073/U$2 ( \19059 , \16334 , RIe2158c8_4535);
and \g454073/U$3 ( \19060 , RIfe7bd38_7753, \16328 );
nor \g454073/U$1 ( \19061 , \19059 , \19060 );
and \g445492/U$2 ( \19062 , \19055 , \19058 , \19061 );
nor \g445492/U$1 ( \19063 , \19062 , \16389 );
and \g446494/U$2 ( \19064 , RIf166178_5621, \16319 );
and \g446494/U$3 ( \19065 , RIe2024d0_4316, \16313 );
and \g448491/U$2 ( \19066 , RIf15b8b8_5501, \16398 );
and \g448491/U$3 ( \19067 , \16341 , RIf15cdd0_5516);
and \g448491/U$4 ( \19068 , RIf1646c0_5602, \16485 );
nor \g448491/U$1 ( \19069 , \19066 , \19067 , \19068 );
and \g454813/U$2 ( \19070 , \16317 , RIf15e2e8_5531);
and \g454813/U$3 ( \19071 , RIf1601d8_5553, \16325 );
nor \g454813/U$1 ( \19072 , \19070 , \19071 );
not \g450534/U$3 ( \19073 , \19072 );
not \g450534/U$4 ( \19074 , \16351 );
and \g450534/U$2 ( \19075 , \19073 , \19074 );
and \g450534/U$5 ( \19076 , \16356 , RIf165368_5611);
nor \g450534/U$1 ( \19077 , \19075 , \19076 );
and \g454121/U$2 ( \19078 , \16361 , RIfca4840_6894);
and \g454121/U$3 ( \19079 , RIf15a7d8_5489, \16364 );
nor \g454121/U$1 ( \19080 , \19078 , \19079 );
and \g454118/U$2 ( \19081 , \16368 , RIfe7bea0_7754);
and \g454118/U$3 ( \19082 , RIfe7ba68_7751, \16371 );
nor \g454118/U$1 ( \19083 , \19081 , \19082 );
nand \g448001/U$1 ( \19084 , \19069 , \19077 , \19080 , \19083 );
nor \g446494/U$1 ( \19085 , \19064 , \19065 , \19084 );
and \g454109/U$2 ( \19086 , \16377 , RIfe7bbd0_7752);
and \g454109/U$3 ( \19087 , RIfcd0a30_7396, \16380 );
nor \g454109/U$1 ( \19088 , \19086 , \19087 );
and \g454106/U$2 ( \19089 , \16334 , RIf1620c8_5575);
and \g454106/U$3 ( \19090 , RIf167258_5633, \16326 );
nor \g454106/U$1 ( \19091 , \19089 , \19090 );
and \g445496/U$2 ( \19092 , \19085 , \19088 , \19091 );
nor \g445496/U$1 ( \19093 , \19092 , \16393 );
or \g444348/U$1 ( \19094 , \18973 , \19033 , \19063 , \19093 );
and \g446471/U$2 ( \19095 , RIe204ac8_4343, \16432 );
and \g446471/U$3 ( \19096 , RIe170ee0_2662, \16361 );
and \g449487/U$2 ( \19097 , RIe1a5d70_3264, \16321 );
and \g449487/U$3 ( \19098 , \16328 , RIe1a8a70_3296);
and \g449487/U$4 ( \19099 , RIe1bba30_3512, \16398 );
nor \g449487/U$1 ( \19100 , \19097 , \19098 , \19099 );
and \g455393/U$2 ( \19101 , \16317 , RIe178d70_2752);
and \g455393/U$3 ( \19102 , RIe18c870_2976, \16325 );
nor \g455393/U$1 ( \19103 , \19101 , \19102 );
not \g450507/U$3 ( \19104 , \19103 );
not \g450507/U$4 ( \19105 , \16330 );
and \g450507/U$2 ( \19106 , \19104 , \19105 );
and \g450507/U$5 ( \19107 , \16341 , RIe1d4f30_3800);
nor \g450507/U$1 ( \19108 , \19106 , \19107 );
and \g454018/U$2 ( \19109 , \16377 , RIe1a0370_3200);
and \g454018/U$3 ( \19110 , RIe1a3070_3232, \16313 );
nor \g454018/U$1 ( \19111 , \19109 , \19110 );
and \g454020/U$2 ( \19112 , \16334 , RIe21b2c8_4599);
and \g454020/U$3 ( \19113 , RIe2266c8_4727, \16380 );
nor \g454020/U$1 ( \19114 , \19112 , \19113 );
nand \g447444/U$1 ( \19115 , \19100 , \19108 , \19111 , \19114 );
nor \g446471/U$1 ( \19116 , \19095 , \19096 , \19115 );
and \g454007/U$2 ( \19117 , \16364 , RIe1ae8a8_3363);
and \g454007/U$3 ( \19118 , RIe1f0a28_4115, \16368 );
nor \g454007/U$1 ( \19119 , \19117 , \19118 );
and \g453884/U$2 ( \19120 , \16371 , RIe1f7ee0_4198);
and \g453884/U$3 ( \19121 , RIe1feb28_4275, \16427 );
nor \g453884/U$1 ( \19122 , \19120 , \19121 );
and \g445477/U$2 ( \19123 , \19116 , \19119 , \19122 );
nor \g445477/U$1 ( \19124 , \19123 , \16586 );
and \g446481/U$2 ( \19125 , RIe1d2230_3768, \16448 );
and \g446481/U$3 ( \19126 , RIe1be730_3544, \16361 );
and \g449494/U$2 ( \19127 , RIe1dd630_3896, \16485 );
and \g449494/U$3 ( \19128 , \16356 , RIe1e0330_3928);
and \g449494/U$4 ( \19129 , RIe1c4130_3608, \16398 );
nor \g449494/U$1 ( \19130 , \19127 , \19128 , \19129 );
and \g454602/U$2 ( \19131 , \16317 , RIe1e8a30_4024);
and \g454602/U$3 ( \19132 , RIe1eb730_4056, \16325 );
nor \g454602/U$1 ( \19133 , \19131 , \19132 );
not \g450516/U$3 ( \19134 , \19133 );
not \g450516/U$4 ( \19135 , \16311 );
and \g450516/U$2 ( \19136 , \19134 , \19135 );
and \g450516/U$5 ( \19137 , \16339 , RIe1c6e30_3640);
nor \g450516/U$1 ( \19138 , \19136 , \19137 );
and \g454052/U$2 ( \19139 , \16377 , RIe1e3030_3960);
and \g454052/U$3 ( \19140 , RIe1e5d30_3992, \16313 );
nor \g454052/U$1 ( \19141 , \19139 , \19140 );
and \g454058/U$2 ( \19142 , \16334 , RIe1d7c30_3832);
and \g454058/U$3 ( \19143 , RIe1da930_3864, \16380 );
nor \g454058/U$1 ( \19144 , \19142 , \19143 );
nand \g447447/U$1 ( \19145 , \19130 , \19138 , \19141 , \19144 );
nor \g446481/U$1 ( \19146 , \19125 , \19126 , \19145 );
and \g454043/U$2 ( \19147 , \16364 , RIe1c1430_3576);
and \g454043/U$3 ( \19148 , RIe1c9b30_3672, \16368 );
nor \g454043/U$1 ( \19149 , \19147 , \19148 );
and \g454038/U$2 ( \19150 , \16371 , RIe1cc830_3704);
and \g454038/U$3 ( \19151 , RIe1cf530_3736, \16427 );
nor \g454038/U$1 ( \19152 , \19150 , \19151 );
and \g445485/U$2 ( \19153 , \19146 , \19149 , \19152 );
nor \g445485/U$1 ( \19154 , \19153 , \16555 );
or \g444231/U$1 ( \19155 , \19094 , \19124 , \19154 );
_DC \g3894/U$1 ( \19156 , \19155 , \16652 );
and \g451170/U$2 ( \19157 , \16361 , RIe170d78_2661);
and \g451170/U$3 ( \19158 , RIe1fe9c0_4274, \16427 );
nor \g451170/U$1 ( \19159 , \19157 , \19158 );
and \g445837/U$2 ( \19160 , RIe204960_4342, \16448 );
and \g445837/U$3 ( \19161 , RIe1f7d78_4197, \16371 );
and \g448671/U$2 ( \19162 , RIe178c08_2751, \16485 );
and \g448671/U$3 ( \19163 , \16356 , RIe18c708_2975);
and \g448671/U$4 ( \19164 , RIe1bb8c8_3511, \16337 );
nor \g448671/U$1 ( \19165 , \19162 , \19163 , \19164 );
and \g454704/U$2 ( \19166 , \16317 , RIe1a5c08_3263);
and \g454704/U$3 ( \19167 , RIe1a8908_3295, \16325 );
nor \g454704/U$1 ( \19168 , \19166 , \19167 );
not \g449696/U$3 ( \19169 , \19168 );
not \g449696/U$4 ( \19170 , \16311 );
and \g449696/U$2 ( \19171 , \19169 , \19170 );
and \g449696/U$5 ( \19172 , \16339 , RIe1d4dc8_3799);
nor \g449696/U$1 ( \19173 , \19171 , \19172 );
and \g451182/U$2 ( \19174 , \16377 , RIe1a0208_3199);
and \g451182/U$3 ( \19175 , RIe1a2f08_3231, \16313 );
nor \g451182/U$1 ( \19176 , \19174 , \19175 );
and \g451185/U$2 ( \19177 , \16334 , RIe21b160_4598);
and \g451185/U$3 ( \19178 , RIe226560_4726, \16380 );
nor \g451185/U$1 ( \19179 , \19177 , \19178 );
nand \g447266/U$1 ( \19180 , \19165 , \19173 , \19176 , \19179 );
nor \g445837/U$1 ( \19181 , \19160 , \19161 , \19180 );
and \g451168/U$2 ( \19182 , \16364 , RIe1ae740_3362);
and \g451168/U$3 ( \19183 , RIe1f08c0_4114, \16368 );
nor \g451168/U$1 ( \19184 , \19182 , \19183 );
nand \g445536/U$1 ( \19185 , \19159 , \19181 , \19184 );
and \g444759/U$2 ( \19186 , \19185 , \16752 );
and \g448660/U$2 ( \19187 , RIe1e88c8_4023, \16321 );
and \g448660/U$3 ( \19188 , \16328 , RIe1eb5c8_4055);
and \g448660/U$4 ( \19189 , RIe1c3fc8_3607, \16337 );
nor \g448660/U$1 ( \19190 , \19187 , \19188 , \19189 );
and \g454196/U$2 ( \19191 , \16317 , RIe1dd4c8_3895);
and \g454196/U$3 ( \19192 , RIe1e01c8_3927, \16325 );
nor \g454196/U$1 ( \19193 , \19191 , \19192 );
not \g449685/U$3 ( \19194 , \19193 );
not \g449685/U$4 ( \19195 , \16330 );
and \g449685/U$2 ( \19196 , \19194 , \19195 );
and \g449685/U$5 ( \19197 , \16339 , RIe1c6cc8_3639);
nor \g449685/U$1 ( \19198 , \19196 , \19197 );
and \g451147/U$2 ( \19199 , \16377 , RIe1e2ec8_3959);
and \g451147/U$3 ( \19200 , RIe1e5bc8_3991, \16313 );
nor \g451147/U$1 ( \19201 , \19199 , \19200 );
and \g451150/U$2 ( \19202 , \16334 , RIe1d7ac8_3831);
and \g451150/U$3 ( \19203 , RIe1da7c8_3863, \16380 );
nor \g451150/U$1 ( \19204 , \19202 , \19203 );
nand \g447263/U$1 ( \19205 , \19190 , \19198 , \19201 , \19204 );
and \g444759/U$3 ( \19206 , \16750 , \19205 );
nor \g444759/U$1 ( \19207 , \19186 , \19206 );
nor \g448322/U$1 ( \19208 , \16555 , \16418 );
and \g446619/U$2 ( \19209 , \19208 , RIe1be5c8_3543);
nor \g448370/U$1 ( \19210 , \16555 , \16440 );
and \g446619/U$3 ( \19211 , RIe1cc6c8_3703, \19210 );
nor \g446619/U$1 ( \19212 , \19209 , \19211 );
nor \g448342/U$1 ( \19213 , \16555 , \16421 );
and \g446623/U$2 ( \19214 , \19213 , RIe1c12c8_3575);
nor \g448323/U$1 ( \19215 , \16555 , \16437 );
and \g446623/U$3 ( \19216 , RIe1c99c8_3671, \19215 );
nor \g446623/U$1 ( \19217 , \19214 , \19216 );
nor \g448358/U$1 ( \19218 , \16555 , \16428 );
and \g446617/U$2 ( \19219 , \19218 , RIe1cf3c8_3735);
nor \g448357/U$1 ( \19220 , \16555 , \16433 );
and \g446617/U$3 ( \19221 , RIe1d20c8_3767, \19220 );
nor \g446617/U$1 ( \19222 , \19219 , \19221 );
nand \g444567/U$1 ( \19223 , \19207 , \19212 , \19217 , \19222 );
and \g451102/U$2 ( \19224 , \16377 , RIfe7e768_7783);
and \g451102/U$3 ( \19225 , RIf154838_5421, \16380 );
nor \g451102/U$1 ( \19226 , \19224 , \19225 );
and \g445821/U$2 ( \19227 , RIf157ad8_5457, \16321 );
and \g445821/U$3 ( \19228 , RIf156e30_5448, \16313 );
and \g448651/U$2 ( \19229 , RIfc52400_5958, \16427 );
and \g448651/U$3 ( \19230 , \16448 , RIf1531b8_5405);
and \g448651/U$4 ( \19231 , RIf1557b0_5432, \16485 );
nor \g448651/U$1 ( \19232 , \19229 , \19230 , \19231 );
and \g454281/U$2 ( \19233 , \16317 , RIf14ecd0_5356);
and \g454281/U$3 ( \19234 , RIf14f978_5365, \16325 );
nor \g454281/U$1 ( \19235 , \19233 , \19234 );
not \g454280/U$1 ( \19236 , \19235 );
and \g449675/U$2 ( \19237 , \19236 , \16336 );
and \g449675/U$3 ( \19238 , RIf1562f0_5440, \16354 );
nor \g449675/U$1 ( \19239 , \19237 , \19238 );
and \g451112/U$2 ( \19240 , \16361 , RIe1ede90_4084);
and \g451112/U$3 ( \19241 , RIf14dec0_5346, \16364 );
nor \g451112/U$1 ( \19242 , \19240 , \19241 );
and \g451109/U$2 ( \19243 , \16368 , RIe1f3188_4143);
and \g451109/U$3 ( \19244 , RIf150a58_5377, \16371 );
nor \g451109/U$1 ( \19245 , \19243 , \19244 );
nand \g448022/U$1 ( \19246 , \19232 , \19239 , \19242 , \19245 );
nor \g445821/U$1 ( \19247 , \19227 , \19228 , \19246 );
and \g451098/U$2 ( \19248 , \16334 , RIfe7e8d0_7784);
and \g451098/U$3 ( \19249 , RIf158e88_5471, \16326 );
nor \g451098/U$1 ( \19250 , \19248 , \19249 );
nand \g445533/U$1 ( \19251 , \19226 , \19247 , \19250 );
and \g444832/U$2 ( \19252 , \19251 , \16481 );
and \g448642/U$2 ( \19253 , RIfca1f78_6865, \16485 );
and \g448642/U$3 ( \19254 , \16354 , RIf14a518_5305);
and \g448642/U$4 ( \19255 , RIf1465d0_5260, \16398 );
nor \g448642/U$1 ( \19256 , \19253 , \19254 , \19255 );
and \g455190/U$2 ( \19257 , \16317 , RIf14b760_5318);
and \g455190/U$3 ( \19258 , RIf14c9a8_5331, \16325 );
nor \g455190/U$1 ( \19259 , \19257 , \19258 );
not \g449667/U$3 ( \19260 , \19259 );
not \g449667/U$4 ( \19261 , \16311 );
and \g449667/U$2 ( \19262 , \19260 , \19261 );
and \g449667/U$5 ( \19263 , \16339 , RIf147278_5269);
nor \g449667/U$1 ( \19264 , \19262 , \19263 );
and \g451083/U$2 ( \19265 , \16377 , RIfe7e600_7782);
and \g451083/U$3 ( \19266 , RIfe7ed08_7787, \16313 );
nor \g451083/U$1 ( \19267 , \19265 , \19266 );
and \g451086/U$2 ( \19268 , \16334 , RIfe7e498_7781);
and \g451086/U$3 ( \19269 , RIfe7eba0_7786, \16380 );
nor \g451086/U$1 ( \19270 , \19268 , \19269 );
nand \g447262/U$1 ( \19271 , \19256 , \19264 , \19267 , \19270 );
and \g444832/U$3 ( \19272 , \16477 , \19271 );
nor \g444832/U$1 ( \19273 , \19252 , \19272 );
and \g446604/U$2 ( \19274 , \17463 , RIe1aac30_3320);
and \g446604/U$3 ( \19275 , RIf147c50_5276, \17465 );
nor \g446604/U$1 ( \19276 , \19274 , \19275 );
and \g446603/U$2 ( \19277 , \17468 , RIe1ac418_3337);
and \g446603/U$3 ( \19278 , RIf148e98_5289, \17470 );
nor \g446603/U$1 ( \19279 , \19277 , \19278 );
and \g446607/U$2 ( \19280 , \17473 , RIe1b0a68_3387);
and \g446607/U$3 ( \19281 , RIfe7e330_7780, \17475 );
nor \g446607/U$1 ( \19282 , \19280 , \19281 );
nand \g444565/U$1 ( \19283 , \19273 , \19276 , \19279 , \19282 );
and \g445800/U$2 ( \19284 , RIe186d08_2911, \16427 );
and \g445800/U$3 ( \19285 , RIe184008_2879, \16368 );
and \g448625/U$2 ( \19286 , RIe194e08_3071, \16485 );
and \g448625/U$3 ( \19287 , \16356 , RIfe7efd8_7789);
and \g448625/U$4 ( \19288 , RIe181308_2847, \16337 );
nor \g448625/U$1 ( \19289 , \19286 , \19287 , \19288 );
and \g454580/U$2 ( \19290 , \16317 , RIe19a808_3135);
and \g454580/U$3 ( \19291 , RIe19d508_3167, \16325 );
nor \g454580/U$1 ( \19292 , \19290 , \19291 );
not \g449650/U$3 ( \19293 , \19292 );
not \g449650/U$4 ( \19294 , \16311 );
and \g449650/U$2 ( \19295 , \19293 , \19294 );
and \g449650/U$5 ( \19296 , \16341 , RIfc4bbf0_5884);
nor \g449650/U$1 ( \19297 , \19295 , \19296 );
and \g451021/U$2 ( \19298 , \16377 , RIe197b08_3103);
and \g451021/U$3 ( \19299 , RIfe7ee70_7788, \16313 );
nor \g451021/U$1 ( \19300 , \19298 , \19299 );
and \g451024/U$2 ( \19301 , \16334 , RIe18f408_3007);
and \g451024/U$3 ( \19302 , RIe192108_3039, \16380 );
nor \g451024/U$1 ( \19303 , \19301 , \19302 );
nand \g447260/U$1 ( \19304 , \19289 , \19297 , \19300 , \19303 );
nor \g445800/U$1 ( \19305 , \19284 , \19285 , \19304 );
and \g451012/U$2 ( \19306 , \16361 , RIe17b908_2783);
and \g451012/U$3 ( \19307 , RIe189a08_2943, \16448 );
nor \g451012/U$1 ( \19308 , \19306 , \19307 );
and \g451007/U$2 ( \19309 , \16364 , RIe17e608_2815);
and \g451007/U$3 ( \19310 , RIf143768_5227, \16371 );
nor \g451007/U$1 ( \19311 , \19309 , \19310 );
and \g444999/U$2 ( \19312 , \19305 , \19308 , \19311 );
nor \g444999/U$1 ( \19313 , \19312 , \16618 );
and \g445806/U$2 ( \19314 , RIee3c280_5143, \16448 );
and \g445806/U$3 ( \19315 , RIfe7f140_7790, \16371 );
and \g448633/U$2 ( \19316 , RIf13f118_5177, \16485 );
and \g448633/U$3 ( \19317 , \16356 , RIfe7f2a8_7791);
and \g448633/U$4 ( \19318 , RIf16f520_5726, \16398 );
nor \g448633/U$1 ( \19319 , \19316 , \19317 , \19318 );
and \g454193/U$2 ( \19320 , \16317 , RIf140d38_5197);
and \g454193/U$3 ( \19321 , RIfe7f410_7792, \16325 );
nor \g454193/U$1 ( \19322 , \19320 , \19321 );
not \g449659/U$3 ( \19323 , \19322 );
not \g449659/U$4 ( \19324 , \16311 );
and \g449659/U$2 ( \19325 , \19323 , \19324 );
and \g449659/U$5 ( \19326 , \16341 , RIf170330_5736);
nor \g449659/U$1 ( \19327 , \19325 , \19326 );
and \g451049/U$2 ( \19328 , \16377 , RIe175ad0_2716);
and \g451049/U$3 ( \19329 , RIe176fe8_2731, \16313 );
nor \g451049/U$1 ( \19330 , \19328 , \19329 );
and \g451054/U$2 ( \19331 , \16334 , RIee3d360_5155);
and \g451054/U$3 ( \19332 , RIee3e440_5167, \16380 );
nor \g451054/U$1 ( \19333 , \19331 , \19332 );
nand \g447261/U$1 ( \19334 , \19319 , \19327 , \19330 , \19333 );
nor \g445806/U$1 ( \19335 , \19314 , \19315 , \19334 );
and \g451038/U$2 ( \19336 , \16364 , RIf16e2d8_5713);
and \g451038/U$3 ( \19337 , RIe173640_2690, \16368 );
nor \g451038/U$1 ( \19338 , \19336 , \19337 );
and \g451043/U$2 ( \19339 , \16361 , RIf16d630_5704);
and \g451043/U$3 ( \19340 , RIee3b1a0_5131, \16427 );
nor \g451043/U$1 ( \19341 , \19339 , \19340 );
and \g445003/U$2 ( \19342 , \19335 , \19338 , \19341 );
nor \g445003/U$1 ( \19343 , \19342 , \16649 );
or \g444385/U$1 ( \19344 , \19223 , \19283 , \19313 , \19343 );
and \g445788/U$2 ( \19345 , RIe223860_4694, \16321 );
and \g445788/U$3 ( \19346 , RIfc9c410_6800, \16313 );
and \g448608/U$2 ( \19347 , RIe20d060_4438, \16398 );
and \g448608/U$3 ( \19348 , \16339 , RIfc873f8_6561);
and \g448608/U$4 ( \19349 , RIe21de60_4630, \16485 );
nor \g448608/U$1 ( \19350 , \19347 , \19348 , \19349 );
and \g455168/U$2 ( \19351 , \16317 , RIe212a60_4502);
and \g455168/U$3 ( \19352 , RIfc9cc80_6806, \16325 );
nor \g455168/U$1 ( \19353 , \19351 , \19352 );
not \g449635/U$3 ( \19354 , \19353 );
not \g449635/U$4 ( \19355 , \16351 );
and \g449635/U$2 ( \19356 , \19354 , \19355 );
and \g449635/U$5 ( \19357 , \16356 , RIfcb8340_7118);
nor \g449635/U$1 ( \19358 , \19356 , \19357 );
and \g450963/U$2 ( \19359 , \16361 , RIe207660_4374);
and \g450963/U$3 ( \19360 , RIe20a360_4406, \16364 );
nor \g450963/U$1 ( \19361 , \19359 , \19360 );
and \g450958/U$2 ( \19362 , \16368 , RIe20fd60_4470);
and \g450958/U$3 ( \19363 , RIfc4ddb0_5908, \16371 );
nor \g450958/U$1 ( \19364 , \19362 , \19363 );
nand \g447513/U$1 ( \19365 , \19350 , \19358 , \19361 , \19364 );
nor \g445788/U$1 ( \19366 , \19345 , \19346 , \19365 );
and \g450949/U$2 ( \19367 , \16377 , RIe220b60_4662);
and \g450949/U$3 ( \19368 , RIe218460_4566, \16380 );
nor \g450949/U$1 ( \19369 , \19367 , \19368 );
and \g450946/U$2 ( \19370 , \16334 , RIe215760_4534);
and \g450946/U$3 ( \19371 , RIfe7ea38_7785, \16328 );
nor \g450946/U$1 ( \19372 , \19370 , \19371 );
and \g444992/U$2 ( \19373 , \19366 , \19369 , \19372 );
nor \g444992/U$1 ( \19374 , \19373 , \16389 );
and \g445792/U$2 ( \19375 , RIfc4e4b8_5913, \16319 );
and \g445792/U$3 ( \19376 , RIe202368_4315, \16313 );
and \g448616/U$2 ( \19377 , RIf15b750_5500, \16337 );
and \g448616/U$3 ( \19378 , \16341 , RIf15cc68_5515);
and \g448616/U$4 ( \19379 , RIf164558_5601, \16485 );
nor \g448616/U$1 ( \19380 , \19377 , \19378 , \19379 );
and \g454330/U$2 ( \19381 , \16317 , RIf15e180_5530);
and \g454330/U$3 ( \19382 , RIf160070_5552, \16325 );
nor \g454330/U$1 ( \19383 , \19381 , \19382 );
not \g449643/U$3 ( \19384 , \19383 );
not \g449643/U$4 ( \19385 , \16351 );
and \g449643/U$2 ( \19386 , \19384 , \19385 );
and \g449643/U$5 ( \19387 , \16354 , RIf165200_5610);
nor \g449643/U$1 ( \19388 , \19386 , \19387 );
and \g450989/U$2 ( \19389 , \16361 , RIf159c98_5481);
and \g450989/U$3 ( \19390 , RIf15a670_5488, \16364 );
nor \g450989/U$1 ( \19391 , \19389 , \19390 );
and \g450984/U$2 ( \19392 , \16368 , RIe1fb9f0_4240);
and \g450984/U$3 ( \19393 , RIe1fcc38_4253, \16371 );
nor \g450984/U$1 ( \19394 , \19392 , \19393 );
nand \g447519/U$1 ( \19395 , \19380 , \19388 , \19391 , \19394 );
nor \g445792/U$1 ( \19396 , \19375 , \19376 , \19395 );
and \g450979/U$2 ( \19397 , \16377 , RIe200a18_4297);
and \g450979/U$3 ( \19398 , RIf163478_5589, \16380 );
nor \g450979/U$1 ( \19399 , \19397 , \19398 );
and \g450978/U$2 ( \19400 , \16334 , RIf161f60_5574);
and \g450978/U$3 ( \19401 , RIfc86750_6552, \16328 );
nor \g450978/U$1 ( \19402 , \19400 , \19401 );
and \g444996/U$2 ( \19403 , \19396 , \19399 , \19402 );
nor \g444996/U$1 ( \19404 , \19403 , \16393 );
or \g444208/U$1 ( \19405 , \19344 , \19374 , \19404 );
_DC \g3919/U$1 ( \19406 , \19405 , \16652 );
and \g452006/U$2 ( \19407 , \16364 , RIe1ae470_3360);
and \g452006/U$3 ( \19408 , RIe1f7aa8_4195, \16371 );
nor \g452006/U$1 ( \19409 , \19407 , \19408 );
and \g446041/U$2 ( \19410 , RIe1fe6f0_4272, \16427 );
and \g446041/U$3 ( \19411 , RIe1f05f0_4112, \16368 );
and \g448945/U$2 ( \19412 , RIe178938_2749, \16485 );
and \g448945/U$3 ( \19413 , \16356 , RIe18c438_2973);
and \g448945/U$4 ( \19414 , RIe1bb5f8_3509, \16337 );
nor \g448945/U$1 ( \19415 , \19412 , \19413 , \19414 );
and \g454279/U$2 ( \19416 , \16317 , RIe1a5938_3261);
and \g454279/U$3 ( \19417 , RIe1a8638_3293, \16325 );
nor \g454279/U$1 ( \19418 , \19416 , \19417 );
not \g449956/U$3 ( \19419 , \19418 );
not \g449956/U$4 ( \19420 , \16311 );
and \g449956/U$2 ( \19421 , \19419 , \19420 );
and \g449956/U$5 ( \19422 , \16339 , RIe1d4af8_3797);
nor \g449956/U$1 ( \19423 , \19421 , \19422 );
and \g452027/U$2 ( \19424 , \16377 , RIe19ff38_3197);
and \g452027/U$3 ( \19425 , RIe1a2c38_3229, \16313 );
nor \g452027/U$1 ( \19426 , \19424 , \19425 );
and \g452030/U$2 ( \19427 , \16334 , RIe21ae90_4596);
and \g452030/U$3 ( \19428 , RIe226290_4724, \16380 );
nor \g452030/U$1 ( \19429 , \19427 , \19428 );
nand \g447324/U$1 ( \19430 , \19415 , \19423 , \19426 , \19429 );
nor \g446041/U$1 ( \19431 , \19410 , \19411 , \19430 );
and \g452013/U$2 ( \19432 , \16361 , RIe170aa8_2659);
and \g452013/U$3 ( \19433 , RIe204690_4340, \16448 );
nor \g452013/U$1 ( \19434 , \19432 , \19433 );
nand \g445584/U$1 ( \19435 , \19409 , \19431 , \19434 );
and \g444865/U$2 ( \19436 , \19435 , \16752 );
and \g448925/U$2 ( \19437 , RIe1cf0f8_3733, \16427 );
and \g448925/U$3 ( \19438 , \16448 , RIe1d1df8_3765);
and \g448925/U$4 ( \19439 , RIe1dd1f8_3893, \16485 );
nor \g448925/U$1 ( \19440 , \19437 , \19438 , \19439 );
and \g454650/U$2 ( \19441 , \16317 , RIe1c3cf8_3605);
and \g454650/U$3 ( \19442 , RIe1c69f8_3637, \16325 );
nor \g454650/U$1 ( \19443 , \19441 , \19442 );
not \g454649/U$1 ( \19444 , \19443 );
and \g449938/U$2 ( \19445 , \19444 , \16336 );
and \g449938/U$3 ( \19446 , RIe1dfef8_3925, \16356 );
nor \g449938/U$1 ( \19447 , \19445 , \19446 );
and \g451975/U$2 ( \19448 , \16361 , RIe1be2f8_3541);
and \g451975/U$3 ( \19449 , RIe1c0ff8_3573, \16364 );
nor \g451975/U$1 ( \19450 , \19448 , \19449 );
and \g451972/U$2 ( \19451 , \16368 , RIe1c96f8_3669);
and \g451972/U$3 ( \19452 , RIe1cc3f8_3701, \16371 );
nor \g451972/U$1 ( \19453 , \19451 , \19452 );
nand \g448060/U$1 ( \19454 , \19440 , \19447 , \19450 , \19453 );
and \g444865/U$3 ( \19455 , \16750 , \19454 );
nor \g444865/U$1 ( \19456 , \19436 , \19455 );
nor \g448354/U$1 ( \19457 , \16555 , \16320 );
and \g446811/U$2 ( \19458 , \19457 , RIe1e85f8_4021);
nor \g448353/U$1 ( \19459 , \16555 , \16327 );
and \g446811/U$3 ( \19460 , RIe1eb2f8_4053, \19459 );
nor \g446811/U$1 ( \19461 , \19458 , \19460 );
nor \g448324/U$1 ( \19462 , \16555 , \16510 );
and \g446810/U$2 ( \19463 , \19462 , RIe1d77f8_3829);
nor \g448356/U$1 ( \19464 , \16555 , \16513 );
and \g446810/U$3 ( \19465 , RIe1da4f8_3861, \19464 );
nor \g446810/U$1 ( \19466 , \19463 , \19465 );
nor \g448325/U$1 ( \19467 , \16555 , \16517 );
and \g446809/U$2 ( \19468 , \19467 , RIe1e2bf8_3957);
nor \g448355/U$1 ( \19469 , \16555 , \16520 );
and \g446809/U$3 ( \19470 , RIe1e58f8_3989, \19469 );
nor \g446809/U$1 ( \19471 , \19468 , \19470 );
nand \g444600/U$1 ( \19472 , \19456 , \19461 , \19466 , \19471 );
and \g451895/U$2 ( \19473 , \16377 , RIfe849d8_7853);
and \g451895/U$3 ( \19474 , RIfe83bc8_7843, \16380 );
nor \g451895/U$1 ( \19475 , \19473 , \19474 );
and \g446014/U$2 ( \19476 , RIf14b5f8_5317, \16321 );
and \g446014/U$3 ( \19477 , RIfe83a60_7842, \16313 );
and \g448905/U$2 ( \19478 , RIf147ae8_5275, \16427 );
and \g448905/U$3 ( \19479 , \16448 , RIf148d30_5288);
and \g448905/U$4 ( \19480 , RIf149b40_5298, \16485 );
nor \g448905/U$1 ( \19481 , \19478 , \19479 , \19480 );
and \g454540/U$2 ( \19482 , \16317 , RIf146300_5258);
and \g454540/U$3 ( \19483 , RIf146fa8_5267, \16325 );
nor \g454540/U$1 ( \19484 , \19482 , \19483 );
not \g454539/U$1 ( \19485 , \19484 );
and \g449923/U$2 ( \19486 , \19485 , \16336 );
and \g449923/U$3 ( \19487 , RIfc74168_6343, \16356 );
nor \g449923/U$1 ( \19488 , \19486 , \19487 );
and \g452338/U$2 ( \19489 , \16361 , RIfe83790_7840);
and \g452338/U$3 ( \19490 , RIfe845a0_7850, \16364 );
nor \g452338/U$1 ( \19491 , \19489 , \19490 );
and \g451917/U$2 ( \19492 , \16368 , RIe1b0900_3386);
and \g451917/U$3 ( \19493 , RIfe84870_7852, \16371 );
nor \g451917/U$1 ( \19494 , \19492 , \19493 );
nand \g448059/U$1 ( \19495 , \19481 , \19488 , \19491 , \19494 );
nor \g446014/U$1 ( \19496 , \19476 , \19477 , \19495 );
and \g453041/U$2 ( \19497 , \16334 , RIfe84708_7851);
and \g453041/U$3 ( \19498 , RIf14c840_5330, \16326 );
nor \g453041/U$1 ( \19499 , \19497 , \19498 );
nand \g445579/U$1 ( \19500 , \19475 , \19496 , \19499 );
and \g444914/U$2 ( \19501 , \19500 , \16477 );
and \g448889/U$2 ( \19502 , RIfc51fc8_5955, \16485 );
and \g448889/U$3 ( \19503 , \16356 , RIf156020_5438);
and \g448889/U$4 ( \19504 , RIf14eb68_5355, \16398 );
nor \g448889/U$1 ( \19505 , \19502 , \19503 , \19504 );
and \g455105/U$2 ( \19506 , \16317 , RIf157970_5456);
and \g455105/U$3 ( \19507 , RIf158d20_5470, \16325 );
nor \g455105/U$1 ( \19508 , \19506 , \19507 );
not \g449904/U$3 ( \19509 , \19508 );
not \g449904/U$4 ( \19510 , \16311 );
and \g449904/U$2 ( \19511 , \19509 , \19510 );
and \g449904/U$5 ( \19512 , \16339 , RIf14f810_5364);
nor \g449904/U$1 ( \19513 , \19511 , \19512 );
and \g451856/U$2 ( \19514 , \16377 , RIfe84438_7849);
and \g451856/U$3 ( \19515 , RIf156cc8_5447, \16313 );
nor \g451856/U$1 ( \19516 , \19514 , \19515 );
and \g452673/U$2 ( \19517 , \16334 , RIe1f51e0_4166);
and \g452673/U$3 ( \19518 , RIf154568_5419, \16380 );
nor \g452673/U$1 ( \19519 , \19517 , \19518 );
nand \g447315/U$1 ( \19520 , \19505 , \19513 , \19516 , \19519 );
and \g444914/U$3 ( \19521 , \16481 , \19520 );
nor \g444914/U$1 ( \19522 , \19501 , \19521 );
and \g446780/U$2 ( \19523 , \17274 , RIf1519d0_5388);
and \g446780/U$3 ( \19524 , RIf153050_5404, \17276 );
nor \g446780/U$1 ( \19525 , \19523 , \19524 );
and \g446787/U$2 ( \19526 , \17279 , RIfe842d0_7848);
and \g446787/U$3 ( \19527 , RIf150788_5375, \17281 );
nor \g446787/U$1 ( \19528 , \19526 , \19527 );
and \g446781/U$2 ( \19529 , \17284 , RIfe84168_7847);
and \g446781/U$3 ( \19530 , RIf14dd58_5345, \17286 );
nor \g446781/U$1 ( \19531 , \19529 , \19530 );
nand \g444597/U$1 ( \19532 , \19522 , \19525 , \19528 , \19531 );
and \g445964/U$2 ( \19533 , RIe223590_4692, \16321 );
and \g445964/U$3 ( \19534 , RIf16bce0_5686, \16313 );
and \g448847/U$2 ( \19535 , RIe212790_4500, \16427 );
and \g448847/U$3 ( \19536 , \16448 , RIf16a228_5667);
and \g448847/U$4 ( \19537 , RIe21db90_4628, \16485 );
nor \g448847/U$1 ( \19538 , \19535 , \19536 , \19537 );
and \g455094/U$2 ( \19539 , \16317 , RIe20cd90_4436);
and \g455094/U$3 ( \19540 , RIf167d98_5641, \16325 );
nor \g455094/U$1 ( \19541 , \19539 , \19540 );
not \g455093/U$1 ( \19542 , \19541 );
and \g449867/U$2 ( \19543 , \19542 , \16336 );
and \g449867/U$3 ( \19544 , RIf16ac00_5674, \16354 );
nor \g449867/U$1 ( \19545 , \19543 , \19544 );
and \g451744/U$2 ( \19546 , \16361 , RIe207390_4372);
and \g451744/U$3 ( \19547 , RIe20a090_4404, \16364 );
nor \g451744/U$1 ( \19548 , \19546 , \19547 );
and \g451736/U$2 ( \19549 , \16368 , RIe20fa90_4468);
and \g451736/U$3 ( \19550 , RIf168fe0_5654, \16371 );
nor \g451736/U$1 ( \19551 , \19549 , \19550 );
nand \g448052/U$1 ( \19552 , \19538 , \19545 , \19548 , \19551 );
nor \g445964/U$1 ( \19553 , \19533 , \19534 , \19552 );
and \g451722/U$2 ( \19554 , \16377 , RIe220890_4660);
and \g451722/U$3 ( \19555 , RIe218190_4564, \16380 );
nor \g451722/U$1 ( \19556 , \19554 , \19555 );
and \g451715/U$2 ( \19557 , \16334 , RIe215490_4532);
and \g451715/U$3 ( \19558 , RIf16caf0_5696, \16328 );
nor \g451715/U$1 ( \19559 , \19557 , \19558 );
and \g445118/U$2 ( \19560 , \19553 , \19556 , \19559 );
nor \g445118/U$1 ( \19561 , \19560 , \16389 );
and \g445991/U$2 ( \19562 , RIf1670f0_5632, \16328 );
and \g445991/U$3 ( \19563 , RIf161df8_5573, \16334 );
and \g448867/U$2 ( \19564 , RIf15e018_5529, \16427 );
and \g448867/U$3 ( \19565 , \16432 , RIf15ff08_5551);
and \g448867/U$4 ( \19566 , RIf1643f0_5600, \16485 );
nor \g448867/U$1 ( \19567 , \19564 , \19565 , \19566 );
and \g454686/U$2 ( \19568 , \16317 , RIf15b5e8_5499);
and \g454686/U$3 ( \19569 , RIf15cb00_5514, \16325 );
nor \g454686/U$1 ( \19570 , \19568 , \19569 );
not \g454685/U$1 ( \19571 , \19570 );
and \g449884/U$2 ( \19572 , \19571 , \16336 );
and \g449884/U$3 ( \19573 , RIf164f30_5608, \16356 );
nor \g449884/U$1 ( \19574 , \19572 , \19573 );
and \g451807/U$2 ( \19575 , \16361 , RIfc887a8_6575);
and \g451807/U$3 ( \19576 , RIf15a508_5487, \16364 );
nor \g451807/U$1 ( \19577 , \19575 , \19576 );
and \g451802/U$2 ( \19578 , \16368 , RIfe84000_7846);
and \g451802/U$3 ( \19579 , RIfe83d30_7844, \16371 );
nor \g451802/U$1 ( \19580 , \19578 , \19579 );
nand \g448055/U$1 ( \19581 , \19567 , \19574 , \19577 , \19580 );
nor \g445991/U$1 ( \19582 , \19562 , \19563 , \19581 );
and \g451782/U$2 ( \19583 , \16377 , RIfe83e98_7845);
and \g451782/U$3 ( \19584 , RIfce8310_7664, \16380 );
nor \g451782/U$1 ( \19585 , \19583 , \19584 );
and \g451778/U$2 ( \19586 , \16313 , RIe202200_4314);
and \g451778/U$3 ( \19587 , RIf165ea8_5619, \16319 );
nor \g451778/U$1 ( \19588 , \19586 , \19587 );
and \g445133/U$2 ( \19589 , \19582 , \19585 , \19588 );
nor \g445133/U$1 ( \19590 , \19589 , \16393 );
or \g444341/U$1 ( \19591 , \19472 , \19532 , \19561 , \19590 );
and \g445937/U$2 ( \19592 , RIe19a538_3133, \16321 );
and \g445937/U$3 ( \19593 , RIf145658_5249, \16313 );
and \g448808/U$2 ( \19594 , RIe186a38_2909, \16427 );
and \g448808/U$3 ( \19595 , \16432 , RIe189738_2941);
and \g448808/U$4 ( \19596 , RIe194b38_3069, \16344 );
nor \g448808/U$1 ( \19597 , \19594 , \19595 , \19596 );
and \g455195/U$2 ( \19598 , \16317 , RIe181038_2845);
and \g455195/U$3 ( \19599 , RIf142c28_5219, \16325 );
nor \g455195/U$1 ( \19600 , \19598 , \19599 );
not \g455194/U$1 ( \19601 , \19600 );
and \g449832/U$2 ( \19602 , \19601 , \16336 );
and \g449832/U$3 ( \19603 , RIf1446e0_5238, \16356 );
nor \g449832/U$1 ( \19604 , \19602 , \19603 );
and \g451629/U$2 ( \19605 , \16361 , RIe17b638_2781);
and \g451629/U$3 ( \19606 , RIe17e338_2813, \16364 );
nor \g451629/U$1 ( \19607 , \19605 , \19606 );
and \g451622/U$2 ( \19608 , \16368 , RIe183d38_2877);
and \g451622/U$3 ( \19609 , RIf143600_5226, \16371 );
nor \g451622/U$1 ( \19610 , \19608 , \19609 );
nand \g448044/U$1 ( \19611 , \19597 , \19604 , \19607 , \19610 );
nor \g445937/U$1 ( \19612 , \19592 , \19593 , \19611 );
and \g451604/U$2 ( \19613 , \16377 , RIe197838_3101);
and \g451604/U$3 ( \19614 , RIe191e38_3037, \16380 );
nor \g451604/U$1 ( \19615 , \19613 , \19614 );
and \g451597/U$2 ( \19616 , \16334 , RIe18f138_3005);
and \g451597/U$3 ( \19617 , RIe19d238_3165, \16328 );
nor \g451597/U$1 ( \19618 , \19616 , \19617 );
and \g445099/U$2 ( \19619 , \19612 , \19615 , \19618 );
nor \g445099/U$1 ( \19620 , \19619 , \16618 );
and \g445951/U$2 ( \19621 , RIee3c118_5142, \16432 );
and \g445951/U$3 ( \19622 , RIee39c88_5116, \16371 );
and \g448823/U$2 ( \19623 , RIf140a68_5195, \16319 );
and \g448823/U$3 ( \19624 , \16328 , RIf1420e8_5211);
and \g448823/U$4 ( \19625 , RIfc5ab00_6054, \16398 );
nor \g448823/U$1 ( \19626 , \19623 , \19624 , \19625 );
and \g454139/U$2 ( \19627 , \16317 , RIf13ee48_5175);
and \g454139/U$3 ( \19628 , RIf13faf0_5184, \16325 );
nor \g454139/U$1 ( \19629 , \19627 , \19628 );
not \g449848/U$3 ( \19630 , \19629 );
not \g449848/U$4 ( \19631 , \16330 );
and \g449848/U$2 ( \19632 , \19630 , \19631 );
and \g449848/U$5 ( \19633 , \16341 , RIf1701c8_5735);
nor \g449848/U$1 ( \19634 , \19632 , \19633 );
and \g451551/U$2 ( \19635 , \16377 , RIfebff10_8304);
and \g451551/U$3 ( \19636 , RIf1401f8_5189, \16313 );
nor \g451551/U$1 ( \19637 , \19635 , \19636 );
and \g451681/U$2 ( \19638 , \16334 , RIee3d1f8_5154);
and \g451681/U$3 ( \19639 , RIee3e2d8_5166, \16380 );
nor \g451681/U$1 ( \19640 , \19638 , \19639 );
nand \g447297/U$1 ( \19641 , \19626 , \19634 , \19637 , \19640 );
nor \g445951/U$1 ( \19642 , \19621 , \19622 , \19641 );
and \g451658/U$2 ( \19643 , \16364 , RIf16e008_5711);
and \g451658/U$3 ( \19644 , RIfe838f8_7841, \16368 );
nor \g451658/U$1 ( \19645 , \19643 , \19644 );
and \g451663/U$2 ( \19646 , \16361 , RIfcb0e88_7035);
and \g451663/U$3 ( \19647 , RIee3b038_5130, \16427 );
nor \g451663/U$1 ( \19648 , \19646 , \19647 );
and \g445110/U$2 ( \19649 , \19642 , \19645 , \19648 );
nor \g445110/U$1 ( \19650 , \19649 , \16649 );
or \g444270/U$1 ( \19651 , \19591 , \19620 , \19650 );
_DC \g399e/U$1 ( \19652 , \19651 , \16652 );
and \g452534/U$2 ( \19653 , \16377 , RIe175800_2714);
and \g452534/U$3 ( \19654 , RIfcc4280_7254, \16380 );
nor \g452534/U$1 ( \19655 , \19653 , \19654 );
and \g446160/U$2 ( \19656 , RIfc9ee40_6830, \16319 );
and \g446160/U$3 ( \19657 , RIe176e80_2730, \16313 );
and \g449087/U$2 ( \19658 , RIee3aed0_5129, \16427 );
and \g449087/U$3 ( \19659 , \16448 , RIee3bfb0_5141);
and \g449087/U$4 ( \19660 , RIfce0cf0_7580, \16485 );
nor \g449087/U$1 ( \19661 , \19658 , \19659 , \19660 );
and \g454902/U$2 ( \19662 , \16317 , RIf16f3b8_5725);
and \g454902/U$3 ( \19663 , RIf170060_5734, \16325 );
nor \g454902/U$1 ( \19664 , \19662 , \19663 );
not \g454901/U$1 ( \19665 , \19664 );
and \g450101/U$2 ( \19666 , \19665 , \16336 );
and \g450101/U$3 ( \19667 , RIfcb70f8_7105, \16354 );
nor \g450101/U$1 ( \19668 , \19666 , \19667 );
and \g452550/U$2 ( \19669 , \16361 , RIf16d4c8_5703);
and \g452550/U$3 ( \19670 , RIf16dea0_5710, \16364 );
nor \g452550/U$1 ( \19671 , \19669 , \19670 );
and \g452544/U$2 ( \19672 , \16368 , RIe173370_2688);
and \g452544/U$3 ( \19673 , RIee39b20_5115, \16371 );
nor \g452544/U$1 ( \19674 , \19672 , \19673 );
nand \g448077/U$1 ( \19675 , \19661 , \19668 , \19671 , \19674 );
nor \g446160/U$1 ( \19676 , \19656 , \19657 , \19675 );
and \g452531/U$2 ( \19677 , \16334 , RIfcba7d0_7144);
and \g452531/U$3 ( \19678 , RIfc9b060_6786, \16328 );
nor \g452531/U$1 ( \19679 , \19677 , \19678 );
nand \g445615/U$1 ( \19680 , \19655 , \19676 , \19679 );
and \g444781/U$2 ( \19681 , \19680 , \17998 );
and \g449079/U$2 ( \19682 , RIe20cc28_4435, \16398 );
and \g449079/U$3 ( \19683 , \16339 , RIf167c30_5640);
and \g449079/U$4 ( \19684 , RIe21da28_4627, \16485 );
nor \g449079/U$1 ( \19685 , \19682 , \19683 , \19684 );
and \g454892/U$2 ( \19686 , \16317 , RIe212628_4499);
and \g454892/U$3 ( \19687 , RIf16a0c0_5666, \16325 );
nor \g454892/U$1 ( \19688 , \19686 , \19687 );
not \g450093/U$3 ( \19689 , \19688 );
not \g450093/U$4 ( \19690 , \16351 );
and \g450093/U$2 ( \19691 , \19689 , \19690 );
and \g450093/U$5 ( \19692 , \16356 , RIf16aa98_5673);
nor \g450093/U$1 ( \19693 , \19691 , \19692 );
and \g452517/U$2 ( \19694 , \16361 , RIe207228_4371);
and \g452517/U$3 ( \19695 , RIe209f28_4403, \16364 );
nor \g452517/U$1 ( \19696 , \19694 , \19695 );
and \g452514/U$2 ( \19697 , \16368 , RIe20f928_4467);
and \g452514/U$3 ( \19698 , RIf168e78_5653, \16371 );
nor \g452514/U$1 ( \19699 , \19697 , \19698 );
nand \g447767/U$1 ( \19700 , \19685 , \19693 , \19696 , \19699 );
and \g444781/U$3 ( \19701 , \16390 , \19700 );
nor \g444781/U$1 ( \19702 , \19681 , \19701 );
and \g446926/U$2 ( \19703 , \18020 , RIe223428_4691);
and \g446926/U$3 ( \19704 , RIf16c988_5695, \18022 );
nor \g446926/U$1 ( \19705 , \19703 , \19704 );
and \g446930/U$2 ( \19706 , \18025 , RIe220728_4659);
and \g446930/U$3 ( \19707 , RIf16bb78_5685, \18027 );
nor \g446930/U$1 ( \19708 , \19706 , \19707 );
and \g446927/U$2 ( \19709 , \18030 , RIe215328_4531);
and \g446927/U$3 ( \19710 , RIe218028_4563, \18032 );
nor \g446927/U$1 ( \19711 , \19709 , \19710 );
nand \g444505/U$1 ( \19712 , \19702 , \19705 , \19708 , \19711 );
and \g452590/U$2 ( \19713 , \16371 , RIe1f7940_4194);
and \g452590/U$3 ( \19714 , RIe1fe588_4271, \16427 );
nor \g452590/U$1 ( \19715 , \19713 , \19714 );
and \g446171/U$2 ( \19716 , RIe204528_4339, \16448 );
and \g446171/U$3 ( \19717 , RIe170940_2658, \16361 );
and \g449103/U$2 ( \19718 , RIe1a57d0_3260, \16319 );
and \g449103/U$3 ( \19719 , \16326 , RIe1a84d0_3292);
and \g449103/U$4 ( \19720 , RIe1bb490_3508, \16337 );
nor \g449103/U$1 ( \19721 , \19718 , \19719 , \19720 );
and \g455396/U$2 ( \19722 , \16317 , RIe1787d0_2748);
and \g455396/U$3 ( \19723 , RIe18c2d0_2972, \16325 );
nor \g455396/U$1 ( \19724 , \19722 , \19723 );
not \g450118/U$3 ( \19725 , \19724 );
not \g450118/U$4 ( \19726 , \16330 );
and \g450118/U$2 ( \19727 , \19725 , \19726 );
and \g450118/U$5 ( \19728 , \16339 , RIe1d4990_3796);
nor \g450118/U$1 ( \19729 , \19727 , \19728 );
and \g452601/U$2 ( \19730 , \16377 , RIe19fdd0_3196);
and \g452601/U$3 ( \19731 , RIe1a2ad0_3228, \16313 );
nor \g452601/U$1 ( \19732 , \19730 , \19731 );
and \g452606/U$2 ( \19733 , \16334 , RIe21ad28_4595);
and \g452606/U$3 ( \19734 , RIe226128_4723, \16380 );
nor \g452606/U$1 ( \19735 , \19733 , \19734 );
nand \g447360/U$1 ( \19736 , \19721 , \19729 , \19732 , \19735 );
nor \g446171/U$1 ( \19737 , \19716 , \19717 , \19736 );
and \g452593/U$2 ( \19738 , \16364 , RIe1ae308_3359);
and \g452593/U$3 ( \19739 , RIe1f0488_4111, \16368 );
nor \g452593/U$1 ( \19740 , \19738 , \19739 );
nand \g445617/U$1 ( \19741 , \19715 , \19737 , \19740 );
and \g444894/U$2 ( \19742 , \19741 , \16752 );
and \g449096/U$2 ( \19743 , RIf147980_5274, \16427 );
and \g449096/U$3 ( \19744 , \16432 , RIf148bc8_5287);
and \g449096/U$4 ( \19745 , RIfc819f8_6497, \16344 );
nor \g449096/U$1 ( \19746 , \19743 , \19744 , \19745 );
and \g454911/U$2 ( \19747 , \16317 , RIf146198_5257);
and \g454911/U$3 ( \19748 , RIfcbb478_7153, \16325 );
nor \g454911/U$1 ( \19749 , \19747 , \19748 );
not \g454910/U$1 ( \19750 , \19749 );
and \g450110/U$2 ( \19751 , \19750 , \16336 );
and \g450110/U$3 ( \19752 , RIf14a248_5303, \16356 );
nor \g450110/U$1 ( \19753 , \19751 , \19752 );
and \g452577/U$2 ( \19754 , \16361 , RIfec08e8_8311);
and \g452577/U$3 ( \19755 , RIfe86058_7869, \16364 );
nor \g452577/U$1 ( \19756 , \19754 , \19755 );
and \g452572/U$2 ( \19757 , \16368 , RIfec0780_8310);
and \g452572/U$3 ( \19758 , RIfe86328_7871, \16371 );
nor \g452572/U$1 ( \19759 , \19757 , \19758 );
nand \g448079/U$1 ( \19760 , \19746 , \19753 , \19756 , \19759 );
and \g444894/U$3 ( \19761 , \16477 , \19760 );
nor \g444894/U$1 ( \19762 , \19742 , \19761 );
and \g446939/U$2 ( \19763 , \18268 , RIf14b490_5316);
and \g446939/U$3 ( \19764 , RIf14c6d8_5329, \18270 );
nor \g446939/U$1 ( \19765 , \19763 , \19764 );
and \g446940/U$2 ( \19766 , \18273 , RIfe86490_7872);
and \g446940/U$3 ( \19767 , RIfe85ef0_7868, \18275 );
nor \g446940/U$1 ( \19768 , \19766 , \19767 );
and \g446941/U$2 ( \19769 , \18278 , RIfe861c0_7870);
and \g446941/U$3 ( \19770 , RIfec0a50_8312, \18280 );
nor \g446941/U$1 ( \19771 , \19769 , \19770 );
nand \g444622/U$1 ( \19772 , \19762 , \19765 , \19768 , \19771 );
and \g446142/U$2 ( \19773 , RIe19a3d0_3132, \16321 );
and \g446142/U$3 ( \19774 , RIf1454f0_5248, \16313 );
and \g449064/U$2 ( \19775 , RIe1868d0_2908, \16427 );
and \g449064/U$3 ( \19776 , \16448 , RIe1895d0_2940);
and \g449064/U$4 ( \19777 , RIe1949d0_3068, \16485 );
nor \g449064/U$1 ( \19778 , \19775 , \19776 , \19777 );
and \g454865/U$2 ( \19779 , \16317 , RIe180ed0_2844);
and \g454865/U$3 ( \19780 , RIfc51758_5949, \16325 );
nor \g454865/U$1 ( \19781 , \19779 , \19780 );
not \g454864/U$1 ( \19782 , \19781 );
and \g450077/U$2 ( \19783 , \19782 , \16336 );
and \g450077/U$3 ( \19784 , RIf144578_5237, \16356 );
nor \g450077/U$1 ( \19785 , \19783 , \19784 );
and \g452461/U$2 ( \19786 , \16361 , RIe17b4d0_2780);
and \g452461/U$3 ( \19787 , RIe17e1d0_2812, \16364 );
nor \g452461/U$1 ( \19788 , \19786 , \19787 );
and \g452458/U$2 ( \19789 , \16368 , RIe183bd0_2876);
and \g452458/U$3 ( \19790 , RIf143498_5225, \16371 );
nor \g452458/U$1 ( \19791 , \19789 , \19790 );
nand \g448073/U$1 ( \19792 , \19778 , \19785 , \19788 , \19791 );
nor \g446142/U$1 ( \19793 , \19773 , \19774 , \19792 );
and \g452452/U$2 ( \19794 , \16377 , RIe1976d0_3100);
and \g452452/U$3 ( \19795 , RIe191cd0_3036, \16380 );
nor \g452452/U$1 ( \19796 , \19794 , \19795 );
and \g452448/U$2 ( \19797 , \16334 , RIe18efd0_3004);
and \g452448/U$3 ( \19798 , RIe19d0d0_3164, \16328 );
nor \g452448/U$1 ( \19799 , \19797 , \19798 );
and \g445251/U$2 ( \19800 , \19793 , \19796 , \19799 );
nor \g445251/U$1 ( \19801 , \19800 , \16618 );
and \g446147/U$2 ( \19802 , RIf15deb0_5528, \16427 );
and \g446147/U$3 ( \19803 , RIfe85d88_7867, \16368 );
and \g449072/U$2 ( \19804 , RIf165d40_5618, \16321 );
and \g449072/U$3 ( \19805 , \16328 , RIf166f88_5631);
and \g449072/U$4 ( \19806 , RIf15b480_5498, \16398 );
nor \g449072/U$1 ( \19807 , \19804 , \19805 , \19806 );
and \g454220/U$2 ( \19808 , \16317 , RIf164288_5599);
and \g454220/U$3 ( \19809 , RIfc52b08_5963, \16325 );
nor \g454220/U$1 ( \19810 , \19808 , \19809 );
not \g450084/U$3 ( \19811 , \19810 );
not \g450084/U$4 ( \19812 , \16330 );
and \g450084/U$2 ( \19813 , \19811 , \19812 );
and \g450084/U$5 ( \19814 , \16341 , RIf15c998_5513);
nor \g450084/U$1 ( \19815 , \19813 , \19814 );
and \g452484/U$2 ( \19816 , \16377 , RIfe86760_7874);
and \g452484/U$3 ( \19817 , RIfec0618_8309, \16313 );
nor \g452484/U$1 ( \19818 , \19816 , \19817 );
and \g452489/U$2 ( \19819 , \16334 , RIf161c90_5572);
and \g452489/U$3 ( \19820 , RIf163310_5588, \16380 );
nor \g452489/U$1 ( \19821 , \19819 , \19820 );
nand \g447353/U$1 ( \19822 , \19807 , \19815 , \19818 , \19821 );
nor \g446147/U$1 ( \19823 , \19802 , \19803 , \19822 );
and \g452476/U$2 ( \19824 , \16361 , RIf159b30_5480);
and \g452476/U$3 ( \19825 , RIf15fda0_5550, \16448 );
nor \g452476/U$1 ( \19826 , \19824 , \19825 );
and \g452472/U$2 ( \19827 , \16364 , RIf15a3a0_5486);
and \g452472/U$3 ( \19828 , RIfe865f8_7873, \16371 );
nor \g452472/U$1 ( \19829 , \19827 , \19828 );
and \g445253/U$2 ( \19830 , \19823 , \19826 , \19829 );
nor \g445253/U$1 ( \19831 , \19830 , \16393 );
or \g444400/U$1 ( \19832 , \19712 , \19772 , \19801 , \19831 );
and \g446129/U$2 ( \19833 , RIf152ee8_5403, \16448 );
and \g446129/U$3 ( \19834 , RIf150620_5374, \16371 );
and \g449049/U$2 ( \19835 , RIfc4ade0_5874, \16321 );
and \g449049/U$3 ( \19836 , \16328 , RIfc83348_6515);
and \g449049/U$4 ( \19837 , RIf14ea00_5354, \16398 );
nor \g449049/U$1 ( \19838 , \19835 , \19836 , \19837 );
and \g454838/U$2 ( \19839 , \16317 , RIfc9f110_6832);
and \g454838/U$3 ( \19840 , RIfc4ac78_5873, \16325 );
nor \g454838/U$1 ( \19841 , \19839 , \19840 );
not \g450062/U$3 ( \19842 , \19841 );
not \g450062/U$4 ( \19843 , \16330 );
and \g450062/U$2 ( \19844 , \19842 , \19843 );
and \g450062/U$5 ( \19845 , \16341 , RIf14f6a8_5363);
nor \g450062/U$1 ( \19846 , \19844 , \19845 );
and \g452400/U$2 ( \19847 , \16377 , RIe1f9f38_4221);
and \g452400/U$3 ( \19848 , RIfc89720_6586, \16313 );
nor \g452400/U$1 ( \19849 , \19847 , \19848 );
and \g452404/U$2 ( \19850 , \16334 , RIe1f5078_4165);
and \g452404/U$3 ( \19851 , RIfc4ab10_5872, \16380 );
nor \g452404/U$1 ( \19852 , \19850 , \19851 );
nand \g447350/U$1 ( \19853 , \19838 , \19846 , \19849 , \19852 );
nor \g446129/U$1 ( \19854 , \19833 , \19834 , \19853 );
and \g452390/U$2 ( \19855 , \16364 , RIf14dbf0_5344);
and \g452390/U$3 ( \19856 , RIe1f2eb8_4141, \16368 );
nor \g452390/U$1 ( \19857 , \19855 , \19856 );
and \g452393/U$2 ( \19858 , \16361 , RIe1edbc0_4082);
and \g452393/U$3 ( \19859 , RIfc899f0_6588, \16427 );
nor \g452393/U$1 ( \19860 , \19858 , \19859 );
and \g445240/U$2 ( \19861 , \19854 , \19857 , \19860 );
nor \g445240/U$1 ( \19862 , \19861 , \16480 );
and \g446135/U$2 ( \19863 , RIe1d1c90_3764, \16448 );
and \g446135/U$3 ( \19864 , RIe1cc290_3700, \16371 );
and \g449057/U$2 ( \19865 , RIe1dd090_3892, \16344 );
and \g449057/U$3 ( \19866 , \16356 , RIe1dfd90_3924);
and \g449057/U$4 ( \19867 , RIe1c3b90_3604, \16398 );
nor \g449057/U$1 ( \19868 , \19865 , \19866 , \19867 );
and \g454856/U$2 ( \19869 , \16317 , RIe1e8490_4020);
and \g454856/U$3 ( \19870 , RIe1eb190_4052, \16325 );
nor \g454856/U$1 ( \19871 , \19869 , \19870 );
not \g450069/U$3 ( \19872 , \19871 );
not \g450069/U$4 ( \19873 , \16311 );
and \g450069/U$2 ( \19874 , \19872 , \19873 );
and \g450069/U$5 ( \19875 , \16339 , RIe1c6890_3636);
nor \g450069/U$1 ( \19876 , \19874 , \19875 );
and \g452426/U$2 ( \19877 , \16377 , RIe1e2a90_3956);
and \g452426/U$3 ( \19878 , RIe1e5790_3988, \16313 );
nor \g452426/U$1 ( \19879 , \19877 , \19878 );
and \g452432/U$2 ( \19880 , \16334 , RIe1d7690_3828);
and \g452432/U$3 ( \19881 , RIe1da390_3860, \16380 );
nor \g452432/U$1 ( \19882 , \19880 , \19881 );
nand \g447351/U$1 ( \19883 , \19868 , \19876 , \19879 , \19882 );
nor \g446135/U$1 ( \19884 , \19863 , \19864 , \19883 );
and \g452416/U$2 ( \19885 , \16364 , RIe1c0e90_3572);
and \g452416/U$3 ( \19886 , RIe1c9590_3668, \16368 );
nor \g452416/U$1 ( \19887 , \19885 , \19886 );
and \g452419/U$2 ( \19888 , \16361 , RIe1be190_3540);
and \g452419/U$3 ( \19889 , RIe1cef90_3732, \16427 );
nor \g452419/U$1 ( \19890 , \19888 , \19889 );
and \g445245/U$2 ( \19891 , \19884 , \19887 , \19890 );
nor \g445245/U$1 ( \19892 , \19891 , \16555 );
or \g444260/U$1 ( \19893 , \19832 , \19862 , \19892 );
_DC \g3a23/U$1 ( \19894 , \19893 , \16652 );
and \g453195/U$2 ( \19895 , \16377 , RIe2205c0_4658);
and \g453195/U$3 ( \19896 , RIe217ec0_4562, \16380 );
nor \g453195/U$1 ( \19897 , \19895 , \19896 );
and \g446298/U$2 ( \19898 , RIe2232c0_4690, \16321 );
and \g446298/U$3 ( \19899 , RIf16ba10_5684, \16313 );
and \g449279/U$2 ( \19900 , RIe20cac0_4434, \16398 );
and \g449279/U$3 ( \19901 , \16341 , RIfc7d240_6446);
and \g449279/U$4 ( \19902 , RIe21d8c0_4626, \16485 );
nor \g449279/U$1 ( \19903 , \19900 , \19901 , \19902 );
and \g454485/U$2 ( \19904 , \16317 , RIe2124c0_4498);
and \g454485/U$3 ( \19905 , RIfebf268_8295, \16325 );
nor \g454485/U$1 ( \19906 , \19904 , \19905 );
not \g450293/U$3 ( \19907 , \19906 );
not \g450293/U$4 ( \19908 , \16351 );
and \g450293/U$2 ( \19909 , \19907 , \19908 );
and \g450293/U$5 ( \19910 , \16354 , RIfcd24e8_7415);
nor \g450293/U$1 ( \19911 , \19909 , \19910 );
and \g453236/U$2 ( \19912 , \16361 , RIe2070c0_4370);
and \g453236/U$3 ( \19913 , RIe209dc0_4402, \16364 );
nor \g453236/U$1 ( \19914 , \19912 , \19913 );
and \g453222/U$2 ( \19915 , \16368 , RIe20f7c0_4466);
and \g453222/U$3 ( \19916 , RIf168d10_5652, \16371 );
nor \g453222/U$1 ( \19917 , \19915 , \19916 );
nand \g447865/U$1 ( \19918 , \19903 , \19911 , \19914 , \19917 );
nor \g446298/U$1 ( \19919 , \19898 , \19899 , \19918 );
and \g453172/U$2 ( \19920 , \16334 , RIe2151c0_4530);
and \g453172/U$3 ( \19921 , RIfe82ae8_7831, \16328 );
nor \g453172/U$1 ( \19922 , \19920 , \19921 );
nand \g445649/U$1 ( \19923 , \19897 , \19919 , \19922 );
and \g444862/U$2 ( \19924 , \19923 , \16390 );
and \g449246/U$2 ( \19925 , RIfebf6a0_8298, \16321 );
and \g449246/U$3 ( \19926 , \16328 , RIf166e20_5630);
and \g449246/U$4 ( \19927 , RIf15b318_5497, \16398 );
nor \g449246/U$1 ( \19928 , \19925 , \19926 , \19927 );
and \g455238/U$2 ( \19929 , \16317 , RIf164120_5598);
and \g455238/U$3 ( \19930 , RIfc8eb80_6646, \16325 );
nor \g455238/U$1 ( \19931 , \19929 , \19930 );
not \g450253/U$3 ( \19932 , \19931 );
not \g450253/U$4 ( \19933 , \16330 );
and \g450253/U$2 ( \19934 , \19932 , \19933 );
and \g450253/U$5 ( \19935 , \16341 , RIfebf3d0_8296);
nor \g450253/U$1 ( \19936 , \19934 , \19935 );
and \g453081/U$2 ( \19937 , \16377 , RIfebf538_8297);
and \g453081/U$3 ( \19938 , RIfebf808_8299, \16313 );
nor \g453081/U$1 ( \19939 , \19937 , \19938 );
and \g453089/U$2 ( \19940 , \16334 , RIf161b28_5571);
and \g453089/U$3 ( \19941 , RIfc453e0_5810, \16380 );
nor \g453089/U$1 ( \19942 , \19940 , \19941 );
nand \g447397/U$1 ( \19943 , \19928 , \19936 , \19939 , \19942 );
and \g444862/U$3 ( \19944 , \16394 , \19943 );
nor \g444862/U$1 ( \19945 , \19924 , \19944 );
and \g447038/U$2 ( \19946 , \16419 , RIfc8f120_6650);
and \g447038/U$3 ( \19947 , RIfca2518_6869, \16422 );
nor \g447038/U$1 ( \19948 , \19946 , \19947 );
and \g447024/U$2 ( \19949 , \16429 , RIf15dd48_5527);
and \g447024/U$3 ( \19950 , RIf15fc38_5549, \16434 );
nor \g447024/U$1 ( \19951 , \19949 , \19950 );
and \g447034/U$2 ( \19952 , \16438 , RIe1fb888_4239);
and \g447034/U$3 ( \19953 , RIe1fc968_4251, \16441 );
nor \g447034/U$1 ( \19954 , \19952 , \19953 );
nand \g444636/U$1 ( \19955 , \19945 , \19948 , \19951 , \19954 );
and \g452858/U$2 ( \19956 , \16380 , RIfc7dc18_6453);
and \g452858/U$3 ( \19957 , RIfcd6700_7462, \16321 );
nor \g452858/U$1 ( \19958 , \19956 , \19957 );
and \g446232/U$2 ( \19959 , RIfc564b0_6004, \16328 );
and \g446232/U$3 ( \19960 , RIe175698_2713, \16377 );
and \g449200/U$2 ( \19961 , RIfcc2a98_7237, \16427 );
and \g449200/U$3 ( \19962 , \16448 , RIfc98630_6756);
and \g449200/U$4 ( \19963 , RIfc45f20_5818, \16485 );
nor \g449200/U$1 ( \19964 , \19961 , \19962 , \19963 );
and \g454958/U$2 ( \19965 , \16317 , RIfc45ae8_5815);
and \g454958/U$3 ( \19966 , RIfc8e478_6641, \16325 );
nor \g454958/U$1 ( \19967 , \19965 , \19966 );
not \g454957/U$1 ( \19968 , \19967 );
and \g450207/U$2 ( \19969 , \19968 , \16336 );
and \g450207/U$3 ( \19970 , RIfc46088_5819, \16356 );
nor \g450207/U$1 ( \19971 , \19969 , \19970 );
and \g452926/U$2 ( \19972 , \16361 , RIfc45980_5814);
and \g452926/U$3 ( \19973 , RIfc8e8b0_6644, \16364 );
nor \g452926/U$1 ( \19974 , \19972 , \19973 );
and \g452910/U$2 ( \19975 , \16368 , RIe173208_2687);
and \g452910/U$3 ( \19976 , RIfc7d510_6448, \16371 );
nor \g452910/U$1 ( \19977 , \19975 , \19976 );
nand \g448093/U$1 ( \19978 , \19964 , \19971 , \19974 , \19977 );
nor \g446232/U$1 ( \19979 , \19959 , \19960 , \19978 );
and \g452865/U$2 ( \19980 , \16334 , RIfcd69d0_7464);
and \g452865/U$3 ( \19981 , RIfc461f0_5820, \16313 );
nor \g452865/U$1 ( \19982 , \19980 , \19981 );
nand \g445632/U$1 ( \19983 , \19958 , \19979 , \19982 );
and \g444710/U$2 ( \19984 , \19983 , \17998 );
and \g449158/U$2 ( \19985 , RIe19a268_3131, \16321 );
and \g449158/U$3 ( \19986 , \16328 , RIe19cf68_3163);
and \g449158/U$4 ( \19987 , RIe180d68_2843, \16398 );
nor \g449158/U$1 ( \19988 , \19985 , \19986 , \19987 );
and \g455024/U$2 ( \19989 , \16317 , RIe194868_3067);
and \g455024/U$3 ( \19990 , RIfc561e0_6002, \16325 );
nor \g455024/U$1 ( \19991 , \19989 , \19990 );
not \g450167/U$3 ( \19992 , \19991 );
not \g450167/U$4 ( \19993 , \16330 );
and \g450167/U$2 ( \19994 , \19992 , \19993 );
and \g450167/U$5 ( \19995 , \16341 , RIfc7d948_6451);
nor \g450167/U$1 ( \19996 , \19994 , \19995 );
and \g452758/U$2 ( \19997 , \16377 , RIe197568_3099);
and \g452758/U$3 ( \19998 , RIfc8d7d0_6632, \16313 );
nor \g452758/U$1 ( \19999 , \19997 , \19998 );
and \g452776/U$2 ( \20000 , \16334 , RIe18ee68_3003);
and \g452776/U$3 ( \20001 , RIe191b68_3035, \16380 );
nor \g452776/U$1 ( \20002 , \20000 , \20001 );
nand \g447377/U$1 ( \20003 , \19988 , \19996 , \19999 , \20002 );
and \g444710/U$3 ( \20004 , \17938 , \20003 );
nor \g444710/U$1 ( \20005 , \19984 , \20004 );
and \g446960/U$2 ( \20006 , \18457 , RIe186768_2907);
and \g446960/U$3 ( \20007 , RIe189468_2939, \18459 );
nor \g446960/U$1 ( \20008 , \20006 , \20007 );
and \g446961/U$2 ( \20009 , \18462 , RIe183a68_2875);
and \g446961/U$3 ( \20010 , RIf143330_5224, \18464 );
nor \g446961/U$1 ( \20011 , \20009 , \20010 );
and \g446971/U$2 ( \20012 , \18467 , RIe17b368_2779);
and \g446971/U$3 ( \20013 , RIe17e068_2811, \18469 );
nor \g446971/U$1 ( \20014 , \20012 , \20013 );
nand \g444511/U$1 ( \20015 , \20005 , \20008 , \20011 , \20014 );
and \g446140/U$2 ( \20016 , RIe1cee28_3731, \16427 );
and \g446140/U$3 ( \20017 , RIe1c9428_3667, \16368 );
and \g449075/U$2 ( \20018 , RIe1e8328_4019, \16319 );
and \g449075/U$3 ( \20019 , \16328 , RIe1eb028_4051);
and \g449075/U$4 ( \20020 , RIe1c3a28_3603, \16398 );
nor \g449075/U$1 ( \20021 , \20018 , \20019 , \20020 );
and \g454879/U$2 ( \20022 , \16317 , RIe1dcf28_3891);
and \g454879/U$3 ( \20023 , RIe1dfc28_3923, \16325 );
nor \g454879/U$1 ( \20024 , \20022 , \20023 );
not \g450086/U$3 ( \20025 , \20024 );
not \g450086/U$4 ( \20026 , \16330 );
and \g450086/U$2 ( \20027 , \20025 , \20026 );
and \g450086/U$5 ( \20028 , \16341 , RIe1c6728_3635);
nor \g450086/U$1 ( \20029 , \20027 , \20028 );
and \g452466/U$2 ( \20030 , \16377 , RIe1e2928_3955);
and \g452466/U$3 ( \20031 , RIe1e5628_3987, \16313 );
nor \g452466/U$1 ( \20032 , \20030 , \20031 );
and \g452481/U$2 ( \20033 , \16334 , RIe1d7528_3827);
and \g452481/U$3 ( \20034 , RIe1da228_3859, \16380 );
nor \g452481/U$1 ( \20035 , \20033 , \20034 );
nand \g447352/U$1 ( \20036 , \20021 , \20029 , \20032 , \20035 );
nor \g446140/U$1 ( \20037 , \20016 , \20017 , \20036 );
and \g452441/U$2 ( \20038 , \16361 , RIe1be028_3539);
and \g452441/U$3 ( \20039 , RIe1d1b28_3763, \16448 );
nor \g452441/U$1 ( \20040 , \20038 , \20039 );
and \g452430/U$2 ( \20041 , \16364 , RIe1c0d28_3571);
and \g452430/U$3 ( \20042 , RIe1cc128_3699, \16371 );
nor \g452430/U$1 ( \20043 , \20041 , \20042 );
and \g445249/U$2 ( \20044 , \20037 , \20040 , \20043 );
nor \g445249/U$1 ( \20045 , \20044 , \16555 );
and \g446165/U$2 ( \20046 , RIe1fe420_4270, \16427 );
and \g446165/U$3 ( \20047 , RIe1f0320_4110, \16368 );
and \g449109/U$2 ( \20048 , RIe178668_2747, \16485 );
and \g449109/U$3 ( \20049 , \16356 , RIe18c168_2971);
and \g449109/U$4 ( \20050 , RIe1bb328_3507, \16398 );
nor \g449109/U$1 ( \20051 , \20048 , \20049 , \20050 );
and \g454936/U$2 ( \20052 , \16317 , RIe1a5668_3259);
and \g454936/U$3 ( \20053 , RIe1a8368_3291, \16325 );
nor \g454936/U$1 ( \20054 , \20052 , \20053 );
not \g450119/U$3 ( \20055 , \20054 );
not \g450119/U$4 ( \20056 , \16311 );
and \g450119/U$2 ( \20057 , \20055 , \20056 );
and \g450119/U$5 ( \20058 , \16341 , RIe1d4828_3795);
nor \g450119/U$1 ( \20059 , \20057 , \20058 );
and \g452582/U$2 ( \20060 , \16377 , RIe19fc68_3195);
and \g452582/U$3 ( \20061 , RIe1a2968_3227, \16313 );
nor \g452582/U$1 ( \20062 , \20060 , \20061 );
and \g452595/U$2 ( \20063 , \16334 , RIe21abc0_4594);
and \g452595/U$3 ( \20064 , RIe225fc0_4722, \16380 );
nor \g452595/U$1 ( \20065 , \20063 , \20064 );
nand \g447359/U$1 ( \20066 , \20051 , \20059 , \20062 , \20065 );
nor \g446165/U$1 ( \20067 , \20046 , \20047 , \20066 );
and \g452555/U$2 ( \20068 , \16361 , RIe1707d8_2657);
and \g452555/U$3 ( \20069 , RIe2043c0_4338, \16448 );
nor \g452555/U$1 ( \20070 , \20068 , \20069 );
and \g452547/U$2 ( \20071 , \16364 , RIe1ae1a0_3358);
and \g452547/U$3 ( \20072 , RIe1f77d8_4193, \16371 );
nor \g452547/U$1 ( \20073 , \20071 , \20072 );
and \g445267/U$2 ( \20074 , \20067 , \20070 , \20073 );
nor \g445267/U$1 ( \20075 , \20074 , \16586 );
or \g444354/U$1 ( \20076 , \19955 , \20015 , \20045 , \20075 );
and \g446085/U$2 ( \20077 , RIfebf970_8300, \16321 );
and \g446085/U$3 ( \20078 , RIfc7cca0_6442, \16313 );
and \g449006/U$2 ( \20079 , RIfc8f828_6655, \16427 );
and \g449006/U$3 ( \20080 , \16356 , RIfe82c50_7832);
and \g449006/U$4 ( \20081 , RIfc8faf8_6657, \16398 );
nor \g449006/U$1 ( \20082 , \20079 , \20080 , \20081 );
and \g452221/U$2 ( \20083 , \16334 , RIe1f4f10_4164);
and \g452221/U$3 ( \20084 , RIfc8f288_6651, \16380 );
nor \g452221/U$1 ( \20085 , \20083 , \20084 );
and \g454772/U$2 ( \20086 , \16331 , RIe1f2d50_4140);
not \g455682/U$1 ( \20087 , \16308 );
and \g454772/U$3 ( \20088 , RIfcb3b88_7067, \20087 );
nor \g454772/U$1 ( \20089 , \20086 , \20088 );
not \g450014/U$3 ( \20090 , \20089 );
not \g450014/U$4 ( \20091 , \16351 );
and \g450014/U$2 ( \20092 , \20090 , \20091 );
and \g450014/U$5 ( \20093 , \16341 , RIfc445d0_5800);
nor \g450014/U$1 ( \20094 , \20092 , \20093 );
and \g452206/U$2 ( \20095 , \16485 , RIf155648_5431);
and \g452206/U$3 ( \20096 , RIf152d80_5402, \16432 );
nor \g452206/U$1 ( \20097 , \20095 , \20096 );
nand \g447338/U$1 ( \20098 , \20082 , \20085 , \20094 , \20097 );
nor \g446085/U$1 ( \20099 , \20077 , \20078 , \20098 );
and \g452163/U$2 ( \20100 , \16364 , RIf14da88_5343);
and \g452163/U$3 ( \20101 , RIe1f9dd0_4220, \16377 );
nor \g452163/U$1 ( \20102 , \20100 , \20101 );
and \g452142/U$2 ( \20103 , \16361 , RIe1eda58_4081);
and \g452142/U$3 ( \20104 , RIfebfad8_8301, \16328 );
nor \g452142/U$1 ( \20105 , \20103 , \20104 );
and \g445203/U$2 ( \20106 , \20099 , \20102 , \20105 );
nor \g445203/U$1 ( \20107 , \20106 , \16480 );
and \g446112/U$2 ( \20108 , RIfc44030_5796, \16321 );
and \g446112/U$3 ( \20109 , RIe1b9000_3482, \16313 );
and \g449045/U$2 ( \20110 , RIfc7ba58_6429, \16398 );
and \g449045/U$3 ( \20111 , \16341 , RIfcdb5c0_7518);
and \g449045/U$4 ( \20112 , RIfc8ff30_6660, \16485 );
nor \g449045/U$1 ( \20113 , \20110 , \20111 , \20112 );
and \g454297/U$2 ( \20114 , \16317 , RIfc43d60_5794);
and \g454297/U$3 ( \20115 , RIfcbe178_7185, \16325 );
nor \g454297/U$1 ( \20116 , \20114 , \20115 );
not \g450052/U$3 ( \20117 , \20116 );
not \g450052/U$4 ( \20118 , \16351 );
and \g450052/U$2 ( \20119 , \20117 , \20118 );
and \g450052/U$5 ( \20120 , \16356 , RIfcbdd40_7182);
nor \g450052/U$1 ( \20121 , \20119 , \20120 );
and \g452359/U$2 ( \20122 , \16361 , RIe1aa960_3318);
and \g452359/U$3 ( \20123 , RIe1ac148_3335, \16364 );
nor \g452359/U$1 ( \20124 , \20122 , \20123 );
and \g452346/U$2 ( \20125 , \16368 , RIe1b0798_3385);
and \g452346/U$3 ( \20126 , RIe1b2520_3406, \16371 );
nor \g452346/U$1 ( \20127 , \20125 , \20126 );
nand \g447744/U$1 ( \20128 , \20113 , \20121 , \20124 , \20127 );
nor \g446112/U$1 ( \20129 , \20108 , \20109 , \20128 );
and \g452310/U$2 ( \20130 , \16377 , RIe1b6fa8_3459);
and \g452310/U$3 ( \20131 , RIe1b50b8_3437, \16380 );
nor \g452310/U$1 ( \20132 , \20130 , \20131 );
and \g452302/U$2 ( \20133 , \16334 , RIe1b3d08_3423);
and \g452302/U$3 ( \20134 , RIfc7bff8_6433, \16328 );
nor \g452302/U$1 ( \20135 , \20133 , \20134 );
and \g445225/U$2 ( \20136 , \20129 , \20132 , \20135 );
nor \g445225/U$1 ( \20137 , \20136 , \16909 );
or \g444181/U$1 ( \20138 , \20076 , \20107 , \20137 );
_DC \g3aa8/U$1 ( \20139 , \20138 , \16652 );
and \g452471/U$2 ( \20140 , \16371 , RIe1f7670_4192);
and \g452471/U$3 ( \20141 , RIe1fe2b8_4269, \16427 );
nor \g452471/U$1 ( \20142 , \20140 , \20141 );
and \g446145/U$2 ( \20143 , RIe204258_4337, \16448 );
and \g446145/U$3 ( \20144 , RIe170670_2656, \16361 );
and \g449077/U$2 ( \20145 , RIe178500_2746, \16485 );
and \g449077/U$3 ( \20146 , \16356 , RIe18c000_2970);
and \g449077/U$4 ( \20147 , RIe1bb1c0_3506, \16398 );
nor \g449077/U$1 ( \20148 , \20145 , \20146 , \20147 );
and \g454882/U$2 ( \20149 , \16317 , RIe1a5500_3258);
and \g454882/U$3 ( \20150 , RIe1a8200_3290, \16325 );
nor \g454882/U$1 ( \20151 , \20149 , \20150 );
not \g450089/U$3 ( \20152 , \20151 );
not \g450089/U$4 ( \20153 , \16311 );
and \g450089/U$2 ( \20154 , \20152 , \20153 );
and \g450089/U$5 ( \20155 , \16341 , RIe1d46c0_3794);
nor \g450089/U$1 ( \20156 , \20154 , \20155 );
and \g452498/U$2 ( \20157 , \16377 , RIe19fb00_3194);
and \g452498/U$3 ( \20158 , RIe1a2800_3226, \16313 );
nor \g452498/U$1 ( \20159 , \20157 , \20158 );
and \g452501/U$2 ( \20160 , \16334 , RIe21aa58_4593);
and \g452501/U$3 ( \20161 , RIe225e58_4721, \16380 );
nor \g452501/U$1 ( \20162 , \20160 , \20161 );
nand \g447355/U$1 ( \20163 , \20148 , \20156 , \20159 , \20162 );
nor \g446145/U$1 ( \20164 , \20143 , \20144 , \20163 );
and \g452474/U$2 ( \20165 , \16364 , RIe1ae038_3357);
and \g452474/U$3 ( \20166 , RIe1f01b8_4109, \16368 );
nor \g452474/U$1 ( \20167 , \20165 , \20166 );
nand \g445610/U$1 ( \20168 , \20142 , \20164 , \20167 );
and \g444893/U$2 ( \20169 , \20168 , \16752 );
and \g449060/U$2 ( \20170 , RIfcc0ba8_7215, \16337 );
and \g449060/U$3 ( \20171 , \16341 , RIfcdd8e8_7543);
and \g449060/U$4 ( \20172 , RIfc94b20_6714, \16485 );
nor \g449060/U$1 ( \20173 , \20170 , \20171 , \20172 );
and \g454862/U$2 ( \20174 , \16317 , RIfceb010_7696);
and \g454862/U$3 ( \20175 , RIfcec3c0_7710, \16325 );
nor \g454862/U$1 ( \20176 , \20174 , \20175 );
not \g450074/U$3 ( \20177 , \20176 );
not \g450074/U$4 ( \20178 , \16351 );
and \g450074/U$2 ( \20179 , \20177 , \20178 );
and \g450074/U$5 ( \20180 , \16356 , RIfc76760_6370);
nor \g450074/U$1 ( \20181 , \20179 , \20180 );
and \g452447/U$2 ( \20182 , \16361 , RIe1aa7f8_3317);
and \g452447/U$3 ( \20183 , RIfe82278_7825, \16364 );
nor \g452447/U$1 ( \20184 , \20182 , \20183 );
and \g452438/U$2 ( \20185 , \16368 , RIfe82110_7824);
and \g452438/U$3 ( \20186 , RIfe823e0_7826, \16371 );
nor \g452438/U$1 ( \20187 , \20185 , \20186 );
nand \g447754/U$1 ( \20188 , \20173 , \20181 , \20184 , \20187 );
and \g444893/U$3 ( \20189 , \16477 , \20188 );
nor \g444893/U$1 ( \20190 , \20169 , \20189 );
and \g446904/U$2 ( \20191 , \18268 , RIf14b328_5315);
and \g446904/U$3 ( \20192 , RIf14c570_5328, \18270 );
nor \g446904/U$1 ( \20193 , \20191 , \20192 );
and \g446908/U$2 ( \20194 , \18273 , RIe1b6e40_3458);
and \g446908/U$3 ( \20195 , RIe1b8e98_3481, \18275 );
nor \g446908/U$1 ( \20196 , \20194 , \20195 );
and \g446911/U$2 ( \20197 , \18278 , RIe1b3ba0_3422);
and \g446911/U$3 ( \20198 , RIe1b4f50_3436, \18280 );
nor \g446911/U$1 ( \20199 , \20197 , \20198 );
nand \g444616/U$1 ( \20200 , \20190 , \20193 , \20196 , \20199 );
and \g452353/U$2 ( \20201 , \16361 , RIe1bdec0_3538);
and \g452353/U$3 ( \20202 , RIe1cecc0_3730, \16427 );
nor \g452353/U$1 ( \20203 , \20201 , \20202 );
and \g446120/U$2 ( \20204 , RIe1d19c0_3762, \16448 );
and \g446120/U$3 ( \20205 , RIe1cbfc0_3698, \16371 );
and \g449043/U$2 ( \20206 , RIe1e81c0_4018, \16321 );
and \g449043/U$3 ( \20207 , \16328 , RIe1eaec0_4050);
and \g449043/U$4 ( \20208 , RIe1c38c0_3602, \16398 );
nor \g449043/U$1 ( \20209 , \20206 , \20207 , \20208 );
and \g454300/U$2 ( \20210 , \16317 , RIe1dcdc0_3890);
and \g454300/U$3 ( \20211 , RIe1dfac0_3922, \16325 );
nor \g454300/U$1 ( \20212 , \20210 , \20211 );
not \g450056/U$3 ( \20213 , \20212 );
not \g450056/U$4 ( \20214 , \16330 );
and \g450056/U$2 ( \20215 , \20213 , \20214 );
and \g450056/U$5 ( \20216 , \16341 , RIe1c65c0_3634);
nor \g450056/U$1 ( \20217 , \20215 , \20216 );
and \g452375/U$2 ( \20218 , \16377 , RIe1e27c0_3954);
and \g452375/U$3 ( \20219 , RIe1e54c0_3986, \16313 );
nor \g452375/U$1 ( \20220 , \20218 , \20219 );
and \g452385/U$2 ( \20221 , \16334 , RIe1d73c0_3826);
and \g452385/U$3 ( \20222 , RIe1da0c0_3858, \16380 );
nor \g452385/U$1 ( \20223 , \20221 , \20222 );
nand \g447349/U$1 ( \20224 , \20209 , \20217 , \20220 , \20223 );
nor \g446120/U$1 ( \20225 , \20204 , \20205 , \20224 );
and \g452348/U$2 ( \20226 , \16364 , RIe1c0bc0_3570);
and \g452348/U$3 ( \20227 , RIe1c92c0_3666, \16368 );
nor \g452348/U$1 ( \20228 , \20226 , \20227 );
nand \g445605/U$1 ( \20229 , \20203 , \20225 , \20228 );
and \g444776/U$2 ( \20230 , \20229 , \16750 );
and \g449026/U$2 ( \20231 , RIfcd7ab0_7476, \16485 );
and \g449026/U$3 ( \20232 , \16356 , RIfcc8a38_7305);
and \g449026/U$4 ( \20233 , RIfc772a0_6378, \16398 );
nor \g449026/U$1 ( \20234 , \20231 , \20232 , \20233 );
and \g454802/U$2 ( \20235 , \16317 , RIf157808_5455);
and \g454802/U$3 ( \20236 , RIf158bb8_5469, \16325 );
nor \g454802/U$1 ( \20237 , \20235 , \20236 );
not \g450037/U$3 ( \20238 , \20237 );
not \g450037/U$4 ( \20239 , \16311 );
and \g450037/U$2 ( \20240 , \20238 , \20239 );
and \g450037/U$5 ( \20241 , \16341 , RIf14f540_5362);
nor \g450037/U$1 ( \20242 , \20240 , \20241 );
and \g452309/U$2 ( \20243 , \16377 , RIfebef98_8293);
and \g452309/U$3 ( \20244 , RIfc5d0f8_6081, \16313 );
nor \g452309/U$1 ( \20245 , \20243 , \20244 );
and \g452313/U$2 ( \20246 , \16334 , RIfeaa0e8_8251);
and \g452313/U$3 ( \20247 , RIfcb1428_7039, \16380 );
nor \g452313/U$1 ( \20248 , \20246 , \20247 );
nand \g447345/U$1 ( \20249 , \20234 , \20242 , \20245 , \20248 );
and \g444776/U$3 ( \20250 , \16481 , \20249 );
nor \g444776/U$1 ( \20251 , \20230 , \20250 );
and \g446877/U$2 ( \20252 , \17274 , RIfce3450_7608);
and \g446877/U$3 ( \20253 , RIfccc548_7347, \17276 );
nor \g446877/U$1 ( \20254 , \20252 , \20253 );
and \g446878/U$2 ( \20255 , \17279 , RIe1f2be8_4139);
and \g446878/U$3 ( \20256 , RIf1504b8_5373, \17281 );
nor \g446878/U$1 ( \20257 , \20255 , \20256 );
and \g446879/U$2 ( \20258 , \17284 , RIe1ed8f0_4080);
and \g446879/U$3 ( \20259 , RIfcec258_7709, \17286 );
nor \g446879/U$1 ( \20260 , \20258 , \20259 );
nand \g444497/U$1 ( \20261 , \20251 , \20254 , \20257 , \20260 );
and \g446069/U$2 ( \20262 , RIe186600_2906, \16427 );
and \g446069/U$3 ( \20263 , RIe183900_2874, \16368 );
and \g448985/U$2 ( \20264 , RIe19a100_3130, \16321 );
and \g448985/U$3 ( \20265 , \16328 , RIe19ce00_3162);
and \g448985/U$4 ( \20266 , RIe180c00_2842, \16337 );
nor \g448985/U$1 ( \20267 , \20264 , \20265 , \20266 );
and \g454430/U$2 ( \20268 , \16317 , RIe194700_3066);
and \g454430/U$3 ( \20269 , RIf144410_5236, \16325 );
nor \g454430/U$1 ( \20270 , \20268 , \20269 );
not \g449987/U$3 ( \20271 , \20270 );
not \g449987/U$4 ( \20272 , \16330 );
and \g449987/U$2 ( \20273 , \20271 , \20272 );
and \g449987/U$5 ( \20274 , \16339 , RIfcdbcc8_7523);
nor \g449987/U$1 ( \20275 , \20273 , \20274 );
and \g452115/U$2 ( \20276 , \16377 , RIe197400_3098);
and \g452115/U$3 ( \20277 , RIfce96c0_7678, \16313 );
nor \g452115/U$1 ( \20278 , \20276 , \20277 );
and \g452161/U$2 ( \20279 , \16334 , RIe18ed00_3002);
and \g452161/U$3 ( \20280 , RIe191a00_3034, \16380 );
nor \g452161/U$1 ( \20281 , \20279 , \20280 );
nand \g447334/U$1 ( \20282 , \20267 , \20275 , \20278 , \20281 );
nor \g446069/U$1 ( \20283 , \20262 , \20263 , \20282 );
and \g452110/U$2 ( \20284 , \16361 , RIe17b200_2778);
and \g452110/U$3 ( \20285 , RIe189300_2938, \16448 );
nor \g452110/U$1 ( \20286 , \20284 , \20285 );
and \g452098/U$2 ( \20287 , \16364 , RIe17df00_2810);
and \g452098/U$3 ( \20288 , RIfebee30_8292, \16371 );
nor \g452098/U$1 ( \20289 , \20287 , \20288 );
and \g445193/U$2 ( \20290 , \20283 , \20286 , \20289 );
nor \g445193/U$1 ( \20291 , \20290 , \16618 );
and \g446090/U$2 ( \20292 , RIf166cb8_5629, \16328 );
and \g446090/U$3 ( \20293 , RIf1619c0_5570, \16334 );
and \g449002/U$2 ( \20294 , RIf15b1b0_5496, \16398 );
and \g449002/U$3 ( \20295 , \16341 , RIf15c830_5512);
and \g449002/U$4 ( \20296 , RIfceb178_7697, \16344 );
nor \g449002/U$1 ( \20297 , \20294 , \20295 , \20296 );
and \g454767/U$2 ( \20298 , \16317 , RIfc77570_6380);
and \g454767/U$3 ( \20299 , RIfccf248_7379, \16325 );
nor \g454767/U$1 ( \20300 , \20298 , \20299 );
not \g450013/U$3 ( \20301 , \20300 );
not \g450013/U$4 ( \20302 , \16351 );
and \g450013/U$2 ( \20303 , \20301 , \20302 );
and \g450013/U$5 ( \20304 , \16356 , RIfc5c888_6075);
nor \g450013/U$1 ( \20305 , \20303 , \20304 );
and \g452237/U$2 ( \20306 , \16361 , RIfccc6b0_7348);
and \g452237/U$3 ( \20307 , RIfcd0fd0_7400, \16364 );
nor \g452237/U$1 ( \20308 , \20306 , \20307 );
and \g452226/U$2 ( \20309 , \16368 , RIe1fb720_4238);
and \g452226/U$3 ( \20310 , RIe1fc800_4250, \16371 );
nor \g452226/U$1 ( \20311 , \20309 , \20310 );
nand \g447725/U$1 ( \20312 , \20297 , \20305 , \20308 , \20311 );
nor \g446090/U$1 ( \20313 , \20292 , \20293 , \20312 );
and \g452207/U$2 ( \20314 , \16377 , RIfe81e40_7822);
and \g452207/U$3 ( \20315 , RIf1631a8_5587, \16380 );
nor \g452207/U$1 ( \20316 , \20314 , \20315 );
and \g452200/U$2 ( \20317 , \16313 , RIfe81fa8_7823);
and \g452200/U$3 ( \20318 , RIf165bd8_5617, \16319 );
nor \g452200/U$1 ( \20319 , \20317 , \20318 );
and \g445210/U$2 ( \20320 , \20313 , \20316 , \20319 );
nor \g445210/U$1 ( \20321 , \20320 , \16393 );
or \g444392/U$1 ( \20322 , \20200 , \20261 , \20291 , \20321 );
and \g446012/U$2 ( \20323 , RIfce7398_7653, \16321 );
and \g446012/U$3 ( \20324 , RIfcb1e00_7046, \16313 );
and \g448912/U$2 ( \20325 , RIfebecc8_8291, \16398 );
and \g448912/U$3 ( \20326 , \16339 , RIf16fef8_5733);
and \g448912/U$4 ( \20327 , RIfcbff00_7206, \16485 );
nor \g448912/U$1 ( \20328 , \20325 , \20326 , \20327 );
and \g454805/U$2 ( \20329 , \16317 , RIfce35b8_7609);
and \g454805/U$3 ( \20330 , RIfc5c180_6070, \16325 );
nor \g454805/U$1 ( \20331 , \20329 , \20330 );
not \g449882/U$3 ( \20332 , \20331 );
not \g449882/U$4 ( \20333 , \16351 );
and \g449882/U$2 ( \20334 , \20332 , \20333 );
and \g449882/U$5 ( \20335 , \16354 , RIfca42a0_6890);
nor \g449882/U$1 ( \20336 , \20334 , \20335 );
and \g452068/U$2 ( \20337 , \16361 , RIfce9288_7675);
and \g452068/U$3 ( \20338 , RIfc5c450_6072, \16364 );
nor \g452068/U$1 ( \20339 , \20337 , \20338 );
and \g451914/U$2 ( \20340 , \16368 , RIfea8a68_8235);
and \g451914/U$3 ( \20341 , RIee399b8_5114, \16371 );
nor \g451914/U$1 ( \20342 , \20340 , \20341 );
nand \g447666/U$1 ( \20343 , \20328 , \20336 , \20339 , \20342 );
nor \g446012/U$1 ( \20344 , \20323 , \20324 , \20343 );
and \g451880/U$2 ( \20345 , \16377 , RIfe82548_7827);
and \g451880/U$3 ( \20346 , RIfcaaee8_6967, \16380 );
nor \g451880/U$1 ( \20347 , \20345 , \20346 );
and \g451870/U$2 ( \20348 , \16334 , RIee3d090_5153);
and \g451870/U$3 ( \20349 , RIf141f80_5210, \16328 );
nor \g451870/U$1 ( \20350 , \20348 , \20349 );
and \g445149/U$2 ( \20351 , \20344 , \20347 , \20350 );
nor \g445149/U$1 ( \20352 , \20351 , \16649 );
and \g446037/U$2 ( \20353 , RIe212358_4497, \16427 );
and \g446037/U$3 ( \20354 , RIe20f658_4465, \16368 );
and \g448854/U$2 ( \20355 , RIe21d758_4625, \16485 );
and \g448854/U$3 ( \20356 , \16356 , RIfce24d8_7597);
and \g448854/U$4 ( \20357 , RIe20c958_4433, \16398 );
nor \g448854/U$1 ( \20358 , \20355 , \20356 , \20357 );
and \g455017/U$2 ( \20359 , \16317 , RIe223158_4689);
and \g455017/U$3 ( \20360 , RIfc40778_5759, \16325 );
nor \g455017/U$1 ( \20361 , \20359 , \20360 );
not \g449959/U$3 ( \20362 , \20361 );
not \g449959/U$4 ( \20363 , \16311 );
and \g449959/U$2 ( \20364 , \20362 , \20363 );
and \g449959/U$5 ( \20365 , \16341 , RIfc77840_6382);
nor \g449959/U$1 ( \20366 , \20364 , \20365 );
and \g452732/U$2 ( \20367 , \16377 , RIe220458_4657);
and \g452732/U$3 ( \20368 , RIfce77d0_7656, \16313 );
nor \g452732/U$1 ( \20369 , \20367 , \20368 );
and \g452031/U$2 ( \20370 , \16334 , RIe215058_4529);
and \g452031/U$3 ( \20371 , RIe217d58_4561, \16380 );
nor \g452031/U$1 ( \20372 , \20370 , \20371 );
nand \g447323/U$1 ( \20373 , \20358 , \20366 , \20369 , \20372 );
nor \g446037/U$1 ( \20374 , \20353 , \20354 , \20373 );
and \g451994/U$2 ( \20375 , \16361 , RIe206f58_4369);
and \g451994/U$3 ( \20376 , RIfce8a18_7669, \16432 );
nor \g451994/U$1 ( \20377 , \20375 , \20376 );
and \g451984/U$2 ( \20378 , \16364 , RIe209c58_4401);
and \g451984/U$3 ( \20379 , RIfce1998_7589, \16371 );
nor \g451984/U$1 ( \20380 , \20378 , \20379 );
and \g445170/U$2 ( \20381 , \20374 , \20377 , \20380 );
nor \g445170/U$1 ( \20382 , \20381 , \16389 );
or \g444215/U$1 ( \20383 , \20322 , \20352 , \20382 );
_DC \g3b2d/U$1 ( \20384 , \20383 , \16652 );
and \g451930/U$2 ( \20385 , \16361 , RIfc62120_6138);
and \g451930/U$3 ( \20386 , RIee3ad68_5128, \16427 );
nor \g451930/U$1 ( \20387 , \20385 , \20386 );
and \g446019/U$2 ( \20388 , RIee3be48_5140, \16432 );
and \g446019/U$3 ( \20389 , RIfc71fa8_6319, \16371 );
and \g448906/U$2 ( \20390 , RIfc726b0_6324, \16485 );
and \g448906/U$3 ( \20391 , \16356 , RIfc72818_6325);
and \g448906/U$4 ( \20392 , RIfccf518_7381, \16337 );
nor \g448906/U$1 ( \20393 , \20390 , \20391 , \20392 );
and \g454388/U$2 ( \20394 , \16317 , RIfca6a00_6918);
and \g454388/U$3 ( \20395 , RIfcaf268_7015, \16325 );
nor \g454388/U$1 ( \20396 , \20394 , \20395 );
not \g449925/U$3 ( \20397 , \20396 );
not \g449925/U$4 ( \20398 , \16311 );
and \g449925/U$2 ( \20399 , \20397 , \20398 );
and \g449925/U$5 ( \20400 , \16341 , RIfcaef98_7013);
nor \g449925/U$1 ( \20401 , \20399 , \20400 );
and \g451889/U$2 ( \20402 , \16377 , RIe175530_2712);
and \g451889/U$3 ( \20403 , RIfcc9b18_7317, \16313 );
nor \g451889/U$1 ( \20404 , \20402 , \20403 );
and \g451933/U$2 ( \20405 , \16334 , RIfc72548_6323);
and \g451933/U$3 ( \20406 , RIfccf7e8_7383, \16380 );
nor \g451933/U$1 ( \20407 , \20405 , \20406 );
nand \g447321/U$1 ( \20408 , \20393 , \20401 , \20404 , \20407 );
nor \g446019/U$1 ( \20409 , \20388 , \20389 , \20408 );
and \g451945/U$2 ( \20410 , \16364 , RIfc71e40_6318);
and \g451945/U$3 ( \20411 , RIe1730a0_2686, \16368 );
nor \g451945/U$1 ( \20412 , \20410 , \20411 );
nand \g445581/U$1 ( \20413 , \20387 , \20409 , \20412 );
and \g444705/U$2 ( \20414 , \20413 , \17998 );
and \g448903/U$2 ( \20415 , RIe194598_3065, \16344 );
and \g448903/U$3 ( \20416 , \16356 , RIf1442a8_5235);
and \g448903/U$4 ( \20417 , RIe180a98_2841, \16398 );
nor \g448903/U$1 ( \20418 , \20415 , \20416 , \20417 );
and \g454531/U$2 ( \20419 , \16317 , RIe199f98_3129);
and \g454531/U$3 ( \20420 , RIe19cc98_3161, \16325 );
nor \g454531/U$1 ( \20421 , \20419 , \20420 );
not \g449924/U$3 ( \20422 , \20421 );
not \g449924/U$4 ( \20423 , \16311 );
and \g449924/U$2 ( \20424 , \20422 , \20423 );
and \g449924/U$5 ( \20425 , \16341 , RIfc61ce8_6135);
nor \g449924/U$1 ( \20426 , \20424 , \20425 );
and \g451928/U$2 ( \20427 , \16377 , RIe197298_3097);
and \g451928/U$3 ( \20428 , RIfc73088_6331, \16313 );
nor \g451928/U$1 ( \20429 , \20427 , \20428 );
and \g451929/U$2 ( \20430 , \16334 , RIe18eb98_3001);
and \g451929/U$3 ( \20431 , RIe191898_3033, \16380 );
nor \g451929/U$1 ( \20432 , \20430 , \20431 );
nand \g447320/U$1 ( \20433 , \20418 , \20426 , \20429 , \20432 );
and \g444705/U$3 ( \20434 , \17938 , \20433 );
nor \g444705/U$1 ( \20435 , \20414 , \20434 );
and \g446803/U$2 ( \20436 , \18457 , RIe186498_2905);
and \g446803/U$3 ( \20437 , RIe189198_2937, \18459 );
nor \g446803/U$1 ( \20438 , \20436 , \20437 );
and \g446804/U$2 ( \20439 , \18462 , RIe183798_2873);
and \g446804/U$3 ( \20440 , RIfc72278_6321, \18464 );
nor \g446804/U$1 ( \20441 , \20439 , \20440 );
and \g446805/U$2 ( \20442 , \18467 , RIe17b098_2777);
and \g446805/U$3 ( \20443 , RIe17dd98_2809, \18469 );
nor \g446805/U$1 ( \20444 , \20442 , \20443 );
nand \g444485/U$1 ( \20445 , \20435 , \20438 , \20441 , \20444 );
and \g451939/U$2 ( \20446 , \16364 , RIe1aded0_3356);
and \g451939/U$3 ( \20447 , RIe1f7508_4191, \16371 );
nor \g451939/U$1 ( \20448 , \20446 , \20447 );
and \g446022/U$2 ( \20449 , RIe1fe150_4268, \16427 );
and \g446022/U$3 ( \20450 , RIe1f0050_4108, \16368 );
and \g448909/U$2 ( \20451 , RIe1a5398_3257, \16321 );
and \g448909/U$3 ( \20452 , \16328 , RIe1a8098_3289);
and \g448909/U$4 ( \20453 , RIe1bb058_3505, \16398 );
nor \g448909/U$1 ( \20454 , \20451 , \20452 , \20453 );
and \g454693/U$2 ( \20455 , \16317 , RIe178398_2745);
and \g454693/U$3 ( \20456 , RIe18be98_2969, \16325 );
nor \g454693/U$1 ( \20457 , \20455 , \20456 );
not \g449929/U$3 ( \20458 , \20457 );
not \g449929/U$4 ( \20459 , \16330 );
and \g449929/U$2 ( \20460 , \20458 , \20459 );
and \g449929/U$5 ( \20461 , \16339 , RIe1d4558_3793);
nor \g449929/U$1 ( \20462 , \20460 , \20461 );
and \g451942/U$2 ( \20463 , \16377 , RIe19f998_3193);
and \g451942/U$3 ( \20464 , RIe1a2698_3225, \16313 );
nor \g451942/U$1 ( \20465 , \20463 , \20464 );
and \g451943/U$2 ( \20466 , \16334 , RIe21a8f0_4592);
and \g451943/U$3 ( \20467 , RIe225cf0_4720, \16380 );
nor \g451943/U$1 ( \20468 , \20466 , \20467 );
nand \g447322/U$1 ( \20469 , \20454 , \20462 , \20465 , \20468 );
nor \g446022/U$1 ( \20470 , \20449 , \20450 , \20469 );
and \g451940/U$2 ( \20471 , \16361 , RIe170508_2655);
and \g451940/U$3 ( \20472 , RIe2040f0_4336, \16432 );
nor \g451940/U$1 ( \20473 , \20471 , \20472 );
nand \g445582/U$1 ( \20474 , \20448 , \20470 , \20473 );
and \g444770/U$2 ( \20475 , \20474 , \16752 );
and \g448907/U$2 ( \20476 , RIe1c3758_3601, \16398 );
and \g448907/U$3 ( \20477 , \16341 , RIe1c6458_3633);
and \g448907/U$4 ( \20478 , RIe1dcc58_3889, \16485 );
nor \g448907/U$1 ( \20479 , \20476 , \20477 , \20478 );
and \g455317/U$2 ( \20480 , \16317 , RIe1ceb58_3729);
and \g455317/U$3 ( \20481 , RIe1d1858_3761, \16325 );
nor \g455317/U$1 ( \20482 , \20480 , \20481 );
not \g449926/U$3 ( \20483 , \20482 );
not \g449926/U$4 ( \20484 , \16351 );
and \g449926/U$2 ( \20485 , \20483 , \20484 );
and \g449926/U$5 ( \20486 , \16356 , RIe1df958_3921);
nor \g449926/U$1 ( \20487 , \20485 , \20486 );
and \g451937/U$2 ( \20488 , \16361 , RIe1bdd58_3537);
and \g451937/U$3 ( \20489 , RIe1c0a58_3569, \16364 );
nor \g451937/U$1 ( \20490 , \20488 , \20489 );
and \g451936/U$2 ( \20491 , \16368 , RIe1c9158_3665);
and \g451936/U$3 ( \20492 , RIe1cbe58_3697, \16371 );
nor \g451936/U$1 ( \20493 , \20491 , \20492 );
nand \g447672/U$1 ( \20494 , \20479 , \20487 , \20490 , \20493 );
and \g444770/U$3 ( \20495 , \16750 , \20494 );
nor \g444770/U$1 ( \20496 , \20475 , \20495 );
and \g446806/U$2 ( \20497 , \19457 , RIe1e8058_4017);
and \g446806/U$3 ( \20498 , RIe1ead58_4049, \19459 );
nor \g446806/U$1 ( \20499 , \20497 , \20498 );
and \g446808/U$2 ( \20500 , \19462 , RIe1d7258_3825);
and \g446808/U$3 ( \20501 , RIe1d9f58_3857, \19464 );
nor \g446808/U$1 ( \20502 , \20500 , \20501 );
and \g446807/U$2 ( \20503 , \19467 , RIe1e2658_3953);
and \g446807/U$3 ( \20504 , RIe1e5358_3985, \19469 );
nor \g446807/U$1 ( \20505 , \20503 , \20504 );
nand \g444602/U$1 ( \20506 , \20496 , \20499 , \20502 , \20505 );
and \g446016/U$2 ( \20507 , RIfc70220_6298, \16448 );
and \g446016/U$3 ( \20508 , RIe1aa690_3316, \16361 );
and \g448899/U$2 ( \20509 , RIf14b1c0_5314, \16321 );
and \g448899/U$3 ( \20510 , \16328 , RIf14c408_5327);
and \g448899/U$4 ( \20511 , RIfc700b8_6297, \16398 );
nor \g448899/U$1 ( \20512 , \20509 , \20510 , \20511 );
and \g454774/U$2 ( \20513 , \16317 , RIfca7c48_6931);
and \g454774/U$3 ( \20514 , RIfc707c0_6302, \16325 );
nor \g454774/U$1 ( \20515 , \20513 , \20514 );
not \g450026/U$3 ( \20516 , \20515 );
not \g450026/U$4 ( \20517 , \16330 );
and \g450026/U$2 ( \20518 , \20516 , \20517 );
and \g450026/U$5 ( \20519 , \16341 , RIfc645b0_6164);
nor \g450026/U$1 ( \20520 , \20518 , \20519 );
and \g451920/U$2 ( \20521 , \16377 , RIe1b6cd8_3457);
and \g451920/U$3 ( \20522 , RIe1b8d30_3480, \16313 );
nor \g451920/U$1 ( \20523 , \20521 , \20522 );
and \g451921/U$2 ( \20524 , \16334 , RIe1b3a38_3421);
and \g451921/U$3 ( \20525 , RIe1b4de8_3435, \16380 );
nor \g451921/U$1 ( \20526 , \20524 , \20525 );
nand \g447318/U$1 ( \20527 , \20512 , \20520 , \20523 , \20526 );
nor \g446016/U$1 ( \20528 , \20507 , \20508 , \20527 );
and \g451919/U$2 ( \20529 , \16364 , RIfeaac28_8259);
and \g451919/U$3 ( \20530 , RIe1b0630_3384, \16368 );
nor \g451919/U$1 ( \20531 , \20529 , \20530 );
and \g451918/U$2 ( \20532 , \16371 , RIe1b23b8_3405);
and \g451918/U$3 ( \20533 , RIfcce870_7372, \16427 );
nor \g451918/U$1 ( \20534 , \20532 , \20533 );
and \g445162/U$2 ( \20535 , \20528 , \20531 , \20534 );
nor \g445162/U$1 ( \20536 , \20535 , \16909 );
and \g446017/U$2 ( \20537 , RIf151868_5387, \16427 );
and \g446017/U$3 ( \20538 , RIe1f2a80_4138, \16368 );
and \g448900/U$2 ( \20539 , RIfcceb40_7374, \16485 );
and \g448900/U$3 ( \20540 , \16356 , RIfc634d0_6152);
and \g448900/U$4 ( \20541 , RIfc63bd8_6157, \16398 );
nor \g448900/U$1 ( \20542 , \20539 , \20540 , \20541 );
and \g454449/U$2 ( \20543 , \16317 , RIf1576a0_5454);
and \g454449/U$3 ( \20544 , RIf158a50_5468, \16325 );
nor \g454449/U$1 ( \20545 , \20543 , \20544 );
not \g449921/U$3 ( \20546 , \20545 );
not \g449921/U$4 ( \20547 , \16311 );
and \g449921/U$2 ( \20548 , \20546 , \20547 );
and \g449921/U$5 ( \20549 , \16341 , RIfc70a90_6304);
nor \g449921/U$1 ( \20550 , \20548 , \20549 );
and \g452088/U$2 ( \20551 , \16377 , RIfe8b620_7930);
and \g452088/U$3 ( \20552 , RIfcdc808_7531, \16313 );
nor \g452088/U$1 ( \20553 , \20551 , \20552 );
and \g451926/U$2 ( \20554 , \16334 , RIe1f4da8_4163);
and \g451926/U$3 ( \20555 , RIf154400_5418, \16380 );
nor \g451926/U$1 ( \20556 , \20554 , \20555 );
nand \g447319/U$1 ( \20557 , \20542 , \20550 , \20553 , \20556 );
nor \g446017/U$1 ( \20558 , \20537 , \20538 , \20557 );
and \g452203/U$2 ( \20559 , \16361 , RIe1ed788_4079);
and \g452203/U$3 ( \20560 , RIf152c18_5401, \16448 );
nor \g452203/U$1 ( \20561 , \20559 , \20560 );
and \g451923/U$2 ( \20562 , \16364 , RIfca7810_6928);
and \g451923/U$3 ( \20563 , RIfc4d108_5899, \16371 );
nor \g451923/U$1 ( \20564 , \20562 , \20563 );
and \g445164/U$2 ( \20565 , \20558 , \20561 , \20564 );
nor \g445164/U$1 ( \20566 , \20565 , \16480 );
or \g444329/U$1 ( \20567 , \20445 , \20506 , \20536 , \20566 );
and \g446013/U$2 ( \20568 , RIe222ff0_4688, \16321 );
and \g446013/U$3 ( \20569 , RIfcc9f50_7320, \16313 );
and \g448896/U$2 ( \20570 , RIe2121f0_4496, \16427 );
and \g448896/U$3 ( \20571 , \16448 , RIfccf3b0_7380);
and \g448896/U$4 ( \20572 , RIe21d5f0_4624, \16485 );
nor \g448896/U$1 ( \20573 , \20570 , \20571 , \20572 );
and \g454923/U$2 ( \20574 , \16317 , RIe20c7f0_4432);
and \g454923/U$3 ( \20575 , RIfc71300_6310, \16325 );
nor \g454923/U$1 ( \20576 , \20574 , \20575 );
not \g454922/U$1 ( \20577 , \20576 );
and \g449917/U$2 ( \20578 , \20577 , \16336 );
and \g449917/U$3 ( \20579 , RIfc4a570_5868, \16356 );
nor \g449917/U$1 ( \20580 , \20578 , \20579 );
and \g451910/U$2 ( \20581 , \16361 , RIe206df0_4368);
and \g451910/U$3 ( \20582 , RIe209af0_4400, \16364 );
nor \g451910/U$1 ( \20583 , \20581 , \20582 );
and \g451908/U$2 ( \20584 , \16368 , RIe20f4f0_4464);
and \g451908/U$3 ( \20585 , RIf168ba8_5651, \16371 );
nor \g451908/U$1 ( \20586 , \20584 , \20585 );
nand \g448058/U$1 ( \20587 , \20573 , \20580 , \20583 , \20586 );
nor \g446013/U$1 ( \20588 , \20568 , \20569 , \20587 );
and \g451906/U$2 ( \20589 , \16377 , RIe2202f0_4656);
and \g451906/U$3 ( \20590 , RIe217bf0_4560, \16380 );
nor \g451906/U$1 ( \20591 , \20589 , \20590 );
and \g451905/U$2 ( \20592 , \16334 , RIe214ef0_4528);
and \g451905/U$3 ( \20593 , RIfe8b350_7928, \16328 );
nor \g451905/U$1 ( \20594 , \20592 , \20593 );
and \g445160/U$2 ( \20595 , \20588 , \20591 , \20594 );
nor \g445160/U$1 ( \20596 , \20595 , \16389 );
and \g446015/U$2 ( \20597 , RIf15fad0_5548, \16448 );
and \g446015/U$3 ( \20598 , RIe1fc698_4249, \16371 );
and \g448898/U$2 ( \20599 , RIfce6588_7643, \16485 );
and \g448898/U$3 ( \20600 , \16356 , RIfc715d0_6312);
and \g448898/U$4 ( \20601 , RIfc63098_6149, \16398 );
nor \g448898/U$1 ( \20602 , \20599 , \20600 , \20601 );
and \g454860/U$2 ( \20603 , \16317 , RIfc71a08_6315);
and \g454860/U$3 ( \20604 , RIfc718a0_6314, \16325 );
nor \g454860/U$1 ( \20605 , \20603 , \20604 );
not \g449919/U$3 ( \20606 , \20605 );
not \g449919/U$4 ( \20607 , \16311 );
and \g449919/U$2 ( \20608 , \20606 , \20607 );
and \g449919/U$5 ( \20609 , \16341 , RIfcae5c0_7006);
nor \g449919/U$1 ( \20610 , \20608 , \20609 );
and \g452490/U$2 ( \20611 , \16377 , RIfe8b1e8_7927);
and \g452490/U$3 ( \20612 , RIe202098_4313, \16313 );
nor \g452490/U$1 ( \20613 , \20611 , \20612 );
and \g451916/U$2 ( \20614 , \16334 , RIf161858_5569);
and \g451916/U$3 ( \20615 , RIfc62c60_6146, \16380 );
nor \g451916/U$1 ( \20616 , \20614 , \20615 );
nand \g447317/U$1 ( \20617 , \20602 , \20610 , \20613 , \20616 );
nor \g446015/U$1 ( \20618 , \20597 , \20598 , \20617 );
and \g452529/U$2 ( \20619 , \16364 , RIfc63200_6150);
and \g452529/U$3 ( \20620 , RIfe8b4b8_7929, \16368 );
nor \g452529/U$1 ( \20621 , \20619 , \20620 );
and \g451912/U$2 ( \20622 , \16361 , RIfc71198_6309);
and \g451912/U$3 ( \20623 , RIf15dbe0_5526, \16427 );
nor \g451912/U$1 ( \20624 , \20622 , \20623 );
and \g445161/U$2 ( \20625 , \20618 , \20621 , \20624 );
nor \g445161/U$1 ( \20626 , \20625 , \16393 );
or \g444214/U$1 ( \20627 , \20567 , \20596 , \20626 );
_DC \g3bb2/U$1 ( \20628 , \20627 , \16652 );
and \g446047/U$2 ( \20629 , RIe1e7ef0_4016, \16321 );
and \g446047/U$3 ( \20630 , RIe1e51f0_3984, \16313 );
and \g448942/U$2 ( \20631 , RIe1c35f0_3600, \16398 );
and \g448942/U$3 ( \20632 , \16341 , RIe1c62f0_3632);
and \g448942/U$4 ( \20633 , RIe1dcaf0_3888, \16485 );
nor \g448942/U$1 ( \20634 , \20631 , \20632 , \20633 );
and \g454500/U$2 ( \20635 , \16317 , RIe1ce9f0_3728);
and \g454500/U$3 ( \20636 , RIe1d16f0_3760, \16325 );
nor \g454500/U$1 ( \20637 , \20635 , \20636 );
not \g449958/U$3 ( \20638 , \20637 );
not \g449958/U$4 ( \20639 , \16351 );
and \g449958/U$2 ( \20640 , \20638 , \20639 );
and \g449958/U$5 ( \20641 , \16354 , RIe1df7f0_3920);
nor \g449958/U$1 ( \20642 , \20640 , \20641 );
and \g452039/U$2 ( \20643 , \16361 , RIe1bdbf0_3536);
and \g452039/U$3 ( \20644 , RIe1c08f0_3568, \16364 );
nor \g452039/U$1 ( \20645 , \20643 , \20644 );
and \g451006/U$2 ( \20646 , \16368 , RIe1c8ff0_3664);
and \g451006/U$3 ( \20647 , RIe1cbcf0_3696, \16371 );
nor \g451006/U$1 ( \20648 , \20646 , \20647 );
nand \g447698/U$1 ( \20649 , \20634 , \20642 , \20645 , \20648 );
nor \g446047/U$1 ( \20650 , \20629 , \20630 , \20649 );
and \g452038/U$2 ( \20651 , \16377 , RIe1e24f0_3952);
and \g452038/U$3 ( \20652 , RIe1d9df0_3856, \16380 );
nor \g452038/U$1 ( \20653 , \20651 , \20652 );
and \g452037/U$2 ( \20654 , \16334 , RIe1d70f0_3824);
and \g452037/U$3 ( \20655 , RIe1eabf0_4048, \16328 );
nor \g452037/U$1 ( \20656 , \20654 , \20655 );
and \g445185/U$2 ( \20657 , \20650 , \20653 , \20656 );
nor \g445185/U$1 ( \20658 , \20657 , \16555 );
and \g446049/U$2 ( \20659 , RIfe89a00_7910, \16427 );
and \g446049/U$3 ( \20660 , RIe1f2918_4137, \16368 );
and \g448943/U$2 ( \20661 , RIf1554e0_5430, \16485 );
and \g448943/U$3 ( \20662 , \16356 , RIfc5bd48_6067);
and \g448943/U$4 ( \20663 , RIfccc818_7349, \16398 );
nor \g448943/U$1 ( \20664 , \20661 , \20662 , \20663 );
and \g455403/U$2 ( \20665 , \16317 , RIfe89cd0_7912);
and \g455403/U$3 ( \20666 , RIf1588e8_5467, \16325 );
nor \g455403/U$1 ( \20667 , \20665 , \20666 );
not \g449961/U$3 ( \20668 , \20667 );
not \g449961/U$4 ( \20669 , \16311 );
and \g449961/U$2 ( \20670 , \20668 , \20669 );
and \g449961/U$5 ( \20671 , \16341 , RIf14f3d8_5361);
nor \g449961/U$1 ( \20672 , \20670 , \20671 );
and \g452047/U$2 ( \20673 , \16377 , RIe1f9c68_4219);
and \g452047/U$3 ( \20674 , RIfc5ba78_6065, \16313 );
nor \g452047/U$1 ( \20675 , \20673 , \20674 );
and \g452049/U$2 ( \20676 , \16334 , RIe1f4c40_4162);
and \g452049/U$3 ( \20677 , RIf154298_5417, \16380 );
nor \g452049/U$1 ( \20678 , \20676 , \20677 );
nand \g447325/U$1 ( \20679 , \20664 , \20672 , \20675 , \20678 );
nor \g446049/U$1 ( \20680 , \20659 , \20660 , \20679 );
and \g452044/U$2 ( \20681 , \16361 , RIe1ed620_4078);
and \g452044/U$3 ( \20682 , RIfe89b68_7911, \16432 );
nor \g452044/U$1 ( \20683 , \20681 , \20682 );
and \g452043/U$2 ( \20684 , \16364 , RIf14d920_5342);
and \g452043/U$3 ( \20685 , RIf150350_5372, \16371 );
nor \g452043/U$1 ( \20686 , \20684 , \20685 );
and \g445187/U$2 ( \20687 , \20680 , \20683 , \20686 );
nor \g445187/U$1 ( \20688 , \20687 , \16480 );
nor \g444670/U$1 ( \20689 , \20658 , \20688 );
and \g446835/U$2 ( \20690 , \18711 , RIfea7af0_8224);
and \g446835/U$3 ( \20691 , RIe176d18_2729, \18713 );
nor \g446835/U$1 ( \20692 , \20690 , \20691 );
not \g444412/U$2 ( \20693 , \20692 );
and \g452087/U$2 ( \20694 , \16377 , RIe197130_3096);
and \g452087/U$3 ( \20695 , RIe191730_3032, \16380 );
nor \g452087/U$1 ( \20696 , \20694 , \20695 );
and \g446060/U$2 ( \20697 , RIe199e30_3128, \16321 );
and \g446060/U$3 ( \20698 , RIf145388_5247, \16313 );
and \g448955/U$2 ( \20699 , RIe180930_2840, \16337 );
and \g448955/U$3 ( \20700 , \16341 , RIfcabcf8_6977);
and \g448955/U$4 ( \20701 , RIe194430_3064, \16485 );
nor \g448955/U$1 ( \20702 , \20699 , \20700 , \20701 );
and \g454468/U$2 ( \20703 , \16317 , RIe186330_2904);
and \g454468/U$3 ( \20704 , RIe189030_2936, \16325 );
nor \g454468/U$1 ( \20705 , \20703 , \20704 );
not \g449972/U$3 ( \20706 , \20705 );
not \g449972/U$4 ( \20707 , \16351 );
and \g449972/U$2 ( \20708 , \20706 , \20707 );
and \g449972/U$5 ( \20709 , \16354 , RIfe8a108_7915);
nor \g449972/U$1 ( \20710 , \20708 , \20709 );
and \g452090/U$2 ( \20711 , \16361 , RIe17af30_2776);
and \g452090/U$3 ( \20712 , RIe17dc30_2808, \16364 );
nor \g452090/U$1 ( \20713 , \20711 , \20712 );
and \g452089/U$2 ( \20714 , \16368 , RIe183630_2872);
and \g452089/U$3 ( \20715 , RIfc6c878_6257, \16371 );
nor \g452089/U$1 ( \20716 , \20714 , \20715 );
nand \g447704/U$1 ( \20717 , \20702 , \20710 , \20713 , \20716 );
nor \g446060/U$1 ( \20718 , \20697 , \20698 , \20717 );
and \g452641/U$2 ( \20719 , \16334 , RIe18ea30_3000);
and \g452641/U$3 ( \20720 , RIe19cb30_3160, \16326 );
nor \g452641/U$1 ( \20721 , \20719 , \20720 );
nand \g445589/U$1 ( \20722 , \20696 , \20718 , \20721 );
and \g444733/U$2 ( \20723 , \20722 , \17938 );
and \g448954/U$2 ( \20724 , RIfceec88_7739, \16321 );
and \g448954/U$3 ( \20725 , \16326 , RIfc6c2d8_6253);
and \g448954/U$4 ( \20726 , RIfe89730_7908, \16337 );
nor \g448954/U$1 ( \20727 , \20724 , \20725 , \20726 );
and \g454822/U$2 ( \20728 , \16317 , RIf163fb8_5597);
and \g454822/U$3 ( \20729 , RIf164dc8_5607, \16325 );
nor \g454822/U$1 ( \20730 , \20728 , \20729 );
not \g449970/U$3 ( \20731 , \20730 );
not \g449970/U$4 ( \20732 , \16330 );
and \g449970/U$2 ( \20733 , \20731 , \20732 );
and \g449970/U$5 ( \20734 , \16339 , RIf15c6c8_5511);
nor \g449970/U$1 ( \20735 , \20733 , \20734 );
and \g452082/U$2 ( \20736 , \16377 , RIe200748_4295);
and \g452082/U$3 ( \20737 , RIe201f30_4312, \16313 );
nor \g452082/U$1 ( \20738 , \20736 , \20737 );
and \g453396/U$2 ( \20739 , \16334 , RIfe895c8_7907);
and \g453396/U$3 ( \20740 , RIf163040_5586, \16380 );
nor \g453396/U$1 ( \20741 , \20739 , \20740 );
nand \g447330/U$1 ( \20742 , \20727 , \20735 , \20738 , \20741 );
and \g444733/U$3 ( \20743 , \16394 , \20742 );
nor \g444733/U$1 ( \20744 , \20723 , \20743 );
and \g446838/U$2 ( \20745 , \16419 , RIf1599c8_5479);
and \g446838/U$3 ( \20746 , RIf15a238_5485, \16422 );
nor \g446838/U$1 ( \20747 , \20745 , \20746 );
and \g446836/U$2 ( \20748 , \16429 , RIfe89898_7909);
and \g446836/U$3 ( \20749 , RIf15f968_5547, \16434 );
nor \g446836/U$1 ( \20750 , \20748 , \20749 );
and \g446837/U$2 ( \20751 , \16438 , RIe1fb5b8_4237);
and \g446837/U$3 ( \20752 , RIfe89460_7906, \16441 );
nor \g446837/U$1 ( \20753 , \20751 , \20752 );
nand \g444492/U$1 ( \20754 , \20744 , \20747 , \20750 , \20753 );
and \g446054/U$2 ( \20755 , RIfcccc50_7352, \16326 );
and \g446054/U$3 ( \20756 , RIfccb738_7337, \16334 );
and \g448950/U$2 ( \20757 , RIf16f250_5724, \16398 );
and \g448950/U$3 ( \20758 , \16339 , RIf16fd90_5732);
and \g448950/U$4 ( \20759 , RIfe89e38_7913, \16485 );
nor \g448950/U$1 ( \20760 , \20757 , \20758 , \20759 );
and \g454484/U$2 ( \20761 , \16317 , RIfcabb90_6976);
and \g454484/U$3 ( \20762 , RIfca9868_6951, \16325 );
nor \g454484/U$1 ( \20763 , \20761 , \20762 );
not \g449967/U$3 ( \20764 , \20763 );
not \g449967/U$4 ( \20765 , \16351 );
and \g449967/U$2 ( \20766 , \20764 , \20765 );
and \g449967/U$5 ( \20767 , \16356 , RIfe89fa0_7914);
nor \g449967/U$1 ( \20768 , \20766 , \20767 );
and \g452070/U$2 ( \20769 , \16361 , RIfcaba28_6975);
and \g452070/U$3 ( \20770 , RIfc6c440_6254, \16364 );
nor \g452070/U$1 ( \20771 , \20769 , \20770 );
and \g452069/U$2 ( \20772 , \16368 , RIe172f38_2685);
and \g452069/U$3 ( \20773 , RIfca99d0_6952, \16371 );
nor \g452069/U$1 ( \20774 , \20772 , \20773 );
nand \g447701/U$1 ( \20775 , \20760 , \20768 , \20771 , \20774 );
nor \g446054/U$1 ( \20776 , \20755 , \20756 , \20775 );
and \g452066/U$2 ( \20777 , \16380 , RIfcdd078_7537);
and \g452066/U$3 ( \20778 , RIfcccdb8_7353, \16321 );
nor \g452066/U$1 ( \20779 , \20777 , \20778 );
and \g445503/U$2 ( \20780 , \20776 , \20779 );
nor \g445503/U$1 ( \20781 , \20780 , \16649 );
and \g446057/U$2 ( \20782 , RIe212088_4495, \16427 );
and \g446057/U$3 ( \20783 , RIe20f388_4463, \16368 );
and \g448951/U$2 ( \20784 , RIe222e88_4687, \16321 );
and \g448951/U$3 ( \20785 , \16326 , RIfc40610_5758);
and \g448951/U$4 ( \20786 , RIe20c688_4431, \16337 );
nor \g448951/U$1 ( \20787 , \20784 , \20785 , \20786 );
and \g454608/U$2 ( \20788 , \16317 , RIe21d488_4623);
and \g454608/U$3 ( \20789 , RIfcab758_6973, \16325 );
nor \g454608/U$1 ( \20790 , \20788 , \20789 );
not \g449968/U$3 ( \20791 , \20790 );
not \g449968/U$4 ( \20792 , \16330 );
and \g449968/U$2 ( \20793 , \20791 , \20792 );
and \g449968/U$5 ( \20794 , \16341 , RIf167ac8_5639);
nor \g449968/U$1 ( \20795 , \20793 , \20794 );
and \g452077/U$2 ( \20796 , \16377 , RIe220188_4655);
and \g452077/U$3 ( \20797 , RIfc5d260_6082, \16313 );
nor \g452077/U$1 ( \20798 , \20796 , \20797 );
and \g452080/U$2 ( \20799 , \16334 , RIe214d88_4527);
and \g452080/U$3 ( \20800 , RIe217a88_4559, \16380 );
nor \g452080/U$1 ( \20801 , \20799 , \20800 );
nand \g447329/U$1 ( \20802 , \20787 , \20795 , \20798 , \20801 );
nor \g446057/U$1 ( \20803 , \20782 , \20783 , \20802 );
and \g452075/U$2 ( \20804 , \16361 , RIe206c88_4367);
and \g452075/U$3 ( \20805 , RIfe892f8_7905, \16432 );
nor \g452075/U$1 ( \20806 , \20804 , \20805 );
and \g452074/U$2 ( \20807 , \16364 , RIe209988_4399);
and \g452074/U$3 ( \20808 , RIf168a40_5650, \16371 );
nor \g452074/U$1 ( \20809 , \20807 , \20808 );
and \g445192/U$2 ( \20810 , \20803 , \20806 , \20809 );
nor \g445192/U$1 ( \20811 , \20810 , \16389 );
nor \g444412/U$1 ( \20812 , \20693 , \20754 , \20781 , \20811 );
and \g452056/U$2 ( \20813 , \16361 , RIe1703a0_2654);
and \g452056/U$3 ( \20814 , RIe1fdfe8_4267, \16427 );
nor \g452056/U$1 ( \20815 , \20813 , \20814 );
and \g446053/U$2 ( \20816 , RIe203f88_4335, \16448 );
and \g446053/U$3 ( \20817 , RIe1f73a0_4190, \16371 );
and \g448947/U$2 ( \20818 , RIe178230_2744, \16485 );
and \g448947/U$3 ( \20819 , \16356 , RIe18bd30_2968);
and \g448947/U$4 ( \20820 , RIe1baef0_3504, \16337 );
nor \g448947/U$1 ( \20821 , \20818 , \20819 , \20820 );
and \g455285/U$2 ( \20822 , \16317 , RIe1a5230_3256);
and \g455285/U$3 ( \20823 , RIe1a7f30_3288, \16325 );
nor \g455285/U$1 ( \20824 , \20822 , \20823 );
not \g449964/U$3 ( \20825 , \20824 );
not \g449964/U$4 ( \20826 , \16311 );
and \g449964/U$2 ( \20827 , \20825 , \20826 );
and \g449964/U$5 ( \20828 , \16341 , RIe1d43f0_3792);
nor \g449964/U$1 ( \20829 , \20827 , \20828 );
and \g452058/U$2 ( \20830 , \16377 , RIe19f830_3192);
and \g452058/U$3 ( \20831 , RIe1a2530_3224, \16313 );
nor \g452058/U$1 ( \20832 , \20830 , \20831 );
and \g452060/U$2 ( \20833 , \16334 , RIe21a788_4591);
and \g452060/U$3 ( \20834 , RIe225b88_4719, \16380 );
nor \g452060/U$1 ( \20835 , \20833 , \20834 );
nand \g447327/U$1 ( \20836 , \20821 , \20829 , \20832 , \20835 );
nor \g446053/U$1 ( \20837 , \20816 , \20817 , \20836 );
and \g452055/U$2 ( \20838 , \16364 , RIe1add68_3355);
and \g452055/U$3 ( \20839 , RIe1efee8_4107, \16368 );
nor \g452055/U$1 ( \20840 , \20838 , \20839 );
nand \g445588/U$1 ( \20841 , \20815 , \20837 , \20840 );
and \g444671/U$2 ( \20842 , \20841 , \16752 );
and \g452051/U$2 ( \20843 , \16361 , RIe1aa528_3315);
and \g452051/U$3 ( \20844 , RIfccdd30_7364, \16427 );
nor \g452051/U$1 ( \20845 , \20843 , \20844 );
and \g446051/U$2 ( \20846 , RIf148a60_5286, \16448 );
and \g446051/U$3 ( \20847 , RIe1b2250_3404, \16371 );
and \g448946/U$2 ( \20848 , RIf1499d8_5297, \16344 );
and \g448946/U$3 ( \20849 , \16356 , RIfcac298_6981);
and \g448946/U$4 ( \20850 , RIfc54728_5983, \16337 );
nor \g448946/U$1 ( \20851 , \20848 , \20849 , \20850 );
and \g454711/U$2 ( \20852 , \16317 , RIf14b058_5313);
and \g454711/U$3 ( \20853 , RIfc680c0_6206, \16325 );
nor \g454711/U$1 ( \20854 , \20852 , \20853 );
not \g449962/U$3 ( \20855 , \20854 );
not \g449962/U$4 ( \20856 , \16311 );
and \g449962/U$2 ( \20857 , \20855 , \20856 );
and \g449962/U$5 ( \20858 , \16339 , RIfc6e768_6279);
nor \g449962/U$1 ( \20859 , \20857 , \20858 );
and \g452376/U$2 ( \20860 , \16377 , RIe1b6b70_3456);
and \g452376/U$3 ( \20861 , RIe1b8bc8_3479, \16313 );
nor \g452376/U$1 ( \20862 , \20860 , \20861 );
and \g452052/U$2 ( \20863 , \16334 , RIfec19c8_8323);
and \g452052/U$3 ( \20864 , RIfe89190_7904, \16380 );
nor \g452052/U$1 ( \20865 , \20863 , \20864 );
nand \g447326/U$1 ( \20866 , \20851 , \20859 , \20862 , \20865 );
nor \g446051/U$1 ( \20867 , \20846 , \20847 , \20866 );
and \g453393/U$2 ( \20868 , \16364 , RIe1abfe0_3334);
and \g453393/U$3 ( \20869 , RIfec1860_8322, \16368 );
nor \g453393/U$1 ( \20870 , \20868 , \20869 );
nand \g445587/U$1 ( \20871 , \20845 , \20867 , \20870 );
and \g444671/U$3 ( \20872 , \16477 , \20871 );
nor \g444671/U$1 ( \20873 , \20842 , \20872 );
nand \g444285/U$1 ( \20874 , \20689 , \20812 , \20873 );
_DC \g3c37/U$1 ( \20875 , \20874 , \16652 );
and \g451521/U$2 ( \20876 , \16380 , RIe217920_4558);
and \g451521/U$3 ( \20877 , RIe222d20_4686, \16321 );
nor \g451521/U$1 ( \20878 , \20876 , \20877 );
and \g445918/U$2 ( \20879 , RIfc404a8_5757, \16328 );
and \g445918/U$3 ( \20880 , RIe220020_4654, \16377 );
and \g448772/U$2 ( \20881 , RIe20c520_4430, \16398 );
and \g448772/U$3 ( \20882 , \16341 , RIfe8e758_7965);
and \g448772/U$4 ( \20883 , RIe21d320_4622, \16344 );
nor \g448772/U$1 ( \20884 , \20881 , \20882 , \20883 );
and \g454611/U$2 ( \20885 , \16317 , RIe211f20_4494);
and \g454611/U$3 ( \20886 , RIfc5b910_6064, \16325 );
nor \g454611/U$1 ( \20887 , \20885 , \20886 );
not \g449800/U$3 ( \20888 , \20887 );
not \g449800/U$4 ( \20889 , \16351 );
and \g449800/U$2 ( \20890 , \20888 , \20889 );
and \g449800/U$5 ( \20891 , \16356 , RIf16a930_5672);
nor \g449800/U$1 ( \20892 , \20890 , \20891 );
and \g451525/U$2 ( \20893 , \16361 , RIe206b20_4366);
and \g451525/U$3 ( \20894 , RIe209820_4398, \16364 );
nor \g451525/U$1 ( \20895 , \20893 , \20894 );
and \g451524/U$2 ( \20896 , \16368 , RIe20f220_4462);
and \g451524/U$3 ( \20897 , RIfe8e8c0_7966, \16371 );
nor \g451524/U$1 ( \20898 , \20896 , \20897 );
nand \g447608/U$1 ( \20899 , \20884 , \20892 , \20895 , \20898 );
nor \g445918/U$1 ( \20900 , \20879 , \20880 , \20899 );
and \g451523/U$2 ( \20901 , \16334 , RIe214c20_4526);
and \g451523/U$3 ( \20902 , RIf16b8a8_5683, \16313 );
nor \g451523/U$1 ( \20903 , \20901 , \20902 );
nand \g445555/U$1 ( \20904 , \20878 , \20900 , \20903 );
and \g444898/U$2 ( \20905 , \20904 , \16390 );
and \g448769/U$2 ( \20906 , RIf15da78_5525, \16427 );
and \g448769/U$3 ( \20907 , \16448 , RIf15f800_5546);
and \g448769/U$4 ( \20908 , RIf163e50_5596, \16485 );
nor \g448769/U$1 ( \20909 , \20906 , \20907 , \20908 );
and \g454564/U$2 ( \20910 , \16317 , RIf15b048_5495);
and \g454564/U$3 ( \20911 , RIf15c560_5510, \16325 );
nor \g454564/U$1 ( \20912 , \20910 , \20911 );
not \g454563/U$1 ( \20913 , \20912 );
and \g449798/U$2 ( \20914 , \20913 , \16336 );
and \g449798/U$3 ( \20915 , RIf164c60_5606, \16354 );
nor \g449798/U$1 ( \20916 , \20914 , \20915 );
and \g451950/U$2 ( \20917 , \16361 , RIf159860_5478);
and \g451950/U$3 ( \20918 , RIfc62828_6143, \16364 );
nor \g451950/U$1 ( \20919 , \20917 , \20918 );
and \g451976/U$2 ( \20920 , \16368 , RIfe8dc18_7957);
and \g451976/U$3 ( \20921 , RIfe8d948_7955, \16371 );
nor \g451976/U$1 ( \20922 , \20920 , \20921 );
nand \g448042/U$1 ( \20923 , \20909 , \20916 , \20919 , \20922 );
and \g444898/U$3 ( \20924 , \16394 , \20923 );
nor \g444898/U$1 ( \20925 , \20905 , \20924 );
and \g446704/U$2 ( \20926 , \16705 , RIf1616f0_5568);
and \g446704/U$3 ( \20927 , RIf162ed8_5585, \16707 );
nor \g446704/U$1 ( \20928 , \20926 , \20927 );
and \g446703/U$2 ( \20929 , \16710 , RIf165a70_5616);
and \g446703/U$3 ( \20930 , RIf166b50_5628, \16712 );
nor \g446703/U$1 ( \20931 , \20929 , \20930 );
and \g446705/U$2 ( \20932 , \16715 , RIfe8dab0_7956);
and \g446705/U$3 ( \20933 , RIfe8dd80_7958, \16717 );
nor \g446705/U$1 ( \20934 , \20932 , \20933 );
nand \g444582/U$1 ( \20935 , \20925 , \20928 , \20931 , \20934 );
and \g451537/U$2 ( \20936 , \16364 , RIf14d7b8_5341);
and \g451537/U$3 ( \20937 , RIf1501e8_5371, \16371 );
nor \g451537/U$1 ( \20938 , \20936 , \20937 );
and \g445920/U$2 ( \20939 , RIf151700_5386, \16427 );
and \g445920/U$3 ( \20940 , RIe1f27b0_4136, \16368 );
and \g448776/U$2 ( \20941 , RIfc61748_6131, \16485 );
and \g448776/U$3 ( \20942 , \16356 , RIfc61e50_6136);
and \g448776/U$4 ( \20943 , RIfc7b620_6426, \16398 );
nor \g448776/U$1 ( \20944 , \20941 , \20942 , \20943 );
and \g454737/U$2 ( \20945 , \16317 , RIf157538_5453);
and \g454737/U$3 ( \20946 , RIf158780_5466, \16325 );
nor \g454737/U$1 ( \20947 , \20945 , \20946 );
not \g449804/U$3 ( \20948 , \20947 );
not \g449804/U$4 ( \20949 , \16311 );
and \g449804/U$2 ( \20950 , \20948 , \20949 );
and \g449804/U$5 ( \20951 , \16341 , RIfc60ed8_6125);
nor \g449804/U$1 ( \20952 , \20950 , \20951 );
and \g451542/U$2 ( \20953 , \16377 , RIe1f9b00_4218);
and \g451542/U$3 ( \20954 , RIfca6e38_6921, \16313 );
nor \g451542/U$1 ( \20955 , \20953 , \20954 );
and \g451543/U$2 ( \20956 , \16334 , RIe1f4ad8_4161);
and \g451543/U$3 ( \20957 , RIf154130_5416, \16380 );
nor \g451543/U$1 ( \20958 , \20956 , \20957 );
nand \g447287/U$1 ( \20959 , \20944 , \20952 , \20955 , \20958 );
nor \g445920/U$1 ( \20960 , \20939 , \20940 , \20959 );
and \g451538/U$2 ( \20961 , \16361 , RIe1ed4b8_4077);
and \g451538/U$3 ( \20962 , RIf152ab0_5400, \16448 );
nor \g451538/U$1 ( \20963 , \20961 , \20962 );
nand \g445557/U$1 ( \20964 , \20938 , \20960 , \20963 );
and \g444833/U$2 ( \20965 , \20964 , \16481 );
and \g448774/U$2 ( \20966 , RIf146030_5256, \16398 );
and \g448774/U$3 ( \20967 , \16341 , RIf146e40_5266);
and \g448774/U$4 ( \20968 , RIfc44fa8_5807, \16344 );
nor \g448774/U$1 ( \20969 , \20966 , \20967 , \20968 );
and \g454585/U$2 ( \20970 , \16317 , RIf147818_5273);
and \g454585/U$3 ( \20971 , RIf1488f8_5285, \16325 );
nor \g454585/U$1 ( \20972 , \20970 , \20971 );
not \g449801/U$3 ( \20973 , \20972 );
not \g449801/U$4 ( \20974 , \16351 );
and \g449801/U$2 ( \20975 , \20973 , \20974 );
and \g449801/U$5 ( \20976 , \16356 , RIfcbd638_7177);
nor \g449801/U$1 ( \20977 , \20975 , \20976 );
and \g451534/U$2 ( \20978 , \16361 , RIfe8e320_7962);
and \g451534/U$3 ( \20979 , RIfe8dee8_7959, \16364 );
nor \g451534/U$1 ( \20980 , \20978 , \20979 );
and \g451532/U$2 ( \20981 , \16368 , RIfe8e488_7963);
and \g451532/U$3 ( \20982 , RIfe8e050_7960, \16371 );
nor \g451532/U$1 ( \20983 , \20981 , \20982 );
nand \g447609/U$1 ( \20984 , \20969 , \20977 , \20980 , \20983 );
and \g444833/U$3 ( \20985 , \16477 , \20984 );
nor \g444833/U$1 ( \20986 , \20965 , \20985 );
and \g446709/U$2 ( \20987 , \18268 , RIfc5ea48_6099);
and \g446709/U$3 ( \20988 , RIfca4de0_6898, \18270 );
nor \g446709/U$1 ( \20989 , \20987 , \20988 );
and \g446710/U$2 ( \20990 , \18273 , RIe1b6a08_3455);
and \g446710/U$3 ( \20991 , RIe1b8a60_3478, \18275 );
nor \g446710/U$1 ( \20992 , \20990 , \20991 );
and \g446711/U$2 ( \20993 , \18278 , RIfe8e1b8_7961);
and \g446711/U$3 ( \20994 , RIfe8e5f0_7964, \18280 );
nor \g446711/U$1 ( \20995 , \20993 , \20994 );
nand \g444583/U$1 ( \20996 , \20986 , \20989 , \20992 , \20995 );
and \g445912/U$2 ( \20997 , RIe1eaa88_4047, \16328 );
and \g445912/U$3 ( \20998 , RIe1e2388_3951, \16377 );
and \g448764/U$2 ( \20999 , RIe1ce888_3727, \16427 );
and \g448764/U$3 ( \21000 , \16448 , RIe1d1588_3759);
and \g448764/U$4 ( \21001 , RIe1dc988_3887, \16485 );
nor \g448764/U$1 ( \21002 , \20999 , \21000 , \21001 );
and \g454552/U$2 ( \21003 , \16317 , RIe1c3488_3599);
and \g454552/U$3 ( \21004 , RIe1c6188_3631, \16325 );
nor \g454552/U$1 ( \21005 , \21003 , \21004 );
not \g454551/U$1 ( \21006 , \21005 );
and \g449794/U$2 ( \21007 , \21006 , \16336 );
and \g449794/U$3 ( \21008 , RIe1df688_3919, \16356 );
nor \g449794/U$1 ( \21009 , \21007 , \21008 );
and \g451500/U$2 ( \21010 , \16361 , RIe1bda88_3535);
and \g451500/U$3 ( \21011 , RIe1c0788_3567, \16364 );
nor \g451500/U$1 ( \21012 , \21010 , \21011 );
and \g451498/U$2 ( \21013 , \16368 , RIe1c8e88_3663);
and \g451498/U$3 ( \21014 , RIe1cbb88_3695, \16371 );
nor \g451498/U$1 ( \21015 , \21013 , \21014 );
nand \g448041/U$1 ( \21016 , \21002 , \21009 , \21012 , \21015 );
nor \g445912/U$1 ( \21017 , \20997 , \20998 , \21016 );
and \g451494/U$2 ( \21018 , \16334 , RIe1d6f88_3823);
and \g451494/U$3 ( \21019 , RIe1e5088_3983, \16313 );
nor \g451494/U$1 ( \21020 , \21018 , \21019 );
and \g451493/U$2 ( \21021 , \16380 , RIe1d9c88_3855);
and \g451493/U$3 ( \21022 , RIe1e7d88_4015, \16321 );
nor \g451493/U$1 ( \21023 , \21021 , \21022 );
and \g445083/U$2 ( \21024 , \21017 , \21020 , \21023 );
nor \g445083/U$1 ( \21025 , \21024 , \16555 );
and \g445914/U$2 ( \21026 , RIe1fde80_4266, \16427 );
and \g445914/U$3 ( \21027 , RIe1efd80_4106, \16368 );
and \g448766/U$2 ( \21028 , RIe1780c8_2743, \16485 );
and \g448766/U$3 ( \21029 , \16354 , RIe18bbc8_2967);
and \g448766/U$4 ( \21030 , RIe1bad88_3503, \16398 );
nor \g448766/U$1 ( \21031 , \21028 , \21029 , \21030 );
and \g454456/U$2 ( \21032 , \16317 , RIe1a50c8_3255);
and \g454456/U$3 ( \21033 , RIe1a7dc8_3287, \16325 );
nor \g454456/U$1 ( \21034 , \21032 , \21033 );
not \g449996/U$3 ( \21035 , \21034 );
not \g449996/U$4 ( \21036 , \16311 );
and \g449996/U$2 ( \21037 , \21035 , \21036 );
and \g449996/U$5 ( \21038 , \16339 , RIe1d4288_3791);
nor \g449996/U$1 ( \21039 , \21037 , \21038 );
and \g451508/U$2 ( \21040 , \16377 , RIe19f6c8_3191);
and \g451508/U$3 ( \21041 , RIe1a23c8_3223, \16313 );
nor \g451508/U$1 ( \21042 , \21040 , \21041 );
and \g451510/U$2 ( \21043 , \16334 , RIe21a620_4590);
and \g451510/U$3 ( \21044 , RIe225a20_4718, \16380 );
nor \g451510/U$1 ( \21045 , \21043 , \21044 );
nand \g447286/U$1 ( \21046 , \21031 , \21039 , \21042 , \21045 );
nor \g445914/U$1 ( \21047 , \21026 , \21027 , \21046 );
and \g451504/U$2 ( \21048 , \16361 , RIe170238_2653);
and \g451504/U$3 ( \21049 , RIe203e20_4334, \16432 );
nor \g451504/U$1 ( \21050 , \21048 , \21049 );
and \g451503/U$2 ( \21051 , \16364 , RIe1adc00_3354);
and \g451503/U$3 ( \21052 , RIe1f7238_4189, \16371 );
nor \g451503/U$1 ( \21053 , \21051 , \21052 );
and \g445087/U$2 ( \21054 , \21047 , \21050 , \21053 );
nor \g445087/U$1 ( \21055 , \21054 , \16586 );
or \g444351/U$1 ( \21056 , \20935 , \20996 , \21025 , \21055 );
and \g445909/U$2 ( \21057 , RIe188ec8_2935, \16448 );
and \g445909/U$3 ( \21058 , RIfc68228_6207, \16371 );
and \g449179/U$2 ( \21059 , RIe199cc8_3127, \16321 );
and \g449179/U$3 ( \21060 , \16326 , RIe19c9c8_3159);
and \g449179/U$4 ( \21061 , RIe1807c8_2839, \16398 );
nor \g449179/U$1 ( \21062 , \21059 , \21060 , \21061 );
and \g455204/U$2 ( \21063 , \16317 , RIe1942c8_3063);
and \g455204/U$3 ( \21064 , RIfec20d0_8328, \16325 );
nor \g455204/U$1 ( \21065 , \21063 , \21064 );
not \g449789/U$3 ( \21066 , \21065 );
not \g449789/U$4 ( \21067 , \16330 );
and \g449789/U$2 ( \21068 , \21066 , \21067 );
and \g449789/U$5 ( \21069 , \16341 , RIfccb5d0_7336);
nor \g449789/U$1 ( \21070 , \21068 , \21069 );
and \g453191/U$2 ( \21071 , \16377 , RIe196fc8_3095);
and \g453191/U$3 ( \21072 , RIfe8ea28_7967, \16313 );
nor \g453191/U$1 ( \21073 , \21071 , \21072 );
and \g453149/U$2 ( \21074 , \16334 , RIe18e8c8_2999);
and \g453149/U$3 ( \21075 , RIe1915c8_3031, \16380 );
nor \g453149/U$1 ( \21076 , \21074 , \21075 );
nand \g447284/U$1 ( \21077 , \21062 , \21070 , \21073 , \21076 );
nor \g445909/U$1 ( \21078 , \21057 , \21058 , \21077 );
and \g451481/U$2 ( \21079 , \16364 , RIe17dac8_2807);
and \g451481/U$3 ( \21080 , RIe1834c8_2871, \16368 );
nor \g451481/U$1 ( \21081 , \21079 , \21080 );
and \g451482/U$2 ( \21082 , \16361 , RIe17adc8_2775);
and \g451482/U$3 ( \21083 , RIe1861c8_2903, \16427 );
nor \g451482/U$1 ( \21084 , \21082 , \21083 );
and \g445081/U$2 ( \21085 , \21078 , \21081 , \21084 );
nor \g445081/U$1 ( \21086 , \21085 , \16618 );
and \g445910/U$2 ( \21087 , RIee3bce0_5139, \16448 );
and \g445910/U$3 ( \21088 , RIee39850_5113, \16371 );
and \g448762/U$2 ( \21089 , RIf140900_5194, \16321 );
and \g448762/U$3 ( \21090 , \16328 , RIf141e18_5209);
and \g448762/U$4 ( \21091 , RIf16f0e8_5723, \16398 );
nor \g448762/U$1 ( \21092 , \21089 , \21090 , \21091 );
and \g455305/U$2 ( \21093 , \16317 , RIf13ece0_5174);
and \g455305/U$3 ( \21094 , RIf13f988_5183, \16325 );
nor \g455305/U$1 ( \21095 , \21093 , \21094 );
not \g449792/U$3 ( \21096 , \21095 );
not \g449792/U$4 ( \21097 , \16330 );
and \g449792/U$2 ( \21098 , \21096 , \21097 );
and \g449792/U$5 ( \21099 , \16341 , RIf16fc28_5731);
nor \g449792/U$1 ( \21100 , \21098 , \21099 );
and \g451490/U$2 ( \21101 , \16377 , RIe1753c8_2711);
and \g451490/U$3 ( \21102 , RIf140090_5188, \16313 );
nor \g451490/U$1 ( \21103 , \21101 , \21102 );
and \g452803/U$2 ( \21104 , \16334 , RIee3cf28_5152);
and \g452803/U$3 ( \21105 , RIee3e170_5165, \16380 );
nor \g452803/U$1 ( \21106 , \21104 , \21105 );
nand \g447285/U$1 ( \21107 , \21092 , \21100 , \21103 , \21106 );
nor \g445910/U$1 ( \21108 , \21087 , \21088 , \21107 );
and \g451488/U$2 ( \21109 , \16364 , RIf16dd38_5709);
and \g451488/U$3 ( \21110 , RIe172dd0_2684, \16368 );
nor \g451488/U$1 ( \21111 , \21109 , \21110 );
and \g451489/U$2 ( \21112 , \16361 , RIfce9120_7674);
and \g451489/U$3 ( \21113 , RIee3ac00_5127, \16427 );
nor \g451489/U$1 ( \21114 , \21112 , \21113 );
and \g445082/U$2 ( \21115 , \21108 , \21111 , \21114 );
nor \g445082/U$1 ( \21116 , \21115 , \16649 );
or \g444272/U$1 ( \21117 , \21056 , \21086 , \21116 );
_DC \g3cbc/U$1 ( \21118 , \21117 , \16652 );
and \g451692/U$2 ( \21119 , \16361 , RIfec1c98_8325);
and \g451692/U$3 ( \21120 , RIf1476b0_5272, \16427 );
nor \g451692/U$1 ( \21121 , \21119 , \21120 );
and \g445957/U$2 ( \21122 , RIf148790_5284, \16432 );
and \g445957/U$3 ( \21123 , RIfe8ba58_7933, \16371 );
and \g448825/U$2 ( \21124 , RIfc4ebc0_5918, \16344 );
and \g448825/U$3 ( \21125 , \16356 , RIfcd4db0_7444);
and \g448825/U$4 ( \21126 , RIfcb8e80_7126, \16398 );
nor \g448825/U$1 ( \21127 , \21124 , \21125 , \21126 );
and \g454405/U$2 ( \21128 , \16317 , RIf14aef0_5312);
and \g454405/U$3 ( \21129 , RIf14c2a0_5326, \16325 );
nor \g454405/U$1 ( \21130 , \21128 , \21129 );
not \g449852/U$3 ( \21131 , \21130 );
not \g449852/U$4 ( \21132 , \16311 );
and \g449852/U$2 ( \21133 , \21131 , \21132 );
and \g449852/U$5 ( \21134 , \16341 , RIfc4e788_5915);
nor \g449852/U$1 ( \21135 , \21133 , \21134 );
and \g451694/U$2 ( \21136 , \16377 , RIe1b68a0_3454);
and \g451694/U$3 ( \21137 , RIe1b88f8_3477, \16313 );
nor \g451694/U$1 ( \21138 , \21136 , \21137 );
and \g451695/U$2 ( \21139 , \16334 , RIfe8bd28_7935);
and \g451695/U$3 ( \21140 , RIfec1e00_8326, \16380 );
nor \g451695/U$1 ( \21141 , \21139 , \21140 );
nand \g447300/U$1 ( \21142 , \21127 , \21135 , \21138 , \21141 );
nor \g445957/U$1 ( \21143 , \21122 , \21123 , \21142 );
and \g451691/U$2 ( \21144 , \16364 , RIfe8bbc0_7934);
and \g451691/U$3 ( \21145 , RIfec1b30_8324, \16368 );
nor \g451691/U$1 ( \21146 , \21144 , \21145 );
nand \g445569/U$1 ( \21147 , \21121 , \21143 , \21146 );
and \g444912/U$2 ( \21148 , \21147 , \16477 );
and \g448822/U$2 ( \21149 , RIe1a4f60_3254, \16321 );
and \g448822/U$3 ( \21150 , \16344 , RIe177f60_2742);
and \g448822/U$4 ( \21151 , RIe18ba60_2966, \16356 );
nor \g448822/U$1 ( \21152 , \21149 , \21150 , \21151 );
and \g451094/U$2 ( \21153 , \16368 , RIe1efc18_4105);
and \g451094/U$3 ( \21154 , RIe1f70d0_4188, \16371 );
nor \g451094/U$1 ( \21155 , \21153 , \21154 );
and \g454643/U$2 ( \21156 , \16317 , RIe1fdd18_4265);
and \g454643/U$3 ( \21157 , RIe203cb8_4333, \16325 );
nor \g454643/U$1 ( \21158 , \21156 , \21157 );
not \g449849/U$3 ( \21159 , \21158 );
not \g449849/U$4 ( \21160 , \16351 );
and \g449849/U$2 ( \21161 , \21159 , \21160 );
and \g449849/U$5 ( \21162 , \16328 , RIe1a7c60_3286);
nor \g449849/U$1 ( \21163 , \21161 , \21162 );
and \g451687/U$2 ( \21164 , \16334 , RIe21a4b8_4589);
and \g451687/U$3 ( \21165 , RIe2258b8_4717, \16380 );
nor \g451687/U$1 ( \21166 , \21164 , \21165 );
nand \g447632/U$1 ( \21167 , \21152 , \21155 , \21163 , \21166 );
and \g444912/U$3 ( \21168 , \16752 , \21167 );
nor \g444912/U$1 ( \21169 , \21148 , \21168 );
and \g446751/U$2 ( \21170 , \17027 , RIe1bac20_3502);
and \g446751/U$3 ( \21171 , RIe1d4120_3790, \17034 );
nor \g446751/U$1 ( \21172 , \21170 , \21171 );
and \g446750/U$2 ( \21173 , \17779 , RIe19f560_3190);
and \g446750/U$3 ( \21174 , RIe1a2260_3222, \17781 );
nor \g446750/U$1 ( \21175 , \21173 , \21174 );
and \g446752/U$2 ( \21176 , \16774 , RIe1700d0_2652);
and \g446752/U$3 ( \21177 , RIe1ada98_3353, \16776 );
nor \g446752/U$1 ( \21178 , \21176 , \21177 );
nand \g444590/U$1 ( \21179 , \21169 , \21172 , \21175 , \21178 );
and \g451682/U$2 ( \21180 , \16361 , RIfe8c160_7938);
and \g451682/U$3 ( \21181 , RIf151598_5385, \16427 );
nor \g451682/U$1 ( \21182 , \21180 , \21181 );
and \g445955/U$2 ( \21183 , RIf152948_5399, \16448 );
and \g445955/U$3 ( \21184 , RIf150080_5370, \16371 );
and \g448820/U$2 ( \21185 , RIf1573d0_5452, \16321 );
and \g448820/U$3 ( \21186 , \16328 , RIf158618_5465);
and \g448820/U$4 ( \21187 , RIfc503a8_5935, \16337 );
nor \g448820/U$1 ( \21188 , \21185 , \21186 , \21187 );
and \g454638/U$2 ( \21189 , \16317 , RIf155378_5429);
and \g454638/U$3 ( \21190 , RIf155eb8_5437, \16325 );
nor \g454638/U$1 ( \21191 , \21189 , \21190 );
not \g449847/U$3 ( \21192 , \21191 );
not \g449847/U$4 ( \21193 , \16330 );
and \g449847/U$2 ( \21194 , \21192 , \21193 );
and \g449847/U$5 ( \21195 , \16339 , RIf14f270_5360);
nor \g449847/U$1 ( \21196 , \21194 , \21195 );
and \g451334/U$2 ( \21197 , \16377 , RIfec1f68_8327);
and \g451334/U$3 ( \21198 , RIf156b60_5446, \16313 );
nor \g451334/U$1 ( \21199 , \21197 , \21198 );
and \g451685/U$2 ( \21200 , \16334 , RIfe8bff8_7937);
and \g451685/U$3 ( \21201 , RIf153fc8_5415, \16380 );
nor \g451685/U$1 ( \21202 , \21200 , \21201 );
nand \g447298/U$1 ( \21203 , \21188 , \21196 , \21199 , \21202 );
nor \g445955/U$1 ( \21204 , \21183 , \21184 , \21203 );
and \g451411/U$2 ( \21205 , \16364 , RIf14d650_5340);
and \g451411/U$3 ( \21206 , RIfe8c2c8_7939, \16368 );
nor \g451411/U$1 ( \21207 , \21205 , \21206 );
nand \g445567/U$1 ( \21208 , \21182 , \21204 , \21207 );
and \g444825/U$2 ( \21209 , \21208 , \16481 );
and \g448818/U$2 ( \21210 , RIe1ce720_3726, \16427 );
and \g448818/U$3 ( \21211 , \16448 , RIe1d1420_3758);
and \g448818/U$4 ( \21212 , RIe1dc820_3886, \16485 );
nor \g448818/U$1 ( \21213 , \21210 , \21211 , \21212 );
and \g454399/U$2 ( \21214 , \16317 , RIe1c3320_3598);
and \g454399/U$3 ( \21215 , RIe1c6020_3630, \16325 );
nor \g454399/U$1 ( \21216 , \21214 , \21215 );
not \g454398/U$1 ( \21217 , \21216 );
and \g449845/U$2 ( \21218 , \21217 , \16336 );
and \g449845/U$3 ( \21219 , RIe1df520_3918, \16356 );
nor \g449845/U$1 ( \21220 , \21218 , \21219 );
and \g451680/U$2 ( \21221 , \16361 , RIe1bd920_3534);
and \g451680/U$3 ( \21222 , RIe1c0620_3566, \16364 );
nor \g451680/U$1 ( \21223 , \21221 , \21222 );
and \g451679/U$2 ( \21224 , \16368 , RIe1c8d20_3662);
and \g451679/U$3 ( \21225 , RIe1cba20_3694, \16371 );
nor \g451679/U$1 ( \21226 , \21224 , \21225 );
nand \g448050/U$1 ( \21227 , \21213 , \21220 , \21223 , \21226 );
and \g444825/U$3 ( \21228 , \16750 , \21227 );
nor \g444825/U$1 ( \21229 , \21209 , \21228 );
and \g446741/U$2 ( \21230 , \19457 , RIe1e7c20_4014);
and \g446741/U$3 ( \21231 , RIe1ea920_4046, \19459 );
nor \g446741/U$1 ( \21232 , \21230 , \21231 );
and \g446743/U$2 ( \21233 , \19462 , RIe1d6e20_3822);
and \g446743/U$3 ( \21234 , RIe1d9b20_3854, \19464 );
nor \g446743/U$1 ( \21235 , \21233 , \21234 );
and \g446742/U$2 ( \21236 , \19467 , RIe1e2220_3950);
and \g446742/U$3 ( \21237 , RIe1e4f20_3982, \19469 );
nor \g446742/U$1 ( \21238 , \21236 , \21237 );
nand \g444589/U$1 ( \21239 , \21229 , \21232 , \21235 , \21238 );
and \g445950/U$2 ( \21240 , RIe186060_2902, \16427 );
and \g445950/U$3 ( \21241 , RIe183360_2870, \16368 );
and \g448815/U$2 ( \21242 , RIe194160_3062, \16485 );
and \g448815/U$3 ( \21243 , \16356 , RIf144140_5234);
and \g448815/U$4 ( \21244 , RIe180660_2838, \16398 );
nor \g448815/U$1 ( \21245 , \21242 , \21243 , \21244 );
and \g454571/U$2 ( \21246 , \16317 , RIe199b60_3126);
and \g454571/U$3 ( \21247 , RIe19c860_3158, \16325 );
nor \g454571/U$1 ( \21248 , \21246 , \21247 );
not \g449841/U$3 ( \21249 , \21248 );
not \g449841/U$4 ( \21250 , \16311 );
and \g449841/U$2 ( \21251 , \21249 , \21250 );
and \g449841/U$5 ( \21252 , \16341 , RIf142ac0_5218);
nor \g449841/U$1 ( \21253 , \21251 , \21252 );
and \g451665/U$2 ( \21254 , \16377 , RIe196e60_3094);
and \g451665/U$3 ( \21255 , RIf145220_5246, \16313 );
nor \g451665/U$1 ( \21256 , \21254 , \21255 );
and \g451666/U$2 ( \21257 , \16334 , RIe18e760_2998);
and \g451666/U$3 ( \21258 , RIe191460_3030, \16380 );
nor \g451666/U$1 ( \21259 , \21257 , \21258 );
nand \g447295/U$1 ( \21260 , \21245 , \21253 , \21256 , \21259 );
nor \g445950/U$1 ( \21261 , \21240 , \21241 , \21260 );
and \g451664/U$2 ( \21262 , \16361 , RIe17ac60_2774);
and \g451664/U$3 ( \21263 , RIe188d60_2934, \16432 );
nor \g451664/U$1 ( \21264 , \21262 , \21263 );
and \g451662/U$2 ( \21265 , \16364 , RIe17d960_2806);
and \g451662/U$3 ( \21266 , RIf1431c8_5223, \16371 );
nor \g451662/U$1 ( \21267 , \21265 , \21266 );
and \g445113/U$2 ( \21268 , \21261 , \21264 , \21267 );
nor \g445113/U$1 ( \21269 , \21268 , \16618 );
and \g445954/U$2 ( \21270 , RIf15d910_5524, \16427 );
and \g445954/U$3 ( \21271 , RIfe8c868_7943, \16368 );
and \g448816/U$2 ( \21272 , RIf163ce8_5595, \16344 );
and \g448816/U$3 ( \21273 , \16356 , RIfc9c578_6801);
and \g448816/U$4 ( \21274 , RIf15aee0_5494, \16398 );
nor \g448816/U$1 ( \21275 , \21272 , \21273 , \21274 );
and \g454630/U$2 ( \21276 , \16317 , RIf165908_5615);
and \g454630/U$3 ( \21277 , RIf1669e8_5627, \16325 );
nor \g454630/U$1 ( \21278 , \21276 , \21277 );
not \g449842/U$3 ( \21279 , \21278 );
not \g449842/U$4 ( \21280 , \16311 );
and \g449842/U$2 ( \21281 , \21279 , \21280 );
and \g449842/U$5 ( \21282 , \16341 , RIf15c3f8_5509);
nor \g449842/U$1 ( \21283 , \21281 , \21282 );
and \g451760/U$2 ( \21284 , \16377 , RIfe8c700_7942);
and \g451760/U$3 ( \21285 , RIfe8c9d0_7944, \16313 );
nor \g451760/U$1 ( \21286 , \21284 , \21285 );
and \g451675/U$2 ( \21287 , \16334 , RIf161588_5567);
and \g451675/U$3 ( \21288 , RIf162d70_5584, \16380 );
nor \g451675/U$1 ( \21289 , \21287 , \21288 );
nand \g447296/U$1 ( \21290 , \21275 , \21283 , \21286 , \21289 );
nor \g445954/U$1 ( \21291 , \21270 , \21271 , \21290 );
and \g451672/U$2 ( \21292 , \16361 , RIf1596f8_5477);
and \g451672/U$3 ( \21293 , RIf15f698_5545, \16448 );
nor \g451672/U$1 ( \21294 , \21292 , \21293 );
and \g451671/U$2 ( \21295 , \16364 , RIf15a0d0_5484);
and \g451671/U$3 ( \21296 , RIfe8c598_7941, \16371 );
nor \g451671/U$1 ( \21297 , \21295 , \21296 );
and \g445114/U$2 ( \21298 , \21291 , \21294 , \21297 );
nor \g445114/U$1 ( \21299 , \21298 , \16393 );
or \g444389/U$1 ( \21300 , \21179 , \21239 , \21269 , \21299 );
and \g445948/U$2 ( \21301 , RIf16c820_5694, \16328 );
and \g445948/U$3 ( \21302 , RIe214ab8_4525, \16334 );
and \g448811/U$2 ( \21303 , RIe211db8_4493, \16427 );
and \g448811/U$3 ( \21304 , \16448 , RIfe8c430_7940);
and \g448811/U$4 ( \21305 , RIe21d1b8_4621, \16485 );
nor \g448811/U$1 ( \21306 , \21303 , \21304 , \21305 );
and \g454357/U$2 ( \21307 , \16317 , RIe20c3b8_4429);
and \g454357/U$3 ( \21308 , RIf167960_5638, \16325 );
nor \g454357/U$1 ( \21309 , \21307 , \21308 );
not \g454356/U$1 ( \21310 , \21309 );
and \g450024/U$2 ( \21311 , \21310 , \16336 );
and \g450024/U$3 ( \21312 , RIf16a7c8_5671, \16356 );
nor \g450024/U$1 ( \21313 , \21311 , \21312 );
and \g451655/U$2 ( \21314 , \16361 , RIe2069b8_4365);
and \g451655/U$3 ( \21315 , RIe2096b8_4397, \16364 );
nor \g451655/U$1 ( \21316 , \21314 , \21315 );
and \g451654/U$2 ( \21317 , \16368 , RIe20f0b8_4461);
and \g451654/U$3 ( \21318 , RIf1688d8_5649, \16371 );
nor \g451654/U$1 ( \21319 , \21317 , \21318 );
nand \g448048/U$1 ( \21320 , \21306 , \21313 , \21316 , \21319 );
nor \g445948/U$1 ( \21321 , \21301 , \21302 , \21320 );
and \g451652/U$2 ( \21322 , \16377 , RIe21feb8_4653);
and \g451652/U$3 ( \21323 , RIe2177b8_4557, \16380 );
nor \g451652/U$1 ( \21324 , \21322 , \21323 );
and \g451651/U$2 ( \21325 , \16313 , RIf16b740_5682);
and \g451651/U$3 ( \21326 , RIe222bb8_4685, \16319 );
nor \g451651/U$1 ( \21327 , \21325 , \21326 );
and \g445111/U$2 ( \21328 , \21321 , \21324 , \21327 );
nor \g445111/U$1 ( \21329 , \21328 , \16389 );
and \g445949/U$2 ( \21330 , RIee3bb78_5138, \16448 );
and \g445949/U$3 ( \21331 , RIfcc4af0_7260, \16361 );
and \g448812/U$2 ( \21332 , RIf140798_5193, \16321 );
and \g448812/U$3 ( \21333 , \16328 , RIf141cb0_5208);
and \g448812/U$4 ( \21334 , RIf16ef80_5722, \16398 );
nor \g448812/U$1 ( \21335 , \21332 , \21333 , \21334 );
and \g454480/U$2 ( \21336 , \16317 , RIf13eb78_5173);
and \g454480/U$3 ( \21337 , RIfceb880_7702, \16325 );
nor \g454480/U$1 ( \21338 , \21336 , \21337 );
not \g449838/U$3 ( \21339 , \21338 );
not \g449838/U$4 ( \21340 , \16330 );
and \g449838/U$2 ( \21341 , \21339 , \21340 );
and \g449838/U$5 ( \21342 , \16341 , RIf16fac0_5730);
nor \g449838/U$1 ( \21343 , \21341 , \21342 );
and \g452131/U$2 ( \21344 , \16377 , RIfe8be90_7936);
and \g452131/U$3 ( \21345 , RIf13ff28_5187, \16313 );
nor \g452131/U$1 ( \21346 , \21344 , \21345 );
and \g451660/U$2 ( \21347 , \16334 , RIee3cdc0_5151);
and \g451660/U$3 ( \21348 , RIee3e008_5164, \16380 );
nor \g451660/U$1 ( \21349 , \21347 , \21348 );
nand \g447294/U$1 ( \21350 , \21335 , \21343 , \21346 , \21349 );
nor \g445949/U$1 ( \21351 , \21330 , \21331 , \21350 );
and \g452183/U$2 ( \21352 , \16364 , RIf16dbd0_5708);
and \g452183/U$3 ( \21353 , RIe172c68_2683, \16368 );
nor \g452183/U$1 ( \21354 , \21352 , \21353 );
and \g452153/U$2 ( \21355 , \16371 , RIee396e8_5112);
and \g452153/U$3 ( \21356 , RIee3aa98_5126, \16427 );
nor \g452153/U$1 ( \21357 , \21355 , \21356 );
and \g445112/U$2 ( \21358 , \21351 , \21354 , \21357 );
nor \g445112/U$1 ( \21359 , \21358 , \16649 );
or \g444209/U$1 ( \21360 , \21300 , \21329 , \21359 );
_DC \g3d41/U$1 ( \21361 , \21360 , \16652 );
and \g446598/U$2 ( \21362 , \19208 , RIe1bd7b8_3533);
and \g446598/U$3 ( \21363 , RIe1c04b8_3565, \19213 );
nor \g446598/U$1 ( \21364 , \21362 , \21363 );
and \g445803/U$2 ( \21365 , RIe1c5eb8_3629, \16341 );
and \g445803/U$3 ( \21366 , RIe1c31b8_3597, \16337 );
and \g448623/U$2 ( \21367 , RIe1e7ab8_4013, \16321 );
and \g448623/U$3 ( \21368 , \16485 , RIe1dc6b8_3885);
and \g448623/U$4 ( \21369 , RIe1df3b8_3917, \16356 );
nor \g448623/U$1 ( \21370 , \21367 , \21368 , \21369 );
and \g451028/U$2 ( \21371 , \16368 , RIe1c8bb8_3661);
and \g451028/U$3 ( \21372 , RIe1cb8b8_3693, \16371 );
nor \g451028/U$1 ( \21373 , \21371 , \21372 );
and \g455382/U$2 ( \21374 , \16317 , RIe1ce5b8_3725);
and \g455382/U$3 ( \21375 , RIe1d12b8_3757, \16325 );
nor \g455382/U$1 ( \21376 , \21374 , \21375 );
not \g449651/U$3 ( \21377 , \21376 );
not \g449651/U$4 ( \21378 , \16351 );
and \g449651/U$2 ( \21379 , \21377 , \21378 );
and \g449651/U$5 ( \21380 , \16328 , RIe1ea7b8_4045);
nor \g449651/U$1 ( \21381 , \21379 , \21380 );
and \g451027/U$2 ( \21382 , \16334 , RIe1d6cb8_3821);
and \g451027/U$3 ( \21383 , RIe1d99b8_3853, \16380 );
nor \g451027/U$1 ( \21384 , \21382 , \21383 );
nand \g447526/U$1 ( \21385 , \21370 , \21373 , \21381 , \21384 );
nor \g445803/U$1 ( \21386 , \21365 , \21366 , \21385 );
not \g444838/U$3 ( \21387 , \21386 );
not \g444838/U$4 ( \21388 , \16555 );
and \g444838/U$2 ( \21389 , \21387 , \21388 );
and \g445805/U$2 ( \21390 , RIf1569f8_5445, \16313 );
and \g445805/U$3 ( \21391 , RIe1ed350_4076, \16361 );
and \g448626/U$2 ( \21392 , RIf151430_5384, \16427 );
and \g448626/U$3 ( \21393 , \16448 , RIf1527e0_5398);
and \g448626/U$4 ( \21394 , RIf157268_5451, \16321 );
nor \g448626/U$1 ( \21395 , \21392 , \21393 , \21394 );
and \g451035/U$2 ( \21396 , \16368 , RIe1f2648_4135);
and \g451035/U$3 ( \21397 , RIfcd2650_7416, \16371 );
nor \g451035/U$1 ( \21398 , \21396 , \21397 );
and \g454342/U$2 ( \21399 , \16317 , RIf155210_5428);
and \g454342/U$3 ( \21400 , RIf155d50_5436, \16325 );
nor \g454342/U$1 ( \21401 , \21399 , \21400 );
not \g449654/U$3 ( \21402 , \21401 );
not \g449654/U$4 ( \21403 , \16330 );
and \g449654/U$2 ( \21404 , \21402 , \21403 );
and \g449654/U$5 ( \21405 , \16328 , RIf1584b0_5464);
nor \g449654/U$1 ( \21406 , \21404 , \21405 );
and \g451033/U$2 ( \21407 , \16334 , RIfe96750_8056);
and \g451033/U$3 ( \21408 , RIf153e60_5414, \16380 );
nor \g451033/U$1 ( \21409 , \21407 , \21408 );
nand \g447528/U$1 ( \21410 , \21395 , \21398 , \21406 , \21409 );
nor \g445805/U$1 ( \21411 , \21390 , \21391 , \21410 );
and \g451032/U$2 ( \21412 , \16364 , RIf14d4e8_5339);
and \g451032/U$3 ( \21413 , RIf14f108_5359, \16341 );
nor \g451032/U$1 ( \21414 , \21412 , \21413 );
and \g451031/U$2 ( \21415 , \16398 , RIfc7f298_6469);
and \g451031/U$3 ( \21416 , RIfe965e8_8055, \16377 );
nor \g451031/U$1 ( \21417 , \21415 , \21416 );
and \g445005/U$2 ( \21418 , \21411 , \21414 , \21417 );
nor \g445005/U$1 ( \21419 , \21418 , \16480 );
nor \g444838/U$1 ( \21420 , \21389 , \21419 );
and \g446599/U$2 ( \21421 , \19467 , RIe1e20b8_3949);
and \g446599/U$3 ( \21422 , RIe1e4db8_3981, \19469 );
nor \g446599/U$1 ( \21423 , \21421 , \21422 );
nand \g444418/U$1 ( \21424 , \21364 , \21420 , \21423 );
and \g451047/U$2 ( \21425 , \16334 , RIe214950_4524);
and \g451047/U$3 ( \21426 , RIf168770_5648, \16371 );
nor \g451047/U$1 ( \21427 , \21425 , \21426 );
and \g445808/U$2 ( \21428 , RIe21d050_4620, \16485 );
and \g445808/U$3 ( \21429 , RIe217650_4556, \16380 );
and \g448630/U$2 ( \21430 , RIe222a50_4684, \16319 );
and \g448630/U$3 ( \21431 , \16326 , RIfe96e58_8061);
and \g448630/U$4 ( \21432 , RIe211c50_4492, \16427 );
nor \g448630/U$1 ( \21433 , \21430 , \21431 , \21432 );
and \g451052/U$2 ( \21434 , \16361 , RIe206850_4364);
and \g451052/U$3 ( \21435 , RIe209550_4396, \16364 );
nor \g451052/U$1 ( \21436 , \21434 , \21435 );
and \g451050/U$2 ( \21437 , \16377 , RIe21fd50_4652);
and \g451050/U$3 ( \21438 , RIfe96cf0_8060, \16313 );
nor \g451050/U$1 ( \21439 , \21437 , \21438 );
and \g454420/U$2 ( \21440 , \16317 , RIe20c250_4428);
and \g454420/U$3 ( \21441 , RIf1677f8_5637, \16325 );
nor \g454420/U$1 ( \21442 , \21440 , \21441 );
not \g454419/U$1 ( \21443 , \21442 );
and \g449657/U$2 ( \21444 , \21443 , \16336 );
and \g449657/U$3 ( \21445 , RIf169f58_5665, \16448 );
nor \g449657/U$1 ( \21446 , \21444 , \21445 );
nand \g448020/U$1 ( \21447 , \21433 , \21436 , \21439 , \21446 );
nor \g445808/U$1 ( \21448 , \21428 , \21429 , \21447 );
and \g451046/U$2 ( \21449 , \16368 , RIe20ef50_4460);
and \g451046/U$3 ( \21450 , RIf16a660_5670, \16354 );
nor \g451046/U$1 ( \21451 , \21449 , \21450 );
nand \g445532/U$1 ( \21452 , \21427 , \21448 , \21451 );
and \g444737/U$2 ( \21453 , \21452 , \16390 );
and \g448628/U$2 ( \21454 , RIee3a930_5125, \16427 );
and \g448628/U$3 ( \21455 , \16448 , RIee3ba10_5137);
and \g448628/U$4 ( \21456 , RIfc542f0_5980, \16321 );
nor \g448628/U$1 ( \21457 , \21454 , \21455 , \21456 );
and \g451041/U$2 ( \21458 , \16368 , RIe172b00_2682);
and \g451041/U$3 ( \21459 , RIfe97290_8064, \16371 );
nor \g451041/U$1 ( \21460 , \21458 , \21459 );
and \g454345/U$2 ( \21461 , \16317 , RIfc48680_5846);
and \g454345/U$3 ( \21462 , RIfca0bc8_6851, \16325 );
nor \g454345/U$1 ( \21463 , \21461 , \21462 );
not \g449656/U$3 ( \21464 , \21463 );
not \g449656/U$4 ( \21465 , \16330 );
and \g449656/U$2 ( \21466 , \21464 , \21465 );
and \g449656/U$5 ( \21467 , \16326 , RIf141b48_5207);
nor \g449656/U$1 ( \21468 , \21466 , \21467 );
and \g451040/U$2 ( \21469 , \16334 , RIfcc6878_7281);
and \g451040/U$3 ( \21470 , RIee3dea0_5163, \16380 );
nor \g451040/U$1 ( \21471 , \21469 , \21470 );
nand \g447529/U$1 ( \21472 , \21457 , \21460 , \21468 , \21471 );
and \g444737/U$3 ( \21473 , \17998 , \21472 );
nor \g444737/U$1 ( \21474 , \21453 , \21473 );
and \g446600/U$2 ( \21475 , \18711 , RIe175260_2710);
and \g446600/U$3 ( \21476 , RIfc800a8_6479, \18713 );
nor \g446600/U$1 ( \21477 , \21475 , \21476 );
and \g446601/U$2 ( \21478 , \18716 , RIf16ee18_5721);
and \g446601/U$3 ( \21479 , RIf16f958_5729, \18718 );
nor \g446601/U$1 ( \21480 , \21478 , \21479 );
and \g446602/U$2 ( \21481 , \18533 , RIf16d360_5702);
and \g446602/U$3 ( \21482 , RIf16da68_5707, \18535 );
nor \g446602/U$1 ( \21483 , \21481 , \21482 );
nand \g444564/U$1 ( \21484 , \21474 , \21477 , \21480 , \21483 );
and \g445799/U$2 ( \21485 , RIe18b8f8_2965, \16356 );
and \g445799/U$3 ( \21486 , RIe21a350_4588, \16334 );
and \g448620/U$2 ( \21487 , RIe1a4df8_3253, \16321 );
and \g448620/U$3 ( \21488 , \16328 , RIe1a7af8_3285);
and \g448620/U$4 ( \21489 , RIe1fdbb0_4264, \16427 );
nor \g448620/U$1 ( \21490 , \21487 , \21488 , \21489 );
and \g451011/U$2 ( \21491 , \16361 , RIe16ff68_2651);
and \g451011/U$3 ( \21492 , RIe1ad930_3352, \16364 );
nor \g451011/U$1 ( \21493 , \21491 , \21492 );
and \g451010/U$2 ( \21494 , \16377 , RIe19f3f8_3189);
and \g451010/U$3 ( \21495 , RIe1a20f8_3221, \16313 );
nor \g451010/U$1 ( \21496 , \21494 , \21495 );
and \g454335/U$2 ( \21497 , \16317 , RIe1baab8_3501);
and \g454335/U$3 ( \21498 , RIe1d3fb8_3789, \16325 );
nor \g454335/U$1 ( \21499 , \21497 , \21498 );
not \g454334/U$1 ( \21500 , \21499 );
and \g449647/U$2 ( \21501 , \21500 , \16336 );
and \g449647/U$3 ( \21502 , RIe203b50_4332, \16448 );
nor \g449647/U$1 ( \21503 , \21501 , \21502 );
nand \g448018/U$1 ( \21504 , \21490 , \21493 , \21496 , \21503 );
nor \g445799/U$1 ( \21505 , \21485 , \21486 , \21504 );
and \g451008/U$2 ( \21506 , \16371 , RIe1f6f68_4187);
and \g451008/U$3 ( \21507 , RIe225750_4716, \16380 );
nor \g451008/U$1 ( \21508 , \21506 , \21507 );
and \g451009/U$2 ( \21509 , \16368 , RIe1efab0_4104);
and \g451009/U$3 ( \21510 , RIe177df8_2741, \16485 );
nor \g451009/U$1 ( \21511 , \21509 , \21510 );
and \g445000/U$2 ( \21512 , \21505 , \21508 , \21511 );
nor \g445000/U$1 ( \21513 , \21512 , \16586 );
and \g445802/U$2 ( \21514 , RIe1b8790_3476, \16313 );
and \g445802/U$3 ( \21515 , RIfe961b0_8052, \16364 );
and \g448621/U$2 ( \21516 , RIfc58d78_6033, \16427 );
and \g448621/U$3 ( \21517 , \16448 , RIf148628_5283);
and \g448621/U$4 ( \21518 , RIf14ad88_5311, \16321 );
nor \g448621/U$1 ( \21519 , \21516 , \21517 , \21518 );
and \g451023/U$2 ( \21520 , \16368 , RIe1b04c8_3383);
and \g451023/U$3 ( \21521 , RIe1b20e8_3403, \16371 );
nor \g451023/U$1 ( \21522 , \21520 , \21521 );
and \g454248/U$2 ( \21523 , \16317 , RIf149870_5296);
and \g454248/U$3 ( \21524 , RIf14a0e0_5302, \16325 );
nor \g454248/U$1 ( \21525 , \21523 , \21524 );
not \g449648/U$3 ( \21526 , \21525 );
not \g449648/U$4 ( \21527 , \16330 );
and \g449648/U$2 ( \21528 , \21526 , \21527 );
and \g449648/U$5 ( \21529 , \16328 , RIf14c138_5325);
nor \g449648/U$1 ( \21530 , \21528 , \21529 );
and \g451020/U$2 ( \21531 , \16334 , RIfe96318_8053);
and \g451020/U$3 ( \21532 , RIfe97128_8063, \16380 );
nor \g451020/U$1 ( \21533 , \21531 , \21532 );
nand \g447525/U$1 ( \21534 , \21519 , \21522 , \21530 , \21533 );
nor \g445802/U$1 ( \21535 , \21514 , \21515 , \21534 );
and \g451017/U$2 ( \21536 , \16339 , RIf146cd8_5265);
and \g451017/U$3 ( \21537 , RIfe96480_8054, \16377 );
nor \g451017/U$1 ( \21538 , \21536 , \21537 );
and \g451019/U$2 ( \21539 , \16361 , RIfe96fc0_8062);
and \g451019/U$3 ( \21540 , RIfc591b0_6036, \16398 );
nor \g451019/U$1 ( \21541 , \21539 , \21540 );
and \g445002/U$2 ( \21542 , \21535 , \21538 , \21541 );
nor \g445002/U$1 ( \21543 , \21542 , \16909 );
or \g444288/U$1 ( \21544 , \21424 , \21484 , \21513 , \21543 );
and \g445794/U$2 ( \21545 , RIf142958_5217, \16341 );
and \g445794/U$3 ( \21546 , RIe196cf8_3093, \16377 );
and \g448617/U$2 ( \21547 , RIe185ef8_2901, \16427 );
and \g448617/U$3 ( \21548 , \16448 , RIe188bf8_2933);
and \g448617/U$4 ( \21549 , RIe1999f8_3125, \16321 );
nor \g448617/U$1 ( \21550 , \21547 , \21548 , \21549 );
and \g450995/U$2 ( \21551 , \16368 , RIe1831f8_2869);
and \g450995/U$3 ( \21552 , RIfe973f8_8065, \16371 );
nor \g450995/U$1 ( \21553 , \21551 , \21552 );
and \g454631/U$2 ( \21554 , \16317 , RIe193ff8_3061);
and \g454631/U$3 ( \21555 , RIf143fd8_5233, \16325 );
nor \g454631/U$1 ( \21556 , \21554 , \21555 );
not \g449644/U$3 ( \21557 , \21556 );
not \g449644/U$4 ( \21558 , \16330 );
and \g449644/U$2 ( \21559 , \21557 , \21558 );
and \g449644/U$5 ( \21560 , \16328 , RIe19c6f8_3157);
nor \g449644/U$1 ( \21561 , \21559 , \21560 );
and \g450994/U$2 ( \21562 , \16334 , RIe18e5f8_2997);
and \g450994/U$3 ( \21563 , RIe1912f8_3029, \16380 );
nor \g450994/U$1 ( \21564 , \21562 , \21563 );
nand \g447520/U$1 ( \21565 , \21550 , \21553 , \21561 , \21564 );
nor \g445794/U$1 ( \21566 , \21545 , \21546 , \21565 );
and \g450991/U$2 ( \21567 , \16361 , RIe17aaf8_2773);
and \g450991/U$3 ( \21568 , RIf1450b8_5245, \16313 );
nor \g450991/U$1 ( \21569 , \21567 , \21568 );
and \g450992/U$2 ( \21570 , \16364 , RIe17d7f8_2805);
and \g450992/U$3 ( \21571 , RIe1804f8_2837, \16337 );
nor \g450992/U$1 ( \21572 , \21570 , \21571 );
and \g444997/U$2 ( \21573 , \21566 , \21569 , \21572 );
nor \g444997/U$1 ( \21574 , \21573 , \16618 );
and \g445797/U$2 ( \21575 , RIf163b80_5594, \16344 );
and \g445797/U$3 ( \21576 , RIf162c08_5583, \16380 );
and \g448618/U$2 ( \21577 , RIf1657a0_5614, \16321 );
and \g448618/U$3 ( \21578 , \16328 , RIf166880_5626);
and \g448618/U$4 ( \21579 , RIf15d7a8_5523, \16427 );
nor \g448618/U$1 ( \21580 , \21577 , \21578 , \21579 );
and \g451003/U$2 ( \21581 , \16361 , RIf159590_5476);
and \g451003/U$3 ( \21582 , RIfc579c8_6019, \16364 );
nor \g451003/U$1 ( \21583 , \21581 , \21582 );
and \g451001/U$2 ( \21584 , \16377 , RIe2005e0_4294);
and \g451001/U$3 ( \21585 , RIe201dc8_4311, \16313 );
nor \g451001/U$1 ( \21586 , \21584 , \21585 );
and \g454332/U$2 ( \21587 , \16317 , RIfc7cf70_6444);
and \g454332/U$3 ( \21588 , RIfcb3fc0_7070, \16325 );
nor \g454332/U$1 ( \21589 , \21587 , \21588 );
not \g454331/U$1 ( \21590 , \21589 );
and \g449645/U$2 ( \21591 , \21590 , \16336 );
and \g449645/U$3 ( \21592 , RIf15f530_5544, \16448 );
nor \g449645/U$1 ( \21593 , \21591 , \21592 );
nand \g448017/U$1 ( \21594 , \21580 , \21583 , \21586 , \21593 );
nor \g445797/U$1 ( \21595 , \21575 , \21576 , \21594 );
and \g450999/U$2 ( \21596 , \16368 , RIfe96a20_8058);
and \g450999/U$3 ( \21597 , RIfe96b88_8059, \16356 );
nor \g450999/U$1 ( \21598 , \21596 , \21597 );
and \g451000/U$2 ( \21599 , \16334 , RIf161420_5566);
and \g451000/U$3 ( \21600 , RIfe968b8_8057, \16371 );
nor \g451000/U$1 ( \21601 , \21599 , \21600 );
and \g444998/U$2 ( \21602 , \21595 , \21598 , \21601 );
nor \g444998/U$1 ( \21603 , \21602 , \16393 );
or \g444197/U$1 ( \21604 , \21544 , \21574 , \21603 );
_DC \g3dc6/U$1 ( \21605 , \21604 , \16652 );
and \g451202/U$2 ( \21606 , \16313 , RIe176bb0_2728);
and \g451202/U$3 ( \21607 , RIf140630_5192, \16321 );
nor \g451202/U$1 ( \21608 , \21606 , \21607 );
and \g445843/U$2 ( \21609 , RIf1419e0_5206, \16328 );
and \g445843/U$3 ( \21610 , RIee3cc58_5150, \16334 );
and \g448674/U$2 ( \21611 , RIf16ecb0_5720, \16398 );
and \g448674/U$3 ( \21612 , \16341 , RIf16f7f0_5728);
and \g448674/U$4 ( \21613 , RIfc5f6f0_6108, \16485 );
nor \g448674/U$1 ( \21614 , \21611 , \21612 , \21613 );
and \g454604/U$2 ( \21615 , \16317 , RIee3a7c8_5124);
and \g454604/U$3 ( \21616 , RIee3b8a8_5136, \16325 );
nor \g454604/U$1 ( \21617 , \21615 , \21616 );
not \g449702/U$3 ( \21618 , \21617 );
not \g449702/U$4 ( \21619 , \16351 );
and \g449702/U$2 ( \21620 , \21618 , \21619 );
and \g449702/U$5 ( \21621 , \16356 , RIfcd1840_7406);
nor \g449702/U$1 ( \21622 , \21620 , \21621 );
and \g451207/U$2 ( \21623 , \16361 , RIfc78ec0_6398);
and \g451207/U$3 ( \21624 , RIf16d900_5706, \16364 );
nor \g451207/U$1 ( \21625 , \21623 , \21624 );
and \g451205/U$2 ( \21626 , \16368 , RIfea9008_8239);
and \g451205/U$3 ( \21627 , RIee39580_5111, \16371 );
nor \g451205/U$1 ( \21628 , \21626 , \21627 );
nand \g447559/U$1 ( \21629 , \21614 , \21622 , \21625 , \21628 );
nor \g445843/U$1 ( \21630 , \21609 , \21610 , \21629 );
and \g451203/U$2 ( \21631 , \16377 , RIe1750f8_2709);
and \g451203/U$3 ( \21632 , RIee3dd38_5162, \16380 );
nor \g451203/U$1 ( \21633 , \21631 , \21632 );
nand \g445537/U$1 ( \21634 , \21608 , \21630 , \21633 );
and \g444750/U$2 ( \21635 , \21634 , \17998 );
and \g448672/U$2 ( \21636 , RIe185d90_2900, \16427 );
and \g448672/U$3 ( \21637 , \16432 , RIe188a90_2932);
and \g448672/U$4 ( \21638 , RIe193e90_3060, \16485 );
nor \g448672/U$1 ( \21639 , \21636 , \21637 , \21638 );
and \g454556/U$2 ( \21640 , \16317 , RIe180390_2836);
and \g454556/U$3 ( \21641 , RIfc76e68_6375, \16325 );
nor \g454556/U$1 ( \21642 , \21640 , \21641 );
not \g454555/U$1 ( \21643 , \21642 );
and \g449700/U$2 ( \21644 , \21643 , \16336 );
and \g449700/U$3 ( \21645 , RIfc76058_6365, \16354 );
nor \g449700/U$1 ( \21646 , \21644 , \21645 );
and \g451197/U$2 ( \21647 , \16361 , RIe17a990_2772);
and \g451197/U$3 ( \21648 , RIe17d690_2804, \16364 );
nor \g451197/U$1 ( \21649 , \21647 , \21648 );
and \g451196/U$2 ( \21650 , \16368 , RIe183090_2868);
and \g451196/U$3 ( \21651 , RIfccd8f8_7361, \16371 );
nor \g451196/U$1 ( \21652 , \21650 , \21651 );
nand \g448024/U$1 ( \21653 , \21639 , \21646 , \21649 , \21652 );
and \g444750/U$3 ( \21654 , \17938 , \21653 );
nor \g444750/U$1 ( \21655 , \21635 , \21654 );
and \g446632/U$2 ( \21656 , \18960 , RIe18e490_2996);
and \g446632/U$3 ( \21657 , RIe191190_3028, \18962 );
nor \g446632/U$1 ( \21658 , \21656 , \21657 );
and \g446631/U$2 ( \21659 , \18965 , RIe199890_3124);
and \g446631/U$3 ( \21660 , RIe19c590_3156, \18967 );
nor \g446631/U$1 ( \21661 , \21659 , \21660 );
and \g446633/U$2 ( \21662 , \18776 , RIe196b90_3092);
and \g446633/U$3 ( \21663 , RIf144f50_5244, \18778 );
nor \g446633/U$1 ( \21664 , \21662 , \21663 );
nand \g444463/U$1 ( \21665 , \21655 , \21658 , \21661 , \21664 );
and \g451221/U$2 ( \21666 , \16364 , RIfe92538_8009);
and \g451221/U$3 ( \21667 , RIfe92808_8011, \16371 );
nor \g451221/U$1 ( \21668 , \21666 , \21667 );
and \g445845/U$2 ( \21669 , RIf15d640_5522, \16427 );
and \g445845/U$3 ( \21670 , RIfe92c40_8014, \16368 );
and \g448678/U$2 ( \21671 , RIfcc6f80_7286, \16319 );
and \g448678/U$3 ( \21672 , \16328 , RIfc45110_5808);
and \g448678/U$4 ( \21673 , RIfe92da8_8015, \16398 );
nor \g448678/U$1 ( \21674 , \21671 , \21672 , \21673 );
and \g454597/U$2 ( \21675 , \16317 , RIf163a18_5593);
and \g454597/U$3 ( \21676 , RIf164af8_5605, \16325 );
nor \g454597/U$1 ( \21677 , \21675 , \21676 );
not \g449829/U$3 ( \21678 , \21677 );
not \g449829/U$4 ( \21679 , \16330 );
and \g449829/U$2 ( \21680 , \21678 , \21679 );
and \g449829/U$5 ( \21681 , \16341 , RIfe926a0_8010);
nor \g449829/U$1 ( \21682 , \21680 , \21681 );
and \g451647/U$2 ( \21683 , \16377 , RIfe92970_8012);
and \g451647/U$3 ( \21684 , RIfe92f10_8016, \16313 );
nor \g451647/U$1 ( \21685 , \21683 , \21684 );
and \g451225/U$2 ( \21686 , \16334 , RIfe92ad8_8013);
and \g451225/U$3 ( \21687 , RIf162aa0_5582, \16380 );
nor \g451225/U$1 ( \21688 , \21686 , \21687 );
nand \g447269/U$1 ( \21689 , \21674 , \21682 , \21685 , \21688 );
nor \g445845/U$1 ( \21690 , \21669 , \21670 , \21689 );
and \g451222/U$2 ( \21691 , \16361 , RIfcb5a78_7089);
and \g451222/U$3 ( \21692 , RIf15f3c8_5543, \16448 );
nor \g451222/U$1 ( \21693 , \21691 , \21692 );
nand \g445539/U$1 ( \21694 , \21668 , \21690 , \21693 );
and \g444761/U$2 ( \21695 , \21694 , \16394 );
and \g448677/U$2 ( \21696 , RIe211ae8_4491, \16427 );
and \g448677/U$3 ( \21697 , \16448 , RIfca2c20_6874);
and \g448677/U$4 ( \21698 , RIe21cee8_4619, \16485 );
nor \g448677/U$1 ( \21699 , \21696 , \21697 , \21698 );
and \g454640/U$2 ( \21700 , \16317 , RIe20c0e8_4427);
and \g454640/U$3 ( \21701 , RIfcc24f8_7233, \16325 );
nor \g454640/U$1 ( \21702 , \21700 , \21701 );
not \g454639/U$1 ( \21703 , \21702 );
and \g449705/U$2 ( \21704 , \21703 , \16336 );
and \g449705/U$3 ( \21705 , RIfc74000_6342, \16356 );
nor \g449705/U$1 ( \21706 , \21704 , \21705 );
and \g451215/U$2 ( \21707 , \16361 , RIe2066e8_4363);
and \g451215/U$3 ( \21708 , RIe2093e8_4395, \16364 );
nor \g451215/U$1 ( \21709 , \21707 , \21708 );
and \g451214/U$2 ( \21710 , \16368 , RIe20ede8_4459);
and \g451214/U$3 ( \21711 , RIfca2950_6872, \16371 );
nor \g451214/U$1 ( \21712 , \21710 , \21711 );
nand \g448025/U$1 ( \21713 , \21699 , \21706 , \21709 , \21712 );
and \g444761/U$3 ( \21714 , \16390 , \21713 );
nor \g444761/U$1 ( \21715 , \21695 , \21714 );
and \g446637/U$2 ( \21716 , \18020 , RIe2228e8_4683);
and \g446637/U$3 ( \21717 , RIfcc8060_7298, \18022 );
nor \g446637/U$1 ( \21718 , \21716 , \21717 );
and \g446638/U$2 ( \21719 , \18025 , RIe21fbe8_4651);
and \g446638/U$3 ( \21720 , RIfc5a3f8_6049, \18027 );
nor \g446638/U$1 ( \21721 , \21719 , \21720 );
and \g446639/U$2 ( \21722 , \18030 , RIe2147e8_4523);
and \g446639/U$3 ( \21723 , RIe2174e8_4555, \18032 );
nor \g446639/U$1 ( \21724 , \21722 , \21723 );
nand \g444464/U$1 ( \21725 , \21715 , \21718 , \21721 , \21724 );
and \g445838/U$2 ( \21726 , RIf158348_5463, \16326 );
and \g445838/U$3 ( \21727 , RIfec3a20_8346, \16334 );
and \g448667/U$2 ( \21728 , RIfec3750_8344, \16427 );
and \g448667/U$3 ( \21729 , \16432 , RIf152678_5397);
and \g448667/U$4 ( \21730 , RIf1550a8_5427, \16485 );
nor \g448667/U$1 ( \21731 , \21728 , \21729 , \21730 );
and \g454741/U$2 ( \21732 , \16317 , RIf14e898_5353);
and \g454741/U$3 ( \21733 , RIf14efa0_5358, \16325 );
nor \g454741/U$1 ( \21734 , \21732 , \21733 );
not \g454740/U$1 ( \21735 , \21734 );
and \g449695/U$2 ( \21736 , \21735 , \16336 );
and \g449695/U$3 ( \21737 , RIfcc5ea0_7274, \16356 );
nor \g449695/U$1 ( \21738 , \21736 , \21737 );
and \g451183/U$2 ( \21739 , \16361 , RIfe92268_8007);
and \g451183/U$3 ( \21740 , RIf14d380_5338, \16364 );
nor \g451183/U$1 ( \21741 , \21739 , \21740 );
and \g451181/U$2 ( \21742 , \16368 , RIfe923d0_8008);
and \g451181/U$3 ( \21743 , RIf14ff18_5369, \16371 );
nor \g451181/U$1 ( \21744 , \21742 , \21743 );
nand \g448023/U$1 ( \21745 , \21731 , \21738 , \21741 , \21744 );
nor \g445838/U$1 ( \21746 , \21726 , \21727 , \21745 );
and \g451180/U$2 ( \21747 , \16377 , RIfec38b8_8345);
and \g451180/U$3 ( \21748 , RIf153cf8_5413, \16380 );
nor \g451180/U$1 ( \21749 , \21747 , \21748 );
and \g451178/U$2 ( \21750 , \16313 , RIfc53be8_5975);
and \g451178/U$3 ( \21751 , RIf157100_5450, \16321 );
nor \g451178/U$1 ( \21752 , \21750 , \21751 );
and \g445029/U$2 ( \21753 , \21746 , \21749 , \21752 );
nor \g445029/U$1 ( \21754 , \21753 , \16480 );
and \g445839/U$2 ( \21755 , RIf147548_5271, \16427 );
and \g445839/U$3 ( \21756 , RIfe91b60_8002, \16368 );
and \g448670/U$2 ( \21757 , RIfc9d220_6810, \16321 );
and \g448670/U$3 ( \21758 , \16328 , RIfcda4e0_7506);
and \g448670/U$4 ( \21759 , RIfc9f548_6835, \16398 );
nor \g448670/U$1 ( \21760 , \21757 , \21758 , \21759 );
and \g454703/U$2 ( \21761 , \16317 , RIfce16c8_7587);
and \g454703/U$3 ( \21762 , RIfc4f2c8_5923, \16325 );
nor \g454703/U$1 ( \21763 , \21761 , \21762 );
not \g449699/U$3 ( \21764 , \21763 );
not \g449699/U$4 ( \21765 , \16330 );
and \g449699/U$2 ( \21766 , \21764 , \21765 );
and \g449699/U$5 ( \21767 , \16341 , RIf146b70_5264);
nor \g449699/U$1 ( \21768 , \21766 , \21767 );
and \g451191/U$2 ( \21769 , \16377 , RIe1b6738_3453);
and \g451191/U$3 ( \21770 , RIe1b8628_3475, \16313 );
nor \g451191/U$1 ( \21771 , \21769 , \21770 );
and \g451192/U$2 ( \21772 , \16334 , RIfe91e30_8004);
and \g451192/U$3 ( \21773 , RIfe91cc8_8003, \16380 );
nor \g451192/U$1 ( \21774 , \21772 , \21773 );
nand \g447267/U$1 ( \21775 , \21760 , \21768 , \21771 , \21774 );
nor \g445839/U$1 ( \21776 , \21755 , \21756 , \21775 );
and \g451187/U$2 ( \21777 , \16361 , RIfe919f8_8001);
and \g451187/U$3 ( \21778 , RIf1484c0_5282, \16448 );
nor \g451187/U$1 ( \21779 , \21777 , \21778 );
and \g451186/U$2 ( \21780 , \16364 , RIfe92100_8006);
and \g451186/U$3 ( \21781 , RIfe91f98_8005, \16371 );
nor \g451186/U$1 ( \21782 , \21780 , \21781 );
and \g445031/U$2 ( \21783 , \21776 , \21779 , \21782 );
nor \g445031/U$1 ( \21784 , \21783 , \16909 );
or \g444328/U$1 ( \21785 , \21665 , \21725 , \21754 , \21784 );
and \g445834/U$2 ( \21786 , RIe1ce450_3724, \16427 );
and \g445834/U$3 ( \21787 , RIe1c8a50_3660, \16368 );
and \g448662/U$2 ( \21788 , RIe1e7950_4012, \16321 );
and \g448662/U$3 ( \21789 , \16326 , RIe1ea650_4044);
and \g448662/U$4 ( \21790 , RIe1c3050_3596, \16337 );
nor \g448662/U$1 ( \21791 , \21788 , \21789 , \21790 );
and \g454841/U$2 ( \21792 , \16317 , RIe1dc550_3884);
and \g454841/U$3 ( \21793 , RIe1df250_3916, \16325 );
nor \g454841/U$1 ( \21794 , \21792 , \21793 );
not \g449690/U$3 ( \21795 , \21794 );
not \g449690/U$4 ( \21796 , \16330 );
and \g449690/U$2 ( \21797 , \21795 , \21796 );
and \g449690/U$5 ( \21798 , \16341 , RIe1c5d50_3628);
nor \g449690/U$1 ( \21799 , \21797 , \21798 );
and \g451164/U$2 ( \21800 , \16377 , RIe1e1f50_3948);
and \g451164/U$3 ( \21801 , RIe1e4c50_3980, \16313 );
nor \g451164/U$1 ( \21802 , \21800 , \21801 );
and \g451165/U$2 ( \21803 , \16334 , RIe1d6b50_3820);
and \g451165/U$3 ( \21804 , RIe1d9850_3852, \16380 );
nor \g451165/U$1 ( \21805 , \21803 , \21804 );
nand \g447264/U$1 ( \21806 , \21791 , \21799 , \21802 , \21805 );
nor \g445834/U$1 ( \21807 , \21786 , \21787 , \21806 );
and \g451161/U$2 ( \21808 , \16361 , RIe1bd650_3532);
and \g451161/U$3 ( \21809 , RIe1d1150_3756, \16448 );
nor \g451161/U$1 ( \21810 , \21808 , \21809 );
and \g451160/U$2 ( \21811 , \16364 , RIe1c0350_3564);
and \g451160/U$3 ( \21812 , RIe1cb750_3692, \16371 );
nor \g451160/U$1 ( \21813 , \21811 , \21812 );
and \g445026/U$2 ( \21814 , \21807 , \21810 , \21813 );
nor \g445026/U$1 ( \21815 , \21814 , \16555 );
and \g445835/U$2 ( \21816 , RIe1fda48_4263, \16427 );
and \g445835/U$3 ( \21817 , RIe1ef948_4103, \16368 );
and \g448665/U$2 ( \21818 , RIe177c90_2740, \16344 );
and \g448665/U$3 ( \21819 , \16354 , RIe18b790_2964);
and \g448665/U$4 ( \21820 , RIe1ba950_3500, \16337 );
nor \g448665/U$1 ( \21821 , \21818 , \21819 , \21820 );
and \g454788/U$2 ( \21822 , \16317 , RIe1a4c90_3252);
and \g454788/U$3 ( \21823 , RIe1a7990_3284, \16325 );
nor \g454788/U$1 ( \21824 , \21822 , \21823 );
not \g449693/U$3 ( \21825 , \21824 );
not \g449693/U$4 ( \21826 , \16311 );
and \g449693/U$2 ( \21827 , \21825 , \21826 );
and \g449693/U$5 ( \21828 , \16339 , RIe1d3e50_3788);
nor \g449693/U$1 ( \21829 , \21827 , \21828 );
and \g451173/U$2 ( \21830 , \16377 , RIe19f290_3188);
and \g451173/U$3 ( \21831 , RIe1a1f90_3220, \16313 );
nor \g451173/U$1 ( \21832 , \21830 , \21831 );
and \g451174/U$2 ( \21833 , \16334 , RIe21a1e8_4587);
and \g451174/U$3 ( \21834 , RIe2255e8_4715, \16380 );
nor \g451174/U$1 ( \21835 , \21833 , \21834 );
nand \g447265/U$1 ( \21836 , \21821 , \21829 , \21832 , \21835 );
nor \g445835/U$1 ( \21837 , \21816 , \21817 , \21836 );
and \g451171/U$2 ( \21838 , \16361 , RIe16fe00_2650);
and \g451171/U$3 ( \21839 , RIe2039e8_4331, \16448 );
nor \g451171/U$1 ( \21840 , \21838 , \21839 );
and \g451169/U$2 ( \21841 , \16364 , RIe1ad7c8_3351);
and \g451169/U$3 ( \21842 , RIe1f6e00_4186, \16371 );
nor \g451169/U$1 ( \21843 , \21841 , \21842 );
and \g445028/U$2 ( \21844 , \21837 , \21840 , \21843 );
nor \g445028/U$1 ( \21845 , \21844 , \16586 );
or \g444223/U$1 ( \21846 , \21785 , \21815 , \21845 );
_DC \g3e4b/U$1 ( \21847 , \21846 , \16652 );
and \g450552/U$2 ( \21848 , \16364 , RIf16eb48_5719);
and \g450552/U$3 ( \21849 , RIee3a660_5123, \16371 );
nor \g450552/U$1 ( \21850 , \21848 , \21849 );
and \g445702/U$2 ( \21851 , RIee3b740_5135, \16427 );
and \g445702/U$3 ( \21852 , RIe174e28_2707, \16368 );
and \g448494/U$2 ( \21853 , RIfe8ff40_7982, \16321 );
and \g448494/U$3 ( \21854 , \16328 , RIfe90210_7984);
and \g448494/U$4 ( \21855 , RIfc5fdf8_6113, \16398 );
nor \g448494/U$1 ( \21856 , \21853 , \21854 , \21855 );
and \g454744/U$2 ( \21857 , \16317 , RIfc61040_6126);
and \g454744/U$3 ( \21858 , RIfcaf6a0_7018, \16325 );
nor \g454744/U$1 ( \21859 , \21857 , \21858 );
not \g449515/U$3 ( \21860 , \21859 );
not \g449515/U$4 ( \21861 , \16330 );
and \g449515/U$2 ( \21862 , \21860 , \21861 );
and \g449515/U$5 ( \21863 , \16341 , RIf170768_5739);
nor \g449515/U$1 ( \21864 , \21862 , \21863 );
and \g450554/U$2 ( \21865 , \16377 , RIe176a48_2727);
and \g450554/U$3 ( \21866 , RIfc72f20_6330, \16313 );
nor \g450554/U$1 ( \21867 , \21865 , \21866 );
and \g450555/U$2 ( \21868 , \16334 , RIfe900a8_7983);
and \g450555/U$3 ( \21869 , RIf13e8a8_5171, \16380 );
nor \g450555/U$1 ( \21870 , \21868 , \21869 );
nand \g447232/U$1 ( \21871 , \21856 , \21864 , \21867 , \21870 );
nor \g445702/U$1 ( \21872 , \21851 , \21852 , \21871 );
and \g450553/U$2 ( \21873 , \16361 , RIfcaaab0_6964);
and \g450553/U$3 ( \21874 , RIee3caf0_5149, \16448 );
nor \g450553/U$1 ( \21875 , \21873 , \21874 );
nand \g445506/U$1 ( \21876 , \21850 , \21872 , \21875 );
and \g444698/U$2 ( \21877 , \21876 , \17998 );
and \g448492/U$2 ( \21878 , RIe19c2c0_3154, \16321 );
and \g448492/U$3 ( \21879 , \16328 , RIe19efc0_3186);
and \g448492/U$4 ( \21880 , RIe182dc0_2866, \16337 );
nor \g448492/U$1 ( \21881 , \21878 , \21879 , \21880 );
and \g454365/U$2 ( \21882 , \16317 , RIe1968c0_3090);
and \g454365/U$3 ( \21883 , RIfc637a0_6154, \16325 );
nor \g454365/U$1 ( \21884 , \21882 , \21883 );
not \g449513/U$3 ( \21885 , \21884 );
not \g449513/U$4 ( \21886 , \16330 );
and \g449513/U$2 ( \21887 , \21885 , \21886 );
and \g449513/U$5 ( \21888 , \16339 , RIfe8fc70_7980);
nor \g449513/U$1 ( \21889 , \21887 , \21888 );
and \g450548/U$2 ( \21890 , \16377 , RIe1995c0_3122);
and \g450548/U$3 ( \21891 , RIf145d60_5254, \16313 );
nor \g450548/U$1 ( \21892 , \21890 , \21891 );
and \g450549/U$2 ( \21893 , \16334 , RIe190ec0_3026);
and \g450549/U$3 ( \21894 , RIe193bc0_3058, \16380 );
nor \g450549/U$1 ( \21895 , \21893 , \21894 );
nand \g447231/U$1 ( \21896 , \21881 , \21889 , \21892 , \21895 );
and \g444698/U$3 ( \21897 , \17938 , \21896 );
nor \g444698/U$1 ( \21898 , \21877 , \21897 );
and \g446500/U$2 ( \21899 , \18457 , RIe1887c0_2930);
and \g446500/U$3 ( \21900 , RIe18b4c0_2962, \18459 );
nor \g446500/U$1 ( \21901 , \21899 , \21900 );
and \g446501/U$2 ( \21902 , \18462 , RIe185ac0_2898);
and \g446501/U$3 ( \21903 , RIfc62af8_6145, \18464 );
nor \g446501/U$1 ( \21904 , \21902 , \21903 );
and \g446502/U$2 ( \21905 , \18467 , RIe17d3c0_2802);
and \g446502/U$3 ( \21906 , RIe1800c0_2834, \18469 );
nor \g446502/U$1 ( \21907 , \21905 , \21906 );
nand \g444445/U$1 ( \21908 , \21898 , \21901 , \21904 , \21907 );
and \g450568/U$2 ( \21909 , \16364 , RIe1b01f8_3381);
and \g450568/U$3 ( \21910 , RIe1f9830_4216, \16371 );
nor \g450568/U$1 ( \21911 , \21909 , \21910 );
and \g445705/U$2 ( \21912 , RIe200478_4293, \16427 );
and \g445705/U$3 ( \21913 , RIe1f2378_4133, \16368 );
and \g448497/U$2 ( \21914 , RIe1a76c0_3282, \16321 );
and \g448497/U$3 ( \21915 , \16328 , RIe1aa3c0_3314);
and \g448497/U$4 ( \21916 , RIe1bd380_3530, \16337 );
nor \g448497/U$1 ( \21917 , \21914 , \21915 , \21916 );
and \g454521/U$2 ( \21918 , \16317 , RIe17a6c0_2770);
and \g454521/U$3 ( \21919 , RIe18e1c0_2994, \16325 );
nor \g454521/U$1 ( \21920 , \21918 , \21919 );
not \g449521/U$3 ( \21921 , \21920 );
not \g449521/U$4 ( \21922 , \16330 );
and \g449521/U$2 ( \21923 , \21921 , \21922 );
and \g449521/U$5 ( \21924 , \16341 , RIe1d6880_3818);
nor \g449521/U$1 ( \21925 , \21923 , \21924 );
and \g450571/U$2 ( \21926 , \16377 , RIe1a1cc0_3218);
and \g450571/U$3 ( \21927 , RIe1a49c0_3250, \16313 );
nor \g450571/U$1 ( \21928 , \21926 , \21927 );
and \g450574/U$2 ( \21929 , \16334 , RIe21cc18_4617);
and \g450574/U$3 ( \21930 , RIe228018_4745, \16380 );
nor \g450574/U$1 ( \21931 , \21929 , \21930 );
nand \g447233/U$1 ( \21932 , \21917 , \21925 , \21928 , \21931 );
nor \g445705/U$1 ( \21933 , \21912 , \21913 , \21932 );
and \g450569/U$2 ( \21934 , \16361 , RIe172830_2680);
and \g450569/U$3 ( \21935 , RIe206418_4361, \16448 );
nor \g450569/U$1 ( \21936 , \21934 , \21935 );
nand \g445507/U$1 ( \21937 , \21911 , \21933 , \21936 );
and \g444751/U$2 ( \21938 , \21937 , \16752 );
and \g448496/U$2 ( \21939 , RIe1c5a80_3626, \16337 );
and \g448496/U$3 ( \21940 , \16341 , RIe1c8780_3658);
and \g448496/U$4 ( \21941 , RIe1def80_3914, \16485 );
nor \g448496/U$1 ( \21942 , \21939 , \21940 , \21941 );
and \g454476/U$2 ( \21943 , \16317 , RIe1d0e80_3754);
and \g454476/U$3 ( \21944 , RIe1d3b80_3786, \16325 );
nor \g454476/U$1 ( \21945 , \21943 , \21944 );
not \g449518/U$3 ( \21946 , \21945 );
not \g449518/U$4 ( \21947 , \16351 );
and \g449518/U$2 ( \21948 , \21946 , \21947 );
and \g449518/U$5 ( \21949 , \16356 , RIe1e1c80_3946);
nor \g449518/U$1 ( \21950 , \21948 , \21949 );
and \g450564/U$2 ( \21951 , \16361 , RIe1c0080_3562);
and \g450564/U$3 ( \21952 , RIe1c2d80_3594, \16364 );
nor \g450564/U$1 ( \21953 , \21951 , \21952 );
and \g450562/U$2 ( \21954 , \16368 , RIe1cb480_3690);
and \g450562/U$3 ( \21955 , RIe1ce180_3722, \16371 );
nor \g450562/U$1 ( \21956 , \21954 , \21955 );
nand \g447455/U$1 ( \21957 , \21942 , \21950 , \21953 , \21956 );
and \g444751/U$3 ( \21958 , \16750 , \21957 );
nor \g444751/U$1 ( \21959 , \21938 , \21958 );
and \g446507/U$2 ( \21960 , \19457 , RIe1ea380_4042);
and \g446507/U$3 ( \21961 , RIe1ed080_4074, \19459 );
nor \g446507/U$1 ( \21962 , \21960 , \21961 );
and \g446509/U$2 ( \21963 , \19462 , RIe1d9580_3850);
and \g446509/U$3 ( \21964 , RIe1dc280_3882, \19464 );
nor \g446509/U$1 ( \21965 , \21963 , \21964 );
and \g446508/U$2 ( \21966 , \19467 , RIe1e4980_3978);
and \g446508/U$3 ( \21967 , RIe1e7680_4010, \19469 );
nor \g446508/U$1 ( \21968 , \21966 , \21967 );
nand \g444549/U$1 ( \21969 , \21959 , \21962 , \21965 , \21968 );
and \g446497/U$2 ( \21970 , RIe225318_4713, \16319 );
and \g446497/U$3 ( \21971 , RIf16c6b8_5693, \16313 );
and \g449512/U$2 ( \21972 , RIe20eb18_4457, \16398 );
and \g449512/U$3 ( \21973 , \16341 , RIfca5a88_6907);
and \g449512/U$4 ( \21974 , RIe21f918_4649, \16344 );
nor \g449512/U$1 ( \21975 , \21972 , \21973 , \21974 );
and \g454868/U$2 ( \21976 , \16317 , RIe214518_4521);
and \g454868/U$3 ( \21977 , RIfca62f8_6913, \16325 );
nor \g454868/U$1 ( \21978 , \21976 , \21977 );
not \g450533/U$3 ( \21979 , \21978 );
not \g450533/U$4 ( \21980 , \16351 );
and \g450533/U$2 ( \21981 , \21979 , \21980 );
and \g450533/U$5 ( \21982 , \16356 , RIf16b5d8_5681);
nor \g450533/U$1 ( \21983 , \21981 , \21982 );
and \g454120/U$2 ( \21984 , \16361 , RIe209118_4393);
and \g454120/U$3 ( \21985 , RIe20be18_4425, \16364 );
nor \g454120/U$1 ( \21986 , \21984 , \21985 );
and \g454119/U$2 ( \21987 , \16368 , RIe211818_4489);
and \g454119/U$3 ( \21988 , RIfcc9578_7313, \16371 );
nor \g454119/U$1 ( \21989 , \21987 , \21988 );
nand \g448002/U$1 ( \21990 , \21975 , \21983 , \21986 , \21989 );
nor \g446497/U$1 ( \21991 , \21970 , \21971 , \21990 );
and \g454117/U$2 ( \21992 , \16377 , RIe222618_4681);
and \g454117/U$3 ( \21993 , RIe219f18_4585, \16380 );
nor \g454117/U$1 ( \21994 , \21992 , \21993 );
and \g454116/U$2 ( \21995 , \16334 , RIe217218_4553);
and \g454116/U$3 ( \21996 , RIf16d1f8_5701, \16326 );
nor \g454116/U$1 ( \21997 , \21995 , \21996 );
and \g445499/U$2 ( \21998 , \21991 , \21994 , \21997 );
nor \g445499/U$1 ( \21999 , \21998 , \16389 );
and \g446499/U$2 ( \22000 , RIf15f260_5542, \16427 );
and \g446499/U$3 ( \22001 , RIe1fc530_4248, \16368 );
and \g448489/U$2 ( \22002 , RIf164990_5604, \16485 );
and \g448489/U$3 ( \22003 , \16356 , RIf165638_5613);
and \g448489/U$4 ( \22004 , RIf15c290_5508, \16337 );
nor \g448489/U$1 ( \22005 , \22002 , \22003 , \22004 );
and \g454827/U$2 ( \22006 , \16317 , RIf166718_5625);
and \g454827/U$3 ( \22007 , RIf167690_5636, \16325 );
nor \g454827/U$1 ( \22008 , \22006 , \22007 );
not \g450536/U$3 ( \22009 , \22008 );
not \g450536/U$4 ( \22010 , \16311 );
and \g450536/U$2 ( \22011 , \22009 , \22010 );
and \g450536/U$5 ( \22012 , \16341 , RIf15d4d8_5521);
nor \g450536/U$1 ( \22013 , \22011 , \22012 );
and \g454130/U$2 ( \22014 , \16377 , RIfe8f838_7977);
and \g454130/U$3 ( \22015 , RIfe8f9a0_7978, \16313 );
nor \g454130/U$1 ( \22016 , \22014 , \22015 );
and \g454131/U$2 ( \22017 , \16334 , RIf1627d0_5580);
and \g454131/U$3 ( \22018 , RIf1638b0_5592, \16380 );
nor \g454131/U$1 ( \22019 , \22017 , \22018 );
nand \g447452/U$1 ( \22020 , \22005 , \22013 , \22016 , \22019 );
nor \g446499/U$1 ( \22021 , \22000 , \22001 , \22020 );
and \g454126/U$2 ( \22022 , \16361 , RIf159f68_5483);
and \g454126/U$3 ( \22023 , RIf161150_5564, \16448 );
nor \g454126/U$1 ( \22024 , \22022 , \22023 );
and \g454125/U$2 ( \22025 , \16364 , RIfca20e0_6866);
and \g454125/U$3 ( \22026 , RIe1fd778_4261, \16371 );
nor \g454125/U$1 ( \22027 , \22025 , \22026 );
and \g445502/U$2 ( \22028 , \22021 , \22024 , \22027 );
nor \g445502/U$1 ( \22029 , \22028 , \16393 );
or \g444349/U$1 ( \22030 , \21908 , \21969 , \21999 , \22029 );
and \g446493/U$2 ( \22031 , RIf1581e0_5462, \16321 );
and \g446493/U$3 ( \22032 , RIfc5ebb0_6100, \16313 );
and \g449506/U$2 ( \22033 , RIfcb1158_7037, \16398 );
and \g449506/U$3 ( \22034 , \16341 , RIfcebe20_7706);
and \g449506/U$4 ( \22035 , RIfc5e8e0_6098, \16485 );
nor \g449506/U$1 ( \22036 , \22033 , \22034 , \22035 );
and \g455366/U$2 ( \22037 , \16317 , RIf1523a8_5395);
and \g455366/U$3 ( \22038 , RIf153b90_5412, \16325 );
nor \g455366/U$1 ( \22039 , \22037 , \22038 );
not \g450529/U$3 ( \22040 , \22039 );
not \g450529/U$4 ( \22041 , \16351 );
and \g450529/U$2 ( \22042 , \22040 , \22041 );
and \g450529/U$5 ( \22043 , \16356 , RIfc69e48_6227);
nor \g450529/U$1 ( \22044 , \22042 , \22043 );
and \g454103/U$2 ( \22045 , \16361 , RIe1ef678_4101);
and \g454103/U$3 ( \22046 , RIf14e730_5352, \16364 );
nor \g454103/U$1 ( \22047 , \22045 , \22046 );
and \g454102/U$2 ( \22048 , \16368 , RIfe8fb08_7979);
and \g454102/U$3 ( \22049 , RIfce88b0_7668, \16371 );
nor \g454102/U$1 ( \22050 , \22048 , \22049 );
nand \g448000/U$1 ( \22051 , \22036 , \22044 , \22047 , \22050 );
nor \g446493/U$1 ( \22052 , \22031 , \22032 , \22051 );
and \g454101/U$2 ( \22053 , \16377 , RIfe8fdd8_7981);
and \g454101/U$3 ( \22054 , RIf154f40_5426, \16380 );
nor \g454101/U$1 ( \22055 , \22053 , \22054 );
and \g454100/U$2 ( \22056 , \16334 , RIe1f6b30_4184);
and \g454100/U$3 ( \22057 , RIf159428_5475, \16328 );
nor \g454100/U$1 ( \22058 , \22056 , \22057 );
and \g445495/U$2 ( \22059 , \22052 , \22055 , \22058 );
nor \g445495/U$1 ( \22060 , \22059 , \16480 );
and \g446495/U$2 ( \22061 , RIf148358_5281, \16427 );
and \g446495/U$3 ( \22062 , RIfec3480_8342, \16368 );
and \g449508/U$2 ( \22063 , RIfc5ce28_6079, \16344 );
and \g449508/U$3 ( \22064 , \16356 , RIfc5cf90_6080);
and \g449508/U$4 ( \22065 , RIfc80be8_6487, \16398 );
nor \g449508/U$1 ( \22066 , \22063 , \22064 , \22065 );
and \g454914/U$2 ( \22067 , \16317 , RIfc5d698_6085);
and \g454914/U$3 ( \22068 , RIfcc8ba0_7306, \16325 );
nor \g454914/U$1 ( \22069 , \22067 , \22068 );
not \g450531/U$3 ( \22070 , \22069 );
not \g450531/U$4 ( \22071 , \16311 );
and \g450531/U$2 ( \22072 , \22070 , \22071 );
and \g450531/U$5 ( \22073 , \16341 , RIfc483b0_5844);
nor \g450531/U$1 ( \22074 , \22072 , \22073 );
and \g454110/U$2 ( \22075 , \16377 , RIfeabd08_8271);
and \g454110/U$3 ( \22076 , RIfec35e8_8343, \16313 );
nor \g454110/U$1 ( \22077 , \22075 , \22076 );
and \g454111/U$2 ( \22078 , \16334 , RIe1b4b18_3433);
and \g454111/U$3 ( \22079 , RIfec31b0_8340, \16380 );
nor \g454111/U$1 ( \22080 , \22078 , \22079 );
nand \g447450/U$1 ( \22081 , \22066 , \22074 , \22077 , \22080 );
nor \g446495/U$1 ( \22082 , \22061 , \22062 , \22081 );
and \g454108/U$2 ( \22083 , \16361 , RIfec3318_8341);
and \g454108/U$3 ( \22084 , RIf149708_5295, \16432 );
nor \g454108/U$1 ( \22085 , \22083 , \22084 );
and \g454107/U$2 ( \22086 , \16364 , RIe1ad4f8_3349);
and \g454107/U$3 ( \22087 , RIe1b3768_3419, \16371 );
nor \g454107/U$1 ( \22088 , \22086 , \22087 );
and \g445497/U$2 ( \22089 , \22082 , \22085 , \22088 );
nor \g445497/U$1 ( \22090 , \22089 , \16909 );
or \g444182/U$1 ( \22091 , \22030 , \22060 , \22090 );
_DC \g3ed0/U$1 ( \22092 , \22091 , \16652 );
and \g450724/U$2 ( \22093 , \16364 , RIfcc65a8_7279);
and \g450724/U$3 ( \22094 , RIfc815c0_6494, \16371 );
nor \g450724/U$1 ( \22095 , \22093 , \22094 );
and \g445739/U$2 ( \22096 , RIfce08b8_7577, \16427 );
and \g445739/U$3 ( \22097 , RIe174cc0_2706, \16368 );
and \g448540/U$2 ( \22098 , RIfc9ff20_6842, \16485 );
and \g448540/U$3 ( \22099 , \16356 , RIfc81e30_6500);
and \g448540/U$4 ( \22100 , RIfc53eb8_5977, \16398 );
nor \g448540/U$1 ( \22101 , \22098 , \22099 , \22100 );
and \g454228/U$2 ( \22102 , \16317 , RIfe8efc8_7971);
and \g454228/U$3 ( \22103 , RIf1427f0_5216, \16325 );
nor \g454228/U$1 ( \22104 , \22102 , \22103 );
not \g449565/U$3 ( \22105 , \22104 );
not \g449565/U$4 ( \22106 , \16311 );
and \g449565/U$2 ( \22107 , \22105 , \22106 );
and \g449565/U$5 ( \22108 , \16341 , RIfca04c0_6846);
nor \g449565/U$1 ( \22109 , \22107 , \22108 );
and \g450729/U$2 ( \22110 , \16377 , RIe1768e0_2726);
and \g450729/U$3 ( \22111 , RIe1779c0_2738, \16313 );
nor \g450729/U$1 ( \22112 , \22110 , \22111 );
and \g450730/U$2 ( \22113 , \16334 , RIfc81b60_6498);
and \g450730/U$3 ( \22114 , RIfca0088_6843, \16380 );
nor \g450730/U$1 ( \22115 , \22113 , \22114 );
nand \g447246/U$1 ( \22116 , \22101 , \22109 , \22112 , \22115 );
nor \g445739/U$1 ( \22117 , \22096 , \22097 , \22116 );
and \g450725/U$2 ( \22118 , \16361 , RIfc80d50_6488);
and \g450725/U$3 ( \22119 , RIfce5778_7633, \16448 );
nor \g450725/U$1 ( \22120 , \22118 , \22119 );
nand \g445515/U$1 ( \22121 , \22095 , \22117 , \22120 );
and \g444701/U$2 ( \22122 , \22121 , \17998 );
and \g448539/U$2 ( \22123 , RIe19c158_3153, \16321 );
and \g448539/U$3 ( \22124 , \16328 , RIe19ee58_3185);
and \g448539/U$4 ( \22125 , RIe182c58_2865, \16398 );
nor \g448539/U$1 ( \22126 , \22123 , \22124 , \22125 );
and \g454226/U$2 ( \22127 , \16317 , RIe196758_3089);
and \g454226/U$3 ( \22128 , RIfe8f298_7973, \16325 );
nor \g454226/U$1 ( \22129 , \22127 , \22128 );
not \g449562/U$3 ( \22130 , \22129 );
not \g449562/U$4 ( \22131 , \16330 );
and \g449562/U$2 ( \22132 , \22130 , \22131 );
and \g449562/U$5 ( \22133 , \16341 , RIfc9f278_6833);
nor \g449562/U$1 ( \22134 , \22132 , \22133 );
and \g450721/U$2 ( \22135 , \16377 , RIe199458_3121);
and \g450721/U$3 ( \22136 , RIf145bf8_5253, \16313 );
nor \g450721/U$1 ( \22137 , \22135 , \22136 );
and \g450722/U$2 ( \22138 , \16334 , RIe190d58_3025);
and \g450722/U$3 ( \22139 , RIe193a58_3057, \16380 );
nor \g450722/U$1 ( \22140 , \22138 , \22139 );
nand \g447245/U$1 ( \22141 , \22126 , \22134 , \22137 , \22140 );
and \g444701/U$3 ( \22142 , \17938 , \22141 );
nor \g444701/U$1 ( \22143 , \22122 , \22142 );
and \g446535/U$2 ( \22144 , \18457 , RIe188658_2929);
and \g446535/U$3 ( \22145 , RIe18b358_2961, \18459 );
nor \g446535/U$1 ( \22146 , \22144 , \22145 );
and \g446536/U$2 ( \22147 , \18462 , RIe185958_2897);
and \g446536/U$3 ( \22148 , RIfe8f130_7972, \18464 );
nor \g446536/U$1 ( \22149 , \22147 , \22148 );
and \g446537/U$2 ( \22150 , \18467 , RIe17d258_2801);
and \g446537/U$3 ( \22151 , RIe17ff58_2833, \18469 );
nor \g446537/U$1 ( \22152 , \22150 , \22151 );
nand \g444450/U$1 ( \22153 , \22143 , \22146 , \22149 , \22152 );
and \g450739/U$2 ( \22154 , \16377 , RIe1b84c0_3474);
and \g450739/U$3 ( \22155 , RIe1b6468_3451, \16380 );
nor \g450739/U$1 ( \22156 , \22154 , \22155 );
and \g445742/U$2 ( \22157 , RIfe8ee60_7970, \16319 );
and \g445742/U$3 ( \22158 , RIfea8090_8228, \16313 );
and \g448544/U$2 ( \22159 , RIfca8ff8_6945, \16398 );
and \g448544/U$3 ( \22160 , \16341 , RIfc67f58_6205);
and \g448544/U$4 ( \22161 , RIfc6c170_6252, \16485 );
nor \g448544/U$1 ( \22162 , \22159 , \22160 , \22161 );
and \g454918/U$2 ( \22163 , \16317 , RIfcaa948_6963);
and \g454918/U$3 ( \22164 , RIfcafad8_7021, \16325 );
nor \g454918/U$1 ( \22165 , \22163 , \22164 );
not \g449569/U$3 ( \22166 , \22165 );
not \g449569/U$4 ( \22167 , \16351 );
and \g449569/U$2 ( \22168 , \22166 , \22167 );
and \g449569/U$5 ( \22169 , \16356 , RIf14aab8_5309);
nor \g449569/U$1 ( \22170 , \22168 , \22169 );
and \g450745/U$2 ( \22171 , \16361 , RIe1abe78_3333);
and \g450745/U$3 ( \22172 , RIfe8eb90_7968, \16364 );
nor \g450745/U$1 ( \22173 , \22171 , \22172 );
and \g450744/U$2 ( \22174 , \16368 , RIfe8f400_7974);
and \g450744/U$3 ( \22175 , RIfe8ecf8_7969, \16371 );
nor \g450744/U$1 ( \22176 , \22174 , \22175 );
nand \g447482/U$1 ( \22177 , \22162 , \22170 , \22173 , \22176 );
nor \g445742/U$1 ( \22178 , \22157 , \22158 , \22177 );
and \g450738/U$2 ( \22179 , \16334 , RIe1b49b0_3432);
and \g450738/U$3 ( \22180 , RIf14d218_5337, \16328 );
nor \g450738/U$1 ( \22181 , \22179 , \22180 );
nand \g445517/U$1 ( \22182 , \22156 , \22178 , \22181 );
and \g444904/U$2 ( \22183 , \22182 , \16477 );
and \g448543/U$2 ( \22184 , RIfc55c40_5998, \16321 );
and \g448543/U$3 ( \22185 , \16326 , RIfc4bd58_5885);
and \g448543/U$4 ( \22186 , RIfc90908_6667, \16398 );
nor \g448543/U$1 ( \22187 , \22184 , \22185 , \22186 );
and \g454230/U$2 ( \22188 , \16317 , RIfcd5ff8_7457);
and \g454230/U$3 ( \22189 , RIf156890_5444, \16325 );
nor \g454230/U$1 ( \22190 , \22188 , \22189 );
not \g449567/U$3 ( \22191 , \22190 );
not \g449567/U$4 ( \22192 , \16330 );
and \g449567/U$2 ( \22193 , \22191 , \22192 );
and \g449567/U$5 ( \22194 , \16341 , RIfc44738_5801);
nor \g449567/U$1 ( \22195 , \22193 , \22194 );
and \g450734/U$2 ( \22196 , \16377 , RIe1fb450_4236);
and \g450734/U$3 ( \22197 , RIfca2ab8_6873, \16313 );
nor \g450734/U$1 ( \22198 , \22196 , \22197 );
and \g450736/U$2 ( \22199 , \16334 , RIfec2aa8_8335);
and \g450736/U$3 ( \22200 , RIf154dd8_5425, \16380 );
nor \g450736/U$1 ( \22201 , \22199 , \22200 );
nand \g447247/U$1 ( \22202 , \22187 , \22195 , \22198 , \22201 );
and \g444904/U$3 ( \22203 , \16481 , \22202 );
nor \g444904/U$1 ( \22204 , \22183 , \22203 );
and \g446541/U$2 ( \22205 , \17274 , RIfcd9400_7494);
and \g446541/U$3 ( \22206 , RIfcb4b00_7078, \17276 );
nor \g446541/U$1 ( \22207 , \22205 , \22206 );
and \g446542/U$2 ( \22208 , \17279 , RIe1f4808_4159);
and \g446542/U$3 ( \22209 , RIf151160_5382, \17281 );
nor \g446542/U$1 ( \22210 , \22208 , \22209 );
and \g446543/U$2 ( \22211 , \17284 , RIe1ef510_4100);
and \g446543/U$3 ( \22212 , RIf14e5c8_5351, \17286 );
nor \g446543/U$1 ( \22213 , \22211 , \22212 );
nand \g444554/U$1 ( \22214 , \22204 , \22207 , \22210 , \22213 );
and \g445734/U$2 ( \22215 , RIe1d0d18_3753, \16427 );
and \g445734/U$3 ( \22216 , RIe1cb318_3689, \16368 );
and \g448535/U$2 ( \22217 , RIe1ea218_4041, \16319 );
and \g448535/U$3 ( \22218 , \16328 , RIe1ecf18_4073);
and \g448535/U$4 ( \22219 , RIe1c5918_3625, \16398 );
nor \g448535/U$1 ( \22220 , \22217 , \22218 , \22219 );
and \g454177/U$2 ( \22221 , \16317 , RIe1dee18_3913);
and \g454177/U$3 ( \22222 , RIe1e1b18_3945, \16325 );
nor \g454177/U$1 ( \22223 , \22221 , \22222 );
not \g449559/U$3 ( \22224 , \22223 );
not \g449559/U$4 ( \22225 , \16330 );
and \g449559/U$2 ( \22226 , \22224 , \22225 );
and \g449559/U$5 ( \22227 , \16341 , RIe1c8618_3657);
nor \g449559/U$1 ( \22228 , \22226 , \22227 );
and \g450709/U$2 ( \22229 , \16377 , RIe1e4818_3977);
and \g450709/U$3 ( \22230 , RIe1e7518_4009, \16313 );
nor \g450709/U$1 ( \22231 , \22229 , \22230 );
and \g450711/U$2 ( \22232 , \16334 , RIe1d9418_3849);
and \g450711/U$3 ( \22233 , RIe1dc118_3881, \16380 );
nor \g450711/U$1 ( \22234 , \22232 , \22233 );
nand \g447244/U$1 ( \22235 , \22220 , \22228 , \22231 , \22234 );
nor \g445734/U$1 ( \22236 , \22215 , \22216 , \22235 );
and \g450708/U$2 ( \22237 , \16361 , RIe1bff18_3561);
and \g450708/U$3 ( \22238 , RIe1d3a18_3785, \16448 );
nor \g450708/U$1 ( \22239 , \22237 , \22238 );
and \g450707/U$2 ( \22240 , \16364 , RIe1c2c18_3593);
and \g450707/U$3 ( \22241 , RIe1ce018_3721, \16371 );
nor \g450707/U$1 ( \22242 , \22240 , \22241 );
and \g444953/U$2 ( \22243 , \22236 , \22239 , \22242 );
nor \g444953/U$1 ( \22244 , \22243 , \16555 );
and \g445737/U$2 ( \22245 , RIe1a4858_3249, \16313 );
and \g445737/U$3 ( \22246 , RIe1726c8_2679, \16361 );
and \g448537/U$2 ( \22247 , RIe1a7558_3281, \16321 );
and \g448537/U$3 ( \22248 , \16485 , RIe17a558_2769);
and \g448537/U$4 ( \22249 , RIe18e058_2993, \16356 );
nor \g448537/U$1 ( \22250 , \22247 , \22248 , \22249 );
and \g450718/U$2 ( \22251 , \16368 , RIe1f2210_4132);
and \g450718/U$3 ( \22252 , RIe1f96c8_4215, \16371 );
nor \g450718/U$1 ( \22253 , \22251 , \22252 );
and \g454221/U$2 ( \22254 , \16317 , RIe200310_4292);
and \g454221/U$3 ( \22255 , RIe2062b0_4360, \16325 );
nor \g454221/U$1 ( \22256 , \22254 , \22255 );
not \g449561/U$3 ( \22257 , \22256 );
not \g449561/U$4 ( \22258 , \16351 );
and \g449561/U$2 ( \22259 , \22257 , \22258 );
and \g449561/U$5 ( \22260 , \16326 , RIe1aa258_3313);
nor \g449561/U$1 ( \22261 , \22259 , \22260 );
and \g453649/U$2 ( \22262 , \16334 , RIe21cab0_4616);
and \g453649/U$3 ( \22263 , RIe227eb0_4744, \16380 );
nor \g453649/U$1 ( \22264 , \22262 , \22263 );
nand \g447477/U$1 ( \22265 , \22250 , \22253 , \22261 , \22264 );
nor \g445737/U$1 ( \22266 , \22245 , \22246 , \22265 );
and \g450715/U$2 ( \22267 , \16364 , RIe1b0090_3380);
and \g450715/U$3 ( \22268 , RIe1d6718_3817, \16339 );
nor \g450715/U$1 ( \22269 , \22267 , \22268 );
and \g450713/U$2 ( \22270 , \16337 , RIe1bd218_3529);
and \g450713/U$3 ( \22271 , RIe1a1b58_3217, \16377 );
nor \g450713/U$1 ( \22272 , \22270 , \22271 );
and \g444954/U$2 ( \22273 , \22266 , \22269 , \22272 );
nor \g444954/U$1 ( \22274 , \22273 , \16586 );
or \g444350/U$1 ( \22275 , \22153 , \22214 , \22244 , \22274 );
and \g445732/U$2 ( \22276 , RIf1665b0_5624, \16321 );
and \g445732/U$3 ( \22277 , RIe203718_4329, \16313 );
and \g448531/U$2 ( \22278 , RIfc87998_6565, \16427 );
and \g448531/U$3 ( \22279 , \16448 , RIfc7e320_6458);
and \g448531/U$4 ( \22280 , RIfcc5360_7266, \16485 );
nor \g448531/U$1 ( \22281 , \22278 , \22279 , \22280 );
and \g454168/U$2 ( \22282 , \16317 , RIf15c128_5507);
and \g454168/U$3 ( \22283 , RIf15d370_5520, \16325 );
nor \g454168/U$1 ( \22284 , \22282 , \22283 );
not \g454167/U$1 ( \22285 , \22284 );
and \g449552/U$2 ( \22286 , \22285 , \16336 );
and \g449552/U$3 ( \22287 , RIfc9da90_6816, \16356 );
nor \g449552/U$1 ( \22288 , \22286 , \22287 );
and \g450695/U$2 ( \22289 , \16361 , RIfce7d70_7660);
and \g450695/U$3 ( \22290 , RIfcc5d38_7273, \16364 );
nor \g450695/U$1 ( \22291 , \22289 , \22290 );
and \g450694/U$2 ( \22292 , \16368 , RIe1fc3c8_4247);
and \g450694/U$3 ( \22293 , RIe1fd610_4260, \16371 );
nor \g450694/U$1 ( \22294 , \22292 , \22293 );
nand \g448008/U$1 ( \22295 , \22281 , \22288 , \22291 , \22294 );
nor \g445732/U$1 ( \22296 , \22276 , \22277 , \22295 );
and \g450692/U$2 ( \22297 , \16377 , RIe201c60_4310);
and \g450692/U$3 ( \22298 , RIf163748_5591, \16380 );
nor \g450692/U$1 ( \22299 , \22297 , \22298 );
and \g450691/U$2 ( \22300 , \16334 , RIf162668_5579);
and \g450691/U$3 ( \22301 , RIf167528_5635, \16328 );
nor \g450691/U$1 ( \22302 , \22300 , \22301 );
and \g444951/U$2 ( \22303 , \22296 , \22299 , \22302 );
nor \g444951/U$1 ( \22304 , \22303 , \16393 );
and \g445733/U$2 ( \22305 , RIe2143b0_4520, \16427 );
and \g445733/U$3 ( \22306 , RIe2116b0_4488, \16368 );
and \g448532/U$2 ( \22307 , RIe21f7b0_4648, \16485 );
and \g448532/U$3 ( \22308 , \16356 , RIfcb5910_7088);
and \g448532/U$4 ( \22309 , RIe20e9b0_4456, \16398 );
nor \g448532/U$1 ( \22310 , \22307 , \22308 , \22309 );
and \g454216/U$2 ( \22311 , \16317 , RIe2251b0_4712);
and \g454216/U$3 ( \22312 , RIfc804e0_6482, \16325 );
nor \g454216/U$1 ( \22313 , \22311 , \22312 );
not \g449554/U$3 ( \22314 , \22313 );
not \g449554/U$4 ( \22315 , \16311 );
and \g449554/U$2 ( \22316 , \22314 , \22315 );
and \g449554/U$5 ( \22317 , \16341 , RIfc7f6d0_6472);
nor \g449554/U$1 ( \22318 , \22316 , \22317 );
and \g454087/U$2 ( \22319 , \16377 , RIe2224b0_4680);
and \g454087/U$3 ( \22320 , RIfc80378_6481, \16313 );
nor \g454087/U$1 ( \22321 , \22319 , \22320 );
and \g450704/U$2 ( \22322 , \16334 , RIe2170b0_4552);
and \g450704/U$3 ( \22323 , RIe219db0_4584, \16380 );
nor \g450704/U$1 ( \22324 , \22322 , \22323 );
nand \g447243/U$1 ( \22325 , \22310 , \22318 , \22321 , \22324 );
nor \g445733/U$1 ( \22326 , \22305 , \22306 , \22325 );
and \g450699/U$2 ( \22327 , \16361 , RIe208fb0_4392);
and \g450699/U$3 ( \22328 , RIfca01f0_6844, \16448 );
nor \g450699/U$1 ( \22329 , \22327 , \22328 );
and \g450698/U$2 ( \22330 , \16364 , RIe20bcb0_4424);
and \g450698/U$3 ( \22331 , RIfc82c40_6510, \16371 );
nor \g450698/U$1 ( \22332 , \22330 , \22331 );
and \g444952/U$2 ( \22333 , \22326 , \22329 , \22332 );
nor \g444952/U$1 ( \22334 , \22333 , \16389 );
or \g444206/U$1 ( \22335 , \22275 , \22304 , \22334 );
_DC \g3f55/U$1 ( \22336 , \22335 , \16652 );
and \g453681/U$2 ( \22337 , \16368 , RIe1f46a0_4158);
and \g453681/U$3 ( \22338 , RIfca3e68_6887, \16485 );
nor \g453681/U$1 ( \22339 , \22337 , \22338 );
and \g446398/U$2 ( \22340 , RIfe9c420_8122, \16354 );
and \g446398/U$3 ( \22341 , RIe1f69c8_4183, \16334 );
and \g449395/U$2 ( \22342 , RIf152240_5394, \16427 );
and \g449395/U$3 ( \22343 , \16398 , RIfc43bf8_5793);
and \g449395/U$4 ( \22344 , RIfca6028_6911, \16341 );
nor \g449395/U$1 ( \22345 , \22342 , \22343 , \22344 );
and \g453684/U$2 ( \22346 , \16361 , RIe1ef3a8_4099);
and \g453684/U$3 ( \22347 , RIf14e460_5350, \16364 );
nor \g453684/U$1 ( \22348 , \22346 , \22347 );
and \g453683/U$2 ( \22349 , \16377 , RIe1fb2e8_4235);
and \g453683/U$3 ( \22350 , RIfcc01d0_7208, \16313 );
nor \g453683/U$1 ( \22351 , \22349 , \22350 );
and \g454927/U$2 ( \22352 , \16317 , RIfe9c2b8_8121);
and \g454927/U$3 ( \22353 , RIfec4290_8352, \16325 );
nor \g454927/U$1 ( \22354 , \22352 , \22353 );
not \g450415/U$3 ( \22355 , \22354 );
not \g450415/U$4 ( \22356 , \16311 );
and \g450415/U$2 ( \22357 , \22355 , \22356 );
and \g450415/U$5 ( \22358 , \16432 , RIf153a28_5411);
nor \g450415/U$1 ( \22359 , \22357 , \22358 );
nand \g447941/U$1 ( \22360 , \22345 , \22348 , \22351 , \22359 );
nor \g446398/U$1 ( \22361 , \22340 , \22341 , \22360 );
and \g453680/U$2 ( \22362 , \16371 , RIf150ff8_5381);
and \g453680/U$3 ( \22363 , RIf154c70_5424, \16380 );
nor \g453680/U$1 ( \22364 , \22362 , \22363 );
nand \g445680/U$1 ( \22365 , \22339 , \22361 , \22364 );
and \g444837/U$2 ( \22366 , \22365 , \16481 );
and \g449391/U$2 ( \22367 , RIf14be68_5323, \16321 );
and \g449391/U$3 ( \22368 , \16328 , RIfc4d6a8_5903);
and \g449391/U$4 ( \22369 , RIf1481f0_5280, \16427 );
nor \g449391/U$1 ( \22370 , \22367 , \22368 , \22369 );
and \g453677/U$2 ( \22371 , \16361 , RIe1abd10_3332);
and \g453677/U$3 ( \22372 , RIfe9bbb0_8116, \16364 );
nor \g453677/U$1 ( \22373 , \22371 , \22372 );
and \g453675/U$2 ( \22374 , \16377 , RIfe9be80_8118);
and \g453675/U$3 ( \22375 , RIe1ba680_3498, \16313 );
nor \g453675/U$1 ( \22376 , \22374 , \22375 );
and \g455128/U$2 ( \22377 , \16317 , RIfcbfac8_7203);
and \g455128/U$3 ( \22378 , RIfc69470_6220, \16325 );
nor \g455128/U$1 ( \22379 , \22377 , \22378 );
not \g455127/U$1 ( \22380 , \22379 );
and \g450412/U$2 ( \22381 , \22380 , \16336 );
and \g450412/U$3 ( \22382 , RIf1495a0_5294, \16448 );
nor \g450412/U$1 ( \22383 , \22381 , \22382 );
nand \g448118/U$1 ( \22384 , \22370 , \22373 , \22376 , \22383 );
and \g444837/U$3 ( \22385 , \16477 , \22384 );
nor \g444837/U$1 ( \22386 , \22366 , \22385 );
and \g447156/U$2 ( \22387 , \17473 , RIe1b1e18_3401);
and \g447156/U$3 ( \22388 , RIe1b3600_3418, \17475 );
nor \g447156/U$1 ( \22389 , \22387 , \22388 );
nor \g448300/U$1 ( \22390 , \16909 , \16484 );
and \g447155/U$2 ( \22391 , \22390 , RIfcd46a8_7439);
nor \g448279/U$1 ( \22392 , \16909 , \16355 );
and \g447155/U$3 ( \22393 , RIfc86e58_6557, \22392 );
nor \g447155/U$1 ( \22394 , \22391 , \22393 );
and \g447157/U$2 ( \22395 , \18278 , RIfe9bd18_8117);
and \g447157/U$3 ( \22396 , RIe1b6300_3450, \18280 );
nor \g447157/U$1 ( \22397 , \22395 , \22396 );
nand \g444658/U$1 ( \22398 , \22386 , \22389 , \22394 , \22397 );
and \g447151/U$2 ( \22399 , \18030 , RIe216f48_4551);
and \g447151/U$3 ( \22400 , RIe219c48_4583, \18032 );
nor \g447151/U$1 ( \22401 , \22399 , \22400 );
and \g446395/U$2 ( \22402 , RIf16b470_5680, \16354 );
and \g446395/U$3 ( \22403 , RIe21f648_4647, \16485 );
and \g449387/U$2 ( \22404 , RIe225048_4711, \16321 );
and \g449387/U$3 ( \22405 , \16328 , RIf16d090_5700);
and \g449387/U$4 ( \22406 , RIe214248_4519, \16427 );
nor \g449387/U$1 ( \22407 , \22404 , \22405 , \22406 );
and \g453663/U$2 ( \22408 , \16361 , RIe208e48_4391);
and \g453663/U$3 ( \22409 , RIe20bb48_4423, \16364 );
nor \g453663/U$1 ( \22410 , \22408 , \22409 );
and \g453662/U$2 ( \22411 , \16377 , RIe222348_4679);
and \g453662/U$3 ( \22412 , RIf16c550_5692, \16313 );
nor \g453662/U$1 ( \22413 , \22411 , \22412 );
and \g455356/U$2 ( \22414 , \16317 , RIe20e848_4455);
and \g455356/U$3 ( \22415 , RIf1684a0_5646, \16325 );
nor \g455356/U$1 ( \22416 , \22414 , \22415 );
not \g455355/U$1 ( \22417 , \22416 );
and \g450408/U$2 ( \22418 , \22417 , \16336 );
and \g450408/U$3 ( \22419 , RIf16a4f8_5669, \16448 );
nor \g450408/U$1 ( \22420 , \22418 , \22419 );
nand \g448117/U$1 ( \22421 , \22407 , \22410 , \22413 , \22420 );
nor \g446395/U$1 ( \22422 , \22402 , \22403 , \22421 );
not \g444821/U$3 ( \22423 , \22422 );
not \g444821/U$4 ( \22424 , \16389 );
and \g444821/U$2 ( \22425 , \22423 , \22424 );
and \g446396/U$2 ( \22426 , RIfe9c6f0_8124, \16313 );
and \g446396/U$3 ( \22427 , RIfc9c848_6803, \16361 );
and \g449389/U$2 ( \22428 , RIf15f0f8_5541, \16427 );
and \g449389/U$3 ( \22429 , \16448 , RIf160fe8_5563);
and \g449389/U$4 ( \22430 , RIf166448_5623, \16321 );
nor \g449389/U$1 ( \22431 , \22428 , \22429 , \22430 );
and \g453669/U$2 ( \22432 , \16368 , RIfe9c588_8123);
and \g453669/U$3 ( \22433 , RIfe9bfe8_8119, \16371 );
nor \g453669/U$1 ( \22434 , \22432 , \22433 );
and \g455104/U$2 ( \22435 , \16317 , RIfcc4550_7256);
and \g455104/U$3 ( \22436 , RIf1654d0_5612, \16325 );
nor \g455104/U$1 ( \22437 , \22435 , \22436 );
not \g450410/U$3 ( \22438 , \22437 );
not \g450410/U$4 ( \22439 , \16330 );
and \g450410/U$2 ( \22440 , \22438 , \22439 );
and \g450410/U$5 ( \22441 , \16328 , RIf1673c0_5634);
nor \g450410/U$1 ( \22442 , \22440 , \22441 );
and \g453668/U$2 ( \22443 , \16334 , RIf162500_5578);
and \g453668/U$3 ( \22444 , RIf1635e0_5590, \16380 );
nor \g453668/U$1 ( \22445 , \22443 , \22444 );
nand \g447939/U$1 ( \22446 , \22431 , \22434 , \22442 , \22445 );
nor \g446396/U$1 ( \22447 , \22426 , \22427 , \22446 );
and \g453666/U$2 ( \22448 , \16364 , RIfc4d540_5902);
and \g453666/U$3 ( \22449 , RIf15d208_5519, \16341 );
nor \g453666/U$1 ( \22450 , \22448 , \22449 );
and \g453665/U$2 ( \22451 , \16398 , RIf15bfc0_5506);
and \g453665/U$3 ( \22452 , RIfe9c150_8120, \16377 );
nor \g453665/U$1 ( \22453 , \22451 , \22452 );
and \g445428/U$2 ( \22454 , \22447 , \22450 , \22453 );
nor \g445428/U$1 ( \22455 , \22454 , \16393 );
nor \g444821/U$1 ( \22456 , \22425 , \22455 );
nor \g448337/U$1 ( \22457 , \16389 , \16437 );
and \g447149/U$2 ( \22458 , \22457 , RIe211548_4487);
nor \g448336/U$1 ( \22459 , \16389 , \16440 );
and \g447149/U$3 ( \22460 , RIf169df0_5664, \22459 );
nor \g447149/U$1 ( \22461 , \22458 , \22460 );
nand \g444436/U$1 ( \22462 , \22401 , \22456 , \22461 );
and \g446391/U$2 ( \22463 , RIe1e73b0_4008, \16313 );
and \g446391/U$3 ( \22464 , RIe1bfdb0_3560, \16361 );
and \g449383/U$2 ( \22465 , RIe1ea0b0_4040, \16319 );
and \g449383/U$3 ( \22466 , \16485 , RIe1decb0_3912);
and \g449383/U$4 ( \22467 , RIe1e19b0_3944, \16354 );
nor \g449383/U$1 ( \22468 , \22465 , \22466 , \22467 );
and \g453547/U$2 ( \22469 , \16368 , RIe1cb1b0_3688);
and \g453547/U$3 ( \22470 , RIe1cdeb0_3720, \16371 );
nor \g453547/U$1 ( \22471 , \22469 , \22470 );
and \g455193/U$2 ( \22472 , \16317 , RIe1d0bb0_3752);
and \g455193/U$3 ( \22473 , RIe1d38b0_3784, \16325 );
nor \g455193/U$1 ( \22474 , \22472 , \22473 );
not \g450402/U$3 ( \22475 , \22474 );
not \g450402/U$4 ( \22476 , \16351 );
and \g450402/U$2 ( \22477 , \22475 , \22476 );
and \g450402/U$5 ( \22478 , \16328 , RIe1ecdb0_4072);
nor \g450402/U$1 ( \22479 , \22477 , \22478 );
and \g453648/U$2 ( \22480 , \16334 , RIe1d92b0_3848);
and \g453648/U$3 ( \22481 , RIe1dbfb0_3880, \16380 );
nor \g453648/U$1 ( \22482 , \22480 , \22481 );
nand \g447937/U$1 ( \22483 , \22468 , \22471 , \22479 , \22482 );
nor \g446391/U$1 ( \22484 , \22463 , \22464 , \22483 );
and \g453644/U$2 ( \22485 , \16364 , RIe1c2ab0_3592);
and \g453644/U$3 ( \22486 , RIe1c84b0_3656, \16341 );
nor \g453644/U$1 ( \22487 , \22485 , \22486 );
and \g453643/U$2 ( \22488 , \16398 , RIe1c57b0_3624);
and \g453643/U$3 ( \22489 , RIe1e46b0_3976, \16377 );
nor \g453643/U$1 ( \22490 , \22488 , \22489 );
and \g445425/U$2 ( \22491 , \22484 , \22487 , \22490 );
nor \g445425/U$1 ( \22492 , \22491 , \16555 );
and \g446393/U$2 ( \22493 , RIe1a46f0_3248, \16313 );
and \g446393/U$3 ( \22494 , RIe172560_2678, \16361 );
and \g449385/U$2 ( \22495 , RIe2001a8_4291, \16427 );
and \g449385/U$3 ( \22496 , \16432 , RIe206148_4359);
and \g449385/U$4 ( \22497 , RIe1a73f0_3280, \16321 );
nor \g449385/U$1 ( \22498 , \22495 , \22496 , \22497 );
and \g453659/U$2 ( \22499 , \16368 , RIe1f20a8_4131);
and \g453659/U$3 ( \22500 , RIe1f9560_4214, \16371 );
nor \g453659/U$1 ( \22501 , \22499 , \22500 );
and \g455314/U$2 ( \22502 , \16317 , RIe17a3f0_2768);
and \g455314/U$3 ( \22503 , RIe18def0_2992, \16325 );
nor \g455314/U$1 ( \22504 , \22502 , \22503 );
not \g450404/U$3 ( \22505 , \22504 );
not \g450404/U$4 ( \22506 , \16330 );
and \g450404/U$2 ( \22507 , \22505 , \22506 );
and \g450404/U$5 ( \22508 , \16328 , RIe1aa0f0_3312);
nor \g450404/U$1 ( \22509 , \22507 , \22508 );
and \g453657/U$2 ( \22510 , \16334 , RIe21c948_4615);
and \g453657/U$3 ( \22511 , RIe227d48_4743, \16380 );
nor \g453657/U$1 ( \22512 , \22510 , \22511 );
nand \g447938/U$1 ( \22513 , \22498 , \22501 , \22509 , \22512 );
nor \g446393/U$1 ( \22514 , \22493 , \22494 , \22513 );
and \g453655/U$2 ( \22515 , \16364 , RIe1aff28_3379);
and \g453655/U$3 ( \22516 , RIe1d65b0_3816, \16341 );
nor \g453655/U$1 ( \22517 , \22515 , \22516 );
and \g453653/U$2 ( \22518 , \16398 , RIe1bd0b0_3528);
and \g453653/U$3 ( \22519 , RIe1a19f0_3216, \16377 );
nor \g453653/U$1 ( \22520 , \22518 , \22519 );
and \g445427/U$2 ( \22521 , \22514 , \22517 , \22520 );
nor \g445427/U$1 ( \22522 , \22521 , \16586 );
or \g444301/U$1 ( \22523 , \22398 , \22462 , \22492 , \22522 );
and \g446387/U$2 ( \22524 , RIf145a90_5252, \16313 );
and \g446387/U$3 ( \22525 , RIe17d0f0_2800, \16361 );
and \g449379/U$2 ( \22526 , RIe1884f0_2928, \16427 );
and \g449379/U$3 ( \22527 , \16432 , RIe18b1f0_2960);
and \g449379/U$4 ( \22528 , RIe19bff0_3152, \16319 );
nor \g449379/U$1 ( \22529 , \22526 , \22527 , \22528 );
and \g453629/U$2 ( \22530 , \16368 , RIe1857f0_2896);
and \g453629/U$3 ( \22531 , RIfc72980_6326, \16371 );
nor \g453629/U$1 ( \22532 , \22530 , \22531 );
and \g455351/U$2 ( \22533 , \16317 , RIe1965f0_3088);
and \g455351/U$3 ( \22534 , RIf144de8_5243, \16325 );
nor \g455351/U$1 ( \22535 , \22533 , \22534 );
not \g450398/U$3 ( \22536 , \22535 );
not \g450398/U$4 ( \22537 , \16330 );
and \g450398/U$2 ( \22538 , \22536 , \22537 );
and \g450398/U$5 ( \22539 , \16326 , RIe19ecf0_3184);
nor \g450398/U$1 ( \22540 , \22538 , \22539 );
and \g453628/U$2 ( \22541 , \16334 , RIe190bf0_3024);
and \g453628/U$3 ( \22542 , RIe1938f0_3056, \16380 );
nor \g453628/U$1 ( \22543 , \22541 , \22542 );
nand \g447933/U$1 ( \22544 , \22529 , \22532 , \22540 , \22543 );
nor \g446387/U$1 ( \22545 , \22524 , \22525 , \22544 );
and \g453626/U$2 ( \22546 , \16364 , RIe17fdf0_2832);
and \g453626/U$3 ( \22547 , RIf143060_5222, \16339 );
nor \g453626/U$1 ( \22548 , \22546 , \22547 );
and \g453625/U$2 ( \22549 , \16337 , RIe182af0_2864);
and \g453625/U$3 ( \22550 , RIe1992f0_3120, \16377 );
nor \g453625/U$1 ( \22551 , \22549 , \22550 );
and \g445423/U$2 ( \22552 , \22545 , \22548 , \22551 );
nor \g445423/U$1 ( \22553 , \22552 , \16618 );
and \g446389/U$2 ( \22554 , RIe177858_2737, \16313 );
and \g446389/U$3 ( \22555 , RIfced608_7723, \16361 );
and \g449382/U$2 ( \22556 , RIf141710_5204, \16321 );
and \g449382/U$3 ( \22557 , \16485 , RIfca54e8_6903);
and \g449382/U$4 ( \22558 , RIfcea638_7689, \16356 );
nor \g449382/U$1 ( \22559 , \22556 , \22557 , \22558 );
and \g453639/U$2 ( \22560 , \16368 , RIe174b58_2705);
and \g453639/U$3 ( \22561 , RIee3a4f8_5122, \16371 );
nor \g453639/U$1 ( \22562 , \22560 , \22561 );
and \g455143/U$2 ( \22563 , \16317 , RIee3b5d8_5134);
and \g455143/U$3 ( \22564 , RIee3c988_5148, \16325 );
nor \g455143/U$1 ( \22565 , \22563 , \22564 );
not \g450401/U$3 ( \22566 , \22565 );
not \g450401/U$4 ( \22567 , \16351 );
and \g450401/U$2 ( \22568 , \22566 , \22567 );
and \g450401/U$5 ( \22569 , \16328 , RIf142688_5215);
nor \g450401/U$1 ( \22570 , \22568 , \22569 );
and \g453638/U$2 ( \22571 , \16334 , RIee3dbd0_5161);
and \g453638/U$3 ( \22572 , RIee3e878_5170, \16380 );
nor \g453638/U$1 ( \22573 , \22571 , \22572 );
nand \g447936/U$1 ( \22574 , \22559 , \22562 , \22570 , \22573 );
nor \g446389/U$1 ( \22575 , \22554 , \22555 , \22574 );
and \g453635/U$2 ( \22576 , \16364 , RIf16e9e0_5718);
and \g453635/U$3 ( \22577 , RIf170600_5738, \16341 );
nor \g453635/U$1 ( \22578 , \22576 , \22577 );
and \g453634/U$2 ( \22579 , \16398 , RIfc76fd0_6376);
and \g453634/U$3 ( \22580 , RIe176778_2725, \16377 );
nor \g453634/U$1 ( \22581 , \22579 , \22580 );
and \g445424/U$2 ( \22582 , \22575 , \22578 , \22581 );
nor \g445424/U$1 ( \22583 , \22582 , \16649 );
or \g444230/U$1 ( \22584 , \22523 , \22553 , \22583 );
_DC \g3fda/U$1 ( \22585 , \22584 , \16652 );
and \g453761/U$2 ( \22586 , \16313 , RIe1a4588_3247);
and \g453761/U$3 ( \22587 , RIe1a7288_3279, \16319 );
nor \g453761/U$1 ( \22588 , \22586 , \22587 );
and \g446416/U$2 ( \22589 , RIe1a9f88_3311, \16328 );
and \g446416/U$3 ( \22590 , RIe21c7e0_4614, \16334 );
and \g449415/U$2 ( \22591 , RIe1bcf48_3527, \16337 );
and \g449415/U$3 ( \22592 , \16341 , RIe1d6448_3815);
and \g449415/U$4 ( \22593 , RIe17a288_2767, \16485 );
nor \g449415/U$1 ( \22594 , \22591 , \22592 , \22593 );
and \g455370/U$2 ( \22595 , \16317 , RIe200040_4290);
and \g455370/U$3 ( \22596 , RIe205fe0_4358, \16325 );
nor \g455370/U$1 ( \22597 , \22595 , \22596 );
not \g450435/U$3 ( \22598 , \22597 );
not \g450435/U$4 ( \22599 , \16351 );
and \g450435/U$2 ( \22600 , \22598 , \22599 );
and \g450435/U$5 ( \22601 , \16354 , RIe18dd88_2991);
nor \g450435/U$1 ( \22602 , \22600 , \22601 );
and \g453768/U$2 ( \22603 , \16361 , RIe1723f8_2677);
and \g453768/U$3 ( \22604 , RIe1afdc0_3378, \16364 );
nor \g453768/U$1 ( \22605 , \22603 , \22604 );
and \g453766/U$2 ( \22606 , \16368 , RIe1f1f40_4130);
and \g453766/U$3 ( \22607 , RIe1f93f8_4213, \16371 );
nor \g453766/U$1 ( \22608 , \22606 , \22607 );
nand \g447957/U$1 ( \22609 , \22594 , \22602 , \22605 , \22608 );
nor \g446416/U$1 ( \22610 , \22589 , \22590 , \22609 );
and \g453763/U$2 ( \22611 , \16377 , RIe1a1888_3215);
and \g453763/U$3 ( \22612 , RIe227be0_4742, \16380 );
nor \g453763/U$1 ( \22613 , \22611 , \22612 );
nand \g445685/U$1 ( \22614 , \22588 , \22610 , \22613 );
and \g444676/U$2 ( \22615 , \22614 , \16752 );
and \g446418/U$2 ( \22616 , RIe1deb48_3911, \16485 );
and \g446418/U$3 ( \22617 , RIe1dbe48_3879, \16380 );
and \g449416/U$2 ( \22618 , RIe1d0a48_3751, \16427 );
and \g449416/U$3 ( \22619 , \16398 , RIe1c5648_3623);
and \g449416/U$4 ( \22620 , RIe1c8348_3655, \16341 );
nor \g449416/U$1 ( \22621 , \22618 , \22619 , \22620 );
and \g453777/U$2 ( \22622 , \16361 , RIe1bfc48_3559);
and \g453777/U$3 ( \22623 , RIe1c2948_3591, \16364 );
nor \g453777/U$1 ( \22624 , \22622 , \22623 );
and \g453776/U$2 ( \22625 , \16377 , RIe1e4548_3975);
and \g453776/U$3 ( \22626 , RIe1e7248_4007, \16313 );
nor \g453776/U$1 ( \22627 , \22625 , \22626 );
and \g455371/U$2 ( \22628 , \16317 , RIe1e9f48_4039);
and \g455371/U$3 ( \22629 , RIe1ecc48_4071, \16325 );
nor \g455371/U$1 ( \22630 , \22628 , \22629 );
not \g450438/U$3 ( \22631 , \22630 );
not \g450438/U$4 ( \22632 , \16311 );
and \g450438/U$2 ( \22633 , \22631 , \22632 );
and \g450438/U$5 ( \22634 , \16448 , RIe1d3748_3783);
nor \g450438/U$1 ( \22635 , \22633 , \22634 );
nand \g447959/U$1 ( \22636 , \22621 , \22624 , \22627 , \22635 );
nor \g446418/U$1 ( \22637 , \22616 , \22617 , \22636 );
and \g453772/U$2 ( \22638 , \16368 , RIe1cb048_3687);
and \g453772/U$3 ( \22639 , RIe1e1848_3943, \16356 );
nor \g453772/U$1 ( \22640 , \22638 , \22639 );
and \g453773/U$2 ( \22641 , \16334 , RIe1d9148_3847);
and \g453773/U$3 ( \22642 , RIe1cdd48_3719, \16371 );
nor \g453773/U$1 ( \22643 , \22641 , \22642 );
and \g445441/U$2 ( \22644 , \22637 , \22640 , \22643 );
nor \g445441/U$1 ( \22645 , \22644 , \16555 );
nor \g444676/U$1 ( \22646 , \22615 , \22645 );
and \g447170/U$2 ( \22647 , \18711 , RIfe9a0f8_8097);
and \g447170/U$3 ( \22648 , RIfe9a260_8098, \18713 );
nor \g447170/U$1 ( \22649 , \22647 , \22648 );
not \g444414/U$2 ( \22650 , \22649 );
and \g453824/U$2 ( \22651 , \16313 , RIf16c3e8_5691);
and \g453824/U$3 ( \22652 , RIe224ee0_4710, \16321 );
nor \g453824/U$1 ( \22653 , \22651 , \22652 );
and \g446429/U$2 ( \22654 , RIfe9aad0_8104, \16328 );
and \g446429/U$3 ( \22655 , RIe216de0_4550, \16334 );
and \g449431/U$2 ( \22656 , RIe20e6e0_4454, \16398 );
and \g449431/U$3 ( \22657 , \16341 , RIf168338_5645);
and \g449431/U$4 ( \22658 , RIe21f4e0_4646, \16344 );
nor \g449431/U$1 ( \22659 , \22656 , \22657 , \22658 );
and \g454505/U$2 ( \22660 , \16317 , RIe2140e0_4518);
and \g454505/U$3 ( \22661 , RIfc880a0_6570, \16325 );
nor \g454505/U$1 ( \22662 , \22660 , \22661 );
not \g450452/U$3 ( \22663 , \22662 );
not \g450452/U$4 ( \22664 , \16351 );
and \g450452/U$2 ( \22665 , \22663 , \22664 );
and \g450452/U$5 ( \22666 , \16356 , RIfcd3898_7429);
nor \g450452/U$1 ( \22667 , \22665 , \22666 );
and \g453828/U$2 ( \22668 , \16361 , RIe208ce0_4390);
and \g453828/U$3 ( \22669 , RIe20b9e0_4422, \16364 );
nor \g453828/U$1 ( \22670 , \22668 , \22669 );
and \g453827/U$2 ( \22671 , \16368 , RIe2113e0_4486);
and \g453827/U$3 ( \22672 , RIf169c88_5663, \16371 );
nor \g453827/U$1 ( \22673 , \22671 , \22672 );
nand \g447964/U$1 ( \22674 , \22659 , \22667 , \22670 , \22673 );
nor \g446429/U$1 ( \22675 , \22654 , \22655 , \22674 );
and \g453825/U$2 ( \22676 , \16377 , RIe2221e0_4678);
and \g453825/U$3 ( \22677 , RIe219ae0_4582, \16380 );
nor \g453825/U$1 ( \22678 , \22676 , \22677 );
nand \g445688/U$1 ( \22679 , \22653 , \22675 , \22678 );
and \g444864/U$2 ( \22680 , \22679 , \16390 );
and \g449429/U$2 ( \22681 , RIf15be58_5505, \16398 );
and \g449429/U$3 ( \22682 , \16339 , RIfca8d28_6943);
and \g449429/U$4 ( \22683 , RIfc85c10_6544, \16485 );
nor \g449429/U$1 ( \22684 , \22681 , \22682 , \22683 );
and \g454483/U$2 ( \22685 , \16317 , RIf15ef90_5540);
and \g454483/U$3 ( \22686 , RIf160e80_5562, \16325 );
nor \g454483/U$1 ( \22687 , \22685 , \22686 );
not \g450450/U$3 ( \22688 , \22687 );
not \g450450/U$4 ( \22689 , \16351 );
and \g450450/U$2 ( \22690 , \22688 , \22689 );
and \g450450/U$5 ( \22691 , \16356 , RIfc500d8_5933);
nor \g450450/U$1 ( \22692 , \22690 , \22691 );
and \g453817/U$2 ( \22693 , \16361 , RIfc6a988_6235);
and \g453817/U$3 ( \22694 , RIfcedba8_7727, \16364 );
nor \g453817/U$1 ( \22695 , \22693 , \22694 );
and \g453816/U$2 ( \22696 , \16368 , RIfe9ac38_8105);
and \g453816/U$3 ( \22697 , RIfe9a968_8103, \16371 );
nor \g453816/U$1 ( \22698 , \22696 , \22697 );
nand \g447963/U$1 ( \22699 , \22684 , \22692 , \22695 , \22698 );
and \g444864/U$3 ( \22700 , \16394 , \22699 );
nor \g444864/U$1 ( \22701 , \22680 , \22700 );
and \g447172/U$2 ( \22702 , \16705 , RIfce9c60_7682);
and \g447172/U$3 ( \22703 , RIfce81a8_7663, \16707 );
nor \g447172/U$1 ( \22704 , \22702 , \22703 );
and \g447171/U$2 ( \22705 , \16710 , RIfc9c6e0_6802);
and \g447171/U$3 ( \22706 , RIfce4c38_7625, \16712 );
nor \g447171/U$1 ( \22707 , \22705 , \22706 );
and \g447173/U$2 ( \22708 , \16715 , RIe201af8_4309);
and \g447173/U$3 ( \22709 , RIe2035b0_4328, \16717 );
nor \g447173/U$1 ( \22710 , \22708 , \22709 );
nand \g444661/U$1 ( \22711 , \22701 , \22704 , \22707 , \22710 );
and \g446425/U$2 ( \22712 , RIfe9a3c8_8099, \16328 );
and \g446425/U$3 ( \22713 , RIfce5340_7630, \16334 );
and \g449423/U$2 ( \22714 , RIfc576f8_6017, \16427 );
and \g449423/U$3 ( \22715 , \16448 , RIfc5cb58_6077);
and \g449423/U$4 ( \22716 , RIf13f820_5182, \16485 );
nor \g449423/U$1 ( \22717 , \22714 , \22715 , \22716 );
and \g455375/U$2 ( \22718 , \16317 , RIfc7c2c8_6435);
and \g455375/U$3 ( \22719 , RIfc7adb0_6420, \16325 );
nor \g455375/U$1 ( \22720 , \22718 , \22719 );
not \g455374/U$1 ( \22721 , \22720 );
and \g450444/U$2 ( \22722 , \22721 , \16336 );
and \g450444/U$3 ( \22723 , RIfcb9150_7128, \16354 );
nor \g450444/U$1 ( \22724 , \22722 , \22723 );
and \g453806/U$2 ( \22725 , \16361 , RIfc7e758_6461);
and \g453806/U$3 ( \22726 , RIfcb2d78_7057, \16364 );
nor \g453806/U$1 ( \22727 , \22725 , \22726 );
and \g453804/U$2 ( \22728 , \16368 , RIe1749f0_2704);
and \g453804/U$3 ( \22729 , RIfc780b0_6388, \16371 );
nor \g453804/U$1 ( \22730 , \22728 , \22729 );
nand \g448121/U$1 ( \22731 , \22717 , \22724 , \22727 , \22730 );
nor \g446425/U$1 ( \22732 , \22712 , \22713 , \22731 );
and \g453801/U$2 ( \22733 , \16380 , RIfc9fc50_6840);
and \g453801/U$3 ( \22734 , RIf1415a8_5203, \16321 );
nor \g453801/U$1 ( \22735 , \22733 , \22734 );
and \g445504/U$2 ( \22736 , \22732 , \22735 );
nor \g445504/U$1 ( \22737 , \22736 , \16649 );
and \g446427/U$2 ( \22738 , RIe18b088_2959, \16448 );
and \g446427/U$3 ( \22739 , RIfe9a800_8102, \16371 );
and \g449426/U$2 ( \22740 , RIe196488_3087, \16485 );
and \g449426/U$3 ( \22741 , \16354 , RIfe9a530_8100);
and \g449426/U$4 ( \22742 , RIe182988_2863, \16398 );
nor \g449426/U$1 ( \22743 , \22740 , \22741 , \22742 );
and \g455084/U$2 ( \22744 , \16317 , RIe19be88_3151);
and \g455084/U$3 ( \22745 , RIe19eb88_3183, \16325 );
nor \g455084/U$1 ( \22746 , \22744 , \22745 );
not \g450448/U$3 ( \22747 , \22746 );
not \g450448/U$4 ( \22748 , \16311 );
and \g450448/U$2 ( \22749 , \22747 , \22748 );
and \g450448/U$5 ( \22750 , \16341 , RIfc8d938_6633);
nor \g450448/U$1 ( \22751 , \22749 , \22750 );
and \g453812/U$2 ( \22752 , \16377 , RIe199188_3119);
and \g453812/U$3 ( \22753 , RIfe9a698_8101, \16313 );
nor \g453812/U$1 ( \22754 , \22752 , \22753 );
and \g453813/U$2 ( \22755 , \16334 , RIe190a88_3023);
and \g453813/U$3 ( \22756 , RIe193788_3055, \16380 );
nor \g453813/U$1 ( \22757 , \22755 , \22756 );
nand \g447428/U$1 ( \22758 , \22743 , \22751 , \22754 , \22757 );
nor \g446427/U$1 ( \22759 , \22738 , \22739 , \22758 );
and \g453808/U$2 ( \22760 , \16364 , RIe17fc88_2831);
and \g453808/U$3 ( \22761 , RIe185688_2895, \16368 );
nor \g453808/U$1 ( \22762 , \22760 , \22761 );
and \g453809/U$2 ( \22763 , \16361 , RIe17cf88_2799);
and \g453809/U$3 ( \22764 , RIe188388_2927, \16427 );
nor \g453809/U$1 ( \22765 , \22763 , \22764 );
and \g445448/U$2 ( \22766 , \22759 , \22762 , \22765 );
nor \g445448/U$1 ( \22767 , \22766 , \16618 );
nor \g444414/U$1 ( \22768 , \22650 , \22711 , \22737 , \22767 );
and \g453791/U$2 ( \22769 , \16364 , RIe1ad390_3348);
and \g453791/U$3 ( \22770 , RIe1b3498_3417, \16371 );
nor \g453791/U$1 ( \22771 , \22769 , \22770 );
and \g446422/U$2 ( \22772 , RIfc55970_5996, \16427 );
and \g446422/U$3 ( \22773 , RIe1b1cb0_3400, \16368 );
and \g449421/U$2 ( \22774 , RIfcc2228_7231, \16485 );
and \g449421/U$3 ( \22775 , \16356 , RIfc598b8_6041);
and \g449421/U$4 ( \22776 , RIfc4b4e8_5879, \16398 );
nor \g449421/U$1 ( \22777 , \22774 , \22775 , \22776 );
and \g455089/U$2 ( \22778 , \16317 , RIfca7ae0_6930);
and \g455089/U$3 ( \22779 , RIfcc70e8_7287, \16325 );
nor \g455089/U$1 ( \22780 , \22778 , \22779 );
not \g450442/U$3 ( \22781 , \22780 );
not \g450442/U$4 ( \22782 , \16311 );
and \g450442/U$2 ( \22783 , \22781 , \22782 );
and \g450442/U$5 ( \22784 , \16341 , RIfcb7698_7109);
nor \g450442/U$1 ( \22785 , \22783 , \22784 );
and \g453795/U$2 ( \22786 , \16377 , RIe1b8358_3473);
and \g453795/U$3 ( \22787 , RIe1ba518_3497, \16313 );
nor \g453795/U$1 ( \22788 , \22786 , \22787 );
and \g453796/U$2 ( \22789 , \16334 , RIe1b4848_3431);
and \g453796/U$3 ( \22790 , RIe1b6198_3449, \16380 );
nor \g453796/U$1 ( \22791 , \22789 , \22790 );
nand \g447427/U$1 ( \22792 , \22777 , \22785 , \22788 , \22791 );
nor \g446422/U$1 ( \22793 , \22772 , \22773 , \22792 );
and \g453792/U$2 ( \22794 , \16361 , RIe1abba8_3331);
and \g453792/U$3 ( \22795 , RIfc82f10_6512, \16448 );
nor \g453792/U$1 ( \22796 , \22794 , \22795 );
nand \g445687/U$1 ( \22797 , \22771 , \22793 , \22796 );
and \g444677/U$2 ( \22798 , \22797 , \16477 );
and \g446419/U$2 ( \22799 , RIfcaee30_7012, \16427 );
and \g446419/U$3 ( \22800 , RIe1f4538_4157, \16368 );
and \g449419/U$2 ( \22801 , RIfccb198_7333, \16319 );
and \g449419/U$3 ( \22802 , \16328 , RIfc71cd8_6317);
and \g449419/U$4 ( \22803 , RIfcaecc8_7011, \16398 );
nor \g449419/U$1 ( \22804 , \22801 , \22802 , \22803 );
and \g455097/U$2 ( \22805 , \16317 , RIfc6d688_6267);
and \g455097/U$3 ( \22806 , RIfc4c730_5892, \16325 );
nor \g455097/U$1 ( \22807 , \22805 , \22806 );
not \g450440/U$3 ( \22808 , \22807 );
not \g450440/U$4 ( \22809 , \16330 );
and \g450440/U$2 ( \22810 , \22808 , \22809 );
and \g450440/U$5 ( \22811 , \16341 , RIfc63ea8_6159);
nor \g450440/U$1 ( \22812 , \22810 , \22811 );
and \g453784/U$2 ( \22813 , \16377 , RIfec3b88_8347);
and \g453784/U$3 ( \22814 , RIfcaa3a8_6959, \16313 );
nor \g453784/U$1 ( \22815 , \22813 , \22814 );
and \g453786/U$2 ( \22816 , \16334 , RIe1f6860_4182);
and \g453786/U$3 ( \22817 , RIfca8e90_6944, \16380 );
nor \g453786/U$1 ( \22818 , \22816 , \22817 );
nand \g447426/U$1 ( \22819 , \22804 , \22812 , \22815 , \22818 );
nor \g446419/U$1 ( \22820 , \22799 , \22800 , \22819 );
and \g453783/U$2 ( \22821 , \16361 , RIfeab1c8_8263);
and \g453783/U$3 ( \22822 , RIfc64e20_6170, \16448 );
nor \g453783/U$1 ( \22823 , \22821 , \22822 );
and \g453782/U$2 ( \22824 , \16364 , RIfcae458_7005);
and \g453782/U$3 ( \22825 , RIfccee10_7376, \16371 );
nor \g453782/U$1 ( \22826 , \22824 , \22825 );
and \g445443/U$2 ( \22827 , \22820 , \22823 , \22826 );
nor \g445443/U$1 ( \22828 , \22827 , \16480 );
nor \g444677/U$1 ( \22829 , \22798 , \22828 );
nand \g444287/U$1 ( \22830 , \22646 , \22768 , \22829 );
_DC \g405f/U$1 ( \22831 , \22830 , \16652 );
and \g453225/U$2 ( \22832 , \16364 , RIe1afc58_3377);
and \g453225/U$3 ( \22833 , RIe1f9290_4212, \16371 );
nor \g453225/U$1 ( \22834 , \22832 , \22833 );
and \g446301/U$2 ( \22835 , RIe1ffed8_4289, \16427 );
and \g446301/U$3 ( \22836 , RIe1f1dd8_4129, \16368 );
and \g449269/U$2 ( \22837 , RIe17a120_2766, \16485 );
and \g449269/U$3 ( \22838 , \16356 , RIe18dc20_2990);
and \g449269/U$4 ( \22839 , RIe1bcde0_3526, \16398 );
nor \g449269/U$1 ( \22840 , \22837 , \22838 , \22839 );
and \g454553/U$2 ( \22841 , \16317 , RIe1a7120_3278);
and \g454553/U$3 ( \22842 , RIe1a9e20_3310, \16325 );
nor \g454553/U$1 ( \22843 , \22841 , \22842 );
not \g450286/U$3 ( \22844 , \22843 );
not \g450286/U$4 ( \22845 , \16311 );
and \g450286/U$2 ( \22846 , \22844 , \22845 );
and \g450286/U$5 ( \22847 , \16341 , RIe1d62e0_3814);
nor \g450286/U$1 ( \22848 , \22846 , \22847 );
and \g453229/U$2 ( \22849 , \16377 , RIe1a1720_3214);
and \g453229/U$3 ( \22850 , RIe1a4420_3246, \16313 );
nor \g453229/U$1 ( \22851 , \22849 , \22850 );
and \g453232/U$2 ( \22852 , \16334 , RIe21c678_4613);
and \g453232/U$3 ( \22853 , RIe227a78_4741, \16380 );
nor \g453232/U$1 ( \22854 , \22852 , \22853 );
nand \g447405/U$1 ( \22855 , \22840 , \22848 , \22851 , \22854 );
nor \g446301/U$1 ( \22856 , \22835 , \22836 , \22855 );
and \g453226/U$2 ( \22857 , \16361 , RIe172290_2676);
and \g453226/U$3 ( \22858 , RIe205e78_4357, \16448 );
nor \g453226/U$1 ( \22859 , \22857 , \22858 );
nand \g445652/U$1 ( \22860 , \22834 , \22856 , \22859 );
and \g444795/U$2 ( \22861 , \22860 , \16752 );
and \g449267/U$2 ( \22862 , RIe1e9de0_4038, \16321 );
and \g449267/U$3 ( \22863 , \16328 , RIe1ecae0_4070);
and \g449267/U$4 ( \22864 , RIe1c54e0_3622, \16398 );
nor \g449267/U$1 ( \22865 , \22862 , \22863 , \22864 );
and \g455294/U$2 ( \22866 , \16317 , RIe1de9e0_3910);
and \g455294/U$3 ( \22867 , RIe1e16e0_3942, \16325 );
nor \g455294/U$1 ( \22868 , \22866 , \22867 );
not \g450285/U$3 ( \22869 , \22868 );
not \g450285/U$4 ( \22870 , \16330 );
and \g450285/U$2 ( \22871 , \22869 , \22870 );
and \g450285/U$5 ( \22872 , \16341 , RIe1c81e0_3654);
nor \g450285/U$1 ( \22873 , \22871 , \22872 );
and \g453220/U$2 ( \22874 , \16377 , RIe1e43e0_3974);
and \g453220/U$3 ( \22875 , RIe1e70e0_4006, \16313 );
nor \g453220/U$1 ( \22876 , \22874 , \22875 );
and \g453221/U$2 ( \22877 , \16334 , RIe1d8fe0_3846);
and \g453221/U$3 ( \22878 , RIe1dbce0_3878, \16380 );
nor \g453221/U$1 ( \22879 , \22877 , \22878 );
nand \g447404/U$1 ( \22880 , \22865 , \22873 , \22876 , \22879 );
and \g444795/U$3 ( \22881 , \16750 , \22880 );
nor \g444795/U$1 ( \22882 , \22861 , \22881 );
and \g447075/U$2 ( \22883 , \19208 , RIe1bfae0_3558);
and \g447075/U$3 ( \22884 , RIe1cdbe0_3718, \19210 );
nor \g447075/U$1 ( \22885 , \22883 , \22884 );
and \g447074/U$2 ( \22886 , \19213 , RIe1c27e0_3590);
and \g447074/U$3 ( \22887 , RIe1caee0_3686, \19215 );
nor \g447074/U$1 ( \22888 , \22886 , \22887 );
and \g447073/U$2 ( \22889 , \19218 , RIe1d08e0_3750);
and \g447073/U$3 ( \22890 , RIe1d35e0_3782, \19220 );
nor \g447073/U$1 ( \22891 , \22889 , \22890 );
nand \g444646/U$1 ( \22892 , \22882 , \22885 , \22888 , \22891 );
and \g453210/U$2 ( \22893 , \16364 , RIfcd4540_7438);
and \g453210/U$3 ( \22894 , RIfe98be0_8082, \16371 );
nor \g453210/U$1 ( \22895 , \22893 , \22894 );
and \g446299/U$2 ( \22896 , RIf15ee28_5539, \16427 );
and \g446299/U$3 ( \22897 , RIfe98eb0_8084, \16368 );
and \g449265/U$2 ( \22898 , RIfc61478_6129, \16319 );
and \g449265/U$3 ( \22899 , \16326 , RIfcd4ae0_7442);
and \g449265/U$4 ( \22900 , RIf15bcf0_5504, \16398 );
nor \g449265/U$1 ( \22901 , \22898 , \22899 , \22900 );
and \g454590/U$2 ( \22902 , \16317 , RIfc70928_6303);
and \g454590/U$3 ( \22903 , RIfc70ec8_6307, \16325 );
nor \g454590/U$1 ( \22904 , \22902 , \22903 );
not \g450281/U$3 ( \22905 , \22904 );
not \g450281/U$4 ( \22906 , \16330 );
and \g450281/U$2 ( \22907 , \22905 , \22906 );
and \g450281/U$5 ( \22908 , \16341 , RIf15d0a0_5518);
nor \g450281/U$1 ( \22909 , \22907 , \22908 );
and \g453213/U$2 ( \22910 , \16377 , RIe201990_4308);
and \g453213/U$3 ( \22911 , RIfeab060_8262, \16313 );
nor \g453213/U$1 ( \22912 , \22910 , \22911 );
and \g453214/U$2 ( \22913 , \16334 , RIfcbe880_7190);
and \g453214/U$3 ( \22914 , RIfcec528_7711, \16380 );
nor \g453214/U$1 ( \22915 , \22913 , \22914 );
nand \g447403/U$1 ( \22916 , \22901 , \22909 , \22912 , \22915 );
nor \g446299/U$1 ( \22917 , \22896 , \22897 , \22916 );
and \g453211/U$2 ( \22918 , \16361 , RIf159e00_5482);
and \g453211/U$3 ( \22919 , RIf160d18_5561, \16448 );
nor \g453211/U$1 ( \22920 , \22918 , \22919 );
nand \g445651/U$1 ( \22921 , \22895 , \22917 , \22920 );
and \g444794/U$2 ( \22922 , \22921 , \16394 );
and \g449264/U$2 ( \22923 , RIe20e578_4453, \16337 );
and \g449264/U$3 ( \22924 , \16341 , RIf1681d0_5644);
and \g449264/U$4 ( \22925 , RIe21f378_4645, \16485 );
nor \g449264/U$1 ( \22926 , \22923 , \22924 , \22925 );
and \g455288/U$2 ( \22927 , \16317 , RIe213f78_4517);
and \g455288/U$3 ( \22928 , RIf16a390_5668, \16325 );
nor \g455288/U$1 ( \22929 , \22927 , \22928 );
not \g450280/U$3 ( \22930 , \22929 );
not \g450280/U$4 ( \22931 , \16351 );
and \g450280/U$2 ( \22932 , \22930 , \22931 );
and \g450280/U$5 ( \22933 , \16356 , RIf16b308_5679);
nor \g450280/U$1 ( \22934 , \22932 , \22933 );
and \g453208/U$2 ( \22935 , \16361 , RIe208b78_4389);
and \g453208/U$3 ( \22936 , RIe20b878_4421, \16364 );
nor \g453208/U$1 ( \22937 , \22935 , \22936 );
and \g453207/U$2 ( \22938 , \16368 , RIe211278_4485);
and \g453207/U$3 ( \22939 , RIf169b20_5662, \16371 );
nor \g453207/U$1 ( \22940 , \22938 , \22939 );
nand \g447864/U$1 ( \22941 , \22926 , \22934 , \22937 , \22940 );
and \g444794/U$3 ( \22942 , \16390 , \22941 );
nor \g444794/U$1 ( \22943 , \22922 , \22942 );
and \g447064/U$2 ( \22944 , \18020 , RIe224d78_4709);
and \g447064/U$3 ( \22945 , RIfe98d48_8083, \18022 );
nor \g447064/U$1 ( \22946 , \22944 , \22945 );
and \g447065/U$2 ( \22947 , \18025 , RIe222078_4677);
and \g447065/U$3 ( \22948 , RIf16c280_5690, \18027 );
nor \g447065/U$1 ( \22949 , \22947 , \22948 );
and \g447066/U$2 ( \22950 , \18030 , RIe216c78_4549);
and \g447066/U$3 ( \22951 , RIe219978_4581, \18032 );
nor \g447066/U$1 ( \22952 , \22950 , \22951 );
nand \g444525/U$1 ( \22953 , \22943 , \22946 , \22949 , \22952 );
and \g446294/U$2 ( \22954 , RIf141440_5202, \16321 );
and \g446294/U$3 ( \22955 , RIe1776f0_2736, \16313 );
and \g449259/U$2 ( \22956 , RIfc68660_6210, \16398 );
and \g449259/U$3 ( \22957 , \16339 , RIf170498_5737);
and \g449259/U$4 ( \22958 , RIfc62dc8_6147, \16485 );
nor \g449259/U$1 ( \22959 , \22956 , \22957 , \22958 );
and \g454644/U$2 ( \22960 , \16317 , RIee3b470_5133);
and \g454644/U$3 ( \22961 , RIee3c820_5147, \16325 );
nor \g454644/U$1 ( \22962 , \22960 , \22961 );
not \g450275/U$3 ( \22963 , \22962 );
not \g450275/U$4 ( \22964 , \16351 );
and \g450275/U$2 ( \22965 , \22963 , \22964 );
and \g450275/U$5 ( \22966 , \16354 , RIfcc5bd0_7272);
nor \g450275/U$1 ( \22967 , \22965 , \22966 );
and \g453193/U$2 ( \22968 , \16361 , RIfc6ea38_6281);
and \g453193/U$3 ( \22969 , RIf16e878_5717, \16364 );
nor \g453193/U$1 ( \22970 , \22968 , \22969 );
and \g453192/U$2 ( \22971 , \16368 , RIe174888_2703);
and \g453192/U$3 ( \22972 , RIee3a390_5121, \16371 );
nor \g453192/U$1 ( \22973 , \22971 , \22972 );
nand \g447862/U$1 ( \22974 , \22959 , \22967 , \22970 , \22973 );
nor \g446294/U$1 ( \22975 , \22954 , \22955 , \22974 );
and \g453189/U$2 ( \22976 , \16377 , RIfeab8d0_8268);
and \g453189/U$3 ( \22977 , RIee3e710_5169, \16380 );
nor \g453189/U$1 ( \22978 , \22976 , \22977 );
and \g453187/U$2 ( \22979 , \16334 , RIfc9cb18_6805);
and \g453187/U$3 ( \22980 , RIf142520_5214, \16328 );
nor \g453187/U$1 ( \22981 , \22979 , \22980 );
and \g445361/U$2 ( \22982 , \22975 , \22978 , \22981 );
nor \g445361/U$1 ( \22983 , \22982 , \16649 );
and \g446297/U$2 ( \22984 , RIe188220_2926, \16427 );
and \g446297/U$3 ( \22985 , RIe185520_2894, \16368 );
and \g449261/U$2 ( \22986 , RIe196320_3086, \16485 );
and \g449261/U$3 ( \22987 , \16356 , RIfe98910_8080);
and \g449261/U$4 ( \22988 , RIe182820_2862, \16398 );
nor \g449261/U$1 ( \22989 , \22986 , \22987 , \22988 );
and \g455291/U$2 ( \22990 , \16317 , RIe19bd20_3150);
and \g455291/U$3 ( \22991 , RIe19ea20_3182, \16325 );
nor \g455291/U$1 ( \22992 , \22990 , \22991 );
not \g450277/U$3 ( \22993 , \22992 );
not \g450277/U$4 ( \22994 , \16311 );
and \g450277/U$2 ( \22995 , \22993 , \22994 );
and \g450277/U$5 ( \22996 , \16339 , RIfc95c00_6726);
nor \g450277/U$1 ( \22997 , \22995 , \22996 );
and \g453202/U$2 ( \22998 , \16377 , RIe199020_3118);
and \g453202/U$3 ( \22999 , RIf145928_5251, \16313 );
nor \g453202/U$1 ( \23000 , \22998 , \22999 );
and \g453203/U$2 ( \23001 , \16334 , RIe190920_3022);
and \g453203/U$3 ( \23002 , RIe193620_3054, \16380 );
nor \g453203/U$1 ( \23003 , \23001 , \23002 );
nand \g447402/U$1 ( \23004 , \22989 , \22997 , \23000 , \23003 );
nor \g446297/U$1 ( \23005 , \22984 , \22985 , \23004 );
and \g453199/U$2 ( \23006 , \16361 , RIe17ce20_2798);
and \g453199/U$3 ( \23007 , RIe18af20_2958, \16448 );
nor \g453199/U$1 ( \23008 , \23006 , \23007 );
and \g453197/U$2 ( \23009 , \16364 , RIe17fb20_2830);
and \g453197/U$3 ( \23010 , RIf143e70_5232, \16371 );
nor \g453197/U$1 ( \23011 , \23009 , \23010 );
and \g445363/U$2 ( \23012 , \23005 , \23008 , \23011 );
nor \g445363/U$1 ( \23013 , \23012 , \16618 );
or \g444406/U$1 ( \23014 , \22892 , \22953 , \22983 , \23013 );
and \g446291/U$2 ( \23015 , RIfcec7f8_7713, \16427 );
and \g446291/U$3 ( \23016 , RIe1b1b48_3399, \16368 );
and \g449255/U$2 ( \23017 , RIf14bd00_5322, \16321 );
and \g449255/U$3 ( \23018 , \16328 , RIfc44b70_5804);
and \g449255/U$4 ( \23019 , RIfcda918_7509, \16398 );
nor \g449255/U$1 ( \23020 , \23017 , \23018 , \23019 );
and \g455274/U$2 ( \23021 , \16317 , RIf149f78_5301);
and \g455274/U$3 ( \23022 , RIf14a950_5308, \16325 );
nor \g455274/U$1 ( \23023 , \23021 , \23022 );
not \g450271/U$3 ( \23024 , \23023 );
not \g450271/U$4 ( \23025 , \16330 );
and \g450271/U$2 ( \23026 , \23024 , \23025 );
and \g450271/U$5 ( \23027 , \16339 , RIfc4b650_5880);
nor \g450271/U$1 ( \23028 , \23026 , \23027 );
and \g453169/U$2 ( \23029 , \16377 , RIfe987a8_8079);
and \g453169/U$3 ( \23030 , RIfe992e8_8087, \16313 );
nor \g453169/U$1 ( \23031 , \23029 , \23030 );
and \g453171/U$2 ( \23032 , \16334 , RIfe98640_8078);
and \g453171/U$3 ( \23033 , RIfe99180_8086, \16380 );
nor \g453171/U$1 ( \23034 , \23032 , \23033 );
nand \g447400/U$1 ( \23035 , \23020 , \23028 , \23031 , \23034 );
nor \g446291/U$1 ( \23036 , \23015 , \23016 , \23035 );
and \g453168/U$2 ( \23037 , \16361 , RIfe99018_8085);
and \g453168/U$3 ( \23038 , RIf149438_5293, \16432 );
nor \g453168/U$1 ( \23039 , \23037 , \23038 );
and \g453167/U$2 ( \23040 , \16364 , RIfe98370_8076);
and \g453167/U$3 ( \23041 , RIfe984d8_8077, \16371 );
nor \g453167/U$1 ( \23042 , \23040 , \23041 );
and \g445357/U$2 ( \23043 , \23036 , \23039 , \23042 );
nor \g445357/U$1 ( \23044 , \23043 , \16909 );
and \g446293/U$2 ( \23045 , RIf1520d8_5393, \16427 );
and \g446293/U$3 ( \23046 , RIe1f43d0_4156, \16368 );
and \g449257/U$2 ( \23047 , RIf155be8_5435, \16485 );
and \g449257/U$3 ( \23048 , \16356 , RIf156728_5443);
and \g449257/U$4 ( \23049 , RIfcd2380_7414, \16398 );
nor \g449257/U$1 ( \23050 , \23047 , \23048 , \23049 );
and \g454652/U$2 ( \23051 , \16317 , RIf158078_5461);
and \g454652/U$3 ( \23052 , RIf1592c0_5474, \16325 );
nor \g454652/U$1 ( \23053 , \23051 , \23052 );
not \g450273/U$3 ( \23054 , \23053 );
not \g450273/U$4 ( \23055 , \16311 );
and \g450273/U$2 ( \23056 , \23054 , \23055 );
and \g450273/U$5 ( \23057 , \16341 , RIf14fdb0_5368);
nor \g450273/U$1 ( \23058 , \23056 , \23057 );
and \g453181/U$2 ( \23059 , \16377 , RIfea7988_8223);
and \g453181/U$3 ( \23060 , RIfca3a30_6884, \16313 );
nor \g453181/U$1 ( \23061 , \23059 , \23060 );
and \g453183/U$2 ( \23062 , \16334 , RIfe98a78_8081);
and \g453183/U$3 ( \23063 , RIf154b08_5423, \16380 );
nor \g453183/U$1 ( \23064 , \23062 , \23063 );
nand \g447401/U$1 ( \23065 , \23050 , \23058 , \23061 , \23064 );
nor \g446293/U$1 ( \23066 , \23045 , \23046 , \23065 );
and \g453177/U$2 ( \23067 , \16361 , RIe1ef240_4098);
and \g453177/U$3 ( \23068 , RIf1538c0_5410, \16448 );
nor \g453177/U$1 ( \23069 , \23067 , \23068 );
and \g453176/U$2 ( \23070 , \16364 , RIf14e2f8_5349);
and \g453176/U$3 ( \23071 , RIf150e90_5380, \16371 );
nor \g453176/U$1 ( \23072 , \23070 , \23071 );
and \g445359/U$2 ( \23073 , \23066 , \23069 , \23072 );
nor \g445359/U$1 ( \23074 , \23073 , \16480 );
or \g444180/U$1 ( \23075 , \23014 , \23044 , \23074 );
_DC \g40e4/U$1 ( \23076 , \23075 , \16652 );
and \g453335/U$2 ( \23077 , \16377 , RIfe97830_8068);
and \g453335/U$3 ( \23078 , RIfc9f980_6838, \16380 );
nor \g453335/U$1 ( \23079 , \23077 , \23078 );
and \g446324/U$2 ( \23080 , RIf1412d8_5201, \16321 );
and \g446324/U$3 ( \23081 , RIfcc4118_7253, \16313 );
and \g449299/U$2 ( \23082 , RIfce27a8_7599, \16398 );
and \g449299/U$3 ( \23083 , \16339 , RIfc4a408_5867);
and \g449299/U$4 ( \23084 , RIf13f6b8_5181, \16485 );
nor \g449299/U$1 ( \23085 , \23082 , \23083 , \23084 );
and \g455244/U$2 ( \23086 , \16317 , RIfc89e28_6591);
and \g455244/U$3 ( \23087 , RIfcc3e48_7251, \16325 );
nor \g455244/U$1 ( \23088 , \23086 , \23087 );
not \g450316/U$3 ( \23089 , \23088 );
not \g450316/U$4 ( \23090 , \16351 );
and \g450316/U$2 ( \23091 , \23089 , \23090 );
and \g450316/U$5 ( \23092 , \16354 , RIfc4a6d8_5869);
nor \g450316/U$1 ( \23093 , \23091 , \23092 );
and \g453337/U$2 ( \23094 , \16361 , RIfcd5d28_7455);
and \g453337/U$3 ( \23095 , RIfc530a8_5967, \16364 );
nor \g453337/U$1 ( \23096 , \23094 , \23095 );
and \g453336/U$2 ( \23097 , \16368 , RIe174720_2702);
and \g453336/U$3 ( \23098 , RIfc89cc0_6590, \16371 );
nor \g453336/U$1 ( \23099 , \23097 , \23098 );
nand \g447883/U$1 ( \23100 , \23085 , \23093 , \23096 , \23099 );
nor \g446324/U$1 ( \23101 , \23080 , \23081 , \23100 );
and \g453334/U$2 ( \23102 , \16334 , RIfc9fae8_6839);
and \g453334/U$3 ( \23103 , RIfcd3730_7428, \16326 );
nor \g453334/U$1 ( \23104 , \23102 , \23103 );
nand \g445659/U$1 ( \23105 , \23079 , \23101 , \23104 );
and \g444796/U$2 ( \23106 , \23105 , \17998 );
and \g449297/U$2 ( \23107 , RIe213e10_4516, \16427 );
and \g449297/U$3 ( \23108 , \16432 , RIfc401d8_5755);
and \g449297/U$4 ( \23109 , RIe21f210_4644, \16485 );
nor \g449297/U$1 ( \23110 , \23107 , \23108 , \23109 );
and \g455249/U$2 ( \23111 , \16317 , RIe20e410_4452);
and \g455249/U$3 ( \23112 , RIfc81cc8_6499, \16325 );
nor \g455249/U$1 ( \23113 , \23111 , \23112 );
not \g455248/U$1 ( \23114 , \23113 );
and \g450315/U$2 ( \23115 , \23114 , \16336 );
and \g450315/U$3 ( \23116 , RIf16b1a0_5678, \16354 );
nor \g450315/U$1 ( \23117 , \23115 , \23116 );
and \g453331/U$2 ( \23118 , \16361 , RIe208a10_4388);
and \g453331/U$3 ( \23119 , RIe20b710_4420, \16364 );
nor \g453331/U$1 ( \23120 , \23118 , \23119 );
and \g453330/U$2 ( \23121 , \16368 , RIe211110_4484);
and \g453330/U$3 ( \23122 , RIf1699b8_5661, \16371 );
nor \g453330/U$1 ( \23123 , \23121 , \23122 );
nand \g448104/U$1 ( \23124 , \23110 , \23117 , \23120 , \23123 );
and \g444796/U$3 ( \23125 , \16390 , \23124 );
nor \g444796/U$1 ( \23126 , \23106 , \23125 );
and \g447088/U$2 ( \23127 , \18020 , RIe224c10_4708);
and \g447088/U$3 ( \23128 , RIf16cf28_5699, \18022 );
nor \g447088/U$1 ( \23129 , \23127 , \23128 );
and \g447089/U$2 ( \23130 , \18025 , RIe221f10_4676);
and \g447089/U$3 ( \23131 , RIfc53210_5968, \18027 );
nor \g447089/U$1 ( \23132 , \23130 , \23131 );
and \g447090/U$2 ( \23133 , \18030 , RIe216b10_4548);
and \g447090/U$3 ( \23134 , RIe219810_4580, \18032 );
nor \g447090/U$1 ( \23135 , \23133 , \23134 );
nand \g444527/U$1 ( \23136 , \23126 , \23129 , \23132 , \23135 );
and \g453352/U$2 ( \23137 , \16377 , RIe1a15b8_3213);
and \g453352/U$3 ( \23138 , RIe227910_4740, \16380 );
nor \g453352/U$1 ( \23139 , \23137 , \23138 );
and \g446328/U$2 ( \23140 , RIe1a6fb8_3277, \16321 );
and \g446328/U$3 ( \23141 , RIe1a42b8_3245, \16313 );
and \g449302/U$2 ( \23142 , RIe1bcc78_3525, \16398 );
and \g449302/U$3 ( \23143 , \16339 , RIe1d6178_3813);
and \g449302/U$4 ( \23144 , RIe179fb8_2765, \16344 );
nor \g449302/U$1 ( \23145 , \23142 , \23143 , \23144 );
and \g455316/U$2 ( \23146 , \16317 , RIe1ffd70_4288);
and \g455316/U$3 ( \23147 , RIe205d10_4356, \16325 );
nor \g455316/U$1 ( \23148 , \23146 , \23147 );
not \g450319/U$3 ( \23149 , \23148 );
not \g450319/U$4 ( \23150 , \16351 );
and \g450319/U$2 ( \23151 , \23149 , \23150 );
and \g450319/U$5 ( \23152 , \16354 , RIe18dab8_2989);
nor \g450319/U$1 ( \23153 , \23151 , \23152 );
and \g453355/U$2 ( \23154 , \16361 , RIe172128_2675);
and \g453355/U$3 ( \23155 , RIe1afaf0_3376, \16364 );
nor \g453355/U$1 ( \23156 , \23154 , \23155 );
and \g453354/U$2 ( \23157 , \16368 , RIe1f1c70_4128);
and \g453354/U$3 ( \23158 , RIe1f9128_4211, \16371 );
nor \g453354/U$1 ( \23159 , \23157 , \23158 );
nand \g447885/U$1 ( \23160 , \23145 , \23153 , \23156 , \23159 );
nor \g446328/U$1 ( \23161 , \23140 , \23141 , \23160 );
and \g453350/U$2 ( \23162 , \16334 , RIe21c510_4612);
and \g453350/U$3 ( \23163 , RIe1a9cb8_3309, \16328 );
nor \g453350/U$1 ( \23164 , \23162 , \23163 );
nand \g445661/U$1 ( \23165 , \23139 , \23161 , \23164 );
and \g444896/U$2 ( \23166 , \23165 , \16752 );
and \g449301/U$2 ( \23167 , RIfcc3a10_7248, \16427 );
and \g449301/U$3 ( \23168 , \16448 , RIfce5610_7632);
and \g449301/U$4 ( \23169 , RIfcbb5e0_7154, \16485 );
nor \g449301/U$1 ( \23170 , \23167 , \23168 , \23169 );
and \g454299/U$2 ( \23171 , \16317 , RIfc81188_6491);
and \g454299/U$3 ( \23172 , RIfc495f8_5857, \16325 );
nor \g454299/U$1 ( \23173 , \23171 , \23172 );
not \g454298/U$1 ( \23174 , \23173 );
and \g450318/U$2 ( \23175 , \23174 , \16336 );
and \g450318/U$3 ( \23176 , RIfce0a20_7578, \16356 );
nor \g450318/U$1 ( \23177 , \23175 , \23176 );
and \g453345/U$2 ( \23178 , \16361 , RIe1aba40_3330);
and \g453345/U$3 ( \23179 , RIe1ad228_3347, \16364 );
nor \g453345/U$1 ( \23180 , \23178 , \23179 );
and \g453344/U$2 ( \23181 , \16368 , RIe1b19e0_3398);
and \g453344/U$3 ( \23182 , RIe1b3330_3416, \16371 );
nor \g453344/U$1 ( \23183 , \23181 , \23182 );
nand \g448106/U$1 ( \23184 , \23170 , \23177 , \23180 , \23183 );
and \g444896/U$3 ( \23185 , \16477 , \23184 );
nor \g444896/U$1 ( \23186 , \23166 , \23185 );
and \g447094/U$2 ( \23187 , \18268 , RIfcb6018_7093);
and \g447094/U$3 ( \23188 , RIfc49a30_5860, \18270 );
nor \g447094/U$1 ( \23189 , \23187 , \23188 );
and \g447095/U$2 ( \23190 , \18273 , RIe1b81f0_3472);
and \g447095/U$3 ( \23191 , RIe1ba3b0_3496, \18275 );
nor \g447095/U$1 ( \23192 , \23190 , \23191 );
and \g447096/U$2 ( \23193 , \18278 , RIfe97998_8069);
and \g447096/U$3 ( \23194 , RIe1b6030_3448, \18280 );
nor \g447096/U$1 ( \23195 , \23193 , \23194 );
nand \g444650/U$1 ( \23196 , \23186 , \23189 , \23192 , \23195 );
and \g446319/U$2 ( \23197 , RIe19bbb8_3149, \16321 );
and \g446319/U$3 ( \23198 , RIfe976c8_8067, \16313 );
and \g449293/U$2 ( \23199 , RIe1880b8_2925, \16427 );
and \g449293/U$3 ( \23200 , \16448 , RIe18adb8_2957);
and \g449293/U$4 ( \23201 , RIe1961b8_3085, \16344 );
nor \g449293/U$1 ( \23202 , \23199 , \23200 , \23201 );
and \g454355/U$2 ( \23203 , \16317 , RIe1826b8_2861);
and \g454355/U$3 ( \23204 , RIfcc3fb0_7252, \16325 );
nor \g454355/U$1 ( \23205 , \23203 , \23204 );
not \g454354/U$1 ( \23206 , \23205 );
and \g450309/U$2 ( \23207 , \23206 , \16336 );
and \g450309/U$3 ( \23208 , RIf144c80_5242, \16356 );
nor \g450309/U$1 ( \23209 , \23207 , \23208 );
and \g453316/U$2 ( \23210 , \16361 , RIe17ccb8_2797);
and \g453316/U$3 ( \23211 , RIe17f9b8_2829, \16364 );
nor \g453316/U$1 ( \23212 , \23210 , \23211 );
and \g453315/U$2 ( \23213 , \16368 , RIe1853b8_2893);
and \g453315/U$3 ( \23214 , RIfe97560_8066, \16371 );
nor \g453315/U$1 ( \23215 , \23213 , \23214 );
nand \g448103/U$1 ( \23216 , \23202 , \23209 , \23212 , \23215 );
nor \g446319/U$1 ( \23217 , \23197 , \23198 , \23216 );
and \g453311/U$2 ( \23218 , \16377 , RIe198eb8_3117);
and \g453311/U$3 ( \23219 , RIe1934b8_3053, \16380 );
nor \g453311/U$1 ( \23220 , \23218 , \23219 );
and \g453310/U$2 ( \23221 , \16334 , RIe1907b8_3021);
and \g453310/U$3 ( \23222 , RIe19e8b8_3181, \16328 );
nor \g453310/U$1 ( \23223 , \23221 , \23222 );
and \g445378/U$2 ( \23224 , \23217 , \23220 , \23223 );
nor \g445378/U$1 ( \23225 , \23224 , \16618 );
and \g446322/U$2 ( \23226 , RIf160bb0_5560, \16448 );
and \g446322/U$3 ( \23227 , RIe1fd4a8_4259, \16371 );
and \g449295/U$2 ( \23228 , RIfc8a3c8_6595, \16485 );
and \g449295/U$3 ( \23229 , \16354 , RIfc53378_5969);
and \g449295/U$4 ( \23230 , RIfe97c68_8071, \16398 );
nor \g449295/U$1 ( \23231 , \23228 , \23229 , \23230 );
and \g455251/U$2 ( \23232 , \16317 , RIfcb6720_7098);
and \g455251/U$3 ( \23233 , RIfc8a0f8_6593, \16325 );
nor \g455251/U$1 ( \23234 , \23232 , \23233 );
not \g450311/U$3 ( \23235 , \23234 );
not \g450311/U$4 ( \23236 , \16311 );
and \g450311/U$2 ( \23237 , \23235 , \23236 );
and \g450311/U$5 ( \23238 , \16341 , RIfc8a530_6596);
nor \g450311/U$1 ( \23239 , \23237 , \23238 );
and \g453324/U$2 ( \23240 , \16377 , RIe201828_4307);
and \g453324/U$3 ( \23241 , RIe203448_4327, \16313 );
nor \g453324/U$1 ( \23242 , \23240 , \23241 );
and \g453325/U$2 ( \23243 , \16334 , RIfc49fd0_5864);
and \g453325/U$3 ( \23244 , RIfcb65b8_7097, \16380 );
nor \g453325/U$1 ( \23245 , \23243 , \23244 );
nand \g447410/U$1 ( \23246 , \23231 , \23239 , \23242 , \23245 );
nor \g446322/U$1 ( \23247 , \23226 , \23227 , \23246 );
and \g453321/U$2 ( \23248 , \16364 , RIfc8a800_6598);
and \g453321/U$3 ( \23249 , RIfe97b00_8070, \16368 );
nor \g453321/U$1 ( \23250 , \23248 , \23249 );
and \g453322/U$2 ( \23251 , \16361 , RIfc8a698_6597);
and \g453322/U$3 ( \23252 , RIf15ecc0_5538, \16427 );
nor \g453322/U$1 ( \23253 , \23251 , \23252 );
and \g445379/U$2 ( \23254 , \23247 , \23250 , \23253 );
nor \g445379/U$1 ( \23255 , \23254 , \16393 );
or \g444408/U$1 ( \23256 , \23136 , \23196 , \23225 , \23255 );
and \g446315/U$2 ( \23257 , RIfcd3460_7426, \16448 );
and \g446315/U$3 ( \23258 , RIfc9a520_6778, \16371 );
and \g449289/U$2 ( \23259 , RIfc81890_6496, \16319 );
and \g449289/U$3 ( \23260 , \16328 , RIfc9a7f0_6780);
and \g449289/U$4 ( \23261 , RIfcd9dd8_7501, \16398 );
nor \g449289/U$1 ( \23262 , \23259 , \23260 , \23261 );
and \g455265/U$2 ( \23263 , \16317 , RIfc81728_6495);
and \g455265/U$3 ( \23264 , RIfc49e68_5863, \16325 );
nor \g455265/U$1 ( \23265 , \23263 , \23264 );
not \g450306/U$3 ( \23266 , \23265 );
not \g450306/U$4 ( \23267 , \16330 );
and \g450306/U$2 ( \23268 , \23266 , \23267 );
and \g450306/U$5 ( \23269 , \16341 , RIfc49d00_5862);
nor \g450306/U$1 ( \23270 , \23268 , \23269 );
and \g453296/U$2 ( \23271 , \16377 , RIe1fb180_4234);
and \g453296/U$3 ( \23272 , RIfcd5e90_7456, \16313 );
nor \g453296/U$1 ( \23273 , \23271 , \23272 );
and \g453297/U$2 ( \23274 , \16334 , RIe1f66f8_4181);
and \g453297/U$3 ( \23275 , RIfcbb1a8_7151, \16380 );
nor \g453297/U$1 ( \23276 , \23274 , \23275 );
nand \g447407/U$1 ( \23277 , \23262 , \23270 , \23273 , \23276 );
nor \g446315/U$1 ( \23278 , \23257 , \23258 , \23277 );
and \g453292/U$2 ( \23279 , \16364 , RIfcbb310_7152);
and \g453292/U$3 ( \23280 , RIe1f4268_4155, \16368 );
nor \g453292/U$1 ( \23281 , \23279 , \23280 );
and \g453295/U$2 ( \23282 , \16361 , RIe1ef0d8_4097);
and \g453295/U$3 ( \23283 , RIfcb62e8_7095, \16427 );
nor \g453295/U$1 ( \23284 , \23282 , \23283 );
and \g445374/U$2 ( \23285 , \23278 , \23281 , \23284 );
nor \g445374/U$1 ( \23286 , \23285 , \16480 );
and \g446317/U$2 ( \23287 , RIe1d0778_3749, \16427 );
and \g446317/U$3 ( \23288 , RIe1cad78_3685, \16368 );
and \g449291/U$2 ( \23289 , RIe1de878_3909, \16344 );
and \g449291/U$3 ( \23290 , \16356 , RIe1e1578_3941);
and \g449291/U$4 ( \23291 , RIe1c5378_3621, \16337 );
nor \g449291/U$1 ( \23292 , \23289 , \23290 , \23291 );
and \g455259/U$2 ( \23293 , \16317 , RIe1e9c78_4037);
and \g455259/U$3 ( \23294 , RIe1ec978_4069, \16325 );
nor \g455259/U$1 ( \23295 , \23293 , \23294 );
not \g450307/U$3 ( \23296 , \23295 );
not \g450307/U$4 ( \23297 , \16311 );
and \g450307/U$2 ( \23298 , \23296 , \23297 );
and \g450307/U$5 ( \23299 , \16339 , RIe1c8078_3653);
nor \g450307/U$1 ( \23300 , \23298 , \23299 );
and \g453305/U$2 ( \23301 , \16377 , RIe1e4278_3973);
and \g453305/U$3 ( \23302 , RIe1e6f78_4005, \16313 );
nor \g453305/U$1 ( \23303 , \23301 , \23302 );
and \g453306/U$2 ( \23304 , \16334 , RIe1d8e78_3845);
and \g453306/U$3 ( \23305 , RIe1dbb78_3877, \16380 );
nor \g453306/U$1 ( \23306 , \23304 , \23305 );
nand \g447408/U$1 ( \23307 , \23292 , \23300 , \23303 , \23306 );
nor \g446317/U$1 ( \23308 , \23287 , \23288 , \23307 );
and \g453303/U$2 ( \23309 , \16361 , RIe1bf978_3557);
and \g453303/U$3 ( \23310 , RIe1d3478_3781, \16448 );
nor \g453303/U$1 ( \23311 , \23309 , \23310 );
and \g453302/U$2 ( \23312 , \16364 , RIe1c2678_3589);
and \g453302/U$3 ( \23313 , RIe1cda78_3717, \16371 );
nor \g453302/U$1 ( \23314 , \23312 , \23313 );
and \g445376/U$2 ( \23315 , \23308 , \23311 , \23314 );
nor \g445376/U$1 ( \23316 , \23315 , \16555 );
or \g444264/U$1 ( \23317 , \23256 , \23286 , \23316 );
_DC \g4169/U$1 ( \23318 , \23317 , \16652 );
and \g448524/U$2 ( \23319 , RIe19ba50_3148, \16321 );
and \g448524/U$3 ( \23320 , \16328 , RIe19e750_3180);
and \g448524/U$4 ( \23321 , RIe182550_2860, \16398 );
nor \g448524/U$1 ( \23322 , \23319 , \23320 , \23321 );
and \g454293/U$2 ( \23323 , \16317 , RIe196050_3084);
and \g454293/U$3 ( \23324 , RIfe9f558_8157, \16325 );
nor \g454293/U$1 ( \23325 , \23323 , \23324 );
not \g449547/U$3 ( \23326 , \23325 );
not \g449547/U$4 ( \23327 , \16330 );
and \g449547/U$2 ( \23328 , \23326 , \23327 );
and \g449547/U$5 ( \23329 , \16339 , RIf142ef8_5221);
nor \g449547/U$1 ( \23330 , \23328 , \23329 );
and \g450668/U$2 ( \23331 , \16377 , RIe198d50_3116);
and \g450668/U$3 ( \23332 , RIfc479d8_5837, \16313 );
nor \g450668/U$1 ( \23333 , \23331 , \23332 );
and \g450670/U$2 ( \23334 , \16334 , RIe190650_3020);
and \g450670/U$3 ( \23335 , RIe193350_3052, \16380 );
nor \g450670/U$1 ( \23336 , \23334 , \23335 );
nand \g447239/U$1 ( \23337 , \23322 , \23330 , \23333 , \23336 );
and \g444700/U$2 ( \23338 , \23337 , \17938 );
and \g445726/U$2 ( \23339 , RIfcb4dd0_7080, \16427 );
and \g445726/U$3 ( \23340 , RIe1fc260_4246, \16368 );
and \g448527/U$2 ( \23341 , RIfc7eb90_6464, \16485 );
and \g448527/U$3 ( \23342 , \16356 , RIfc98ea0_6762);
and \g448527/U$4 ( \23343 , RIfe9f120_8154, \16337 );
nor \g448527/U$1 ( \23344 , \23341 , \23342 , \23343 );
and \g454269/U$2 ( \23345 , \16317 , RIfcd6598_7461);
and \g454269/U$3 ( \23346 , RIfc46bc8_5827, \16325 );
nor \g454269/U$1 ( \23347 , \23345 , \23346 );
not \g449548/U$3 ( \23348 , \23347 );
not \g449548/U$4 ( \23349 , \16311 );
and \g449548/U$2 ( \23350 , \23348 , \23349 );
and \g449548/U$5 ( \23351 , \16341 , RIf15cf38_5517);
nor \g449548/U$1 ( \23352 , \23350 , \23351 );
and \g450673/U$2 ( \23353 , \16377 , RIe2016c0_4306);
and \g450673/U$3 ( \23354 , RIe2032e0_4326, \16313 );
nor \g450673/U$1 ( \23355 , \23353 , \23354 );
and \g450674/U$2 ( \23356 , \16334 , RIfcbcaf8_7169);
and \g450674/U$3 ( \23357 , RIfce0318_7573, \16380 );
nor \g450674/U$1 ( \23358 , \23356 , \23357 );
nand \g447240/U$1 ( \23359 , \23344 , \23352 , \23355 , \23358 );
nor \g445726/U$1 ( \23360 , \23339 , \23340 , \23359 );
and \g450672/U$2 ( \23361 , \16361 , RIfc8d0c8_6627);
and \g450672/U$3 ( \23362 , RIfc8cf60_6626, \16448 );
nor \g450672/U$1 ( \23363 , \23361 , \23362 );
and \g450671/U$2 ( \23364 , \16364 , RIfc7ea28_6463);
and \g450671/U$3 ( \23365 , RIe1fd340_4258, \16371 );
nor \g450671/U$1 ( \23366 , \23364 , \23365 );
and \g444948/U$2 ( \23367 , \23360 , \23363 , \23366 );
nor \g444948/U$1 ( \23368 , \23367 , \16393 );
nor \g444700/U$1 ( \23369 , \23338 , \23368 );
and \g446526/U$2 ( \23370 , \18457 , RIe187f50_2924);
and \g446526/U$3 ( \23371 , RIe18ac50_2956, \18459 );
nor \g446526/U$1 ( \23372 , \23370 , \23371 );
and \g446527/U$2 ( \23373 , \18462 , RIe185250_2892);
and \g446527/U$3 ( \23374 , RIfc47870_5836, \18464 );
nor \g446527/U$1 ( \23375 , \23373 , \23374 );
and \g446528/U$2 ( \23376 , \18467 , RIe17cb50_2796);
and \g446528/U$3 ( \23377 , RIe17f850_2828, \18469 );
nor \g446528/U$1 ( \23378 , \23376 , \23377 );
nand \g444447/U$1 ( \23379 , \23369 , \23372 , \23375 , \23378 );
and \g450684/U$2 ( \23380 , \16364 , RIe1c2510_3588);
and \g450684/U$3 ( \23381 , RIe1cd910_3716, \16371 );
nor \g450684/U$1 ( \23382 , \23380 , \23381 );
and \g445729/U$2 ( \23383 , RIe1d0610_3748, \16427 );
and \g445729/U$3 ( \23384 , RIe1cac10_3684, \16368 );
and \g448529/U$2 ( \23385 , RIe1e9b10_4036, \16319 );
and \g448529/U$3 ( \23386 , \16326 , RIe1ec810_4068);
and \g448529/U$4 ( \23387 , RIe1c5210_3620, \16398 );
nor \g448529/U$1 ( \23388 , \23385 , \23386 , \23387 );
and \g454215/U$2 ( \23389 , \16317 , RIe1de710_3908);
and \g454215/U$3 ( \23390 , RIe1e1410_3940, \16325 );
nor \g454215/U$1 ( \23391 , \23389 , \23390 );
not \g449551/U$3 ( \23392 , \23391 );
not \g449551/U$4 ( \23393 , \16330 );
and \g449551/U$2 ( \23394 , \23392 , \23393 );
and \g449551/U$5 ( \23395 , \16341 , RIe1c7f10_3652);
nor \g449551/U$1 ( \23396 , \23394 , \23395 );
and \g450688/U$2 ( \23397 , \16377 , RIe1e4110_3972);
and \g450688/U$3 ( \23398 , RIe1e6e10_4004, \16313 );
nor \g450688/U$1 ( \23399 , \23397 , \23398 );
and \g450689/U$2 ( \23400 , \16334 , RIe1d8d10_3844);
and \g450689/U$3 ( \23401 , RIe1dba10_3876, \16380 );
nor \g450689/U$1 ( \23402 , \23400 , \23401 );
nand \g447241/U$1 ( \23403 , \23388 , \23396 , \23399 , \23402 );
nor \g445729/U$1 ( \23404 , \23383 , \23384 , \23403 );
and \g450686/U$2 ( \23405 , \16361 , RIe1bf810_3556);
and \g450686/U$3 ( \23406 , RIe1d3310_3780, \16432 );
nor \g450686/U$1 ( \23407 , \23405 , \23406 );
nand \g445513/U$1 ( \23408 , \23382 , \23404 , \23407 );
and \g444753/U$2 ( \23409 , \23408 , \16750 );
and \g448528/U$2 ( \23410 , RIfc8d398_6629, \16337 );
and \g448528/U$3 ( \23411 , \16339 , RIfceedf0_7740);
and \g448528/U$4 ( \23412 , RIfc7e8c0_6462, \16485 );
nor \g448528/U$1 ( \23413 , \23410 , \23411 , \23412 );
and \g454236/U$2 ( \23414 , \16317 , RIfc468f8_5825);
and \g454236/U$3 ( \23415 , RIfce58e0_7634, \16325 );
nor \g454236/U$1 ( \23416 , \23414 , \23415 );
not \g449549/U$3 ( \23417 , \23416 );
not \g449549/U$4 ( \23418 , \16351 );
and \g449549/U$2 ( \23419 , \23417 , \23418 );
and \g449549/U$5 ( \23420 , \16354 , RIfc55f10_6000);
nor \g449549/U$1 ( \23421 , \23419 , \23420 );
and \g450680/U$2 ( \23422 , \16361 , RIe1eef70_4096);
and \g450680/U$3 ( \23423 , RIfc8d500_6630, \16364 );
nor \g450680/U$1 ( \23424 , \23422 , \23423 );
and \g450679/U$2 ( \23425 , \16368 , RIe1f4100_4154);
and \g450679/U$3 ( \23426 , RIfcc2ed0_7240, \16371 );
nor \g450679/U$1 ( \23427 , \23425 , \23426 );
nand \g447471/U$1 ( \23428 , \23413 , \23421 , \23424 , \23427 );
and \g444753/U$3 ( \23429 , \16481 , \23428 );
nor \g444753/U$1 ( \23430 , \23409 , \23429 );
and \g446530/U$2 ( \23431 , \16505 , RIfc98bd0_6760);
and \g446530/U$3 ( \23432 , RIfcbcc60_7170, \16507 );
nor \g446530/U$1 ( \23433 , \23431 , \23432 );
and \g446531/U$2 ( \23434 , \16511 , RIe1f6590_4180);
and \g446531/U$3 ( \23435 , RIfc8d230_6628, \16514 );
nor \g446531/U$1 ( \23436 , \23434 , \23435 );
and \g446529/U$2 ( \23437 , \16518 , RIe1fb018_4233);
and \g446529/U$3 ( \23438 , RIfce2d48_7603, \16521 );
nor \g446529/U$1 ( \23439 , \23437 , \23438 );
nand \g444448/U$1 ( \23440 , \23430 , \23433 , \23436 , \23439 );
and \g445722/U$2 ( \23441 , RIe224aa8_4707, \16319 );
and \g445722/U$3 ( \23442 , RIfc55808_5995, \16313 );
and \g448521/U$2 ( \23443 , RIe213ca8_4515, \16427 );
and \g448521/U$3 ( \23444 , \16448 , RIfcbc828_7167);
and \g448521/U$4 ( \23445 , RIe21f0a8_4643, \16485 );
nor \g448521/U$1 ( \23446 , \23443 , \23444 , \23445 );
and \g454201/U$2 ( \23447 , \16317 , RIe20e2a8_4451);
and \g454201/U$3 ( \23448 , RIfcbc990_7168, \16325 );
nor \g454201/U$1 ( \23449 , \23447 , \23448 );
not \g454200/U$1 ( \23450 , \23449 );
and \g449543/U$2 ( \23451 , \23450 , \16336 );
and \g449543/U$3 ( \23452 , RIfcb50a0_7082, \16356 );
nor \g449543/U$1 ( \23453 , \23451 , \23452 );
and \g450655/U$2 ( \23454 , \16361 , RIe2088a8_4387);
and \g450655/U$3 ( \23455 , RIe20b5a8_4419, \16364 );
nor \g450655/U$1 ( \23456 , \23454 , \23455 );
and \g450654/U$2 ( \23457 , \16368 , RIe210fa8_4483);
and \g450654/U$3 ( \23458 , RIfc47000_5830, \16371 );
nor \g450654/U$1 ( \23459 , \23457 , \23458 );
nand \g448007/U$1 ( \23460 , \23446 , \23453 , \23456 , \23459 );
nor \g445722/U$1 ( \23461 , \23441 , \23442 , \23460 );
and \g450653/U$2 ( \23462 , \16377 , RIe221da8_4675);
and \g450653/U$3 ( \23463 , RIe2196a8_4579, \16380 );
nor \g450653/U$1 ( \23464 , \23462 , \23463 );
and \g450652/U$2 ( \23465 , \16334 , RIe2169a8_4547);
and \g450652/U$3 ( \23466 , RIfe9f288_8155, \16328 );
nor \g450652/U$1 ( \23467 , \23465 , \23466 );
and \g444944/U$2 ( \23468 , \23461 , \23464 , \23467 );
nor \g444944/U$1 ( \23469 , \23468 , \16389 );
and \g445725/U$2 ( \23470 , RIfca15a0_6858, \16427 );
and \g445725/U$3 ( \23471 , RIe1745b8_2701, \16368 );
and \g448522/U$2 ( \23472 , RIfcbc6c0_7166, \16321 );
and \g448522/U$3 ( \23473 , \16326 , RIfcb5208_7083);
and \g448522/U$4 ( \23474 , RIfc556a0_5994, \16398 );
nor \g448522/U$1 ( \23475 , \23472 , \23473 , \23474 );
and \g454203/U$2 ( \23476 , \16317 , RIfe9f3f0_8156);
and \g454203/U$3 ( \23477 , RIf13fdc0_5186, \16325 );
nor \g454203/U$1 ( \23478 , \23476 , \23477 );
not \g449544/U$3 ( \23479 , \23478 );
not \g449544/U$4 ( \23480 , \16330 );
and \g449544/U$2 ( \23481 , \23479 , \23480 );
and \g449544/U$5 ( \23482 , \16339 , RIfc8cc90_6624);
nor \g449544/U$1 ( \23483 , \23481 , \23482 );
and \g450662/U$2 ( \23484 , \16377 , RIe176610_2724);
and \g450662/U$3 ( \23485 , RIe177588_2735, \16313 );
nor \g450662/U$1 ( \23486 , \23484 , \23485 );
and \g450663/U$2 ( \23487 , \16334 , RIfc47708_5835);
and \g450663/U$3 ( \23488 , RIfce40f8_7617, \16380 );
nor \g450663/U$1 ( \23489 , \23487 , \23488 );
nand \g447237/U$1 ( \23490 , \23475 , \23483 , \23486 , \23489 );
nor \g445725/U$1 ( \23491 , \23470 , \23471 , \23490 );
and \g450659/U$2 ( \23492 , \16361 , RIfce8e50_7672);
and \g450659/U$3 ( \23493 , RIfc47438_5833, \16448 );
nor \g450659/U$1 ( \23494 , \23492 , \23493 );
and \g450658/U$2 ( \23495 , \16364 , RIfc7ee60_6466);
and \g450658/U$3 ( \23496 , RIfc99170_6764, \16371 );
nor \g450658/U$1 ( \23497 , \23495 , \23496 );
and \g444946/U$2 ( \23498 , \23491 , \23494 , \23497 );
nor \g444946/U$1 ( \23499 , \23498 , \16649 );
or \g444338/U$1 ( \23500 , \23379 , \23440 , \23469 , \23499 );
and \g445720/U$2 ( \23501 , RIfcb4c68_7079, \16427 );
and \g445720/U$3 ( \23502 , RIfe9ee50_8152, \16368 );
and \g448517/U$2 ( \23503 , RIfe9efb8_8153, \16321 );
and \g448517/U$3 ( \23504 , \16328 , RIf14d0b0_5336);
and \g448517/U$4 ( \23505 , RIfc46358_5821, \16337 );
nor \g448517/U$1 ( \23506 , \23503 , \23504 , \23505 );
and \g454194/U$2 ( \23507 , \16317 , RIfec50a0_8362);
and \g454194/U$3 ( \23508 , RIfec4dd0_8360, \16325 );
nor \g454194/U$1 ( \23509 , \23507 , \23508 );
not \g449539/U$3 ( \23510 , \23509 );
not \g449539/U$4 ( \23511 , \16330 );
and \g449539/U$2 ( \23512 , \23510 , \23511 );
and \g449539/U$5 ( \23513 , \16341 , RIfcbcdc8_7171);
nor \g449539/U$1 ( \23514 , \23512 , \23513 );
and \g450642/U$2 ( \23515 , \16377 , RIe1b8088_3471);
and \g450642/U$3 ( \23516 , RIe1ba248_3495, \16313 );
nor \g450642/U$1 ( \23517 , \23515 , \23516 );
and \g450643/U$2 ( \23518 , \16334 , RIe1b46e0_3430);
and \g450643/U$3 ( \23519 , RIe1b5ec8_3447, \16380 );
nor \g450643/U$1 ( \23520 , \23518 , \23519 );
nand \g447235/U$1 ( \23521 , \23506 , \23514 , \23517 , \23520 );
nor \g445720/U$1 ( \23522 , \23501 , \23502 , \23521 );
and \g450640/U$2 ( \23523 , \16361 , RIfec4f38_8361);
and \g450640/U$3 ( \23524 , RIfcb4998_7077, \16448 );
nor \g450640/U$1 ( \23525 , \23523 , \23524 );
and \g450639/U$2 ( \23526 , \16364 , RIfec5208_8363);
and \g450639/U$3 ( \23527 , RIfec5370_8364, \16371 );
nor \g450639/U$1 ( \23528 , \23526 , \23527 );
and \g444942/U$2 ( \23529 , \23522 , \23525 , \23528 );
nor \g444942/U$1 ( \23530 , \23529 , \16909 );
and \g445721/U$2 ( \23531 , RIe1ffc08_4287, \16427 );
and \g445721/U$3 ( \23532 , RIe1f1b08_4127, \16368 );
and \g448520/U$2 ( \23533 , RIe1a6e50_3276, \16319 );
and \g448520/U$3 ( \23534 , \16328 , RIe1a9b50_3308);
and \g448520/U$4 ( \23535 , RIe1bcb10_3524, \16398 );
nor \g448520/U$1 ( \23536 , \23533 , \23534 , \23535 );
and \g454376/U$2 ( \23537 , \16317 , RIe179e50_2764);
and \g454376/U$3 ( \23538 , RIe18d950_2988, \16325 );
nor \g454376/U$1 ( \23539 , \23537 , \23538 );
not \g449542/U$3 ( \23540 , \23539 );
not \g449542/U$4 ( \23541 , \16330 );
and \g449542/U$2 ( \23542 , \23540 , \23541 );
and \g449542/U$5 ( \23543 , \16339 , RIe1d6010_3812);
nor \g449542/U$1 ( \23544 , \23542 , \23543 );
and \g450649/U$2 ( \23545 , \16377 , RIe1a1450_3212);
and \g450649/U$3 ( \23546 , RIe1a4150_3244, \16313 );
nor \g450649/U$1 ( \23547 , \23545 , \23546 );
and \g450650/U$2 ( \23548 , \16334 , RIe21c3a8_4611);
and \g450650/U$3 ( \23549 , RIe2277a8_4739, \16380 );
nor \g450650/U$1 ( \23550 , \23548 , \23549 );
nand \g447236/U$1 ( \23551 , \23536 , \23544 , \23547 , \23550 );
nor \g445721/U$1 ( \23552 , \23531 , \23532 , \23551 );
and \g450646/U$2 ( \23553 , \16361 , RIe171fc0_2674);
and \g450646/U$3 ( \23554 , RIe205ba8_4355, \16448 );
nor \g450646/U$1 ( \23555 , \23553 , \23554 );
and \g450645/U$2 ( \23556 , \16364 , RIe1af988_3375);
and \g450645/U$3 ( \23557 , RIe1f8fc0_4210, \16371 );
nor \g450645/U$1 ( \23558 , \23556 , \23557 );
and \g444943/U$2 ( \23559 , \23552 , \23555 , \23558 );
nor \g444943/U$1 ( \23560 , \23559 , \16586 );
or \g444165/U$1 ( \23561 , \23500 , \23530 , \23560 );
_DC \g41ee/U$1 ( \23562 , \23561 , \16652 );
and \g452586/U$2 ( \23563 , \16371 , RIe1f8b88_4207);
and \g452586/U$3 ( \23564 , RIe1ff7d0_4284, \16427 );
nor \g452586/U$1 ( \23565 , \23563 , \23564 );
and \g445946/U$2 ( \23566 , RIe205770_4352, \16432 );
and \g445946/U$3 ( \23567 , RIe171b88_2671, \16361 );
and \g448809/U$2 ( \23568 , RIe179a18_2761, \16485 );
and \g448809/U$3 ( \23569 , \16354 , RIe18d518_2985);
and \g448809/U$4 ( \23570 , RIe1bc6d8_3521, \16337 );
nor \g448809/U$1 ( \23571 , \23568 , \23569 , \23570 );
and \g454870/U$2 ( \23572 , \16317 , RIe1a6a18_3273);
and \g454870/U$3 ( \23573 , RIe1a9718_3305, \16325 );
nor \g454870/U$1 ( \23574 , \23572 , \23573 );
not \g449837/U$3 ( \23575 , \23574 );
not \g449837/U$4 ( \23576 , \16311 );
and \g449837/U$2 ( \23577 , \23575 , \23576 );
and \g449837/U$5 ( \23578 , \16341 , RIe1d5bd8_3809);
nor \g449837/U$1 ( \23579 , \23577 , \23578 );
and \g451646/U$2 ( \23580 , \16377 , RIe1a1018_3209);
and \g451646/U$3 ( \23581 , RIe1a3d18_3241, \16313 );
nor \g451646/U$1 ( \23582 , \23580 , \23581 );
and \g451648/U$2 ( \23583 , \16334 , RIe21bf70_4608);
and \g451648/U$3 ( \23584 , RIe227370_4736, \16380 );
nor \g451648/U$1 ( \23585 , \23583 , \23584 );
nand \g447293/U$1 ( \23586 , \23571 , \23579 , \23582 , \23585 );
nor \g445946/U$1 ( \23587 , \23566 , \23567 , \23586 );
and \g451644/U$2 ( \23588 , \16364 , RIe1af550_3372);
and \g451644/U$3 ( \23589 , RIe1f16d0_4124, \16368 );
nor \g451644/U$1 ( \23590 , \23588 , \23589 );
nand \g445563/U$1 ( \23591 , \23565 , \23587 , \23590 );
and \g444888/U$2 ( \23592 , \23591 , \16752 );
and \g448806/U$2 ( \23593 , RIfcdfd78_7569, \16427 );
and \g448806/U$3 ( \23594 , \16448 , RIfc90bd8_6669);
and \g448806/U$4 ( \23595 , RIf149e10_5300, \16485 );
nor \g448806/U$1 ( \23596 , \23593 , \23594 , \23595 );
and \g454619/U$2 ( \23597 , \16317 , RIfcc7520_7290);
and \g454619/U$3 ( \23598 , RIfc973e8_6743, \16325 );
nor \g454619/U$1 ( \23599 , \23597 , \23598 );
not \g454618/U$1 ( \23600 , \23599 );
and \g449835/U$2 ( \23601 , \23600 , \16336 );
and \g449835/U$3 ( \23602 , RIfcd6f70_7468, \16354 );
nor \g449835/U$1 ( \23603 , \23601 , \23602 );
and \g451642/U$2 ( \23604 , \16361 , RIe1ab608_3327);
and \g451642/U$3 ( \23605 , RIe1acdf0_3344, \16364 );
nor \g451642/U$1 ( \23606 , \23604 , \23605 );
and \g451641/U$2 ( \23607 , \16368 , RIe1b15a8_3395);
and \g451641/U$3 ( \23608 , RIe1b2ef8_3413, \16371 );
nor \g451641/U$1 ( \23609 , \23607 , \23608 );
nand \g448047/U$1 ( \23610 , \23596 , \23603 , \23606 , \23609 );
and \g444888/U$3 ( \23611 , \16477 , \23610 );
nor \g444888/U$1 ( \23612 , \23592 , \23611 );
and \g446729/U$2 ( \23613 , \18268 , RIfce3cc0_7614);
and \g446729/U$3 ( \23614 , RIfcc73b8_7289, \18270 );
nor \g446729/U$1 ( \23615 , \23613 , \23614 );
and \g446730/U$2 ( \23616 , \18273 , RIe1b7c50_3468);
and \g446730/U$3 ( \23617 , RIe1b9e10_3492, \18275 );
nor \g446730/U$1 ( \23618 , \23616 , \23617 );
and \g446731/U$2 ( \23619 , \18278 , RIfea0200_8166);
and \g446731/U$3 ( \23620 , RIe1b5a90_3444, \18280 );
nor \g446731/U$1 ( \23621 , \23619 , \23620 );
nand \g444586/U$1 ( \23622 , \23612 , \23615 , \23618 , \23621 );
and \g451635/U$2 ( \23623 , \16377 , RIe198918_3113);
and \g451635/U$3 ( \23624 , RIe192f18_3049, \16380 );
nor \g451635/U$1 ( \23625 , \23623 , \23624 );
and \g445943/U$2 ( \23626 , RIe19b618_3145, \16321 );
and \g445943/U$3 ( \23627 , RIfc8f3f0_6652, \16313 );
and \g448805/U$2 ( \23628 , RIe187b18_2921, \16427 );
and \g448805/U$3 ( \23629 , \16432 , RIe18a818_2953);
and \g448805/U$4 ( \23630 , RIe195c18_3081, \16344 );
nor \g448805/U$1 ( \23631 , \23628 , \23629 , \23630 );
and \g454617/U$2 ( \23632 , \16317 , RIe182118_2857);
and \g454617/U$3 ( \23633 , RIfcb3cf0_7068, \16325 );
nor \g454617/U$1 ( \23634 , \23632 , \23633 );
not \g454616/U$1 ( \23635 , \23634 );
and \g449833/U$2 ( \23636 , \23635 , \16336 );
and \g449833/U$3 ( \23637 , RIf144b18_5241, \16354 );
nor \g449833/U$1 ( \23638 , \23636 , \23637 );
and \g452863/U$2 ( \23639 , \16361 , RIe17c718_2793);
and \g452863/U$3 ( \23640 , RIe17f418_2825, \16364 );
nor \g452863/U$1 ( \23641 , \23639 , \23640 );
and \g451636/U$2 ( \23642 , \16368 , RIe184e18_2889);
and \g451636/U$3 ( \23643 , RIf143d08_5231, \16371 );
nor \g451636/U$1 ( \23644 , \23642 , \23643 );
nand \g448046/U$1 ( \23645 , \23631 , \23638 , \23641 , \23644 );
nor \g445943/U$1 ( \23646 , \23626 , \23627 , \23645 );
and \g451634/U$2 ( \23647 , \16334 , RIe190218_3017);
and \g451634/U$3 ( \23648 , RIe19e318_3177, \16326 );
nor \g451634/U$1 ( \23649 , \23647 , \23648 );
nand \g445562/U$1 ( \23650 , \23625 , \23646 , \23649 );
and \g444732/U$2 ( \23651 , \23650 , \17938 );
and \g448803/U$2 ( \23652 , RIfc97820_6746, \16319 );
and \g448803/U$3 ( \23653 , \16328 , RIfc8fc60_6658);
and \g448803/U$4 ( \23654 , RIf15bb88_5503, \16398 );
nor \g448803/U$1 ( \23655 , \23652 , \23653 , \23654 );
and \g454905/U$2 ( \23656 , \16317 , RIfcdfee0_7570);
and \g454905/U$3 ( \23657 , RIfcc27c8_7235, \16325 );
nor \g454905/U$1 ( \23658 , \23656 , \23657 );
not \g449830/U$3 ( \23659 , \23658 );
not \g449830/U$4 ( \23660 , \16330 );
and \g449830/U$2 ( \23661 , \23659 , \23660 );
and \g449830/U$5 ( \23662 , \16341 , RIfc7be90_6432);
nor \g449830/U$1 ( \23663 , \23661 , \23662 );
and \g453028/U$2 ( \23664 , \16377 , RIe201288_4303);
and \g453028/U$3 ( \23665 , RIe202ea8_4323, \16313 );
nor \g453028/U$1 ( \23666 , \23664 , \23665 );
and \g451633/U$2 ( \23667 , \16334 , RIfc58670_6028);
and \g451633/U$3 ( \23668 , RIfc44198_5797, \16380 );
nor \g451633/U$1 ( \23669 , \23667 , \23668 );
nand \g447291/U$1 ( \23670 , \23655 , \23663 , \23666 , \23669 );
and \g444732/U$3 ( \23671 , \16394 , \23670 );
nor \g444732/U$1 ( \23672 , \23651 , \23671 );
and \g446728/U$2 ( \23673 , \16419 , RIfcd8e60_7490);
and \g446728/U$3 ( \23674 , RIfcd8cf8_7489, \16422 );
nor \g446728/U$1 ( \23675 , \23673 , \23674 );
and \g446725/U$2 ( \23676 , \16429 , RIf15e9f0_5536);
and \g446725/U$3 ( \23677 , RIf1608e0_5558, \16434 );
nor \g446725/U$1 ( \23678 , \23676 , \23677 );
and \g446726/U$2 ( \23679 , \16438 , RIe1fc0f8_4245);
and \g446726/U$3 ( \23680 , RIfe9ff30_8164, \16441 );
nor \g446726/U$1 ( \23681 , \23679 , \23680 );
nand \g444477/U$1 ( \23682 , \23672 , \23675 , \23678 , \23681 );
and \g445940/U$2 ( \23683 , RIf16cdc0_5698, \16328 );
and \g445940/U$3 ( \23684 , RIe221970_4672, \16377 );
and \g448800/U$2 ( \23685 , RIe213870_4512, \16427 );
and \g448800/U$3 ( \23686 , \16448 , RIfc3ff08_5753);
and \g448800/U$4 ( \23687 , RIe21ec70_4640, \16485 );
nor \g448800/U$1 ( \23688 , \23685 , \23686 , \23687 );
and \g455268/U$2 ( \23689 , \16317 , RIe20de70_4448);
and \g455268/U$3 ( \23690 , RIfc58940_6030, \16325 );
nor \g455268/U$1 ( \23691 , \23689 , \23690 );
not \g455267/U$1 ( \23692 , \23691 );
and \g449827/U$2 ( \23693 , \23692 , \16336 );
and \g449827/U$3 ( \23694 , RIfc58508_6027, \16356 );
nor \g449827/U$1 ( \23695 , \23693 , \23694 );
and \g451621/U$2 ( \23696 , \16361 , RIe208470_4384);
and \g451621/U$3 ( \23697 , RIe20b170_4416, \16364 );
nor \g451621/U$1 ( \23698 , \23696 , \23697 );
and \g453341/U$2 ( \23699 , \16368 , RIe210b70_4480);
and \g453341/U$3 ( \23700 , RIf1696e8_5659, \16371 );
nor \g453341/U$1 ( \23701 , \23699 , \23700 );
nand \g448045/U$1 ( \23702 , \23688 , \23695 , \23698 , \23701 );
nor \g445940/U$1 ( \23703 , \23683 , \23684 , \23702 );
and \g451620/U$2 ( \23704 , \16334 , RIe216570_4544);
and \g451620/U$3 ( \23705 , RIf16c118_5689, \16313 );
nor \g451620/U$1 ( \23706 , \23704 , \23705 );
and \g451619/U$2 ( \23707 , \16380 , RIe219270_4576);
and \g451619/U$3 ( \23708 , RIe224670_4704, \16321 );
nor \g451619/U$1 ( \23709 , \23707 , \23708 );
and \g445105/U$2 ( \23710 , \23703 , \23706 , \23709 );
nor \g445105/U$1 ( \23711 , \23710 , \16389 );
and \g445942/U$2 ( \23712 , RIfc8f6c0_6654, \16448 );
and \g445942/U$3 ( \23713 , RIfc583a0_6026, \16361 );
and \g448802/U$2 ( \23714 , RIf13f550_5180, \16485 );
and \g448802/U$3 ( \23715 , \16356 , RIfc57e00_6022);
and \g448802/U$4 ( \23716 , RIfc8f990_6656, \16337 );
nor \g448802/U$1 ( \23717 , \23714 , \23715 , \23716 );
and \g454610/U$2 ( \23718 , \16317 , RIf141170_5200);
and \g454610/U$3 ( \23719 , RIfc448a0_5802, \16325 );
nor \g454610/U$1 ( \23720 , \23718 , \23719 );
not \g449828/U$3 ( \23721 , \23720 );
not \g449828/U$4 ( \23722 , \16311 );
and \g449828/U$2 ( \23723 , \23721 , \23722 );
and \g449828/U$5 ( \23724 , \16341 , RIfc7c700_6438);
nor \g449828/U$1 ( \23725 , \23723 , \23724 );
and \g451627/U$2 ( \23726 , \16377 , RIfea0098_8165);
and \g451627/U$3 ( \23727 , RIfc7c9d0_6440, \16313 );
nor \g451627/U$1 ( \23728 , \23726 , \23727 );
and \g451628/U$2 ( \23729 , \16334 , RIee3d900_5159);
and \g451628/U$3 ( \23730 , RIfcd6e08_7467, \16380 );
nor \g451628/U$1 ( \23731 , \23729 , \23730 );
nand \g447290/U$1 ( \23732 , \23717 , \23725 , \23728 , \23731 );
nor \g445942/U$1 ( \23733 , \23712 , \23713 , \23732 );
and \g451625/U$2 ( \23734 , \16364 , RIfce9828_7679);
and \g451625/U$3 ( \23735 , RIe1742e8_2699, \16368 );
nor \g451625/U$1 ( \23736 , \23734 , \23735 );
and \g451624/U$2 ( \23737 , \16371 , RIfca27e8_6871);
and \g451624/U$3 ( \23738 , RIfce0048_7571, \16427 );
nor \g451624/U$1 ( \23739 , \23737 , \23738 );
and \g445108/U$2 ( \23740 , \23733 , \23736 , \23739 );
nor \g445108/U$1 ( \23741 , \23740 , \16649 );
or \g444342/U$1 ( \23742 , \23622 , \23682 , \23711 , \23741 );
and \g445935/U$2 ( \23743 , RIfca2d88_6875, \16328 );
and \g445935/U$3 ( \23744 , RIe1f6158_4177, \16334 );
and \g448797/U$2 ( \23745 , RIfc907a0_6666, \16337 );
and \g448797/U$3 ( \23746 , \16341 , RIfc59048_6035);
and \g448797/U$4 ( \23747 , RIfc90200_6662, \16485 );
nor \g448797/U$1 ( \23748 , \23745 , \23746 , \23747 );
and \g455147/U$2 ( \23749 , \16317 , RIfca2ef0_6876);
and \g455147/U$3 ( \23750 , RIfc904d0_6664, \16325 );
nor \g455147/U$1 ( \23751 , \23749 , \23750 );
not \g449824/U$3 ( \23752 , \23751 );
not \g449824/U$4 ( \23753 , \16351 );
and \g449824/U$2 ( \23754 , \23752 , \23753 );
and \g449824/U$5 ( \23755 , \16356 , RIfc90098_6661);
nor \g449824/U$1 ( \23756 , \23754 , \23755 );
and \g451610/U$2 ( \23757 , \16361 , RIe1eeb38_4093);
and \g451610/U$3 ( \23758 , RIfc90638_6665, \16364 );
nor \g451610/U$1 ( \23759 , \23757 , \23758 );
and \g451609/U$2 ( \23760 , \16368 , RIe1f3e30_4152);
and \g451609/U$3 ( \23761 , RIfc97550_6744, \16371 );
nor \g451609/U$1 ( \23762 , \23760 , \23761 );
nand \g447624/U$1 ( \23763 , \23748 , \23756 , \23759 , \23762 );
nor \g445935/U$1 ( \23764 , \23743 , \23744 , \23763 );
and \g451606/U$2 ( \23765 , \16377 , RIe1fabe0_4230);
and \g451606/U$3 ( \23766 , RIfcd20b0_7412, \16380 );
nor \g451606/U$1 ( \23767 , \23765 , \23766 );
and \g453729/U$2 ( \23768 , \16313 , RIfcb3a20_7066);
and \g453729/U$3 ( \23769 , RIfcbdea8_7183, \16321 );
nor \g453729/U$1 ( \23770 , \23768 , \23769 );
and \g445103/U$2 ( \23771 , \23764 , \23767 , \23770 );
nor \g445103/U$1 ( \23772 , \23771 , \16480 );
and \g445939/U$2 ( \23773 , RIe1d2ed8_3777, \16448 );
and \g445939/U$3 ( \23774 , RIe1bf3d8_3553, \16361 );
and \g448798/U$2 ( \23775 , RIe1de2d8_3905, \16485 );
and \g448798/U$3 ( \23776 , \16356 , RIe1e0fd8_3937);
and \g448798/U$4 ( \23777 , RIe1c4dd8_3617, \16398 );
nor \g448798/U$1 ( \23778 , \23775 , \23776 , \23777 );
and \g455200/U$2 ( \23779 , \16317 , RIe1e96d8_4033);
and \g455200/U$3 ( \23780 , RIe1ec3d8_4065, \16325 );
nor \g455200/U$1 ( \23781 , \23779 , \23780 );
not \g449825/U$3 ( \23782 , \23781 );
not \g449825/U$4 ( \23783 , \16311 );
and \g449825/U$2 ( \23784 , \23782 , \23783 );
and \g449825/U$5 ( \23785 , \16341 , RIe1c7ad8_3649);
nor \g449825/U$1 ( \23786 , \23784 , \23785 );
and \g451615/U$2 ( \23787 , \16377 , RIe1e3cd8_3969);
and \g451615/U$3 ( \23788 , RIe1e69d8_4001, \16313 );
nor \g451615/U$1 ( \23789 , \23787 , \23788 );
and \g451616/U$2 ( \23790 , \16334 , RIe1d88d8_3841);
and \g451616/U$3 ( \23791 , RIe1db5d8_3873, \16380 );
nor \g451616/U$1 ( \23792 , \23790 , \23791 );
nand \g447289/U$1 ( \23793 , \23778 , \23786 , \23789 , \23792 );
nor \g445939/U$1 ( \23794 , \23773 , \23774 , \23793 );
and \g451614/U$2 ( \23795 , \16364 , RIe1c20d8_3585);
and \g451614/U$3 ( \23796 , RIe1ca7d8_3681, \16368 );
nor \g451614/U$1 ( \23797 , \23795 , \23796 );
and \g451612/U$2 ( \23798 , \16371 , RIe1cd4d8_3713);
and \g451612/U$3 ( \23799 , RIe1d01d8_3745, \16427 );
nor \g451612/U$1 ( \23800 , \23798 , \23799 );
and \g445104/U$2 ( \23801 , \23794 , \23797 , \23800 );
nor \g445104/U$1 ( \23802 , \23801 , \16555 );
or \g444258/U$1 ( \23803 , \23742 , \23772 , \23802 );
_DC \g4273/U$1 ( \23804 , \23803 , \16652 );
and \g450727/U$2 ( \23805 , \16364 , RIf16e170_5712);
and \g450727/U$3 ( \23806 , RIfcd7678_7473, \16398 );
nor \g450727/U$1 ( \23807 , \23805 , \23806 );
and \g445735/U$2 ( \23808 , RIfcd7948_7475, \16341 );
and \g445735/U$3 ( \23809 , RIe175968_2715, \16377 );
and \g448559/U$2 ( \23810 , RIf140bd0_5196, \16321 );
and \g448559/U$3 ( \23811 , \16485 , RIf13efb0_5176);
and \g448559/U$4 ( \23812 , RIfc79b68_6407, \16356 );
nor \g448559/U$1 ( \23813 , \23810 , \23811 , \23812 );
and \g450757/U$2 ( \23814 , \16368 , RIe1734d8_2689);
and \g450757/U$3 ( \23815 , RIfc79898_6405, \16371 );
nor \g450757/U$1 ( \23816 , \23814 , \23815 );
and \g454615/U$2 ( \23817 , \16317 , RIfcea200_7686);
and \g454615/U$3 ( \23818 , RIfcd8320_7482, \16325 );
nor \g454615/U$1 ( \23819 , \23817 , \23818 );
not \g449580/U$3 ( \23820 , \23819 );
not \g449580/U$4 ( \23821 , \16351 );
and \g449580/U$2 ( \23822 , \23820 , \23821 );
and \g449580/U$5 ( \23823 , \16326 , RIf142250_5212);
nor \g449580/U$1 ( \23824 , \23822 , \23823 );
and \g450743/U$2 ( \23825 , \16334 , RIfcb2aa8_7055);
and \g450743/U$3 ( \23826 , RIfc92528_6687, \16380 );
nor \g450743/U$1 ( \23827 , \23825 , \23826 );
nand \g447481/U$1 ( \23828 , \23813 , \23816 , \23824 , \23827 );
nor \g445735/U$1 ( \23829 , \23808 , \23809 , \23828 );
and \g450706/U$2 ( \23830 , \16361 , RIfc927f8_6689);
and \g450706/U$3 ( \23831 , RIfec43f8_8353, \16313 );
nor \g450706/U$1 ( \23832 , \23830 , \23831 );
nand \g445512/U$1 ( \23833 , \23807 , \23829 , \23832 );
and \g444699/U$2 ( \23834 , \23833 , \17998 );
and \g448523/U$2 ( \23835 , RIe186ba0_2910, \16427 );
and \g448523/U$3 ( \23836 , \16448 , RIe1898a0_2942);
and \g448523/U$4 ( \23837 , RIe19a6a0_3134, \16321 );
nor \g448523/U$1 ( \23838 , \23835 , \23836 , \23837 );
and \g450634/U$2 ( \23839 , \16368 , RIe183ea0_2878);
and \g450634/U$3 ( \23840 , RIfc422a8_5775, \16371 );
nor \g450634/U$1 ( \23841 , \23839 , \23840 );
and \g454202/U$2 ( \23842 , \16317 , RIe194ca0_3070);
and \g454202/U$3 ( \23843 , RIfc923c0_6686, \16325 );
nor \g454202/U$1 ( \23844 , \23842 , \23843 );
not \g449540/U$3 ( \23845 , \23844 );
not \g449540/U$4 ( \23846 , \16330 );
and \g449540/U$2 ( \23847 , \23845 , \23846 );
and \g449540/U$5 ( \23848 , \16328 , RIe19d3a0_3166);
nor \g449540/U$1 ( \23849 , \23847 , \23848 );
and \g450614/U$2 ( \23850 , \16334 , RIe18f2a0_3006);
and \g450614/U$3 ( \23851 , RIe191fa0_3038, \16380 );
nor \g450614/U$1 ( \23852 , \23850 , \23851 );
nand \g447465/U$1 ( \23853 , \23838 , \23841 , \23849 , \23852 );
and \g444699/U$3 ( \23854 , \17938 , \23853 );
nor \g444699/U$1 ( \23855 , \23834 , \23854 );
and \g446504/U$2 ( \23856 , \18776 , RIe1979a0_3102);
and \g446504/U$3 ( \23857 , RIfcb2c10_7056, \18778 );
nor \g446504/U$1 ( \23858 , \23856 , \23857 );
and \g446513/U$2 ( \23859 , \18781 , RIe1811a0_2846);
and \g446513/U$3 ( \23860 , RIfcbecb8_7193, \18783 );
nor \g446513/U$1 ( \23861 , \23859 , \23860 );
and \g446514/U$2 ( \23862 , \18467 , RIe17b7a0_2782);
and \g446514/U$3 ( \23863 , RIe17e4a0_2814, \18469 );
nor \g446514/U$1 ( \23864 , \23862 , \23863 );
nand \g444449/U$1 ( \23865 , \23855 , \23858 , \23861 , \23864 );
and \g447176/U$2 ( \23866 , \19215 , RIe1c9860_3670);
and \g447176/U$3 ( \23867 , RIe1cc560_3702, \19210 );
nor \g447176/U$1 ( \23868 , \23866 , \23867 );
and \g446447/U$2 ( \23869 , RIe1e0060_3926, \16356 );
and \g446447/U$3 ( \23870 , RIe1dd360_3894, \16485 );
and \g449471/U$2 ( \23871 , RIe1cf260_3734, \16427 );
and \g449471/U$3 ( \23872 , \16337 , RIe1c3e60_3606);
and \g449471/U$4 ( \23873 , RIe1c6b60_3638, \16341 );
nor \g449471/U$1 ( \23874 , \23871 , \23872 , \23873 );
and \g453929/U$2 ( \23875 , \16361 , RIe1be460_3542);
and \g453929/U$3 ( \23876 , RIe1c1160_3574, \16364 );
nor \g453929/U$1 ( \23877 , \23875 , \23876 );
and \g453925/U$2 ( \23878 , \16377 , RIe1e2d60_3958);
and \g453925/U$3 ( \23879 , RIe1e5a60_3990, \16313 );
nor \g453925/U$1 ( \23880 , \23878 , \23879 );
and \g454285/U$2 ( \23881 , \16317 , RIe1e8760_4022);
and \g454285/U$3 ( \23882 , RIe1eb460_4054, \16325 );
nor \g454285/U$1 ( \23883 , \23881 , \23882 );
not \g450488/U$3 ( \23884 , \23883 );
not \g450488/U$4 ( \23885 , \16311 );
and \g450488/U$2 ( \23886 , \23884 , \23885 );
and \g450488/U$5 ( \23887 , \16448 , RIe1d1f60_3766);
nor \g450488/U$1 ( \23888 , \23886 , \23887 );
nand \g447979/U$1 ( \23889 , \23874 , \23877 , \23880 , \23888 );
nor \g446447/U$1 ( \23890 , \23869 , \23870 , \23889 );
not \g444897/U$3 ( \23891 , \23890 );
not \g444897/U$4 ( \23892 , \16555 );
and \g444897/U$2 ( \23893 , \23891 , \23892 );
and \g446475/U$2 ( \23894 , RIe18c5a0_2974, \16354 );
and \g446475/U$3 ( \23895 , RIe1f0758_4113, \16368 );
and \g449509/U$2 ( \23896 , RIe1a5aa0_3262, \16321 );
and \g449509/U$3 ( \23897 , \16326 , RIe1a87a0_3294);
and \g449509/U$4 ( \23898 , RIe1fe858_4273, \16427 );
nor \g449509/U$1 ( \23899 , \23896 , \23897 , \23898 );
and \g454083/U$2 ( \23900 , \16361 , RIe170c10_2660);
and \g454083/U$3 ( \23901 , RIe1ae5d8_3361, \16364 );
nor \g454083/U$1 ( \23902 , \23900 , \23901 );
and \g454065/U$2 ( \23903 , \16377 , RIe1a00a0_3198);
and \g454065/U$3 ( \23904 , RIe1a2da0_3230, \16313 );
nor \g454065/U$1 ( \23905 , \23903 , \23904 );
and \g454963/U$2 ( \23906 , \16317 , RIe1bb760_3510);
and \g454963/U$3 ( \23907 , RIe1d4c60_3798, \16325 );
nor \g454963/U$1 ( \23908 , \23906 , \23907 );
not \g454962/U$1 ( \23909 , \23908 );
and \g450525/U$2 ( \23910 , \23909 , \16336 );
and \g450525/U$3 ( \23911 , RIe2047f8_4341, \16448 );
nor \g450525/U$1 ( \23912 , \23910 , \23911 );
nand \g448127/U$1 ( \23913 , \23899 , \23902 , \23905 , \23912 );
nor \g446475/U$1 ( \23914 , \23894 , \23895 , \23913 );
and \g454023/U$2 ( \23915 , \16334 , RIe21aff8_4597);
and \g454023/U$3 ( \23916 , RIe1f7c10_4196, \16371 );
nor \g454023/U$1 ( \23917 , \23915 , \23916 );
and \g454012/U$2 ( \23918 , \16380 , RIe2263f8_4725);
and \g454012/U$3 ( \23919 , RIe178aa0_2750, \16344 );
nor \g454012/U$1 ( \23920 , \23918 , \23919 );
and \g445482/U$2 ( \23921 , \23914 , \23917 , \23920 );
nor \g445482/U$1 ( \23922 , \23921 , \16586 );
nor \g444897/U$1 ( \23923 , \23893 , \23922 );
and \g447188/U$2 ( \23924 , \19462 , RIe1d7960_3830);
and \g447188/U$3 ( \23925 , RIe1da660_3862, \19464 );
nor \g447188/U$1 ( \23926 , \23924 , \23925 );
nand \g444437/U$1 ( \23927 , \23868 , \23923 , \23926 );
and \g446388/U$2 ( \23928 , RIfc79028_6399, \16339 );
and \g446388/U$3 ( \23929 , RIe2008b0_4296, \16377 );
and \g449392/U$2 ( \23930 , RIf166010_5620, \16319 );
and \g449392/U$3 ( \23931 , \16344 , RIfc41ba0_5770);
and \g449392/U$4 ( \23932 , RIf165098_5609, \16356 );
nor \g449392/U$1 ( \23933 , \23930 , \23931 , \23932 );
and \g453647/U$2 ( \23934 , \16368 , RIfec4560_8354);
and \g453647/U$3 ( \23935 , RIe1fcad0_4252, \16371 );
nor \g453647/U$1 ( \23936 , \23934 , \23935 );
and \g454977/U$2 ( \23937 , \16317 , RIfc79190_6400);
and \g454977/U$3 ( \23938 , RIfc418d0_5768, \16325 );
nor \g454977/U$1 ( \23939 , \23937 , \23938 );
not \g450406/U$3 ( \23940 , \23939 );
not \g450406/U$4 ( \23941 , \16351 );
and \g450406/U$2 ( \23942 , \23940 , \23941 );
and \g450406/U$5 ( \23943 , \16328 , RIfcd7510_7472);
nor \g450406/U$1 ( \23944 , \23942 , \23943 );
and \g453637/U$2 ( \23945 , \16334 , RIfc92c30_6692);
and \g453637/U$3 ( \23946 , RIfc41a38_5769, \16380 );
nor \g453637/U$1 ( \23947 , \23945 , \23946 );
nand \g447934/U$1 ( \23948 , \23933 , \23936 , \23944 , \23947 );
nor \g446388/U$1 ( \23949 , \23928 , \23929 , \23948 );
and \g453589/U$2 ( \23950 , \16361 , RIfcd81b8_7481);
and \g453589/U$3 ( \23951 , RIfe9d230_8132, \16313 );
nor \g453589/U$1 ( \23952 , \23950 , \23951 );
and \g453603/U$2 ( \23953 , \16364 , RIfcc1df0_7228);
and \g453603/U$3 ( \23954 , RIfcbf258_7197, \16398 );
nor \g453603/U$1 ( \23955 , \23953 , \23954 );
and \g445413/U$2 ( \23956 , \23949 , \23952 , \23955 );
nor \g445413/U$1 ( \23957 , \23956 , \16393 );
and \g446408/U$2 ( \23958 , RIf16ad68_5675, \16356 );
and \g446408/U$3 ( \23959 , RIe20fbf8_4469, \16368 );
and \g449428/U$2 ( \23960 , RIe2128f8_4501, \16427 );
and \g449428/U$3 ( \23961 , \16337 , RIe20cef8_4437);
and \g449428/U$4 ( \23962 , RIfc41d08_5771, \16339 );
nor \g449428/U$1 ( \23963 , \23960 , \23961 , \23962 );
and \g453779/U$2 ( \23964 , \16361 , RIe2074f8_4373);
and \g453779/U$3 ( \23965 , RIe20a1f8_4405, \16364 );
nor \g453779/U$1 ( \23966 , \23964 , \23965 );
and \g453769/U$2 ( \23967 , \16377 , RIe2209f8_4661);
and \g453769/U$3 ( \23968 , RIfc795c8_6403, \16313 );
nor \g453769/U$1 ( \23969 , \23967 , \23968 );
and \g455081/U$2 ( \23970 , \16317 , RIe2236f8_4693);
and \g455081/U$3 ( \23971 , RIfc92960_6690, \16325 );
nor \g455081/U$1 ( \23972 , \23970 , \23971 );
not \g450446/U$3 ( \23973 , \23972 );
not \g450446/U$4 ( \23974 , \16311 );
and \g450446/U$2 ( \23975 , \23973 , \23974 );
and \g450446/U$5 ( \23976 , \16448 , RIfe9d398_8133);
nor \g450446/U$1 ( \23977 , \23975 , \23976 );
nand \g447955/U$1 ( \23978 , \23963 , \23966 , \23969 , \23977 );
nor \g446408/U$1 ( \23979 , \23958 , \23959 , \23978 );
and \g453727/U$2 ( \23980 , \16334 , RIe2155f8_4533);
and \g453727/U$3 ( \23981 , RIfcdb9f8_7521, \16371 );
nor \g453727/U$1 ( \23982 , \23980 , \23981 );
and \g453720/U$2 ( \23983 , \16380 , RIe2182f8_4565);
and \g453720/U$3 ( \23984 , RIe21dcf8_4629, \16344 );
nor \g453720/U$1 ( \23985 , \23983 , \23984 );
and \g445433/U$2 ( \23986 , \23979 , \23982 , \23985 );
nor \g445433/U$1 ( \23987 , \23986 , \16389 );
or \g444299/U$1 ( \23988 , \23865 , \23927 , \23957 , \23987 );
and \g446325/U$2 ( \23989 , RIfce3180_7606, \16339 );
and \g446325/U$3 ( \23990 , RIe1fa0a0_4222, \16377 );
and \g449319/U$2 ( \23991 , RIfec46c8_8355, \16427 );
and \g449319/U$3 ( \23992 , \16448 , RIfec4830_8356);
and \g449319/U$4 ( \23993 , RIfc5b4d8_6061, \16321 );
nor \g449319/U$1 ( \23994 , \23991 , \23992 , \23993 );
and \g453365/U$2 ( \23995 , \16368 , RIe1f3020_4142);
and \g453365/U$3 ( \23996 , RIf1508f0_5376, \16371 );
nor \g453365/U$1 ( \23997 , \23995 , \23996 );
and \g455225/U$2 ( \23998 , \16317 , RIfe9d500_8134);
and \g455225/U$3 ( \23999 , RIf156188_5439, \16325 );
nor \g455225/U$1 ( \24000 , \23998 , \23999 );
not \g450327/U$3 ( \24001 , \24000 );
not \g450327/U$4 ( \24002 , \16330 );
and \g450327/U$2 ( \24003 , \24001 , \24002 );
and \g450327/U$5 ( \24004 , \16328 , RIfc92d98_6693);
nor \g450327/U$1 ( \24005 , \24003 , \24004 );
and \g453351/U$2 ( \24006 , \16334 , RIe1f5348_4167);
and \g453351/U$3 ( \24007 , RIf1546d0_5420, \16380 );
nor \g453351/U$1 ( \24008 , \24006 , \24007 );
nand \g447884/U$1 ( \24009 , \23994 , \23997 , \24005 , \24008 );
nor \g446325/U$1 ( \24010 , \23989 , \23990 , \24009 );
and \g453299/U$2 ( \24011 , \16361 , RIe1edd28_4083);
and \g453299/U$3 ( \24012 , RIfcd77e0_7474, \16313 );
nor \g453299/U$1 ( \24013 , \24011 , \24012 );
and \g453317/U$2 ( \24014 , \16364 , RIfcbf690_7200);
and \g453317/U$3 ( \24015 , RIfce8fb8_7673, \16398 );
nor \g453317/U$1 ( \24016 , \24014 , \24015 );
and \g445371/U$2 ( \24017 , \24010 , \24013 , \24016 );
nor \g445371/U$1 ( \24018 , \24017 , \16480 );
and \g446355/U$2 ( \24019 , RIf147110_5268, \16341 );
and \g446355/U$3 ( \24020 , RIe1b7110_3460, \16377 );
and \g449358/U$2 ( \24021 , RIfe9cc90_8128, \16319 );
and \g449358/U$3 ( \24022 , \16485 , RIfe9cb28_8127);
and \g449358/U$4 ( \24023 , RIf14a3b0_5304, \16356 );
nor \g449358/U$1 ( \24024 , \24021 , \24022 , \24023 );
and \g453506/U$2 ( \24025 , \16368 , RIfe9cdf8_8129);
and \g453506/U$3 ( \24026 , RIfe9c858_8125, \16371 );
nor \g453506/U$1 ( \24027 , \24025 , \24026 );
and \g454736/U$2 ( \24028 , \16317 , RIfce9558_7677);
and \g454736/U$3 ( \24029 , RIfce2208_7595, \16325 );
nor \g454736/U$1 ( \24030 , \24028 , \24029 );
not \g450371/U$3 ( \24031 , \24030 );
not \g450371/U$4 ( \24032 , \16351 );
and \g450371/U$2 ( \24033 , \24031 , \24032 );
and \g450371/U$5 ( \24034 , \16328 , RIfe9d0c8_8131);
nor \g450371/U$1 ( \24035 , \24033 , \24034 );
and \g453490/U$2 ( \24036 , \16334 , RIfe9c9c0_8126);
and \g453490/U$3 ( \24037 , RIfe9cf60_8130, \16380 );
nor \g453490/U$1 ( \24038 , \24036 , \24037 );
nand \g447907/U$1 ( \24039 , \24024 , \24027 , \24035 , \24038 );
nor \g446355/U$1 ( \24040 , \24019 , \24020 , \24039 );
and \g453440/U$2 ( \24041 , \16361 , RIe1aaac8_3319);
and \g453440/U$3 ( \24042 , RIe1b9168_3483, \16313 );
nor \g453440/U$1 ( \24043 , \24041 , \24042 );
and \g453470/U$2 ( \24044 , \16364 , RIe1ac2b0_3336);
and \g453470/U$3 ( \24045 , RIf146468_5259, \16337 );
nor \g453470/U$1 ( \24046 , \24044 , \24045 );
and \g445397/U$2 ( \24047 , \24040 , \24043 , \24046 );
nor \g445397/U$1 ( \24048 , \24047 , \16909 );
or \g444161/U$1 ( \24049 , \23988 , \24018 , \24048 );
_DC \g42f8/U$1 ( \24050 , \24049 , \16652 );
and \g447103/U$2 ( \24051 , \18030 , RIe214680_4522);
and \g447103/U$3 ( \24052 , RIe217380_4554, \18032 );
nor \g447103/U$1 ( \24053 , \24051 , \24052 );
and \g446335/U$2 ( \24054 , RIfcd0b98_7397, \16354 );
and \g446335/U$3 ( \24055 , RIe21cd80_4618, \16485 );
and \g449316/U$2 ( \24056 , RIe222780_4682, \16319 );
and \g449316/U$3 ( \24057 , \16328 , RIfc40340_5756);
and \g449316/U$4 ( \24058 , RIe211980_4490, \16427 );
nor \g449316/U$1 ( \24059 , \24056 , \24057 , \24058 );
and \g453397/U$2 ( \24060 , \16361 , RIe206580_4362);
and \g453397/U$3 ( \24061 , RIe209280_4394, \16364 );
nor \g453397/U$1 ( \24062 , \24060 , \24061 );
and \g453391/U$2 ( \24063 , \16377 , RIe21fa80_4650);
and \g453391/U$3 ( \24064 , RIfcdd618_7541, \16313 );
nor \g453391/U$1 ( \24065 , \24063 , \24064 );
and \g455329/U$2 ( \24066 , \16317 , RIe20bf80_4426);
and \g455329/U$3 ( \24067 , RIfcc0770_7212, \16325 );
nor \g455329/U$1 ( \24068 , \24066 , \24067 );
not \g455328/U$1 ( \24069 , \24068 );
and \g450334/U$2 ( \24070 , \24069 , \16336 );
and \g450334/U$3 ( \24071 , RIfec4998_8357, \16432 );
nor \g450334/U$1 ( \24072 , \24070 , \24071 );
nand \g448109/U$1 ( \24073 , \24059 , \24062 , \24065 , \24072 );
nor \g446335/U$1 ( \24074 , \24054 , \24055 , \24073 );
not \g444820/U$3 ( \24075 , \24074 );
not \g444820/U$4 ( \24076 , \16389 );
and \g444820/U$2 ( \24077 , \24075 , \24076 );
and \g446344/U$2 ( \24078 , RIfec4c68_8359, \16313 );
and \g446344/U$3 ( \24079 , RIfccc3e0_7346, \16361 );
and \g449327/U$2 ( \24080 , RIfcc08d8_7213, \16427 );
and \g449327/U$3 ( \24081 , \16448 , RIfccd088_7355);
and \g449327/U$4 ( \24082 , RIfcee580_7734, \16321 );
nor \g449327/U$1 ( \24083 , \24080 , \24081 , \24082 );
and \g453436/U$2 ( \24084 , \16368 , RIfe9e1a8_8143);
and \g453436/U$3 ( \24085 , RIfe9e040_8142, \16371 );
nor \g453436/U$1 ( \24086 , \24084 , \24085 );
and \g455018/U$2 ( \24087 , \16317 , RIfcebcb8_7705);
and \g455018/U$3 ( \24088 , RIfc949b8_6713, \16325 );
nor \g455018/U$1 ( \24089 , \24087 , \24088 );
not \g450344/U$3 ( \24090 , \24089 );
not \g450344/U$4 ( \24091 , \16330 );
and \g450344/U$2 ( \24092 , \24090 , \24091 );
and \g450344/U$5 ( \24093 , \16326 , RIfce2370_7596);
nor \g450344/U$1 ( \24094 , \24092 , \24093 );
and \g453432/U$2 ( \24095 , \16334 , RIf1612b8_5565);
and \g453432/U$3 ( \24096 , RIf162938_5581, \16380 );
nor \g453432/U$1 ( \24097 , \24095 , \24096 );
nand \g447897/U$1 ( \24098 , \24083 , \24086 , \24094 , \24097 );
nor \g446344/U$1 ( \24099 , \24078 , \24079 , \24098 );
and \g453420/U$2 ( \24100 , \16364 , RIfc94c88_6715);
and \g453420/U$3 ( \24101 , RIfcead40_7694, \16341 );
nor \g453420/U$1 ( \24102 , \24100 , \24101 );
and \g453419/U$2 ( \24103 , \16398 , RIf15ad78_5493);
and \g453419/U$3 ( \24104 , RIfec4b00_8358, \16377 );
nor \g453419/U$1 ( \24105 , \24103 , \24104 );
and \g445389/U$2 ( \24106 , \24099 , \24102 , \24105 );
nor \g445389/U$1 ( \24107 , \24106 , \16393 );
nor \g444820/U$1 ( \24108 , \24077 , \24107 );
and \g447100/U$2 ( \24109 , \22457 , RIe20ec80_4458);
and \g447100/U$3 ( \24110 , RIf168608_5647, \22459 );
nor \g447100/U$1 ( \24111 , \24109 , \24110 );
nand \g444431/U$1 ( \24112 , \24053 , \24108 , \24111 );
and \g453494/U$2 ( \24113 , \16334 , RIe1b38d0_3420);
and \g453494/U$3 ( \24114 , RIe1b1f80_3402, \16371 );
nor \g453494/U$1 ( \24115 , \24113 , \24114 );
and \g446362/U$2 ( \24116 , RIfc76490_6368, \16485 );
and \g446362/U$3 ( \24117 , RIe1b4c80_3434, \16380 );
and \g449347/U$2 ( \24118 , RIf14ac20_5310, \16321 );
and \g449347/U$3 ( \24119 , \16328 , RIf14bfd0_5324);
and \g449347/U$4 ( \24120 , RIfceaea8_7695, \16427 );
nor \g449347/U$1 ( \24121 , \24118 , \24119 , \24120 );
and \g453512/U$2 ( \24122 , \16361 , RIfe9dd70_8140);
and \g453512/U$3 ( \24123 , RIfe9e5e0_8146, \16364 );
nor \g453512/U$1 ( \24124 , \24122 , \24123 );
and \g453503/U$2 ( \24125 , \16377 , RIe1b65d0_3452);
and \g453503/U$3 ( \24126 , RIfe9ded8_8141, \16313 );
nor \g453503/U$1 ( \24127 , \24125 , \24126 );
and \g454898/U$2 ( \24128 , \16317 , RIf145ec8_5255);
and \g454898/U$3 ( \24129 , RIfcd0760_7394, \16325 );
nor \g454898/U$1 ( \24130 , \24128 , \24129 );
not \g454897/U$1 ( \24131 , \24130 );
and \g450367/U$2 ( \24132 , \24131 , \16336 );
and \g450367/U$3 ( \24133 , RIfcc0fe0_7218, \16448 );
nor \g450367/U$1 ( \24134 , \24132 , \24133 );
nand \g448113/U$1 ( \24135 , \24121 , \24124 , \24127 , \24134 );
nor \g446362/U$1 ( \24136 , \24116 , \24117 , \24135 );
and \g453491/U$2 ( \24137 , \16368 , RIe1b0360_3382);
and \g453491/U$3 ( \24138 , RIfcecd98_7717, \16356 );
nor \g453491/U$1 ( \24139 , \24137 , \24138 );
nand \g445669/U$1 ( \24140 , \24115 , \24136 , \24139 );
and \g444922/U$2 ( \24141 , \24140 , \16477 );
and \g449338/U$2 ( \24142 , RIfc94df0_6716, \16319 );
and \g449338/U$3 ( \24143 , \16328 , RIfc765f8_6369);
and \g449338/U$4 ( \24144 , RIf1512c8_5383, \16427 );
nor \g449338/U$1 ( \24145 , \24142 , \24143 , \24144 );
and \g453473/U$2 ( \24146 , \16361 , RIe1ed1e8_4075);
and \g453473/U$3 ( \24147 , RIfcc0e78_7217, \16364 );
nor \g453473/U$1 ( \24148 , \24146 , \24147 );
and \g453471/U$2 ( \24149 , \16377 , RIe1f9998_4217);
and \g453471/U$3 ( \24150 , RIfcc0a40_7214, \16313 );
nor \g453471/U$1 ( \24151 , \24149 , \24150 );
and \g454528/U$2 ( \24152 , \16317 , RIfc950c0_6718);
and \g454528/U$3 ( \24153 , RIfc761c0_6366, \16325 );
nor \g454528/U$1 ( \24154 , \24152 , \24153 );
not \g454527/U$1 ( \24155 , \24154 );
and \g450355/U$2 ( \24156 , \24155 , \16336 );
and \g450355/U$3 ( \24157 , RIf152510_5396, \16448 );
nor \g450355/U$1 ( \24158 , \24156 , \24157 );
nand \g448112/U$1 ( \24159 , \24145 , \24148 , \24151 , \24158 );
and \g444922/U$3 ( \24160 , \16481 , \24159 );
nor \g444922/U$1 ( \24161 , \24141 , \24160 );
and \g447115/U$2 ( \24162 , \16511 , RIe1f4970_4160);
and \g447115/U$3 ( \24163 , RIfceb2e0_7698, \16514 );
nor \g447115/U$1 ( \24164 , \24162 , \24163 );
nor \g448456/U$1 ( \24165 , \16480 , \16484 );
and \g447113/U$2 ( \24166 , \24165 , RIfce8748_7667);
nor \g448447/U$1 ( \24167 , \16480 , \16355 );
and \g447113/U$3 ( \24168 , RIfcc8d08_7307, \24167 );
nor \g447113/U$1 ( \24169 , \24166 , \24168 );
and \g447114/U$2 ( \24170 , \17279 , RIe1f24e0_4134);
and \g447114/U$3 ( \24171 , RIfcb0ff0_7036, \17281 );
nor \g447114/U$1 ( \24172 , \24170 , \24171 );
nand \g444653/U$1 ( \24173 , \24161 , \24164 , \24169 , \24172 );
and \g446320/U$2 ( \24174 , RIe1a1e28_3219, \16313 );
and \g446320/U$3 ( \24175 , RIe1ad660_3350, \16364 );
and \g449298/U$2 ( \24176 , RIe1a4b28_3251, \16321 );
and \g449298/U$3 ( \24177 , \16344 , RIe177b28_2739);
and \g449298/U$4 ( \24178 , RIe18b628_2963, \16354 );
nor \g449298/U$1 ( \24179 , \24176 , \24177 , \24178 );
and \g453329/U$2 ( \24180 , \16368 , RIe1ef7e0_4102);
and \g453329/U$3 ( \24181 , RIe1f6c98_4185, \16371 );
nor \g453329/U$1 ( \24182 , \24180 , \24181 );
and \g455246/U$2 ( \24183 , \16317 , RIe1fd8e0_4262);
and \g455246/U$3 ( \24184 , RIe203880_4330, \16325 );
nor \g455246/U$1 ( \24185 , \24183 , \24184 );
not \g450314/U$3 ( \24186 , \24185 );
not \g450314/U$4 ( \24187 , \16351 );
and \g450314/U$2 ( \24188 , \24186 , \24187 );
and \g450314/U$5 ( \24189 , \16328 , RIe1a7828_3283);
nor \g450314/U$1 ( \24190 , \24188 , \24189 );
and \g453327/U$2 ( \24191 , \16334 , RIe21a080_4586);
and \g453327/U$3 ( \24192 , RIe225480_4714, \16380 );
nor \g453327/U$1 ( \24193 , \24191 , \24192 );
nand \g447882/U$1 ( \24194 , \24179 , \24182 , \24190 , \24193 );
nor \g446320/U$1 ( \24195 , \24174 , \24175 , \24194 );
and \g453314/U$2 ( \24196 , \16341 , RIe1d3ce8_3787);
and \g453314/U$3 ( \24197 , RIe19f128_3187, \16377 );
nor \g453314/U$1 ( \24198 , \24196 , \24197 );
and \g453318/U$2 ( \24199 , \16361 , RIe16fc98_2649);
and \g453318/U$3 ( \24200 , RIe1ba7e8_3499, \16398 );
nor \g453318/U$1 ( \24201 , \24199 , \24200 );
and \g445377/U$2 ( \24202 , \24195 , \24198 , \24201 );
nor \g445377/U$1 ( \24203 , \24202 , \16586 );
and \g446327/U$2 ( \24204 , RIe1dc3e8_3883, \16485 );
and \g446327/U$3 ( \24205 , RIe1d96e8_3851, \16380 );
and \g449306/U$2 ( \24206 , RIe1ce2e8_3723, \16427 );
and \g449306/U$3 ( \24207 , \16337 , RIe1c2ee8_3595);
and \g449306/U$4 ( \24208 , RIe1c5be8_3627, \16341 );
nor \g449306/U$1 ( \24209 , \24206 , \24207 , \24208 );
and \g453360/U$2 ( \24210 , \16361 , RIe1bd4e8_3531);
and \g453360/U$3 ( \24211 , RIe1c01e8_3563, \16364 );
nor \g453360/U$1 ( \24212 , \24210 , \24211 );
and \g453358/U$2 ( \24213 , \16377 , RIe1e1de8_3947);
and \g453358/U$3 ( \24214 , RIe1e4ae8_3979, \16313 );
nor \g453358/U$1 ( \24215 , \24213 , \24214 );
and \g454270/U$2 ( \24216 , \16317 , RIe1e77e8_4011);
and \g454270/U$3 ( \24217 , RIe1ea4e8_4043, \16325 );
nor \g454270/U$1 ( \24218 , \24216 , \24217 );
not \g450322/U$3 ( \24219 , \24218 );
not \g450322/U$4 ( \24220 , \16311 );
and \g450322/U$2 ( \24221 , \24219 , \24220 );
and \g450322/U$5 ( \24222 , \16448 , RIe1d0fe8_3755);
nor \g450322/U$1 ( \24223 , \24221 , \24222 );
nand \g447886/U$1 ( \24224 , \24209 , \24212 , \24215 , \24223 );
nor \g446327/U$1 ( \24225 , \24204 , \24205 , \24224 );
and \g453343/U$2 ( \24226 , \16368 , RIe1c88e8_3659);
and \g453343/U$3 ( \24227 , RIe1df0e8_3915, \16356 );
nor \g453343/U$1 ( \24228 , \24226 , \24227 );
and \g453347/U$2 ( \24229 , \16334 , RIe1d69e8_3819);
and \g453347/U$3 ( \24230 , RIe1cb5e8_3691, \16371 );
nor \g453347/U$1 ( \24231 , \24229 , \24230 );
and \g445382/U$2 ( \24232 , \24225 , \24228 , \24231 );
nor \g445382/U$1 ( \24233 , \24232 , \16555 );
or \g444300/U$1 ( \24234 , \24112 , \24173 , \24203 , \24233 );
and \g446307/U$2 ( \24235 , RIfe9e478_8145, \16341 );
and \g446307/U$3 ( \24236 , RIe196a28_3091, \16377 );
and \g449282/U$2 ( \24237 , RIe199728_3123, \16321 );
and \g449282/U$3 ( \24238 , \16485 , RIe193d28_3059);
and \g449282/U$4 ( \24239 , RIfcc04a0_7210, \16356 );
nor \g449282/U$1 ( \24240 , \24237 , \24238 , \24239 );
and \g453265/U$2 ( \24241 , \16368 , RIe182f28_2867);
and \g453265/U$3 ( \24242 , RIfce1830_7588, \16371 );
nor \g453265/U$1 ( \24243 , \24241 , \24242 );
and \g455272/U$2 ( \24244 , \16317 , RIe185c28_2899);
and \g455272/U$3 ( \24245 , RIe188928_2931, \16325 );
nor \g455272/U$1 ( \24246 , \24244 , \24245 );
not \g450297/U$3 ( \24247 , \24246 );
not \g450297/U$4 ( \24248 , \16351 );
and \g450297/U$2 ( \24249 , \24247 , \24248 );
and \g450297/U$5 ( \24250 , \16328 , RIe19c428_3155);
nor \g450297/U$1 ( \24251 , \24249 , \24250 );
and \g453263/U$2 ( \24252 , \16334 , RIe18e328_2995);
and \g453263/U$3 ( \24253 , RIe191028_3027, \16380 );
nor \g453263/U$1 ( \24254 , \24252 , \24253 );
nand \g447872/U$1 ( \24255 , \24240 , \24243 , \24251 , \24254 );
nor \g446307/U$1 ( \24256 , \24235 , \24236 , \24255 );
and \g453251/U$2 ( \24257 , \16361 , RIe17a828_2771);
and \g453251/U$3 ( \24258 , RIfe9e310_8144, \16313 );
nor \g453251/U$1 ( \24259 , \24257 , \24258 );
and \g453254/U$2 ( \24260 , \16364 , RIe17d528_2803);
and \g453254/U$3 ( \24261 , RIe180228_2835, \16398 );
nor \g453254/U$1 ( \24262 , \24260 , \24261 );
and \g445367/U$2 ( \24263 , \24256 , \24259 , \24262 );
nor \g445367/U$1 ( \24264 , \24263 , \16618 );
and \g446312/U$2 ( \24265 , RIfc77408_6379, \16356 );
and \g446312/U$3 ( \24266 , RIe172998_2681, \16368 );
and \g449290/U$2 ( \24267 , RIfced338_7721, \16427 );
and \g449290/U$3 ( \24268 , \16398 , RIfcddff0_7548);
and \g449290/U$4 ( \24269 , RIfcdc268_7527, \16341 );
nor \g449290/U$1 ( \24270 , \24267 , \24268 , \24269 );
and \g453294/U$2 ( \24271 , \16361 , RIfce7230_7652);
and \g453294/U$3 ( \24272 , RIfcc0608_7211, \16364 );
nor \g453294/U$1 ( \24273 , \24271 , \24272 );
and \g453288/U$2 ( \24274 , \16377 , RIe174f90_2708);
and \g453288/U$3 ( \24275 , RIfc94418_6709, \16313 );
nor \g453288/U$1 ( \24276 , \24274 , \24275 );
and \g454391/U$2 ( \24277 , \16317 , RIfcb12c0_7038);
and \g454391/U$3 ( \24278 , RIf141878_5205, \16325 );
nor \g454391/U$1 ( \24279 , \24277 , \24278 );
not \g450305/U$3 ( \24280 , \24279 );
not \g450305/U$4 ( \24281 , \16311 );
and \g450305/U$2 ( \24282 , \24280 , \24281 );
and \g450305/U$5 ( \24283 , \16432 , RIfc946e8_6711);
nor \g450305/U$1 ( \24284 , \24282 , \24283 );
nand \g447878/U$1 ( \24285 , \24270 , \24273 , \24276 , \24284 );
nor \g446312/U$1 ( \24286 , \24265 , \24266 , \24285 );
and \g453281/U$2 ( \24287 , \16334 , RIfc94580_6710);
and \g453281/U$3 ( \24288 , RIfce5fe8_7639, \16371 );
nor \g453281/U$1 ( \24289 , \24287 , \24288 );
and \g453278/U$2 ( \24290 , \16380 , RIfcdc100_7526);
and \g453278/U$3 ( \24291 , RIf13ea10_5172, \16485 );
nor \g453278/U$1 ( \24292 , \24290 , \24291 );
and \g445372/U$2 ( \24293 , \24286 , \24289 , \24292 );
nor \g445372/U$1 ( \24294 , \24293 , \16649 );
or \g444228/U$1 ( \24295 , \24234 , \24264 , \24294 );
_DC \g437d/U$1 ( \24296 , \24295 , \16652 );
and \g453831/U$2 ( \24297 , \16361 , RIfe9ea18_8149);
and \g453831/U$3 ( \24298 , RIfceda40_7726, \16427 );
nor \g453831/U$1 ( \24299 , \24297 , \24298 );
and \g446003/U$2 ( \24300 , RIfc95d68_6727, \16448 );
and \g446003/U$3 ( \24301 , RIfe9eb80_8150, \16371 );
and \g448887/U$2 ( \24302 , RIdf273d0_1823, \16485 );
and \g448887/U$3 ( \24303 , \16356 , RIdf296f8_1848);
and \g448887/U$4 ( \24304 , RIdf1eb68_1726, \16398 );
nor \g448887/U$1 ( \24305 , \24302 , \24303 , \24304 );
and \g454574/U$2 ( \24306 , \16317 , RIfcd0328_7391);
and \g454574/U$3 ( \24307 , RIfc5e778_6097, \16325 );
nor \g454574/U$1 ( \24308 , \24306 , \24307 );
not \g450382/U$3 ( \24309 , \24308 );
not \g450382/U$4 ( \24310 , \16311 );
and \g450382/U$2 ( \24311 , \24309 , \24310 );
and \g450382/U$5 ( \24312 , \16341 , RIfcd01c0_7390);
nor \g450382/U$1 ( \24313 , \24311 , \24312 );
and \g451882/U$2 ( \24314 , \16377 , RIfcee6e8_7735);
and \g451882/U$3 ( \24315 , RIfc757e8_6359, \16313 );
nor \g451882/U$1 ( \24316 , \24314 , \24315 );
and \g451883/U$2 ( \24317 , \16334 , RIdf23b90_1783);
and \g451883/U$3 ( \24318 , RIdf257b0_1803, \16380 );
nor \g451883/U$1 ( \24319 , \24317 , \24318 );
nand \g447316/U$1 ( \24320 , \24305 , \24313 , \24316 , \24319 );
nor \g446003/U$1 ( \24321 , \24300 , \24301 , \24320 );
and \g451871/U$2 ( \24322 , \16364 , RIfe9ece8_8151);
and \g451871/U$3 ( \24323 , RIfc75518_6357, \16368 );
nor \g451871/U$1 ( \24324 , \24322 , \24323 );
nand \g445578/U$1 ( \24325 , \24299 , \24321 , \24324 );
and \g444834/U$2 ( \24326 , \24325 , \16481 );
and \g448880/U$2 ( \24327 , RIfc96308_6731, \16319 );
and \g448880/U$3 ( \24328 , \16328 , RIfc961a0_6730);
and \g448880/U$4 ( \24329 , RIded6610_903, \16398 );
nor \g448880/U$1 ( \24330 , \24327 , \24328 , \24329 );
and \g454976/U$2 ( \24331 , \16317 , RIdee1e48_1034);
and \g454976/U$3 ( \24332 , RIdee42d8_1060, \16325 );
nor \g454976/U$1 ( \24333 , \24331 , \24332 );
not \g449900/U$3 ( \24334 , \24333 );
not \g449900/U$4 ( \24335 , \16330 );
and \g449900/U$2 ( \24336 , \24334 , \24335 );
and \g449900/U$5 ( \24337 , \16341 , RIded8938_928);
nor \g449900/U$1 ( \24338 , \24336 , \24337 );
and \g451858/U$2 ( \24339 , \16377 , RIfce6150_7640);
and \g451858/U$3 ( \24340 , RIfc5ee80_6102, \16313 );
nor \g451858/U$1 ( \24341 , \24339 , \24340 );
and \g451860/U$2 ( \24342 , \16334 , RIdeddac8_986);
and \g451860/U$3 ( \24343 , RIdee00c0_1013, \16380 );
nor \g451860/U$1 ( \24344 , \24342 , \24343 );
nand \g447234/U$1 ( \24345 , \24330 , \24338 , \24341 , \24344 );
and \g444834/U$3 ( \24346 , \16477 , \24345 );
nor \g444834/U$1 ( \24347 , \24326 , \24346 );
and \g446786/U$2 ( \24348 , \17463 , RIded2290_855);
and \g446786/U$3 ( \24349 , RIfc75248_6355, \17465 );
nor \g446786/U$1 ( \24350 , \24348 , \24349 );
and \g446785/U$2 ( \24351 , \17468 , RIded4450_879);
and \g446785/U$3 ( \24352 , RIfc96470_6732, \17470 );
nor \g446785/U$1 ( \24353 , \24351 , \24352 );
and \g446790/U$2 ( \24354 , \17473 , RIfcb0618_7029);
and \g446790/U$3 ( \24355 , RIfc74ca8_6351, \17475 );
nor \g446790/U$1 ( \24356 , \24354 , \24355 );
nand \g444598/U$1 ( \24357 , \24347 , \24350 , \24353 , \24356 );
and \g448865/U$2 ( \24358 , RIde8c1c8_273, \16485 );
and \g448865/U$3 ( \24359 , \16354 , RIfe9e8b0_8148);
and \g448865/U$4 ( \24360 , RIe16a9a0_2590, \16398 );
nor \g448865/U$1 ( \24361 , \24358 , \24359 , \24360 );
and \g454692/U$2 ( \24362 , \16317 , RIfc957c8_6723);
and \g454692/U$3 ( \24363 , RIee1c840_4783, \16325 );
nor \g454692/U$1 ( \24364 , \24362 , \24363 );
not \g449887/U$3 ( \24365 , \24364 );
not \g449887/U$4 ( \24366 , \16311 );
and \g449887/U$2 ( \24367 , \24365 , \24366 );
and \g449887/U$5 ( \24368 , \16341 , RIfc95390_6720);
nor \g449887/U$1 ( \24369 , \24367 , \24368 );
and \g451823/U$2 ( \24370 , \16377 , RIfc5e610_6096);
and \g451823/U$3 ( \24371 , RIfcc8e70_7308, \16313 );
nor \g451823/U$1 ( \24372 , \24370 , \24371 );
and \g451824/U$2 ( \24373 , \16334 , RIde83b40_232);
and \g451824/U$3 ( \24374 , RIde88028_253, \16380 );
nor \g451824/U$1 ( \24375 , \24373 , \24374 );
nand \g447311/U$1 ( \24376 , \24361 , \24369 , \24372 , \24375 );
and \g444678/U$2 ( \24377 , \24376 , \17998 );
and \g445994/U$2 ( \24378 , RIfcebb50_7704, \16448 );
and \g445994/U$3 ( \24379 , RIde9a778_343, \16361 );
and \g448873/U$2 ( \24380 , RIdec1490_663, \16321 );
and \g448873/U$3 ( \24381 , \16328 , RIdec4190_695);
and \g448873/U$4 ( \24382 , RIdea7978_407, \16398 );
nor \g448873/U$1 ( \24383 , \24380 , \24381 , \24382 );
and \g454589/U$2 ( \24384 , \16317 , RIdebba90_599);
and \g454589/U$3 ( \24385 , RIfc954f8_6721, \16325 );
nor \g454589/U$1 ( \24386 , \24384 , \24385 );
not \g449895/U$3 ( \24387 , \24386 );
not \g449895/U$4 ( \24388 , \16330 );
and \g449895/U$2 ( \24389 , \24387 , \24388 );
and \g449895/U$5 ( \24390 , \16341 , RIfcdf0d0_7560);
nor \g449895/U$1 ( \24391 , \24389 , \24390 );
and \g451200/U$2 ( \24392 , \16377 , RIdebe790_631);
and \g451200/U$3 ( \24393 , RIfceaa70_7692, \16313 );
nor \g451200/U$1 ( \24394 , \24392 , \24393 );
and \g451846/U$2 ( \24395 , \16334 , RIdeb6090_535);
and \g451846/U$3 ( \24396 , RIdeb8d90_567, \16380 );
nor \g451846/U$1 ( \24397 , \24395 , \24396 );
nand \g447314/U$1 ( \24398 , \24383 , \24391 , \24394 , \24397 );
nor \g445994/U$1 ( \24399 , \24378 , \24379 , \24398 );
and \g451838/U$2 ( \24400 , \16364 , RIdea1078_375);
and \g451838/U$3 ( \24401 , RIdead990_439, \16368 );
nor \g451838/U$1 ( \24402 , \24400 , \24401 );
and \g451836/U$2 ( \24403 , \16371 , RIee1e190_4801);
and \g451836/U$3 ( \24404 , RIdeb0690_471, \16427 );
nor \g451836/U$1 ( \24405 , \24403 , \24404 );
and \g445143/U$2 ( \24406 , \24399 , \24402 , \24405 );
nor \g445143/U$1 ( \24407 , \24406 , \16618 );
nor \g444678/U$1 ( \24408 , \24377 , \24407 );
and \g446774/U$2 ( \24409 , \18523 , RIfca4c78_6897);
and \g446774/U$3 ( \24410 , RIfcb0bb8_7033, \18525 );
nor \g446774/U$1 ( \24411 , \24409 , \24410 );
and \g446775/U$2 ( \24412 , \18528 , RIfc75d88_6363);
and \g446775/U$3 ( \24413 , RIfca4b10_6896, \18530 );
nor \g446775/U$1 ( \24414 , \24412 , \24413 );
and \g446776/U$2 ( \24415 , \18533 , RIe166e90_2548);
and \g446776/U$3 ( \24416 , RIfcc8fd8_7309, \18535 );
nor \g446776/U$1 ( \24417 , \24415 , \24416 );
nand \g444481/U$1 ( \24418 , \24408 , \24411 , \24414 , \24417 );
and \g445977/U$2 ( \24419 , RIdef9b60_1305, \16427 );
and \g445977/U$3 ( \24420 , RIdef4160_1241, \16368 );
and \g448852/U$2 ( \24421 , RIdf13060_1593, \16321 );
and \g448852/U$3 ( \24422 , \16328 , RIdf15d60_1625);
and \g448852/U$4 ( \24423 , RIdeee760_1177, \16398 );
nor \g448852/U$1 ( \24424 , \24421 , \24422 , \24423 );
and \g455069/U$2 ( \24425 , \16317 , RIdf07c60_1465);
and \g455069/U$3 ( \24426 , RIdf0a960_1497, \16325 );
nor \g455069/U$1 ( \24427 , \24425 , \24426 );
not \g449876/U$3 ( \24428 , \24427 );
not \g449876/U$4 ( \24429 , \16330 );
and \g449876/U$2 ( \24430 , \24428 , \24429 );
and \g449876/U$5 ( \24431 , \16339 , RIdef1460_1209);
nor \g449876/U$1 ( \24432 , \24430 , \24431 );
and \g453077/U$2 ( \24433 , \16377 , RIdf0d660_1529);
and \g453077/U$3 ( \24434 , RIdf10360_1561, \16313 );
nor \g453077/U$1 ( \24435 , \24433 , \24434 );
and \g451780/U$2 ( \24436 , \16334 , RIdf02260_1401);
and \g451780/U$3 ( \24437 , RIdf04f60_1433, \16380 );
nor \g451780/U$1 ( \24438 , \24436 , \24437 );
nand \g447307/U$1 ( \24439 , \24424 , \24432 , \24435 , \24438 );
nor \g445977/U$1 ( \24440 , \24419 , \24420 , \24439 );
and \g451775/U$2 ( \24441 , \16361 , RIdee8d60_1113);
and \g451775/U$3 ( \24442 , RIdefc860_1337, \16432 );
nor \g451775/U$1 ( \24443 , \24441 , \24442 );
and \g451774/U$2 ( \24444 , \16364 , RIdeeba60_1145);
and \g451774/U$3 ( \24445 , RIdef6e60_1273, \16371 );
nor \g451774/U$1 ( \24446 , \24444 , \24445 );
and \g445131/U$2 ( \24447 , \24440 , \24443 , \24446 );
nor \g445131/U$1 ( \24448 , \24447 , \16555 );
and \g445984/U$2 ( \24449 , RIdf36f88_2002, \16427 );
and \g445984/U$3 ( \24450 , RIdf1be68_1694, \16368 );
and \g448936/U$2 ( \24451 , RIde93e78_311, \16485 );
and \g448936/U$3 ( \24452 , \16356 , RIdeb3390_503);
and \g448936/U$4 ( \24453 , RIdee6060_1081, \16398 );
nor \g448936/U$1 ( \24454 , \24451 , \24452 , \24453 );
and \g454738/U$2 ( \24455 , \16317 , RIdecc890_791);
and \g454738/U$3 ( \24456 , RIdecf590_823, \16325 );
nor \g454738/U$1 ( \24457 , \24455 , \24456 );
not \g449880/U$3 ( \24458 , \24457 );
not \g449880/U$4 ( \24459 , \16311 );
and \g449880/U$2 ( \24460 , \24458 , \24459 );
and \g449880/U$5 ( \24461 , \16341 , RIdeff560_1369);
nor \g449880/U$1 ( \24462 , \24460 , \24461 );
and \g451800/U$2 ( \24463 , \16377 , RIdec6e90_727);
and \g451800/U$3 ( \24464 , RIdec9b90_759, \16313 );
nor \g451800/U$1 ( \24465 , \24463 , \24464 );
and \g451804/U$2 ( \24466 , \16334 , RIe158d90_2388);
and \g451804/U$3 ( \24467 , RIe16cf98_2617, \16380 );
nor \g451804/U$1 ( \24468 , \24466 , \24467 );
nand \g447309/U$1 ( \24469 , \24454 , \24462 , \24465 , \24468 );
nor \g445984/U$1 ( \24470 , \24449 , \24450 , \24469 );
and \g451794/U$2 ( \24471 , \16361 , RIde79dc0_184);
and \g451794/U$3 ( \24472 , RIe142590_2132, \16448 );
nor \g451794/U$1 ( \24473 , \24471 , \24472 );
and \g452701/U$2 ( \24474 , \16364 , RIdedadc8_954);
and \g452701/U$3 ( \24475 , RIdf2b5e8_1870, \16371 );
nor \g452701/U$1 ( \24476 , \24474 , \24475 );
and \g445139/U$2 ( \24477 , \24470 , \24473 , \24476 );
nor \g445139/U$1 ( \24478 , \24477 , \16586 );
or \g444353/U$1 ( \24479 , \24357 , \24418 , \24448 , \24478 );
and \g445967/U$2 ( \24480 , RIe164190_2516, \16326 );
and \g445967/U$3 ( \24481 , RIe153390_2324, \16334 );
and \g448838/U$2 ( \24482 , RIe150690_2292, \16427 );
and \g448838/U$3 ( \24483 , \16448 , RIfc3ecc0_5740);
and \g448838/U$4 ( \24484 , RIe15ba90_2420, \16485 );
nor \g448838/U$1 ( \24485 , \24482 , \24483 , \24484 );
and \g454381/U$2 ( \24486 , \16317 , RIe14ac90_2228);
and \g454381/U$3 ( \24487 , RIfca6730_6916, \16325 );
nor \g454381/U$1 ( \24488 , \24486 , \24487 );
not \g454380/U$1 ( \24489 , \24488 );
and \g449862/U$2 ( \24490 , \24489 , \16336 );
and \g449862/U$3 ( \24491 , RIfc74f78_6353, \16356 );
nor \g449862/U$1 ( \24492 , \24490 , \24491 );
and \g451735/U$2 ( \24493 , \16361 , RIe145290_2164);
and \g451735/U$3 ( \24494 , RIe147f90_2196, \16364 );
nor \g451735/U$1 ( \24495 , \24493 , \24494 );
and \g451734/U$2 ( \24496 , \16368 , RIe14d990_2260);
and \g451734/U$3 ( \24497 , RIfce8b80_7670, \16371 );
nor \g451734/U$1 ( \24498 , \24496 , \24497 );
nand \g448053/U$1 ( \24499 , \24485 , \24492 , \24495 , \24498 );
nor \g445967/U$1 ( \24500 , \24480 , \24481 , \24499 );
and \g451727/U$2 ( \24501 , \16377 , RIe15e790_2452);
and \g451727/U$3 ( \24502 , RIe156090_2356, \16380 );
nor \g451727/U$1 ( \24503 , \24501 , \24502 );
and \g451726/U$2 ( \24504 , \16313 , RIfe9e748_8147);
and \g451726/U$3 ( \24505 , RIe161490_2484, \16321 );
nor \g451726/U$1 ( \24506 , \24504 , \24505 );
and \g445122/U$2 ( \24507 , \24500 , \24503 , \24506 );
nor \g445122/U$1 ( \24508 , \24507 , \16389 );
and \g445972/U$2 ( \24509 , RIfc5f2b8_6105, \16321 );
and \g445972/U$3 ( \24510 , RIfc753b0_6356, \16313 );
and \g448844/U$2 ( \24511 , RIdf327d0_1951, \16398 );
and \g448844/U$3 ( \24512 , \16341 , RIdf34828_1974);
and \g448844/U$4 ( \24513 , RIdf3e170_2083, \16485 );
nor \g448844/U$1 ( \24514 , \24511 , \24512 , \24513 );
and \g455377/U$2 ( \24515 , \16317 , RIfcc1850_7224);
and \g455377/U$3 ( \24516 , RIfcc1c88_7227, \16325 );
nor \g455377/U$1 ( \24517 , \24515 , \24516 );
not \g449869/U$3 ( \24518 , \24517 );
not \g449869/U$4 ( \24519 , \16351 );
and \g449869/U$2 ( \24520 , \24518 , \24519 );
and \g449869/U$5 ( \24521 , \16356 , RIe140268_2107);
nor \g449869/U$1 ( \24522 , \24520 , \24521 );
and \g451763/U$2 ( \24523 , \16361 , RIdf2e2e8_1902);
and \g451763/U$3 ( \24524 , RIdf301d8_1924, \16364 );
nor \g451763/U$1 ( \24525 , \24523 , \24524 );
and \g451758/U$2 ( \24526 , \16368 , RIfc96038_6729);
and \g451758/U$3 ( \24527 , RIfc965d8_6733, \16371 );
nor \g451758/U$1 ( \24528 , \24526 , \24527 );
nand \g447642/U$1 ( \24529 , \24514 , \24522 , \24525 , \24528 );
nor \g445972/U$1 ( \24530 , \24509 , \24510 , \24529 );
and \g451751/U$2 ( \24531 , \16377 , RIfc74b40_6350);
and \g451751/U$3 ( \24532 , RIdf3be48_2058, \16380 );
nor \g451751/U$1 ( \24533 , \24531 , \24532 );
and \g454042/U$2 ( \24534 , \16334 , RIdf39c88_2034);
and \g454042/U$3 ( \24535 , RIfcee2b0_7732, \16326 );
nor \g454042/U$1 ( \24536 , \24534 , \24535 );
and \g445125/U$2 ( \24537 , \24530 , \24533 , \24536 );
nor \g445125/U$1 ( \24538 , \24537 , \16393 );
or \g444212/U$1 ( \24539 , \24479 , \24508 , \24538 );
_DC \g44da/U$1 ( \24540 , \24539 , \16652 );
and \g449177/U$2 ( \24541 , RIe209280_4394, \8319 );
and \g449177/U$3 ( \24542 , \8326 , RIe20bf80_4426);
and \g449177/U$4 ( \24543 , RIe211980_4490, \8488 );
nor \g449177/U$1 ( \24544 , \24541 , \24542 , \24543 );
and \g452890/U$2 ( \24545 , \8335 , RIe206580_4362);
and \g452890/U$3 ( \24546 , RIfcc0770_7212, \8340 );
nor \g452890/U$1 ( \24547 , \24545 , \24546 );
and \g452889/U$2 ( \24548 , \8404 , RIe21fa80_4650);
and \g452889/U$3 ( \24549 , RIfc40340_5756, \8351 );
nor \g452889/U$1 ( \24550 , \24548 , \24549 );
and \g455082/U$2 ( \24551 , \8313 , RIfcdd618_7541);
and \g455082/U$3 ( \24552 , RIe222780_4682, \8323 );
nor \g455082/U$1 ( \24553 , \24551 , \24552 );
not \g450194/U$3 ( \24554 , \24553 );
not \g450194/U$4 ( \24555 , \8328 );
and \g450194/U$2 ( \24556 , \24554 , \24555 );
and \g450194/U$5 ( \24557 , \8359 , RIfec4998_8357);
nor \g450194/U$1 ( \24558 , \24556 , \24557 );
nand \g447813/U$1 ( \24559 , \24544 , \24547 , \24550 , \24558 );
and \g444788/U$2 ( \24560 , \24559 , \8369 );
and \g446234/U$2 ( \24561 , RIfec4c68_8359, \8371 );
and \g446234/U$3 ( \24562 , RIfc94c88_6715, \8319 );
and \g449182/U$2 ( \24563 , RIfe9e040_8142, \8531 );
and \g449182/U$3 ( \24564 , \8488 , RIfcc08d8_7213);
and \g449182/U$4 ( \24565 , RIfcee580_7734, \8330 );
nor \g449182/U$1 ( \24566 , \24563 , \24564 , \24565 );
and \g452902/U$2 ( \24567 , \8356 , RIfe9e1a8_8143);
and \g452902/U$3 ( \24568 , RIfccd088_7355, \8359 );
nor \g452902/U$1 ( \24569 , \24567 , \24568 );
and \g455091/U$2 ( \24570 , \8313 , RIf162938_5581);
and \g455091/U$3 ( \24571 , RIfcebcb8_7705, \8323 );
nor \g455091/U$1 ( \24572 , \24570 , \24571 );
not \g450198/U$3 ( \24573 , \24572 );
not \g450198/U$4 ( \24574 , \8376 );
and \g450198/U$2 ( \24575 , \24573 , \24574 );
and \g450198/U$5 ( \24576 , \8351 , RIfce2370_7596);
nor \g450198/U$1 ( \24577 , \24575 , \24576 );
and \g452901/U$2 ( \24578 , \8378 , RIf1612b8_5565);
and \g452901/U$3 ( \24579 , RIfc949b8_6713, \8417 );
nor \g452901/U$1 ( \24580 , \24578 , \24579 );
nand \g447815/U$1 ( \24581 , \24566 , \24569 , \24577 , \24580 );
nor \g446234/U$1 ( \24582 , \24561 , \24562 , \24581 );
and \g452896/U$2 ( \24583 , \8335 , RIfccc3e0_7346);
and \g452896/U$3 ( \24584 , RIfcead40_7694, \8340 );
nor \g452896/U$1 ( \24585 , \24583 , \24584 );
and \g452894/U$2 ( \24586 , \8326 , RIf15ad78_5493);
and \g452894/U$3 ( \24587 , RIfec4b00_8358, \8404 );
nor \g452894/U$1 ( \24588 , \24586 , \24587 );
and \g445314/U$2 ( \24589 , \24582 , \24585 , \24588 );
nor \g445314/U$1 ( \24590 , \24589 , \8422 );
nor \g444788/U$1 ( \24591 , \24560 , \24590 );
and \g447003/U$2 ( \24592 , \8438 , RIe214680_4522);
and \g447003/U$3 ( \24593 , RIe217380_4554, \8440 );
nor \g447003/U$1 ( \24594 , \24592 , \24593 );
and \g447004/U$2 ( \24595 , \8431 , RIe21cd80_4618);
and \g447004/U$3 ( \24596 , RIfcd0b98_7397, \8434 );
nor \g447004/U$1 ( \24597 , \24595 , \24596 );
and \g447005/U$2 ( \24598 , \8717 , RIe20ec80_4458);
and \g447005/U$3 ( \24599 , RIf168608_5647, \8719 );
nor \g447005/U$1 ( \24600 , \24598 , \24599 );
nand \g444514/U$1 ( \24601 , \24591 , \24594 , \24597 , \24600 );
and \g452919/U$2 ( \24602 , \8326 , RIe1ba7e8_3499);
and \g452919/U$3 ( \24603 , RIe19f128_3187, \8404 );
nor \g452919/U$1 ( \24604 , \24602 , \24603 );
and \g446239/U$2 ( \24605 , RIe1a1e28_3219, \8371 );
and \g446239/U$3 ( \24606 , RIe1ad660_3350, \8317 );
and \g449188/U$2 ( \24607 , RIe1f6c98_4185, \8531 );
and \g449188/U$3 ( \24608 , \8488 , RIe1fd8e0_4262);
and \g449188/U$4 ( \24609 , RIe1a4b28_3251, \8383 );
nor \g449188/U$1 ( \24610 , \24607 , \24608 , \24609 );
and \g452929/U$2 ( \24611 , \8356 , RIe1ef7e0_4102);
and \g452929/U$3 ( \24612 , RIe203880_4330, \8359 );
nor \g452929/U$1 ( \24613 , \24611 , \24612 );
and \g455000/U$2 ( \24614 , \8313 , RIe225480_4714);
and \g455000/U$3 ( \24615 , RIe177b28_2739, \8323 );
nor \g455000/U$1 ( \24616 , \24614 , \24615 );
not \g450204/U$3 ( \24617 , \24616 );
not \g450204/U$4 ( \24618 , \8376 );
and \g450204/U$2 ( \24619 , \24617 , \24618 );
and \g450204/U$5 ( \24620 , \8351 , RIe1a7828_3283);
nor \g450204/U$1 ( \24621 , \24619 , \24620 );
and \g452927/U$2 ( \24622 , \8378 , RIe21a080_4586);
and \g452927/U$3 ( \24623 , RIe18b628_2963, \8417 );
nor \g452927/U$1 ( \24624 , \24622 , \24623 );
nand \g447820/U$1 ( \24625 , \24610 , \24613 , \24621 , \24624 );
nor \g446239/U$1 ( \24626 , \24605 , \24606 , \24625 );
and \g452921/U$2 ( \24627 , \8335 , RIe16fc98_2649);
and \g452921/U$3 ( \24628 , RIe1d3ce8_3787, \8340 );
nor \g452921/U$1 ( \24629 , \24627 , \24628 );
nand \g445639/U$1 ( \24630 , \24604 , \24626 , \24629 );
and \g444881/U$2 ( \24631 , \24630 , \9010 );
and \g449185/U$2 ( \24632 , RIfcc0e78_7217, \8319 );
and \g449185/U$3 ( \24633 , \8326 , RIfc950c0_6718);
and \g449185/U$4 ( \24634 , RIf1512c8_5383, \8486 );
nor \g449185/U$1 ( \24635 , \24632 , \24633 , \24634 );
and \g452914/U$2 ( \24636 , \8335 , RIe1ed1e8_4075);
and \g452914/U$3 ( \24637 , RIfc761c0_6366, \8340 );
nor \g452914/U$1 ( \24638 , \24636 , \24637 );
and \g452911/U$2 ( \24639 , \8404 , RIe1f9998_4217);
and \g452911/U$3 ( \24640 , RIfc765f8_6369, \8351 );
nor \g452911/U$1 ( \24641 , \24639 , \24640 );
and \g455289/U$2 ( \24642 , \8313 , RIfcc0a40_7214);
and \g455289/U$3 ( \24643 , RIfc94df0_6716, \8323 );
nor \g455289/U$1 ( \24644 , \24642 , \24643 );
not \g450201/U$3 ( \24645 , \24644 );
not \g450201/U$4 ( \24646 , \8328 );
and \g450201/U$2 ( \24647 , \24645 , \24646 );
and \g450201/U$5 ( \24648 , \8359 , RIf152510_5396);
nor \g450201/U$1 ( \24649 , \24647 , \24648 );
nand \g447817/U$1 ( \24650 , \24635 , \24638 , \24641 , \24649 );
and \g444881/U$3 ( \24651 , \8752 , \24650 );
nor \g444881/U$1 ( \24652 , \24631 , \24651 );
and \g447009/U$2 ( \24653 , \11516 , RIfce8748_7667);
and \g447009/U$3 ( \24654 , RIfcc8d08_7307, \11518 );
nor \g447009/U$1 ( \24655 , \24653 , \24654 );
and \g447010/U$2 ( \24656 , \13486 , RIe1f24e0_4134);
and \g447010/U$3 ( \24657 , RIfcb0ff0_7036, \13488 );
nor \g447010/U$1 ( \24658 , \24656 , \24657 );
and \g447011/U$2 ( \24659 , \11521 , RIe1f4970_4160);
and \g447011/U$3 ( \24660 , RIfceb2e0_7698, \11523 );
nor \g447011/U$1 ( \24661 , \24659 , \24660 );
nand \g444637/U$1 ( \24662 , \24652 , \24655 , \24658 , \24661 );
and \g446226/U$2 ( \24663 , RIe193d28_3059, \8409 );
and \g446226/U$3 ( \24664 , RIe18e328_2995, \8378 );
and \g449172/U$2 ( \24665 , RIfe9e310_8144, \8373 );
and \g449172/U$3 ( \24666 , \8383 , RIe199728_3123);
and \g449172/U$4 ( \24667 , RIe185c28_2899, \8486 );
nor \g449172/U$1 ( \24668 , \24665 , \24666 , \24667 );
and \g452868/U$2 ( \24669 , \8335 , RIe17a828_2771);
and \g452868/U$3 ( \24670 , RIfe9e478_8145, \8340 );
nor \g452868/U$1 ( \24671 , \24669 , \24670 );
and \g452866/U$2 ( \24672 , \8404 , RIe196a28_3091);
and \g452866/U$3 ( \24673 , RIe19c428_3155, \8351 );
nor \g452866/U$1 ( \24674 , \24672 , \24673 );
and \g455059/U$2 ( \24675 , \8313 , RIe17d528_2803);
and \g455059/U$3 ( \24676 , RIe180228_2835, \8323 );
nor \g455059/U$1 ( \24677 , \24675 , \24676 );
not \g455058/U$1 ( \24678 , \24677 );
and \g450187/U$2 ( \24679 , \24678 , \8316 );
and \g450187/U$3 ( \24680 , RIe188928_2931, \8359 );
nor \g450187/U$1 ( \24681 , \24679 , \24680 );
nand \g448206/U$1 ( \24682 , \24668 , \24671 , \24674 , \24681 );
nor \g446226/U$1 ( \24683 , \24663 , \24664 , \24682 );
and \g452861/U$2 ( \24684 , \8356 , RIe182f28_2867);
and \g452861/U$3 ( \24685 , RIfcc04a0_7210, \8417 );
nor \g452861/U$1 ( \24686 , \24684 , \24685 );
and \g452859/U$2 ( \24687 , \8523 , RIfce1830_7588);
and \g452859/U$3 ( \24688 , RIe191028_3027, \8412 );
nor \g452859/U$1 ( \24689 , \24687 , \24688 );
and \g445309/U$2 ( \24690 , \24683 , \24686 , \24689 );
nor \g445309/U$1 ( \24691 , \24690 , \8589 );
and \g446229/U$2 ( \24692 , RIfc94418_6709, \8373 );
and \g446229/U$3 ( \24693 , RIfce7230_7652, \8335 );
and \g449174/U$2 ( \24694 , RIfce5fe8_7639, \8531 );
and \g449174/U$3 ( \24695 , \8486 , RIfced338_7721);
and \g449174/U$4 ( \24696 , RIfcb12c0_7038, \8383 );
nor \g449174/U$1 ( \24697 , \24694 , \24695 , \24696 );
and \g452880/U$2 ( \24698 , \8356 , RIe172998_2681);
and \g452880/U$3 ( \24699 , RIfc946e8_6711, \8359 );
nor \g452880/U$1 ( \24700 , \24698 , \24699 );
and \g455133/U$2 ( \24701 , \8313 , RIfcdc100_7526);
and \g455133/U$3 ( \24702 , RIf13ea10_5172, \8323 );
nor \g455133/U$1 ( \24703 , \24701 , \24702 );
not \g450191/U$3 ( \24704 , \24703 );
not \g450191/U$4 ( \24705 , \8376 );
and \g450191/U$2 ( \24706 , \24704 , \24705 );
and \g450191/U$5 ( \24707 , \8351 , RIf141878_5205);
nor \g450191/U$1 ( \24708 , \24706 , \24707 );
and \g452879/U$2 ( \24709 , \8378 , RIfc94580_6710);
and \g452879/U$3 ( \24710 , RIfc77408_6379, \8417 );
nor \g452879/U$1 ( \24711 , \24709 , \24710 );
nand \g447811/U$1 ( \24712 , \24697 , \24700 , \24708 , \24711 );
nor \g446229/U$1 ( \24713 , \24692 , \24693 , \24712 );
and \g452872/U$2 ( \24714 , \8340 , RIfcdc268_7527);
and \g452872/U$3 ( \24715 , RIe174f90_2708, \8404 );
nor \g452872/U$1 ( \24716 , \24714 , \24715 );
and \g452875/U$2 ( \24717 , \8319 , RIfcc0608_7211);
and \g452875/U$3 ( \24718 , RIfcddff0_7548, \8326 );
nor \g452875/U$1 ( \24719 , \24717 , \24718 );
and \g445311/U$2 ( \24720 , \24713 , \24716 , \24719 );
nor \g445311/U$1 ( \24721 , \24720 , \8558 );
or \g444404/U$1 ( \24722 , \24601 , \24662 , \24691 , \24721 );
and \g446220/U$2 ( \24723 , RIfcd0760_7394, \8340 );
and \g446220/U$3 ( \24724 , RIe1b65d0_3452, \8404 );
and \g449166/U$2 ( \24725 , RIe1b1f80_3402, \8531 );
and \g449166/U$3 ( \24726 , \8488 , RIfceaea8_7695);
and \g449166/U$4 ( \24727 , RIf14ac20_5310, \8383 );
nor \g449166/U$1 ( \24728 , \24725 , \24726 , \24727 );
and \g452839/U$2 ( \24729 , \8356 , RIe1b0360_3382);
and \g452839/U$3 ( \24730 , RIfcc0fe0_7218, \8359 );
nor \g452839/U$1 ( \24731 , \24729 , \24730 );
and \g455047/U$2 ( \24732 , \8313 , RIe1b4c80_3434);
and \g455047/U$3 ( \24733 , RIfc76490_6368, \8323 );
nor \g455047/U$1 ( \24734 , \24732 , \24733 );
not \g450181/U$3 ( \24735 , \24734 );
not \g450181/U$4 ( \24736 , \8376 );
and \g450181/U$2 ( \24737 , \24735 , \24736 );
and \g450181/U$5 ( \24738 , \8351 , RIf14bfd0_5324);
nor \g450181/U$1 ( \24739 , \24737 , \24738 );
and \g452838/U$2 ( \24740 , \8378 , RIe1b38d0_3420);
and \g452838/U$3 ( \24741 , RIfcecd98_7717, \8417 );
nor \g452838/U$1 ( \24742 , \24740 , \24741 );
nand \g447808/U$1 ( \24743 , \24728 , \24731 , \24739 , \24742 );
nor \g446220/U$1 ( \24744 , \24723 , \24724 , \24743 );
and \g452832/U$2 ( \24745 , \8335 , RIfe9dd70_8140);
and \g452832/U$3 ( \24746 , RIfe9ded8_8141, \8373 );
nor \g452832/U$1 ( \24747 , \24745 , \24746 );
and \g452834/U$2 ( \24748 , \8319 , RIfe9e5e0_8146);
and \g452834/U$3 ( \24749 , RIf145ec8_5255, \8326 );
nor \g452834/U$1 ( \24750 , \24748 , \24749 );
and \g445304/U$2 ( \24751 , \24744 , \24747 , \24750 );
nor \g445304/U$1 ( \24752 , \24751 , \8481 );
and \g446222/U$2 ( \24753 , RIe1dc3e8_3883, \8407 );
and \g446222/U$3 ( \24754 , RIe1d69e8_3819, \8378 );
and \g449168/U$2 ( \24755 , RIe1c01e8_3563, \8319 );
and \g449168/U$3 ( \24756 , \8326 , RIe1c2ee8_3595);
and \g449168/U$4 ( \24757 , RIe1ce2e8_3723, \8486 );
nor \g449168/U$1 ( \24758 , \24755 , \24756 , \24757 );
and \g452853/U$2 ( \24759 , \8335 , RIe1bd4e8_3531);
and \g452853/U$3 ( \24760 , RIe1c5be8_3627, \8340 );
nor \g452853/U$1 ( \24761 , \24759 , \24760 );
and \g452851/U$2 ( \24762 , \8404 , RIe1e1de8_3947);
and \g452851/U$3 ( \24763 , RIe1ea4e8_4043, \8351 );
nor \g452851/U$1 ( \24764 , \24762 , \24763 );
and \g455209/U$2 ( \24765 , \8313 , RIe1e4ae8_3979);
and \g455209/U$3 ( \24766 , RIe1e77e8_4011, \8323 );
nor \g455209/U$1 ( \24767 , \24765 , \24766 );
not \g450183/U$3 ( \24768 , \24767 );
not \g450183/U$4 ( \24769 , \8328 );
and \g450183/U$2 ( \24770 , \24768 , \24769 );
and \g450183/U$5 ( \24771 , \8359 , RIe1d0fe8_3755);
nor \g450183/U$1 ( \24772 , \24770 , \24771 );
nand \g447809/U$1 ( \24773 , \24758 , \24761 , \24764 , \24772 );
nor \g446222/U$1 ( \24774 , \24753 , \24754 , \24773 );
and \g452848/U$2 ( \24775 , \8356 , RIe1c88e8_3659);
and \g452848/U$3 ( \24776 , RIe1df0e8_3915, \8417 );
nor \g452848/U$1 ( \24777 , \24775 , \24776 );
and \g452844/U$2 ( \24778 , \8531 , RIe1cb5e8_3691);
and \g452844/U$3 ( \24779 , RIe1d96e8_3851, \8414 );
nor \g452844/U$1 ( \24780 , \24778 , \24779 );
and \g445307/U$2 ( \24781 , \24774 , \24777 , \24780 );
nor \g445307/U$1 ( \24782 , \24781 , \8477 );
or \g444201/U$1 ( \24783 , \24722 , \24752 , \24782 );
_DC \g455e/U$1 ( \24784 , \24783 , \8654 );
and \g449480/U$2 ( \24785 , RIdf13fd8_1604, \16321 );
and \g449480/U$3 ( \24786 , \16328 , RIdf16cd8_1636);
and \g449480/U$4 ( \24787 , RIdeef6d8_1188, \16337 );
nor \g449480/U$1 ( \24788 , \24785 , \24786 , \24787 );
and \g455385/U$2 ( \24789 , \16317 , RIdf08bd8_1476);
and \g455385/U$3 ( \24790 , RIdf0b8d8_1508, \16325 );
nor \g455385/U$1 ( \24791 , \24789 , \24790 );
not \g450501/U$3 ( \24792 , \24791 );
not \g450501/U$4 ( \24793 , \16330 );
and \g450501/U$2 ( \24794 , \24792 , \24793 );
and \g450501/U$5 ( \24795 , \16341 , RIdef23d8_1220);
nor \g450501/U$1 ( \24796 , \24794 , \24795 );
and \g454000/U$2 ( \24797 , \16377 , RIdf0e5d8_1540);
and \g454000/U$3 ( \24798 , RIdf112d8_1572, \16313 );
nor \g454000/U$1 ( \24799 , \24797 , \24798 );
and \g454004/U$2 ( \24800 , \16334 , RIdf031d8_1412);
and \g454004/U$3 ( \24801 , RIdf05ed8_1444, \16380 );
nor \g454004/U$1 ( \24802 , \24800 , \24801 );
nand \g447443/U$1 ( \24803 , \24788 , \24796 , \24799 , \24802 );
and \g444719/U$2 ( \24804 , \24803 , \16750 );
and \g446472/U$2 ( \24805 , RIfcb1c98_7045, \16448 );
and \g446472/U$3 ( \24806 , RIfe9d938_8137, \16361 );
and \g449485/U$2 ( \24807 , RIfea8bd0_8236, \16485 );
and \g449485/U$3 ( \24808 , \16354 , RIfe9d668_8135);
and \g449485/U$4 ( \24809 , RIdf1f6a8_1734, \16337 );
nor \g449485/U$1 ( \24810 , \24807 , \24808 , \24809 );
and \g455014/U$2 ( \24811 , \16317 , RIfc93ba8_6703);
and \g455014/U$3 ( \24812 , RIee2ba20_4955, \16325 );
nor \g455014/U$1 ( \24813 , \24811 , \24812 );
not \g450505/U$3 ( \24814 , \24813 );
not \g450505/U$4 ( \24815 , \16311 );
and \g450505/U$2 ( \24816 , \24814 , \24815 );
and \g450505/U$5 ( \24817 , \16341 , RIdf21598_1756);
nor \g450505/U$1 ( \24818 , \24816 , \24817 );
and \g454019/U$2 ( \24819 , \16377 , RIee27ad8_4910);
and \g454019/U$3 ( \24820 , RIfc77de0_6386, \16313 );
nor \g454019/U$1 ( \24821 , \24819 , \24820 );
and \g454021/U$2 ( \24822 , \16334 , RIfe9d7d0_8136);
and \g454021/U$3 ( \24823 , RIdf26458_1812, \16380 );
nor \g454021/U$1 ( \24824 , \24822 , \24823 );
nand \g447445/U$1 ( \24825 , \24810 , \24818 , \24821 , \24824 );
nor \g446472/U$1 ( \24826 , \24805 , \24806 , \24825 );
and \g454013/U$2 ( \24827 , \16364 , RIdf1aef0_1683);
and \g454013/U$3 ( \24828 , RIfcc0068_7207, \16368 );
nor \g454013/U$1 ( \24829 , \24827 , \24828 );
and \g454011/U$2 ( \24830 , \16371 , RIdf22ab0_1771);
and \g454011/U$3 ( \24831 , RIee26cc8_4900, \16427 );
nor \g454011/U$1 ( \24832 , \24830 , \24831 );
and \g445480/U$2 ( \24833 , \24826 , \24829 , \24832 );
nor \g445480/U$1 ( \24834 , \24833 , \16480 );
nor \g444719/U$1 ( \24835 , \24804 , \24834 );
and \g447211/U$2 ( \24836 , \19208 , RIdee9cd8_1124);
and \g447211/U$3 ( \24837 , RIdef7dd8_1284, \19210 );
nor \g447211/U$1 ( \24838 , \24836 , \24837 );
and \g447212/U$2 ( \24839 , \19213 , RIdeec9d8_1156);
and \g447212/U$3 ( \24840 , RIdef50d8_1252, \19215 );
nor \g447212/U$1 ( \24841 , \24839 , \24840 );
and \g447210/U$2 ( \24842 , \19218 , RIdefaad8_1316);
and \g447210/U$3 ( \24843 , RIdefd7d8_1348, \19220 );
nor \g447210/U$1 ( \24844 , \24842 , \24843 );
nand \g444665/U$1 ( \24845 , \24835 , \24838 , \24841 , \24844 );
and \g449469/U$2 ( \24846 , RIdebca08_610, \16485 );
and \g449469/U$3 ( \24847 , \16354 , RIfc934a0_6698);
and \g449469/U$4 ( \24848 , RIdea9d90_418, \16398 );
nor \g449469/U$1 ( \24849 , \24846 , \24847 , \24848 );
and \g454237/U$2 ( \24850 , \16317 , RIdec2408_674);
and \g454237/U$3 ( \24851 , RIdec5108_706, \16325 );
nor \g454237/U$1 ( \24852 , \24850 , \24851 );
not \g450492/U$3 ( \24853 , \24852 );
not \g450492/U$4 ( \24854 , \16311 );
and \g450492/U$2 ( \24855 , \24853 , \24854 );
and \g450492/U$5 ( \24856 , \16341 , RIfcc8498_7301);
nor \g450492/U$1 ( \24857 , \24855 , \24856 );
and \g453961/U$2 ( \24858 , \16377 , RIdebf708_642);
and \g453961/U$3 ( \24859 , RIfc93608_6699, \16313 );
nor \g453961/U$1 ( \24860 , \24858 , \24859 );
and \g453964/U$2 ( \24861 , \16334 , RIdeb7008_546);
and \g453964/U$3 ( \24862 , RIdeb9d08_578, \16380 );
nor \g453964/U$1 ( \24863 , \24861 , \24862 );
nand \g447439/U$1 ( \24864 , \24849 , \24857 , \24860 , \24863 );
and \g444713/U$2 ( \24865 , \24864 , \17938 );
and \g446464/U$2 ( \24866 , RIfceb718_7701, \16328 );
and \g446464/U$3 ( \24867 , RIfe9daa0_8138, \16334 );
and \g449475/U$2 ( \24868 , RIfcdbf98_7525, \16427 );
and \g449475/U$3 ( \24869 , \16448 , RIfce8478_7665);
and \g449475/U$4 ( \24870 , RIdf3ecb0_2091, \16485 );
nor \g449475/U$1 ( \24871 , \24868 , \24869 , \24870 );
and \g455398/U$2 ( \24872 , \16317 , RIdf33040_1957);
and \g455398/U$3 ( \24873 , RIdf354d0_1983, \16325 );
nor \g455398/U$1 ( \24874 , \24872 , \24873 );
not \g455397/U$1 ( \24875 , \24874 );
and \g450495/U$2 ( \24876 , \24875 , \16336 );
and \g450495/U$3 ( \24877 , RIe140da8_2115, \16356 );
nor \g450495/U$1 ( \24878 , \24876 , \24877 );
and \g453984/U$2 ( \24879 , \16361 , RIdf2ee28_1910);
and \g453984/U$3 ( \24880 , RIdf30fe8_1934, \16364 );
nor \g453984/U$1 ( \24881 , \24879 , \24880 );
and \g453981/U$2 ( \24882 , \16368 , RIfc93fe0_6706);
and \g453981/U$3 ( \24883 , RIfc776d8_6381, \16371 );
nor \g453981/U$1 ( \24884 , \24882 , \24883 );
nand \g448125/U$1 ( \24885 , \24871 , \24878 , \24881 , \24884 );
nor \g446464/U$1 ( \24886 , \24866 , \24867 , \24885 );
and \g453976/U$2 ( \24887 , \16377 , RIfce7938_7657);
and \g453976/U$3 ( \24888 , RIdf3c988_2066, \16380 );
nor \g453976/U$1 ( \24889 , \24887 , \24888 );
and \g453972/U$2 ( \24890 , \16313 , RIfc93e78_6705);
and \g453972/U$3 ( \24891 , RIfcb19c8_7043, \16319 );
nor \g453972/U$1 ( \24892 , \24890 , \24891 );
and \g445473/U$2 ( \24893 , \24886 , \24889 , \24892 );
nor \g445473/U$1 ( \24894 , \24893 , \16393 );
nor \g444713/U$1 ( \24895 , \24865 , \24894 );
and \g447200/U$2 ( \24896 , \18457 , RIdeb1608_482);
and \g447200/U$3 ( \24897 , RIfcdf7d8_7565, \18459 );
nor \g447200/U$1 ( \24898 , \24896 , \24897 );
and \g447205/U$2 ( \24899 , \18462 , RIdeae908_450);
and \g447205/U$3 ( \24900 , RIfc78218_6389, \18464 );
nor \g447205/U$1 ( \24901 , \24899 , \24900 );
and \g447204/U$2 ( \24902 , \18467 , RIde9cb90_354);
and \g447204/U$3 ( \24903 , RIdea3490_386, \18469 );
nor \g447204/U$1 ( \24904 , \24902 , \24903 );
nand \g444544/U$1 ( \24905 , \24895 , \24898 , \24901 , \24904 );
and \g446453/U$2 ( \24906 , RIee1cc78_4786, \16328 );
and \g446453/U$3 ( \24907 , RIde85238_239, \16334 );
and \g449460/U$2 ( \24908 , RIfc938d8_6701, \16427 );
and \g449460/U$3 ( \24909 , \16432 , RIde813e0_220);
and \g449460/U$4 ( \24910 , RIde8d578_279, \16344 );
nor \g449460/U$1 ( \24911 , \24908 , \24909 , \24910 );
and \g454544/U$2 ( \24912 , \16317 , RIe16b4e0_2598);
and \g454544/U$3 ( \24913 , RIfce8ce8_7671, \16325 );
nor \g454544/U$1 ( \24914 , \24912 , \24913 );
not \g454543/U$1 ( \24915 , \24914 );
and \g450480/U$2 ( \24916 , \24915 , \16336 );
and \g450480/U$3 ( \24917 , RIde909f8_295, \16354 );
nor \g450480/U$1 ( \24918 , \24916 , \24917 );
and \g453932/U$2 ( \24919 , \16361 , RIfea9f80_8250);
and \g453932/U$3 ( \24920 , RIfea8d38_8237, \16364 );
nor \g453932/U$1 ( \24921 , \24919 , \24920 );
and \g453928/U$2 ( \24922 , \16368 , RIfcbfd98_7205);
and \g453928/U$3 ( \24923 , RIfce5e80_7638, \16371 );
nor \g453928/U$1 ( \24924 , \24922 , \24923 );
nand \g448123/U$1 ( \24925 , \24911 , \24918 , \24921 , \24924 );
nor \g446453/U$1 ( \24926 , \24906 , \24907 , \24925 );
and \g453922/U$2 ( \24927 , \16377 , RIee1aab8_4762);
and \g453922/U$3 ( \24928 , RIfea8ea0_8238, \16380 );
nor \g453922/U$1 ( \24929 , \24927 , \24928 );
and \g453921/U$2 ( \24930 , \16313 , RIee1b328_4768);
and \g453921/U$3 ( \24931 , RIee1bb98_4774, \16319 );
nor \g453921/U$1 ( \24932 , \24930 , \24931 );
and \g445467/U$2 ( \24933 , \24926 , \24929 , \24932 );
nor \g445467/U$1 ( \24934 , \24933 , \16649 );
and \g446458/U$2 ( \24935 , RIe165108_2527, \16328 );
and \g446458/U$3 ( \24936 , RIe154308_2335, \16334 );
and \g449464/U$2 ( \24937 , RIe151608_2303, \16427 );
and \g449464/U$3 ( \24938 , \16448 , RIfea7550_8220);
and \g449464/U$4 ( \24939 , RIe15ca08_2431, \16485 );
nor \g449464/U$1 ( \24940 , \24937 , \24938 , \24939 );
and \g454390/U$2 ( \24941 , \16317 , RIe14bc08_2239);
and \g454390/U$3 ( \24942 , RIfcd1408_7403, \16325 );
nor \g454390/U$1 ( \24943 , \24941 , \24942 );
not \g454389/U$1 ( \24944 , \24943 );
and \g450483/U$2 ( \24945 , \24944 , \16336 );
and \g450483/U$3 ( \24946 , RIfe9dc08_8139, \16354 );
nor \g450483/U$1 ( \24947 , \24945 , \24946 );
and \g453949/U$2 ( \24948 , \16361 , RIe146208_2175);
and \g453949/U$3 ( \24949 , RIe148f08_2207, \16364 );
nor \g453949/U$1 ( \24950 , \24948 , \24949 );
and \g453948/U$2 ( \24951 , \16368 , RIe14e908_2271);
and \g453948/U$3 ( \24952 , RIfcd6160_7458, \16371 );
nor \g453948/U$1 ( \24953 , \24951 , \24952 );
nand \g448124/U$1 ( \24954 , \24940 , \24947 , \24950 , \24953 );
nor \g446458/U$1 ( \24955 , \24935 , \24936 , \24954 );
and \g453940/U$2 ( \24956 , \16377 , RIe15f708_2463);
and \g453940/U$3 ( \24957 , RIe157008_2367, \16380 );
nor \g453940/U$1 ( \24958 , \24956 , \24957 );
and \g453938/U$2 ( \24959 , \16313 , RIfc779a8_6383);
and \g453938/U$3 ( \24960 , RIe162408_2495, \16321 );
nor \g453938/U$1 ( \24961 , \24959 , \24960 );
and \g445469/U$2 ( \24962 , \24955 , \24958 , \24961 );
nor \g445469/U$1 ( \24963 , \24962 , \16389 );
or \g444347/U$1 ( \24964 , \24845 , \24905 , \24934 , \24963 );
and \g446444/U$2 ( \24965 , RIfc5c9f0_6076, \16432 );
and \g446444/U$3 ( \24966 , RIfea76b8_8221, \16361 );
and \g449450/U$2 ( \24967 , RIdee2af0_1043, \16485 );
and \g449450/U$3 ( \24968 , \16356 , RIdee4878_1064);
and \g449450/U$4 ( \24969 , RIded7150_911, \16398 );
nor \g449450/U$1 ( \24970 , \24967 , \24968 , \24969 );
and \g454718/U$2 ( \24971 , \16317 , RIfcde6f8_7553);
and \g454718/U$3 ( \24972 , RIfc942b0_6708, \16325 );
nor \g454718/U$1 ( \24973 , \24971 , \24972 );
not \g450470/U$3 ( \24974 , \24973 );
not \g450470/U$4 ( \24975 , \16311 );
and \g450470/U$2 ( \24976 , \24974 , \24975 );
and \g450470/U$5 ( \24977 , \16339 , RIded95e0_937);
nor \g450470/U$1 ( \24978 , \24976 , \24977 );
and \g453893/U$2 ( \24979 , \16377 , RIfcde860_7554);
and \g453893/U$3 ( \24980 , RIfcd1138_7401, \16313 );
nor \g453893/U$1 ( \24981 , \24979 , \24980 );
and \g453896/U$2 ( \24982 , \16334 , RIdede8d8_996);
and \g453896/U$3 ( \24983 , RIdee0a98_1020, \16380 );
nor \g453896/U$1 ( \24984 , \24982 , \24983 );
nand \g447434/U$1 ( \24985 , \24970 , \24978 , \24981 , \24984 );
nor \g446444/U$1 ( \24986 , \24965 , \24966 , \24985 );
and \g453889/U$2 ( \24987 , \16364 , RIded5260_889);
and \g453889/U$3 ( \24988 , RIee21160_4835, \16368 );
nor \g453889/U$1 ( \24989 , \24987 , \24988 );
and \g453886/U$2 ( \24990 , \16371 , RIfcc8768_7303);
and \g453886/U$3 ( \24991 , RIee22240_4847, \16427 );
nor \g453886/U$1 ( \24992 , \24990 , \24991 );
and \g445461/U$2 ( \24993 , \24986 , \24989 , \24992 );
nor \g445461/U$1 ( \24994 , \24993 , \16909 );
and \g446450/U$2 ( \24995 , RIe143508_2143, \16448 );
and \g446450/U$3 ( \24996 , RIdf2c560_1881, \16371 );
and \g449455/U$2 ( \24997 , RIde96290_322, \16485 );
and \g449455/U$3 ( \24998 , \16356 , RIdeb4308_514);
and \g449455/U$4 ( \24999 , RIdee6fd8_1092, \16398 );
nor \g449455/U$1 ( \25000 , \24997 , \24998 , \24999 );
and \g454662/U$2 ( \25001 , \16317 , RIdecd808_802);
and \g454662/U$3 ( \25002 , RIded0508_834, \16325 );
nor \g454662/U$1 ( \25003 , \25001 , \25002 );
not \g450475/U$3 ( \25004 , \25003 );
not \g450475/U$4 ( \25005 , \16311 );
and \g450475/U$2 ( \25006 , \25004 , \25005 );
and \g450475/U$5 ( \25007 , \16341 , RIdf004d8_1380);
nor \g450475/U$1 ( \25008 , \25006 , \25007 );
and \g453912/U$2 ( \25009 , \16377 , RIdec7e08_738);
and \g453912/U$3 ( \25010 , RIdecab08_770, \16313 );
nor \g453912/U$1 ( \25011 , \25009 , \25010 );
and \g453913/U$2 ( \25012 , \16334 , RIe159d08_2399);
and \g453913/U$3 ( \25013 , RIe16df10_2628, \16380 );
nor \g453913/U$1 ( \25014 , \25012 , \25013 );
nand \g447435/U$1 ( \25015 , \25000 , \25008 , \25011 , \25014 );
nor \g446450/U$1 ( \25016 , \24995 , \24996 , \25015 );
and \g453905/U$2 ( \25017 , \16364 , RIdedbd40_965);
and \g453905/U$3 ( \25018 , RIdf1cde0_1705, \16368 );
nor \g453905/U$1 ( \25019 , \25017 , \25018 );
and \g453907/U$2 ( \25020 , \16361 , RIde7c1d8_195);
and \g453907/U$3 ( \25021 , RIdf37f00_2013, \16427 );
nor \g453907/U$1 ( \25022 , \25020 , \25021 );
and \g445464/U$2 ( \25023 , \25016 , \25019 , \25022 );
nor \g445464/U$1 ( \25024 , \25023 , \16586 );
or \g444168/U$1 ( \25025 , \24964 , \24994 , \25024 );
_DC \g45e3/U$1 ( \25026 , \25025 , \16652 );
and \g448669/U$2 ( \25027 , RIe2182f8_4565, \8412 );
and \g448669/U$3 ( \25028 , \8409 , RIe21dcf8_4629);
and \g448669/U$4 ( \25029 , RIe20cef8_4437, \8326 );
nor \g448669/U$1 ( \25030 , \25027 , \25028 , \25029 );
and \g451190/U$2 ( \25031 , \8356 , RIe20fbf8_4469);
and \g451190/U$3 ( \25032 , RIfe9d398_8133, \8359 );
nor \g451190/U$1 ( \25033 , \25031 , \25032 );
and \g454408/U$2 ( \25034 , \8313 , RIfcdb9f8_7521);
and \g454408/U$3 ( \25035 , RIe2128f8_4501, \8323 );
nor \g454408/U$1 ( \25036 , \25034 , \25035 );
not \g449698/U$3 ( \25037 , \25036 );
not \g449698/U$4 ( \25038 , \8347 );
and \g449698/U$2 ( \25039 , \25037 , \25038 );
and \g449698/U$5 ( \25040 , \8340 , RIfc41d08_5771);
nor \g449698/U$1 ( \25041 , \25039 , \25040 );
and \g451189/U$2 ( \25042 , \8378 , RIe2155f8_4533);
and \g451189/U$3 ( \25043 , RIf16ad68_5675, \8417 );
nor \g451189/U$1 ( \25044 , \25042 , \25043 );
nand \g447556/U$1 ( \25045 , \25030 , \25033 , \25041 , \25044 );
and \g444760/U$2 ( \25046 , \25045 , \8369 );
and \g445840/U$2 ( \25047 , RIfe9d230_8132, \8371 );
and \g445840/U$3 ( \25048 , RIf166010_5620, \8383 );
and \g448673/U$2 ( \25049 , RIfc41a38_5769, \8412 );
and \g448673/U$3 ( \25050 , \8409 , RIfc41ba0_5770);
and \g448673/U$4 ( \25051 , RIfcbf258_7197, \8326 );
nor \g448673/U$1 ( \25052 , \25049 , \25050 , \25051 );
and \g451199/U$2 ( \25053 , \8356 , RIfec4560_8354);
and \g451199/U$3 ( \25054 , RIfc418d0_5768, \8359 );
nor \g451199/U$1 ( \25055 , \25053 , \25054 );
and \g454572/U$2 ( \25056 , \8313 , RIe1fcad0_4252);
and \g454572/U$3 ( \25057 , RIfc79190_6400, \8323 );
nor \g454572/U$1 ( \25058 , \25056 , \25057 );
not \g449701/U$3 ( \25059 , \25058 );
not \g449701/U$4 ( \25060 , \8347 );
and \g449701/U$2 ( \25061 , \25059 , \25060 );
and \g449701/U$5 ( \25062 , \8340 , RIfc79028_6399);
nor \g449701/U$1 ( \25063 , \25061 , \25062 );
and \g451198/U$2 ( \25064 , \8378 , RIfc92c30_6692);
and \g451198/U$3 ( \25065 , RIf165098_5609, \8417 );
nor \g451198/U$1 ( \25066 , \25064 , \25065 );
nand \g447557/U$1 ( \25067 , \25052 , \25055 , \25063 , \25066 );
nor \g445840/U$1 ( \25068 , \25047 , \25048 , \25067 );
and \g451194/U$2 ( \25069 , \8335 , RIfcd81b8_7481);
and \g451194/U$3 ( \25070 , RIfcd7510_7472, \8351 );
nor \g451194/U$1 ( \25071 , \25069 , \25070 );
and \g451195/U$2 ( \25072 , \8319 , RIfcc1df0_7228);
and \g451195/U$3 ( \25073 , RIe2008b0_4296, \8404 );
nor \g451195/U$1 ( \25074 , \25072 , \25073 );
and \g445032/U$2 ( \25075 , \25068 , \25071 , \25074 );
nor \g445032/U$1 ( \25076 , \25075 , \8422 );
nor \g444760/U$1 ( \25077 , \25046 , \25076 );
and \g446629/U$2 ( \25078 , \8426 , RIe2209f8_4661);
and \g446629/U$3 ( \25079 , RIfc795c8_6403, \8428 );
nor \g446629/U$1 ( \25080 , \25078 , \25079 );
and \g446628/U$2 ( \25081 , \13735 , RIe2236f8_4693);
and \g446628/U$3 ( \25082 , RIfc92960_6690, \13737 );
nor \g446628/U$1 ( \25083 , \25081 , \25082 );
and \g446630/U$2 ( \25084 , \8707 , RIe2074f8_4373);
and \g446630/U$3 ( \25085 , RIe20a1f8_4405, \8709 );
nor \g446630/U$1 ( \25086 , \25084 , \25085 );
nand \g444462/U$1 ( \25087 , \25077 , \25080 , \25083 , \25086 );
and \g451220/U$2 ( \25088 , \8319 , RIfcbf690_7200);
and \g451220/U$3 ( \25089 , RIe1fa0a0_4222, \8404 );
nor \g451220/U$1 ( \25090 , \25088 , \25089 );
and \g445844/U$2 ( \25091 , RIfcd77e0_7474, \8371 );
and \g445844/U$3 ( \25092 , RIfc5b4d8_6061, \8330 );
and \g448679/U$2 ( \25093 , RIf1546d0_5420, \8412 );
and \g448679/U$3 ( \25094 , \8409 , RIfe9d500_8134);
and \g448679/U$4 ( \25095 , RIfce8fb8_7673, \8326 );
nor \g448679/U$1 ( \25096 , \25093 , \25094 , \25095 );
and \g451224/U$2 ( \25097 , \8356 , RIe1f3020_4142);
and \g451224/U$3 ( \25098 , RIfec4830_8356, \8359 );
nor \g451224/U$1 ( \25099 , \25097 , \25098 );
and \g454425/U$2 ( \25100 , \8313 , RIf1508f0_5376);
and \g454425/U$3 ( \25101 , RIfec46c8_8355, \8323 );
nor \g454425/U$1 ( \25102 , \25100 , \25101 );
not \g449707/U$3 ( \25103 , \25102 );
not \g449707/U$4 ( \25104 , \8347 );
and \g449707/U$2 ( \25105 , \25103 , \25104 );
and \g449707/U$5 ( \25106 , \8340 , RIfce3180_7606);
nor \g449707/U$1 ( \25107 , \25105 , \25106 );
and \g451223/U$2 ( \25108 , \8378 , RIe1f5348_4167);
and \g451223/U$3 ( \25109 , RIf156188_5439, \8417 );
nor \g451223/U$1 ( \25110 , \25108 , \25109 );
nand \g447561/U$1 ( \25111 , \25096 , \25099 , \25107 , \25110 );
nor \g445844/U$1 ( \25112 , \25091 , \25092 , \25111 );
and \g451219/U$2 ( \25113 , \8335 , RIe1edd28_4083);
and \g451219/U$3 ( \25114 , RIfc92d98_6693, \8351 );
nor \g451219/U$1 ( \25115 , \25113 , \25114 );
nand \g445538/U$1 ( \25116 , \25090 , \25112 , \25115 );
and \g444841/U$2 ( \25117 , \25116 , \8752 );
and \g448676/U$2 ( \25118 , RIe1bb760_3510, \8326 );
and \g448676/U$3 ( \25119 , \8531 , RIe1f7c10_4196);
and \g448676/U$4 ( \25120 , RIe1fe858_4273, \8486 );
nor \g448676/U$1 ( \25121 , \25118 , \25119 , \25120 );
and \g451211/U$2 ( \25122 , \8356 , RIe1f0758_4113);
and \g451211/U$3 ( \25123 , RIe2047f8_4341, \8359 );
nor \g451211/U$1 ( \25124 , \25122 , \25123 );
and \g454651/U$2 ( \25125 , \8313 , RIe2263f8_4725);
and \g454651/U$3 ( \25126 , RIe178aa0_2750, \8323 );
nor \g454651/U$1 ( \25127 , \25125 , \25126 );
not \g449704/U$3 ( \25128 , \25127 );
not \g449704/U$4 ( \25129 , \8376 );
and \g449704/U$2 ( \25130 , \25128 , \25129 );
and \g449704/U$5 ( \25131 , \8340 , RIe1d4c60_3798);
nor \g449704/U$1 ( \25132 , \25130 , \25131 );
and \g451210/U$2 ( \25133 , \8378 , RIe21aff8_4597);
and \g451210/U$3 ( \25134 , RIe18c5a0_2974, \8417 );
nor \g451210/U$1 ( \25135 , \25133 , \25134 );
nand \g447560/U$1 ( \25136 , \25121 , \25124 , \25132 , \25135 );
and \g444841/U$3 ( \25137 , \9010 , \25136 );
nor \g444841/U$1 ( \25138 , \25117 , \25137 );
and \g446635/U$2 ( \25139 , \9041 , RIe1a00a0_3198);
and \g446635/U$3 ( \25140 , RIe1a2da0_3230, \9043 );
nor \g446635/U$1 ( \25141 , \25139 , \25140 );
and \g446634/U$2 ( \25142 , \14956 , RIe1a5aa0_3262);
and \g446634/U$3 ( \25143 , RIe1a87a0_3294, \14958 );
nor \g446634/U$1 ( \25144 , \25142 , \25143 );
and \g446636/U$2 ( \25145 , \13244 , RIe170c10_2660);
and \g446636/U$3 ( \25146 , RIe1ae5d8_3361, \13246 );
nor \g446636/U$1 ( \25147 , \25145 , \25146 );
nand \g444569/U$1 ( \25148 , \25138 , \25141 , \25144 , \25147 );
and \g445833/U$2 ( \25149 , RIfcb2c10_7056, \8373 );
and \g445833/U$3 ( \25150 , RIe19a6a0_3134, \8383 );
and \g448664/U$2 ( \25151 , RIe1811a0_2846, \8324 );
and \g448664/U$3 ( \25152 , \8523 , RIfc422a8_5775);
and \g448664/U$4 ( \25153 , RIe186ba0_2910, \8488 );
nor \g448664/U$1 ( \25154 , \25151 , \25152 , \25153 );
and \g451167/U$2 ( \25155 , \8356 , RIe183ea0_2878);
and \g451167/U$3 ( \25156 , RIe1898a0_2942, \8359 );
nor \g451167/U$1 ( \25157 , \25155 , \25156 );
and \g454318/U$2 ( \25158 , \8313 , RIe191fa0_3038);
and \g454318/U$3 ( \25159 , RIe194ca0_3070, \8323 );
nor \g454318/U$1 ( \25160 , \25158 , \25159 );
not \g449691/U$3 ( \25161 , \25160 );
not \g449691/U$4 ( \25162 , \8376 );
and \g449691/U$2 ( \25163 , \25161 , \25162 );
and \g449691/U$5 ( \25164 , \8340 , RIfcbecb8_7193);
nor \g449691/U$1 ( \25165 , \25163 , \25164 );
and \g451166/U$2 ( \25166 , \8378 , RIe18f2a0_3006);
and \g451166/U$3 ( \25167 , RIfc923c0_6686, \8417 );
nor \g451166/U$1 ( \25168 , \25166 , \25167 );
nand \g447554/U$1 ( \25169 , \25154 , \25157 , \25165 , \25168 );
nor \g445833/U$1 ( \25170 , \25149 , \25150 , \25169 );
and \g451162/U$2 ( \25171 , \8335 , RIe17b7a0_2782);
and \g451162/U$3 ( \25172 , RIe19d3a0_3166, \8351 );
nor \g451162/U$1 ( \25173 , \25171 , \25172 );
and \g451163/U$2 ( \25174 , \8317 , RIe17e4a0_2814);
and \g451163/U$3 ( \25175 , RIe1979a0_3102, \8404 );
nor \g451163/U$1 ( \25176 , \25174 , \25175 );
and \g445025/U$2 ( \25177 , \25170 , \25173 , \25176 );
nor \g445025/U$1 ( \25178 , \25177 , \8589 );
and \g445836/U$2 ( \25179 , RIfec43f8_8353, \8371 );
and \g445836/U$3 ( \25180 , RIf140bd0_5196, \8383 );
and \g448666/U$2 ( \25181 , RIfcd7678_7473, \8326 );
and \g448666/U$3 ( \25182 , \8523 , RIfc79898_6405);
and \g448666/U$4 ( \25183 , RIfcea200_7686, \8488 );
nor \g448666/U$1 ( \25184 , \25181 , \25182 , \25183 );
and \g451179/U$2 ( \25185 , \8356 , RIe1734d8_2689);
and \g451179/U$3 ( \25186 , RIfcd8320_7482, \8359 );
nor \g451179/U$1 ( \25187 , \25185 , \25186 );
and \g454754/U$2 ( \25188 , \8313 , RIfc92528_6687);
and \g454754/U$3 ( \25189 , RIf13efb0_5176, \8323 );
nor \g454754/U$1 ( \25190 , \25188 , \25189 );
not \g449694/U$3 ( \25191 , \25190 );
not \g449694/U$4 ( \25192 , \8376 );
and \g449694/U$2 ( \25193 , \25191 , \25192 );
and \g449694/U$5 ( \25194 , \8340 , RIfcd7948_7475);
nor \g449694/U$1 ( \25195 , \25193 , \25194 );
and \g451176/U$2 ( \25196 , \8378 , RIfcb2aa8_7055);
and \g451176/U$3 ( \25197 , RIfc79b68_6407, \8417 );
nor \g451176/U$1 ( \25198 , \25196 , \25197 );
nand \g447555/U$1 ( \25199 , \25184 , \25187 , \25195 , \25198 );
nor \g445836/U$1 ( \25200 , \25179 , \25180 , \25199 );
and \g451172/U$2 ( \25201 , \8335 , RIfc927f8_6689);
and \g451172/U$3 ( \25202 , RIf142250_5212, \8351 );
nor \g451172/U$1 ( \25203 , \25201 , \25202 );
and \g451175/U$2 ( \25204 , \8319 , RIf16e170_5712);
and \g451175/U$3 ( \25205 , RIe175968_2715, \8404 );
nor \g451175/U$1 ( \25206 , \25204 , \25205 );
and \g445027/U$2 ( \25207 , \25200 , \25203 , \25206 );
nor \g445027/U$1 ( \25208 , \25207 , \8558 );
or \g444386/U$1 ( \25209 , \25087 , \25148 , \25178 , \25208 );
and \g445829/U$2 ( \25210 , RIe1da660_3862, \8414 );
and \g445829/U$3 ( \25211 , RIe1c9860_3670, \8356 );
and \g448656/U$2 ( \25212 , RIe1c1160_3574, \8319 );
and \g448656/U$3 ( \25213 , \8324 , RIe1c3e60_3606);
and \g448656/U$4 ( \25214 , RIe1dd360_3894, \8409 );
nor \g448656/U$1 ( \25215 , \25212 , \25213 , \25214 );
and \g451141/U$2 ( \25216 , \8335 , RIe1be460_3542);
and \g451141/U$3 ( \25217 , RIe1c6b60_3638, \8340 );
nor \g451141/U$1 ( \25218 , \25216 , \25217 );
and \g451140/U$2 ( \25219 , \8404 , RIe1e2d60_3958);
and \g451140/U$3 ( \25220 , RIe1eb460_4054, \8351 );
nor \g451140/U$1 ( \25221 , \25219 , \25220 );
and \g454969/U$2 ( \25222 , \8313 , RIe1e5a60_3990);
and \g454969/U$3 ( \25223 , RIe1e8760_4022, \8323 );
nor \g454969/U$1 ( \25224 , \25222 , \25223 );
not \g449681/U$3 ( \25225 , \25224 );
not \g449681/U$4 ( \25226 , \8328 );
and \g449681/U$2 ( \25227 , \25225 , \25226 );
and \g449681/U$5 ( \25228 , \8417 , RIe1e0060_3926);
nor \g449681/U$1 ( \25229 , \25227 , \25228 );
nand \g447548/U$1 ( \25230 , \25215 , \25218 , \25221 , \25229 );
nor \g445829/U$1 ( \25231 , \25210 , \25211 , \25230 );
and \g451135/U$2 ( \25232 , \8378 , RIe1d7960_3830);
and \g451135/U$3 ( \25233 , RIe1d1f60_3766, \8359 );
nor \g451135/U$1 ( \25234 , \25232 , \25233 );
and \g451134/U$2 ( \25235 , \8531 , RIe1cc560_3702);
and \g451134/U$3 ( \25236 , RIe1cf260_3734, \8486 );
nor \g451134/U$1 ( \25237 , \25235 , \25236 );
and \g445022/U$2 ( \25238 , \25231 , \25234 , \25237 );
nor \g445022/U$1 ( \25239 , \25238 , \8477 );
and \g445832/U$2 ( \25240 , RIfe9cf60_8130, \8414 );
and \g445832/U$3 ( \25241 , RIfe9cdf8_8129, \8356 );
and \g448659/U$2 ( \25242 , RIe1ac2b0_3336, \8319 );
and \g448659/U$3 ( \25243 , \8324 , RIf146468_5259);
and \g448659/U$4 ( \25244 , RIfe9cb28_8127, \8409 );
nor \g448659/U$1 ( \25245 , \25242 , \25243 , \25244 );
and \g451155/U$2 ( \25246 , \8335 , RIe1aaac8_3319);
and \g451155/U$3 ( \25247 , RIf147110_5268, \8340 );
nor \g451155/U$1 ( \25248 , \25246 , \25247 );
and \g451154/U$2 ( \25249 , \8404 , RIe1b7110_3460);
and \g451154/U$3 ( \25250 , RIfe9d0c8_8131, \8351 );
nor \g451154/U$1 ( \25251 , \25249 , \25250 );
and \g454883/U$2 ( \25252 , \8313 , RIe1b9168_3483);
and \g454883/U$3 ( \25253 , RIfe9cc90_8128, \8323 );
nor \g454883/U$1 ( \25254 , \25252 , \25253 );
not \g449686/U$3 ( \25255 , \25254 );
not \g449686/U$4 ( \25256 , \8328 );
and \g449686/U$2 ( \25257 , \25255 , \25256 );
and \g449686/U$5 ( \25258 , \8417 , RIf14a3b0_5304);
nor \g449686/U$1 ( \25259 , \25257 , \25258 );
nand \g447550/U$1 ( \25260 , \25245 , \25248 , \25251 , \25259 );
nor \g445832/U$1 ( \25261 , \25240 , \25241 , \25260 );
and \g451151/U$2 ( \25262 , \8378 , RIfe9c9c0_8126);
and \g451151/U$3 ( \25263 , RIfce2208_7595, \8359 );
nor \g451151/U$1 ( \25264 , \25262 , \25263 );
and \g451149/U$2 ( \25265 , \8531 , RIfe9c858_8125);
and \g451149/U$3 ( \25266 , RIfce9558_7677, \8486 );
nor \g451149/U$1 ( \25267 , \25265 , \25266 );
and \g445024/U$2 ( \25268 , \25261 , \25264 , \25267 );
nor \g445024/U$1 ( \25269 , \25268 , \8481 );
or \g444195/U$1 ( \25270 , \25209 , \25239 , \25269 );
_DC \g4667/U$1 ( \25271 , \25270 , \8654 );
and \g448931/U$2 ( \25272 , RIdeb2580_493, \16427 );
and \g448931/U$3 ( \25273 , \16448 , RIfcbe448_7187);
and \g448931/U$4 ( \25274 , RIdec3380_685, \16321 );
nor \g448931/U$1 ( \25275 , \25272 , \25273 , \25274 );
and \g452009/U$2 ( \25276 , \16368 , RIdeaf880_461);
and \g452009/U$3 ( \25277 , RIfcb3480_7062, \16371 );
nor \g452009/U$1 ( \25278 , \25276 , \25277 );
and \g455402/U$2 ( \25279 , \16317 , RIdebd980_621);
and \g455402/U$3 ( \25280 , RIfcd70d8_7469, \16325 );
nor \g455402/U$1 ( \25281 , \25279 , \25280 );
not \g450356/U$3 ( \25282 , \25281 );
not \g450356/U$4 ( \25283 , \16330 );
and \g450356/U$2 ( \25284 , \25282 , \25283 );
and \g450356/U$5 ( \25285 , \16328 , RIdec6080_717);
nor \g450356/U$1 ( \25286 , \25284 , \25285 );
and \g452007/U$2 ( \25287 , \16334 , RIdeb7f80_557);
and \g452007/U$3 ( \25288 , RIdebac80_589, \16380 );
nor \g452007/U$1 ( \25289 , \25287 , \25288 );
nand \g447687/U$1 ( \25290 , \25275 , \25278 , \25286 , \25289 );
and \g444706/U$2 ( \25291 , \25290 , \17938 );
and \g446043/U$2 ( \25292 , RIfc5a560_6050, \16313 );
and \g446043/U$3 ( \25293 , RIdf2fda0_1921, \16361 );
and \g448937/U$2 ( \25294 , RIfc7a270_6412, \16321 );
and \g448937/U$3 ( \25295 , \16485 , RIe13f5c0_2098);
and \g448937/U$4 ( \25296 , RIfea6fb0_8216, \16356 );
nor \g448937/U$1 ( \25297 , \25294 , \25295 , \25296 );
and \g452022/U$2 ( \25298 , \16368 , RIee2d910_4977);
and \g452022/U$3 ( \25299 , RIfc91cb8_6681, \16371 );
nor \g452022/U$1 ( \25300 , \25298 , \25299 );
and \g454933/U$2 ( \25301 , \16317 , RIee2fc38_5002);
and \g454933/U$3 ( \25302 , RIfce5bb0_7636, \16325 );
nor \g454933/U$1 ( \25303 , \25301 , \25302 );
not \g449950/U$3 ( \25304 , \25303 );
not \g449950/U$4 ( \25305 , \16351 );
and \g449950/U$2 ( \25306 , \25304 , \25305 );
and \g449950/U$5 ( \25307 , \16328 , RIfc42b18_5781);
nor \g449950/U$1 ( \25308 , \25306 , \25307 );
and \g453112/U$2 ( \25309 , \16334 , RIdf3b038_2048);
and \g453112/U$3 ( \25310 , RIdf3d4c8_2074, \16380 );
nor \g453112/U$1 ( \25311 , \25309 , \25310 );
nand \g447692/U$1 ( \25312 , \25297 , \25300 , \25308 , \25311 );
nor \g446043/U$1 ( \25313 , \25292 , \25293 , \25312 );
and \g452018/U$2 ( \25314 , \16364 , RIdf31c90_1943);
and \g452018/U$3 ( \25315 , RIdf362e0_1993, \16341 );
nor \g452018/U$1 ( \25316 , \25314 , \25315 );
and \g453551/U$2 ( \25317 , \16337 , RIdf33e50_1967);
and \g453551/U$3 ( \25318 , RIfc96b78_6737, \16377 );
nor \g453551/U$1 ( \25319 , \25317 , \25318 );
and \g445181/U$2 ( \25320 , \25313 , \25316 , \25319 );
nor \g445181/U$1 ( \25321 , \25320 , \16393 );
nor \g444706/U$1 ( \25322 , \25291 , \25321 );
and \g446820/U$2 ( \25323 , \18776 , RIdec0680_653);
and \g446820/U$3 ( \25324 , RIee204b8_4826, \18778 );
nor \g446820/U$1 ( \25325 , \25323 , \25324 );
and \g446821/U$2 ( \25326 , \18781 , RIdeac1a8_429);
and \g446821/U$3 ( \25327 , RIfc43928_5791, \18783 );
nor \g446821/U$1 ( \25328 , \25326 , \25327 );
and \g446822/U$2 ( \25329 , \18467 , RIde9efa8_365);
and \g446822/U$3 ( \25330 , RIdea58a8_397, \18469 );
nor \g446822/U$1 ( \25331 , \25329 , \25330 );
nand \g444487/U$1 ( \25332 , \25322 , \25325 , \25328 , \25331 );
and \g452041/U$2 ( \25333 , \16368 , RIdef6050_1263);
and \g452041/U$3 ( \25334 , RIdf09b50_1487, \16485 );
nor \g452041/U$1 ( \25335 , \25333 , \25334 );
and \g446048/U$2 ( \25336 , RIdf0c850_1519, \16356 );
and \g446048/U$3 ( \25337 , RIdf04150_1423, \16334 );
and \g448944/U$2 ( \25338 , RIdf14f50_1615, \16321 );
and \g448944/U$3 ( \25339 , \16326 , RIdf17c50_1647);
and \g448944/U$4 ( \25340 , RIdefba50_1327, \16427 );
nor \g448944/U$1 ( \25341 , \25338 , \25339 , \25340 );
and \g452048/U$2 ( \25342 , \16361 , RIdeeac50_1135);
and \g452048/U$3 ( \25343 , RIdeed950_1167, \16364 );
nor \g452048/U$1 ( \25344 , \25342 , \25343 );
and \g452046/U$2 ( \25345 , \16377 , RIdf0f550_1551);
and \g452046/U$3 ( \25346 , RIdf12250_1583, \16313 );
nor \g452046/U$1 ( \25347 , \25345 , \25346 );
and \g455136/U$2 ( \25348 , \16317 , RIdef0650_1199);
and \g455136/U$3 ( \25349 , RIdef3350_1231, \16325 );
nor \g455136/U$1 ( \25350 , \25348 , \25349 );
not \g455135/U$1 ( \25351 , \25350 );
and \g449960/U$2 ( \25352 , \25351 , \16336 );
and \g449960/U$3 ( \25353 , RIdefe750_1359, \16448 );
nor \g449960/U$1 ( \25354 , \25352 , \25353 );
nand \g448063/U$1 ( \25355 , \25341 , \25344 , \25347 , \25354 );
nor \g446048/U$1 ( \25356 , \25336 , \25337 , \25355 );
and \g452040/U$2 ( \25357 , \16371 , RIdef8d50_1295);
and \g452040/U$3 ( \25358 , RIdf06e50_1455, \16380 );
nor \g452040/U$1 ( \25359 , \25357 , \25358 );
nand \g445586/U$1 ( \25360 , \25335 , \25356 , \25359 );
and \g444772/U$2 ( \25361 , \25360 , \16750 );
and \g448939/U$2 ( \25362 , RIfcb3318_7061, \16427 );
and \g448939/U$3 ( \25363 , \16398 , RIdf20350_1743);
and \g448939/U$4 ( \25364 , RIfc430b8_5785, \16341 );
nor \g448939/U$1 ( \25365 , \25362 , \25363 , \25364 );
and \g451480/U$2 ( \25366 , \16361 , RIdf19e10_1671);
and \g451480/U$3 ( \25367 , RIfc7a978_6417, \16364 );
nor \g451480/U$1 ( \25368 , \25366 , \25367 );
and \g451724/U$2 ( \25369 , \16377 , RIfc7ac48_6419);
and \g451724/U$3 ( \25370 , RIfc96fb0_6740, \16313 );
nor \g451724/U$1 ( \25371 , \25369 , \25370 );
and \g455152/U$2 ( \25372 , \16317 , RIfc59e58_6045);
and \g455152/U$3 ( \25373 , RIfc43658_5789, \16325 );
nor \g455152/U$1 ( \25374 , \25372 , \25373 );
not \g449954/U$3 ( \25375 , \25374 );
not \g449954/U$4 ( \25376 , \16311 );
and \g449954/U$2 ( \25377 , \25375 , \25376 );
and \g449954/U$5 ( \25378 , \16448 , RIfc91718_6677);
nor \g449954/U$1 ( \25379 , \25377 , \25378 );
nand \g447696/U$1 ( \25380 , \25365 , \25368 , \25371 , \25379 );
and \g444772/U$3 ( \25381 , \16481 , \25380 );
nor \g444772/U$1 ( \25382 , \25361 , \25381 );
and \g446834/U$2 ( \25383 , \16511 , RIdf25210_1799);
and \g446834/U$3 ( \25384 , RIdf26cc8_1818, \16514 );
nor \g446834/U$1 ( \25385 , \25383 , \25384 );
and \g446829/U$2 ( \25386 , \24165 , RIdf28bb8_1840);
and \g446829/U$3 ( \25387 , RIfea0368_8167, \24167 );
nor \g446829/U$1 ( \25388 , \25386 , \25387 );
and \g446830/U$2 ( \25389 , \17279 , RIfc91880_6678);
and \g446830/U$3 ( \25390 , RIfc919e8_6679, \17281 );
nor \g446830/U$1 ( \25391 , \25389 , \25390 );
nand \g444489/U$1 ( \25392 , \25382 , \25385 , \25388 , \25391 );
and \g446032/U$2 ( \25393 , RIfea99e0_8246, \16356 );
and \g446032/U$3 ( \25394 , RIdedf2b0_1003, \16334 );
and \g448921/U$2 ( \25395 , RIfc968a8_6735, \16321 );
and \g448921/U$3 ( \25396 , \16326 , RIfcd1b10_7408);
and \g448921/U$4 ( \25397 , RIfcd85f0_7484, \16427 );
nor \g448921/U$1 ( \25398 , \25395 , \25396 , \25397 );
and \g451981/U$2 ( \25399 , \16361 , RIded37a8_870);
and \g451981/U$3 ( \25400 , RIded5f08_898, \16364 );
nor \g451981/U$1 ( \25401 , \25399 , \25400 );
and \g451980/U$2 ( \25402 , \16377 , RIfcdfc10_7568);
and \g451980/U$3 ( \25403 , RIfc91f88_6683, \16313 );
nor \g451980/U$1 ( \25404 , \25402 , \25403 );
and \g454190/U$2 ( \25405 , \16317 , RIfea9878_8245);
and \g454190/U$3 ( \25406 , RIdeda3f0_947, \16325 );
nor \g454190/U$1 ( \25407 , \25405 , \25406 );
not \g454189/U$1 ( \25408 , \25407 );
and \g449937/U$2 ( \25409 , \25408 , \16336 );
and \g449937/U$3 ( \25410 , RIfcc7d90_7296, \16448 );
nor \g449937/U$1 ( \25411 , \25409 , \25410 );
nand \g448061/U$1 ( \25412 , \25398 , \25401 , \25404 , \25411 );
nor \g446032/U$1 ( \25413 , \25393 , \25394 , \25412 );
and \g451973/U$2 ( \25414 , \16371 , RIfce3888_7611);
and \g451973/U$3 ( \25415 , RIdee1308_1026, \16380 );
nor \g451973/U$1 ( \25416 , \25414 , \25415 );
and \g451974/U$2 ( \25417 , \16368 , RIfc5a830_6052);
and \g451974/U$3 ( \25418 , RIdee3630_1051, \16485 );
nor \g451974/U$1 ( \25419 , \25417 , \25418 );
and \g445174/U$2 ( \25420 , \25413 , \25416 , \25419 );
nor \g445174/U$1 ( \25421 , \25420 , \16909 );
and \g446035/U$2 ( \25422 , RIdeb5280_525, \16356 );
and \g446035/U$3 ( \25423 , RIe15ac80_2410, \16334 );
and \g448926/U$2 ( \25424 , RIdf38e78_2024, \16427 );
and \g448926/U$3 ( \25425 , \16398 , RIdee7f50_1103);
and \g448926/U$4 ( \25426 , RIdf01450_1391, \16341 );
nor \g448926/U$1 ( \25427 , \25424 , \25425 , \25426 );
and \g451995/U$2 ( \25428 , \16361 , RIde7e5f0_206);
and \g451995/U$3 ( \25429 , RIdedccb8_976, \16364 );
nor \g451995/U$1 ( \25430 , \25428 , \25429 );
and \g451993/U$2 ( \25431 , \16377 , RIdec8d80_749);
and \g451993/U$3 ( \25432 , RIdecba80_781, \16313 );
nor \g451993/U$1 ( \25433 , \25431 , \25432 );
and \g454723/U$2 ( \25434 , \16317 , RIdece780_813);
and \g454723/U$3 ( \25435 , RIded1480_845, \16325 );
nor \g454723/U$1 ( \25436 , \25434 , \25435 );
not \g449941/U$3 ( \25437 , \25436 );
not \g449941/U$4 ( \25438 , \16311 );
and \g449941/U$2 ( \25439 , \25437 , \25438 );
and \g449941/U$5 ( \25440 , \16448 , RIe144480_2154);
nor \g449941/U$1 ( \25441 , \25439 , \25440 );
nand \g447684/U$1 ( \25442 , \25427 , \25430 , \25433 , \25441 );
nor \g446035/U$1 ( \25443 , \25422 , \25423 , \25442 );
and \g451987/U$2 ( \25444 , \16371 , RIdf2d4d8_1892);
and \g451987/U$3 ( \25445 , RIe16ee88_2639, \16380 );
nor \g451987/U$1 ( \25446 , \25444 , \25445 );
and \g451989/U$2 ( \25447 , \16368 , RIdf1dd58_1716);
and \g451989/U$3 ( \25448 , RIde986a8_333, \16485 );
nor \g451989/U$1 ( \25449 , \25447 , \25448 );
and \g445176/U$2 ( \25450 , \25443 , \25446 , \25449 );
nor \g445176/U$1 ( \25451 , \25450 , \16586 );
or \g444317/U$1 ( \25452 , \25332 , \25392 , \25421 , \25451 );
and \g446024/U$2 ( \25453 , RIfcc77f0_7292, \16313 );
and \g446024/U$3 ( \25454 , RIe168948_2567, \16361 );
and \g448913/U$2 ( \25455 , RIee1c408_4780, \16321 );
and \g448913/U$3 ( \25456 , \16344 , RIde8ec70_286);
and \g448913/U$4 ( \25457 , RIde92438_303, \16356 );
nor \g448913/U$1 ( \25458 , \25455 , \25456 , \25457 );
and \g451954/U$2 ( \25459 , \16368 , RIfc91448_6675);
and \g451954/U$3 ( \25460 , RIfcd1de0_7410, \16371 );
nor \g451954/U$1 ( \25461 , \25459 , \25460 );
and \g454474/U$2 ( \25462 , \16317 , RIfc59a20_6042);
and \g454474/U$3 ( \25463 , RIfca31c0_6878, \16325 );
nor \g454474/U$1 ( \25464 , \25462 , \25463 );
not \g449931/U$3 ( \25465 , \25464 );
not \g449931/U$4 ( \25466 , \16351 );
and \g449931/U$2 ( \25467 , \25465 , \25466 );
and \g449931/U$5 ( \25468 , \16326 , RIfcd88c0_7486);
nor \g449931/U$1 ( \25469 , \25467 , \25468 );
and \g451952/U$2 ( \25470 , \16334 , RIde86930_246);
and \g451952/U$3 ( \25471 , RIde8aad0_266, \16380 );
nor \g451952/U$1 ( \25472 , \25470 , \25471 );
nand \g447675/U$1 ( \25473 , \25458 , \25461 , \25469 , \25472 );
nor \g446024/U$1 ( \25474 , \25453 , \25454 , \25473 );
and \g451948/U$2 ( \25475 , \16364 , RIfc97118_6741);
and \g451948/U$3 ( \25476 , RIfc97280_6742, \16339 );
nor \g451948/U$1 ( \25477 , \25475 , \25476 );
and \g451946/U$2 ( \25478 , \16398 , RIe16c188_2607);
and \g451946/U$3 ( \25479 , RIfea04d0_8168, \16377 );
nor \g451946/U$1 ( \25480 , \25478 , \25479 );
and \g445166/U$2 ( \25481 , \25474 , \25477 , \25480 );
nor \g445166/U$1 ( \25482 , \25481 , \16649 );
and \g446028/U$2 ( \25483 , RIfcd1c78_7409, \16356 );
and \g446028/U$3 ( \25484 , RIe155280_2346, \16334 );
and \g448918/U$2 ( \25485 , RIe152580_2314, \16427 );
and \g448918/U$3 ( \25486 , \16398 , RIe14cb80_2250);
and \g448918/U$4 ( \25487 , RIfc7a3d8_6413, \16341 );
nor \g448918/U$1 ( \25488 , \25485 , \25486 , \25487 );
and \g451967/U$2 ( \25489 , \16361 , RIe147180_2186);
and \g451967/U$3 ( \25490 , RIe149e80_2218, \16364 );
nor \g451967/U$1 ( \25491 , \25489 , \25490 );
and \g451966/U$2 ( \25492 , \16377 , RIe160680_2474);
and \g451966/U$3 ( \25493 , RIee37ac8_5092, \16313 );
nor \g451966/U$1 ( \25494 , \25492 , \25493 );
and \g454694/U$2 ( \25495 , \16317 , RIe163380_2506);
and \g454694/U$3 ( \25496 , RIe166080_2538, \16325 );
nor \g454694/U$1 ( \25497 , \25495 , \25496 );
not \g449934/U$3 ( \25498 , \25497 );
not \g449934/U$4 ( \25499 , \16311 );
and \g449934/U$2 ( \25500 , \25498 , \25499 );
and \g449934/U$5 ( \25501 , \16448 , RIfc3f530_5746);
nor \g449934/U$1 ( \25502 , \25500 , \25501 );
nand \g447678/U$1 ( \25503 , \25488 , \25491 , \25494 , \25502 );
nor \g446028/U$1 ( \25504 , \25483 , \25484 , \25503 );
and \g451090/U$2 ( \25505 , \16371 , RIee35368_5064);
and \g451090/U$3 ( \25506 , RIe157f80_2378, \16380 );
nor \g451090/U$1 ( \25507 , \25505 , \25506 );
and \g451963/U$2 ( \25508 , \16368 , RIe14f880_2282);
and \g451963/U$3 ( \25509 , RIe15d980_2442, \16344 );
nor \g451963/U$1 ( \25510 , \25508 , \25509 );
and \g445171/U$2 ( \25511 , \25504 , \25507 , \25510 );
nor \g445171/U$1 ( \25512 , \25511 , \16389 );
or \g444213/U$1 ( \25513 , \25452 , \25482 , \25512 );
_DC \g46ec/U$1 ( \25514 , \25513 , \16652 );
and \g446901/U$2 ( \25515 , \10230 , RIe1fc0f8_4245);
and \g446901/U$3 ( \25516 , RIfe9ff30_8164, \10232 );
nor \g446901/U$1 ( \25517 , \25515 , \25516 );
and \g446131/U$2 ( \25518 , RIfcc27c8_7235, \8417 );
and \g446131/U$3 ( \25519 , RIfcdfee0_7570, \8409 );
and \g449046/U$2 ( \25520 , RIfcd8cf8_7489, \8319 );
and \g449046/U$3 ( \25521 , \8326 , RIf15bb88_5503);
and \g449046/U$4 ( \25522 , RIf15e9f0_5536, \8488 );
nor \g449046/U$1 ( \25523 , \25520 , \25521 , \25522 );
and \g452401/U$2 ( \25524 , \8335 , RIfcd8e60_7490);
and \g452401/U$3 ( \25525 , RIfc7be90_6432, \8340 );
nor \g452401/U$1 ( \25526 , \25524 , \25525 );
and \g452399/U$2 ( \25527 , \8404 , RIe201288_4303);
and \g452399/U$3 ( \25528 , RIfc8fc60_6658, \8351 );
nor \g452399/U$1 ( \25529 , \25527 , \25528 );
and \g454837/U$2 ( \25530 , \8313 , RIe202ea8_4323);
and \g454837/U$3 ( \25531 , RIfc97820_6746, \8323 );
nor \g454837/U$1 ( \25532 , \25530 , \25531 );
not \g450060/U$3 ( \25533 , \25532 );
not \g450060/U$4 ( \25534 , \8328 );
and \g450060/U$2 ( \25535 , \25533 , \25534 );
and \g450060/U$5 ( \25536 , \8359 , RIf1608e0_5558);
nor \g450060/U$1 ( \25537 , \25535 , \25536 );
nand \g447748/U$1 ( \25538 , \25523 , \25526 , \25529 , \25537 );
nor \g446131/U$1 ( \25539 , \25518 , \25519 , \25538 );
not \g444869/U$3 ( \25540 , \25539 );
not \g444869/U$4 ( \25541 , \8422 );
and \g444869/U$2 ( \25542 , \25540 , \25541 );
and \g446132/U$2 ( \25543 , RIfc58508_6027, \8417 );
and \g446132/U$3 ( \25544 , RIe210b70_4480, \8356 );
and \g449048/U$2 ( \25545 , RIe20b170_4416, \8319 );
and \g449048/U$3 ( \25546 , \8326 , RIe20de70_4448);
and \g449048/U$4 ( \25547 , RIe213870_4512, \8486 );
nor \g449048/U$1 ( \25548 , \25545 , \25546 , \25547 );
and \g452409/U$2 ( \25549 , \8335 , RIe208470_4384);
and \g452409/U$3 ( \25550 , RIfc58940_6030, \8340 );
nor \g452409/U$1 ( \25551 , \25549 , \25550 );
and \g452408/U$2 ( \25552 , \8404 , RIe221970_4672);
and \g452408/U$3 ( \25553 , RIf16cdc0_5698, \8351 );
nor \g452408/U$1 ( \25554 , \25552 , \25553 );
and \g454839/U$2 ( \25555 , \8313 , RIf16c118_5689);
and \g454839/U$3 ( \25556 , RIe224670_4704, \8323 );
nor \g454839/U$1 ( \25557 , \25555 , \25556 );
not \g450063/U$3 ( \25558 , \25557 );
not \g450063/U$4 ( \25559 , \8328 );
and \g450063/U$2 ( \25560 , \25558 , \25559 );
and \g450063/U$5 ( \25561 , \8359 , RIfc3ff08_5753);
nor \g450063/U$1 ( \25562 , \25560 , \25561 );
nand \g447749/U$1 ( \25563 , \25548 , \25551 , \25554 , \25562 );
nor \g446132/U$1 ( \25564 , \25543 , \25544 , \25563 );
and \g452406/U$2 ( \25565 , \8378 , RIe216570_4544);
and \g452406/U$3 ( \25566 , RIf1696e8_5659, \8531 );
nor \g452406/U$1 ( \25567 , \25565 , \25566 );
and \g452405/U$2 ( \25568 , \8414 , RIe219270_4576);
and \g452405/U$3 ( \25569 , RIe21ec70_4640, \8409 );
nor \g452405/U$1 ( \25570 , \25568 , \25569 );
and \g445243/U$2 ( \25571 , \25564 , \25567 , \25570 );
nor \g445243/U$1 ( \25572 , \25571 , \8368 );
nor \g444869/U$1 ( \25573 , \25542 , \25572 );
and \g446902/U$2 ( \25574 , \14165 , RIfc58670_6028);
and \g446902/U$3 ( \25575 , RIfc44198_5797, \14167 );
nor \g446902/U$1 ( \25576 , \25574 , \25575 );
nand \g444428/U$1 ( \25577 , \25517 , \25573 , \25576 );
and \g452418/U$2 ( \25578 , \8319 , RIe1c20d8_3585);
and \g452418/U$3 ( \25579 , RIe1c4dd8_3617, \8324 );
nor \g452418/U$1 ( \25580 , \25578 , \25579 );
and \g446134/U$2 ( \25581 , RIe1c7ad8_3649, \8340 );
and \g446134/U$3 ( \25582 , RIe1e3cd8_3969, \8404 );
and \g449052/U$2 ( \25583 , RIe1db5d8_3873, \8414 );
and \g449052/U$3 ( \25584 , \8409 , RIe1de2d8_3905);
and \g449052/U$4 ( \25585 , RIe1e96d8_4033, \8330 );
nor \g449052/U$1 ( \25586 , \25583 , \25584 , \25585 );
and \g452421/U$2 ( \25587 , \8356 , RIe1ca7d8_3681);
and \g452421/U$3 ( \25588 , RIe1d2ed8_3777, \8359 );
nor \g452421/U$1 ( \25589 , \25587 , \25588 );
and \g454852/U$2 ( \25590 , \8313 , RIe1cd4d8_3713);
and \g454852/U$3 ( \25591 , RIe1d01d8_3745, \8323 );
nor \g454852/U$1 ( \25592 , \25590 , \25591 );
not \g450066/U$3 ( \25593 , \25592 );
not \g450066/U$4 ( \25594 , \8347 );
and \g450066/U$2 ( \25595 , \25593 , \25594 );
and \g450066/U$5 ( \25596 , \8351 , RIe1ec3d8_4065);
nor \g450066/U$1 ( \25597 , \25595 , \25596 );
and \g452420/U$2 ( \25598 , \8378 , RIe1d88d8_3841);
and \g452420/U$3 ( \25599 , RIe1e0fd8_3937, \8417 );
nor \g452420/U$1 ( \25600 , \25598 , \25599 );
nand \g447751/U$1 ( \25601 , \25586 , \25589 , \25597 , \25600 );
nor \g446134/U$1 ( \25602 , \25581 , \25582 , \25601 );
and \g452417/U$2 ( \25603 , \8335 , RIe1bf3d8_3553);
and \g452417/U$3 ( \25604 , RIe1e69d8_4001, \8373 );
nor \g452417/U$1 ( \25605 , \25603 , \25604 );
nand \g445608/U$1 ( \25606 , \25580 , \25602 , \25605 );
and \g444778/U$2 ( \25607 , \25606 , \8478 );
and \g449050/U$2 ( \25608 , RIe1b2ef8_3413, \8523 );
and \g449050/U$3 ( \25609 , \8486 , RIfcdfd78_7569);
and \g449050/U$4 ( \25610 , RIfce3cc0_7614, \8383 );
nor \g449050/U$1 ( \25611 , \25608 , \25609 , \25610 );
and \g452413/U$2 ( \25612 , \8356 , RIe1b15a8_3395);
and \g452413/U$3 ( \25613 , RIfc90bd8_6669, \8359 );
nor \g452413/U$1 ( \25614 , \25612 , \25613 );
and \g454848/U$2 ( \25615 , \8313 , RIe1b5a90_3444);
and \g454848/U$3 ( \25616 , RIf149e10_5300, \8323 );
nor \g454848/U$1 ( \25617 , \25615 , \25616 );
not \g450064/U$3 ( \25618 , \25617 );
not \g450064/U$4 ( \25619 , \8376 );
and \g450064/U$2 ( \25620 , \25618 , \25619 );
and \g450064/U$5 ( \25621 , \8351 , RIfcc73b8_7289);
nor \g450064/U$1 ( \25622 , \25620 , \25621 );
and \g452412/U$2 ( \25623 , \8378 , RIfea0200_8166);
and \g452412/U$3 ( \25624 , RIfcd6f70_7468, \8417 );
nor \g452412/U$1 ( \25625 , \25623 , \25624 );
nand \g447750/U$1 ( \25626 , \25611 , \25614 , \25622 , \25625 );
and \g444778/U$3 ( \25627 , \8482 , \25626 );
nor \g444778/U$1 ( \25628 , \25607 , \25627 );
and \g446906/U$2 ( \25629 , \8509 , RIe1ab608_3327);
and \g446906/U$3 ( \25630 , RIe1acdf0_3344, \8511 );
nor \g446906/U$1 ( \25631 , \25629 , \25630 );
and \g446905/U$2 ( \25632 , \8514 , RIfcc7520_7290);
and \g446905/U$3 ( \25633 , RIfc973e8_6743, \8517 );
nor \g446905/U$1 ( \25634 , \25632 , \25633 );
and \g446907/U$2 ( \25635 , \8969 , RIe1b7c50_3468);
and \g446907/U$3 ( \25636 , RIe1b9e10_3492, \8971 );
nor \g446907/U$1 ( \25637 , \25635 , \25636 );
nand \g444502/U$1 ( \25638 , \25628 , \25631 , \25634 , \25637 );
and \g446127/U$2 ( \25639 , RIfcb3a20_7066, \8373 );
and \g446127/U$3 ( \25640 , RIe1eeb38_4093, \8335 );
and \g449041/U$2 ( \25641 , RIfc97550_6744, \8531 );
and \g449041/U$3 ( \25642 , \8488 , RIfca2ef0_6876);
and \g449041/U$4 ( \25643 , RIfcbdea8_7183, \8383 );
nor \g449041/U$1 ( \25644 , \25641 , \25642 , \25643 );
and \g452388/U$2 ( \25645 , \8356 , RIe1f3e30_4152);
and \g452388/U$3 ( \25646 , RIfc904d0_6664, \8359 );
nor \g452388/U$1 ( \25647 , \25645 , \25646 );
and \g454306/U$2 ( \25648 , \8313 , RIfcd20b0_7412);
and \g454306/U$3 ( \25649 , RIfc90200_6662, \8323 );
nor \g454306/U$1 ( \25650 , \25648 , \25649 );
not \g450055/U$3 ( \25651 , \25650 );
not \g450055/U$4 ( \25652 , \8376 );
and \g450055/U$2 ( \25653 , \25651 , \25652 );
and \g450055/U$5 ( \25654 , \8351 , RIfca2d88_6875);
nor \g450055/U$1 ( \25655 , \25653 , \25654 );
and \g452386/U$2 ( \25656 , \8378 , RIe1f6158_4177);
and \g452386/U$3 ( \25657 , RIfc90098_6661, \8417 );
nor \g452386/U$1 ( \25658 , \25656 , \25657 );
nand \g447746/U$1 ( \25659 , \25644 , \25647 , \25655 , \25658 );
nor \g446127/U$1 ( \25660 , \25639 , \25640 , \25659 );
and \g452383/U$2 ( \25661 , \8340 , RIfc59048_6035);
and \g452383/U$3 ( \25662 , RIe1fabe0_4230, \8404 );
nor \g452383/U$1 ( \25663 , \25661 , \25662 );
and \g452384/U$2 ( \25664 , \8319 , RIfc90638_6665);
and \g452384/U$3 ( \25665 , RIfc907a0_6666, \8326 );
nor \g452384/U$1 ( \25666 , \25664 , \25665 );
and \g445239/U$2 ( \25667 , \25660 , \25663 , \25666 );
nor \g445239/U$1 ( \25668 , \25667 , \8621 );
and \g446128/U$2 ( \25669 , RIe18d518_2985, \8417 );
and \g446128/U$3 ( \25670 , RIe1f16d0_4124, \8356 );
and \g449044/U$2 ( \25671 , RIe1af550_3372, \8319 );
and \g449044/U$3 ( \25672 , \8326 , RIe1bc6d8_3521);
and \g449044/U$4 ( \25673 , RIe1ff7d0_4284, \8488 );
nor \g449044/U$1 ( \25674 , \25671 , \25672 , \25673 );
and \g452395/U$2 ( \25675 , \8335 , RIe171b88_2671);
and \g452395/U$3 ( \25676 , RIe1d5bd8_3809, \8340 );
nor \g452395/U$1 ( \25677 , \25675 , \25676 );
and \g452394/U$2 ( \25678 , \8404 , RIe1a1018_3209);
and \g452394/U$3 ( \25679 , RIe1a9718_3305, \8351 );
nor \g452394/U$1 ( \25680 , \25678 , \25679 );
and \g454834/U$2 ( \25681 , \8313 , RIe1a3d18_3241);
and \g454834/U$3 ( \25682 , RIe1a6a18_3273, \8323 );
nor \g454834/U$1 ( \25683 , \25681 , \25682 );
not \g450058/U$3 ( \25684 , \25683 );
not \g450058/U$4 ( \25685 , \8328 );
and \g450058/U$2 ( \25686 , \25684 , \25685 );
and \g450058/U$5 ( \25687 , \8359 , RIe205770_4352);
nor \g450058/U$1 ( \25688 , \25686 , \25687 );
nand \g447747/U$1 ( \25689 , \25674 , \25677 , \25680 , \25688 );
nor \g446128/U$1 ( \25690 , \25669 , \25670 , \25689 );
and \g452392/U$2 ( \25691 , \8378 , RIe21bf70_4608);
and \g452392/U$3 ( \25692 , RIe1f8b88_4207, \8523 );
nor \g452392/U$1 ( \25693 , \25691 , \25692 );
and \g452391/U$2 ( \25694 , \8414 , RIe227370_4736);
and \g452391/U$3 ( \25695 , RIe179a18_2761, \8409 );
nor \g452391/U$1 ( \25696 , \25694 , \25695 );
and \g445241/U$2 ( \25697 , \25690 , \25693 , \25696 );
nor \g445241/U$1 ( \25698 , \25697 , \8651 );
or \g444292/U$1 ( \25699 , \25577 , \25638 , \25668 , \25698 );
and \g446123/U$2 ( \25700 , RIe192f18_3049, \8414 );
and \g446123/U$3 ( \25701 , RIf144b18_5241, \8417 );
and \g449037/U$2 ( \25702 , RIfc8f3f0_6652, \8373 );
and \g449037/U$3 ( \25703 , \8383 , RIe19b618_3145);
and \g449037/U$4 ( \25704 , RIe187b18_2921, \8488 );
nor \g449037/U$1 ( \25705 , \25702 , \25703 , \25704 );
and \g452372/U$2 ( \25706 , \8335 , RIe17c718_2793);
and \g452372/U$3 ( \25707 , RIfcb3cf0_7068, \8340 );
nor \g452372/U$1 ( \25708 , \25706 , \25707 );
and \g452371/U$2 ( \25709 , \8404 , RIe198918_3113);
and \g452371/U$3 ( \25710 , RIe19e318_3177, \8351 );
nor \g452371/U$1 ( \25711 , \25709 , \25710 );
and \g454821/U$2 ( \25712 , \8313 , RIe17f418_2825);
and \g454821/U$3 ( \25713 , RIe182118_2857, \8323 );
nor \g454821/U$1 ( \25714 , \25712 , \25713 );
not \g454820/U$1 ( \25715 , \25714 );
and \g450050/U$2 ( \25716 , \25715 , \8316 );
and \g450050/U$3 ( \25717 , RIe18a818_2953, \8359 );
nor \g450050/U$1 ( \25718 , \25716 , \25717 );
nand \g448195/U$1 ( \25719 , \25705 , \25708 , \25711 , \25718 );
nor \g446123/U$1 ( \25720 , \25700 , \25701 , \25719 );
and \g452367/U$2 ( \25721 , \8378 , RIe190218_3017);
and \g452367/U$3 ( \25722 , RIf143d08_5231, \8531 );
nor \g452367/U$1 ( \25723 , \25721 , \25722 );
and \g452368/U$2 ( \25724 , \8356 , RIe184e18_2889);
and \g452368/U$3 ( \25725 , RIe195c18_3081, \8409 );
nor \g452368/U$1 ( \25726 , \25724 , \25725 );
and \g445236/U$2 ( \25727 , \25720 , \25723 , \25726 );
nor \g445236/U$1 ( \25728 , \25727 , \8589 );
and \g446124/U$2 ( \25729 , RIfc57e00_6022, \8417 );
and \g446124/U$3 ( \25730 , RIe1742e8_2699, \8356 );
and \g449040/U$2 ( \25731 , RIfc7c9d0_6440, \8373 );
and \g449040/U$3 ( \25732 , \8330 , RIf141170_5200);
and \g449040/U$4 ( \25733 , RIfce0048_7571, \8488 );
nor \g449040/U$1 ( \25734 , \25731 , \25732 , \25733 );
and \g452380/U$2 ( \25735 , \8335 , RIfc583a0_6026);
and \g452380/U$3 ( \25736 , RIfc7c700_6438, \8340 );
nor \g452380/U$1 ( \25737 , \25735 , \25736 );
and \g452379/U$2 ( \25738 , \8404 , RIfea0098_8165);
and \g452379/U$3 ( \25739 , RIfc448a0_5802, \8351 );
nor \g452379/U$1 ( \25740 , \25738 , \25739 );
and \g454829/U$2 ( \25741 , \8313 , RIfce9828_7679);
and \g454829/U$3 ( \25742 , RIfc8f990_6656, \8323 );
nor \g454829/U$1 ( \25743 , \25741 , \25742 );
not \g454828/U$1 ( \25744 , \25743 );
and \g450054/U$2 ( \25745 , \25744 , \8316 );
and \g450054/U$3 ( \25746 , RIfc8f6c0_6654, \8359 );
nor \g450054/U$1 ( \25747 , \25745 , \25746 );
nand \g448196/U$1 ( \25748 , \25734 , \25737 , \25740 , \25747 );
nor \g446124/U$1 ( \25749 , \25729 , \25730 , \25748 );
and \g452378/U$2 ( \25750 , \8378 , RIee3d900_5159);
and \g452378/U$3 ( \25751 , RIfca27e8_6871, \8531 );
nor \g452378/U$1 ( \25752 , \25750 , \25751 );
and \g452377/U$2 ( \25753 , \8414 , RIfcd6e08_7467);
and \g452377/U$3 ( \25754 , RIf13f550_5180, \8407 );
nor \g452377/U$1 ( \25755 , \25753 , \25754 );
and \g445237/U$2 ( \25756 , \25749 , \25752 , \25755 );
nor \g445237/U$1 ( \25757 , \25756 , \8558 );
or \g444234/U$1 ( \25758 , \25699 , \25728 , \25757 );
_DC \g4770/U$1 ( \25759 , \25758 , \8654 );
and \g452904/U$2 ( \25760 , \16364 , RIdf31f60_1945);
and \g452904/U$3 ( \25761 , RIfc8ece8_6647, \16371 );
nor \g452904/U$1 ( \25762 , \25760 , \25761 );
and \g446236/U$2 ( \25763 , RIee2ff08_5004, \16427 );
and \g446236/U$3 ( \25764 , RIee2dd48_4980, \16368 );
and \g449183/U$2 ( \25765 , RIe13f9f8_2101, \16485 );
and \g449183/U$3 ( \25766 , \16356 , RIe141d20_2126);
and \g449183/U$4 ( \25767 , RIdf34120_1969, \16398 );
nor \g449183/U$1 ( \25768 , \25765 , \25766 , \25767 );
and \g455050/U$2 ( \25769 , \16317 , RIfc45278_5809);
and \g455050/U$3 ( \25770 , RIfc8ee50_6648, \16325 );
nor \g455050/U$1 ( \25771 , \25769 , \25770 );
not \g450200/U$3 ( \25772 , \25771 );
not \g450200/U$4 ( \25773 , \16311 );
and \g450200/U$2 ( \25774 , \25772 , \25773 );
and \g450200/U$5 ( \25775 , \16341 , RIdf36718_1996);
nor \g450200/U$1 ( \25776 , \25774 , \25775 );
and \g452907/U$2 ( \25777 , \16377 , RIfca2248_6867);
and \g452907/U$3 ( \25778 , RIfc98360_6754, \16313 );
nor \g452907/U$1 ( \25779 , \25777 , \25778 );
and \g452909/U$2 ( \25780 , \16334 , RIdf3b470_2051);
and \g452909/U$3 ( \25781 , RIdf3d900_2077, \16380 );
nor \g452909/U$1 ( \25782 , \25780 , \25781 );
nand \g447391/U$1 ( \25783 , \25768 , \25776 , \25779 , \25782 );
nor \g446236/U$1 ( \25784 , \25763 , \25764 , \25783 );
and \g452905/U$2 ( \25785 , \16361 , RIfe9f6c0_8158);
and \g452905/U$3 ( \25786 , RIfcd6ca0_7466, \16448 );
nor \g452905/U$1 ( \25787 , \25785 , \25786 );
nand \g445638/U$1 ( \25788 , \25762 , \25784 , \25787 );
and \g444789/U$2 ( \25789 , \25788 , \16394 );
and \g449181/U$2 ( \25790 , RIe14cfb8_2253, \16398 );
and \g449181/U$3 ( \25791 , \16341 , RIfcbd368_7175);
and \g449181/U$4 ( \25792 , RIe15ddb8_2445, \16344 );
nor \g449181/U$1 ( \25793 , \25790 , \25791 , \25792 );
and \g455129/U$2 ( \25794 , \16317 , RIe1529b8_2317);
and \g455129/U$3 ( \25795 , RIfe9f828_8159, \16325 );
nor \g455129/U$1 ( \25796 , \25794 , \25795 );
not \g450197/U$3 ( \25797 , \25796 );
not \g450197/U$4 ( \25798 , \16351 );
and \g450197/U$2 ( \25799 , \25797 , \25798 );
and \g450197/U$5 ( \25800 , \16354 , RIfc8ea18_6645);
nor \g450197/U$1 ( \25801 , \25799 , \25800 );
and \g452900/U$2 ( \25802 , \16361 , RIe1475b8_2189);
and \g452900/U$3 ( \25803 , RIe14a2b8_2221, \16364 );
nor \g452900/U$1 ( \25804 , \25802 , \25803 );
and \g452898/U$2 ( \25805 , \16368 , RIe14fcb8_2285);
and \g452898/U$3 ( \25806 , RIfe9f990_8160, \16371 );
nor \g452898/U$1 ( \25807 , \25805 , \25806 );
nand \g447814/U$1 ( \25808 , \25793 , \25801 , \25804 , \25807 );
and \g444789/U$3 ( \25809 , \16390 , \25808 );
nor \g444789/U$1 ( \25810 , \25789 , \25809 );
and \g447006/U$2 ( \25811 , \18020 , RIe1637b8_2509);
and \g447006/U$3 ( \25812 , RIe1664b8_2541, \18022 );
nor \g447006/U$1 ( \25813 , \25811 , \25812 );
and \g447007/U$2 ( \25814 , \18025 , RIe160ab8_2477);
and \g447007/U$3 ( \25815 , RIee37f00_5095, \18027 );
nor \g447007/U$1 ( \25816 , \25814 , \25815 );
and \g447008/U$2 ( \25817 , \18030 , RIe1556b8_2349);
and \g447008/U$3 ( \25818 , RIe1583b8_2381, \18032 );
nor \g447008/U$1 ( \25819 , \25817 , \25818 );
nand \g444516/U$1 ( \25820 , \25810 , \25813 , \25816 , \25819 );
and \g452887/U$2 ( \25821 , \16364 , RIe16a298_2585);
and \g452887/U$3 ( \25822 , RIfcd96d0_7496, \16371 );
nor \g452887/U$1 ( \25823 , \25821 , \25822 );
and \g446231/U$2 ( \25824 , RIfc8e040_6638, \16427 );
and \g446231/U$3 ( \25825 , RIfca1e10_6864, \16368 );
and \g449178/U$2 ( \25826 , RIfc8ded8_6637, \16321 );
and \g449178/U$3 ( \25827 , \16328 , RIfcd6868_7463);
and \g449178/U$4 ( \25828 , RIe16c5c0_2610, \16337 );
nor \g449178/U$1 ( \25829 , \25826 , \25827 , \25828 );
and \g455083/U$2 ( \25830 , \16317 , RIde8f300_288);
and \g455083/U$3 ( \25831 , RIde92e10_306, \16325 );
nor \g455083/U$1 ( \25832 , \25830 , \25831 );
not \g450196/U$3 ( \25833 , \25832 );
not \g450196/U$4 ( \25834 , \16330 );
and \g450196/U$2 ( \25835 , \25833 , \25834 );
and \g450196/U$5 ( \25836 , \16341 , RIfcbd200_7174);
nor \g450196/U$1 ( \25837 , \25835 , \25836 );
and \g452891/U$2 ( \25838 , \16377 , RIfc56618_6005);
and \g452891/U$3 ( \25839 , RIfc7dd80_6454, \16313 );
nor \g452891/U$1 ( \25840 , \25838 , \25839 );
and \g452892/U$2 ( \25841 , \16334 , RIde86fc0_248);
and \g452892/U$3 ( \25842 , RIde8b160_268, \16380 );
nor \g452892/U$1 ( \25843 , \25841 , \25842 );
nand \g447390/U$1 ( \25844 , \25829 , \25837 , \25840 , \25843 );
nor \g446231/U$1 ( \25845 , \25824 , \25825 , \25844 );
and \g452888/U$2 ( \25846 , \16361 , RIe168ab0_2568);
and \g452888/U$3 ( \25847 , RIde82ad8_227, \16448 );
nor \g452888/U$1 ( \25848 , \25846 , \25847 );
nand \g445636/U$1 ( \25849 , \25823 , \25845 , \25848 );
and \g444711/U$2 ( \25850 , \25849 , \17998 );
and \g449175/U$2 ( \25851 , RIdec37b8_688, \16321 );
and \g449175/U$3 ( \25852 , \16326 , RIdec64b8_720);
and \g449175/U$4 ( \25853 , RIdeacb80_432, \16398 );
nor \g449175/U$1 ( \25854 , \25851 , \25852 , \25853 );
and \g455072/U$2 ( \25855 , \16317 , RIdebddb8_624);
and \g455072/U$3 ( \25856 , RIfc56348_6003, \16325 );
nor \g455072/U$1 ( \25857 , \25855 , \25856 );
not \g450192/U$3 ( \25858 , \25857 );
not \g450192/U$4 ( \25859 , \16330 );
and \g450192/U$2 ( \25860 , \25858 , \25859 );
and \g450192/U$5 ( \25861 , \16339 , RIfc8dc08_6635);
nor \g450192/U$1 ( \25862 , \25860 , \25861 );
and \g452884/U$2 ( \25863 , \16377 , RIdec0ab8_656);
and \g452884/U$3 ( \25864 , RIfc8daa0_6634, \16313 );
nor \g452884/U$1 ( \25865 , \25863 , \25864 );
and \g452886/U$2 ( \25866 , \16334 , RIdeb83b8_560);
and \g452886/U$3 ( \25867 , RIdebb0b8_592, \16380 );
nor \g452886/U$1 ( \25868 , \25866 , \25867 );
nand \g447389/U$1 ( \25869 , \25854 , \25862 , \25865 , \25868 );
and \g444711/U$3 ( \25870 , \17938 , \25869 );
nor \g444711/U$1 ( \25871 , \25850 , \25870 );
and \g447001/U$2 ( \25872 , \18457 , RIdeb29b8_496);
and \g447001/U$3 ( \25873 , RIfc98798_6757, \18459 );
nor \g447001/U$1 ( \25874 , \25872 , \25873 );
and \g447000/U$2 ( \25875 , \18462 , RIdeafcb8_464);
and \g447000/U$3 ( \25876 , RIfcbd098_7173, \18464 );
nor \g447000/U$1 ( \25877 , \25875 , \25876 );
and \g447002/U$2 ( \25878 , \18467 , RIde9f980_368);
and \g447002/U$3 ( \25879 , RIdea6280_400, \18469 );
nor \g447002/U$1 ( \25880 , \25878 , \25879 );
nand \g444515/U$1 ( \25881 , \25871 , \25874 , \25877 , \25880 );
and \g446227/U$2 ( \25882 , RIfc44e40_5806, \16321 );
and \g446227/U$3 ( \25883 , RIfc57860_6018, \16313 );
and \g449171/U$2 ( \25884 , RIee22678_4850, \16427 );
and \g449171/U$3 ( \25885 , \16448 , RIfcbd4d0_7176);
and \g449171/U$4 ( \25886 , RIdee3900_1053, \16485 );
nor \g449171/U$1 ( \25887 , \25884 , \25885 , \25886 );
and \g455180/U$2 ( \25888 , \16317 , RIded80c8_922);
and \g455180/U$3 ( \25889 , RIfe9fc60_8162, \16325 );
nor \g455180/U$1 ( \25890 , \25888 , \25889 );
not \g455179/U$1 ( \25891 , \25890 );
and \g450186/U$2 ( \25892 , \25891 , \16336 );
and \g450186/U$3 ( \25893 , RIfe9faf8_8161, \16356 );
nor \g450186/U$1 ( \25894 , \25892 , \25893 );
and \g452867/U$2 ( \25895 , \16361 , RIded3be0_873);
and \g452867/U$3 ( \25896 , RIfe9fdc8_8163, \16364 );
nor \g452867/U$1 ( \25897 , \25895 , \25896 );
and \g452864/U$2 ( \25898 , \16368 , RIee21598_4838);
and \g452864/U$3 ( \25899 , RIfc98090_6752, \16371 );
nor \g452864/U$1 ( \25900 , \25898 , \25899 );
nand \g448092/U$1 ( \25901 , \25887 , \25894 , \25897 , \25900 );
nor \g446227/U$1 ( \25902 , \25882 , \25883 , \25901 );
and \g452862/U$2 ( \25903 , \16377 , RIfca23b0_6868);
and \g452862/U$3 ( \25904 , RIdee1740_1029, \16380 );
nor \g452862/U$1 ( \25905 , \25903 , \25904 );
and \g452860/U$2 ( \25906 , \16334 , RIdedf6e8_1006);
and \g452860/U$3 ( \25907 , RIfc8efb8_6649, \16328 );
nor \g452860/U$1 ( \25908 , \25906 , \25907 );
and \g445310/U$2 ( \25909 , \25902 , \25905 , \25908 );
nor \g445310/U$1 ( \25910 , \25909 , \16909 );
and \g446228/U$2 ( \25911 , RIfc8e748_6643, \16427 );
and \g446228/U$3 ( \25912 , RIfcc2c00_7238, \16368 );
and \g449173/U$2 ( \25913 , RIfc45db8_5817, \16319 );
and \g449173/U$3 ( \25914 , \16328 , RIfcb4560_7074);
and \g449173/U$4 ( \25915 , RIdf20788_1746, \16337 );
nor \g449173/U$1 ( \25916 , \25913 , \25914 , \25915 );
and \g455065/U$2 ( \25917 , \16317 , RIdf28ff0_1843);
and \g455065/U$3 ( \25918 , RIdf2aee0_1865, \16325 );
nor \g455065/U$1 ( \25919 , \25917 , \25918 );
not \g450188/U$3 ( \25920 , \25919 );
not \g450188/U$4 ( \25921 , \16330 );
and \g450188/U$2 ( \25922 , \25920 , \25921 );
and \g450188/U$5 ( \25923 , \16341 , RIdf21e08_1762);
nor \g450188/U$1 ( \25924 , \25922 , \25923 );
and \g452874/U$2 ( \25925 , \16377 , RIfc7d678_6449);
and \g452874/U$3 ( \25926 , RIfc8e1a8_6639, \16313 );
nor \g452874/U$1 ( \25927 , \25925 , \25926 );
and \g452876/U$2 ( \25928 , \16334 , RIdf25378_1800);
and \g452876/U$3 ( \25929 , RIdf26e30_1819, \16380 );
nor \g452876/U$1 ( \25930 , \25928 , \25929 );
nand \g447388/U$1 ( \25931 , \25916 , \25924 , \25927 , \25930 );
nor \g446228/U$1 ( \25932 , \25911 , \25912 , \25931 );
and \g452870/U$2 ( \25933 , \16361 , RIdf1a248_1674);
and \g452870/U$3 ( \25934 , RIfcb43f8_7073, \16432 );
nor \g452870/U$1 ( \25935 , \25933 , \25934 );
and \g452869/U$2 ( \25936 , \16364 , RIdf1b760_1689);
and \g452869/U$3 ( \25937 , RIdf23488_1778, \16371 );
nor \g452869/U$1 ( \25938 , \25936 , \25937 );
and \g445312/U$2 ( \25939 , \25932 , \25935 , \25938 );
nor \g445312/U$1 ( \25940 , \25939 , \16480 );
or \g444332/U$1 ( \25941 , \25820 , \25881 , \25910 , \25940 );
and \g446221/U$2 ( \25942 , RIdf15388_1618, \16321 );
and \g446221/U$3 ( \25943 , RIdf12688_1586, \16313 );
and \g449167/U$2 ( \25944 , RIdefbe88_1330, \16427 );
and \g449167/U$3 ( \25945 , \16448 , RIdefeb88_1362);
and \g449167/U$4 ( \25946 , RIdf09f88_1490, \16485 );
nor \g449167/U$1 ( \25947 , \25944 , \25945 , \25946 );
and \g455231/U$2 ( \25948 , \16317 , RIdef0a88_1202);
and \g455231/U$3 ( \25949 , RIdef3788_1234, \16325 );
nor \g455231/U$1 ( \25950 , \25948 , \25949 );
not \g455230/U$1 ( \25951 , \25950 );
and \g450182/U$2 ( \25952 , \25951 , \16336 );
and \g450182/U$3 ( \25953 , RIdf0cc88_1522, \16356 );
nor \g450182/U$1 ( \25954 , \25952 , \25953 );
and \g452843/U$2 ( \25955 , \16361 , RIdeeb088_1138);
and \g452843/U$3 ( \25956 , RIdeedd88_1170, \16364 );
nor \g452843/U$1 ( \25957 , \25955 , \25956 );
and \g452842/U$2 ( \25958 , \16368 , RIdef6488_1266);
and \g452842/U$3 ( \25959 , RIdef9188_1298, \16371 );
nor \g452842/U$1 ( \25960 , \25958 , \25959 );
nand \g448091/U$1 ( \25961 , \25947 , \25954 , \25957 , \25960 );
nor \g446221/U$1 ( \25962 , \25942 , \25943 , \25961 );
and \g452841/U$2 ( \25963 , \16377 , RIdf0f988_1554);
and \g452841/U$3 ( \25964 , RIdf07288_1458, \16380 );
nor \g452841/U$1 ( \25965 , \25963 , \25964 );
and \g452840/U$2 ( \25966 , \16334 , RIdf04588_1426);
and \g452840/U$3 ( \25967 , RIdf18088_1650, \16328 );
nor \g452840/U$1 ( \25968 , \25966 , \25967 );
and \g445305/U$2 ( \25969 , \25962 , \25965 , \25968 );
nor \g445305/U$1 ( \25970 , \25969 , \16555 );
and \g446224/U$2 ( \25971 , RIdf392b0_2027, \16427 );
and \g446224/U$3 ( \25972 , RIdf1e190_1719, \16368 );
and \g449169/U$2 ( \25973 , RIde99080_336, \16344 );
and \g449169/U$3 ( \25974 , \16356 , RIdeb56b8_528);
and \g449169/U$4 ( \25975 , RIdee8388_1106, \16398 );
nor \g449169/U$1 ( \25976 , \25973 , \25974 , \25975 );
and \g455051/U$2 ( \25977 , \16317 , RIdecebb8_816);
and \g455051/U$3 ( \25978 , RIded18b8_848, \16325 );
nor \g455051/U$1 ( \25979 , \25977 , \25978 );
not \g450184/U$3 ( \25980 , \25979 );
not \g450184/U$4 ( \25981 , \16311 );
and \g450184/U$2 ( \25982 , \25980 , \25981 );
and \g450184/U$5 ( \25983 , \16341 , RIdf01888_1394);
nor \g450184/U$1 ( \25984 , \25982 , \25983 );
and \g452854/U$2 ( \25985 , \16377 , RIdec91b8_752);
and \g452854/U$3 ( \25986 , RIdecbeb8_784, \16313 );
nor \g452854/U$1 ( \25987 , \25985 , \25986 );
and \g452855/U$2 ( \25988 , \16334 , RIe15b0b8_2413);
and \g452855/U$3 ( \25989 , RIe16f2c0_2642, \16380 );
nor \g452855/U$1 ( \25990 , \25988 , \25989 );
nand \g447386/U$1 ( \25991 , \25976 , \25984 , \25987 , \25990 );
nor \g446224/U$1 ( \25992 , \25971 , \25972 , \25991 );
and \g452852/U$2 ( \25993 , \16361 , RIde7efc8_209);
and \g452852/U$3 ( \25994 , RIe1448b8_2157, \16448 );
nor \g452852/U$1 ( \25995 , \25993 , \25994 );
and \g452850/U$2 ( \25996 , \16364 , RIdedd0f0_979);
and \g452850/U$3 ( \25997 , RIdf2d910_1895, \16371 );
nor \g452850/U$1 ( \25998 , \25996 , \25997 );
and \g445308/U$2 ( \25999 , \25992 , \25995 , \25998 );
nor \g445308/U$1 ( \26000 , \25999 , \16586 );
or \g444227/U$1 ( \26001 , \25941 , \25970 , \26000 );
_DC \g47f5/U$1 ( \26002 , \26001 , \16652 );
and \g449212/U$2 ( \26003 , RIfc47000_5830, \8531 );
and \g449212/U$3 ( \26004 , \8488 , RIe213ca8_4515);
and \g449212/U$4 ( \26005 , RIe224aa8_4707, \8330 );
nor \g449212/U$1 ( \26006 , \26003 , \26004 , \26005 );
and \g453006/U$2 ( \26007 , \8335 , RIe2088a8_4387);
and \g453006/U$3 ( \26008 , RIfcbc990_7168, \8340 );
nor \g453006/U$1 ( \26009 , \26007 , \26008 );
and \g455158/U$2 ( \26010 , \8313 , RIe20b5a8_4419);
and \g455158/U$3 ( \26011 , RIe20e2a8_4451, \8323 );
nor \g455158/U$1 ( \26012 , \26010 , \26011 );
not \g455157/U$1 ( \26013 , \26012 );
and \g450228/U$2 ( \26014 , \26013 , \8316 );
and \g450228/U$3 ( \26015 , RIfe9f288_8155, \8351 );
nor \g450228/U$1 ( \26016 , \26014 , \26015 );
and \g453005/U$2 ( \26017 , \8356 , RIe210fa8_4483);
and \g453005/U$3 ( \26018 , RIfcbc828_7167, \8359 );
nor \g453005/U$1 ( \26019 , \26017 , \26018 );
nand \g448211/U$1 ( \26020 , \26006 , \26009 , \26016 , \26019 );
and \g444792/U$2 ( \26021 , \26020 , \8369 );
and \g446258/U$2 ( \26022 , RIe1fd340_4258, \8531 );
and \g446258/U$3 ( \26023 , RIfc7ea28_6463, \8319 );
and \g449213/U$2 ( \26024 , RIe2032e0_4326, \8373 );
and \g449213/U$3 ( \26025 , \8383 , RIfcd6598_7461);
and \g449213/U$4 ( \26026 , RIfcb4dd0_7080, \8488 );
nor \g449213/U$1 ( \26027 , \26024 , \26025 , \26026 );
and \g454295/U$2 ( \26028 , \8313 , RIfce0318_7573);
and \g454295/U$3 ( \26029 , RIfc7eb90_6464, \8323 );
nor \g454295/U$1 ( \26030 , \26028 , \26029 );
not \g450230/U$3 ( \26031 , \26030 );
not \g450230/U$4 ( \26032 , \8376 );
and \g450230/U$2 ( \26033 , \26031 , \26032 );
and \g450230/U$5 ( \26034 , \8359 , RIfc8cf60_6626);
nor \g450230/U$1 ( \26035 , \26033 , \26034 );
and \g453011/U$2 ( \26036 , \8404 , RIe2016c0_4306);
and \g453011/U$3 ( \26037 , RIfc46bc8_5827, \8351 );
nor \g453011/U$1 ( \26038 , \26036 , \26037 );
and \g453013/U$2 ( \26039 , \8378 , RIfcbcaf8_7169);
and \g453013/U$3 ( \26040 , RIfc98ea0_6762, \8417 );
nor \g453013/U$1 ( \26041 , \26039 , \26040 );
nand \g447836/U$1 ( \26042 , \26027 , \26035 , \26038 , \26041 );
nor \g446258/U$1 ( \26043 , \26022 , \26023 , \26042 );
and \g453009/U$2 ( \26044 , \8335 , RIfc8d0c8_6627);
and \g453009/U$3 ( \26045 , RIf15cf38_5517, \8340 );
nor \g453009/U$1 ( \26046 , \26044 , \26045 );
and \g453008/U$2 ( \26047 , \8324 , RIfe9f120_8154);
and \g453008/U$3 ( \26048 , RIe1fc260_4246, \8356 );
nor \g453008/U$1 ( \26049 , \26047 , \26048 );
and \g445334/U$2 ( \26050 , \26043 , \26046 , \26049 );
nor \g445334/U$1 ( \26051 , \26050 , \8422 );
nor \g444792/U$1 ( \26052 , \26021 , \26051 );
and \g447027/U$2 ( \26053 , \8426 , RIe221da8_4675);
and \g447027/U$3 ( \26054 , RIfc55808_5995, \8428 );
nor \g447027/U$1 ( \26055 , \26053 , \26054 );
and \g447026/U$2 ( \26056 , \8431 , RIe21f0a8_4643);
and \g447026/U$3 ( \26057 , RIfcb50a0_7082, \8434 );
nor \g447026/U$1 ( \26058 , \26056 , \26057 );
and \g447028/U$2 ( \26059 , \8438 , RIe2169a8_4547);
and \g447028/U$3 ( \26060 , RIe2196a8_4579, \8440 );
nor \g447028/U$1 ( \26061 , \26059 , \26060 );
nand \g444520/U$1 ( \26062 , \26052 , \26055 , \26058 , \26061 );
and \g453026/U$2 ( \26063 , \8404 , RIe1e4110_3972);
and \g453026/U$3 ( \26064 , RIe1de710_3908, \8409 );
nor \g453026/U$1 ( \26065 , \26063 , \26064 );
and \g446260/U$2 ( \26066 , RIe1e6e10_4004, \8373 );
and \g446260/U$3 ( \26067 , RIe1d8d10_3844, \8378 );
and \g449219/U$2 ( \26068 , RIe1c2510_3588, \8319 );
and \g449219/U$3 ( \26069 , \8326 , RIe1c5210_3620);
and \g449219/U$4 ( \26070 , RIe1e9b10_4036, \8383 );
nor \g449219/U$1 ( \26071 , \26068 , \26069 , \26070 );
and \g453032/U$2 ( \26072 , \8335 , RIe1bf810_3556);
and \g453032/U$3 ( \26073 , RIe1c7f10_3652, \8340 );
nor \g453032/U$1 ( \26074 , \26072 , \26073 );
and \g455178/U$2 ( \26075 , \8313 , RIe1cd910_3716);
and \g455178/U$3 ( \26076 , RIe1d0610_3748, \8323 );
nor \g455178/U$1 ( \26077 , \26075 , \26076 );
not \g450235/U$3 ( \26078 , \26077 );
not \g450235/U$4 ( \26079 , \8347 );
and \g450235/U$2 ( \26080 , \26078 , \26079 );
and \g450235/U$5 ( \26081 , \8351 , RIe1ec810_4068);
nor \g450235/U$1 ( \26082 , \26080 , \26081 );
and \g453030/U$2 ( \26083 , \8356 , RIe1cac10_3684);
and \g453030/U$3 ( \26084 , RIe1d3310_3780, \8359 );
nor \g453030/U$1 ( \26085 , \26083 , \26084 );
nand \g447838/U$1 ( \26086 , \26071 , \26074 , \26082 , \26085 );
nor \g446260/U$1 ( \26087 , \26066 , \26067 , \26086 );
and \g453025/U$2 ( \26088 , \8414 , RIe1dba10_3876);
and \g453025/U$3 ( \26089 , RIe1e1410_3940, \8417 );
nor \g453025/U$1 ( \26090 , \26088 , \26089 );
nand \g445641/U$1 ( \26091 , \26065 , \26087 , \26090 );
and \g444793/U$2 ( \26092 , \26091 , \8478 );
and \g449217/U$2 ( \26093 , RIfc8d500_6630, \8319 );
and \g449217/U$3 ( \26094 , \8326 , RIfc8d398_6629);
and \g449217/U$4 ( \26095 , RIfc98bd0_6760, \8383 );
nor \g449217/U$1 ( \26096 , \26093 , \26094 , \26095 );
and \g453021/U$2 ( \26097 , \8335 , RIe1eef70_4096);
and \g453021/U$3 ( \26098 , RIfceedf0_7740, \8340 );
nor \g453021/U$1 ( \26099 , \26097 , \26098 );
and \g454315/U$2 ( \26100 , \8313 , RIfcc2ed0_7240);
and \g454315/U$3 ( \26101 , RIfc468f8_5825, \8323 );
nor \g454315/U$1 ( \26102 , \26100 , \26101 );
not \g450232/U$3 ( \26103 , \26102 );
not \g450232/U$4 ( \26104 , \8347 );
and \g450232/U$2 ( \26105 , \26103 , \26104 );
and \g450232/U$5 ( \26106 , \8351 , RIfcbcc60_7170);
nor \g450232/U$1 ( \26107 , \26105 , \26106 );
and \g453020/U$2 ( \26108 , \8356 , RIe1f4100_4154);
and \g453020/U$3 ( \26109 , RIfce58e0_7634, \8359 );
nor \g453020/U$1 ( \26110 , \26108 , \26109 );
nand \g447837/U$1 ( \26111 , \26096 , \26099 , \26107 , \26110 );
and \g444793/U$3 ( \26112 , \8752 , \26111 );
nor \g444793/U$1 ( \26113 , \26092 , \26112 );
and \g447036/U$2 ( \26114 , \11511 , RIe1fb018_4233);
and \g447036/U$3 ( \26115 , RIfce2d48_7603, \11513 );
nor \g447036/U$1 ( \26116 , \26114 , \26115 );
and \g447035/U$2 ( \26117 , \11516 , RIfc7e8c0_6462);
and \g447035/U$3 ( \26118 , RIfc55f10_6000, \11518 );
nor \g447035/U$1 ( \26119 , \26117 , \26118 );
and \g447037/U$2 ( \26120 , \11521 , RIe1f6590_4180);
and \g447037/U$3 ( \26121 , RIfc8d230_6628, \11523 );
nor \g447037/U$1 ( \26122 , \26120 , \26121 );
nand \g444521/U$1 ( \26123 , \26113 , \26116 , \26119 , \26122 );
and \g446254/U$2 ( \26124 , RIfec4dd0_8360, \8417 );
and \g446254/U$3 ( \26125 , RIe1b8088_3471, \8404 );
and \g449207/U$2 ( \26126 , RIfec5370_8364, \8531 );
and \g449207/U$3 ( \26127 , \8486 , RIfcb4c68_7079);
and \g449207/U$4 ( \26128 , RIfe9efb8_8153, \8383 );
nor \g449207/U$1 ( \26129 , \26126 , \26127 , \26128 );
and \g452992/U$2 ( \26130 , \8335 , RIfec4f38_8361);
and \g452992/U$3 ( \26131 , RIfcbcdc8_7171, \8340 );
nor \g452992/U$1 ( \26132 , \26130 , \26131 );
and \g454887/U$2 ( \26133 , \8313 , RIfec5208_8363);
and \g454887/U$3 ( \26134 , RIfc46358_5821, \8323 );
nor \g454887/U$1 ( \26135 , \26133 , \26134 );
not \g454886/U$1 ( \26136 , \26135 );
and \g450222/U$2 ( \26137 , \26136 , \8316 );
and \g450222/U$3 ( \26138 , RIf14d0b0_5336, \8351 );
nor \g450222/U$1 ( \26139 , \26137 , \26138 );
and \g452990/U$2 ( \26140 , \8356 , RIfe9ee50_8152);
and \g452990/U$3 ( \26141 , RIfcb4998_7077, \8359 );
nor \g452990/U$1 ( \26142 , \26140 , \26141 );
nand \g448209/U$1 ( \26143 , \26129 , \26132 , \26139 , \26142 );
nor \g446254/U$1 ( \26144 , \26124 , \26125 , \26143 );
and \g452987/U$2 ( \26145 , \8378 , RIe1b46e0_3430);
and \g452987/U$3 ( \26146 , RIe1ba248_3495, \8373 );
nor \g452987/U$1 ( \26147 , \26145 , \26146 );
and \g452986/U$2 ( \26148 , \8414 , RIe1b5ec8_3447);
and \g452986/U$3 ( \26149 , RIfec50a0_8362, \8409 );
nor \g452986/U$1 ( \26150 , \26148 , \26149 );
and \g445332/U$2 ( \26151 , \26144 , \26147 , \26150 );
nor \g445332/U$1 ( \26152 , \26151 , \8481 );
and \g446255/U$2 ( \26153 , RIe1a4150_3244, \8371 );
and \g446255/U$3 ( \26154 , RIe21c3a8_4611, \8378 );
and \g449210/U$2 ( \26155 , RIe1f8fc0_4210, \8531 );
and \g449210/U$3 ( \26156 , \8488 , RIe1ffc08_4287);
and \g449210/U$4 ( \26157 , RIe1a6e50_3276, \8383 );
nor \g449210/U$1 ( \26158 , \26155 , \26156 , \26157 );
and \g452999/U$2 ( \26159 , \8335 , RIe171fc0_2674);
and \g452999/U$3 ( \26160 , RIe1d6010_3812, \8340 );
nor \g452999/U$1 ( \26161 , \26159 , \26160 );
and \g454873/U$2 ( \26162 , \8313 , RIe1af988_3375);
and \g454873/U$3 ( \26163 , RIe1bcb10_3524, \8323 );
nor \g454873/U$1 ( \26164 , \26162 , \26163 );
not \g454872/U$1 ( \26165 , \26164 );
and \g450225/U$2 ( \26166 , \26165 , \8316 );
and \g450225/U$3 ( \26167 , RIe1a9b50_3308, \8351 );
nor \g450225/U$1 ( \26168 , \26166 , \26167 );
and \g452997/U$2 ( \26169 , \8356 , RIe1f1b08_4127);
and \g452997/U$3 ( \26170 , RIe205ba8_4355, \8359 );
nor \g452997/U$1 ( \26171 , \26169 , \26170 );
nand \g448210/U$1 ( \26172 , \26158 , \26161 , \26168 , \26171 );
nor \g446255/U$1 ( \26173 , \26153 , \26154 , \26172 );
and \g452996/U$2 ( \26174 , \8404 , RIe1a1450_3212);
and \g452996/U$3 ( \26175 , RIe179e50_2764, \8409 );
nor \g452996/U$1 ( \26176 , \26174 , \26175 );
and \g452995/U$2 ( \26177 , \8412 , RIe2277a8_4739);
and \g452995/U$3 ( \26178 , RIe18d950_2988, \8417 );
nor \g452995/U$1 ( \26179 , \26177 , \26178 );
and \g445333/U$2 ( \26180 , \26173 , \26176 , \26179 );
nor \g445333/U$1 ( \26181 , \26180 , \8651 );
or \g444325/U$1 ( \26182 , \26062 , \26123 , \26152 , \26181 );
and \g446250/U$2 ( \26183 , RIfe9f558_8157, \8417 );
and \g446250/U$3 ( \26184 , RIe198d50_3116, \8404 );
and \g449202/U$2 ( \26185 , RIe17f850_2828, \8319 );
and \g449202/U$3 ( \26186 , \8326 , RIe182550_2860);
and \g449202/U$4 ( \26187 , RIe19ba50_3148, \8330 );
nor \g449202/U$1 ( \26188 , \26185 , \26186 , \26187 );
and \g452973/U$2 ( \26189 , \8335 , RIe17cb50_2796);
and \g452973/U$3 ( \26190 , RIf142ef8_5221, \8340 );
nor \g452973/U$1 ( \26191 , \26189 , \26190 );
and \g454919/U$2 ( \26192 , \8313 , RIfc47870_5836);
and \g454919/U$3 ( \26193 , RIe187f50_2924, \8323 );
nor \g454919/U$1 ( \26194 , \26192 , \26193 );
not \g450218/U$3 ( \26195 , \26194 );
not \g450218/U$4 ( \26196 , \8347 );
and \g450218/U$2 ( \26197 , \26195 , \26196 );
and \g450218/U$5 ( \26198 , \8351 , RIe19e750_3180);
nor \g450218/U$1 ( \26199 , \26197 , \26198 );
and \g452972/U$2 ( \26200 , \8356 , RIe185250_2892);
and \g452972/U$3 ( \26201 , RIe18ac50_2956, \8359 );
nor \g452972/U$1 ( \26202 , \26200 , \26201 );
nand \g447830/U$1 ( \26203 , \26188 , \26191 , \26199 , \26202 );
nor \g446250/U$1 ( \26204 , \26183 , \26184 , \26203 );
and \g452971/U$2 ( \26205 , \8378 , RIe190650_3020);
and \g452971/U$3 ( \26206 , RIfc479d8_5837, \8373 );
nor \g452971/U$1 ( \26207 , \26205 , \26206 );
and \g452969/U$2 ( \26208 , \8414 , RIe193350_3052);
and \g452969/U$3 ( \26209 , RIe196050_3084, \8409 );
nor \g452969/U$1 ( \26210 , \26208 , \26209 );
and \g445328/U$2 ( \26211 , \26204 , \26207 , \26210 );
nor \g445328/U$1 ( \26212 , \26211 , \8589 );
and \g446252/U$2 ( \26213 , RIe177588_2735, \8373 );
and \g446252/U$3 ( \26214 , RIfc7ee60_6466, \8319 );
and \g449205/U$2 ( \26215 , RIfce40f8_7617, \8414 );
and \g449205/U$3 ( \26216 , \8409 , RIfe9f3f0_8156);
and \g449205/U$4 ( \26217 , RIfcbc6c0_7166, \8383 );
nor \g449205/U$1 ( \26218 , \26215 , \26216 , \26217 );
and \g452984/U$2 ( \26219 , \8356 , RIe1745b8_2701);
and \g452984/U$3 ( \26220 , RIfc47438_5833, \8359 );
nor \g452984/U$1 ( \26221 , \26219 , \26220 );
and \g455138/U$2 ( \26222 , \8313 , RIfc99170_6764);
and \g455138/U$3 ( \26223 , RIfca15a0_6858, \8323 );
nor \g455138/U$1 ( \26224 , \26222 , \26223 );
not \g450221/U$3 ( \26225 , \26224 );
not \g450221/U$4 ( \26226 , \8347 );
and \g450221/U$2 ( \26227 , \26225 , \26226 );
and \g450221/U$5 ( \26228 , \8351 , RIfcb5208_7083);
nor \g450221/U$1 ( \26229 , \26227 , \26228 );
and \g452983/U$2 ( \26230 , \8378 , RIfc47708_5835);
and \g452983/U$3 ( \26231 , RIf13fdc0_5186, \8417 );
nor \g452983/U$1 ( \26232 , \26230 , \26231 );
nand \g447831/U$1 ( \26233 , \26218 , \26221 , \26229 , \26232 );
nor \g446252/U$1 ( \26234 , \26213 , \26214 , \26233 );
and \g452979/U$2 ( \26235 , \8335 , RIfce8e50_7672);
and \g452979/U$3 ( \26236 , RIfc8cc90_6624, \8340 );
nor \g452979/U$1 ( \26237 , \26235 , \26236 );
and \g452978/U$2 ( \26238 , \8324 , RIfc556a0_5994);
and \g452978/U$3 ( \26239 , RIe176610_2724, \8404 );
nor \g452978/U$1 ( \26240 , \26238 , \26239 );
and \g445331/U$2 ( \26241 , \26234 , \26237 , \26240 );
nor \g445331/U$1 ( \26242 , \26241 , \8558 );
or \g444280/U$1 ( \26243 , \26182 , \26212 , \26242 );
_DC \g4879/U$1 ( \26244 , \26243 , \8654 );
and \g447101/U$2 ( \26245 , \16438 , RIee2deb0_4981);
and \g447101/U$3 ( \26246 , RIee2eb58_4990, \16441 );
nor \g447101/U$1 ( \26247 , \26245 , \26246 );
and \g446334/U$2 ( \26248 , RIe141e88_2127, \16356 );
and \g446334/U$3 ( \26249 , RIe13fb60_2102, \16344 );
and \g449312/U$2 ( \26250 , RIee30070_5005, \16427 );
and \g449312/U$3 ( \26251 , \16398 , RIdf34288_1970);
and \g449312/U$4 ( \26252 , RIdf36880_1997, \16341 );
nor \g449312/U$1 ( \26253 , \26250 , \26251 , \26252 );
and \g453383/U$2 ( \26254 , \16361 , RIfe97dd0_8072);
and \g453383/U$3 ( \26255 , RIdf320c8_1946, \16364 );
nor \g453383/U$1 ( \26256 , \26254 , \26255 );
and \g453382/U$2 ( \26257 , \16377 , RIfc99878_6769);
and \g453382/U$3 ( \26258 , RIfc480e0_5842, \16313 );
nor \g453382/U$1 ( \26259 , \26257 , \26258 );
and \g455325/U$2 ( \26260 , \16317 , RIfc7fb08_6475);
and \g455325/U$3 ( \26261 , RIfc8be80_6614, \16325 );
nor \g455325/U$1 ( \26262 , \26260 , \26261 );
not \g450330/U$3 ( \26263 , \26262 );
not \g450330/U$4 ( \26264 , \16311 );
and \g450330/U$2 ( \26265 , \26263 , \26264 );
and \g450330/U$5 ( \26266 , \16448 , RIfe97f38_8073);
nor \g450330/U$1 ( \26267 , \26265 , \26266 );
nand \g447889/U$1 ( \26268 , \26253 , \26256 , \26259 , \26267 );
nor \g446334/U$1 ( \26269 , \26248 , \26249 , \26268 );
not \g444899/U$3 ( \26270 , \26269 );
not \g444899/U$4 ( \26271 , \16393 );
and \g444899/U$2 ( \26272 , \26270 , \26271 );
and \g446337/U$2 ( \26273 , RIee38068_5096, \16313 );
and \g446337/U$3 ( \26274 , RIe147720_2190, \16361 );
and \g449313/U$2 ( \26275 , RIe152b20_2318, \16427 );
and \g449313/U$3 ( \26276 , \16448 , RIfcbbe50_7160);
and \g449313/U$4 ( \26277 , RIe163920_2510, \16321 );
nor \g449313/U$1 ( \26278 , \26275 , \26276 , \26277 );
and \g453390/U$2 ( \26279 , \16368 , RIe14fe20_2286);
and \g453390/U$3 ( \26280 , RIfc47e10_5840, \16371 );
nor \g453390/U$1 ( \26281 , \26279 , \26280 );
and \g455326/U$2 ( \26282 , \16317 , RIe15df20_2446);
and \g455326/U$3 ( \26283 , RIfc48248_5843, \16325 );
nor \g455326/U$1 ( \26284 , \26282 , \26283 );
not \g450331/U$3 ( \26285 , \26284 );
not \g450331/U$4 ( \26286 , \16330 );
and \g450331/U$2 ( \26287 , \26285 , \26286 );
and \g450331/U$5 ( \26288 , \16328 , RIe166620_2542);
nor \g450331/U$1 ( \26289 , \26287 , \26288 );
and \g453389/U$2 ( \26290 , \16334 , RIe155820_2350);
and \g453389/U$3 ( \26291 , RIe158520_2382, \16380 );
nor \g453389/U$1 ( \26292 , \26290 , \26291 );
nand \g447890/U$1 ( \26293 , \26278 , \26281 , \26289 , \26292 );
nor \g446337/U$1 ( \26294 , \26273 , \26274 , \26293 );
and \g453388/U$2 ( \26295 , \16364 , RIe14a420_2222);
and \g453388/U$3 ( \26296 , RIfca0e98_6853, \16341 );
nor \g453388/U$1 ( \26297 , \26295 , \26296 );
and \g453387/U$2 ( \26298 , \16398 , RIe14d120_2254);
and \g453387/U$3 ( \26299 , RIe160c20_2478, \16377 );
nor \g453387/U$1 ( \26300 , \26298 , \26299 );
and \g445388/U$2 ( \26301 , \26294 , \26297 , \26300 );
nor \g445388/U$1 ( \26302 , \26301 , \16389 );
nor \g444899/U$1 ( \26303 , \26272 , \26302 );
and \g447102/U$2 ( \26304 , \16705 , RIdf3b5d8_2052);
and \g447102/U$3 ( \26305 , RIdf3da68_2078, \16707 );
nor \g447102/U$1 ( \26306 , \26304 , \26305 );
nand \g444432/U$1 ( \26307 , \26247 , \26303 , \26306 );
and \g453401/U$2 ( \26308 , \16377 , RIfc80210_6480);
and \g453401/U$3 ( \26309 , RIdf26f98_1820, \16380 );
nor \g453401/U$1 ( \26310 , \26308 , \26309 );
and \g446339/U$2 ( \26311 , RIfc48ab8_5849, \16321 );
and \g446339/U$3 ( \26312 , RIfce05e8_7575, \16313 );
and \g449317/U$2 ( \26313 , RIfc48950_5848, \16427 );
and \g449317/U$3 ( \26314 , \16448 , RIfc8bbb0_6612);
and \g449317/U$4 ( \26315 , RIdf29158_1844, \16485 );
nor \g449317/U$1 ( \26316 , \26313 , \26314 , \26315 );
and \g455331/U$2 ( \26317 , \16317 , RIdf208f0_1747);
and \g455331/U$3 ( \26318 , RIdf21f70_1763, \16325 );
nor \g455331/U$1 ( \26319 , \26317 , \26318 );
not \g455330/U$1 ( \26320 , \26319 );
and \g450335/U$2 ( \26321 , \26320 , \16336 );
and \g450335/U$3 ( \26322 , RIdf2b048_1866, \16356 );
nor \g450335/U$1 ( \26323 , \26321 , \26322 );
and \g453404/U$2 ( \26324 , \16361 , RIdf1a3b0_1675);
and \g453404/U$3 ( \26325 , RIdf1b8c8_1690, \16364 );
nor \g453404/U$1 ( \26326 , \26324 , \26325 );
and \g453403/U$2 ( \26327 , \16368 , RIfc8bd18_6613);
and \g453403/U$3 ( \26328 , RIdf235f0_1779, \16371 );
nor \g453403/U$1 ( \26329 , \26327 , \26328 );
nand \g448110/U$1 ( \26330 , \26316 , \26323 , \26326 , \26329 );
nor \g446339/U$1 ( \26331 , \26311 , \26312 , \26330 );
and \g453400/U$2 ( \26332 , \16334 , RIdf254e0_1801);
and \g453400/U$3 ( \26333 , RIfcc3740_7246, \16326 );
nor \g453400/U$1 ( \26334 , \26332 , \26333 );
nand \g445663/U$1 ( \26335 , \26310 , \26331 , \26334 );
and \g444835/U$2 ( \26336 , \26335 , \16481 );
and \g449314/U$2 ( \26337 , RIfcb5370_7084, \16427 );
and \g449314/U$3 ( \26338 , \16398 , RIded8230_923);
and \g449314/U$4 ( \26339 , RIdeda6c0_949, \16341 );
nor \g449314/U$1 ( \26340 , \26337 , \26338 , \26339 );
and \g453399/U$2 ( \26341 , \16361 , RIded3d48_874);
and \g453399/U$3 ( \26342 , RIded6070_899, \16364 );
nor \g453399/U$1 ( \26343 , \26341 , \26342 );
and \g453398/U$2 ( \26344 , \16377 , RIfca1168_6855);
and \g453398/U$3 ( \26345 , RIfc99710_6768, \16313 );
nor \g453398/U$1 ( \26346 , \26344 , \26345 );
and \g455327/U$2 ( \26347 , \16317 , RIfcd9838_7497);
and \g455327/U$3 ( \26348 , RIfcbc120_7162, \16325 );
nor \g455327/U$1 ( \26349 , \26347 , \26348 );
not \g450333/U$3 ( \26350 , \26349 );
not \g450333/U$4 ( \26351 , \16311 );
and \g450333/U$2 ( \26352 , \26350 , \26351 );
and \g450333/U$5 ( \26353 , \16432 , RIfc549f8_5985);
nor \g450333/U$1 ( \26354 , \26352 , \26353 );
nand \g447892/U$1 ( \26355 , \26340 , \26343 , \26346 , \26354 );
and \g444835/U$3 ( \26356 , \16477 , \26355 );
nor \g444835/U$1 ( \26357 , \26336 , \26356 );
and \g447105/U$2 ( \26358 , \17473 , RIfce0480_7574);
and \g447105/U$3 ( \26359 , RIfce43c8_7619, \17475 );
nor \g447105/U$1 ( \26360 , \26358 , \26359 );
and \g447104/U$2 ( \26361 , \22390 , RIdee3a68_1054);
and \g447104/U$3 ( \26362 , RIdee57f0_1075, \22392 );
nor \g447104/U$1 ( \26363 , \26361 , \26362 );
and \g447106/U$2 ( \26364 , \18278 , RIdedf850_1007);
and \g447106/U$3 ( \26365 , RIdee18a8_1030, \18280 );
nor \g447106/U$1 ( \26366 , \26364 , \26365 );
nand \g444652/U$1 ( \26367 , \26357 , \26360 , \26363 , \26366 );
and \g446332/U$2 ( \26368 , RIfce4698_7621, \16313 );
and \g446332/U$3 ( \26369 , RIe16a400_2586, \16364 );
and \g449307/U$2 ( \26370 , RIfcbba18_7157, \16427 );
and \g449307/U$3 ( \26371 , \16448 , RIde82e20_228);
and \g449307/U$4 ( \26372 , RIfe98208_8075, \16321 );
nor \g449307/U$1 ( \26373 , \26370 , \26371 , \26372 );
and \g453374/U$2 ( \26374 , \16368 , RIfc99f80_6774);
and \g453374/U$3 ( \26375 , RIfc48d88_5851, \16371 );
nor \g453374/U$1 ( \26376 , \26374 , \26375 );
and \g455226/U$2 ( \26377 , \16317 , RIde8f648_289);
and \g455226/U$3 ( \26378 , RIde93158_307, \16325 );
nor \g455226/U$1 ( \26379 , \26377 , \26378 );
not \g450326/U$3 ( \26380 , \26379 );
not \g450326/U$4 ( \26381 , \16330 );
and \g450326/U$2 ( \26382 , \26380 , \26381 );
and \g450326/U$5 ( \26383 , \16328 , RIfcd9c70_7500);
nor \g450326/U$1 ( \26384 , \26382 , \26383 );
and \g453373/U$2 ( \26385 , \16334 , RIde87308_249);
and \g453373/U$3 ( \26386 , RIde8b4a8_269, \16380 );
nor \g453373/U$1 ( \26387 , \26385 , \26386 );
nand \g447887/U$1 ( \26388 , \26373 , \26376 , \26384 , \26387 );
nor \g446332/U$1 ( \26389 , \26368 , \26369 , \26388 );
and \g453371/U$2 ( \26390 , \16341 , RIfc8b4a8_6607);
and \g453371/U$3 ( \26391 , RIfe980a0_8074, \16377 );
nor \g453371/U$1 ( \26392 , \26390 , \26391 );
and \g453372/U$2 ( \26393 , \16361 , RIe168c18_2569);
and \g453372/U$3 ( \26394 , RIe16c728_2611, \16398 );
nor \g453372/U$1 ( \26395 , \26393 , \26394 );
and \g445385/U$2 ( \26396 , \26389 , \26392 , \26395 );
nor \g445385/U$1 ( \26397 , \26396 , \16649 );
and \g446333/U$2 ( \26398 , RIfc80eb8_6489, \16356 );
and \g446333/U$3 ( \26399 , RIdeb8520_561, \16334 );
and \g449309/U$2 ( \26400 , RIdeb2b20_497, \16427 );
and \g449309/U$3 ( \26401 , \16337 , RIdeacec8_433);
and \g449309/U$4 ( \26402 , RIfc491c0_5854, \16341 );
nor \g449309/U$1 ( \26403 , \26400 , \26401 , \26402 );
and \g453380/U$2 ( \26404 , \16361 , RIde9fcc8_369);
and \g453380/U$3 ( \26405 , RIdea65c8_401, \16364 );
nor \g453380/U$1 ( \26406 , \26404 , \26405 );
and \g453379/U$2 ( \26407 , \16377 , RIdec0c20_657);
and \g453379/U$3 ( \26408 , RIfc49328_5855, \16313 );
nor \g453379/U$1 ( \26409 , \26407 , \26408 );
and \g455321/U$2 ( \26410 , \16317 , RIdec3920_689);
and \g455321/U$3 ( \26411 , RIdec6620_721, \16325 );
nor \g455321/U$1 ( \26412 , \26410 , \26411 );
not \g450329/U$3 ( \26413 , \26412 );
not \g450329/U$4 ( \26414 , \16311 );
and \g450329/U$2 ( \26415 , \26413 , \26414 );
and \g450329/U$5 ( \26416 , \16448 , RIfc80648_6483);
nor \g450329/U$1 ( \26417 , \26415 , \26416 );
nand \g447888/U$1 ( \26418 , \26403 , \26406 , \26409 , \26417 );
nor \g446333/U$1 ( \26419 , \26398 , \26399 , \26418 );
and \g453376/U$2 ( \26420 , \16371 , RIfc8b340_6606);
and \g453376/U$3 ( \26421 , RIdebb220_593, \16380 );
nor \g453376/U$1 ( \26422 , \26420 , \26421 );
and \g453377/U$2 ( \26423 , \16368 , RIdeafe20_465);
and \g453377/U$3 ( \26424 , RIdebdf20_625, \16485 );
nor \g453377/U$1 ( \26425 , \26423 , \26424 );
and \g445387/U$2 ( \26426 , \26419 , \26422 , \26425 );
nor \g445387/U$1 ( \26427 , \26426 , \16618 );
or \g444311/U$1 ( \26428 , \26307 , \26367 , \26397 , \26427 );
and \g446330/U$2 ( \26429 , RIdefbff0_1331, \16427 );
and \g446330/U$3 ( \26430 , RIdef65f0_1267, \16368 );
and \g449304/U$2 ( \26431 , RIdf154f0_1619, \16321 );
and \g449304/U$3 ( \26432 , \16328 , RIdf181f0_1651);
and \g449304/U$4 ( \26433 , RIdef0bf0_1203, \16398 );
nor \g449304/U$1 ( \26434 , \26431 , \26432 , \26433 );
and \g455319/U$2 ( \26435 , \16317 , RIdf0a0f0_1491);
and \g455319/U$3 ( \26436 , RIdf0cdf0_1523, \16325 );
nor \g455319/U$1 ( \26437 , \26435 , \26436 );
not \g450321/U$3 ( \26438 , \26437 );
not \g450321/U$4 ( \26439 , \16330 );
and \g450321/U$2 ( \26440 , \26438 , \26439 );
and \g450321/U$5 ( \26441 , \16341 , RIdef38f0_1235);
nor \g450321/U$1 ( \26442 , \26440 , \26441 );
and \g453363/U$2 ( \26443 , \16377 , RIdf0faf0_1555);
and \g453363/U$3 ( \26444 , RIdf127f0_1587, \16313 );
nor \g453363/U$1 ( \26445 , \26443 , \26444 );
and \g453364/U$2 ( \26446 , \16334 , RIdf046f0_1427);
and \g453364/U$3 ( \26447 , RIdf073f0_1459, \16380 );
nor \g453364/U$1 ( \26448 , \26446 , \26447 );
nand \g447413/U$1 ( \26449 , \26434 , \26442 , \26445 , \26448 );
nor \g446330/U$1 ( \26450 , \26429 , \26430 , \26449 );
and \g453362/U$2 ( \26451 , \16361 , RIdeeb1f0_1139);
and \g453362/U$3 ( \26452 , RIdefecf0_1363, \16448 );
nor \g453362/U$1 ( \26453 , \26451 , \26452 );
and \g453361/U$2 ( \26454 , \16364 , RIdeedef0_1171);
and \g453361/U$3 ( \26455 , RIdef92f0_1299, \16371 );
nor \g453361/U$1 ( \26456 , \26454 , \26455 );
and \g445383/U$2 ( \26457 , \26450 , \26453 , \26456 );
nor \g445383/U$1 ( \26458 , \26457 , \16555 );
and \g446331/U$2 ( \26459 , RIdf39418_2028, \16427 );
and \g446331/U$3 ( \26460 , RIdf1e2f8_1720, \16368 );
and \g449305/U$2 ( \26461 , RIde993c8_337, \16485 );
and \g449305/U$3 ( \26462 , \16356 , RIdeb5820_529);
and \g449305/U$4 ( \26463 , RIdee84f0_1107, \16398 );
nor \g449305/U$1 ( \26464 , \26461 , \26462 , \26463 );
and \g455229/U$2 ( \26465 , \16317 , RIdeced20_817);
and \g455229/U$3 ( \26466 , RIded1a20_849, \16325 );
nor \g455229/U$1 ( \26467 , \26465 , \26466 );
not \g450324/U$3 ( \26468 , \26467 );
not \g450324/U$4 ( \26469 , \16311 );
and \g450324/U$2 ( \26470 , \26468 , \26469 );
and \g450324/U$5 ( \26471 , \16341 , RIdf019f0_1395);
nor \g450324/U$1 ( \26472 , \26470 , \26471 );
and \g453369/U$2 ( \26473 , \16377 , RIdec9320_753);
and \g453369/U$3 ( \26474 , RIdecc020_785, \16313 );
nor \g453369/U$1 ( \26475 , \26473 , \26474 );
and \g453370/U$2 ( \26476 , \16334 , RIe15b220_2414);
and \g453370/U$3 ( \26477 , RIe16f428_2643, \16380 );
nor \g453370/U$1 ( \26478 , \26476 , \26477 );
nand \g447414/U$1 ( \26479 , \26464 , \26472 , \26475 , \26478 );
nor \g446331/U$1 ( \26480 , \26459 , \26460 , \26479 );
and \g453368/U$2 ( \26481 , \16361 , RIde7f310_210);
and \g453368/U$3 ( \26482 , RIe144a20_2158, \16448 );
nor \g453368/U$1 ( \26483 , \26481 , \26482 );
and \g453367/U$2 ( \26484 , \16364 , RIdedd258_980);
and \g453367/U$3 ( \26485 , RIdf2da78_1896, \16371 );
nor \g453367/U$1 ( \26486 , \26484 , \26485 );
and \g445384/U$2 ( \26487 , \26480 , \26483 , \26486 );
nor \g445384/U$1 ( \26488 , \26487 , \16586 );
or \g444221/U$1 ( \26489 , \26428 , \26458 , \26488 );
_DC \g48fe/U$1 ( \26490 , \26489 , \16652 );
and \g453441/U$2 ( \26491 , \8414 , RIe1934b8_3053);
and \g453441/U$3 ( \26492 , RIe1961b8_3085, \8407 );
nor \g453441/U$1 ( \26493 , \26491 , \26492 );
and \g446347/U$2 ( \26494 , RIf144c80_5242, \8417 );
and \g446347/U$3 ( \26495 , RIe1853b8_2893, \8356 );
and \g449328/U$2 ( \26496 , RIe17f9b8_2829, \8319 );
and \g449328/U$3 ( \26497 , \8326 , RIe1826b8_2861);
and \g449328/U$4 ( \26498 , RIe1880b8_2925, \8488 );
nor \g449328/U$1 ( \26499 , \26496 , \26497 , \26498 );
and \g453445/U$2 ( \26500 , \8335 , RIe17ccb8_2797);
and \g453445/U$3 ( \26501 , RIfcc3fb0_7252, \8340 );
nor \g453445/U$1 ( \26502 , \26500 , \26501 );
and \g453444/U$2 ( \26503 , \8404 , RIe198eb8_3117);
and \g453444/U$3 ( \26504 , RIe19e8b8_3181, \8351 );
nor \g453444/U$1 ( \26505 , \26503 , \26504 );
and \g455207/U$2 ( \26506 , \8313 , RIfe976c8_8067);
and \g455207/U$3 ( \26507 , RIe19bbb8_3149, \8323 );
nor \g455207/U$1 ( \26508 , \26506 , \26507 );
not \g450345/U$3 ( \26509 , \26508 );
not \g450345/U$4 ( \26510 , \8328 );
and \g450345/U$2 ( \26511 , \26509 , \26510 );
and \g450345/U$5 ( \26512 , \8359 , RIe18adb8_2957);
nor \g450345/U$1 ( \26513 , \26511 , \26512 );
nand \g447900/U$1 ( \26514 , \26499 , \26502 , \26505 , \26513 );
nor \g446347/U$1 ( \26515 , \26494 , \26495 , \26514 );
and \g453442/U$2 ( \26516 , \8378 , RIe1907b8_3021);
and \g453442/U$3 ( \26517 , RIfe97560_8066, \8531 );
nor \g453442/U$1 ( \26518 , \26516 , \26517 );
nand \g445664/U$1 ( \26519 , \26493 , \26515 , \26518 );
and \g444730/U$2 ( \26520 , \26519 , \9702 );
and \g449326/U$2 ( \26521 , RIfcc4118_7253, \8373 );
and \g449326/U$3 ( \26522 , \8330 , RIf1412d8_5201);
and \g449326/U$4 ( \26523 , RIfc89e28_6591, \8488 );
nor \g449326/U$1 ( \26524 , \26521 , \26522 , \26523 );
and \g453439/U$2 ( \26525 , \8335 , RIfcd5d28_7455);
and \g453439/U$3 ( \26526 , RIfc4a408_5867, \8340 );
nor \g453439/U$1 ( \26527 , \26525 , \26526 );
and \g453438/U$2 ( \26528 , \8404 , RIfe97830_8068);
and \g453438/U$3 ( \26529 , RIfcd3730_7428, \8351 );
nor \g453438/U$1 ( \26530 , \26528 , \26529 );
and \g455406/U$2 ( \26531 , \8313 , RIfc530a8_5967);
and \g455406/U$3 ( \26532 , RIfce27a8_7599, \8323 );
nor \g455406/U$1 ( \26533 , \26531 , \26532 );
not \g455405/U$1 ( \26534 , \26533 );
and \g450343/U$2 ( \26535 , \26534 , \8316 );
and \g450343/U$3 ( \26536 , RIfcc3e48_7251, \8359 );
nor \g450343/U$1 ( \26537 , \26535 , \26536 );
nand \g448225/U$1 ( \26538 , \26524 , \26527 , \26530 , \26537 );
and \g444730/U$3 ( \26539 , \9700 , \26538 );
nor \g444730/U$1 ( \26540 , \26520 , \26539 );
and \g447108/U$2 ( \26541 , \12254 , RIfc9fae8_6839);
and \g447108/U$3 ( \26542 , RIfc9f980_6838, \12256 );
nor \g447108/U$1 ( \26543 , \26541 , \26542 );
nor \g448302/U$1 ( \26544 , \8558 , \8408 );
and \g447107/U$2 ( \26545 , \26544 , RIf13f6b8_5181);
nor \g448301/U$1 ( \26546 , \8558 , \8433 );
and \g447107/U$3 ( \26547 , RIfc4a6d8_5869, \26546 );
nor \g447107/U$1 ( \26548 , \26545 , \26547 );
and \g447109/U$2 ( \26549 , \12264 , RIe174720_2702);
and \g447109/U$3 ( \26550 , RIfc89cc0_6590, \12266 );
nor \g447109/U$1 ( \26551 , \26549 , \26550 );
nand \g444529/U$1 ( \26552 , \26540 , \26543 , \26548 , \26551 );
and \g453453/U$2 ( \26553 , \8326 , RIe1bcc78_3525);
and \g453453/U$3 ( \26554 , RIe1a15b8_3213, \8404 );
nor \g453453/U$1 ( \26555 , \26553 , \26554 );
and \g446350/U$2 ( \26556 , RIe1a42b8_3245, \8371 );
and \g446350/U$3 ( \26557 , RIe1afaf0_3376, \8319 );
and \g449331/U$2 ( \26558 , RIe227910_4740, \8412 );
and \g449331/U$3 ( \26559 , \8409 , RIe179fb8_2765);
and \g449331/U$4 ( \26560 , RIe1a6fb8_3277, \8383 );
nor \g449331/U$1 ( \26561 , \26558 , \26559 , \26560 );
and \g453457/U$2 ( \26562 , \8356 , RIe1f1c70_4128);
and \g453457/U$3 ( \26563 , RIe205d10_4356, \8359 );
nor \g453457/U$1 ( \26564 , \26562 , \26563 );
and \g455202/U$2 ( \26565 , \8313 , RIe1f9128_4211);
and \g455202/U$3 ( \26566 , RIe1ffd70_4288, \8323 );
nor \g455202/U$1 ( \26567 , \26565 , \26566 );
not \g450348/U$3 ( \26568 , \26567 );
not \g450348/U$4 ( \26569 , \8347 );
and \g450348/U$2 ( \26570 , \26568 , \26569 );
and \g450348/U$5 ( \26571 , \8351 , RIe1a9cb8_3309);
nor \g450348/U$1 ( \26572 , \26570 , \26571 );
and \g453456/U$2 ( \26573 , \8378 , RIe21c510_4612);
and \g453456/U$3 ( \26574 , RIe18dab8_2989, \8417 );
nor \g453456/U$1 ( \26575 , \26573 , \26574 );
nand \g447903/U$1 ( \26576 , \26561 , \26564 , \26572 , \26575 );
nor \g446350/U$1 ( \26577 , \26556 , \26557 , \26576 );
and \g453454/U$2 ( \26578 , \8335 , RIe172128_2675);
and \g453454/U$3 ( \26579 , RIe1d6178_3813, \8340 );
nor \g453454/U$1 ( \26580 , \26578 , \26579 );
nand \g445665/U$1 ( \26581 , \26555 , \26577 , \26580 );
and \g444885/U$2 ( \26582 , \26581 , \9010 );
and \g449329/U$2 ( \26583 , RIe1ad228_3347, \8319 );
and \g449329/U$3 ( \26584 , \8326 , RIfc81188_6491);
and \g449329/U$4 ( \26585 , RIfcc3a10_7248, \8486 );
nor \g449329/U$1 ( \26586 , \26583 , \26584 , \26585 );
and \g453449/U$2 ( \26587 , \8335 , RIe1aba40_3330);
and \g453449/U$3 ( \26588 , RIfc495f8_5857, \8340 );
nor \g453449/U$1 ( \26589 , \26587 , \26588 );
and \g453448/U$2 ( \26590 , \8404 , RIe1b81f0_3472);
and \g453448/U$3 ( \26591 , RIfc49a30_5860, \8351 );
nor \g453448/U$1 ( \26592 , \26590 , \26591 );
and \g455205/U$2 ( \26593 , \8313 , RIe1ba3b0_3496);
and \g455205/U$3 ( \26594 , RIfcb6018_7093, \8323 );
nor \g455205/U$1 ( \26595 , \26593 , \26594 );
not \g450346/U$3 ( \26596 , \26595 );
not \g450346/U$4 ( \26597 , \8328 );
and \g450346/U$2 ( \26598 , \26596 , \26597 );
and \g450346/U$5 ( \26599 , \8359 , RIfce5610_7632);
nor \g450346/U$1 ( \26600 , \26598 , \26599 );
nand \g447901/U$1 ( \26601 , \26586 , \26589 , \26592 , \26600 );
and \g444885/U$3 ( \26602 , \8482 , \26601 );
nor \g444885/U$1 ( \26603 , \26582 , \26602 );
and \g447110/U$2 ( \26604 , \8964 , RIfcbb5e0_7154);
and \g447110/U$3 ( \26605 , RIfce0a20_7578, \8966 );
nor \g447110/U$1 ( \26606 , \26604 , \26605 );
and \g447111/U$2 ( \26607 , \8521 , RIe1b19e0_3398);
and \g447111/U$3 ( \26608 , RIe1b3330_3416, \8525 );
nor \g447111/U$1 ( \26609 , \26607 , \26608 );
and \g447112/U$2 ( \26610 , \8974 , RIfe97998_8069);
and \g447112/U$3 ( \26611 , RIe1b6030_3448, \8976 );
nor \g447112/U$1 ( \26612 , \26610 , \26611 );
nand \g444654/U$1 ( \26613 , \26603 , \26606 , \26609 , \26612 );
and \g446343/U$2 ( \26614 , RIfcd5e90_7456, \8373 );
and \g446343/U$3 ( \26615 , RIfcbb310_7152, \8319 );
and \g449322/U$2 ( \26616 , RIfc9a520_6778, \8531 );
and \g449322/U$3 ( \26617 , \8488 , RIfcb62e8_7095);
and \g449322/U$4 ( \26618 , RIfc81890_6496, \8383 );
nor \g449322/U$1 ( \26619 , \26616 , \26617 , \26618 );
and \g453425/U$2 ( \26620 , \8356 , RIe1f4268_4155);
and \g453425/U$3 ( \26621 , RIfcd3460_7426, \8359 );
nor \g453425/U$1 ( \26622 , \26620 , \26621 );
and \g455213/U$2 ( \26623 , \8313 , RIfcbb1a8_7151);
and \g455213/U$3 ( \26624 , RIfc81728_6495, \8323 );
nor \g455213/U$1 ( \26625 , \26623 , \26624 );
not \g450340/U$3 ( \26626 , \26625 );
not \g450340/U$4 ( \26627 , \8376 );
and \g450340/U$2 ( \26628 , \26626 , \26627 );
and \g450340/U$5 ( \26629 , \8351 , RIfc9a7f0_6780);
nor \g450340/U$1 ( \26630 , \26628 , \26629 );
and \g453424/U$2 ( \26631 , \8378 , RIe1f66f8_4181);
and \g453424/U$3 ( \26632 , RIfc49e68_5863, \8417 );
nor \g453424/U$1 ( \26633 , \26631 , \26632 );
nand \g447896/U$1 ( \26634 , \26619 , \26622 , \26630 , \26633 );
nor \g446343/U$1 ( \26635 , \26614 , \26615 , \26634 );
and \g453422/U$2 ( \26636 , \8335 , RIe1ef0d8_4097);
and \g453422/U$3 ( \26637 , RIfc49d00_5862, \8340 );
nor \g453422/U$1 ( \26638 , \26636 , \26637 );
and \g453421/U$2 ( \26639 , \8326 , RIfcd9dd8_7501);
and \g453421/U$3 ( \26640 , RIe1fb180_4234, \8404 );
nor \g453421/U$1 ( \26641 , \26639 , \26640 );
and \g445394/U$2 ( \26642 , \26635 , \26638 , \26641 );
nor \g445394/U$1 ( \26643 , \26642 , \8621 );
and \g446346/U$2 ( \26644 , RIe1d8e78_3845, \8378 );
and \g446346/U$3 ( \26645 , RIe1c8078_3653, \8340 );
and \g449324/U$2 ( \26646 , RIe1de878_3909, \8409 );
and \g449324/U$3 ( \26647 , \8373 , RIe1e6f78_4005);
and \g449324/U$4 ( \26648 , RIe1e9c78_4037, \8330 );
nor \g449324/U$1 ( \26649 , \26646 , \26647 , \26648 );
and \g454147/U$2 ( \26650 , \8313 , RIe1cda78_3717);
and \g454147/U$3 ( \26651 , RIe1d0778_3749, \8323 );
nor \g454147/U$1 ( \26652 , \26650 , \26651 );
not \g450341/U$3 ( \26653 , \26652 );
not \g450341/U$4 ( \26654 , \8347 );
and \g450341/U$2 ( \26655 , \26653 , \26654 );
and \g450341/U$5 ( \26656 , \8417 , RIe1e1578_3941);
nor \g450341/U$1 ( \26657 , \26655 , \26656 );
and \g453430/U$2 ( \26658 , \8404 , RIe1e4278_3973);
and \g453430/U$3 ( \26659 , RIe1ec978_4069, \8351 );
nor \g453430/U$1 ( \26660 , \26658 , \26659 );
and \g453431/U$2 ( \26661 , \8356 , RIe1cad78_3685);
and \g453431/U$3 ( \26662 , RIe1d3478_3781, \8359 );
nor \g453431/U$1 ( \26663 , \26661 , \26662 );
nand \g447898/U$1 ( \26664 , \26649 , \26657 , \26660 , \26663 );
nor \g446346/U$1 ( \26665 , \26644 , \26645 , \26664 );
and \g453429/U$2 ( \26666 , \8335 , RIe1bf978_3557);
and \g453429/U$3 ( \26667 , RIe1dbb78_3877, \8414 );
nor \g453429/U$1 ( \26668 , \26666 , \26667 );
and \g453428/U$2 ( \26669 , \8317 , RIe1c2678_3589);
and \g453428/U$3 ( \26670 , RIe1c5378_3621, \8326 );
nor \g453428/U$1 ( \26671 , \26669 , \26670 );
and \g445395/U$2 ( \26672 , \26665 , \26668 , \26671 );
nor \g445395/U$1 ( \26673 , \26672 , \8477 );
or \g444378/U$1 ( \26674 , \26552 , \26613 , \26643 , \26673 );
and \g446341/U$2 ( \26675 , RIfc53210_5968, \8371 );
and \g446341/U$3 ( \26676 , RIe20b710_4420, \8319 );
and \g449318/U$2 ( \26677 , RIf1699b8_5661, \8531 );
and \g449318/U$3 ( \26678 , \8488 , RIe213e10_4516);
and \g449318/U$4 ( \26679 , RIe224c10_4708, \8330 );
nor \g449318/U$1 ( \26680 , \26677 , \26678 , \26679 );
and \g453411/U$2 ( \26681 , \8356 , RIe211110_4484);
and \g453411/U$3 ( \26682 , RIfc401d8_5755, \8359 );
nor \g453411/U$1 ( \26683 , \26681 , \26682 );
and \g455332/U$2 ( \26684 , \8313 , RIe219810_4580);
and \g455332/U$3 ( \26685 , RIe21f210_4644, \8323 );
nor \g455332/U$1 ( \26686 , \26684 , \26685 );
not \g450336/U$3 ( \26687 , \26686 );
not \g450336/U$4 ( \26688 , \8376 );
and \g450336/U$2 ( \26689 , \26687 , \26688 );
and \g450336/U$5 ( \26690 , \8351 , RIf16cf28_5699);
nor \g450336/U$1 ( \26691 , \26689 , \26690 );
and \g453410/U$2 ( \26692 , \8378 , RIe216b10_4548);
and \g453410/U$3 ( \26693 , RIf16b1a0_5678, \8417 );
nor \g453410/U$1 ( \26694 , \26692 , \26693 );
nand \g447893/U$1 ( \26695 , \26680 , \26683 , \26691 , \26694 );
nor \g446341/U$1 ( \26696 , \26675 , \26676 , \26695 );
and \g453408/U$2 ( \26697 , \8335 , RIe208a10_4388);
and \g453408/U$3 ( \26698 , RIfc81cc8_6499, \8340 );
nor \g453408/U$1 ( \26699 , \26697 , \26698 );
and \g453407/U$2 ( \26700 , \8326 , RIe20e410_4452);
and \g453407/U$3 ( \26701 , RIe221f10_4676, \8404 );
nor \g453407/U$1 ( \26702 , \26700 , \26701 );
and \g445391/U$2 ( \26703 , \26696 , \26699 , \26702 );
nor \g445391/U$1 ( \26704 , \26703 , \8368 );
and \g446342/U$2 ( \26705 , RIfc53378_5969, \8417 );
and \g446342/U$3 ( \26706 , RIfe97b00_8070, \8356 );
and \g449321/U$2 ( \26707 , RIfc8a800_6598, \8319 );
and \g449321/U$3 ( \26708 , \8326 , RIfe97c68_8071);
and \g449321/U$4 ( \26709 , RIf15ecc0_5538, \8488 );
nor \g449321/U$1 ( \26710 , \26707 , \26708 , \26709 );
and \g453417/U$2 ( \26711 , \8335 , RIfc8a698_6597);
and \g453417/U$3 ( \26712 , RIfc8a530_6596, \8340 );
nor \g453417/U$1 ( \26713 , \26711 , \26712 );
and \g453416/U$2 ( \26714 , \8404 , RIe201828_4307);
and \g453416/U$3 ( \26715 , RIfc8a0f8_6593, \8351 );
nor \g453416/U$1 ( \26716 , \26714 , \26715 );
and \g455217/U$2 ( \26717 , \8313 , RIe203448_4327);
and \g455217/U$3 ( \26718 , RIfcb6720_7098, \8323 );
nor \g455217/U$1 ( \26719 , \26717 , \26718 );
not \g450338/U$3 ( \26720 , \26719 );
not \g450338/U$4 ( \26721 , \8328 );
and \g450338/U$2 ( \26722 , \26720 , \26721 );
and \g450338/U$5 ( \26723 , \8359 , RIf160bb0_5560);
nor \g450338/U$1 ( \26724 , \26722 , \26723 );
nand \g447895/U$1 ( \26725 , \26710 , \26713 , \26716 , \26724 );
nor \g446342/U$1 ( \26726 , \26705 , \26706 , \26725 );
and \g453415/U$2 ( \26727 , \8378 , RIfc49fd0_5864);
and \g453415/U$3 ( \26728 , RIe1fd4a8_4259, \8531 );
nor \g453415/U$1 ( \26729 , \26727 , \26728 );
and \g453414/U$2 ( \26730 , \8414 , RIfcb65b8_7097);
and \g453414/U$3 ( \26731 , RIfc8a3c8_6595, \8409 );
nor \g453414/U$1 ( \26732 , \26730 , \26731 );
and \g445392/U$2 ( \26733 , \26726 , \26729 , \26732 );
nor \g445392/U$1 ( \26734 , \26733 , \8422 );
or \g444249/U$1 ( \26735 , \26674 , \26704 , \26734 );
_DC \g4982/U$1 ( \26736 , \26735 , \8654 );
and \g444434/U$2 ( \26737 , RIfe99cc0_8094, \17284 );
and \g444434/U$3 ( \26738 , RIdf1ba30_1691, \17286 );
and \g446360/U$2 ( \26739 , RIdf0cf58_1524, \16356 );
and \g446360/U$3 ( \26740 , RIdf04858_1428, \16334 );
and \g449340/U$2 ( \26741 , RIdefc158_1332, \16427 );
and \g449340/U$3 ( \26742 , \16398 , RIdef0d58_1204);
and \g449340/U$4 ( \26743 , RIdef3a58_1236, \16339 );
nor \g449340/U$1 ( \26744 , \26741 , \26742 , \26743 );
and \g453493/U$2 ( \26745 , \16361 , RIdeeb358_1140);
and \g453493/U$3 ( \26746 , RIdeee058_1172, \16364 );
nor \g453493/U$1 ( \26747 , \26745 , \26746 );
and \g453492/U$2 ( \26748 , \16377 , RIdf0fc58_1556);
and \g453492/U$3 ( \26749 , RIdf12958_1588, \16313 );
nor \g453492/U$1 ( \26750 , \26748 , \26749 );
and \g455054/U$2 ( \26751 , \16317 , RIdf15658_1620);
and \g455054/U$3 ( \26752 , RIdf18358_1652, \16325 );
nor \g455054/U$1 ( \26753 , \26751 , \26752 );
not \g450361/U$3 ( \26754 , \26753 );
not \g450361/U$4 ( \26755 , \16311 );
and \g450361/U$2 ( \26756 , \26754 , \26755 );
and \g450361/U$5 ( \26757 , \16432 , RIdefee58_1364);
nor \g450361/U$1 ( \26758 , \26756 , \26757 );
nand \g447911/U$1 ( \26759 , \26744 , \26747 , \26750 , \26758 );
nor \g446360/U$1 ( \26760 , \26739 , \26740 , \26759 );
and \g453489/U$2 ( \26761 , \16368 , RIdef6758_1268);
and \g453489/U$3 ( \26762 , RIdf0a258_1492, \16344 );
nor \g453489/U$1 ( \26763 , \26761 , \26762 );
and \g453024/U$2 ( \26764 , \16371 , RIdef9458_1300);
and \g453024/U$3 ( \26765 , RIdf07558_1460, \16380 );
nor \g453024/U$1 ( \26766 , \26764 , \26765 );
and \g445670/U$1 ( \26767 , \26760 , \26763 , \26766 );
or \g444668/U$2 ( \26768 , \26767 , \16555 );
and \g446358/U$2 ( \26769 , RIdf220d8_1764, \16339 );
and \g446358/U$3 ( \26770 , RIdf20a58_1748, \16398 );
and \g449339/U$2 ( \26771 , RIfcb6e28_7103, \16321 );
and \g449339/U$3 ( \26772 , \16485 , RIdf292c0_1845);
and \g449339/U$4 ( \26773 , RIdf2b1b0_1867, \16356 );
nor \g449339/U$1 ( \26774 , \26771 , \26772 , \26773 );
and \g453484/U$2 ( \26775 , \16368 , RIfc82da8_6511);
and \g453484/U$3 ( \26776 , RIdf23758_1780, \16371 );
nor \g453484/U$1 ( \26777 , \26775 , \26776 );
and \g455212/U$2 ( \26778 , \16317 , RIfc4a9a8_5871);
and \g455212/U$3 ( \26779 , RIfc9ac28_6783, \16325 );
nor \g455212/U$1 ( \26780 , \26778 , \26779 );
not \g450359/U$3 ( \26781 , \26780 );
not \g450359/U$4 ( \26782 , \16351 );
and \g450359/U$2 ( \26783 , \26781 , \26782 );
and \g450359/U$5 ( \26784 , \16328 , RIfc83078_6513);
nor \g450359/U$1 ( \26785 , \26783 , \26784 );
and \g453483/U$2 ( \26786 , \16334 , RIfe999f0_8092);
and \g453483/U$3 ( \26787 , RIfe99b58_8093, \16380 );
nor \g453483/U$1 ( \26788 , \26786 , \26787 );
nand \g447909/U$1 ( \26789 , \26774 , \26777 , \26785 , \26788 );
nor \g446358/U$1 ( \26790 , \26769 , \26770 , \26789 );
or \g444668/U$3 ( \26791 , \16480 , \26790 );
and \g447118/U$2 ( \26792 , \16518 , RIfcbad70_7148);
and \g447118/U$3 ( \26793 , RIfc9ad90_6784, \16521 );
nor \g447118/U$1 ( \26794 , \26792 , \26793 );
nand \g444668/U$1 ( \26795 , \26768 , \26791 , \26794 );
nor \g444434/U$1 ( \26796 , \26737 , \26738 , \26795 );
and \g453459/U$2 ( \26797 , \16334 , RIe155988_2351);
and \g453459/U$3 ( \26798 , RIfc895b8_6585, \16371 );
nor \g453459/U$1 ( \26799 , \26797 , \26798 );
and \g446351/U$2 ( \26800 , RIe15e088_2447, \16485 );
and \g446351/U$3 ( \26801 , RIe158688_2383, \16380 );
and \g449332/U$2 ( \26802 , RIe163a88_2511, \16321 );
and \g449332/U$3 ( \26803 , \16328 , RIe166788_2543);
and \g449332/U$4 ( \26804 , RIe152c88_2319, \16427 );
nor \g449332/U$1 ( \26805 , \26802 , \26803 , \26804 );
and \g453462/U$2 ( \26806 , \16361 , RIe147888_2191);
and \g453462/U$3 ( \26807 , RIe14a588_2223, \16364 );
nor \g453462/U$1 ( \26808 , \26806 , \26807 );
and \g453461/U$2 ( \26809 , \16377 , RIe160d88_2479);
and \g453461/U$3 ( \26810 , RIfc83618_6517, \16313 );
nor \g453461/U$1 ( \26811 , \26809 , \26810 );
and \g455345/U$2 ( \26812 , \16317 , RIe14d288_2255);
and \g455345/U$3 ( \26813 , RIfc51cf8_5953, \16325 );
nor \g455345/U$1 ( \26814 , \26812 , \26813 );
not \g455344/U$1 ( \26815 , \26814 );
and \g450349/U$2 ( \26816 , \26815 , \16336 );
and \g450349/U$3 ( \26817 , RIfc3f800_5748, \16448 );
nor \g450349/U$1 ( \26818 , \26816 , \26817 );
nand \g448111/U$1 ( \26819 , \26805 , \26808 , \26811 , \26818 );
nor \g446351/U$1 ( \26820 , \26800 , \26801 , \26819 );
and \g453458/U$2 ( \26821 , \16368 , RIe14ff88_2287);
and \g453458/U$3 ( \26822 , RIee36718_5078, \16356 );
nor \g453458/U$1 ( \26823 , \26821 , \26822 );
nand \g445666/U$1 ( \26824 , \26799 , \26820 , \26823 );
and \g444674/U$2 ( \26825 , \26824 , \16390 );
and \g446353/U$2 ( \26826 , RIfe99888_8091, \16354 );
and \g446353/U$3 ( \26827 , RIfe995b8_8089, \16334 );
and \g449334/U$2 ( \26828 , RIfcc43e8_7255, \16427 );
and \g449334/U$3 ( \26829 , \16398 , RIe16c890_2612);
and \g449334/U$4 ( \26830 , RIfcc5798_7269, \16341 );
nor \g449334/U$1 ( \26831 , \26828 , \26829 , \26830 );
and \g453469/U$2 ( \26832 , \16361 , RIe168d80_2570);
and \g453469/U$3 ( \26833 , RIe16a568_2587, \16364 );
nor \g453469/U$1 ( \26834 , \26832 , \26833 );
and \g453467/U$2 ( \26835 , \16377 , RIee1aef0_4765);
and \g453467/U$3 ( \26836 , RIee1b5f8_4770, \16313 );
nor \g453467/U$1 ( \26837 , \26835 , \26836 );
and \g455360/U$2 ( \26838 , \16317 , RIee1c570_4781);
and \g455360/U$3 ( \26839 , RIee1d650_4793, \16325 );
nor \g455360/U$1 ( \26840 , \26838 , \26839 );
not \g450351/U$3 ( \26841 , \26840 );
not \g450351/U$4 ( \26842 , \16311 );
and \g450351/U$2 ( \26843 , \26841 , \26842 );
and \g450351/U$5 ( \26844 , \16448 , RIde83168_229);
nor \g450351/U$1 ( \26845 , \26843 , \26844 );
nand \g447904/U$1 ( \26846 , \26831 , \26834 , \26837 , \26845 );
nor \g446353/U$1 ( \26847 , \26826 , \26827 , \26846 );
and \g453465/U$2 ( \26848 , \16371 , RIfcd5a58_7453);
and \g453465/U$3 ( \26849 , RIfe99720_8090, \16380 );
nor \g453465/U$1 ( \26850 , \26848 , \26849 );
and \g453466/U$2 ( \26851 , \16368 , RIfc89450_6584);
and \g453466/U$3 ( \26852 , RIfe99450_8088, \16344 );
nor \g453466/U$1 ( \26853 , \26851 , \26852 );
and \g445400/U$2 ( \26854 , \26847 , \26850 , \26853 );
nor \g445400/U$1 ( \26855 , \26854 , \16649 );
nor \g444674/U$1 ( \26856 , \26825 , \26855 );
and \g453478/U$2 ( \26857 , \16398 , RIdee8658_1108);
and \g453478/U$3 ( \26858 , RIdec9488_754, \16377 );
nor \g453478/U$1 ( \26859 , \26857 , \26858 );
and \g446356/U$2 ( \26860 , RIdecc188_786, \16313 );
and \g446356/U$3 ( \26861 , RIde7f658_211, \16361 );
and \g449337/U$2 ( \26862 , RIdf39580_2029, \16427 );
and \g449337/U$3 ( \26863 , \16448 , RIe144b88_2159);
and \g449337/U$4 ( \26864 , RIdecee88_818, \16321 );
nor \g449337/U$1 ( \26865 , \26862 , \26863 , \26864 );
and \g453481/U$2 ( \26866 , \16368 , RIdf1e460_1721);
and \g453481/U$3 ( \26867 , RIdf2dbe0_1897, \16371 );
nor \g453481/U$1 ( \26868 , \26866 , \26867 );
and \g455297/U$2 ( \26869 , \16317 , RIde99710_338);
and \g455297/U$3 ( \26870 , RIdeb5988_530, \16325 );
nor \g455297/U$1 ( \26871 , \26869 , \26870 );
not \g450357/U$3 ( \26872 , \26871 );
not \g450357/U$4 ( \26873 , \16330 );
and \g450357/U$2 ( \26874 , \26872 , \26873 );
and \g450357/U$5 ( \26875 , \16326 , RIded1b88_850);
nor \g450357/U$1 ( \26876 , \26874 , \26875 );
and \g453480/U$2 ( \26877 , \16334 , RIe15b388_2415);
and \g453480/U$3 ( \26878 , RIe16f590_2644, \16380 );
nor \g453480/U$1 ( \26879 , \26877 , \26878 );
nand \g447908/U$1 ( \26880 , \26865 , \26868 , \26876 , \26879 );
nor \g446356/U$1 ( \26881 , \26860 , \26861 , \26880 );
and \g453479/U$2 ( \26882 , \16364 , RIdedd3c0_981);
and \g453479/U$3 ( \26883 , RIdf01b58_1396, \16341 );
nor \g453479/U$1 ( \26884 , \26882 , \26883 );
nand \g445668/U$1 ( \26885 , \26859 , \26881 , \26884 );
and \g444675/U$2 ( \26886 , \26885 , \16752 );
and \g453474/U$2 ( \26887 , \16398 , RIded8398_924);
and \g453474/U$3 ( \26888 , RIfc826a0_6506, \16377 );
nor \g453474/U$1 ( \26889 , \26887 , \26888 );
and \g446354/U$2 ( \26890 , RIfc52568_5959, \16313 );
and \g446354/U$3 ( \26891 , RIded3eb0_875, \16361 );
and \g449336/U$2 ( \26892 , RIfc89b58_6589, \16427 );
and \g449336/U$3 ( \26893 , \16448 , RIfce4800_7622);
and \g449336/U$4 ( \26894 , RIee24b08_4876, \16319 );
nor \g449336/U$1 ( \26895 , \26892 , \26893 , \26894 );
and \g453477/U$2 ( \26896 , \16368 , RIfc82538_6505);
and \g453477/U$3 ( \26897 , RIfc9f3e0_6834, \16371 );
nor \g453477/U$1 ( \26898 , \26896 , \26897 );
and \g455239/U$2 ( \26899 , \16317 , RIdee3bd0_1055);
and \g455239/U$3 ( \26900 , RIdee5958_1076, \16325 );
nor \g455239/U$1 ( \26901 , \26899 , \26900 );
not \g450354/U$3 ( \26902 , \26901 );
not \g450354/U$4 ( \26903 , \16330 );
and \g450354/U$2 ( \26904 , \26902 , \26903 );
and \g450354/U$5 ( \26905 , \16326 , RIee25918_4886);
nor \g450354/U$1 ( \26906 , \26904 , \26905 );
and \g453476/U$2 ( \26907 , \16334 , RIdedf9b8_1008);
and \g453476/U$3 ( \26908 , RIfe99f90_8096, \16380 );
nor \g453476/U$1 ( \26909 , \26907 , \26908 );
nand \g447906/U$1 ( \26910 , \26895 , \26898 , \26906 , \26909 );
nor \g446354/U$1 ( \26911 , \26890 , \26891 , \26910 );
and \g453475/U$2 ( \26912 , \16364 , RIfeabe70_8272);
and \g453475/U$3 ( \26913 , RIdeda828_950, \16341 );
nor \g453475/U$1 ( \26914 , \26912 , \26913 );
nand \g445667/U$1 ( \26915 , \26889 , \26911 , \26914 );
and \g444675/U$3 ( \26916 , \16477 , \26915 );
nor \g444675/U$1 ( \26917 , \26886 , \26916 );
and \g444435/U$2 ( \26918 , RIfe99e28_8095, \16419 );
and \g444435/U$3 ( \26919 , RIdf32230_1947, \16422 );
and \g446363/U$2 ( \26920 , RIfc892e8_6583, \16341 );
and \g446363/U$3 ( \26921 , RIdec0d88_658, \16377 );
and \g449344/U$2 ( \26922 , RIdec3a88_690, \16321 );
and \g449344/U$3 ( \26923 , \16485 , RIdebe088_626);
and \g449344/U$4 ( \26924 , RIee1f810_4817, \16356 );
nor \g449344/U$1 ( \26925 , \26922 , \26923 , \26924 );
and \g453505/U$2 ( \26926 , \16368 , RIdeaff88_466);
and \g453505/U$3 ( \26927 , RIfce1f38_7593, \16371 );
nor \g453505/U$1 ( \26928 , \26926 , \26927 );
and \g454973/U$2 ( \26929 , \16317 , RIdeb2c88_498);
and \g454973/U$3 ( \26930 , RIfc9b1c8_6787, \16325 );
nor \g454973/U$1 ( \26931 , \26929 , \26930 );
not \g450363/U$3 ( \26932 , \26931 );
not \g450363/U$4 ( \26933 , \16351 );
and \g450363/U$2 ( \26934 , \26932 , \26933 );
and \g450363/U$5 ( \26935 , \16328 , RIdec6788_722);
nor \g450363/U$1 ( \26936 , \26934 , \26935 );
and \g453504/U$2 ( \26937 , \16334 , RIdeb8688_562);
and \g453504/U$3 ( \26938 , RIdebb388_594, \16380 );
nor \g453504/U$1 ( \26939 , \26937 , \26938 );
nand \g447913/U$1 ( \26940 , \26925 , \26928 , \26936 , \26939 );
nor \g446363/U$1 ( \26941 , \26920 , \26921 , \26940 );
and \g453501/U$2 ( \26942 , \16364 , RIdea6910_402);
and \g453501/U$3 ( \26943 , RIdead210_434, \16398 );
nor \g453501/U$1 ( \26944 , \26942 , \26943 );
and \g453500/U$2 ( \26945 , \16361 , RIdea0010_370);
and \g453500/U$3 ( \26946 , RIee20788_4828, \16313 );
nor \g453500/U$1 ( \26947 , \26945 , \26946 );
and \g445671/U$1 ( \26948 , \26941 , \26944 , \26947 );
or \g444669/U$2 ( \26949 , \26948 , \16618 );
and \g446361/U$2 ( \26950 , RIdf369e8_1998, \16341 );
and \g446361/U$3 ( \26951 , RIdf343f0_1971, \16398 );
and \g449343/U$2 ( \26952 , RIee301d8_5006, \16427 );
and \g449343/U$3 ( \26953 , \16448 , RIfcb6f90_7104);
and \g449343/U$4 ( \26954 , RIee338b0_5045, \16321 );
nor \g449343/U$1 ( \26955 , \26952 , \26953 , \26954 );
and \g453496/U$2 ( \26956 , \16368 , RIee2e018_4982);
and \g453496/U$3 ( \26957 , RIfcba938_7145, \16371 );
nor \g453496/U$1 ( \26958 , \26956 , \26957 );
and \g455339/U$2 ( \26959 , \16317 , RIe13fcc8_2103);
and \g455339/U$3 ( \26960 , RIe141ff0_2128, \16325 );
nor \g455339/U$1 ( \26961 , \26959 , \26960 );
not \g450362/U$3 ( \26962 , \26961 );
not \g450362/U$4 ( \26963 , \16330 );
and \g450362/U$2 ( \26964 , \26962 , \26963 );
and \g450362/U$5 ( \26965 , \16328 , RIee34990_5057);
nor \g450362/U$1 ( \26966 , \26964 , \26965 );
and \g453495/U$2 ( \26967 , \16334 , RIdf3b740_2053);
and \g453495/U$3 ( \26968 , RIdf3dbd0_2079, \16380 );
nor \g453495/U$1 ( \26969 , \26967 , \26968 );
nand \g447912/U$1 ( \26970 , \26955 , \26958 , \26966 , \26969 );
nor \g446361/U$1 ( \26971 , \26950 , \26951 , \26970 );
or \g444669/U$3 ( \26972 , \16393 , \26971 );
and \g447119/U$2 ( \26973 , \16715 , RIfcd3b68_7431);
and \g447119/U$3 ( \26974 , RIfc831e0_6514, \16717 );
nor \g447119/U$1 ( \26975 , \26973 , \26974 );
nand \g444669/U$1 ( \26976 , \26949 , \26972 , \26975 );
nor \g444435/U$1 ( \26977 , \26918 , \26919 , \26976 );
nand \g444160/U$1 ( \26978 , \26796 , \26856 , \26917 , \26977 );
_DC \g4a07/U$1 ( \26979 , \26978 , \16652 );
and \g453542/U$2 ( \26980 , \8531 , RIe1cdbe0_3718);
and \g453542/U$3 ( \26981 , RIe1dbce0_3878, \8414 );
nor \g453542/U$1 ( \26982 , \26980 , \26981 );
and \g446371/U$2 ( \26983 , RIe1de9e0_3910, \8409 );
and \g446371/U$3 ( \26984 , RIe1d8fe0_3846, \8378 );
and \g449354/U$2 ( \26985 , RIe1e70e0_4006, \8373 );
and \g449354/U$3 ( \26986 , \8383 , RIe1e9de0_4038);
and \g449354/U$4 ( \26987 , RIe1d08e0_3750, \8488 );
nor \g449354/U$1 ( \26988 , \26985 , \26986 , \26987 );
and \g453546/U$2 ( \26989 , \8335 , RIe1bfae0_3558);
and \g453546/U$3 ( \26990 , RIe1c81e0_3654, \8340 );
nor \g453546/U$1 ( \26991 , \26989 , \26990 );
and \g453544/U$2 ( \26992 , \8404 , RIe1e43e0_3974);
and \g453544/U$3 ( \26993 , RIe1ecae0_4070, \8351 );
nor \g453544/U$1 ( \26994 , \26992 , \26993 );
and \g455343/U$2 ( \26995 , \8313 , RIe1c27e0_3590);
and \g455343/U$3 ( \26996 , RIe1c54e0_3622, \8323 );
nor \g455343/U$1 ( \26997 , \26995 , \26996 );
not \g455342/U$1 ( \26998 , \26997 );
and \g450376/U$2 ( \26999 , \26998 , \8316 );
and \g450376/U$3 ( \27000 , RIe1d35e0_3782, \8359 );
nor \g450376/U$1 ( \27001 , \26999 , \27000 );
nand \g448229/U$1 ( \27002 , \26988 , \26991 , \26994 , \27001 );
nor \g446371/U$1 ( \27003 , \26983 , \26984 , \27002 );
and \g453543/U$2 ( \27004 , \8356 , RIe1caee0_3686);
and \g453543/U$3 ( \27005 , RIe1e16e0_3942, \8417 );
nor \g453543/U$1 ( \27006 , \27004 , \27005 );
nand \g445673/U$1 ( \27007 , \26982 , \27003 , \27006 );
and \g444800/U$2 ( \27008 , \27007 , \8478 );
and \g449353/U$2 ( \27009 , RIfca3a30_6884, \8373 );
and \g449353/U$3 ( \27010 , \8383 , RIf158078_5461);
and \g449353/U$4 ( \27011 , RIf1520d8_5393, \8488 );
nor \g449353/U$1 ( \27012 , \27009 , \27010 , \27011 );
and \g453538/U$2 ( \27013 , \8335 , RIe1ef240_4098);
and \g453538/U$3 ( \27014 , RIf14fdb0_5368, \8340 );
nor \g453538/U$1 ( \27015 , \27013 , \27014 );
and \g453537/U$2 ( \27016 , \8404 , RIfea7988_8223);
and \g453537/U$3 ( \27017 , RIf1592c0_5474, \8351 );
nor \g453537/U$1 ( \27018 , \27016 , \27017 );
and \g455182/U$2 ( \27019 , \8313 , RIf14e2f8_5349);
and \g455182/U$3 ( \27020 , RIfcd2380_7414, \8323 );
nor \g455182/U$1 ( \27021 , \27019 , \27020 );
not \g455181/U$1 ( \27022 , \27021 );
and \g450374/U$2 ( \27023 , \27022 , \8316 );
and \g450374/U$3 ( \27024 , RIf1538c0_5410, \8359 );
nor \g450374/U$1 ( \27025 , \27023 , \27024 );
nand \g448227/U$1 ( \27026 , \27012 , \27015 , \27018 , \27025 );
and \g444800/U$3 ( \27027 , \8752 , \27026 );
nor \g444800/U$1 ( \27028 , \27008 , \27027 );
and \g447124/U$2 ( \27029 , \11516 , RIf155be8_5435);
and \g447124/U$3 ( \27030 , RIf156728_5443, \11518 );
nor \g447124/U$1 ( \27031 , \27029 , \27030 );
and \g447125/U$2 ( \27032 , \13486 , RIe1f43d0_4156);
and \g447125/U$3 ( \27033 , RIf150e90_5380, \13488 );
nor \g447125/U$1 ( \27034 , \27032 , \27033 );
and \g447127/U$2 ( \27035 , \11521 , RIfe98a78_8081);
and \g447127/U$3 ( \27036 , RIf154b08_5423, \11523 );
nor \g447127/U$1 ( \27037 , \27035 , \27036 );
nand \g444532/U$1 ( \27038 , \27028 , \27031 , \27034 , \27037 );
and \g453553/U$2 ( \27039 , \8356 , RIe1b1b48_3399);
and \g453553/U$3 ( \27040 , RIf149f78_5301, \8409 );
nor \g453553/U$1 ( \27041 , \27039 , \27040 );
and \g446373/U$2 ( \27042 , RIfe99180_8086, \8412 );
and \g446373/U$3 ( \27043 , RIf14a950_5308, \8417 );
and \g449359/U$2 ( \27044 , RIfe992e8_8087, \8373 );
and \g449359/U$3 ( \27045 , \8383 , RIf14bd00_5322);
and \g449359/U$4 ( \27046 , RIfcec7f8_7713, \8488 );
nor \g449359/U$1 ( \27047 , \27044 , \27045 , \27046 );
and \g453557/U$2 ( \27048 , \8335 , RIfe99018_8085);
and \g453557/U$3 ( \27049 , RIfc4b650_5880, \8340 );
nor \g453557/U$1 ( \27050 , \27048 , \27049 );
and \g453555/U$2 ( \27051 , \8404 , RIfe987a8_8079);
and \g453555/U$3 ( \27052 , RIfc44b70_5804, \8351 );
nor \g453555/U$1 ( \27053 , \27051 , \27052 );
and \g455171/U$2 ( \27054 , \8313 , RIfe98370_8076);
and \g455171/U$3 ( \27055 , RIfcda918_7509, \8323 );
nor \g455171/U$1 ( \27056 , \27054 , \27055 );
not \g455170/U$1 ( \27057 , \27056 );
and \g450379/U$2 ( \27058 , \27057 , \8316 );
and \g450379/U$3 ( \27059 , RIf149438_5293, \8359 );
nor \g450379/U$1 ( \27060 , \27058 , \27059 );
nand \g448230/U$1 ( \27061 , \27047 , \27050 , \27053 , \27060 );
nor \g446373/U$1 ( \27062 , \27042 , \27043 , \27061 );
and \g453552/U$2 ( \27063 , \8378 , RIfe98640_8078);
and \g453552/U$3 ( \27064 , RIfe984d8_8077, \8523 );
nor \g453552/U$1 ( \27065 , \27063 , \27064 );
nand \g445674/U$1 ( \27066 , \27041 , \27062 , \27065 );
and \g444923/U$2 ( \27067 , \27066 , \8482 );
and \g449357/U$2 ( \27068 , RIe227a78_4741, \8414 );
and \g449357/U$3 ( \27069 , \8407 , RIe17a120_2766);
and \g449357/U$4 ( \27070 , RIe1a7120_3278, \8330 );
nor \g449357/U$1 ( \27071 , \27068 , \27069 , \27070 );
and \g453550/U$2 ( \27072 , \8356 , RIe1f1dd8_4129);
and \g453550/U$3 ( \27073 , RIe205e78_4357, \8359 );
nor \g453550/U$1 ( \27074 , \27072 , \27073 );
and \g454687/U$2 ( \27075 , \8313 , RIe1f9290_4212);
and \g454687/U$3 ( \27076 , RIe1ffed8_4289, \8323 );
nor \g454687/U$1 ( \27077 , \27075 , \27076 );
not \g450378/U$3 ( \27078 , \27077 );
not \g450378/U$4 ( \27079 , \8347 );
and \g450378/U$2 ( \27080 , \27078 , \27079 );
and \g450378/U$5 ( \27081 , \8351 , RIe1a9e20_3310);
nor \g450378/U$1 ( \27082 , \27080 , \27081 );
and \g453549/U$2 ( \27083 , \8378 , RIe21c678_4613);
and \g453549/U$3 ( \27084 , RIe18dc20_2990, \8417 );
nor \g453549/U$1 ( \27085 , \27083 , \27084 );
nand \g447921/U$1 ( \27086 , \27071 , \27074 , \27082 , \27085 );
and \g444923/U$3 ( \27087 , \9010 , \27086 );
nor \g444923/U$1 ( \27088 , \27067 , \27087 );
and \g447128/U$2 ( \27089 , \9041 , RIe1a1720_3214);
and \g447128/U$3 ( \27090 , RIe1a4420_3246, \9043 );
nor \g447128/U$1 ( \27091 , \27089 , \27090 );
and \g447129/U$2 ( \27092 , \13239 , RIe1bcde0_3526);
and \g447129/U$3 ( \27093 , RIe1d62e0_3814, \13241 );
nor \g447129/U$1 ( \27094 , \27092 , \27093 );
and \g447130/U$2 ( \27095 , \13244 , RIe172290_2676);
and \g447130/U$3 ( \27096 , RIe1afc58_3377, \13246 );
nor \g447130/U$1 ( \27097 , \27095 , \27096 );
nand \g444656/U$1 ( \27098 , \27088 , \27091 , \27094 , \27097 );
and \g446367/U$2 ( \27099 , RIe21f378_4645, \8409 );
and \g446367/U$3 ( \27100 , RIe216c78_4549, \8378 );
and \g449350/U$2 ( \27101 , RIf16c280_5690, \8373 );
and \g449350/U$3 ( \27102 , \8383 , RIe224d78_4709);
and \g449350/U$4 ( \27103 , RIe213f78_4517, \8488 );
nor \g449350/U$1 ( \27104 , \27101 , \27102 , \27103 );
and \g453523/U$2 ( \27105 , \8335 , RIe208b78_4389);
and \g453523/U$3 ( \27106 , RIf1681d0_5644, \8340 );
nor \g453523/U$1 ( \27107 , \27105 , \27106 );
and \g453522/U$2 ( \27108 , \8404 , RIe222078_4677);
and \g453522/U$3 ( \27109 , RIfe98d48_8083, \8351 );
nor \g453522/U$1 ( \27110 , \27108 , \27109 );
and \g455187/U$2 ( \27111 , \8313 , RIe20b878_4421);
and \g455187/U$3 ( \27112 , RIe20e578_4453, \8323 );
nor \g455187/U$1 ( \27113 , \27111 , \27112 );
not \g455186/U$1 ( \27114 , \27113 );
and \g450369/U$2 ( \27115 , \27114 , \8316 );
and \g450369/U$3 ( \27116 , RIf16a390_5668, \8359 );
nor \g450369/U$1 ( \27117 , \27115 , \27116 );
nand \g448226/U$1 ( \27118 , \27104 , \27107 , \27110 , \27117 );
nor \g446367/U$1 ( \27119 , \27099 , \27100 , \27118 );
and \g453521/U$2 ( \27120 , \8356 , RIe211278_4485);
and \g453521/U$3 ( \27121 , RIf16b308_5679, \8417 );
nor \g453521/U$1 ( \27122 , \27120 , \27121 );
and \g453520/U$2 ( \27123 , \8531 , RIf169b20_5662);
and \g453520/U$3 ( \27124 , RIe219978_4581, \8414 );
nor \g453520/U$1 ( \27125 , \27123 , \27124 );
and \g445405/U$2 ( \27126 , \27119 , \27122 , \27125 );
nor \g445405/U$1 ( \27127 , \27126 , \8368 );
and \g446368/U$2 ( \27128 , RIfc70ec8_6307, \8417 );
and \g446368/U$3 ( \27129 , RIfe98eb0_8084, \8356 );
and \g449351/U$2 ( \27130 , RIfcd4540_7438, \8319 );
and \g449351/U$3 ( \27131 , \8324 , RIf15bcf0_5504);
and \g449351/U$4 ( \27132 , RIf15ee28_5539, \8488 );
nor \g449351/U$1 ( \27133 , \27130 , \27131 , \27132 );
and \g453531/U$2 ( \27134 , \8335 , RIf159e00_5482);
and \g453531/U$3 ( \27135 , RIf15d0a0_5518, \8340 );
nor \g453531/U$1 ( \27136 , \27134 , \27135 );
and \g453530/U$2 ( \27137 , \8404 , RIe201990_4308);
and \g453530/U$3 ( \27138 , RIfcd4ae0_7442, \8351 );
nor \g453530/U$1 ( \27139 , \27137 , \27138 );
and \g455183/U$2 ( \27140 , \8313 , RIfeab060_8262);
and \g455183/U$3 ( \27141 , RIfc61478_6129, \8323 );
nor \g455183/U$1 ( \27142 , \27140 , \27141 );
not \g450372/U$3 ( \27143 , \27142 );
not \g450372/U$4 ( \27144 , \8328 );
and \g450372/U$2 ( \27145 , \27143 , \27144 );
and \g450372/U$5 ( \27146 , \8359 , RIf160d18_5561);
nor \g450372/U$1 ( \27147 , \27145 , \27146 );
nand \g447918/U$1 ( \27148 , \27133 , \27136 , \27139 , \27147 );
nor \g446368/U$1 ( \27149 , \27128 , \27129 , \27148 );
and \g453527/U$2 ( \27150 , \8378 , RIfcbe880_7190);
and \g453527/U$3 ( \27151 , RIfe98be0_8082, \8523 );
nor \g453527/U$1 ( \27152 , \27150 , \27151 );
and \g453526/U$2 ( \27153 , \8414 , RIfcec528_7711);
and \g453526/U$3 ( \27154 , RIfc70928_6303, \8407 );
nor \g453526/U$1 ( \27155 , \27153 , \27154 );
and \g445407/U$2 ( \27156 , \27149 , \27152 , \27155 );
nor \g445407/U$1 ( \27157 , \27156 , \8422 );
or \g444373/U$1 ( \27158 , \27038 , \27098 , \27127 , \27157 );
and \g446364/U$2 ( \27159 , RIf145928_5251, \8373 );
and \g446364/U$3 ( \27160 , RIe17fb20_2830, \8319 );
and \g449346/U$2 ( \27161 , RIf143e70_5232, \8531 );
and \g449346/U$3 ( \27162 , \8488 , RIe188220_2926);
and \g449346/U$4 ( \27163 , RIe19bd20_3150, \8330 );
nor \g449346/U$1 ( \27164 , \27161 , \27162 , \27163 );
and \g453514/U$2 ( \27165 , \8356 , RIe185520_2894);
and \g453514/U$3 ( \27166 , RIe18af20_2958, \8359 );
nor \g453514/U$1 ( \27167 , \27165 , \27166 );
and \g454138/U$2 ( \27168 , \8313 , RIe193620_3054);
and \g454138/U$3 ( \27169 , RIe196320_3086, \8323 );
nor \g454138/U$1 ( \27170 , \27168 , \27169 );
not \g450365/U$3 ( \27171 , \27170 );
not \g450365/U$4 ( \27172 , \8376 );
and \g450365/U$2 ( \27173 , \27171 , \27172 );
and \g450365/U$5 ( \27174 , \8351 , RIe19ea20_3182);
nor \g450365/U$1 ( \27175 , \27173 , \27174 );
and \g453513/U$2 ( \27176 , \8378 , RIe190920_3022);
and \g453513/U$3 ( \27177 , RIfe98910_8080, \8417 );
nor \g453513/U$1 ( \27178 , \27176 , \27177 );
nand \g447915/U$1 ( \27179 , \27164 , \27167 , \27175 , \27178 );
nor \g446364/U$1 ( \27180 , \27159 , \27160 , \27179 );
and \g453511/U$2 ( \27181 , \8335 , RIe17ce20_2798);
and \g453511/U$3 ( \27182 , RIfc95c00_6726, \8340 );
nor \g453511/U$1 ( \27183 , \27181 , \27182 );
and \g453510/U$2 ( \27184 , \8326 , RIe182820_2862);
and \g453510/U$3 ( \27185 , RIe199020_3118, \8404 );
nor \g453510/U$1 ( \27186 , \27184 , \27185 );
and \g445403/U$2 ( \27187 , \27180 , \27183 , \27186 );
nor \g445403/U$1 ( \27188 , \27187 , \8589 );
and \g446366/U$2 ( \27189 , RIe1776f0_2736, \8373 );
and \g446366/U$3 ( \27190 , RIf16e878_5717, \8317 );
and \g449349/U$2 ( \27191 , RIee3e710_5169, \8414 );
and \g449349/U$3 ( \27192 , \8407 , RIfc62dc8_6147);
and \g449349/U$4 ( \27193 , RIf141440_5202, \8383 );
nor \g449349/U$1 ( \27194 , \27191 , \27192 , \27193 );
and \g453518/U$2 ( \27195 , \8356 , RIe174888_2703);
and \g453518/U$3 ( \27196 , RIee3c820_5147, \8359 );
nor \g453518/U$1 ( \27197 , \27195 , \27196 );
and \g455192/U$2 ( \27198 , \8313 , RIee3a390_5121);
and \g455192/U$3 ( \27199 , RIee3b470_5133, \8323 );
nor \g455192/U$1 ( \27200 , \27198 , \27199 );
not \g450368/U$3 ( \27201 , \27200 );
not \g450368/U$4 ( \27202 , \8347 );
and \g450368/U$2 ( \27203 , \27201 , \27202 );
and \g450368/U$5 ( \27204 , \8351 , RIf142520_5214);
nor \g450368/U$1 ( \27205 , \27203 , \27204 );
and \g453517/U$2 ( \27206 , \8378 , RIfc9cb18_6805);
and \g453517/U$3 ( \27207 , RIfcc5bd0_7272, \8417 );
nor \g453517/U$1 ( \27208 , \27206 , \27207 );
nand \g447916/U$1 ( \27209 , \27194 , \27197 , \27205 , \27208 );
nor \g446366/U$1 ( \27210 , \27189 , \27190 , \27209 );
and \g453516/U$2 ( \27211 , \8335 , RIfc6ea38_6281);
and \g453516/U$3 ( \27212 , RIf170498_5737, \8340 );
nor \g453516/U$1 ( \27213 , \27211 , \27212 );
and \g453515/U$2 ( \27214 , \8326 , RIfc68660_6210);
and \g453515/U$3 ( \27215 , RIfeab8d0_8268, \8404 );
nor \g453515/U$1 ( \27216 , \27214 , \27215 );
and \g445404/U$2 ( \27217 , \27210 , \27213 , \27216 );
nor \g445404/U$1 ( \27218 , \27217 , \8558 );
or \g444283/U$1 ( \27219 , \27158 , \27188 , \27218 );
_DC \g4a8b/U$1 ( \27220 , \27219 , \8654 );
and \g453878/U$2 ( \27221 , \16371 , RIdef95c0_1301);
and \g453878/U$3 ( \27222 , RIdefc2c0_1333, \16427 );
nor \g453878/U$1 ( \27223 , \27221 , \27222 );
and \g446442/U$2 ( \27224 , RIdefefc0_1365, \16448 );
and \g446442/U$3 ( \27225 , RIdeeb4c0_1141, \16361 );
and \g449446/U$2 ( \27226 , RIdf0a3c0_1493, \16485 );
and \g449446/U$3 ( \27227 , \16356 , RIdf0d0c0_1525);
and \g449446/U$4 ( \27228 , RIdef0ec0_1205, \16398 );
nor \g449446/U$1 ( \27229 , \27226 , \27227 , \27228 );
and \g455388/U$2 ( \27230 , \16317 , RIdf157c0_1621);
and \g455388/U$3 ( \27231 , RIdf184c0_1653, \16325 );
nor \g455388/U$1 ( \27232 , \27230 , \27231 );
not \g450467/U$3 ( \27233 , \27232 );
not \g450467/U$4 ( \27234 , \16311 );
and \g450467/U$2 ( \27235 , \27233 , \27234 );
and \g450467/U$5 ( \27236 , \16341 , RIdef3bc0_1237);
nor \g450467/U$1 ( \27237 , \27235 , \27236 );
and \g453880/U$2 ( \27238 , \16377 , RIdf0fdc0_1557);
and \g453880/U$3 ( \27239 , RIdf12ac0_1589, \16313 );
nor \g453880/U$1 ( \27240 , \27238 , \27239 );
and \g453881/U$2 ( \27241 , \16334 , RIdf049c0_1429);
and \g453881/U$3 ( \27242 , RIdf076c0_1461, \16380 );
nor \g453881/U$1 ( \27243 , \27241 , \27242 );
nand \g447433/U$1 ( \27244 , \27229 , \27237 , \27240 , \27243 );
nor \g446442/U$1 ( \27245 , \27224 , \27225 , \27244 );
and \g453879/U$2 ( \27246 , \16364 , RIdeee1c0_1173);
and \g453879/U$3 ( \27247 , RIdef68c0_1269, \16368 );
nor \g453879/U$1 ( \27248 , \27246 , \27247 );
nand \g445691/U$1 ( \27249 , \27223 , \27245 , \27248 );
and \g444807/U$2 ( \27250 , \27249 , \16750 );
and \g449444/U$2 ( \27251 , RIdeceff0_819, \16321 );
and \g449444/U$3 ( \27252 , \16328 , RIded1cf0_851);
and \g449444/U$4 ( \27253 , RIdee87c0_1109, \16398 );
nor \g449444/U$1 ( \27254 , \27251 , \27252 , \27253 );
and \g454890/U$2 ( \27255 , \16317 , RIde99a58_339);
and \g454890/U$3 ( \27256 , RIdeb5af0_531, \16325 );
nor \g454890/U$1 ( \27257 , \27255 , \27256 );
not \g450464/U$3 ( \27258 , \27257 );
not \g450464/U$4 ( \27259 , \16330 );
and \g450464/U$2 ( \27260 , \27258 , \27259 );
and \g450464/U$5 ( \27261 , \16341 , RIdf01cc0_1397);
nor \g450464/U$1 ( \27262 , \27260 , \27261 );
and \g453871/U$2 ( \27263 , \16377 , RIdec95f0_755);
and \g453871/U$3 ( \27264 , RIdecc2f0_787, \16313 );
nor \g453871/U$1 ( \27265 , \27263 , \27264 );
and \g453872/U$2 ( \27266 , \16334 , RIe15b4f0_2416);
and \g453872/U$3 ( \27267 , RIe16f6f8_2645, \16380 );
nor \g453872/U$1 ( \27268 , \27266 , \27267 );
nand \g447432/U$1 ( \27269 , \27254 , \27262 , \27265 , \27268 );
and \g444807/U$3 ( \27270 , \16752 , \27269 );
nor \g444807/U$1 ( \27271 , \27250 , \27270 );
and \g447187/U$2 ( \27272 , \16774 , RIde7f9a0_212);
and \g447187/U$3 ( \27273 , RIdedd528_982, \16776 );
nor \g447187/U$1 ( \27274 , \27272 , \27273 );
and \g447186/U$2 ( \27275 , \16779 , RIdf1e5c8_1722);
and \g447186/U$3 ( \27276 , RIdf2dd48_1898, \16781 );
nor \g447186/U$1 ( \27277 , \27275 , \27276 );
and \g447185/U$2 ( \27278 , \16784 , RIdf396e8_2030);
and \g447185/U$3 ( \27279 , RIe144cf0_2160, \16786 );
nor \g447185/U$1 ( \27280 , \27278 , \27279 );
nand \g444541/U$1 ( \27281 , \27271 , \27274 , \27277 , \27280 );
and \g453863/U$2 ( \27282 , \16371 , RIfcb5640_7086);
and \g453863/U$3 ( \27283 , RIfca4408_6891, \16427 );
nor \g453863/U$1 ( \27284 , \27282 , \27283 );
and \g446439/U$2 ( \27285 , RIfc7ff40_6478, \16448 );
and \g446439/U$3 ( \27286 , RIded4018_876, \16361 );
and \g449443/U$2 ( \27287 , RIfc6b900_6246, \16321 );
and \g449443/U$3 ( \27288 , \16326 , RIfc69b78_6225);
and \g449443/U$4 ( \27289 , RIded8500_925, \16398 );
nor \g449443/U$1 ( \27290 , \27287 , \27288 , \27289 );
and \g455043/U$2 ( \27291 , \16317 , RIdee3d38_1056);
and \g455043/U$3 ( \27292 , RIdee5ac0_1077, \16325 );
nor \g455043/U$1 ( \27293 , \27291 , \27292 );
not \g450463/U$3 ( \27294 , \27293 );
not \g450463/U$4 ( \27295 , \16330 );
and \g450463/U$2 ( \27296 , \27294 , \27295 );
and \g450463/U$5 ( \27297 , \16341 , RIdeda990_951);
nor \g450463/U$1 ( \27298 , \27296 , \27297 );
and \g453866/U$2 ( \27299 , \16377 , RIfced770_7724);
and \g453866/U$3 ( \27300 , RIfc4d270_5900, \16313 );
nor \g453866/U$1 ( \27301 , \27299 , \27300 );
and \g453867/U$2 ( \27302 , \16334 , RIdedfb20_1009);
and \g453867/U$3 ( \27303 , RIdee1a10_1031, \16380 );
nor \g453867/U$1 ( \27304 , \27302 , \27303 );
nand \g447431/U$1 ( \27305 , \27290 , \27298 , \27301 , \27304 );
nor \g446439/U$1 ( \27306 , \27285 , \27286 , \27305 );
and \g453865/U$2 ( \27307 , \16364 , RIded61d8_900);
and \g453865/U$3 ( \27308 , RIee21700_4839, \16368 );
nor \g453865/U$1 ( \27309 , \27307 , \27308 );
nand \g445689/U$1 ( \27310 , \27284 , \27306 , \27309 );
and \g444925/U$2 ( \27311 , \27310 , \16477 );
and \g449441/U$2 ( \27312 , RIdf20bc0_1749, \16398 );
and \g449441/U$3 ( \27313 , \16341 , RIfcaad80_6966);
and \g449441/U$4 ( \27314 , RIdf29428_1846, \16344 );
nor \g449441/U$1 ( \27315 , \27312 , \27313 , \27314 );
and \g455060/U$2 ( \27316 , \16317 , RIfcdcda8_7535);
and \g455060/U$3 ( \27317 , RIfc5e1d8_6093, \16325 );
nor \g455060/U$1 ( \27318 , \27316 , \27317 );
not \g450461/U$3 ( \27319 , \27318 );
not \g450461/U$4 ( \27320 , \16351 );
and \g450461/U$2 ( \27321 , \27319 , \27320 );
and \g450461/U$5 ( \27322 , \16356 , RIdf2b318_1868);
nor \g450461/U$1 ( \27323 , \27321 , \27322 );
and \g453861/U$2 ( \27324 , \16361 , RIdf1a518_1676);
and \g453861/U$3 ( \27325 , RIfc61b80_6134, \16364 );
nor \g453861/U$1 ( \27326 , \27324 , \27325 );
and \g453860/U$2 ( \27327 , \16368 , RIfc691a0_6218);
and \g453860/U$3 ( \27328 , RIfcac400_6982, \16371 );
nor \g453860/U$1 ( \27329 , \27327 , \27328 );
nand \g447970/U$1 ( \27330 , \27315 , \27323 , \27326 , \27329 );
and \g444925/U$3 ( \27331 , \16481 , \27330 );
nor \g444925/U$1 ( \27332 , \27311 , \27331 );
and \g447179/U$2 ( \27333 , \16505 , RIfca1b40_6862);
and \g447179/U$3 ( \27334 , RIfcb1860_7042, \16507 );
nor \g447179/U$1 ( \27335 , \27333 , \27334 );
and \g447182/U$2 ( \27336 , \16511 , RIfe9af08_8107);
and \g447182/U$3 ( \27337 , RIdf27100_1821, \16514 );
nor \g447182/U$1 ( \27338 , \27336 , \27337 );
and \g447180/U$2 ( \27339 , \16518 , RIfe9ada0_8106);
and \g447180/U$3 ( \27340 , RIfc5c018_6069, \16521 );
nor \g447180/U$1 ( \27341 , \27339 , \27340 );
nand \g444663/U$1 ( \27342 , \27332 , \27335 , \27338 , \27341 );
and \g446436/U$2 ( \27343 , RIe163bf0_2512, \16321 );
and \g446436/U$3 ( \27344 , RIee381d0_5097, \16313 );
and \g449436/U$2 ( \27345 , RIe152df0_2320, \16427 );
and \g449436/U$3 ( \27346 , \16448 , RIfc3f968_5749);
and \g449436/U$4 ( \27347 , RIe15e1f0_2448, \16485 );
nor \g449436/U$1 ( \27348 , \27345 , \27346 , \27347 );
and \g455380/U$2 ( \27349 , \16317 , RIe14d3f0_2256);
and \g455380/U$3 ( \27350 , RIfc84b30_6532, \16325 );
nor \g455380/U$1 ( \27351 , \27349 , \27350 );
not \g455379/U$1 ( \27352 , \27351 );
and \g450458/U$2 ( \27353 , \27352 , \16336 );
and \g450458/U$3 ( \27354 , RIfcdfaa8_7567, \16356 );
nor \g450458/U$1 ( \27355 , \27353 , \27354 );
and \g453851/U$2 ( \27356 , \16361 , RIe1479f0_2192);
and \g453851/U$3 ( \27357 , RIe14a6f0_2224, \16364 );
nor \g453851/U$1 ( \27358 , \27356 , \27357 );
and \g453850/U$2 ( \27359 , \16368 , RIe1500f0_2288);
and \g453850/U$3 ( \27360 , RIfcd5080_7446, \16371 );
nor \g453850/U$1 ( \27361 , \27359 , \27360 );
nand \g448122/U$1 ( \27362 , \27348 , \27355 , \27358 , \27361 );
nor \g446436/U$1 ( \27363 , \27343 , \27344 , \27362 );
and \g453849/U$2 ( \27364 , \16377 , RIe160ef0_2480);
and \g453849/U$3 ( \27365 , RIe1587f0_2384, \16380 );
nor \g453849/U$1 ( \27366 , \27364 , \27365 );
and \g453848/U$2 ( \27367 , \16334 , RIe155af0_2352);
and \g453848/U$3 ( \27368 , RIe1668f0_2544, \16328 );
nor \g453848/U$1 ( \27369 , \27367 , \27368 );
and \g445457/U$2 ( \27370 , \27363 , \27366 , \27369 );
nor \g445457/U$1 ( \27371 , \27370 , \16389 );
and \g446437/U$2 ( \27372 , RIfc57590_6016, \16448 );
and \g446437/U$3 ( \27373 , RIfe9b070_8108, \16361 );
and \g449439/U$2 ( \27374 , RIfc92f00_6694, \16319 );
and \g449439/U$3 ( \27375 , \16328 , RIfcea098_7685);
and \g449439/U$4 ( \27376 , RIdf34558_1972, \16398 );
nor \g449439/U$1 ( \27377 , \27374 , \27375 , \27376 );
and \g455381/U$2 ( \27378 , \16317 , RIe13fe30_2104);
and \g455381/U$3 ( \27379 , RIe142158_2129, \16325 );
nor \g455381/U$1 ( \27380 , \27378 , \27379 );
not \g450460/U$3 ( \27381 , \27380 );
not \g450460/U$4 ( \27382 , \16330 );
and \g450460/U$2 ( \27383 , \27381 , \27382 );
and \g450460/U$5 ( \27384 , \16341 , RIdf36b50_1999);
nor \g450460/U$1 ( \27385 , \27383 , \27384 );
and \g453857/U$2 ( \27386 , \16377 , RIfcdcc40_7534);
and \g453857/U$3 ( \27387 , RIfc54890_5984, \16313 );
nor \g453857/U$1 ( \27388 , \27386 , \27387 );
and \g453858/U$2 ( \27389 , \16334 , RIdf3b8a8_2054);
and \g453858/U$3 ( \27390 , RIdf3dd38_2080, \16380 );
nor \g453858/U$1 ( \27391 , \27389 , \27390 );
nand \g447430/U$1 ( \27392 , \27377 , \27385 , \27388 , \27391 );
nor \g446437/U$1 ( \27393 , \27372 , \27373 , \27392 );
and \g453856/U$2 ( \27394 , \16364 , RIdf32398_1948);
and \g453856/U$3 ( \27395 , RIee2e180_4983, \16368 );
nor \g453856/U$1 ( \27396 , \27394 , \27395 );
and \g453855/U$2 ( \27397 , \16371 , RIfcd0490_7392);
and \g453855/U$3 ( \27398 , RIee30340_5007, \16427 );
nor \g453855/U$1 ( \27399 , \27397 , \27398 );
and \g445458/U$2 ( \27400 , \27393 , \27396 , \27399 );
nor \g445458/U$1 ( \27401 , \27400 , \16393 );
or \g444346/U$1 ( \27402 , \27281 , \27342 , \27371 , \27401 );
and \g446433/U$2 ( \27403 , RIdec68f0_723, \16328 );
and \g446433/U$3 ( \27404 , RIdeb87f0_563, \16334 );
and \g449432/U$2 ( \27405 , RIdead3f0_435, \16398 );
and \g449432/U$3 ( \27406 , \16341 , RIfc5ff60_6114);
and \g449432/U$4 ( \27407 , RIdebe1f0_627, \16485 );
nor \g449432/U$1 ( \27408 , \27405 , \27406 , \27407 );
and \g455070/U$2 ( \27409 , \16317 , RIdeb2df0_499);
and \g455070/U$3 ( \27410 , RIfc9b8d0_6792, \16325 );
nor \g455070/U$1 ( \27411 , \27409 , \27410 );
not \g450453/U$3 ( \27412 , \27411 );
not \g450453/U$4 ( \27413 , \16351 );
and \g450453/U$2 ( \27414 , \27412 , \27413 );
and \g450453/U$5 ( \27415 , \16354 , RIfc7ce08_6443);
nor \g450453/U$1 ( \27416 , \27414 , \27415 );
and \g453836/U$2 ( \27417 , \16361 , RIdea0358_371);
and \g453836/U$3 ( \27418 , RIdea6c58_403, \16364 );
nor \g453836/U$1 ( \27419 , \27417 , \27418 );
and \g453835/U$2 ( \27420 , \16368 , RIdeb00f0_467);
and \g453835/U$3 ( \27421 , RIfcc6710_7280, \16371 );
nor \g453835/U$1 ( \27422 , \27420 , \27421 );
nand \g447967/U$1 ( \27423 , \27408 , \27416 , \27419 , \27422 );
nor \g446433/U$1 ( \27424 , \27403 , \27404 , \27423 );
and \g453834/U$2 ( \27425 , \16377 , RIdec0ef0_659);
and \g453834/U$3 ( \27426 , RIdebb4f0_595, \16380 );
nor \g453834/U$1 ( \27427 , \27425 , \27426 );
and \g453832/U$2 ( \27428 , \16313 , RIee208f0_4829);
and \g453832/U$3 ( \27429 , RIdec3bf0_691, \16321 );
nor \g453832/U$1 ( \27430 , \27428 , \27429 );
and \g445454/U$2 ( \27431 , \27424 , \27427 , \27430 );
nor \g445454/U$1 ( \27432 , \27431 , \16618 );
and \g446434/U$2 ( \27433 , RIfcb2238_7049, \16427 );
and \g446434/U$3 ( \27434 , RIfcdb020_7514, \16368 );
and \g449434/U$2 ( \27435 , RIfe9b1d8_8109, \16485 );
and \g449434/U$3 ( \27436 , \16354 , RIde934a0_308);
and \g449434/U$4 ( \27437 , RIe16c9f8_2613, \16398 );
nor \g449434/U$1 ( \27438 , \27435 , \27436 , \27437 );
and \g455066/U$2 ( \27439 , \16317 , RIee1c6d8_4782);
and \g455066/U$3 ( \27440 , RIfce5070_7628, \16325 );
nor \g455066/U$1 ( \27441 , \27439 , \27440 );
not \g450456/U$3 ( \27442 , \27441 );
not \g450456/U$4 ( \27443 , \16311 );
and \g450456/U$2 ( \27444 , \27442 , \27443 );
and \g450456/U$5 ( \27445 , \16341 , RIfc511b8_5945);
nor \g450456/U$1 ( \27446 , \27444 , \27445 );
and \g453843/U$2 ( \27447 , \16377 , RIee1b058_4766);
and \g453843/U$3 ( \27448 , RIfce70c8_7651, \16313 );
nor \g453843/U$1 ( \27449 , \27447 , \27448 );
and \g453844/U$2 ( \27450 , \16334 , RIfe9b340_8110);
and \g453844/U$3 ( \27451 , RIde8b7f0_270, \16380 );
nor \g453844/U$1 ( \27452 , \27450 , \27451 );
nand \g447429/U$1 ( \27453 , \27438 , \27446 , \27449 , \27452 );
nor \g446434/U$1 ( \27454 , \27433 , \27434 , \27453 );
and \g453841/U$2 ( \27455 , \16361 , RIe168ee8_2571);
and \g453841/U$3 ( \27456 , RIfc6b798_6245, \16448 );
nor \g453841/U$1 ( \27457 , \27455 , \27456 );
and \g453840/U$2 ( \27458 , \16364 , RIfcb27d8_7053);
and \g453840/U$3 ( \27459 , RIfcd3a00_7430, \16371 );
nor \g453840/U$1 ( \27460 , \27458 , \27459 );
and \g445455/U$2 ( \27461 , \27454 , \27457 , \27460 );
nor \g445455/U$1 ( \27462 , \27461 , \16649 );
or \g444284/U$1 ( \27463 , \27402 , \27432 , \27462 );
_DC \g4b10/U$1 ( \27464 , \27463 , \16652 );
and \g453917/U$2 ( \27465 , \8531 , RIfc780b0_6388);
and \g453917/U$3 ( \27466 , RIfc9fc50_6840, \8414 );
nor \g453917/U$1 ( \27467 , \27465 , \27466 );
and \g446451/U$2 ( \27468 , RIf13f820_5182, \8409 );
and \g446451/U$3 ( \27469 , RIfce5340_7630, \8378 );
and \g449456/U$2 ( \27470 , RIfe9a260_8098, \8373 );
and \g449456/U$3 ( \27471 , \8383 , RIf1415a8_5203);
and \g449456/U$4 ( \27472 , RIfc576f8_6017, \8486 );
nor \g449456/U$1 ( \27473 , \27470 , \27471 , \27472 );
and \g453920/U$2 ( \27474 , \8335 , RIfc7e758_6461);
and \g453920/U$3 ( \27475 , RIfc7adb0_6420, \8340 );
nor \g453920/U$1 ( \27476 , \27474 , \27475 );
and \g453919/U$2 ( \27477 , \8404 , RIfe9a0f8_8097);
and \g453919/U$3 ( \27478 , RIfe9a3c8_8099, \8351 );
nor \g453919/U$1 ( \27479 , \27477 , \27478 );
and \g454654/U$2 ( \27480 , \8313 , RIfcb2d78_7057);
and \g454654/U$3 ( \27481 , RIfc7c2c8_6435, \8323 );
nor \g454654/U$1 ( \27482 , \27480 , \27481 );
not \g454653/U$1 ( \27483 , \27482 );
and \g450477/U$2 ( \27484 , \27483 , \8316 );
and \g450477/U$3 ( \27485 , RIfc5cb58_6077, \8359 );
nor \g450477/U$1 ( \27486 , \27484 , \27485 );
nand \g448244/U$1 ( \27487 , \27473 , \27476 , \27479 , \27486 );
nor \g446451/U$1 ( \27488 , \27468 , \27469 , \27487 );
and \g453918/U$2 ( \27489 , \8356 , RIe1749f0_2704);
and \g453918/U$3 ( \27490 , RIfcb9150_7128, \8417 );
nor \g453918/U$1 ( \27491 , \27489 , \27490 );
nand \g445692/U$1 ( \27492 , \27467 , \27488 , \27491 );
and \g444748/U$2 ( \27493 , \27492 , \9700 );
and \g449453/U$2 ( \27494 , RIfe9a698_8101, \8373 );
and \g449453/U$3 ( \27495 , \8330 , RIe19be88_3151);
and \g449453/U$4 ( \27496 , RIe188388_2927, \8488 );
nor \g449453/U$1 ( \27497 , \27494 , \27495 , \27496 );
and \g453915/U$2 ( \27498 , \8335 , RIe17cf88_2799);
and \g453915/U$3 ( \27499 , RIfc8d938_6633, \8340 );
nor \g453915/U$1 ( \27500 , \27498 , \27499 );
and \g453914/U$2 ( \27501 , \8404 , RIe199188_3119);
and \g453914/U$3 ( \27502 , RIe19eb88_3183, \8351 );
nor \g453914/U$1 ( \27503 , \27501 , \27502 );
and \g454671/U$2 ( \27504 , \8313 , RIe17fc88_2831);
and \g454671/U$3 ( \27505 , RIe182988_2863, \8323 );
nor \g454671/U$1 ( \27506 , \27504 , \27505 );
not \g454670/U$1 ( \27507 , \27506 );
and \g450474/U$2 ( \27508 , \27507 , \8316 );
and \g450474/U$3 ( \27509 , RIe18b088_2959, \8359 );
nor \g450474/U$1 ( \27510 , \27508 , \27509 );
nand \g448243/U$1 ( \27511 , \27497 , \27500 , \27503 , \27510 );
and \g444748/U$3 ( \27512 , \9702 , \27511 );
nor \g444748/U$1 ( \27513 , \27493 , \27512 );
and \g447189/U$2 ( \27514 , \11700 , RIe196488_3087);
and \g447189/U$3 ( \27515 , RIfe9a530_8100, \11702 );
nor \g447189/U$1 ( \27516 , \27514 , \27515 );
and \g447190/U$2 ( \27517 , \9230 , RIe185688_2895);
and \g447190/U$3 ( \27518 , RIfe9a800_8102, \9232 );
nor \g447190/U$1 ( \27519 , \27517 , \27518 );
and \g447191/U$2 ( \27520 , \9170 , RIe190a88_3023);
and \g447191/U$3 ( \27521 , RIe193788_3055, \9172 );
nor \g447191/U$1 ( \27522 , \27520 , \27521 );
nand \g444542/U$1 ( \27523 , \27513 , \27516 , \27519 , \27522 );
and \g453926/U$2 ( \27524 , \8523 , RIfccee10_7376);
and \g453926/U$3 ( \27525 , RIfca8e90_6944, \8412 );
nor \g453926/U$1 ( \27526 , \27524 , \27525 );
and \g446454/U$2 ( \27527 , RIfc6d688_6267, \8409 );
and \g446454/U$3 ( \27528 , RIe1f6860_4182, \8378 );
and \g449459/U$2 ( \27529 , RIfcae458_7005, \8317 );
and \g449459/U$3 ( \27530 , \8326 , RIfcaecc8_7011);
and \g449459/U$4 ( \27531 , RIfcaee30_7012, \8488 );
nor \g449459/U$1 ( \27532 , \27529 , \27530 , \27531 );
and \g453931/U$2 ( \27533 , \8335 , RIfeab1c8_8263);
and \g453931/U$3 ( \27534 , RIfc63ea8_6159, \8340 );
nor \g453931/U$1 ( \27535 , \27533 , \27534 );
and \g453930/U$2 ( \27536 , \8404 , RIfec3b88_8347);
and \g453930/U$3 ( \27537 , RIfc71cd8_6317, \8351 );
nor \g453930/U$1 ( \27538 , \27536 , \27537 );
and \g454554/U$2 ( \27539 , \8313 , RIfcaa3a8_6959);
and \g454554/U$3 ( \27540 , RIfccb198_7333, \8323 );
nor \g454554/U$1 ( \27541 , \27539 , \27540 );
not \g450479/U$3 ( \27542 , \27541 );
not \g450479/U$4 ( \27543 , \8328 );
and \g450479/U$2 ( \27544 , \27542 , \27543 );
and \g450479/U$5 ( \27545 , \8359 , RIfc64e20_6170);
nor \g450479/U$1 ( \27546 , \27544 , \27545 );
nand \g447981/U$1 ( \27547 , \27532 , \27535 , \27538 , \27546 );
nor \g446454/U$1 ( \27548 , \27527 , \27528 , \27547 );
and \g453927/U$2 ( \27549 , \8356 , RIe1f4538_4157);
and \g453927/U$3 ( \27550 , RIfc4c730_5892, \8417 );
nor \g453927/U$1 ( \27551 , \27549 , \27550 );
nand \g445693/U$1 ( \27552 , \27526 , \27548 , \27551 );
and \g444845/U$2 ( \27553 , \27552 , \8752 );
and \g449458/U$2 ( \27554 , RIe227be0_4742, \8414 );
and \g449458/U$3 ( \27555 , \8409 , RIe17a288_2767);
and \g449458/U$4 ( \27556 , RIe1a7288_3279, \8383 );
nor \g449458/U$1 ( \27557 , \27554 , \27555 , \27556 );
and \g453924/U$2 ( \27558 , \8356 , RIe1f1f40_4130);
and \g453924/U$3 ( \27559 , RIe205fe0_4358, \8359 );
nor \g453924/U$1 ( \27560 , \27558 , \27559 );
and \g454621/U$2 ( \27561 , \8313 , RIe1f93f8_4213);
and \g454621/U$3 ( \27562 , RIe200040_4290, \8323 );
nor \g454621/U$1 ( \27563 , \27561 , \27562 );
not \g450478/U$3 ( \27564 , \27563 );
not \g450478/U$4 ( \27565 , \8347 );
and \g450478/U$2 ( \27566 , \27564 , \27565 );
and \g450478/U$5 ( \27567 , \8351 , RIe1a9f88_3311);
nor \g450478/U$1 ( \27568 , \27566 , \27567 );
and \g453923/U$2 ( \27569 , \8378 , RIe21c7e0_4614);
and \g453923/U$3 ( \27570 , RIe18dd88_2991, \8417 );
nor \g453923/U$1 ( \27571 , \27569 , \27570 );
nand \g447980/U$1 ( \27572 , \27557 , \27560 , \27568 , \27571 );
and \g444845/U$3 ( \27573 , \9010 , \27572 );
nor \g444845/U$1 ( \27574 , \27553 , \27573 );
and \g447193/U$2 ( \27575 , \9041 , RIe1a1888_3215);
and \g447193/U$3 ( \27576 , RIe1a4588_3247, \9043 );
nor \g447193/U$1 ( \27577 , \27575 , \27576 );
and \g447194/U$2 ( \27578 , \13239 , RIe1bcf48_3527);
and \g447194/U$3 ( \27579 , RIe1d6448_3815, \13241 );
nor \g447194/U$1 ( \27580 , \27578 , \27579 );
and \g447195/U$2 ( \27581 , \13244 , RIe1723f8_2677);
and \g447195/U$3 ( \27582 , RIe1afdc0_3378, \13246 );
nor \g447195/U$1 ( \27583 , \27581 , \27582 );
nand \g444664/U$1 ( \27584 , \27574 , \27577 , \27580 , \27583 );
and \g446446/U$2 ( \27585 , RIe1e7248_4007, \8371 );
and \g446446/U$3 ( \27586 , RIe1c2948_3591, \8317 );
and \g449451/U$2 ( \27587 , RIe1cdd48_3719, \8531 );
and \g449451/U$3 ( \27588 , \8486 , RIe1d0a48_3751);
and \g449451/U$4 ( \27589 , RIe1e9f48_4039, \8383 );
nor \g449451/U$1 ( \27590 , \27587 , \27588 , \27589 );
and \g453903/U$2 ( \27591 , \8356 , RIe1cb048_3687);
and \g453903/U$3 ( \27592 , RIe1d3748_3783, \8359 );
nor \g453903/U$1 ( \27593 , \27591 , \27592 );
and \g454708/U$2 ( \27594 , \8313 , RIe1dbe48_3879);
and \g454708/U$3 ( \27595 , RIe1deb48_3911, \8323 );
nor \g454708/U$1 ( \27596 , \27594 , \27595 );
not \g450471/U$3 ( \27597 , \27596 );
not \g450471/U$4 ( \27598 , \8376 );
and \g450471/U$2 ( \27599 , \27597 , \27598 );
and \g450471/U$5 ( \27600 , \8351 , RIe1ecc48_4071);
nor \g450471/U$1 ( \27601 , \27599 , \27600 );
and \g453902/U$2 ( \27602 , \8378 , RIe1d9148_3847);
and \g453902/U$3 ( \27603 , RIe1e1848_3943, \8417 );
nor \g453902/U$1 ( \27604 , \27602 , \27603 );
nand \g447976/U$1 ( \27605 , \27590 , \27593 , \27601 , \27604 );
nor \g446446/U$1 ( \27606 , \27585 , \27586 , \27605 );
and \g453900/U$2 ( \27607 , \8335 , RIe1bfc48_3559);
and \g453900/U$3 ( \27608 , RIe1c8348_3655, \8340 );
nor \g453900/U$1 ( \27609 , \27607 , \27608 );
and \g453899/U$2 ( \27610 , \8326 , RIe1c5648_3623);
and \g453899/U$3 ( \27611 , RIe1e4548_3975, \8404 );
nor \g453899/U$1 ( \27612 , \27610 , \27611 );
and \g445465/U$2 ( \27613 , \27606 , \27609 , \27612 );
nor \g445465/U$1 ( \27614 , \27613 , \8477 );
and \g446449/U$2 ( \27615 , RIfcc2228_7231, \8409 );
and \g446449/U$3 ( \27616 , RIe1b4848_3431, \8378 );
and \g449452/U$2 ( \27617 , RIe1ad390_3348, \8319 );
and \g449452/U$3 ( \27618 , \8324 , RIfc4b4e8_5879);
and \g449452/U$4 ( \27619 , RIfc55970_5996, \8488 );
nor \g449452/U$1 ( \27620 , \27617 , \27618 , \27619 );
and \g453909/U$2 ( \27621 , \8335 , RIe1abba8_3331);
and \g453909/U$3 ( \27622 , RIfcb7698_7109, \8340 );
nor \g453909/U$1 ( \27623 , \27621 , \27622 );
and \g453908/U$2 ( \27624 , \8404 , RIe1b8358_3473);
and \g453908/U$3 ( \27625 , RIfcc70e8_7287, \8351 );
nor \g453908/U$1 ( \27626 , \27624 , \27625 );
and \g455391/U$2 ( \27627 , \8313 , RIe1ba518_3497);
and \g455391/U$3 ( \27628 , RIfca7ae0_6930, \8323 );
nor \g455391/U$1 ( \27629 , \27627 , \27628 );
not \g450473/U$3 ( \27630 , \27629 );
not \g450473/U$4 ( \27631 , \8328 );
and \g450473/U$2 ( \27632 , \27630 , \27631 );
and \g450473/U$5 ( \27633 , \8359 , RIfc82f10_6512);
nor \g450473/U$1 ( \27634 , \27632 , \27633 );
nand \g447977/U$1 ( \27635 , \27620 , \27623 , \27626 , \27634 );
nor \g446449/U$1 ( \27636 , \27615 , \27616 , \27635 );
and \g453906/U$2 ( \27637 , \8356 , RIe1b1cb0_3400);
and \g453906/U$3 ( \27638 , RIfc598b8_6041, \8417 );
nor \g453906/U$1 ( \27639 , \27637 , \27638 );
and \g453904/U$2 ( \27640 , \8531 , RIe1b3498_3417);
and \g453904/U$3 ( \27641 , RIe1b6198_3449, \8414 );
nor \g453904/U$1 ( \27642 , \27640 , \27641 );
and \g445466/U$2 ( \27643 , \27636 , \27639 , \27642 );
nor \g445466/U$1 ( \27644 , \27643 , \8481 );
or \g444337/U$1 ( \27645 , \27523 , \27584 , \27614 , \27644 );
and \g446443/U$2 ( \27646 , RIf16c3e8_5691, \8373 );
and \g446443/U$3 ( \27647 , RIe20b9e0_4422, \8319 );
and \g449448/U$2 ( \27648 , RIf169c88_5663, \8523 );
and \g449448/U$3 ( \27649 , \8488 , RIe2140e0_4518);
and \g449448/U$4 ( \27650 , RIe224ee0_4710, \8383 );
nor \g449448/U$1 ( \27651 , \27648 , \27649 , \27650 );
and \g453888/U$2 ( \27652 , \8356 , RIe2113e0_4486);
and \g453888/U$3 ( \27653 , RIfc880a0_6570, \8359 );
nor \g453888/U$1 ( \27654 , \27652 , \27653 );
and \g455389/U$2 ( \27655 , \8313 , RIe219ae0_4582);
and \g455389/U$3 ( \27656 , RIe21f4e0_4646, \8323 );
nor \g455389/U$1 ( \27657 , \27655 , \27656 );
not \g450468/U$3 ( \27658 , \27657 );
not \g450468/U$4 ( \27659 , \8376 );
and \g450468/U$2 ( \27660 , \27658 , \27659 );
and \g450468/U$5 ( \27661 , \8351 , RIfe9aad0_8104);
nor \g450468/U$1 ( \27662 , \27660 , \27661 );
and \g453887/U$2 ( \27663 , \8378 , RIe216de0_4550);
and \g453887/U$3 ( \27664 , RIfcd3898_7429, \8417 );
nor \g453887/U$1 ( \27665 , \27663 , \27664 );
nand \g447974/U$1 ( \27666 , \27651 , \27654 , \27662 , \27665 );
nor \g446443/U$1 ( \27667 , \27646 , \27647 , \27666 );
and \g453885/U$2 ( \27668 , \8335 , RIe208ce0_4390);
and \g453885/U$3 ( \27669 , RIf168338_5645, \8340 );
nor \g453885/U$1 ( \27670 , \27668 , \27669 );
and \g453883/U$2 ( \27671 , \8326 , RIe20e6e0_4454);
and \g453883/U$3 ( \27672 , RIe2221e0_4678, \8404 );
nor \g453883/U$1 ( \27673 , \27671 , \27672 );
and \g445462/U$2 ( \27674 , \27667 , \27670 , \27673 );
nor \g445462/U$1 ( \27675 , \27674 , \8368 );
and \g446445/U$2 ( \27676 , RIfca8d28_6943, \8340 );
and \g446445/U$3 ( \27677 , RIe201af8_4309, \8404 );
and \g449449/U$2 ( \27678 , RIfce81a8_7663, \8412 );
and \g449449/U$3 ( \27679 , \8407 , RIfc85c10_6544);
and \g449449/U$4 ( \27680 , RIfc9c6e0_6802, \8383 );
nor \g449449/U$1 ( \27681 , \27678 , \27679 , \27680 );
and \g453895/U$2 ( \27682 , \8356 , RIfe9ac38_8105);
and \g453895/U$3 ( \27683 , RIf160e80_5562, \8359 );
nor \g453895/U$1 ( \27684 , \27682 , \27683 );
and \g455390/U$2 ( \27685 , \8313 , RIfe9a968_8103);
and \g455390/U$3 ( \27686 , RIf15ef90_5540, \8323 );
nor \g455390/U$1 ( \27687 , \27685 , \27686 );
not \g450469/U$3 ( \27688 , \27687 );
not \g450469/U$4 ( \27689 , \8347 );
and \g450469/U$2 ( \27690 , \27688 , \27689 );
and \g450469/U$5 ( \27691 , \8351 , RIfce4c38_7625);
nor \g450469/U$1 ( \27692 , \27690 , \27691 );
and \g453894/U$2 ( \27693 , \8378 , RIfce9c60_7682);
and \g453894/U$3 ( \27694 , RIfc500d8_5933, \8417 );
nor \g453894/U$1 ( \27695 , \27693 , \27694 );
nand \g447975/U$1 ( \27696 , \27681 , \27684 , \27692 , \27695 );
nor \g446445/U$1 ( \27697 , \27676 , \27677 , \27696 );
and \g453891/U$2 ( \27698 , \8335 , RIfc6a988_6235);
and \g453891/U$3 ( \27699 , RIe2035b0_4328, \8371 );
nor \g453891/U$1 ( \27700 , \27698 , \27699 );
and \g453892/U$2 ( \27701 , \8319 , RIfcedba8_7727);
and \g453892/U$3 ( \27702 , RIf15be58_5505, \8326 );
nor \g453892/U$1 ( \27703 , \27701 , \27702 );
and \g445463/U$2 ( \27704 , \27697 , \27700 , \27703 );
nor \g445463/U$1 ( \27705 , \27704 , \8422 );
or \g444251/U$1 ( \27706 , \27645 , \27675 , \27705 );
_DC \g4b94/U$1 ( \27707 , \27706 , \8654 );
and \g453960/U$2 ( \27708 , \16371 , RIfc65960_6178);
and \g453960/U$3 ( \27709 , RIfc42c80_5782, \16427 );
nor \g453960/U$1 ( \27710 , \27708 , \27709 );
and \g446461/U$2 ( \27711 , RIde834b0_230, \16448 );
and \g446461/U$3 ( \27712 , RIe169050_2572, \16361 );
and \g449468/U$2 ( \27713 , RIfc83780_6518, \16321 );
and \g449468/U$3 ( \27714 , \16326 , RIfc81458_6493);
and \g449468/U$4 ( \27715 , RIe16cb60_2614, \16398 );
nor \g449468/U$1 ( \27716 , \27713 , \27714 , \27715 );
and \g454267/U$2 ( \27717 , \16317 , RIde8f990_290);
and \g454267/U$3 ( \27718 , RIde937e8_309, \16325 );
nor \g454267/U$1 ( \27719 , \27717 , \27718 );
not \g450491/U$3 ( \27720 , \27719 );
not \g450491/U$4 ( \27721 , \16330 );
and \g450491/U$2 ( \27722 , \27720 , \27721 );
and \g450491/U$5 ( \27723 , \16341 , RIee392b0_5109);
nor \g450491/U$1 ( \27724 , \27722 , \27723 );
and \g453965/U$2 ( \27725 , \16377 , RIfcd3e38_7433);
and \g453965/U$3 ( \27726 , RIfc4e620_5914, \16313 );
nor \g453965/U$1 ( \27727 , \27725 , \27726 );
and \g453966/U$2 ( \27728 , \16334 , RIde87650_250);
and \g453966/U$3 ( \27729 , RIde8bb38_271, \16380 );
nor \g453966/U$1 ( \27730 , \27728 , \27729 );
nand \g447440/U$1 ( \27731 , \27716 , \27724 , \27727 , \27730 );
nor \g446461/U$1 ( \27732 , \27711 , \27712 , \27731 );
and \g453962/U$2 ( \27733 , \16364 , RIe16a6d0_2588);
and \g453962/U$3 ( \27734 , RIfc6c710_6256, \16368 );
nor \g453962/U$1 ( \27735 , \27733 , \27734 );
nand \g445695/U$1 ( \27736 , \27710 , \27732 , \27735 );
and \g444809/U$2 ( \27737 , \27736 , \17998 );
and \g449467/U$2 ( \27738 , RIe14d558_2257, \16337 );
and \g449467/U$3 ( \27739 , \16339 , RIfcb9b28_7135);
and \g449467/U$4 ( \27740 , RIe15e358_2449, \16344 );
nor \g449467/U$1 ( \27741 , \27738 , \27739 , \27740 );
and \g455032/U$2 ( \27742 , \16317 , RIe152f58_2321);
and \g455032/U$3 ( \27743 , RIfe9ba48_8115, \16325 );
nor \g455032/U$1 ( \27744 , \27742 , \27743 );
not \g450490/U$3 ( \27745 , \27744 );
not \g450490/U$4 ( \27746 , \16351 );
and \g450490/U$2 ( \27747 , \27745 , \27746 );
and \g450490/U$5 ( \27748 , \16356 , RIfcd54b8_7449);
nor \g450490/U$1 ( \27749 , \27747 , \27748 );
and \g453959/U$2 ( \27750 , \16361 , RIe147b58_2193);
and \g453959/U$3 ( \27751 , RIe14a858_2225, \16364 );
nor \g453959/U$1 ( \27752 , \27750 , \27751 );
and \g453958/U$2 ( \27753 , \16368 , RIe150258_2289);
and \g453958/U$3 ( \27754 , RIfec4128_8351, \16371 );
nor \g453958/U$1 ( \27755 , \27753 , \27754 );
nand \g447984/U$1 ( \27756 , \27741 , \27749 , \27752 , \27755 );
and \g444809/U$3 ( \27757 , \16390 , \27756 );
nor \g444809/U$1 ( \27758 , \27737 , \27757 );
and \g447201/U$2 ( \27759 , \18020 , RIe163d58_2513);
and \g447201/U$3 ( \27760 , RIe166a58_2545, \18022 );
nor \g447201/U$1 ( \27761 , \27759 , \27760 );
and \g447202/U$2 ( \27762 , \18025 , RIe161058_2481);
and \g447202/U$3 ( \27763 , RIfec3cf0_8348, \18027 );
nor \g447202/U$1 ( \27764 , \27762 , \27763 );
and \g447203/U$2 ( \27765 , \18030 , RIe155c58_2353);
and \g447203/U$3 ( \27766 , RIe158958_2385, \18032 );
nor \g447203/U$1 ( \27767 , \27765 , \27766 );
nand \g444545/U$1 ( \27768 , \27758 , \27761 , \27764 , \27767 );
and \g453973/U$2 ( \27769 , \16371 , RIfce1c68_7591);
and \g453973/U$3 ( \27770 , RIdeb2f58_500, \16427 );
nor \g453973/U$1 ( \27771 , \27769 , \27770 );
and \g446465/U$2 ( \27772 , RIfcb96f0_7132, \16432 );
and \g446465/U$3 ( \27773 , RIdea06a0_372, \16361 );
and \g449473/U$2 ( \27774 , RIdec3d58_692, \16321 );
and \g449473/U$3 ( \27775 , \16328 , RIdec6a58_724);
and \g449473/U$4 ( \27776 , RIdead558_436, \16398 );
nor \g449473/U$1 ( \27777 , \27774 , \27775 , \27776 );
and \g455026/U$2 ( \27778 , \16317 , RIdebe358_628);
and \g455026/U$3 ( \27779 , RIfc59fc0_6046, \16325 );
nor \g455026/U$1 ( \27780 , \27778 , \27779 );
not \g450494/U$3 ( \27781 , \27780 );
not \g450494/U$4 ( \27782 , \16330 );
and \g450494/U$2 ( \27783 , \27781 , \27782 );
and \g450494/U$5 ( \27784 , \16341 , RIfc9b498_6789);
nor \g450494/U$1 ( \27785 , \27783 , \27784 );
and \g453977/U$2 ( \27786 , \16377 , RIdec1058_660);
and \g453977/U$3 ( \27787 , RIfc723e0_6322, \16313 );
nor \g453977/U$1 ( \27788 , \27786 , \27787 );
and \g453978/U$2 ( \27789 , \16334 , RIdeb8958_564);
and \g453978/U$3 ( \27790 , RIdebb658_596, \16380 );
nor \g453978/U$1 ( \27791 , \27789 , \27790 );
nand \g447442/U$1 ( \27792 , \27777 , \27785 , \27788 , \27791 );
nor \g446465/U$1 ( \27793 , \27772 , \27773 , \27792 );
and \g453974/U$2 ( \27794 , \16364 , RIdea6fa0_404);
and \g453974/U$3 ( \27795 , RIdeb0258_468, \16368 );
nor \g453974/U$1 ( \27796 , \27794 , \27795 );
nand \g445696/U$1 ( \27797 , \27771 , \27793 , \27796 );
and \g444736/U$2 ( \27798 , \27797 , \17938 );
and \g449472/U$2 ( \27799 , RIfc553d0_5992, \16321 );
and \g449472/U$3 ( \27800 , \16326 , RIfcdb2f0_7516);
and \g449472/U$4 ( \27801 , RIfec3fc0_8350, \16398 );
nor \g449472/U$1 ( \27802 , \27799 , \27800 , \27801 );
and \g454212/U$2 ( \27803 , \16317 , RIe13ff98_2105);
and \g454212/U$3 ( \27804 , RIe1422c0_2130, \16325 );
nor \g454212/U$1 ( \27805 , \27803 , \27804 );
not \g450493/U$3 ( \27806 , \27805 );
not \g450493/U$4 ( \27807 , \16330 );
and \g450493/U$2 ( \27808 , \27806 , \27807 );
and \g450493/U$5 ( \27809 , \16341 , RIdf36cb8_2000);
nor \g450493/U$1 ( \27810 , \27808 , \27809 );
and \g453970/U$2 ( \27811 , \16377 , RIfcbd908_7179);
and \g453970/U$3 ( \27812 , RIfc9a0e8_6775, \16313 );
nor \g453970/U$1 ( \27813 , \27811 , \27812 );
and \g453971/U$2 ( \27814 , \16334 , RIdf3ba10_2055);
and \g453971/U$3 ( \27815 , RIdf3dea0_2081, \16380 );
nor \g453971/U$1 ( \27816 , \27814 , \27815 );
nand \g447441/U$1 ( \27817 , \27802 , \27810 , \27813 , \27816 );
and \g444736/U$3 ( \27818 , \16394 , \27817 );
nor \g444736/U$1 ( \27819 , \27798 , \27818 );
and \g447209/U$2 ( \27820 , \16419 , RIfec3e58_8349);
and \g447209/U$3 ( \27821 , RIdf32500_1949, \16422 );
nor \g447209/U$1 ( \27822 , \27820 , \27821 );
and \g447207/U$2 ( \27823 , \16429 , RIee304a8_5008);
and \g447207/U$3 ( \27824 , RIfc87128_6559, \16434 );
nor \g447207/U$1 ( \27825 , \27823 , \27824 );
and \g447208/U$2 ( \27826 , \16438 , RIee2e2e8_4984);
and \g447208/U$3 ( \27827 , RIfcc51f8_7265, \16441 );
nor \g447208/U$1 ( \27828 , \27826 , \27827 );
nand \g444546/U$1 ( \27829 , \27819 , \27822 , \27825 , \27828 );
and \g446459/U$2 ( \27830 , RIe144e58_2161, \16448 );
and \g446459/U$3 ( \27831 , RIde7fce8_213, \16361 );
and \g449463/U$2 ( \27832 , RIdecf158_820, \16319 );
and \g449463/U$3 ( \27833 , \16326 , RIded1e58_852);
and \g449463/U$4 ( \27834 , RIdee8928_1110, \16398 );
nor \g449463/U$1 ( \27835 , \27832 , \27833 , \27834 );
and \g454402/U$2 ( \27836 , \16317 , RIde99da0_340);
and \g454402/U$3 ( \27837 , RIdeb5c58_532, \16325 );
nor \g454402/U$1 ( \27838 , \27836 , \27837 );
not \g450484/U$3 ( \27839 , \27838 );
not \g450484/U$4 ( \27840 , \16330 );
and \g450484/U$2 ( \27841 , \27839 , \27840 );
and \g450484/U$5 ( \27842 , \16341 , RIdf01e28_1398);
nor \g450484/U$1 ( \27843 , \27841 , \27842 );
and \g453950/U$2 ( \27844 , \16377 , RIdec9758_756);
and \g453950/U$3 ( \27845 , RIdecc458_788, \16313 );
nor \g453950/U$1 ( \27846 , \27844 , \27845 );
and \g453951/U$2 ( \27847 , \16334 , RIe15b658_2417);
and \g453951/U$3 ( \27848 , RIe16f860_2646, \16380 );
nor \g453951/U$1 ( \27849 , \27847 , \27848 );
nand \g447437/U$1 ( \27850 , \27835 , \27843 , \27846 , \27849 );
nor \g446459/U$1 ( \27851 , \27830 , \27831 , \27850 );
and \g453947/U$2 ( \27852 , \16364 , RIdedd690_983);
and \g453947/U$3 ( \27853 , RIdf1e730_1723, \16368 );
nor \g453947/U$1 ( \27854 , \27852 , \27853 );
and \g453946/U$2 ( \27855 , \16371 , RIdf2deb0_1899);
and \g453946/U$3 ( \27856 , RIdf39850_2031, \16427 );
nor \g453946/U$1 ( \27857 , \27855 , \27856 );
and \g445471/U$2 ( \27858 , \27851 , \27854 , \27857 );
nor \g445471/U$1 ( \27859 , \27858 , \16586 );
and \g446460/U$2 ( \27860 , RIee227e0_4851, \16427 );
and \g446460/U$3 ( \27861 , RIee21868_4840, \16368 );
and \g449465/U$2 ( \27862 , RIdee3ea0_1057, \16485 );
and \g449465/U$3 ( \27863 , \16354 , RIdee5c28_1078);
and \g449465/U$4 ( \27864 , RIded8668_926, \16398 );
nor \g449465/U$1 ( \27865 , \27862 , \27863 , \27864 );
and \g455036/U$2 ( \27866 , \16317 , RIee24c70_4877);
and \g455036/U$3 ( \27867 , RIee25a80_4887, \16325 );
nor \g455036/U$1 ( \27868 , \27866 , \27867 );
not \g450487/U$3 ( \27869 , \27868 );
not \g450487/U$4 ( \27870 , \16311 );
and \g450487/U$2 ( \27871 , \27869 , \27870 );
and \g450487/U$5 ( \27872 , \16341 , RIdedaaf8_952);
nor \g450487/U$1 ( \27873 , \27871 , \27872 );
and \g453956/U$2 ( \27874 , \16377 , RIfccc110_7344);
and \g453956/U$3 ( \27875 , RIfcddd20_7546, \16313 );
nor \g453956/U$1 ( \27876 , \27874 , \27875 );
and \g453957/U$2 ( \27877 , \16334 , RIdedfc88_1010);
and \g453957/U$3 ( \27878 , RIdee1b78_1032, \16380 );
nor \g453957/U$1 ( \27879 , \27877 , \27878 );
nand \g447438/U$1 ( \27880 , \27865 , \27873 , \27876 , \27879 );
nor \g446460/U$1 ( \27881 , \27860 , \27861 , \27880 );
and \g453955/U$2 ( \27882 , \16361 , RIded4180_877);
and \g453955/U$3 ( \27883 , RIfc6a6b8_6233, \16432 );
nor \g453955/U$1 ( \27884 , \27882 , \27883 );
and \g453954/U$2 ( \27885 , \16364 , RIded6340_901);
and \g453954/U$3 ( \27886 , RIfc88be0_6578, \16371 );
nor \g453954/U$1 ( \27887 , \27885 , \27886 );
and \g445472/U$2 ( \27888 , \27881 , \27884 , \27887 );
nor \g445472/U$1 ( \27889 , \27888 , \16909 );
or \g444321/U$1 ( \27890 , \27768 , \27829 , \27859 , \27889 );
and \g446455/U$2 ( \27891 , RIdf18628_1654, \16328 );
and \g446455/U$3 ( \27892 , RIdf04b28_1430, \16334 );
and \g449461/U$2 ( \27893 , RIdef1028_1206, \16398 );
and \g449461/U$3 ( \27894 , \16341 , RIdef3d28_1238);
and \g449461/U$4 ( \27895 , RIdf0a528_1494, \16485 );
nor \g449461/U$1 ( \27896 , \27893 , \27894 , \27895 );
and \g455392/U$2 ( \27897 , \16317 , RIdefc428_1334);
and \g455392/U$3 ( \27898 , RIdeff128_1366, \16325 );
nor \g455392/U$1 ( \27899 , \27897 , \27898 );
not \g450481/U$3 ( \27900 , \27899 );
not \g450481/U$4 ( \27901 , \16351 );
and \g450481/U$2 ( \27902 , \27900 , \27901 );
and \g450481/U$5 ( \27903 , \16356 , RIdf0d228_1526);
nor \g450481/U$1 ( \27904 , \27902 , \27903 );
and \g453936/U$2 ( \27905 , \16361 , RIdeeb628_1142);
and \g453936/U$3 ( \27906 , RIdeee328_1174, \16364 );
nor \g453936/U$1 ( \27907 , \27905 , \27906 );
and \g453935/U$2 ( \27908 , \16368 , RIdef6a28_1270);
and \g453935/U$3 ( \27909 , RIdef9728_1302, \16371 );
nor \g453935/U$1 ( \27910 , \27908 , \27909 );
nand \g447982/U$1 ( \27911 , \27896 , \27904 , \27907 , \27910 );
nor \g446455/U$1 ( \27912 , \27891 , \27892 , \27911 );
and \g453934/U$2 ( \27913 , \16377 , RIdf0ff28_1558);
and \g453934/U$3 ( \27914 , RIdf07828_1462, \16380 );
nor \g453934/U$1 ( \27915 , \27913 , \27914 );
and \g453933/U$2 ( \27916 , \16313 , RIdf12c28_1590);
and \g453933/U$3 ( \27917 , RIdf15928_1622, \16321 );
nor \g453933/U$1 ( \27918 , \27916 , \27917 );
and \g445468/U$2 ( \27919 , \27912 , \27915 , \27918 );
nor \g445468/U$1 ( \27920 , \27919 , \16555 );
and \g446457/U$2 ( \27921 , RIfcb7c38_7113, \16448 );
and \g446457/U$3 ( \27922 , RIdf238c0_1781, \16371 );
and \g449462/U$2 ( \27923 , RIfe9b610_8112, \16485 );
and \g449462/U$3 ( \27924 , \16356 , RIfe9b8e0_8114);
and \g449462/U$4 ( \27925 , RIfeaa3b8_8253, \16398 );
nor \g449462/U$1 ( \27926 , \27923 , \27924 , \27925 );
and \g454460/U$2 ( \27927 , \16317 , RIee2ad78_4946);
and \g454460/U$3 ( \27928 , RIee2c830_4965, \16325 );
nor \g454460/U$1 ( \27929 , \27927 , \27928 );
not \g450482/U$3 ( \27930 , \27929 );
not \g450482/U$4 ( \27931 , \16311 );
and \g450482/U$2 ( \27932 , \27930 , \27931 );
and \g450482/U$5 ( \27933 , \16339 , RIdf22240_1765);
nor \g450482/U$1 ( \27934 , \27932 , \27933 );
and \g453942/U$2 ( \27935 , \16377 , RIee284b0_4917);
and \g453942/U$3 ( \27936 , RIee296f8_4930, \16313 );
nor \g453942/U$1 ( \27937 , \27935 , \27936 );
and \g453943/U$2 ( \27938 , \16334 , RIfe9b4a8_8111);
and \g453943/U$3 ( \27939 , RIfe9b778_8113, \16380 );
nor \g453943/U$1 ( \27940 , \27938 , \27939 );
nand \g447436/U$1 ( \27941 , \27926 , \27934 , \27937 , \27940 );
nor \g446457/U$1 ( \27942 , \27921 , \27922 , \27941 );
and \g453939/U$2 ( \27943 , \16364 , RIdf1bb98_1692);
and \g453939/U$3 ( \27944 , RIfc75ab8_6361, \16368 );
nor \g453939/U$1 ( \27945 , \27943 , \27944 );
and \g453941/U$2 ( \27946 , \16361 , RIdf1a680_1677);
and \g453941/U$3 ( \27947 , RIfc86b88_6555, \16427 );
nor \g453941/U$1 ( \27948 , \27946 , \27947 );
and \g445470/U$2 ( \27949 , \27942 , \27945 , \27948 );
nor \g445470/U$1 ( \27950 , \27949 , \16480 );
or \g444265/U$1 ( \27951 , \27890 , \27920 , \27950 );
_DC \g4c19/U$1 ( \27952 , \27951 , \16652 );
and \g447214/U$2 ( \27953 , \11511 , RIe1fb2e8_4235);
and \g447214/U$3 ( \27954 , RIfcc01d0_7208, \11513 );
nor \g447214/U$1 ( \27955 , \27953 , \27954 );
and \g446470/U$2 ( \27956 , RIfc43bf8_5793, \8326 );
and \g446470/U$3 ( \27957 , RIfca6028_6911, \8340 );
and \g449482/U$2 ( \27958 , RIf150ff8_5381, \8531 );
and \g449482/U$3 ( \27959 , \8488 , RIf152240_5394);
and \g449482/U$4 ( \27960 , RIfe9c2b8_8121, \8383 );
nor \g449482/U$1 ( \27961 , \27958 , \27959 , \27960 );
and \g454009/U$2 ( \27962 , \8356 , RIe1f46a0_4158);
and \g454009/U$3 ( \27963 , RIf153a28_5411, \8359 );
nor \g454009/U$1 ( \27964 , \27962 , \27963 );
and \g455350/U$2 ( \27965 , \8313 , RIf154c70_5424);
and \g455350/U$3 ( \27966 , RIfca3e68_6887, \8323 );
nor \g455350/U$1 ( \27967 , \27965 , \27966 );
not \g450503/U$3 ( \27968 , \27967 );
not \g450503/U$4 ( \27969 , \8376 );
and \g450503/U$2 ( \27970 , \27968 , \27969 );
and \g450503/U$5 ( \27971 , \8351 , RIfec4290_8352);
nor \g450503/U$1 ( \27972 , \27970 , \27971 );
and \g454008/U$2 ( \27973 , \8378 , RIe1f69c8_4183);
and \g454008/U$3 ( \27974 , RIfe9c420_8122, \8417 );
nor \g454008/U$1 ( \27975 , \27973 , \27974 );
nand \g447990/U$1 ( \27976 , \27961 , \27964 , \27972 , \27975 );
nor \g446470/U$1 ( \27977 , \27956 , \27957 , \27976 );
not \g444823/U$3 ( \27978 , \27977 );
not \g444823/U$4 ( \27979 , \8621 );
and \g444823/U$2 ( \27980 , \27978 , \27979 );
and \g446473/U$2 ( \27981 , RIe1dbfb0_3880, \8412 );
and \g446473/U$3 ( \27982 , RIe1e19b0_3944, \8417 );
and \g449483/U$2 ( \27983 , RIe1c2ab0_3592, \8319 );
and \g449483/U$3 ( \27984 , \8326 , RIe1c57b0_3624);
and \g449483/U$4 ( \27985 , RIe1d0bb0_3752, \8488 );
nor \g449483/U$1 ( \27986 , \27983 , \27984 , \27985 );
and \g454017/U$2 ( \27987 , \8335 , RIe1bfdb0_3560);
and \g454017/U$3 ( \27988 , RIe1c84b0_3656, \8340 );
nor \g454017/U$1 ( \27989 , \27987 , \27988 );
and \g454016/U$2 ( \27990 , \8404 , RIe1e46b0_3976);
and \g454016/U$3 ( \27991 , RIe1ecdb0_4072, \8351 );
nor \g454016/U$1 ( \27992 , \27990 , \27991 );
and \g454493/U$2 ( \27993 , \8313 , RIe1e73b0_4008);
and \g454493/U$3 ( \27994 , RIe1ea0b0_4040, \8323 );
nor \g454493/U$1 ( \27995 , \27993 , \27994 );
not \g450504/U$3 ( \27996 , \27995 );
not \g450504/U$4 ( \27997 , \8328 );
and \g450504/U$2 ( \27998 , \27996 , \27997 );
and \g450504/U$5 ( \27999 , \8359 , RIe1d38b0_3784);
nor \g450504/U$1 ( \28000 , \27998 , \27999 );
nand \g447991/U$1 ( \28001 , \27986 , \27989 , \27992 , \28000 );
nor \g446473/U$1 ( \28002 , \27981 , \27982 , \28001 );
and \g454014/U$2 ( \28003 , \8378 , RIe1d92b0_3848);
and \g454014/U$3 ( \28004 , RIe1cdeb0_3720, \8531 );
nor \g454014/U$1 ( \28005 , \28003 , \28004 );
and \g454015/U$2 ( \28006 , \8356 , RIe1cb1b0_3688);
and \g454015/U$3 ( \28007 , RIe1decb0_3912, \8407 );
nor \g454015/U$1 ( \28008 , \28006 , \28007 );
and \g445479/U$2 ( \28009 , \28002 , \28005 , \28008 );
nor \g445479/U$1 ( \28010 , \28009 , \8477 );
nor \g444823/U$1 ( \28011 , \27980 , \28010 );
and \g447213/U$2 ( \28012 , \11762 , RIe1ef3a8_4099);
and \g447213/U$3 ( \28013 , RIf14e460_5350, \11764 );
nor \g447213/U$1 ( \28014 , \28012 , \28013 );
nand \g444441/U$1 ( \28015 , \27955 , \28011 , \28014 );
and \g454025/U$2 ( \28016 , \8324 , RIe1bd0b0_3528);
and \g454025/U$3 ( \28017 , RIe1a19f0_3216, \8404 );
nor \g454025/U$1 ( \28018 , \28016 , \28017 );
and \g446474/U$2 ( \28019 , RIe1a46f0_3248, \8373 );
and \g446474/U$3 ( \28020 , RIe1aff28_3379, \8319 );
and \g449486/U$2 ( \28021 , RIe227d48_4743, \8412 );
and \g449486/U$3 ( \28022 , \8407 , RIe17a3f0_2768);
and \g449486/U$4 ( \28023 , RIe1a73f0_3280, \8383 );
nor \g449486/U$1 ( \28024 , \28021 , \28022 , \28023 );
and \g454028/U$2 ( \28025 , \8356 , RIe1f20a8_4131);
and \g454028/U$3 ( \28026 , RIe206148_4359, \8359 );
nor \g454028/U$1 ( \28027 , \28025 , \28026 );
and \g455395/U$2 ( \28028 , \8313 , RIe1f9560_4214);
and \g455395/U$3 ( \28029 , RIe2001a8_4291, \8323 );
nor \g455395/U$1 ( \28030 , \28028 , \28029 );
not \g450508/U$3 ( \28031 , \28030 );
not \g450508/U$4 ( \28032 , \8347 );
and \g450508/U$2 ( \28033 , \28031 , \28032 );
and \g450508/U$5 ( \28034 , \8351 , RIe1aa0f0_3312);
nor \g450508/U$1 ( \28035 , \28033 , \28034 );
and \g454027/U$2 ( \28036 , \8378 , RIe21c948_4615);
and \g454027/U$3 ( \28037 , RIe18def0_2992, \8417 );
nor \g454027/U$1 ( \28038 , \28036 , \28037 );
nand \g447992/U$1 ( \28039 , \28024 , \28027 , \28035 , \28038 );
nor \g446474/U$1 ( \28040 , \28019 , \28020 , \28039 );
and \g454026/U$2 ( \28041 , \8335 , RIe172560_2678);
and \g454026/U$3 ( \28042 , RIe1d65b0_3816, \8340 );
nor \g454026/U$1 ( \28043 , \28041 , \28042 );
nand \g445697/U$1 ( \28044 , \28018 , \28040 , \28043 );
and \g444886/U$2 ( \28045 , \28044 , \9010 );
and \g449484/U$2 ( \28046 , RIe1ba680_3498, \8373 );
and \g449484/U$3 ( \28047 , \8383 , RIf14be68_5323);
and \g449484/U$4 ( \28048 , RIf1481f0_5280, \8488 );
nor \g449484/U$1 ( \28049 , \28046 , \28047 , \28048 );
and \g454024/U$2 ( \28050 , \8335 , RIe1abd10_3332);
and \g454024/U$3 ( \28051 , RIfc69470_6220, \8340 );
nor \g454024/U$1 ( \28052 , \28050 , \28051 );
and \g454022/U$2 ( \28053 , \8404 , RIfe9be80_8118);
and \g454022/U$3 ( \28054 , RIfc4d6a8_5903, \8351 );
nor \g454022/U$1 ( \28055 , \28053 , \28054 );
and \g455016/U$2 ( \28056 , \8313 , RIfe9bbb0_8116);
and \g455016/U$3 ( \28057 , RIfcbfac8_7203, \8323 );
nor \g455016/U$1 ( \28058 , \28056 , \28057 );
not \g455015/U$1 ( \28059 , \28058 );
and \g450506/U$2 ( \28060 , \28059 , \8316 );
and \g450506/U$3 ( \28061 , RIf1495a0_5294, \8359 );
nor \g450506/U$1 ( \28062 , \28060 , \28061 );
nand \g448248/U$1 ( \28063 , \28049 , \28052 , \28055 , \28062 );
and \g444886/U$3 ( \28064 , \8482 , \28063 );
nor \g444886/U$1 ( \28065 , \28045 , \28064 );
and \g447215/U$2 ( \28066 , \8964 , RIfcd46a8_7439);
and \g447215/U$3 ( \28067 , RIfc86e58_6557, \8966 );
nor \g447215/U$1 ( \28068 , \28066 , \28067 );
and \g447216/U$2 ( \28069 , \8521 , RIe1b1e18_3401);
and \g447216/U$3 ( \28070 , RIe1b3600_3418, \8525 );
nor \g447216/U$1 ( \28071 , \28069 , \28070 );
and \g447217/U$2 ( \28072 , \8974 , RIfe9bd18_8117);
and \g447217/U$3 ( \28073 , RIe1b6300_3450, \8976 );
nor \g447217/U$1 ( \28074 , \28072 , \28073 );
nand \g444666/U$1 ( \28075 , \28065 , \28068 , \28071 , \28074 );
and \g446468/U$2 ( \28076 , RIe177858_2737, \8371 );
and \g446468/U$3 ( \28077 , RIf16e9e0_5718, \8319 );
and \g449478/U$2 ( \28078 , RIee3e878_5170, \8414 );
and \g449478/U$3 ( \28079 , \8409 , RIfca54e8_6903);
and \g449478/U$4 ( \28080 , RIf141710_5204, \8383 );
nor \g449478/U$1 ( \28081 , \28078 , \28079 , \28080 );
and \g453999/U$2 ( \28082 , \8356 , RIe174b58_2705);
and \g453999/U$3 ( \28083 , RIee3c988_5148, \8359 );
nor \g453999/U$1 ( \28084 , \28082 , \28083 );
and \g455260/U$2 ( \28085 , \8313 , RIee3a4f8_5122);
and \g455260/U$3 ( \28086 , RIee3b5d8_5134, \8323 );
nor \g455260/U$1 ( \28087 , \28085 , \28086 );
not \g450499/U$3 ( \28088 , \28087 );
not \g450499/U$4 ( \28089 , \8347 );
and \g450499/U$2 ( \28090 , \28088 , \28089 );
and \g450499/U$5 ( \28091 , \8351 , RIf142688_5215);
nor \g450499/U$1 ( \28092 , \28090 , \28091 );
and \g453998/U$2 ( \28093 , \8378 , RIee3dbd0_5161);
and \g453998/U$3 ( \28094 , RIfcea638_7689, \8417 );
nor \g453998/U$1 ( \28095 , \28093 , \28094 );
nand \g447988/U$1 ( \28096 , \28081 , \28084 , \28092 , \28095 );
nor \g446468/U$1 ( \28097 , \28076 , \28077 , \28096 );
and \g453997/U$2 ( \28098 , \8335 , RIfced608_7723);
and \g453997/U$3 ( \28099 , RIf170600_5738, \8340 );
nor \g453997/U$1 ( \28100 , \28098 , \28099 );
and \g453996/U$2 ( \28101 , \8324 , RIfc76fd0_6376);
and \g453996/U$3 ( \28102 , RIe176778_2725, \8404 );
nor \g453996/U$1 ( \28103 , \28101 , \28102 );
and \g445476/U$2 ( \28104 , \28097 , \28100 , \28103 );
nor \g445476/U$1 ( \28105 , \28104 , \8558 );
and \g446469/U$2 ( \28106 , RIf144de8_5243, \8417 );
and \g446469/U$3 ( \28107 , RIe1857f0_2896, \8356 );
and \g449479/U$2 ( \28108 , RIe17fdf0_2832, \8319 );
and \g449479/U$3 ( \28109 , \8326 , RIe182af0_2864);
and \g449479/U$4 ( \28110 , RIe1884f0_2928, \8488 );
nor \g449479/U$1 ( \28111 , \28108 , \28109 , \28110 );
and \g454006/U$2 ( \28112 , \8335 , RIe17d0f0_2800);
and \g454006/U$3 ( \28113 , RIf143060_5222, \8340 );
nor \g454006/U$1 ( \28114 , \28112 , \28113 );
and \g454005/U$2 ( \28115 , \8404 , RIe1992f0_3120);
and \g454005/U$3 ( \28116 , RIe19ecf0_3184, \8351 );
nor \g454005/U$1 ( \28117 , \28115 , \28116 );
and \g455019/U$2 ( \28118 , \8313 , RIf145a90_5252);
and \g455019/U$3 ( \28119 , RIe19bff0_3152, \8323 );
nor \g455019/U$1 ( \28120 , \28118 , \28119 );
not \g450502/U$3 ( \28121 , \28120 );
not \g450502/U$4 ( \28122 , \8328 );
and \g450502/U$2 ( \28123 , \28121 , \28122 );
and \g450502/U$5 ( \28124 , \8359 , RIe18b1f0_2960);
nor \g450502/U$1 ( \28125 , \28123 , \28124 );
nand \g447989/U$1 ( \28126 , \28111 , \28114 , \28117 , \28125 );
nor \g446469/U$1 ( \28127 , \28106 , \28107 , \28126 );
and \g454002/U$2 ( \28128 , \8378 , RIe190bf0_3024);
and \g454002/U$3 ( \28129 , RIfc72980_6326, \8531 );
nor \g454002/U$1 ( \28130 , \28128 , \28129 );
and \g454001/U$2 ( \28131 , \8412 , RIe1938f0_3056);
and \g454001/U$3 ( \28132 , RIe1965f0_3088, \8409 );
nor \g454001/U$1 ( \28133 , \28131 , \28132 );
and \g445478/U$2 ( \28134 , \28127 , \28130 , \28133 );
nor \g445478/U$1 ( \28135 , \28134 , \8589 );
or \g444312/U$1 ( \28136 , \28015 , \28075 , \28105 , \28135 );
and \g446466/U$2 ( \28137 , RIe21f648_4647, \8407 );
and \g446466/U$3 ( \28138 , RIe216f48_4551, \8378 );
and \g449474/U$2 ( \28139 , RIf16c550_5692, \8373 );
and \g449474/U$3 ( \28140 , \8383 , RIe225048_4711);
and \g449474/U$4 ( \28141 , RIe214248_4519, \8488 );
nor \g449474/U$1 ( \28142 , \28139 , \28140 , \28141 );
and \g453988/U$2 ( \28143 , \8335 , RIe208e48_4391);
and \g453988/U$3 ( \28144 , RIf1684a0_5646, \8340 );
nor \g453988/U$1 ( \28145 , \28143 , \28144 );
and \g453987/U$2 ( \28146 , \8404 , RIe222348_4679);
and \g453987/U$3 ( \28147 , RIf16d090_5700, \8351 );
nor \g453987/U$1 ( \28148 , \28146 , \28147 );
and \g455411/U$2 ( \28149 , \8313 , RIe20bb48_4423);
and \g455411/U$3 ( \28150 , RIe20e848_4455, \8323 );
nor \g455411/U$1 ( \28151 , \28149 , \28150 );
not \g455410/U$1 ( \28152 , \28151 );
and \g450496/U$2 ( \28153 , \28152 , \8316 );
and \g450496/U$3 ( \28154 , RIf16a4f8_5669, \8359 );
nor \g450496/U$1 ( \28155 , \28153 , \28154 );
nand \g448247/U$1 ( \28156 , \28142 , \28145 , \28148 , \28155 );
nor \g446466/U$1 ( \28157 , \28137 , \28138 , \28156 );
and \g453983/U$2 ( \28158 , \8356 , RIe211548_4487);
and \g453983/U$3 ( \28159 , RIf16b470_5680, \8417 );
nor \g453983/U$1 ( \28160 , \28158 , \28159 );
and \g453982/U$2 ( \28161 , \8523 , RIf169df0_5664);
and \g453982/U$3 ( \28162 , RIe219c48_4583, \8414 );
nor \g453982/U$1 ( \28163 , \28161 , \28162 );
and \g445474/U$2 ( \28164 , \28157 , \28160 , \28163 );
nor \g445474/U$1 ( \28165 , \28164 , \8368 );
and \g446467/U$2 ( \28166 , RIfcc4550_7256, \8409 );
and \g446467/U$3 ( \28167 , RIf162500_5578, \8378 );
and \g449477/U$2 ( \28168 , RIfc4d540_5902, \8319 );
and \g449477/U$3 ( \28169 , \8324 , RIf15bfc0_5506);
and \g449477/U$4 ( \28170 , RIf15f0f8_5541, \8488 );
nor \g449477/U$1 ( \28171 , \28168 , \28169 , \28170 );
and \g453992/U$2 ( \28172 , \8335 , RIfc9c848_6803);
and \g453992/U$3 ( \28173 , RIf15d208_5519, \8340 );
nor \g453992/U$1 ( \28174 , \28172 , \28173 );
and \g453993/U$2 ( \28175 , \8404 , RIfe9c150_8120);
and \g453993/U$3 ( \28176 , RIf1673c0_5634, \8351 );
nor \g453993/U$1 ( \28177 , \28175 , \28176 );
and \g455394/U$2 ( \28178 , \8313 , RIfe9c6f0_8124);
and \g455394/U$3 ( \28179 , RIf166448_5623, \8323 );
nor \g455394/U$1 ( \28180 , \28178 , \28179 );
not \g450498/U$3 ( \28181 , \28180 );
not \g450498/U$4 ( \28182 , \8328 );
and \g450498/U$2 ( \28183 , \28181 , \28182 );
and \g450498/U$5 ( \28184 , \8359 , RIf160fe8_5563);
nor \g450498/U$1 ( \28185 , \28183 , \28184 );
nand \g447987/U$1 ( \28186 , \28171 , \28174 , \28177 , \28185 );
nor \g446467/U$1 ( \28187 , \28166 , \28167 , \28186 );
and \g453991/U$2 ( \28188 , \8356 , RIfe9c588_8123);
and \g453991/U$3 ( \28189 , RIf1654d0_5612, \8417 );
nor \g453991/U$1 ( \28190 , \28188 , \28189 );
and \g453990/U$2 ( \28191 , \8531 , RIfe9bfe8_8119);
and \g453990/U$3 ( \28192 , RIf1635e0_5590, \8414 );
nor \g453990/U$1 ( \28193 , \28191 , \28192 );
and \g445475/U$2 ( \28194 , \28187 , \28190 , \28193 );
nor \g445475/U$1 ( \28195 , \28194 , \8422 );
or \g444236/U$1 ( \28196 , \28136 , \28165 , \28195 );
_DC \g4c9d/U$1 ( \28197 , \28196 , \8654 );
and \g450789/U$2 ( \28198 , \16313 , RIee23fc8_4868);
and \g450789/U$3 ( \28199 , RIfc6af28_6239, \16319 );
nor \g450789/U$1 ( \28200 , \28198 , \28199 );
and \g445753/U$2 ( \28201 , RIee25be8_4888, \16326 );
and \g445753/U$3 ( \28202 , RIdedfdf0_1011, \16334 );
and \g448558/U$2 ( \28203 , RIded87d0_927, \16398 );
and \g448558/U$3 ( \28204 , \16339 , RIfe8f6d0_7976);
and \g448558/U$4 ( \28205 , RIdee4008_1058, \16485 );
nor \g448558/U$1 ( \28206 , \28203 , \28204 , \28205 );
and \g454499/U$2 ( \28207 , \16317 , RIfc534e0_5970);
and \g454499/U$3 ( \28208 , RIfc6b090_6240, \16325 );
nor \g454499/U$1 ( \28209 , \28207 , \28208 );
not \g449585/U$3 ( \28210 , \28209 );
not \g449585/U$4 ( \28211 , \16351 );
and \g449585/U$2 ( \28212 , \28210 , \28211 );
and \g449585/U$5 ( \28213 , \16354 , RIdee5d90_1079);
nor \g449585/U$1 ( \28214 , \28212 , \28213 );
and \g450793/U$2 ( \28215 , \16361 , RIded42e8_878);
and \g450793/U$3 ( \28216 , RIfe8f568_7975, \16364 );
nor \g450793/U$1 ( \28217 , \28215 , \28216 );
and \g450792/U$2 ( \28218 , \16368 , RIfc66770_6188);
and \g450792/U$3 ( \28219 , RIfca5920_6906, \16371 );
nor \g450792/U$1 ( \28220 , \28218 , \28219 );
nand \g447486/U$1 ( \28221 , \28206 , \28214 , \28217 , \28220 );
nor \g445753/U$1 ( \28222 , \28201 , \28202 , \28221 );
and \g450790/U$2 ( \28223 , \16377 , RIfccf680_7382);
and \g450790/U$3 ( \28224 , RIdee1ce0_1033, \16380 );
nor \g450790/U$1 ( \28225 , \28223 , \28224 );
nand \g445518/U$1 ( \28226 , \28200 , \28222 , \28225 );
and \g444905/U$2 ( \28227 , \28226 , \16477 );
and \g448557/U$2 ( \28228 , RIde9a0e8_341, \16485 );
and \g448557/U$3 ( \28229 , \16356 , RIdeb5dc0_533);
and \g448557/U$4 ( \28230 , RIdee8a90_1111, \16398 );
nor \g448557/U$1 ( \28231 , \28228 , \28229 , \28230 );
and \g454251/U$2 ( \28232 , \16317 , RIdecf2c0_821);
and \g454251/U$3 ( \28233 , RIded1fc0_853, \16325 );
nor \g454251/U$1 ( \28234 , \28232 , \28233 );
not \g449584/U$3 ( \28235 , \28234 );
not \g449584/U$4 ( \28236 , \16311 );
and \g449584/U$2 ( \28237 , \28235 , \28236 );
and \g449584/U$5 ( \28238 , \16339 , RIdf01f90_1399);
nor \g449584/U$1 ( \28239 , \28237 , \28238 );
and \g450784/U$2 ( \28240 , \16377 , RIdec98c0_757);
and \g450784/U$3 ( \28241 , RIdecc5c0_789, \16313 );
nor \g450784/U$1 ( \28242 , \28240 , \28241 );
and \g450785/U$2 ( \28243 , \16334 , RIe15b7c0_2418);
and \g450785/U$3 ( \28244 , RIe16f9c8_2647, \16380 );
nor \g450785/U$1 ( \28245 , \28243 , \28244 );
nand \g447252/U$1 ( \28246 , \28231 , \28239 , \28242 , \28245 );
and \g444905/U$3 ( \28247 , \16752 , \28246 );
nor \g444905/U$1 ( \28248 , \28227 , \28247 );
and \g446549/U$2 ( \28249 , \16774 , RIde80030_214);
and \g446549/U$3 ( \28250 , RIdedd7f8_984, \16776 );
nor \g446549/U$1 ( \28251 , \28249 , \28250 );
and \g446548/U$2 ( \28252 , \16779 , RIdf1e898_1724);
and \g446548/U$3 ( \28253 , RIdf2e018_1900, \16781 );
nor \g446548/U$1 ( \28254 , \28252 , \28253 );
and \g446547/U$2 ( \28255 , \16784 , RIdf399b8_2032);
and \g446547/U$3 ( \28256 , RIe144fc0_2162, \16786 );
nor \g446547/U$1 ( \28257 , \28255 , \28256 );
nand \g444555/U$1 ( \28258 , \28248 , \28251 , \28254 , \28257 );
and \g448552/U$2 ( \28259 , RIdebe4c0_629, \16485 );
and \g448552/U$3 ( \28260 , \16356 , RIee1f978_4818);
and \g448552/U$4 ( \28261 , RIdead6c0_437, \16337 );
nor \g448552/U$1 ( \28262 , \28259 , \28260 , \28261 );
and \g454669/U$2 ( \28263 , \16317 , RIdec3ec0_693);
and \g454669/U$3 ( \28264 , RIdec6bc0_725, \16325 );
nor \g454669/U$1 ( \28265 , \28263 , \28264 );
not \g449581/U$3 ( \28266 , \28265 );
not \g449581/U$4 ( \28267 , \16311 );
and \g449581/U$2 ( \28268 , \28266 , \28267 );
and \g449581/U$5 ( \28269 , \16341 , RIfc5e4a8_6095);
nor \g449581/U$1 ( \28270 , \28268 , \28269 );
and \g450774/U$2 ( \28271 , \16377 , RIdec11c0_661);
and \g450774/U$3 ( \28272 , RIee20a58_4830, \16313 );
nor \g450774/U$1 ( \28273 , \28271 , \28272 );
and \g450775/U$2 ( \28274 , \16334 , RIdeb8ac0_565);
and \g450775/U$3 ( \28275 , RIdebb7c0_597, \16380 );
nor \g450775/U$1 ( \28276 , \28274 , \28275 );
nand \g447250/U$1 ( \28277 , \28262 , \28270 , \28273 , \28276 );
and \g444702/U$2 ( \28278 , \28277 , \17938 );
and \g445750/U$2 ( \28279 , RIee34af8_5058, \16328 );
and \g445750/U$3 ( \28280 , RIfcbcf30_7172, \16377 );
and \g448556/U$2 ( \28281 , RIee30610_5009, \16427 );
and \g448556/U$3 ( \28282 , \16448 , RIfc731f0_6332);
and \g448556/U$4 ( \28283 , RIe140100_2106, \16485 );
nor \g448556/U$1 ( \28284 , \28281 , \28282 , \28283 );
and \g454247/U$2 ( \28285 , \16317 , RIfec3048_8339);
and \g454247/U$3 ( \28286 , RIfec2ee0_8338, \16325 );
nor \g454247/U$1 ( \28287 , \28285 , \28286 );
not \g454246/U$1 ( \28288 , \28287 );
and \g449583/U$2 ( \28289 , \28288 , \16336 );
and \g449583/U$3 ( \28290 , RIe142428_2131, \16354 );
nor \g449583/U$1 ( \28291 , \28289 , \28290 );
and \g450782/U$2 ( \28292 , \16361 , RIfec2d78_8337);
and \g450782/U$3 ( \28293 , RIfec2c10_8336, \16364 );
nor \g450782/U$1 ( \28294 , \28292 , \28293 );
and \g450781/U$2 ( \28295 , \16368 , RIee2e450_4985);
and \g450781/U$3 ( \28296 , RIfcbe010_7184, \16371 );
nor \g450781/U$1 ( \28297 , \28295 , \28296 );
nand \g448011/U$1 ( \28298 , \28284 , \28291 , \28294 , \28297 );
nor \g445750/U$1 ( \28299 , \28279 , \28280 , \28298 );
and \g450779/U$2 ( \28300 , \16334 , RIdf3bb78_2056);
and \g450779/U$3 ( \28301 , RIee327d0_5033, \16313 );
nor \g450779/U$1 ( \28302 , \28300 , \28301 );
and \g450778/U$2 ( \28303 , \16380 , RIfea7280_8218);
and \g450778/U$3 ( \28304 , RIee33a18_5046, \16321 );
nor \g450778/U$1 ( \28305 , \28303 , \28304 );
and \g444964/U$2 ( \28306 , \28299 , \28302 , \28305 );
nor \g444964/U$1 ( \28307 , \28306 , \16393 );
nor \g444702/U$1 ( \28308 , \28278 , \28307 );
and \g446544/U$2 ( \28309 , \18457 , RIdeb30c0_501);
and \g446544/U$3 ( \28310 , RIee1efa0_4811, \18459 );
nor \g446544/U$1 ( \28311 , \28309 , \28310 );
and \g446545/U$2 ( \28312 , \18462 , RIdeb03c0_469);
and \g446545/U$3 ( \28313 , RIfcb04b0_7028, \18464 );
nor \g446545/U$1 ( \28314 , \28312 , \28313 );
and \g446546/U$2 ( \28315 , \18467 , RIdea09e8_373);
and \g446546/U$3 ( \28316 , RIdea72e8_405, \18469 );
nor \g446546/U$1 ( \28317 , \28315 , \28316 );
nand \g444452/U$1 ( \28318 , \28308 , \28311 , \28314 , \28317 );
and \g445747/U$2 ( \28319 , RIe166bc0_2546, \16326 );
and \g445747/U$3 ( \28320 , RIe155dc0_2354, \16334 );
and \g448548/U$2 ( \28321 , RIe1530c0_2322, \16427 );
and \g448548/U$3 ( \28322 , \16448 , RIee35a70_5069);
and \g448548/U$4 ( \28323 , RIe15e4c0_2450, \16485 );
nor \g448548/U$1 ( \28324 , \28321 , \28322 , \28323 );
and \g454240/U$2 ( \28325 , \16317 , RIe14d6c0_2258);
and \g454240/U$3 ( \28326 , RIfc9fdb8_6841, \16325 );
nor \g454240/U$1 ( \28327 , \28325 , \28326 );
not \g454239/U$1 ( \28328 , \28327 );
and \g449574/U$2 ( \28329 , \28328 , \16336 );
and \g449574/U$3 ( \28330 , RIfc54b60_5986, \16356 );
nor \g449574/U$1 ( \28331 , \28329 , \28330 );
and \g450767/U$2 ( \28332 , \16361 , RIe147cc0_2194);
and \g450767/U$3 ( \28333 , RIe14a9c0_2226, \16364 );
nor \g450767/U$1 ( \28334 , \28332 , \28333 );
and \g450766/U$2 ( \28335 , \16368 , RIe1503c0_2290);
and \g450766/U$3 ( \28336 , RIee357a0_5067, \16371 );
nor \g450766/U$1 ( \28337 , \28335 , \28336 );
nand \g448010/U$1 ( \28338 , \28324 , \28331 , \28334 , \28337 );
nor \g445747/U$1 ( \28339 , \28319 , \28320 , \28338 );
and \g450764/U$2 ( \28340 , \16377 , RIe1611c0_2482);
and \g450764/U$3 ( \28341 , RIe158ac0_2386, \16380 );
nor \g450764/U$1 ( \28342 , \28340 , \28341 );
and \g450763/U$2 ( \28343 , \16313 , RIee38338_5098);
and \g450763/U$3 ( \28344 , RIe163ec0_2514, \16321 );
nor \g450763/U$1 ( \28345 , \28343 , \28344 );
and \g444961/U$2 ( \28346 , \28339 , \28342 , \28345 );
nor \g444961/U$1 ( \28347 , \28346 , \16389 );
and \g445748/U$2 ( \28348 , RIfc7bd28_6431, \16427 );
and \g445748/U$3 ( \28349 , RIfc7a108_6411, \16368 );
and \g448550/U$2 ( \28350 , RIfea7820_8222, \16485 );
and \g448550/U$3 ( \28351 , \16356 , RIde93b30_310);
and \g448550/U$4 ( \28352 , RIe16ccc8_2615, \16398 );
nor \g448550/U$1 ( \28353 , \28350 , \28351 , \28352 );
and \g454243/U$2 ( \28354 , \16317 , RIfcd16d8_7405);
and \g454243/U$3 ( \28355 , RIfcb2508_7051, \16325 );
nor \g454243/U$1 ( \28356 , \28354 , \28355 );
not \g449579/U$3 ( \28357 , \28356 );
not \g449579/U$4 ( \28358 , \16311 );
and \g449579/U$2 ( \28359 , \28357 , \28358 );
and \g449579/U$5 ( \28360 , \16339 , RIfc7a6a8_6415);
nor \g449579/U$1 ( \28361 , \28359 , \28360 );
and \g450770/U$2 ( \28362 , \16377 , RIfc63d40_6158);
and \g450770/U$3 ( \28363 , RIfc5d800_6086, \16313 );
nor \g450770/U$1 ( \28364 , \28362 , \28363 );
and \g450771/U$2 ( \28365 , \16334 , RIde87998_251);
and \g450771/U$3 ( \28366 , RIfea73e8_8219, \16380 );
nor \g450771/U$1 ( \28367 , \28365 , \28366 );
nand \g447249/U$1 ( \28368 , \28353 , \28361 , \28364 , \28367 );
nor \g445748/U$1 ( \28369 , \28348 , \28349 , \28368 );
and \g450769/U$2 ( \28370 , \16361 , RIe1691b8_2573);
and \g450769/U$3 ( \28371 , RIde837f8_231, \16448 );
nor \g450769/U$1 ( \28372 , \28370 , \28371 );
and \g450768/U$2 ( \28373 , \16364 , RIe16a838_2589);
and \g450768/U$3 ( \28374 , RIfcc7ef8_7297, \16371 );
nor \g450768/U$1 ( \28375 , \28373 , \28374 );
and \g444962/U$2 ( \28376 , \28369 , \28372 , \28375 );
nor \g444962/U$1 ( \28377 , \28376 , \16649 );
or \g444339/U$1 ( \28378 , \28258 , \28318 , \28347 , \28377 );
and \g445743/U$2 ( \28379 , RIdf18790_1655, \16328 );
and \g445743/U$3 ( \28380 , RIdf04c90_1431, \16334 );
and \g448546/U$2 ( \28381 , RIdefc590_1335, \16427 );
and \g448546/U$3 ( \28382 , \16448 , RIdeff290_1367);
and \g448546/U$4 ( \28383 , RIdf0a690_1495, \16485 );
nor \g448546/U$1 ( \28384 , \28381 , \28382 , \28383 );
and \g454288/U$2 ( \28385 , \16317 , RIdef1190_1207);
and \g454288/U$3 ( \28386 , RIdef3e90_1239, \16325 );
nor \g454288/U$1 ( \28387 , \28385 , \28386 );
not \g454287/U$1 ( \28388 , \28387 );
and \g449571/U$2 ( \28389 , \28388 , \16336 );
and \g449571/U$3 ( \28390 , RIdf0d390_1527, \16356 );
nor \g449571/U$1 ( \28391 , \28389 , \28390 );
and \g450752/U$2 ( \28392 , \16361 , RIdeeb790_1143);
and \g450752/U$3 ( \28393 , RIdeee490_1175, \16364 );
nor \g450752/U$1 ( \28394 , \28392 , \28393 );
and \g450750/U$2 ( \28395 , \16368 , RIdef6b90_1271);
and \g450750/U$3 ( \28396 , RIdef9890_1303, \16371 );
nor \g450750/U$1 ( \28397 , \28395 , \28396 );
nand \g448009/U$1 ( \28398 , \28384 , \28391 , \28394 , \28397 );
nor \g445743/U$1 ( \28399 , \28379 , \28380 , \28398 );
and \g450749/U$2 ( \28400 , \16377 , RIdf10090_1559);
and \g450749/U$3 ( \28401 , RIdf07990_1463, \16380 );
nor \g450749/U$1 ( \28402 , \28400 , \28401 );
and \g450748/U$2 ( \28403 , \16313 , RIdf12d90_1591);
and \g450748/U$3 ( \28404 , RIdf15a90_1623, \16321 );
nor \g450748/U$1 ( \28405 , \28403 , \28404 );
and \g444958/U$2 ( \28406 , \28399 , \28402 , \28405 );
nor \g444958/U$1 ( \28407 , \28406 , \16555 );
and \g445746/U$2 ( \28408 , RIfcc9de8_7319, \16432 );
and \g445746/U$3 ( \28409 , RIdf1a7e8_1678, \16361 );
and \g448547/U$2 ( \28410 , RIfcb4830_7076, \16319 );
and \g448547/U$3 ( \28411 , \16326 , RIfcb46c8_7075);
and \g448547/U$4 ( \28412 , RIdf20d28_1750, \16398 );
nor \g448547/U$1 ( \28413 , \28410 , \28411 , \28412 );
and \g454238/U$2 ( \28414 , \16317 , RIdf29590_1847);
and \g454238/U$3 ( \28415 , RIdf2b480_1869, \16325 );
nor \g454238/U$1 ( \28416 , \28414 , \28415 );
not \g449572/U$3 ( \28417 , \28416 );
not \g449572/U$4 ( \28418 , \16330 );
and \g449572/U$2 ( \28419 , \28417 , \28418 );
and \g449572/U$5 ( \28420 , \16339 , RIdf223a8_1766);
nor \g449572/U$1 ( \28421 , \28419 , \28420 );
and \g450758/U$2 ( \28422 , \16377 , RIfcb88e0_7122);
and \g450758/U$3 ( \28423 , RIee29860_4931, \16313 );
nor \g450758/U$1 ( \28424 , \28422 , \28423 );
and \g452253/U$2 ( \28425 , \16334 , RIdf25648_1802);
and \g452253/U$3 ( \28426 , RIdf27268_1822, \16380 );
nor \g452253/U$1 ( \28427 , \28425 , \28426 );
nand \g447248/U$1 ( \28428 , \28413 , \28421 , \28424 , \28427 );
nor \g445746/U$1 ( \28429 , \28408 , \28409 , \28428 );
and \g450756/U$2 ( \28430 , \16364 , RIdf1bd00_1693);
and \g450756/U$3 ( \28431 , RIfc823d0_6504, \16368 );
nor \g450756/U$1 ( \28432 , \28430 , \28431 );
and \g450755/U$2 ( \28433 , \16371 , RIdf23a28_1782);
and \g450755/U$3 ( \28434 , RIfc53648_5971, \16427 );
nor \g450755/U$1 ( \28435 , \28433 , \28434 );
and \g444959/U$2 ( \28436 , \28429 , \28432 , \28435 );
nor \g444959/U$1 ( \28437 , \28436 , \16480 );
or \g444257/U$1 ( \28438 , \28378 , \28407 , \28437 );
_DC \g4d22/U$1 ( \28439 , \28438 , \16652 );
and \g446557/U$2 ( \28440 , \11511 , RIe1fb450_4236);
and \g446557/U$3 ( \28441 , RIfca2ab8_6873, \11513 );
nor \g446557/U$1 ( \28442 , \28440 , \28441 );
and \g445759/U$2 ( \28443 , RIfc90908_6667, \8324 );
and \g445759/U$3 ( \28444 , RIfc44738_5801, \8340 );
and \g448567/U$2 ( \28445 , RIf151160_5382, \8531 );
and \g448567/U$3 ( \28446 , \8488 , RIfcd9400_7494);
and \g448567/U$4 ( \28447 , RIfc55c40_5998, \8383 );
nor \g448567/U$1 ( \28448 , \28445 , \28446 , \28447 );
and \g450819/U$2 ( \28449 , \8356 , RIe1f4808_4159);
and \g450819/U$3 ( \28450 , RIfcb4b00_7078, \8359 );
nor \g450819/U$1 ( \28451 , \28449 , \28450 );
and \g454171/U$2 ( \28452 , \8313 , RIf154dd8_5425);
and \g454171/U$3 ( \28453 , RIfcd5ff8_7457, \8323 );
nor \g454171/U$1 ( \28454 , \28452 , \28453 );
not \g449593/U$3 ( \28455 , \28454 );
not \g449593/U$4 ( \28456 , \8376 );
and \g449593/U$2 ( \28457 , \28455 , \28456 );
and \g449593/U$5 ( \28458 , \8351 , RIfc4bd58_5885);
nor \g449593/U$1 ( \28459 , \28457 , \28458 );
and \g450818/U$2 ( \28460 , \8378 , RIfec2aa8_8335);
and \g450818/U$3 ( \28461 , RIf156890_5444, \8417 );
nor \g450818/U$1 ( \28462 , \28460 , \28461 );
nand \g447489/U$1 ( \28463 , \28448 , \28451 , \28459 , \28462 );
nor \g445759/U$1 ( \28464 , \28443 , \28444 , \28463 );
not \g444811/U$3 ( \28465 , \28464 );
not \g444811/U$4 ( \28466 , \8621 );
and \g444811/U$2 ( \28467 , \28465 , \28466 );
and \g445760/U$2 ( \28468 , RIe1dee18_3913, \8409 );
and \g445760/U$3 ( \28469 , RIe1d9418_3849, \8378 );
and \g448568/U$2 ( \28470 , RIe1e7518_4009, \8373 );
and \g448568/U$3 ( \28471 , \8383 , RIe1ea218_4041);
and \g448568/U$4 ( \28472 , RIe1d0d18_3753, \8488 );
nor \g448568/U$1 ( \28473 , \28470 , \28471 , \28472 );
and \g450825/U$2 ( \28474 , \8335 , RIe1bff18_3561);
and \g450825/U$3 ( \28475 , RIe1c8618_3657, \8340 );
nor \g450825/U$1 ( \28476 , \28474 , \28475 );
and \g450824/U$2 ( \28477 , \8404 , RIe1e4818_3977);
and \g450824/U$3 ( \28478 , RIe1ecf18_4073, \8351 );
nor \g450824/U$1 ( \28479 , \28477 , \28478 );
and \g454283/U$2 ( \28480 , \8313 , RIe1c2c18_3593);
and \g454283/U$3 ( \28481 , RIe1c5918_3625, \8323 );
nor \g454283/U$1 ( \28482 , \28480 , \28481 );
not \g454282/U$1 ( \28483 , \28482 );
and \g449594/U$2 ( \28484 , \28483 , \8316 );
and \g449594/U$3 ( \28485 , RIe1d3a18_3785, \8359 );
nor \g449594/U$1 ( \28486 , \28484 , \28485 );
nand \g448141/U$1 ( \28487 , \28473 , \28476 , \28479 , \28486 );
nor \g445760/U$1 ( \28488 , \28468 , \28469 , \28487 );
and \g450822/U$2 ( \28489 , \8356 , RIe1cb318_3689);
and \g450822/U$3 ( \28490 , RIe1e1b18_3945, \8417 );
nor \g450822/U$1 ( \28491 , \28489 , \28490 );
and \g450821/U$2 ( \28492 , \8531 , RIe1ce018_3721);
and \g450821/U$3 ( \28493 , RIe1dc118_3881, \8414 );
nor \g450821/U$1 ( \28494 , \28492 , \28493 );
and \g444974/U$2 ( \28495 , \28488 , \28491 , \28494 );
nor \g444974/U$1 ( \28496 , \28495 , \8477 );
nor \g444811/U$1 ( \28497 , \28467 , \28496 );
and \g446556/U$2 ( \28498 , \11762 , RIe1ef510_4100);
and \g446556/U$3 ( \28499 , RIf14e5c8_5351, \11764 );
nor \g446556/U$1 ( \28500 , \28498 , \28499 );
nand \g444417/U$1 ( \28501 , \28442 , \28497 , \28500 );
and \g448570/U$2 ( \28502 , RIfcc65a8_7279, \8319 );
and \g448570/U$3 ( \28503 , \8326 , RIfc53eb8_5977);
and \g448570/U$4 ( \28504 , RIfce08b8_7577, \8486 );
nor \g448570/U$1 ( \28505 , \28502 , \28503 , \28504 );
and \g450831/U$2 ( \28506 , \8335 , RIfc80d50_6488);
and \g450831/U$3 ( \28507 , RIfca04c0_6846, \8340 );
nor \g450831/U$1 ( \28508 , \28506 , \28507 );
and \g450830/U$2 ( \28509 , \8404 , RIe1768e0_2726);
and \g450830/U$3 ( \28510 , RIf1427f0_5216, \8351 );
nor \g450830/U$1 ( \28511 , \28509 , \28510 );
and \g455198/U$2 ( \28512 , \8313 , RIe1779c0_2738);
and \g455198/U$3 ( \28513 , RIfe8efc8_7971, \8323 );
nor \g455198/U$1 ( \28514 , \28512 , \28513 );
not \g449596/U$3 ( \28515 , \28514 );
not \g449596/U$4 ( \28516 , \8328 );
and \g449596/U$2 ( \28517 , \28515 , \28516 );
and \g449596/U$5 ( \28518 , \8359 , RIfce5778_7633);
nor \g449596/U$1 ( \28519 , \28517 , \28518 );
nand \g447490/U$1 ( \28520 , \28505 , \28508 , \28511 , \28519 );
and \g444679/U$2 ( \28521 , \28520 , \9700 );
and \g445761/U$2 ( \28522 , RIe193a58_3057, \8414 );
and \g445761/U$3 ( \28523 , RIfe8f298_7973, \8417 );
and \g448571/U$2 ( \28524 , RIf145bf8_5253, \8373 );
and \g448571/U$3 ( \28525 , \8383 , RIe19c158_3153);
and \g448571/U$4 ( \28526 , RIe188658_2929, \8486 );
nor \g448571/U$1 ( \28527 , \28524 , \28525 , \28526 );
and \g450837/U$2 ( \28528 , \8335 , RIe17d258_2801);
and \g450837/U$3 ( \28529 , RIfc9f278_6833, \8340 );
nor \g450837/U$1 ( \28530 , \28528 , \28529 );
and \g450836/U$2 ( \28531 , \8404 , RIe199458_3121);
and \g450836/U$3 ( \28532 , RIe19ee58_3185, \8351 );
nor \g450836/U$1 ( \28533 , \28531 , \28532 );
and \g454272/U$2 ( \28534 , \8313 , RIe17ff58_2833);
and \g454272/U$3 ( \28535 , RIe182c58_2865, \8323 );
nor \g454272/U$1 ( \28536 , \28534 , \28535 );
not \g454271/U$1 ( \28537 , \28536 );
and \g449599/U$2 ( \28538 , \28537 , \8316 );
and \g449599/U$3 ( \28539 , RIe18b358_2961, \8359 );
nor \g449599/U$1 ( \28540 , \28538 , \28539 );
nand \g448142/U$1 ( \28541 , \28527 , \28530 , \28533 , \28540 );
nor \g445761/U$1 ( \28542 , \28522 , \28523 , \28541 );
and \g450834/U$2 ( \28543 , \8378 , RIe190d58_3025);
and \g450834/U$3 ( \28544 , RIfe8f130_7972, \8531 );
nor \g450834/U$1 ( \28545 , \28543 , \28544 );
and \g450833/U$2 ( \28546 , \8356 , RIe185958_2897);
and \g450833/U$3 ( \28547 , RIe196758_3089, \8409 );
nor \g450833/U$1 ( \28548 , \28546 , \28547 );
and \g444975/U$2 ( \28549 , \28542 , \28545 , \28548 );
nor \g444975/U$1 ( \28550 , \28549 , \8589 );
nor \g444679/U$1 ( \28551 , \28521 , \28550 );
and \g446563/U$2 ( \28552 , \12254 , RIfc81b60_6498);
and \g446563/U$3 ( \28553 , RIfca0088_6843, \12256 );
nor \g446563/U$1 ( \28554 , \28552 , \28553 );
and \g446562/U$2 ( \28555 , \26544 , RIfc9ff20_6842);
and \g446562/U$3 ( \28556 , RIfc81e30_6500, \26546 );
nor \g446562/U$1 ( \28557 , \28555 , \28556 );
and \g446564/U$2 ( \28558 , \12264 , RIe174cc0_2706);
and \g446564/U$3 ( \28559 , RIfc815c0_6494, \12266 );
nor \g446564/U$1 ( \28560 , \28558 , \28559 );
nand \g444454/U$1 ( \28561 , \28551 , \28554 , \28557 , \28560 );
and \g445757/U$2 ( \28562 , RIfc6c170_6252, \8409 );
and \g445757/U$3 ( \28563 , RIe1b49b0_3432, \8378 );
and \g448564/U$2 ( \28564 , RIfea8090_8228, \8371 );
and \g448564/U$3 ( \28565 , \8330 , RIfe8ee60_7970);
and \g448564/U$4 ( \28566 , RIfcaa948_6963, \8488 );
nor \g448564/U$1 ( \28567 , \28564 , \28565 , \28566 );
and \g450810/U$2 ( \28568 , \8335 , RIe1abe78_3333);
and \g450810/U$3 ( \28569 , RIfc67f58_6205, \8340 );
nor \g450810/U$1 ( \28570 , \28568 , \28569 );
and \g450809/U$2 ( \28571 , \8404 , RIe1b84c0_3474);
and \g450809/U$3 ( \28572 , RIf14d218_5337, \8351 );
nor \g450809/U$1 ( \28573 , \28571 , \28572 );
and \g454310/U$2 ( \28574 , \8313 , RIfe8eb90_7968);
and \g454310/U$3 ( \28575 , RIfca8ff8_6945, \8323 );
nor \g454310/U$1 ( \28576 , \28574 , \28575 );
not \g454309/U$1 ( \28577 , \28576 );
and \g449590/U$2 ( \28578 , \28577 , \8316 );
and \g449590/U$3 ( \28579 , RIfcafad8_7021, \8359 );
nor \g449590/U$1 ( \28580 , \28578 , \28579 );
nand \g448137/U$1 ( \28581 , \28567 , \28570 , \28573 , \28580 );
nor \g445757/U$1 ( \28582 , \28562 , \28563 , \28581 );
and \g450808/U$2 ( \28583 , \8356 , RIfe8f400_7974);
and \g450808/U$3 ( \28584 , RIf14aab8_5309, \8417 );
nor \g450808/U$1 ( \28585 , \28583 , \28584 );
and \g450807/U$2 ( \28586 , \8531 , RIfe8ecf8_7969);
and \g450807/U$3 ( \28587 , RIe1b6468_3451, \8412 );
nor \g450807/U$1 ( \28588 , \28586 , \28587 );
and \g444970/U$2 ( \28589 , \28582 , \28585 , \28588 );
nor \g444970/U$1 ( \28590 , \28589 , \8481 );
and \g445758/U$2 ( \28591 , RIe227eb0_4744, \8412 );
and \g445758/U$3 ( \28592 , RIe18e058_2993, \8417 );
and \g448566/U$2 ( \28593 , RIe1a4858_3249, \8373 );
and \g448566/U$3 ( \28594 , \8383 , RIe1a7558_3281);
and \g448566/U$4 ( \28595 , RIe200310_4292, \8488 );
nor \g448566/U$1 ( \28596 , \28593 , \28594 , \28595 );
and \g450817/U$2 ( \28597 , \8335 , RIe1726c8_2679);
and \g450817/U$3 ( \28598 , RIe1d6718_3817, \8340 );
nor \g450817/U$1 ( \28599 , \28597 , \28598 );
and \g450816/U$2 ( \28600 , \8404 , RIe1a1b58_3217);
and \g450816/U$3 ( \28601 , RIe1aa258_3313, \8351 );
nor \g450816/U$1 ( \28602 , \28600 , \28601 );
and \g454305/U$2 ( \28603 , \8313 , RIe1b0090_3380);
and \g454305/U$3 ( \28604 , RIe1bd218_3529, \8323 );
nor \g454305/U$1 ( \28605 , \28603 , \28604 );
not \g454304/U$1 ( \28606 , \28605 );
and \g449592/U$2 ( \28607 , \28606 , \8316 );
and \g449592/U$3 ( \28608 , RIe2062b0_4360, \8359 );
nor \g449592/U$1 ( \28609 , \28607 , \28608 );
nand \g448138/U$1 ( \28610 , \28596 , \28599 , \28602 , \28609 );
nor \g445758/U$1 ( \28611 , \28591 , \28592 , \28610 );
and \g450814/U$2 ( \28612 , \8378 , RIe21cab0_4616);
and \g450814/U$3 ( \28613 , RIe1f96c8_4215, \8531 );
nor \g450814/U$1 ( \28614 , \28612 , \28613 );
and \g450815/U$2 ( \28615 , \8356 , RIe1f2210_4132);
and \g450815/U$3 ( \28616 , RIe17a558_2769, \8409 );
nor \g450815/U$1 ( \28617 , \28615 , \28616 );
and \g444972/U$2 ( \28618 , \28611 , \28614 , \28617 );
nor \g444972/U$1 ( \28619 , \28618 , \8651 );
or \g444289/U$1 ( \28620 , \28501 , \28561 , \28590 , \28619 );
and \g445754/U$2 ( \28621 , RIfc80378_6481, \8373 );
and \g445754/U$3 ( \28622 , RIe20bcb0_4424, \8319 );
and \g448561/U$2 ( \28623 , RIfc82c40_6510, \8523 );
and \g448561/U$3 ( \28624 , \8488 , RIe2143b0_4520);
and \g448561/U$4 ( \28625 , RIe2251b0_4712, \8383 );
nor \g448561/U$1 ( \28626 , \28623 , \28624 , \28625 );
and \g450800/U$2 ( \28627 , \8356 , RIe2116b0_4488);
and \g450800/U$3 ( \28628 , RIfca01f0_6844, \8359 );
nor \g450800/U$1 ( \28629 , \28627 , \28628 );
and \g454259/U$2 ( \28630 , \8313 , RIe219db0_4584);
and \g454259/U$3 ( \28631 , RIe21f7b0_4648, \8323 );
nor \g454259/U$1 ( \28632 , \28630 , \28631 );
not \g449588/U$3 ( \28633 , \28632 );
not \g449588/U$4 ( \28634 , \8376 );
and \g449588/U$2 ( \28635 , \28633 , \28634 );
and \g449588/U$5 ( \28636 , \8351 , RIfc804e0_6482);
nor \g449588/U$1 ( \28637 , \28635 , \28636 );
and \g450799/U$2 ( \28638 , \8378 , RIe2170b0_4552);
and \g450799/U$3 ( \28639 , RIfcb5910_7088, \8417 );
nor \g450799/U$1 ( \28640 , \28638 , \28639 );
nand \g447487/U$1 ( \28641 , \28626 , \28629 , \28637 , \28640 );
nor \g445754/U$1 ( \28642 , \28621 , \28622 , \28641 );
and \g450798/U$2 ( \28643 , \8335 , RIe208fb0_4392);
and \g450798/U$3 ( \28644 , RIfc7f6d0_6472, \8340 );
nor \g450798/U$1 ( \28645 , \28643 , \28644 );
and \g450797/U$2 ( \28646 , \8326 , RIe20e9b0_4456);
and \g450797/U$3 ( \28647 , RIe2224b0_4680, \8404 );
nor \g450797/U$1 ( \28648 , \28646 , \28647 );
and \g444968/U$2 ( \28649 , \28642 , \28645 , \28648 );
nor \g444968/U$1 ( \28650 , \28649 , \8368 );
and \g445755/U$2 ( \28651 , RIe203718_4329, \8371 );
and \g445755/U$3 ( \28652 , RIfcc5d38_7273, \8317 );
and \g448563/U$2 ( \28653 , RIe1fd610_4260, \8531 );
and \g448563/U$3 ( \28654 , \8488 , RIfc87998_6565);
and \g448563/U$4 ( \28655 , RIf1665b0_5624, \8383 );
nor \g448563/U$1 ( \28656 , \28653 , \28654 , \28655 );
and \g450804/U$2 ( \28657 , \8356 , RIe1fc3c8_4247);
and \g450804/U$3 ( \28658 , RIfc7e320_6458, \8359 );
nor \g450804/U$1 ( \28659 , \28657 , \28658 );
and \g454374/U$2 ( \28660 , \8313 , RIf163748_5591);
and \g454374/U$3 ( \28661 , RIfcc5360_7266, \8323 );
nor \g454374/U$1 ( \28662 , \28660 , \28661 );
not \g449589/U$3 ( \28663 , \28662 );
not \g449589/U$4 ( \28664 , \8376 );
and \g449589/U$2 ( \28665 , \28663 , \28664 );
and \g449589/U$5 ( \28666 , \8351 , RIf167528_5635);
nor \g449589/U$1 ( \28667 , \28665 , \28666 );
and \g450803/U$2 ( \28668 , \8378 , RIf162668_5579);
and \g450803/U$3 ( \28669 , RIfc9da90_6816, \8417 );
nor \g450803/U$1 ( \28670 , \28668 , \28669 );
nand \g447488/U$1 ( \28671 , \28656 , \28659 , \28667 , \28670 );
nor \g445755/U$1 ( \28672 , \28651 , \28652 , \28671 );
and \g450802/U$2 ( \28673 , \8335 , RIfce7d70_7660);
and \g450802/U$3 ( \28674 , RIf15d370_5520, \8340 );
nor \g450802/U$1 ( \28675 , \28673 , \28674 );
and \g450801/U$2 ( \28676 , \8326 , RIf15c128_5507);
and \g450801/U$3 ( \28677 , RIe201c60_4310, \8404 );
nor \g450801/U$1 ( \28678 , \28676 , \28677 );
and \g444969/U$2 ( \28679 , \28672 , \28675 , \28678 );
nor \g444969/U$1 ( \28680 , \28679 , \8422 );
or \g444176/U$1 ( \28681 , \28620 , \28650 , \28680 );
_DC \g4da6/U$1 ( \28682 , \28681 , \8654 );
and \g450870/U$2 ( \28683 , \16313 , RIfcba668_7143);
and \g450870/U$3 ( \28684 , RIfc55538_5993, \16321 );
nor \g450870/U$1 ( \28685 , \28683 , \28684 );
and \g445769/U$2 ( \28686 , RIfcbac08_7147, \16328 );
and \g445769/U$3 ( \28687 , RIde87ce0_252, \16334 );
and \g448583/U$2 ( \28688 , RIe16ce30_2616, \16398 );
and \g448583/U$3 ( \28689 , \16341 , RIee39418_5110);
and \g448583/U$4 ( \28690 , RIfe91458_7997, \16485 );
nor \g448583/U$1 ( \28691 , \28688 , \28689 , \28690 );
and \g454286/U$2 ( \28692 , \16317 , RIfc88640_6574);
and \g454286/U$3 ( \28693 , RIfc85238_6537, \16325 );
nor \g454286/U$1 ( \28694 , \28692 , \28693 );
not \g449608/U$3 ( \28695 , \28694 );
not \g449608/U$4 ( \28696 , \16351 );
and \g449608/U$2 ( \28697 , \28695 , \28696 );
and \g449608/U$5 ( \28698 , \16354 , RIfe912f0_7996);
nor \g449608/U$1 ( \28699 , \28697 , \28698 );
and \g450874/U$2 ( \28700 , \16361 , RIe169320_2574);
and \g450874/U$3 ( \28701 , RIfc884d8_6573, \16364 );
nor \g450874/U$1 ( \28702 , \28700 , \28701 );
and \g450873/U$2 ( \28703 , \16368 , RIfcd5788_7451);
and \g450873/U$3 ( \28704 , RIfcda210_7504, \16371 );
nor \g450873/U$1 ( \28705 , \28703 , \28704 );
nand \g447494/U$1 ( \28706 , \28691 , \28699 , \28702 , \28705 );
nor \g445769/U$1 ( \28707 , \28686 , \28687 , \28706 );
and \g451343/U$2 ( \28708 , \16377 , RIfc4af48_5875);
and \g451343/U$3 ( \28709 , RIde8be80_272, \16380 );
nor \g451343/U$1 ( \28710 , \28708 , \28709 );
nand \g445523/U$1 ( \28711 , \28685 , \28707 , \28710 );
and \g444756/U$2 ( \28712 , \28711 , \17998 );
and \g448580/U$2 ( \28713 , RIe153228_2323, \16427 );
and \g448580/U$3 ( \28714 , \16432 , RIfe91188_7995);
and \g448580/U$4 ( \28715 , RIe15e628_2451, \16485 );
nor \g448580/U$1 ( \28716 , \28713 , \28714 , \28715 );
and \g454668/U$2 ( \28717 , \16317 , RIe14d828_2259);
and \g454668/U$3 ( \28718 , RIfcda378_7505, \16325 );
nor \g454668/U$1 ( \28719 , \28717 , \28718 );
not \g454667/U$1 ( \28720 , \28719 );
and \g449607/U$2 ( \28721 , \28720 , \16336 );
and \g449607/U$3 ( \28722 , RIee36880_5079, \16356 );
nor \g449607/U$1 ( \28723 , \28721 , \28722 );
and \g450868/U$2 ( \28724 , \16361 , RIe147e28_2195);
and \g450868/U$3 ( \28725 , RIe14ab28_2227, \16364 );
nor \g450868/U$1 ( \28726 , \28724 , \28725 );
and \g450867/U$2 ( \28727 , \16368 , RIe150528_2291);
and \g450867/U$3 ( \28728 , RIfe91020_7994, \16371 );
nor \g450867/U$1 ( \28729 , \28727 , \28728 );
nand \g448015/U$1 ( \28730 , \28716 , \28723 , \28726 , \28729 );
and \g444756/U$3 ( \28731 , \16390 , \28730 );
nor \g444756/U$1 ( \28732 , \28712 , \28731 );
and \g446568/U$2 ( \28733 , \18020 , RIe164028_2515);
and \g446568/U$3 ( \28734 , RIe166d28_2547, \18022 );
nor \g446568/U$1 ( \28735 , \28733 , \28734 );
and \g446569/U$2 ( \28736 , \18025 , RIe161328_2483);
and \g446569/U$3 ( \28737 , RIfe90918_7989, \18027 );
nor \g446569/U$1 ( \28738 , \28736 , \28737 );
and \g446570/U$2 ( \28739 , \18030 , RIe155f28_2355);
and \g446570/U$3 ( \28740 , RIe158c28_2387, \18032 );
nor \g446570/U$1 ( \28741 , \28739 , \28740 );
nand \g444456/U$1 ( \28742 , \28732 , \28735 , \28738 , \28741 );
and \g448584/U$2 ( \28743 , RIdf15bf8_1624, \16321 );
and \g448584/U$3 ( \28744 , \16326 , RIdf188f8_1656);
and \g448584/U$4 ( \28745 , RIdef12f8_1208, \16398 );
nor \g448584/U$1 ( \28746 , \28743 , \28744 , \28745 );
and \g454289/U$2 ( \28747 , \16317 , RIdf0a7f8_1496);
and \g454289/U$3 ( \28748 , RIdf0d4f8_1528, \16325 );
nor \g454289/U$1 ( \28749 , \28747 , \28748 );
not \g449610/U$3 ( \28750 , \28749 );
not \g449610/U$4 ( \28751 , \16330 );
and \g449610/U$2 ( \28752 , \28750 , \28751 );
and \g449610/U$5 ( \28753 , \16341 , RIdef3ff8_1240);
nor \g449610/U$1 ( \28754 , \28752 , \28753 );
and \g450877/U$2 ( \28755 , \16377 , RIdf101f8_1560);
and \g450877/U$3 ( \28756 , RIdf12ef8_1592, \16313 );
nor \g450877/U$1 ( \28757 , \28755 , \28756 );
and \g450878/U$2 ( \28758 , \16334 , RIdf04df8_1432);
and \g450878/U$3 ( \28759 , RIdf07af8_1464, \16380 );
nor \g450878/U$1 ( \28760 , \28758 , \28759 );
nand \g447258/U$1 ( \28761 , \28746 , \28754 , \28757 , \28760 );
and \g444714/U$2 ( \28762 , \28761 , \16750 );
and \g445772/U$2 ( \28763 , RIfc9d928_6815, \16432 );
and \g445772/U$3 ( \28764 , RIdf1a950_1679, \16361 );
and \g448586/U$2 ( \28765 , RIee2aee0_4947, \16319 );
and \g448586/U$3 ( \28766 , \16328 , RIee2c998_4966);
and \g448586/U$4 ( \28767 , RIdf20e90_1751, \16398 );
nor \g448586/U$1 ( \28768 , \28765 , \28766 , \28767 );
and \g454955/U$2 ( \28769 , \16317 , RIfe907b0_7988);
and \g454955/U$3 ( \28770 , RIfe90378_7985, \16325 );
nor \g454955/U$1 ( \28771 , \28769 , \28770 );
not \g449612/U$3 ( \28772 , \28771 );
not \g449612/U$4 ( \28773 , \16330 );
and \g449612/U$2 ( \28774 , \28772 , \28773 );
and \g449612/U$5 ( \28775 , \16341 , RIfc86a20_6554);
nor \g449612/U$1 ( \28776 , \28774 , \28775 );
and \g450882/U$2 ( \28777 , \16377 , RIee28618_4918);
and \g450882/U$3 ( \28778 , RIee299c8_4932, \16313 );
nor \g450882/U$1 ( \28779 , \28777 , \28778 );
and \g450883/U$2 ( \28780 , \16334 , RIfe90648_7987);
and \g450883/U$3 ( \28781 , RIfe904e0_7986, \16380 );
nor \g450883/U$1 ( \28782 , \28780 , \28781 );
nand \g447259/U$1 ( \28783 , \28768 , \28776 , \28779 , \28782 );
nor \g445772/U$1 ( \28784 , \28763 , \28764 , \28783 );
and \g450881/U$2 ( \28785 , \16364 , RIfcb8fe8_7127);
and \g450881/U$3 ( \28786 , RIfc4ee90_5920, \16368 );
nor \g450881/U$1 ( \28787 , \28785 , \28786 );
and \g450880/U$2 ( \28788 , \16371 , RIfcb92b8_7129);
and \g450880/U$3 ( \28789 , RIfc86048_6547, \16427 );
nor \g450880/U$1 ( \28790 , \28788 , \28789 );
and \g444980/U$2 ( \28791 , \28784 , \28787 , \28790 );
nor \g444980/U$1 ( \28792 , \28791 , \16480 );
nor \g444714/U$1 ( \28793 , \28762 , \28792 );
and \g446572/U$2 ( \28794 , \19208 , RIdeeb8f8_1144);
and \g446572/U$3 ( \28795 , RIdef99f8_1304, \19210 );
nor \g446572/U$1 ( \28796 , \28794 , \28795 );
and \g446573/U$2 ( \28797 , \19213 , RIdeee5f8_1176);
and \g446573/U$3 ( \28798 , RIdef6cf8_1272, \19215 );
nor \g446573/U$1 ( \28799 , \28797 , \28798 );
and \g446571/U$2 ( \28800 , \19218 , RIdefc6f8_1336);
and \g446571/U$3 ( \28801 , RIdeff3f8_1368, \19220 );
nor \g446571/U$1 ( \28802 , \28800 , \28801 );
nand \g444558/U$1 ( \28803 , \28793 , \28796 , \28799 , \28802 );
and \g445766/U$2 ( \28804 , RIee24dd8_4878, \16319 );
and \g445766/U$3 ( \28805 , RIfc4ff70_5932, \16313 );
and \g448577/U$2 ( \28806 , RIfe91728_7999, \16398 );
and \g448577/U$3 ( \28807 , \16339 , RIdedac60_953);
and \g448577/U$4 ( \28808 , RIdee4170_1059, \16485 );
nor \g448577/U$1 ( \28809 , \28806 , \28807 , \28808 );
and \g454277/U$2 ( \28810 , \16317 , RIee22948_4852);
and \g454277/U$3 ( \28811 , RIfcd4810_7440, \16325 );
nor \g454277/U$1 ( \28812 , \28810 , \28811 );
not \g449603/U$3 ( \28813 , \28812 );
not \g449603/U$4 ( \28814 , \16351 );
and \g449603/U$2 ( \28815 , \28813 , \28814 );
and \g449603/U$5 ( \28816 , \16356 , RIdee5ef8_1080);
nor \g449603/U$1 ( \28817 , \28815 , \28816 );
and \g450857/U$2 ( \28818 , \16361 , RIfe91890_8000);
and \g450857/U$3 ( \28819 , RIded64a8_902, \16364 );
nor \g450857/U$1 ( \28820 , \28818 , \28819 );
and \g450856/U$2 ( \28821 , \16368 , RIee219d0_4841);
and \g450856/U$3 ( \28822 , RIfce1560_7586, \16371 );
nor \g450856/U$1 ( \28823 , \28821 , \28822 );
nand \g447491/U$1 ( \28824 , \28809 , \28817 , \28820 , \28823 );
nor \g445766/U$1 ( \28825 , \28804 , \28805 , \28824 );
and \g450854/U$2 ( \28826 , \16377 , RIfc50240_5934);
and \g450854/U$3 ( \28827 , RIfe915c0_7998, \16380 );
nor \g450854/U$1 ( \28828 , \28826 , \28827 );
and \g450853/U$2 ( \28829 , \16334 , RIdedff58_1012);
and \g450853/U$3 ( \28830 , RIfc857d8_6541, \16328 );
nor \g450853/U$1 ( \28831 , \28829 , \28830 );
and \g444978/U$2 ( \28832 , \28825 , \28828 , \28831 );
nor \g444978/U$1 ( \28833 , \28832 , \16909 );
and \g445768/U$2 ( \28834 , RIdecc728_790, \16313 );
and \g445768/U$3 ( \28835 , RIdedd960_985, \16364 );
and \g448578/U$2 ( \28836 , RIdecf428_822, \16321 );
and \g448578/U$3 ( \28837 , \16485 , RIde9a430_342);
and \g448578/U$4 ( \28838 , RIdeb5f28_534, \16356 );
nor \g448578/U$1 ( \28839 , \28836 , \28837 , \28838 );
and \g450863/U$2 ( \28840 , \16368 , RIdf1ea00_1725);
and \g450863/U$3 ( \28841 , RIdf2e180_1901, \16371 );
nor \g450863/U$1 ( \28842 , \28840 , \28841 );
and \g454217/U$2 ( \28843 , \16317 , RIdf39b20_2033);
and \g454217/U$3 ( \28844 , RIe145128_2163, \16325 );
nor \g454217/U$1 ( \28845 , \28843 , \28844 );
not \g449604/U$3 ( \28846 , \28845 );
not \g449604/U$4 ( \28847 , \16351 );
and \g449604/U$2 ( \28848 , \28846 , \28847 );
and \g449604/U$5 ( \28849 , \16328 , RIded2128_854);
nor \g449604/U$1 ( \28850 , \28848 , \28849 );
and \g450862/U$2 ( \28851 , \16334 , RIe15b928_2419);
and \g450862/U$3 ( \28852 , RIe16fb30_2648, \16380 );
nor \g450862/U$1 ( \28853 , \28851 , \28852 );
nand \g447493/U$1 ( \28854 , \28839 , \28842 , \28850 , \28853 );
nor \g445768/U$1 ( \28855 , \28834 , \28835 , \28854 );
and \g450859/U$2 ( \28856 , \16341 , RIdf020f8_1400);
and \g450859/U$3 ( \28857 , RIdec9a28_758, \16377 );
nor \g450859/U$1 ( \28858 , \28856 , \28857 );
and \g450860/U$2 ( \28859 , \16361 , RIde80378_215);
and \g450860/U$3 ( \28860 , RIdee8bf8_1112, \16398 );
nor \g450860/U$1 ( \28861 , \28859 , \28860 );
and \g444979/U$2 ( \28862 , \28855 , \28858 , \28861 );
nor \g444979/U$1 ( \28863 , \28862 , \16586 );
or \g444315/U$1 ( \28864 , \28742 , \28803 , \28833 , \28863 );
and \g445763/U$2 ( \28865 , RIfc412b8_5767, \16448 );
and \g445763/U$3 ( \28866 , RIdea0d30_374, \16361 );
and \g448573/U$2 ( \28867 , RIdec4028_694, \16321 );
and \g448573/U$3 ( \28868 , \16328 , RIdec6d28_726);
and \g448573/U$4 ( \28869 , RIdead828_438, \16337 );
nor \g448573/U$1 ( \28870 , \28867 , \28868 , \28869 );
and \g454609/U$2 ( \28871 , \16317 , RIdebe628_630);
and \g454609/U$3 ( \28872 , RIfcbaed8_7149, \16325 );
nor \g454609/U$1 ( \28873 , \28871 , \28872 );
not \g449600/U$3 ( \28874 , \28873 );
not \g449600/U$4 ( \28875 , \16330 );
and \g449600/U$2 ( \28876 , \28874 , \28875 );
and \g449600/U$5 ( \28877 , \16341 , RIee1e028_4800);
nor \g449600/U$1 ( \28878 , \28876 , \28877 );
and \g450842/U$2 ( \28879 , \16377 , RIdec1328_662);
and \g450842/U$3 ( \28880 , RIee20bc0_4831, \16313 );
nor \g450842/U$1 ( \28881 , \28879 , \28880 );
and \g450843/U$2 ( \28882 , \16334 , RIdeb8c28_566);
and \g450843/U$3 ( \28883 , RIdebb928_598, \16380 );
nor \g450843/U$1 ( \28884 , \28882 , \28883 );
nand \g447255/U$1 ( \28885 , \28870 , \28878 , \28881 , \28884 );
nor \g445763/U$1 ( \28886 , \28865 , \28866 , \28885 );
and \g450841/U$2 ( \28887 , \16364 , RIdea7630_406);
and \g450841/U$3 ( \28888 , RIdeb0528_470, \16368 );
nor \g450841/U$1 ( \28889 , \28887 , \28888 );
and \g450840/U$2 ( \28890 , \16371 , RIfc9ea08_6827);
and \g450840/U$3 ( \28891 , RIdeb3228_502, \16427 );
nor \g450840/U$1 ( \28892 , \28890 , \28891 );
and \g444976/U$2 ( \28893 , \28886 , \28889 , \28892 );
nor \g444976/U$1 ( \28894 , \28893 , \16618 );
and \g445764/U$2 ( \28895 , RIfe90eb8_7993, \16328 );
and \g445764/U$3 ( \28896 , RIdf3bce0_2057, \16334 );
and \g448575/U$2 ( \28897 , RIee30778_5010, \16427 );
and \g448575/U$3 ( \28898 , \16448 , RIfcec690_7712);
and \g448575/U$4 ( \28899 , RIfe90a80_7990, \16344 );
nor \g448575/U$1 ( \28900 , \28897 , \28898 , \28899 );
and \g454397/U$2 ( \28901 , \16317 , RIdf346c0_1973);
and \g454397/U$3 ( \28902 , RIdf36e20_2001, \16325 );
nor \g454397/U$1 ( \28903 , \28901 , \28902 );
not \g454396/U$1 ( \28904 , \28903 );
and \g449602/U$2 ( \28905 , \28904 , \16336 );
and \g449602/U$3 ( \28906 , RIfe90be8_7991, \16356 );
nor \g449602/U$1 ( \28907 , \28905 , \28906 );
and \g450850/U$2 ( \28908 , \16361 , RIdf30070_1923);
and \g450850/U$3 ( \28909 , RIdf32668_1950, \16364 );
nor \g450850/U$1 ( \28910 , \28908 , \28909 );
and \g450851/U$2 ( \28911 , \16368 , RIee2e5b8_4986);
and \g450851/U$3 ( \28912 , RIfc87dd0_6568, \16371 );
nor \g450851/U$1 ( \28913 , \28911 , \28912 );
nand \g448014/U$1 ( \28914 , \28900 , \28907 , \28910 , \28913 );
nor \g445764/U$1 ( \28915 , \28895 , \28896 , \28914 );
and \g450849/U$2 ( \28916 , \16377 , RIfc9c2a8_6799);
and \g450849/U$3 ( \28917 , RIdf3e008_2082, \16380 );
nor \g450849/U$1 ( \28918 , \28916 , \28917 );
and \g450848/U$2 ( \28919 , \16313 , RIfcb99c0_7134);
and \g450848/U$3 ( \28920 , RIfe90d50_7992, \16321 );
nor \g450848/U$1 ( \28921 , \28919 , \28920 );
and \g444977/U$2 ( \28922 , \28915 , \28918 , \28921 );
nor \g444977/U$1 ( \28923 , \28922 , \16393 );
or \g444267/U$1 ( \28924 , \28864 , \28894 , \28923 );
_DC \g4e2b/U$1 ( \28925 , \28924 , \16652 );
and \g450916/U$2 ( \28926 , \8326 , RIfc5fdf8_6113);
and \g450916/U$3 ( \28927 , RIe176a48_2727, \8404 );
nor \g450916/U$1 ( \28928 , \28926 , \28927 );
and \g445779/U$2 ( \28929 , RIfc72f20_6330, \8373 );
and \g445779/U$3 ( \28930 , RIf16eb48_5719, \8319 );
and \g448596/U$2 ( \28931 , RIf13e8a8_5171, \8414 );
and \g448596/U$3 ( \28932 , \8409 , RIfc61040_6126);
and \g448596/U$4 ( \28933 , RIfe8ff40_7982, \8330 );
nor \g448596/U$1 ( \28934 , \28931 , \28932 , \28933 );
and \g450919/U$2 ( \28935 , \8356 , RIe174e28_2707);
and \g450919/U$3 ( \28936 , RIee3caf0_5149, \8359 );
nor \g450919/U$1 ( \28937 , \28935 , \28936 );
and \g454517/U$2 ( \28938 , \8313 , RIee3a660_5123);
and \g454517/U$3 ( \28939 , RIee3b740_5135, \8323 );
nor \g454517/U$1 ( \28940 , \28938 , \28939 );
not \g449623/U$3 ( \28941 , \28940 );
not \g449623/U$4 ( \28942 , \8347 );
and \g449623/U$2 ( \28943 , \28941 , \28942 );
and \g449623/U$5 ( \28944 , \8351 , RIfe90210_7984);
nor \g449623/U$1 ( \28945 , \28943 , \28944 );
and \g450918/U$2 ( \28946 , \8378 , RIfe900a8_7983);
and \g450918/U$3 ( \28947 , RIfcaf6a0_7018, \8417 );
nor \g450918/U$1 ( \28948 , \28946 , \28947 );
nand \g447503/U$1 ( \28949 , \28934 , \28937 , \28945 , \28948 );
nor \g445779/U$1 ( \28950 , \28929 , \28930 , \28949 );
and \g450917/U$2 ( \28951 , \8335 , RIfcaaab0_6964);
and \g450917/U$3 ( \28952 , RIf170768_5739, \8340 );
nor \g450917/U$1 ( \28953 , \28951 , \28952 );
nand \g445524/U$1 ( \28954 , \28928 , \28950 , \28953 );
and \g444690/U$2 ( \28955 , \28954 , \9700 );
and \g448594/U$2 ( \28956 , RIe1800c0_2834, \8317 );
and \g448594/U$3 ( \28957 , \8326 , RIe182dc0_2866);
and \g448594/U$4 ( \28958 , RIe1887c0_2930, \8488 );
nor \g448594/U$1 ( \28959 , \28956 , \28957 , \28958 );
and \g450914/U$2 ( \28960 , \8335 , RIe17d3c0_2802);
and \g450914/U$3 ( \28961 , RIfe8fc70_7980, \8340 );
nor \g450914/U$1 ( \28962 , \28960 , \28961 );
and \g450912/U$2 ( \28963 , \8404 , RIe1995c0_3122);
and \g450912/U$3 ( \28964 , RIe19efc0_3186, \8351 );
nor \g450912/U$1 ( \28965 , \28963 , \28964 );
and \g454303/U$2 ( \28966 , \8313 , RIf145d60_5254);
and \g454303/U$3 ( \28967 , RIe19c2c0_3154, \8323 );
nor \g454303/U$1 ( \28968 , \28966 , \28967 );
not \g449621/U$3 ( \28969 , \28968 );
not \g449621/U$4 ( \28970 , \8328 );
and \g449621/U$2 ( \28971 , \28969 , \28970 );
and \g449621/U$5 ( \28972 , \8359 , RIe18b4c0_2962);
nor \g449621/U$1 ( \28973 , \28971 , \28972 );
nand \g447502/U$1 ( \28974 , \28959 , \28962 , \28965 , \28973 );
and \g444690/U$3 ( \28975 , \9702 , \28974 );
nor \g444690/U$1 ( \28976 , \28955 , \28975 );
and \g446578/U$2 ( \28977 , \11700 , RIe1968c0_3090);
and \g446578/U$3 ( \28978 , RIfc637a0_6154, \11702 );
nor \g446578/U$1 ( \28979 , \28977 , \28978 );
and \g446577/U$2 ( \28980 , \9230 , RIe185ac0_2898);
and \g446577/U$3 ( \28981 , RIfc62af8_6145, \9232 );
nor \g446577/U$1 ( \28982 , \28980 , \28981 );
and \g446579/U$2 ( \28983 , \9170 , RIe190ec0_3026);
and \g446579/U$3 ( \28984 , RIe193bc0_3058, \9172 );
nor \g446579/U$1 ( \28985 , \28983 , \28984 );
nand \g444457/U$1 ( \28986 , \28976 , \28979 , \28982 , \28985 );
and \g450927/U$2 ( \28987 , \8356 , RIfe8fb08_7979);
and \g450927/U$3 ( \28988 , RIfc5e8e0_6098, \8409 );
nor \g450927/U$1 ( \28989 , \28987 , \28988 );
and \g445782/U$2 ( \28990 , RIf154f40_5426, \8414 );
and \g445782/U$3 ( \28991 , RIfc69e48_6227, \8417 );
and \g448598/U$2 ( \28992 , RIf14e730_5352, \8319 );
and \g448598/U$3 ( \28993 , \8324 , RIfcb1158_7037);
and \g448598/U$4 ( \28994 , RIf1523a8_5395, \8486 );
nor \g448598/U$1 ( \28995 , \28992 , \28993 , \28994 );
and \g450931/U$2 ( \28996 , \8335 , RIe1ef678_4101);
and \g450931/U$3 ( \28997 , RIfcebe20_7706, \8340 );
nor \g450931/U$1 ( \28998 , \28996 , \28997 );
and \g450930/U$2 ( \28999 , \8404 , RIfe8fdd8_7981);
and \g450930/U$3 ( \29000 , RIf159428_5475, \8351 );
nor \g450930/U$1 ( \29001 , \28999 , \29000 );
and \g454896/U$2 ( \29002 , \8313 , RIfc5ebb0_6100);
and \g454896/U$3 ( \29003 , RIf1581e0_5462, \8323 );
nor \g454896/U$1 ( \29004 , \29002 , \29003 );
not \g449625/U$3 ( \29005 , \29004 );
not \g449625/U$4 ( \29006 , \8328 );
and \g449625/U$2 ( \29007 , \29005 , \29006 );
and \g449625/U$5 ( \29008 , \8359 , RIf153b90_5412);
nor \g449625/U$1 ( \29009 , \29007 , \29008 );
nand \g447506/U$1 ( \29010 , \28995 , \28998 , \29001 , \29009 );
nor \g445782/U$1 ( \29011 , \28990 , \28991 , \29010 );
and \g450926/U$2 ( \29012 , \8378 , RIe1f6b30_4184);
and \g450926/U$3 ( \29013 , RIfce88b0_7668, \8531 );
nor \g450926/U$1 ( \29014 , \29012 , \29013 );
nand \g445526/U$1 ( \29015 , \28989 , \29011 , \29014 );
and \g444722/U$2 ( \29016 , \29015 , \8752 );
and \g448597/U$2 ( \29017 , RIe1c5a80_3626, \8326 );
and \g448597/U$3 ( \29018 , \8523 , RIe1ce180_3722);
and \g448597/U$4 ( \29019 , RIe1d0e80_3754, \8486 );
nor \g448597/U$1 ( \29020 , \29017 , \29018 , \29019 );
and \g454211/U$2 ( \29021 , \8313 , RIe1e7680_4010);
and \g454211/U$3 ( \29022 , RIe1ea380_4042, \8323 );
nor \g454211/U$1 ( \29023 , \29021 , \29022 );
not \g449624/U$3 ( \29024 , \29023 );
not \g449624/U$4 ( \29025 , \8328 );
and \g449624/U$2 ( \29026 , \29024 , \29025 );
and \g449624/U$5 ( \29027 , \8340 , RIe1c8780_3658);
nor \g449624/U$1 ( \29028 , \29026 , \29027 );
and \g450923/U$2 ( \29029 , \8404 , RIe1e4980_3978);
and \g450923/U$3 ( \29030 , RIe1ed080_4074, \8351 );
nor \g450923/U$1 ( \29031 , \29029 , \29030 );
and \g450924/U$2 ( \29032 , \8356 , RIe1cb480_3690);
and \g450924/U$3 ( \29033 , RIe1d3b80_3786, \8359 );
nor \g450924/U$1 ( \29034 , \29032 , \29033 );
nand \g447504/U$1 ( \29035 , \29020 , \29028 , \29031 , \29034 );
and \g444722/U$3 ( \29036 , \8478 , \29035 );
nor \g444722/U$1 ( \29037 , \29016 , \29036 );
and \g446580/U$2 ( \29038 , \10534 , RIe1def80_3914);
and \g446580/U$3 ( \29039 , RIe1e1c80_3946, \10536 );
nor \g446580/U$1 ( \29040 , \29038 , \29039 );
and \g446581/U$2 ( \29041 , \10539 , RIe1d9580_3850);
and \g446581/U$3 ( \29042 , RIe1dc280_3882, \10541 );
nor \g446581/U$1 ( \29043 , \29041 , \29042 );
and \g446582/U$2 ( \29044 , \8785 , RIe1c0080_3562);
and \g446582/U$3 ( \29045 , RIe1c2d80_3594, \8787 );
nor \g446582/U$1 ( \29046 , \29044 , \29045 );
nand \g444560/U$1 ( \29047 , \29037 , \29040 , \29043 , \29046 );
and \g445776/U$2 ( \29048 , RIf15d4d8_5521, \8340 );
and \g445776/U$3 ( \29049 , RIfe8f838_7977, \8404 );
and \g448590/U$2 ( \29050 , RIf1638b0_5592, \8412 );
and \g448590/U$3 ( \29051 , \8409 , RIf164990_5604);
and \g448590/U$4 ( \29052 , RIf166718_5625, \8383 );
nor \g448590/U$1 ( \29053 , \29050 , \29051 , \29052 );
and \g454094/U$2 ( \29054 , \8356 , RIe1fc530_4248);
and \g454094/U$3 ( \29055 , RIf161150_5564, \8359 );
nor \g454094/U$1 ( \29056 , \29054 , \29055 );
and \g454296/U$2 ( \29057 , \8313 , RIe1fd778_4261);
and \g454296/U$3 ( \29058 , RIf15f260_5542, \8323 );
nor \g454296/U$1 ( \29059 , \29057 , \29058 );
not \g449618/U$3 ( \29060 , \29059 );
not \g449618/U$4 ( \29061 , \8347 );
and \g449618/U$2 ( \29062 , \29060 , \29061 );
and \g449618/U$5 ( \29063 , \8351 , RIf167690_5636);
nor \g449618/U$1 ( \29064 , \29062 , \29063 );
and \g450904/U$2 ( \29065 , \8378 , RIf1627d0_5580);
and \g450904/U$3 ( \29066 , RIf165638_5613, \8417 );
nor \g450904/U$1 ( \29067 , \29065 , \29066 );
nand \g447499/U$1 ( \29068 , \29053 , \29056 , \29064 , \29067 );
nor \g445776/U$1 ( \29069 , \29048 , \29049 , \29068 );
and \g450901/U$2 ( \29070 , \8335 , RIf159f68_5483);
and \g450901/U$3 ( \29071 , RIfe8f9a0_7978, \8373 );
nor \g450901/U$1 ( \29072 , \29070 , \29071 );
and \g450902/U$2 ( \29073 , \8317 , RIfca20e0_6866);
and \g450902/U$3 ( \29074 , RIf15c290_5508, \8326 );
nor \g450902/U$1 ( \29075 , \29073 , \29074 );
and \g444984/U$2 ( \29076 , \29069 , \29072 , \29075 );
nor \g444984/U$1 ( \29077 , \29076 , \8422 );
and \g445777/U$2 ( \29078 , RIe219f18_4585, \8412 );
and \g445777/U$3 ( \29079 , RIf16b5d8_5681, \8417 );
and \g448592/U$2 ( \29080 , RIe20be18_4425, \8319 );
and \g448592/U$3 ( \29081 , \8326 , RIe20eb18_4457);
and \g448592/U$4 ( \29082 , RIe214518_4521, \8488 );
nor \g448592/U$1 ( \29083 , \29080 , \29081 , \29082 );
and \g450910/U$2 ( \29084 , \8335 , RIe209118_4393);
and \g450910/U$3 ( \29085 , RIfca5a88_6907, \8340 );
nor \g450910/U$1 ( \29086 , \29084 , \29085 );
and \g450909/U$2 ( \29087 , \8404 , RIe222618_4681);
and \g450909/U$3 ( \29088 , RIf16d1f8_5701, \8351 );
nor \g450909/U$1 ( \29089 , \29087 , \29088 );
and \g454851/U$2 ( \29090 , \8313 , RIf16c6b8_5693);
and \g454851/U$3 ( \29091 , RIe225318_4713, \8323 );
nor \g454851/U$1 ( \29092 , \29090 , \29091 );
not \g449619/U$3 ( \29093 , \29092 );
not \g449619/U$4 ( \29094 , \8328 );
and \g449619/U$2 ( \29095 , \29093 , \29094 );
and \g449619/U$5 ( \29096 , \8359 , RIfca62f8_6913);
nor \g449619/U$1 ( \29097 , \29095 , \29096 );
nand \g447500/U$1 ( \29098 , \29083 , \29086 , \29089 , \29097 );
nor \g445777/U$1 ( \29099 , \29078 , \29079 , \29098 );
and \g450905/U$2 ( \29100 , \8378 , RIe217218_4553);
and \g450905/U$3 ( \29101 , RIfcc9578_7313, \8531 );
nor \g450905/U$1 ( \29102 , \29100 , \29101 );
and \g450907/U$2 ( \29103 , \8356 , RIe211818_4489);
and \g450907/U$3 ( \29104 , RIe21f918_4649, \8409 );
nor \g450907/U$1 ( \29105 , \29103 , \29104 );
and \g444985/U$2 ( \29106 , \29099 , \29102 , \29105 );
nor \g444985/U$1 ( \29107 , \29106 , \8368 );
or \g444359/U$1 ( \29108 , \28986 , \29047 , \29077 , \29107 );
and \g445773/U$2 ( \29109 , RIfc483b0_5844, \8340 );
and \g445773/U$3 ( \29110 , RIfeabd08_8271, \8404 );
and \g448587/U$2 ( \29111 , RIe1b3768_3419, \8531 );
and \g448587/U$3 ( \29112 , \8488 , RIf148358_5281);
and \g448587/U$4 ( \29113 , RIfc5d698_6085, \8383 );
nor \g448587/U$1 ( \29114 , \29111 , \29112 , \29113 );
and \g450889/U$2 ( \29115 , \8356 , RIfec3480_8342);
and \g450889/U$3 ( \29116 , RIf149708_5295, \8359 );
nor \g450889/U$1 ( \29117 , \29115 , \29116 );
and \g454294/U$2 ( \29118 , \8313 , RIfec31b0_8340);
and \g454294/U$3 ( \29119 , RIfc5ce28_6079, \8323 );
nor \g454294/U$1 ( \29120 , \29118 , \29119 );
not \g449613/U$3 ( \29121 , \29120 );
not \g449613/U$4 ( \29122 , \8376 );
and \g449613/U$2 ( \29123 , \29121 , \29122 );
and \g449613/U$5 ( \29124 , \8351 , RIfcc8ba0_7306);
nor \g449613/U$1 ( \29125 , \29123 , \29124 );
and \g450888/U$2 ( \29126 , \8378 , RIe1b4b18_3433);
and \g450888/U$3 ( \29127 , RIfc5cf90_6080, \8417 );
nor \g450888/U$1 ( \29128 , \29126 , \29127 );
nand \g447496/U$1 ( \29129 , \29114 , \29117 , \29125 , \29128 );
nor \g445773/U$1 ( \29130 , \29109 , \29110 , \29129 );
and \g450884/U$2 ( \29131 , \8335 , RIfec3318_8341);
and \g450884/U$3 ( \29132 , RIfec35e8_8343, \8373 );
nor \g450884/U$1 ( \29133 , \29131 , \29132 );
and \g450886/U$2 ( \29134 , \8319 , RIe1ad4f8_3349);
and \g450886/U$3 ( \29135 , RIfc80be8_6487, \8326 );
nor \g450886/U$1 ( \29136 , \29134 , \29135 );
and \g444981/U$2 ( \29137 , \29130 , \29133 , \29136 );
nor \g444981/U$1 ( \29138 , \29137 , \8481 );
and \g445775/U$2 ( \29139 , RIe1a49c0_3250, \8373 );
and \g445775/U$3 ( \29140 , RIe172830_2680, \8335 );
and \g448588/U$2 ( \29141 , RIe1f9830_4216, \8531 );
and \g448588/U$3 ( \29142 , \8488 , RIe200478_4293);
and \g448588/U$4 ( \29143 , RIe1a76c0_3282, \8330 );
nor \g448588/U$1 ( \29144 , \29141 , \29142 , \29143 );
and \g450899/U$2 ( \29145 , \8356 , RIe1f2378_4133);
and \g450899/U$3 ( \29146 , RIe206418_4361, \8359 );
nor \g450899/U$1 ( \29147 , \29145 , \29146 );
and \g454855/U$2 ( \29148 , \8313 , RIe228018_4745);
and \g454855/U$3 ( \29149 , RIe17a6c0_2770, \8323 );
nor \g454855/U$1 ( \29150 , \29148 , \29149 );
not \g449614/U$3 ( \29151 , \29150 );
not \g449614/U$4 ( \29152 , \8376 );
and \g449614/U$2 ( \29153 , \29151 , \29152 );
and \g449614/U$5 ( \29154 , \8351 , RIe1aa3c0_3314);
nor \g449614/U$1 ( \29155 , \29153 , \29154 );
and \g450897/U$2 ( \29156 , \8378 , RIe21cc18_4617);
and \g450897/U$3 ( \29157 , RIe18e1c0_2994, \8417 );
nor \g450897/U$1 ( \29158 , \29156 , \29157 );
nand \g447498/U$1 ( \29159 , \29144 , \29147 , \29155 , \29158 );
nor \g445775/U$1 ( \29160 , \29139 , \29140 , \29159 );
and \g450893/U$2 ( \29161 , \8340 , RIe1d6880_3818);
and \g450893/U$3 ( \29162 , RIe1a1cc0_3218, \8404 );
nor \g450893/U$1 ( \29163 , \29161 , \29162 );
and \g450894/U$2 ( \29164 , \8319 , RIe1b01f8_3381);
and \g450894/U$3 ( \29165 , RIe1bd380_3530, \8326 );
nor \g450894/U$1 ( \29166 , \29164 , \29165 );
and \g444983/U$2 ( \29167 , \29160 , \29163 , \29166 );
nor \g444983/U$1 ( \29168 , \29167 , \8651 );
or \g444169/U$1 ( \29169 , \29108 , \29138 , \29168 );
_DC \g4eaf/U$1 ( \29170 , \29169 , \8654 );
and \g451265/U$2 ( \29171 , \16377 , RIee22c18_4854);
and \g451265/U$3 ( \29172 , RIdee0228_1014, \16380 );
nor \g451265/U$1 ( \29173 , \29171 , \29172 );
and \g445856/U$2 ( \29174 , RIee24130_4869, \16321 );
and \g445856/U$3 ( \29175 , RIee235f0_4861, \16313 );
and \g448690/U$2 ( \29176 , RIee21ca0_4843, \16427 );
and \g448690/U$3 ( \29177 , \16432 , RIfc684f8_6209);
and \g448690/U$4 ( \29178 , RIdee1fb0_1035, \16485 );
nor \g448690/U$1 ( \29179 , \29176 , \29177 , \29178 );
and \g454347/U$2 ( \29180 , \16317 , RIfe93ff0_8028);
and \g454347/U$3 ( \29181 , RIded8aa0_929, \16325 );
nor \g454347/U$1 ( \29182 , \29180 , \29181 );
not \g454346/U$1 ( \29183 , \29182 );
and \g449719/U$2 ( \29184 , \29183 , \16336 );
and \g449719/U$3 ( \29185 , RIfe93d20_8026, \16354 );
nor \g449719/U$1 ( \29186 , \29184 , \29185 );
and \g451267/U$2 ( \29187 , \16361 , RIfe93e88_8027);
and \g451267/U$3 ( \29188 , RIded45b8_880, \16364 );
nor \g451267/U$1 ( \29189 , \29187 , \29188 );
and \g451139/U$2 ( \29190 , \16368 , RIee20d28_4832);
and \g451139/U$3 ( \29191 , RIfc68390_6208, \16371 );
nor \g451139/U$1 ( \29192 , \29190 , \29191 );
nand \g448029/U$1 ( \29193 , \29179 , \29186 , \29189 , \29192 );
nor \g445856/U$1 ( \29194 , \29174 , \29175 , \29193 );
and \g451184/U$2 ( \29195 , \16334 , RIdeddc30_987);
and \g451184/U$3 ( \29196 , RIee24f40_4879, \16328 );
nor \g451184/U$1 ( \29197 , \29195 , \29196 );
nand \g445540/U$1 ( \29198 , \29173 , \29194 , \29197 );
and \g444908/U$2 ( \29199 , \29198 , \16477 );
and \g448689/U$2 ( \29200 , RIdf1ecd0_1727, \16398 );
and \g448689/U$3 ( \29201 , \16341 , RIdf20ff8_1752);
and \g448689/U$4 ( \29202 , RIfe931e0_8018, \16485 );
nor \g448689/U$1 ( \29203 , \29200 , \29201 , \29202 );
and \g454403/U$2 ( \29204 , \16317 , RIfca8788_6939);
and \g454403/U$3 ( \29205 , RIfc672b0_6196, \16325 );
nor \g454403/U$1 ( \29206 , \29204 , \29205 );
not \g449717/U$3 ( \29207 , \29206 );
not \g449717/U$4 ( \29208 , \16351 );
and \g449717/U$2 ( \29209 , \29207 , \29208 );
and \g449717/U$5 ( \29210 , \16354 , RIdf29860_1849);
nor \g449717/U$1 ( \29211 , \29209 , \29210 );
and \g451260/U$2 ( \29212 , \16361 , RIfea7c58_8225);
and \g451260/U$3 ( \29213 , RIdf1aab8_1680, \16364 );
nor \g451260/U$1 ( \29214 , \29212 , \29213 );
and \g451259/U$2 ( \29215 , \16368 , RIfcea7a0_7690);
and \g451259/U$3 ( \29216 , RIdf22510_1767, \16371 );
nor \g451259/U$1 ( \29217 , \29215 , \29216 );
nand \g447565/U$1 ( \29218 , \29203 , \29211 , \29214 , \29217 );
and \g444908/U$3 ( \29219 , \16481 , \29218 );
nor \g444908/U$1 ( \29220 , \29199 , \29219 );
and \g446640/U$2 ( \29221 , \16505 , RIee29b30_4933);
and \g446640/U$3 ( \29222 , RIee2b048_4948, \16507 );
nor \g446640/U$1 ( \29223 , \29221 , \29222 );
and \g446642/U$2 ( \29224 , \16511 , RIfe93078_8017);
and \g446642/U$3 ( \29225 , RIfe93348_8019, \16514 );
nor \g446642/U$1 ( \29226 , \29224 , \29225 );
and \g446641/U$2 ( \29227 , \16518 , RIfc6fb18_6293);
and \g446641/U$3 ( \29228 , RIfc67148_6195, \16521 );
nor \g446641/U$1 ( \29229 , \29227 , \29228 );
nand \g444570/U$1 ( \29230 , \29220 , \29223 , \29226 , \29229 );
and \g451277/U$2 ( \29231 , \16377 , RIe15e8f8_2453);
and \g451277/U$3 ( \29232 , RIe1561f8_2357, \16380 );
nor \g451277/U$1 ( \29233 , \29231 , \29232 );
and \g445859/U$2 ( \29234 , RIe1615f8_2485, \16319 );
and \g445859/U$3 ( \29235 , RIee369e8_5080, \16313 );
and \g448693/U$2 ( \29236 , RIe1507f8_2293, \16427 );
and \g448693/U$3 ( \29237 , \16448 , RIfc3ee28_5741);
and \g448693/U$4 ( \29238 , RIe15bbf8_2421, \16485 );
nor \g448693/U$1 ( \29239 , \29236 , \29237 , \29238 );
and \g454445/U$2 ( \29240 , \16317 , RIe14adf8_2229);
and \g454445/U$3 ( \29241 , RIfcca7c0_7326, \16325 );
nor \g454445/U$1 ( \29242 , \29240 , \29241 );
not \g454444/U$1 ( \29243 , \29242 );
and \g449724/U$2 ( \29244 , \29243 , \16336 );
and \g449724/U$3 ( \29245 , RIee35bd8_5070, \16356 );
nor \g449724/U$1 ( \29246 , \29244 , \29245 );
and \g450955/U$2 ( \29247 , \16361 , RIe1453f8_2165);
and \g450955/U$3 ( \29248 , RIe1480f8_2197, \16364 );
nor \g450955/U$1 ( \29249 , \29247 , \29248 );
and \g451279/U$2 ( \29250 , \16368 , RIe14daf8_2261);
and \g451279/U$3 ( \29251 , RIfce6c90_7648, \16371 );
nor \g451279/U$1 ( \29252 , \29250 , \29251 );
nand \g448030/U$1 ( \29253 , \29239 , \29246 , \29249 , \29252 );
nor \g445859/U$1 ( \29254 , \29234 , \29235 , \29253 );
and \g451276/U$2 ( \29255 , \16334 , RIe1534f8_2325);
and \g451276/U$3 ( \29256 , RIe1642f8_2517, \16328 );
nor \g451276/U$1 ( \29257 , \29255 , \29256 );
nand \g445541/U$1 ( \29258 , \29233 , \29254 , \29257 );
and \g444856/U$2 ( \29259 , \29258 , \16390 );
and \g448692/U$2 ( \29260 , RIee32938_5034, \16319 );
and \g448692/U$3 ( \29261 , \16328 , RIee33b80_5047);
and \g448692/U$4 ( \29262 , RIdf32938_1952, \16337 );
nor \g448692/U$1 ( \29263 , \29260 , \29261 , \29262 );
and \g455130/U$2 ( \29264 , \16317 , RIfe93618_8021);
and \g455130/U$3 ( \29265 , RIe1403d0_2108, \16325 );
nor \g455130/U$1 ( \29266 , \29264 , \29265 );
not \g449721/U$3 ( \29267 , \29266 );
not \g449721/U$4 ( \29268 , \16330 );
and \g449721/U$2 ( \29269 , \29267 , \29268 );
and \g449721/U$5 ( \29270 , \16339 , RIfe93bb8_8025);
nor \g449721/U$1 ( \29271 , \29269 , \29270 );
and \g451271/U$2 ( \29272 , \16377 , RIee30bb0_5013);
and \g451271/U$3 ( \29273 , RIee316f0_5021, \16313 );
nor \g451271/U$1 ( \29274 , \29272 , \29273 );
and \g451273/U$2 ( \29275 , \16334 , RIfe934b0_8020);
and \g451273/U$3 ( \29276 , RIdf3bfb0_2059, \16380 );
nor \g451273/U$1 ( \29277 , \29275 , \29276 );
nand \g447274/U$1 ( \29278 , \29263 , \29271 , \29274 , \29277 );
and \g444856/U$3 ( \29279 , \16394 , \29278 );
nor \g444856/U$1 ( \29280 , \29259 , \29279 );
and \g446645/U$2 ( \29281 , \16419 , RIdf2e450_1903);
and \g446645/U$3 ( \29282 , RIdf30340_1925, \16422 );
nor \g446645/U$1 ( \29283 , \29281 , \29282 );
and \g446643/U$2 ( \29284 , \16429 , RIee2ecc0_4991);
and \g446643/U$3 ( \29285 , RIfcd0d00_7398, \16434 );
nor \g446643/U$1 ( \29286 , \29284 , \29285 );
and \g446644/U$2 ( \29287 , \16438 , RIee2cb00_4967);
and \g446644/U$3 ( \29288 , RIee2e720_4987, \16441 );
nor \g446644/U$1 ( \29289 , \29287 , \29288 );
nand \g444571/U$1 ( \29290 , \29280 , \29283 , \29286 , \29289 );
and \g445850/U$2 ( \29291 , RIdec42f8_696, \16328 );
and \g445850/U$3 ( \29292 , RIdeb61f8_536, \16334 );
and \g448685/U$2 ( \29293 , RIdeb07f8_472, \16427 );
and \g448685/U$3 ( \29294 , \16448 , RIee1ea00_4807);
and \g448685/U$4 ( \29295 , RIdebbbf8_600, \16485 );
nor \g448685/U$1 ( \29296 , \29293 , \29294 , \29295 );
and \g454478/U$2 ( \29297 , \16317 , RIdea7cc0_408);
and \g454478/U$3 ( \29298 , RIfc5d3c8_6083, \16325 );
nor \g454478/U$1 ( \29299 , \29297 , \29298 );
not \g454477/U$1 ( \29300 , \29299 );
and \g449714/U$2 ( \29301 , \29300 , \16336 );
and \g449714/U$3 ( \29302 , RIfe93780_8022, \16356 );
nor \g449714/U$1 ( \29303 , \29301 , \29302 );
and \g451249/U$2 ( \29304 , \16361 , RIde9aac0_344);
and \g451249/U$3 ( \29305 , RIdea13c0_376, \16364 );
nor \g451249/U$1 ( \29306 , \29304 , \29305 );
and \g451248/U$2 ( \29307 , \16368 , RIdeadaf8_440);
and \g451248/U$3 ( \29308 , RIee1e2f8_4802, \16371 );
nor \g451248/U$1 ( \29309 , \29307 , \29308 );
nand \g448027/U$1 ( \29310 , \29296 , \29303 , \29306 , \29309 );
nor \g445850/U$1 ( \29311 , \29291 , \29292 , \29310 );
and \g451245/U$2 ( \29312 , \16377 , RIdebe8f8_632);
and \g451245/U$3 ( \29313 , RIdeb8ef8_568, \16380 );
nor \g451245/U$1 ( \29314 , \29312 , \29313 );
and \g451244/U$2 ( \29315 , \16313 , RIfcc6cb0_7284);
and \g451244/U$3 ( \29316 , RIdec15f8_664, \16321 );
nor \g451244/U$1 ( \29317 , \29315 , \29316 );
and \g445040/U$2 ( \29318 , \29311 , \29314 , \29317 );
nor \g445040/U$1 ( \29319 , \29318 , \16618 );
and \g445852/U$2 ( \29320 , RIfcc3b78_7249, \16321 );
and \g445852/U$3 ( \29321 , RIfc7d0d8_6445, \16313 );
and \g448686/U$2 ( \29322 , RIe16ab08_2591, \16398 );
and \g448686/U$3 ( \29323 , \16341 , RIee38a40_5103);
and \g448686/U$4 ( \29324 , RIfe938e8_8023, \16485 );
nor \g448686/U$1 ( \29325 , \29322 , \29323 , \29324 );
and \g454454/U$2 ( \29326 , \16317 , RIfc976b8_6745);
and \g454454/U$3 ( \29327 , RIfc5f420_6106, \16325 );
nor \g454454/U$1 ( \29328 , \29326 , \29327 );
not \g449716/U$3 ( \29329 , \29328 );
not \g449716/U$4 ( \29330 , \16351 );
and \g449716/U$2 ( \29331 , \29329 , \29330 );
and \g449716/U$5 ( \29332 , \16354 , RIfe93a50_8024);
nor \g449716/U$1 ( \29333 , \29331 , \29332 );
and \g451254/U$2 ( \29334 , \16361 , RIe166ff8_2549);
and \g451254/U$3 ( \29335 , RIe169488_2575, \16364 );
nor \g451254/U$1 ( \29336 , \29334 , \29335 );
and \g451253/U$2 ( \29337 , \16368 , RIfc60500_6118);
and \g451253/U$3 ( \29338 , RIfc90a70_6668, \16371 );
nor \g451253/U$1 ( \29339 , \29337 , \29338 );
nand \g447563/U$1 ( \29340 , \29325 , \29333 , \29336 , \29339 );
nor \g445852/U$1 ( \29341 , \29320 , \29321 , \29340 );
and \g451251/U$2 ( \29342 , \16377 , RIfc59750_6040);
and \g451251/U$3 ( \29343 , RIde88370_254, \16380 );
nor \g451251/U$1 ( \29344 , \29342 , \29343 );
and \g451330/U$2 ( \29345 , \16334 , RIde83e88_233);
and \g451330/U$3 ( \29346 , RIfc58238_6025, \16328 );
nor \g451330/U$1 ( \29347 , \29345 , \29346 );
and \g445042/U$2 ( \29348 , \29341 , \29344 , \29347 );
nor \g445042/U$1 ( \29349 , \29348 , \16649 );
or \g444388/U$1 ( \29350 , \29230 , \29290 , \29319 , \29349 );
and \g445847/U$2 ( \29351 , RIdf131c8_1594, \16321 );
and \g445847/U$3 ( \29352 , RIdf104c8_1562, \16313 );
and \g448680/U$2 ( \29353 , RIdef9cc8_1306, \16427 );
and \g448680/U$3 ( \29354 , \16448 , RIdefc9c8_1338);
and \g448680/U$4 ( \29355 , RIdf07dc8_1466, \16485 );
nor \g448680/U$1 ( \29356 , \29353 , \29354 , \29355 );
and \g454546/U$2 ( \29357 , \16317 , RIdeee8c8_1178);
and \g454546/U$3 ( \29358 , RIdef15c8_1210, \16325 );
nor \g454546/U$1 ( \29359 , \29357 , \29358 );
not \g454545/U$1 ( \29360 , \29359 );
and \g449709/U$2 ( \29361 , \29360 , \16336 );
and \g449709/U$3 ( \29362 , RIdf0aac8_1498, \16356 );
nor \g449709/U$1 ( \29363 , \29361 , \29362 );
and \g451233/U$2 ( \29364 , \16361 , RIdee8ec8_1114);
and \g451233/U$3 ( \29365 , RIdeebbc8_1146, \16364 );
nor \g451233/U$1 ( \29366 , \29364 , \29365 );
and \g451232/U$2 ( \29367 , \16368 , RIdef42c8_1242);
and \g451232/U$3 ( \29368 , RIdef6fc8_1274, \16371 );
nor \g451232/U$1 ( \29369 , \29367 , \29368 );
nand \g448026/U$1 ( \29370 , \29356 , \29363 , \29366 , \29369 );
nor \g445847/U$1 ( \29371 , \29351 , \29352 , \29370 );
and \g451229/U$2 ( \29372 , \16377 , RIdf0d7c8_1530);
and \g451229/U$3 ( \29373 , RIdf050c8_1434, \16380 );
nor \g451229/U$1 ( \29374 , \29372 , \29373 );
and \g451228/U$2 ( \29375 , \16334 , RIdf023c8_1402);
and \g451228/U$3 ( \29376 , RIdf15ec8_1626, \16328 );
nor \g451228/U$1 ( \29377 , \29375 , \29376 );
and \g445035/U$2 ( \29378 , \29371 , \29374 , \29377 );
nor \g445035/U$1 ( \29379 , \29378 , \16555 );
and \g445849/U$2 ( \29380 , RIdecf6f8_824, \16328 );
and \g445849/U$3 ( \29381 , RIe158ef8_2389, \16334 );
and \g448681/U$2 ( \29382 , RIdee61c8_1082, \16337 );
and \g448681/U$3 ( \29383 , \16339 , RIdeff6c8_1370);
and \g448681/U$4 ( \29384 , RIde941c0_312, \16485 );
nor \g448681/U$1 ( \29385 , \29382 , \29383 , \29384 );
and \g454501/U$2 ( \29386 , \16317 , RIdf370f0_2003);
and \g454501/U$3 ( \29387 , RIe1426f8_2133, \16325 );
nor \g454501/U$1 ( \29388 , \29386 , \29387 );
not \g449711/U$3 ( \29389 , \29388 );
not \g449711/U$4 ( \29390 , \16351 );
and \g449711/U$2 ( \29391 , \29389 , \29390 );
and \g449711/U$5 ( \29392 , \16354 , RIdeb34f8_504);
nor \g449711/U$1 ( \29393 , \29391 , \29392 );
and \g451242/U$2 ( \29394 , \16361 , RIde7a108_185);
and \g451242/U$3 ( \29395 , RIdedaf30_955, \16364 );
nor \g451242/U$1 ( \29396 , \29394 , \29395 );
and \g451241/U$2 ( \29397 , \16368 , RIdf1bfd0_1695);
and \g451241/U$3 ( \29398 , RIdf2b750_1871, \16371 );
nor \g451241/U$1 ( \29399 , \29397 , \29398 );
nand \g447562/U$1 ( \29400 , \29385 , \29393 , \29396 , \29399 );
nor \g445849/U$1 ( \29401 , \29380 , \29381 , \29400 );
and \g451240/U$2 ( \29402 , \16377 , RIdec6ff8_728);
and \g451240/U$3 ( \29403 , RIe16d100_2618, \16380 );
nor \g451240/U$1 ( \29404 , \29402 , \29403 );
and \g451237/U$2 ( \29405 , \16313 , RIdec9cf8_760);
and \g451237/U$3 ( \29406 , RIdecc9f8_792, \16321 );
nor \g451237/U$1 ( \29407 , \29405 , \29406 );
and \g445037/U$2 ( \29408 , \29401 , \29404 , \29407 );
nor \g445037/U$1 ( \29409 , \29408 , \16586 );
or \g444224/U$1 ( \29410 , \29350 , \29379 , \29409 );
_DC \g4f34/U$1 ( \29411 , \29410 , \16652 );
and \g451308/U$2 ( \29412 , \8523 , RIee39580_5111);
and \g451308/U$3 ( \29413 , RIee3dd38_5162, \8412 );
nor \g451308/U$1 ( \29414 , \29412 , \29413 );
and \g445866/U$2 ( \29415 , RIfc5f6f0_6108, \8409 );
and \g445866/U$3 ( \29416 , RIee3cc58_5150, \8378 );
and \g448705/U$2 ( \29417 , RIe176bb0_2728, \8373 );
and \g448705/U$3 ( \29418 , \8330 , RIf140630_5192);
and \g448705/U$4 ( \29419 , RIee3a7c8_5124, \8488 );
nor \g448705/U$1 ( \29420 , \29417 , \29418 , \29419 );
and \g451312/U$2 ( \29421 , \8335 , RIfc78ec0_6398);
and \g451312/U$3 ( \29422 , RIf16f7f0_5728, \8340 );
nor \g451312/U$1 ( \29423 , \29421 , \29422 );
and \g451311/U$2 ( \29424 , \8404 , RIe1750f8_2709);
and \g451311/U$3 ( \29425 , RIf1419e0_5206, \8351 );
nor \g451311/U$1 ( \29426 , \29424 , \29425 );
and \g454459/U$2 ( \29427 , \8313 , RIf16d900_5706);
and \g454459/U$3 ( \29428 , RIf16ecb0_5720, \8323 );
nor \g454459/U$1 ( \29429 , \29427 , \29428 );
not \g454458/U$1 ( \29430 , \29429 );
and \g449735/U$2 ( \29431 , \29430 , \8316 );
and \g449735/U$3 ( \29432 , RIee3b8a8_5136, \8359 );
nor \g449735/U$1 ( \29433 , \29431 , \29432 );
nand \g448153/U$1 ( \29434 , \29420 , \29423 , \29426 , \29433 );
nor \g445866/U$1 ( \29435 , \29415 , \29416 , \29434 );
and \g451309/U$2 ( \29436 , \8356 , RIfea9008_8239);
and \g451309/U$3 ( \29437 , RIfcd1840_7406, \8417 );
nor \g451309/U$1 ( \29438 , \29436 , \29437 );
nand \g445542/U$1 ( \29439 , \29414 , \29435 , \29438 );
and \g444692/U$2 ( \29440 , \29439 , \9700 );
and \g448702/U$2 ( \29441 , RIe191190_3028, \8412 );
and \g448702/U$3 ( \29442 , \8407 , RIe193e90_3060);
and \g448702/U$4 ( \29443 , RIe199890_3124, \8383 );
nor \g448702/U$1 ( \29444 , \29441 , \29442 , \29443 );
and \g451306/U$2 ( \29445 , \8356 , RIe183090_2868);
and \g451306/U$3 ( \29446 , RIe188a90_2932, \8359 );
nor \g451306/U$1 ( \29447 , \29445 , \29446 );
and \g455211/U$2 ( \29448 , \8313 , RIfccd8f8_7361);
and \g455211/U$3 ( \29449 , RIe185d90_2900, \8323 );
nor \g455211/U$1 ( \29450 , \29448 , \29449 );
not \g449516/U$3 ( \29451 , \29450 );
not \g449516/U$4 ( \29452 , \8347 );
and \g449516/U$2 ( \29453 , \29451 , \29452 );
and \g449516/U$5 ( \29454 , \8351 , RIe19c590_3156);
nor \g449516/U$1 ( \29455 , \29453 , \29454 );
and \g450559/U$2 ( \29456 , \8378 , RIe18e490_2996);
and \g450559/U$3 ( \29457 , RIfc76058_6365, \8417 );
nor \g450559/U$1 ( \29458 , \29456 , \29457 );
nand \g447571/U$1 ( \29459 , \29444 , \29447 , \29455 , \29458 );
and \g444692/U$3 ( \29460 , \9702 , \29459 );
nor \g444692/U$1 ( \29461 , \29440 , \29460 );
and \g446655/U$2 ( \29462 , \9724 , RIe196b90_3092);
and \g446655/U$3 ( \29463 , RIf144f50_5244, \9726 );
nor \g446655/U$1 ( \29464 , \29462 , \29463 );
and \g446652/U$2 ( \29465 , \9729 , RIe17a990_2772);
and \g446652/U$3 ( \29466 , RIe17d690_2804, \9731 );
nor \g446652/U$1 ( \29467 , \29465 , \29466 );
and \g446651/U$2 ( \29468 , \9734 , RIe180390_2836);
and \g446651/U$3 ( \29469 , RIfc76e68_6375, \9736 );
nor \g446651/U$1 ( \29470 , \29468 , \29469 );
nand \g444467/U$1 ( \29471 , \29461 , \29464 , \29467 , \29470 );
and \g451319/U$2 ( \29472 , \8356 , RIe1c8a50_3660);
and \g451319/U$3 ( \29473 , RIe1dc550_3884, \8409 );
nor \g451319/U$1 ( \29474 , \29472 , \29473 );
and \g445868/U$2 ( \29475 , RIe1d9850_3852, \8414 );
and \g445868/U$3 ( \29476 , RIe1df250_3916, \8417 );
and \g448709/U$2 ( \29477 , RIe1e4c50_3980, \8373 );
and \g448709/U$3 ( \29478 , \8330 , RIe1e7950_4012);
and \g448709/U$4 ( \29479 , RIe1ce450_3724, \8486 );
nor \g448709/U$1 ( \29480 , \29477 , \29478 , \29479 );
and \g451321/U$2 ( \29481 , \8335 , RIe1bd650_3532);
and \g451321/U$3 ( \29482 , RIe1c5d50_3628, \8340 );
nor \g451321/U$1 ( \29483 , \29481 , \29482 );
and \g453597/U$2 ( \29484 , \8404 , RIe1e1f50_3948);
and \g453597/U$3 ( \29485 , RIe1ea650_4044, \8351 );
nor \g453597/U$1 ( \29486 , \29484 , \29485 );
and \g454250/U$2 ( \29487 , \8313 , RIe1c0350_3564);
and \g454250/U$3 ( \29488 , RIe1c3050_3596, \8323 );
nor \g454250/U$1 ( \29489 , \29487 , \29488 );
not \g454249/U$1 ( \29490 , \29489 );
and \g449739/U$2 ( \29491 , \29490 , \8316 );
and \g449739/U$3 ( \29492 , RIe1d1150_3756, \8359 );
nor \g449739/U$1 ( \29493 , \29491 , \29492 );
nand \g448154/U$1 ( \29494 , \29480 , \29483 , \29486 , \29493 );
nor \g445868/U$1 ( \29495 , \29475 , \29476 , \29494 );
and \g453645/U$2 ( \29496 , \8378 , RIe1d6b50_3820);
and \g453645/U$3 ( \29497 , RIe1cb750_3692, \8531 );
nor \g453645/U$1 ( \29498 , \29496 , \29497 );
nand \g445545/U$1 ( \29499 , \29474 , \29495 , \29498 );
and \g444762/U$2 ( \29500 , \29499 , \8478 );
and \g448707/U$2 ( \29501 , RIfe91cc8_8003, \8414 );
and \g448707/U$3 ( \29502 , \8409 , RIfce16c8_7587);
and \g448707/U$4 ( \29503 , RIfc9d220_6810, \8330 );
nor \g448707/U$1 ( \29504 , \29501 , \29502 , \29503 );
and \g451316/U$2 ( \29505 , \8356 , RIfe91b60_8002);
and \g451316/U$3 ( \29506 , RIf1484c0_5282, \8359 );
nor \g451316/U$1 ( \29507 , \29505 , \29506 );
and \g454470/U$2 ( \29508 , \8313 , RIfe91f98_8005);
and \g454470/U$3 ( \29509 , RIf147548_5271, \8323 );
nor \g454470/U$1 ( \29510 , \29508 , \29509 );
not \g449736/U$3 ( \29511 , \29510 );
not \g449736/U$4 ( \29512 , \8347 );
and \g449736/U$2 ( \29513 , \29511 , \29512 );
and \g449736/U$5 ( \29514 , \8351 , RIfcda4e0_7506);
nor \g449736/U$1 ( \29515 , \29513 , \29514 );
and \g451315/U$2 ( \29516 , \8378 , RIfe91e30_8004);
and \g451315/U$3 ( \29517 , RIfc4f2c8_5923, \8417 );
nor \g451315/U$1 ( \29518 , \29516 , \29517 );
nand \g447573/U$1 ( \29519 , \29504 , \29507 , \29515 , \29518 );
and \g444762/U$3 ( \29520 , \8482 , \29519 );
nor \g444762/U$1 ( \29521 , \29500 , \29520 );
and \g446659/U$2 ( \29522 , \8509 , RIfe919f8_8001);
and \g446659/U$3 ( \29523 , RIfe92100_8006, \8511 );
nor \g446659/U$1 ( \29524 , \29522 , \29523 );
and \g446658/U$2 ( \29525 , \8514 , RIfc9f548_6835);
and \g446658/U$3 ( \29526 , RIf146b70_5264, \8517 );
nor \g446658/U$1 ( \29527 , \29525 , \29526 );
and \g446660/U$2 ( \29528 , \8969 , RIe1b6738_3453);
and \g446660/U$3 ( \29529 , RIe1b8628_3475, \8971 );
nor \g446660/U$1 ( \29530 , \29528 , \29529 );
nand \g444468/U$1 ( \29531 , \29521 , \29524 , \29527 , \29530 );
and \g445863/U$2 ( \29532 , RIe21cee8_4619, \8407 );
and \g445863/U$3 ( \29533 , RIe2147e8_4523, \8378 );
and \g448699/U$2 ( \29534 , RIfc5a3f8_6049, \8373 );
and \g448699/U$3 ( \29535 , \8330 , RIe2228e8_4683);
and \g448699/U$4 ( \29536 , RIe211ae8_4491, \8486 );
nor \g448699/U$1 ( \29537 , \29534 , \29535 , \29536 );
and \g451300/U$2 ( \29538 , \8335 , RIe2066e8_4363);
and \g451300/U$3 ( \29539 , RIfcc24f8_7233, \8340 );
nor \g451300/U$1 ( \29540 , \29538 , \29539 );
and \g451298/U$2 ( \29541 , \8404 , RIe21fbe8_4651);
and \g451298/U$3 ( \29542 , RIfcc8060_7298, \8351 );
nor \g451298/U$1 ( \29543 , \29541 , \29542 );
and \g454482/U$2 ( \29544 , \8313 , RIe2093e8_4395);
and \g454482/U$3 ( \29545 , RIe20c0e8_4427, \8323 );
nor \g454482/U$1 ( \29546 , \29544 , \29545 );
not \g454481/U$1 ( \29547 , \29546 );
and \g449729/U$2 ( \29548 , \29547 , \8316 );
and \g449729/U$3 ( \29549 , RIfca2c20_6874, \8359 );
nor \g449729/U$1 ( \29550 , \29548 , \29549 );
nand \g448152/U$1 ( \29551 , \29537 , \29540 , \29543 , \29550 );
nor \g445863/U$1 ( \29552 , \29532 , \29533 , \29551 );
and \g451295/U$2 ( \29553 , \8356 , RIe20ede8_4459);
and \g451295/U$3 ( \29554 , RIfc74000_6342, \8417 );
nor \g451295/U$1 ( \29555 , \29553 , \29554 );
and \g451294/U$2 ( \29556 , \8531 , RIfca2950_6872);
and \g451294/U$3 ( \29557 , RIe2174e8_4555, \8414 );
nor \g451294/U$1 ( \29558 , \29556 , \29557 );
and \g445050/U$2 ( \29559 , \29552 , \29555 , \29558 );
nor \g445050/U$1 ( \29560 , \29559 , \8368 );
and \g445865/U$2 ( \29561 , RIfe92f10_8016, \8373 );
and \g445865/U$3 ( \29562 , RIfe92538_8009, \8319 );
and \g448701/U$2 ( \29563 , RIfe92808_8011, \8523 );
and \g448701/U$3 ( \29564 , \8488 , RIf15d640_5522);
and \g448701/U$4 ( \29565 , RIfcc6f80_7286, \8330 );
nor \g448701/U$1 ( \29566 , \29563 , \29564 , \29565 );
and \g450612/U$2 ( \29567 , \8356 , RIfe92c40_8014);
and \g450612/U$3 ( \29568 , RIf15f3c8_5543, \8359 );
nor \g450612/U$1 ( \29569 , \29567 , \29568 );
and \g454452/U$2 ( \29570 , \8313 , RIf162aa0_5582);
and \g454452/U$3 ( \29571 , RIf163a18_5593, \8323 );
nor \g454452/U$1 ( \29572 , \29570 , \29571 );
not \g449733/U$3 ( \29573 , \29572 );
not \g449733/U$4 ( \29574 , \8376 );
and \g449733/U$2 ( \29575 , \29573 , \29574 );
and \g449733/U$5 ( \29576 , \8351 , RIfc45110_5808);
nor \g449733/U$1 ( \29577 , \29575 , \29576 );
and \g451305/U$2 ( \29578 , \8378 , RIfe92ad8_8013);
and \g451305/U$3 ( \29579 , RIf164af8_5605, \8417 );
nor \g451305/U$1 ( \29580 , \29578 , \29579 );
nand \g447570/U$1 ( \29581 , \29566 , \29569 , \29577 , \29580 );
nor \g445865/U$1 ( \29582 , \29561 , \29562 , \29581 );
and \g451303/U$2 ( \29583 , \8335 , RIfcb5a78_7089);
and \g451303/U$3 ( \29584 , RIfe926a0_8010, \8340 );
nor \g451303/U$1 ( \29585 , \29583 , \29584 );
and \g451302/U$2 ( \29586 , \8326 , RIfe92da8_8015);
and \g451302/U$3 ( \29587 , RIfe92970_8012, \8404 );
nor \g451302/U$1 ( \29588 , \29586 , \29587 );
and \g445051/U$2 ( \29589 , \29582 , \29585 , \29588 );
nor \g445051/U$1 ( \29590 , \29589 , \8422 );
or \g444361/U$1 ( \29591 , \29471 , \29531 , \29560 , \29590 );
and \g445861/U$2 ( \29592 , RIfc53be8_5975, \8373 );
and \g445861/U$3 ( \29593 , RIfe92268_8007, \8335 );
and \g448695/U$2 ( \29594 , RIf14ff18_5369, \8531 );
and \g448695/U$3 ( \29595 , \8488 , RIfec3750_8344);
and \g448695/U$4 ( \29596 , RIf157100_5450, \8383 );
nor \g448695/U$1 ( \29597 , \29594 , \29595 , \29596 );
and \g451286/U$2 ( \29598 , \8356 , RIfe923d0_8008);
and \g451286/U$3 ( \29599 , RIf152678_5397, \8359 );
nor \g451286/U$1 ( \29600 , \29598 , \29599 );
and \g454833/U$2 ( \29601 , \8313 , RIf153cf8_5413);
and \g454833/U$3 ( \29602 , RIf1550a8_5427, \8323 );
nor \g454833/U$1 ( \29603 , \29601 , \29602 );
not \g449725/U$3 ( \29604 , \29603 );
not \g449725/U$4 ( \29605 , \8376 );
and \g449725/U$2 ( \29606 , \29604 , \29605 );
and \g449725/U$5 ( \29607 , \8351 , RIf158348_5463);
nor \g449725/U$1 ( \29608 , \29606 , \29607 );
and \g451285/U$2 ( \29609 , \8378 , RIfec3a20_8346);
and \g451285/U$3 ( \29610 , RIfcc5ea0_7274, \8417 );
nor \g451285/U$1 ( \29611 , \29609 , \29610 );
nand \g447567/U$1 ( \29612 , \29597 , \29600 , \29608 , \29611 );
nor \g445861/U$1 ( \29613 , \29592 , \29593 , \29612 );
and \g451282/U$2 ( \29614 , \8340 , RIf14efa0_5358);
and \g451282/U$3 ( \29615 , RIfec38b8_8345, \8404 );
nor \g451282/U$1 ( \29616 , \29614 , \29615 );
and \g451283/U$2 ( \29617 , \8319 , RIf14d380_5338);
and \g451283/U$3 ( \29618 , RIf14e898_5353, \8324 );
nor \g451283/U$1 ( \29619 , \29617 , \29618 );
and \g445047/U$2 ( \29620 , \29613 , \29616 , \29619 );
nor \g445047/U$1 ( \29621 , \29620 , \8621 );
and \g445862/U$2 ( \29622 , RIe177c90_2740, \8409 );
and \g445862/U$3 ( \29623 , RIe21a1e8_4587, \8378 );
and \g448696/U$2 ( \29624 , RIe1ad7c8_3351, \8319 );
and \g448696/U$3 ( \29625 , \8326 , RIe1ba950_3500);
and \g448696/U$4 ( \29626 , RIe1fda48_4263, \8488 );
nor \g448696/U$1 ( \29627 , \29624 , \29625 , \29626 );
and \g451292/U$2 ( \29628 , \8335 , RIe16fe00_2650);
and \g451292/U$3 ( \29629 , RIe1d3e50_3788, \8340 );
nor \g451292/U$1 ( \29630 , \29628 , \29629 );
and \g451291/U$2 ( \29631 , \8404 , RIe19f290_3188);
and \g451291/U$3 ( \29632 , RIe1a7990_3284, \8351 );
nor \g451291/U$1 ( \29633 , \29631 , \29632 );
and \g454284/U$2 ( \29634 , \8313 , RIe1a1f90_3220);
and \g454284/U$3 ( \29635 , RIe1a4c90_3252, \8323 );
nor \g454284/U$1 ( \29636 , \29634 , \29635 );
not \g449727/U$3 ( \29637 , \29636 );
not \g449727/U$4 ( \29638 , \8328 );
and \g449727/U$2 ( \29639 , \29637 , \29638 );
and \g449727/U$5 ( \29640 , \8359 , RIe2039e8_4331);
nor \g449727/U$1 ( \29641 , \29639 , \29640 );
nand \g447569/U$1 ( \29642 , \29627 , \29630 , \29633 , \29641 );
nor \g445862/U$1 ( \29643 , \29622 , \29623 , \29642 );
and \g450827/U$2 ( \29644 , \8356 , RIe1ef948_4103);
and \g450827/U$3 ( \29645 , RIe18b790_2964, \8417 );
nor \g450827/U$1 ( \29646 , \29644 , \29645 );
and \g451288/U$2 ( \29647 , \8531 , RIe1f6e00_4186);
and \g451288/U$3 ( \29648 , RIe2255e8_4715, \8412 );
nor \g451288/U$1 ( \29649 , \29647 , \29648 );
and \g445048/U$2 ( \29650 , \29643 , \29646 , \29649 );
nor \g445048/U$1 ( \29651 , \29650 , \8651 );
or \g444186/U$1 ( \29652 , \29591 , \29621 , \29651 );
_DC \g4fb8/U$1 ( \29653 , \29652 , \8654 );
and \g451353/U$2 ( \29654 , \16377 , RIe15ea60_2454);
and \g451353/U$3 ( \29655 , RIe156360_2358, \16380 );
nor \g451353/U$1 ( \29656 , \29654 , \29655 );
and \g445877/U$2 ( \29657 , RIe161760_2486, \16321 );
and \g445877/U$3 ( \29658 , RIfe942c0_8030, \16313 );
and \g448721/U$2 ( \29659 , RIe150960_2294, \16427 );
and \g448721/U$3 ( \29660 , \16448 , RIfe94428_8031);
and \g448721/U$4 ( \29661 , RIe15bd60_2422, \16485 );
nor \g448721/U$1 ( \29662 , \29659 , \29660 , \29661 );
and \g454199/U$2 ( \29663 , \16317 , RIe14af60_2230);
and \g454199/U$3 ( \29664 , RIfc5c2e8_6071, \16325 );
nor \g454199/U$1 ( \29665 , \29663 , \29664 );
not \g454198/U$1 ( \29666 , \29665 );
and \g449751/U$2 ( \29667 , \29666 , \16336 );
and \g449751/U$3 ( \29668 , RIfe94158_8029, \16356 );
nor \g449751/U$1 ( \29669 , \29667 , \29668 );
and \g451357/U$2 ( \29670 , \16361 , RIe145560_2166);
and \g451357/U$3 ( \29671 , RIe148260_2198, \16364 );
nor \g451357/U$1 ( \29672 , \29670 , \29671 );
and \g451356/U$2 ( \29673 , \16368 , RIe14dc60_2262);
and \g451356/U$3 ( \29674 , RIfe94590_8032, \16371 );
nor \g451356/U$1 ( \29675 , \29673 , \29674 );
nand \g448034/U$1 ( \29676 , \29662 , \29669 , \29672 , \29675 );
nor \g445877/U$1 ( \29677 , \29657 , \29658 , \29676 );
and \g452633/U$2 ( \29678 , \16334 , RIe153660_2326);
and \g452633/U$3 ( \29679 , RIe164460_2518, \16328 );
nor \g452633/U$1 ( \29680 , \29678 , \29679 );
nand \g445546/U$1 ( \29681 , \29656 , \29677 , \29680 );
and \g444739/U$2 ( \29682 , \29681 , \16390 );
and \g448719/U$2 ( \29683 , RIfe95508_8043, \16319 );
and \g448719/U$3 ( \29684 , \16328 , RIfe957d8_8045);
and \g448719/U$4 ( \29685 , RIfe95c10_8048, \16337 );
nor \g448719/U$1 ( \29686 , \29683 , \29684 , \29685 );
and \g454479/U$2 ( \29687 , \16317 , RIfe95238_8041);
and \g454479/U$3 ( \29688 , RIfe95aa8_8047, \16325 );
nor \g454479/U$1 ( \29689 , \29687 , \29688 );
not \g449749/U$3 ( \29690 , \29689 );
not \g449749/U$4 ( \29691 , \16330 );
and \g449749/U$2 ( \29692 , \29690 , \29691 );
and \g449749/U$5 ( \29693 , \16341 , RIee38ba8_5104);
nor \g449749/U$1 ( \29694 , \29692 , \29693 );
and \g451348/U$2 ( \29695 , \16377 , RIee1a7e8_4760);
and \g451348/U$3 ( \29696 , RIfe95670_8044, \16313 );
nor \g451348/U$1 ( \29697 , \29695 , \29696 );
and \g451350/U$2 ( \29698 , \16334 , RIfe953a0_8042);
and \g451350/U$3 ( \29699 , RIfe95940_8046, \16380 );
nor \g451350/U$1 ( \29700 , \29698 , \29699 );
nand \g447282/U$1 ( \29701 , \29686 , \29694 , \29697 , \29700 );
and \g444739/U$3 ( \29702 , \17998 , \29701 );
nor \g444739/U$1 ( \29703 , \29682 , \29702 );
and \g446668/U$2 ( \29704 , \18523 , RIee19438_4746);
and \g446668/U$3 ( \29705 , RIee1a0e0_4755, \18525 );
nor \g446668/U$1 ( \29706 , \29704 , \29705 );
and \g446667/U$2 ( \29707 , \18528 , RIee19870_4749);
and \g446667/U$3 ( \29708 , RIee19ca8_4752, \18530 );
nor \g446667/U$1 ( \29709 , \29707 , \29708 );
and \g446670/U$2 ( \29710 , \18533 , RIfea9440_8242);
and \g446670/U$3 ( \29711 , RIee384a0_5099, \18535 );
nor \g446670/U$1 ( \29712 , \29710 , \29711 );
nand \g444575/U$1 ( \29713 , \29703 , \29706 , \29709 , \29712 );
and \g451365/U$2 ( \29714 , \16313 , RIfcb2940_7054);
and \g451365/U$3 ( \29715 , RIfe946f8_8033, \16321 );
nor \g451365/U$1 ( \29716 , \29714 , \29715 );
and \g445879/U$2 ( \29717 , RIee2b1b0_4949, \16328 );
and \g445879/U$3 ( \29718 , RIfe94860_8034, \16334 );
and \g448724/U$2 ( \29719 , RIee269f8_4898, \16427 );
and \g448724/U$3 ( \29720 , \16432 , RIee26f98_4902);
and \g448724/U$4 ( \29721 , RIdf27538_1824, \16485 );
nor \g448724/U$1 ( \29722 , \29719 , \29720 , \29721 );
and \g454490/U$2 ( \29723 , \16317 , RIfe94c98_8037);
and \g454490/U$3 ( \29724 , RIee26188_4892, \16325 );
nor \g454490/U$1 ( \29725 , \29723 , \29724 );
not \g454489/U$1 ( \29726 , \29725 );
and \g449755/U$2 ( \29727 , \29726 , \16336 );
and \g449755/U$3 ( \29728 , RIfe949c8_8035, \16356 );
nor \g449755/U$1 ( \29729 , \29727 , \29728 );
and \g451370/U$2 ( \29730 , \16361 , RIfea9170_8240);
and \g451370/U$3 ( \29731 , RIee25d50_4889, \16364 );
nor \g451370/U$1 ( \29732 , \29730 , \29731 );
and \g451369/U$2 ( \29733 , \16368 , RIee26458_4894);
and \g451369/U$3 ( \29734 , RIee26728_4896, \16371 );
nor \g451369/U$1 ( \29735 , \29733 , \29734 );
nand \g448036/U$1 ( \29736 , \29722 , \29729 , \29732 , \29735 );
nor \g445879/U$1 ( \29737 , \29717 , \29718 , \29736 );
and \g451366/U$2 ( \29738 , \16377 , RIee273d0_4905);
and \g451366/U$3 ( \29739 , RIfe94b30_8036, \16380 );
nor \g451366/U$1 ( \29740 , \29738 , \29739 );
nand \g445548/U$1 ( \29741 , \29716 , \29737 , \29740 );
and \g444824/U$2 ( \29742 , \29741 , \16481 );
and \g448722/U$2 ( \29743 , RIdef9e30_1307, \16427 );
and \g448722/U$3 ( \29744 , \16448 , RIdefcb30_1339);
and \g448722/U$4 ( \29745 , RIdf07f30_1467, \16344 );
nor \g448722/U$1 ( \29746 , \29743 , \29744 , \29745 );
and \g454321/U$2 ( \29747 , \16317 , RIdeeea30_1179);
and \g454321/U$3 ( \29748 , RIdef1730_1211, \16325 );
nor \g454321/U$1 ( \29749 , \29747 , \29748 );
not \g454320/U$1 ( \29750 , \29749 );
and \g449753/U$2 ( \29751 , \29750 , \16336 );
and \g449753/U$3 ( \29752 , RIdf0ac30_1499, \16356 );
nor \g449753/U$1 ( \29753 , \29751 , \29752 );
and \g451362/U$2 ( \29754 , \16361 , RIdee9030_1115);
and \g451362/U$3 ( \29755 , RIdeebd30_1147, \16364 );
nor \g451362/U$1 ( \29756 , \29754 , \29755 );
and \g451361/U$2 ( \29757 , \16368 , RIdef4430_1243);
and \g451361/U$3 ( \29758 , RIdef7130_1275, \16371 );
nor \g451361/U$1 ( \29759 , \29757 , \29758 );
nand \g448035/U$1 ( \29760 , \29746 , \29753 , \29756 , \29759 );
and \g444824/U$3 ( \29761 , \16750 , \29760 );
nor \g444824/U$1 ( \29762 , \29742 , \29761 );
and \g446671/U$2 ( \29763 , \19457 , RIdf13330_1595);
and \g446671/U$3 ( \29764 , RIdf16030_1627, \19459 );
nor \g446671/U$1 ( \29765 , \29763 , \29764 );
and \g446673/U$2 ( \29766 , \19462 , RIdf02530_1403);
and \g446673/U$3 ( \29767 , RIdf05230_1435, \19464 );
nor \g446673/U$1 ( \29768 , \29766 , \29767 );
and \g446672/U$2 ( \29769 , \19467 , RIdf0d930_1531);
and \g446672/U$3 ( \29770 , RIdf10630_1563, \19469 );
nor \g446672/U$1 ( \29771 , \29769 , \29770 );
nand \g444576/U$1 ( \29772 , \29762 , \29765 , \29768 , \29771 );
and \g445873/U$2 ( \29773 , RIe142860_2134, \16448 );
and \g445873/U$3 ( \29774 , RIdf2b8b8_1872, \16371 );
and \g448715/U$2 ( \29775 , RIdeccb60_793, \16321 );
and \g448715/U$3 ( \29776 , \16328 , RIdecf860_825);
and \g448715/U$4 ( \29777 , RIdee6330_1083, \16398 );
nor \g448715/U$1 ( \29778 , \29775 , \29776 , \29777 );
and \g454830/U$2 ( \29779 , \16317 , RIde94508_313);
and \g454830/U$3 ( \29780 , RIdeb3660_505, \16325 );
nor \g454830/U$1 ( \29781 , \29779 , \29780 );
not \g449744/U$3 ( \29782 , \29781 );
not \g449744/U$4 ( \29783 , \16330 );
and \g449744/U$2 ( \29784 , \29782 , \29783 );
and \g449744/U$5 ( \29785 , \16341 , RIdeff830_1371);
nor \g449744/U$1 ( \29786 , \29784 , \29785 );
and \g451341/U$2 ( \29787 , \16377 , RIdec7160_729);
and \g451341/U$3 ( \29788 , RIdec9e60_761, \16313 );
nor \g451341/U$1 ( \29789 , \29787 , \29788 );
and \g452989/U$2 ( \29790 , \16334 , RIe159060_2390);
and \g452989/U$3 ( \29791 , RIe16d268_2619, \16380 );
nor \g452989/U$1 ( \29792 , \29790 , \29791 );
nand \g447280/U$1 ( \29793 , \29778 , \29786 , \29789 , \29792 );
nor \g445873/U$1 ( \29794 , \29773 , \29774 , \29793 );
and \g451338/U$2 ( \29795 , \16364 , RIdedb098_956);
and \g451338/U$3 ( \29796 , RIdf1c138_1696, \16368 );
nor \g451338/U$1 ( \29797 , \29795 , \29796 );
and \g451339/U$2 ( \29798 , \16361 , RIde7a450_186);
and \g451339/U$3 ( \29799 , RIdf37258_2004, \16427 );
nor \g451339/U$1 ( \29800 , \29798 , \29799 );
and \g445056/U$2 ( \29801 , \29794 , \29797 , \29800 );
nor \g445056/U$1 ( \29802 , \29801 , \16586 );
and \g445875/U$2 ( \29803 , RIee21e08_4844, \16427 );
and \g445875/U$3 ( \29804 , RIfc5dad0_6088, \16368 );
and \g448718/U$2 ( \29805 , RIfe94f68_8039, \16485 );
and \g448718/U$3 ( \29806 , \16356 , RIfe950d0_8040);
and \g448718/U$4 ( \29807 , RIfe96048_8051, \16337 );
nor \g448718/U$1 ( \29808 , \29805 , \29806 , \29807 );
and \g455003/U$2 ( \29809 , \16317 , RIee24298_4870);
and \g455003/U$3 ( \29810 , RIee250a8_4880, \16325 );
nor \g455003/U$1 ( \29811 , \29809 , \29810 );
not \g449746/U$3 ( \29812 , \29811 );
not \g449746/U$4 ( \29813 , \16311 );
and \g449746/U$2 ( \29814 , \29812 , \29813 );
and \g449746/U$5 ( \29815 , \16341 , RIfeaa250_8252);
nor \g449746/U$1 ( \29816 , \29814 , \29815 );
and \g452882/U$2 ( \29817 , \16377 , RIee22d80_4855);
and \g452882/U$3 ( \29818 , RIee23758_4862, \16313 );
nor \g452882/U$1 ( \29819 , \29817 , \29818 );
and \g451347/U$2 ( \29820 , \16334 , RIdeddd98_988);
and \g451347/U$3 ( \29821 , RIfe94e00_8038, \16380 );
nor \g451347/U$1 ( \29822 , \29820 , \29821 );
nand \g447281/U$1 ( \29823 , \29808 , \29816 , \29819 , \29822 );
nor \g445875/U$1 ( \29824 , \29803 , \29804 , \29823 );
and \g451345/U$2 ( \29825 , \16361 , RIfe95ee0_8050);
and \g451345/U$3 ( \29826 , RIee22ab0_4853, \16448 );
nor \g451345/U$1 ( \29827 , \29825 , \29826 );
and \g453002/U$2 ( \29828 , \16364 , RIfe95d78_8049);
and \g453002/U$3 ( \29829 , RIfca46d8_6893, \16371 );
nor \g453002/U$1 ( \29830 , \29828 , \29829 );
and \g445057/U$2 ( \29831 , \29824 , \29827 , \29830 );
nor \g445057/U$1 ( \29832 , \29831 , \16909 );
or \g444316/U$1 ( \29833 , \29713 , \29772 , \29802 , \29832 );
and \g445870/U$2 ( \29834 , RIee33ce8_5048, \16326 );
and \g445870/U$3 ( \29835 , RIdf39df0_2035, \16334 );
and \g448711/U$2 ( \29836 , RIee2ee28_4992, \16427 );
and \g448711/U$3 ( \29837 , \16448 , RIfcdd780_7542);
and \g448711/U$4 ( \29838 , RIdf3e2d8_2084, \16485 );
nor \g448711/U$1 ( \29839 , \29836 , \29837 , \29838 );
and \g454466/U$2 ( \29840 , \16317 , RIdf32aa0_1953);
and \g454466/U$3 ( \29841 , RIdf34990_1975, \16325 );
nor \g454466/U$1 ( \29842 , \29840 , \29841 );
not \g454465/U$1 ( \29843 , \29842 );
and \g449740/U$2 ( \29844 , \29843 , \16336 );
and \g449740/U$3 ( \29845 , RIe140538_2109, \16354 );
nor \g449740/U$1 ( \29846 , \29844 , \29845 );
and \g451329/U$2 ( \29847 , \16361 , RIdf2e5b8_1904);
and \g451329/U$3 ( \29848 , RIdf304a8_1926, \16364 );
nor \g451329/U$1 ( \29849 , \29847 , \29848 );
and \g451327/U$2 ( \29850 , \16368 , RIee2cc68_4968);
and \g451327/U$3 ( \29851 , RIfcc88d0_7304, \16371 );
nor \g451327/U$1 ( \29852 , \29850 , \29851 );
nand \g448033/U$1 ( \29853 , \29839 , \29846 , \29849 , \29852 );
nor \g445870/U$1 ( \29854 , \29834 , \29835 , \29853 );
and \g451325/U$2 ( \29855 , \16377 , RIfc5d530_6084);
and \g451325/U$3 ( \29856 , RIdf3c118_2060, \16380 );
nor \g451325/U$1 ( \29857 , \29855 , \29856 );
and \g451324/U$2 ( \29858 , \16313 , RIee31858_5022);
and \g451324/U$3 ( \29859 , RIee32aa0_5035, \16321 );
nor \g451324/U$1 ( \29860 , \29858 , \29859 );
and \g445052/U$2 ( \29861 , \29854 , \29857 , \29860 );
nor \g445052/U$1 ( \29862 , \29861 , \16393 );
and \g445871/U$2 ( \29863 , RIee1eb68_4808, \16448 );
and \g445871/U$3 ( \29864 , RIde9ae08_345, \16361 );
and \g448713/U$2 ( \29865 , RIdebbd60_601, \16485 );
and \g448713/U$3 ( \29866 , \16356 , RIee1f108_4812);
and \g448713/U$4 ( \29867 , RIdea8008_409, \16337 );
nor \g448713/U$1 ( \29868 , \29865 , \29866 , \29867 );
and \g455293/U$2 ( \29869 , \16317 , RIdec1760_665);
and \g455293/U$3 ( \29870 , RIdec4460_697, \16325 );
nor \g455293/U$1 ( \29871 , \29869 , \29870 );
not \g449742/U$3 ( \29872 , \29871 );
not \g449742/U$4 ( \29873 , \16311 );
and \g449742/U$2 ( \29874 , \29872 , \29873 );
and \g449742/U$5 ( \29875 , \16341 , RIee1d7b8_4794);
nor \g449742/U$1 ( \29876 , \29874 , \29875 );
and \g451337/U$2 ( \29877 , \16377 , RIdebea60_633);
and \g451337/U$3 ( \29878 , RIee1fae0_4819, \16313 );
nor \g451337/U$1 ( \29879 , \29877 , \29878 );
and \g453206/U$2 ( \29880 , \16334 , RIdeb6360_537);
and \g453206/U$3 ( \29881 , RIdeb9060_569, \16380 );
nor \g453206/U$1 ( \29882 , \29880 , \29881 );
nand \g447279/U$1 ( \29883 , \29868 , \29876 , \29879 , \29882 );
nor \g445871/U$1 ( \29884 , \29863 , \29864 , \29883 );
and \g451333/U$2 ( \29885 , \16364 , RIdea1708_377);
and \g451333/U$3 ( \29886 , RIdeadc60_441, \16368 );
nor \g451333/U$1 ( \29887 , \29885 , \29886 );
and \g453332/U$2 ( \29888 , \16371 , RIee1e460_4803);
and \g453332/U$3 ( \29889 , RIdeb0960_473, \16427 );
nor \g453332/U$1 ( \29890 , \29888 , \29889 );
and \g445054/U$2 ( \29891 , \29884 , \29887 , \29890 );
nor \g445054/U$1 ( \29892 , \29891 , \16618 );
or \g444269/U$1 ( \29893 , \29833 , \29862 , \29892 );
_DC \g503d/U$1 ( \29894 , \29893 , \16652 );
and \g451405/U$2 ( \29895 , \8523 , RIfe97290_8064);
and \g451405/U$3 ( \29896 , RIee3dea0_5163, \8414 );
nor \g451405/U$1 ( \29897 , \29895 , \29896 );
and \g445889/U$2 ( \29898 , RIfc48680_5846, \8407 );
and \g445889/U$3 ( \29899 , RIfcc6878_7281, \8378 );
and \g448735/U$2 ( \29900 , RIf16da68_5707, \8319 );
and \g448735/U$3 ( \29901 , \8326 , RIf16ee18_5721);
and \g448735/U$4 ( \29902 , RIee3a930_5125, \8488 );
nor \g448735/U$1 ( \29903 , \29900 , \29901 , \29902 );
and \g451404/U$2 ( \29904 , \8335 , RIf16d360_5702);
and \g451404/U$3 ( \29905 , RIf16f958_5729, \8340 );
nor \g451404/U$1 ( \29906 , \29904 , \29905 );
and \g451403/U$2 ( \29907 , \8404 , RIe175260_2710);
and \g451403/U$3 ( \29908 , RIf141b48_5207, \8351 );
nor \g451403/U$1 ( \29909 , \29907 , \29908 );
and \g454509/U$2 ( \29910 , \8313 , RIfc800a8_6479);
and \g454509/U$3 ( \29911 , RIfc542f0_5980, \8323 );
nor \g454509/U$1 ( \29912 , \29910 , \29911 );
not \g449747/U$3 ( \29913 , \29912 );
not \g449747/U$4 ( \29914 , \8328 );
and \g449747/U$2 ( \29915 , \29913 , \29914 );
and \g449747/U$5 ( \29916 , \8359 , RIee3ba10_5137);
nor \g449747/U$1 ( \29917 , \29915 , \29916 );
nand \g447584/U$1 ( \29918 , \29903 , \29906 , \29909 , \29917 );
nor \g445889/U$1 ( \29919 , \29898 , \29899 , \29918 );
and \g451398/U$2 ( \29920 , \8356 , RIe172b00_2682);
and \g451398/U$3 ( \29921 , RIfca0bc8_6851, \8417 );
nor \g451398/U$1 ( \29922 , \29920 , \29921 );
nand \g445550/U$1 ( \29923 , \29897 , \29919 , \29922 );
and \g444693/U$2 ( \29924 , \29923 , \9700 );
and \g448734/U$2 ( \29925 , RIe1912f8_3029, \8414 );
and \g448734/U$3 ( \29926 , \8407 , RIe193ff8_3061);
and \g448734/U$4 ( \29927 , RIe1999f8_3125, \8383 );
nor \g448734/U$1 ( \29928 , \29925 , \29926 , \29927 );
and \g451469/U$2 ( \29929 , \8356 , RIe1831f8_2869);
and \g451469/U$3 ( \29930 , RIe188bf8_2933, \8359 );
nor \g451469/U$1 ( \29931 , \29929 , \29930 );
and \g454584/U$2 ( \29932 , \8313 , RIfe973f8_8065);
and \g454584/U$3 ( \29933 , RIe185ef8_2901, \8323 );
nor \g454584/U$1 ( \29934 , \29932 , \29933 );
not \g449764/U$3 ( \29935 , \29934 );
not \g449764/U$4 ( \29936 , \8347 );
and \g449764/U$2 ( \29937 , \29935 , \29936 );
and \g449764/U$5 ( \29938 , \8351 , RIe19c6f8_3157);
nor \g449764/U$1 ( \29939 , \29937 , \29938 );
and \g451526/U$2 ( \29940 , \8378 , RIe18e5f8_2997);
and \g451526/U$3 ( \29941 , RIf143fd8_5233, \8417 );
nor \g451526/U$1 ( \29942 , \29940 , \29941 );
nand \g447581/U$1 ( \29943 , \29928 , \29931 , \29939 , \29942 );
and \g444693/U$3 ( \29944 , \9702 , \29943 );
nor \g444693/U$1 ( \29945 , \29924 , \29944 );
and \g446680/U$2 ( \29946 , \9724 , RIe196cf8_3093);
and \g446680/U$3 ( \29947 , RIf1450b8_5245, \9726 );
nor \g446680/U$1 ( \29948 , \29946 , \29947 );
and \g446678/U$2 ( \29949 , \9729 , RIe17aaf8_2773);
and \g446678/U$3 ( \29950 , RIe17d7f8_2805, \9731 );
nor \g446678/U$1 ( \29951 , \29949 , \29950 );
and \g446677/U$2 ( \29952 , \9734 , RIe1804f8_2837);
and \g446677/U$3 ( \29953 , RIf142958_5217, \9736 );
nor \g446677/U$1 ( \29954 , \29952 , \29953 );
nand \g444470/U$1 ( \29955 , \29945 , \29948 , \29951 , \29954 );
and \g451412/U$2 ( \29956 , \8319 , RIf14d4e8_5339);
and \g451412/U$3 ( \29957 , RIfc7f298_6469, \8326 );
nor \g451412/U$1 ( \29958 , \29956 , \29957 );
and \g445892/U$2 ( \29959 , RIf14f108_5359, \8340 );
and \g445892/U$3 ( \29960 , RIfe965e8_8055, \8404 );
and \g448738/U$2 ( \29961 , RIfcd2650_7416, \8531 );
and \g448738/U$3 ( \29962 , \8488 , RIf151430_5384);
and \g448738/U$4 ( \29963 , RIf157268_5451, \8383 );
nor \g448738/U$1 ( \29964 , \29961 , \29962 , \29963 );
and \g451416/U$2 ( \29965 , \8356 , RIe1f2648_4135);
and \g451416/U$3 ( \29966 , RIf1527e0_5398, \8359 );
nor \g451416/U$1 ( \29967 , \29965 , \29966 );
and \g454325/U$2 ( \29968 , \8313 , RIf153e60_5414);
and \g454325/U$3 ( \29969 , RIf155210_5428, \8323 );
nor \g454325/U$1 ( \29970 , \29968 , \29969 );
not \g449769/U$3 ( \29971 , \29970 );
not \g449769/U$4 ( \29972 , \8376 );
and \g449769/U$2 ( \29973 , \29971 , \29972 );
and \g449769/U$5 ( \29974 , \8351 , RIf1584b0_5464);
nor \g449769/U$1 ( \29975 , \29973 , \29974 );
and \g451415/U$2 ( \29976 , \8378 , RIfe96750_8056);
and \g451415/U$3 ( \29977 , RIf155d50_5436, \8417 );
nor \g451415/U$1 ( \29978 , \29976 , \29977 );
nand \g447587/U$1 ( \29979 , \29964 , \29967 , \29975 , \29978 );
nor \g445892/U$1 ( \29980 , \29959 , \29960 , \29979 );
and \g451048/U$2 ( \29981 , \8335 , RIe1ed350_4076);
and \g451048/U$3 ( \29982 , RIf1569f8_5445, \8371 );
nor \g451048/U$1 ( \29983 , \29981 , \29982 );
nand \g445551/U$1 ( \29984 , \29958 , \29980 , \29983 );
and \g444842/U$2 ( \29985 , \29984 , \8752 );
and \g448737/U$2 ( \29986 , RIe1ad930_3352, \8319 );
and \g448737/U$3 ( \29987 , \8324 , RIe1baab8_3501);
and \g448737/U$4 ( \29988 , RIe1fdbb0_4264, \8488 );
nor \g448737/U$1 ( \29989 , \29986 , \29987 , \29988 );
and \g451408/U$2 ( \29990 , \8335 , RIe16ff68_2651);
and \g451408/U$3 ( \29991 , RIe1d3fb8_3789, \8340 );
nor \g451408/U$1 ( \29992 , \29990 , \29991 );
and \g451407/U$2 ( \29993 , \8404 , RIe19f3f8_3189);
and \g451407/U$3 ( \29994 , RIe1a7af8_3285, \8351 );
nor \g451407/U$1 ( \29995 , \29993 , \29994 );
and \g454404/U$2 ( \29996 , \8313 , RIe1a20f8_3221);
and \g454404/U$3 ( \29997 , RIe1a4df8_3253, \8323 );
nor \g454404/U$1 ( \29998 , \29996 , \29997 );
not \g449767/U$3 ( \29999 , \29998 );
not \g449767/U$4 ( \30000 , \8328 );
and \g449767/U$2 ( \30001 , \29999 , \30000 );
and \g449767/U$5 ( \30002 , \8359 , RIe203b50_4332);
nor \g449767/U$1 ( \30003 , \30001 , \30002 );
nand \g447585/U$1 ( \30004 , \29989 , \29992 , \29995 , \30003 );
and \g444842/U$3 ( \30005 , \9010 , \30004 );
nor \g444842/U$1 ( \30006 , \29985 , \30005 );
and \g446684/U$2 ( \30007 , \9031 , RIe21a350_4588);
and \g446684/U$3 ( \30008 , RIe225750_4716, \9033 );
nor \g446684/U$1 ( \30009 , \30007 , \30008 );
and \g446683/U$2 ( \30010 , \9036 , RIe177df8_2741);
and \g446683/U$3 ( \30011 , RIe18b8f8_2965, \9038 );
nor \g446683/U$1 ( \30012 , \30010 , \30011 );
and \g446685/U$2 ( \30013 , \11213 , RIe1efab0_4104);
and \g446685/U$3 ( \30014 , RIe1f6f68_4187, \11215 );
nor \g446685/U$1 ( \30015 , \30013 , \30014 );
nand \g444577/U$1 ( \30016 , \30006 , \30009 , \30012 , \30015 );
and \g445884/U$2 ( \30017 , RIe21d050_4620, \8409 );
and \g445884/U$3 ( \30018 , RIe214950_4524, \8378 );
and \g448731/U$2 ( \30019 , RIe209550_4396, \8319 );
and \g448731/U$3 ( \30020 , \8326 , RIe20c250_4428);
and \g448731/U$4 ( \30021 , RIe211c50_4492, \8488 );
nor \g448731/U$1 ( \30022 , \30019 , \30020 , \30021 );
and \g451389/U$2 ( \30023 , \8335 , RIe206850_4364);
and \g451389/U$3 ( \30024 , RIf1677f8_5637, \8340 );
nor \g451389/U$1 ( \30025 , \30023 , \30024 );
and \g451388/U$2 ( \30026 , \8404 , RIe21fd50_4652);
and \g451388/U$3 ( \30027 , RIfe96e58_8061, \8351 );
nor \g451388/U$1 ( \30028 , \30026 , \30027 );
and \g454659/U$2 ( \30029 , \8313 , RIfe96cf0_8060);
and \g454659/U$3 ( \30030 , RIe222a50_4684, \8323 );
nor \g454659/U$1 ( \30031 , \30029 , \30030 );
not \g449761/U$3 ( \30032 , \30031 );
not \g449761/U$4 ( \30033 , \8328 );
and \g449761/U$2 ( \30034 , \30032 , \30033 );
and \g449761/U$5 ( \30035 , \8359 , RIf169f58_5665);
nor \g449761/U$1 ( \30036 , \30034 , \30035 );
nand \g447578/U$1 ( \30037 , \30022 , \30025 , \30028 , \30036 );
nor \g445884/U$1 ( \30038 , \30017 , \30018 , \30037 );
and \g451385/U$2 ( \30039 , \8356 , RIe20ef50_4460);
and \g451385/U$3 ( \30040 , RIf16a660_5670, \8417 );
nor \g451385/U$1 ( \30041 , \30039 , \30040 );
and \g451384/U$2 ( \30042 , \8531 , RIf168770_5648);
and \g451384/U$3 ( \30043 , RIe217650_4556, \8414 );
nor \g451384/U$1 ( \30044 , \30042 , \30043 );
and \g445062/U$2 ( \30045 , \30038 , \30041 , \30044 );
nor \g445062/U$1 ( \30046 , \30045 , \8368 );
and \g445886/U$2 ( \30047 , RIf162c08_5583, \8414 );
and \g445886/U$3 ( \30048 , RIfe96b88_8059, \8417 );
and \g448732/U$2 ( \30049 , RIfc579c8_6019, \8319 );
and \g448732/U$3 ( \30050 , \8326 , RIfc7cf70_6444);
and \g448732/U$4 ( \30051 , RIf15d7a8_5523, \8486 );
nor \g448732/U$1 ( \30052 , \30049 , \30050 , \30051 );
and \g451649/U$2 ( \30053 , \8335 , RIf159590_5476);
and \g451649/U$3 ( \30054 , RIfcb3fc0_7070, \8340 );
nor \g451649/U$1 ( \30055 , \30053 , \30054 );
and \g451394/U$2 ( \30056 , \8404 , RIe2005e0_4294);
and \g451394/U$3 ( \30057 , RIf166880_5626, \8351 );
nor \g451394/U$1 ( \30058 , \30056 , \30057 );
and \g454504/U$2 ( \30059 , \8313 , RIe201dc8_4311);
and \g454504/U$3 ( \30060 , RIf1657a0_5614, \8323 );
nor \g454504/U$1 ( \30061 , \30059 , \30060 );
not \g449763/U$3 ( \30062 , \30061 );
not \g449763/U$4 ( \30063 , \8328 );
and \g449763/U$2 ( \30064 , \30062 , \30063 );
and \g449763/U$5 ( \30065 , \8359 , RIf15f530_5544);
nor \g449763/U$1 ( \30066 , \30064 , \30065 );
nand \g447580/U$1 ( \30067 , \30052 , \30055 , \30058 , \30066 );
nor \g445886/U$1 ( \30068 , \30047 , \30048 , \30067 );
and \g451391/U$2 ( \30069 , \8378 , RIf161420_5566);
and \g451391/U$3 ( \30070 , RIfe968b8_8057, \8531 );
nor \g451391/U$1 ( \30071 , \30069 , \30070 );
and \g451392/U$2 ( \30072 , \8356 , RIfe96a20_8058);
and \g451392/U$3 ( \30073 , RIf163b80_5594, \8409 );
nor \g451392/U$1 ( \30074 , \30072 , \30073 );
and \g445064/U$2 ( \30075 , \30068 , \30071 , \30074 );
nor \g445064/U$1 ( \30076 , \30075 , \8422 );
or \g444362/U$1 ( \30077 , \29955 , \30016 , \30046 , \30076 );
and \g445881/U$2 ( \30078 , RIe1dc6b8_3885, \8409 );
and \g445881/U$3 ( \30079 , RIe1d6cb8_3821, \8378 );
and \g448726/U$2 ( \30080 , RIe1e4db8_3981, \8373 );
and \g448726/U$3 ( \30081 , \8383 , RIe1e7ab8_4013);
and \g448726/U$4 ( \30082 , RIe1ce5b8_3725, \8488 );
nor \g448726/U$1 ( \30083 , \30080 , \30081 , \30082 );
and \g451375/U$2 ( \30084 , \8335 , RIe1bd7b8_3533);
and \g451375/U$3 ( \30085 , RIe1c5eb8_3629, \8340 );
nor \g451375/U$1 ( \30086 , \30084 , \30085 );
and \g451374/U$2 ( \30087 , \8404 , RIe1e20b8_3949);
and \g451374/U$3 ( \30088 , RIe1ea7b8_4045, \8351 );
nor \g451374/U$1 ( \30089 , \30087 , \30088 );
and \g454702/U$2 ( \30090 , \8313 , RIe1c04b8_3565);
and \g454702/U$3 ( \30091 , RIe1c31b8_3597, \8323 );
nor \g454702/U$1 ( \30092 , \30090 , \30091 );
not \g454701/U$1 ( \30093 , \30092 );
and \g449944/U$2 ( \30094 , \30093 , \8316 );
and \g449944/U$3 ( \30095 , RIe1d12b8_3757, \8359 );
nor \g449944/U$1 ( \30096 , \30094 , \30095 );
nand \g448157/U$1 ( \30097 , \30083 , \30086 , \30089 , \30096 );
nor \g445881/U$1 ( \30098 , \30078 , \30079 , \30097 );
and \g451373/U$2 ( \30099 , \8356 , RIe1c8bb8_3661);
and \g451373/U$3 ( \30100 , RIe1df3b8_3917, \8417 );
nor \g451373/U$1 ( \30101 , \30099 , \30100 );
and \g451372/U$2 ( \30102 , \8523 , RIe1cb8b8_3693);
and \g451372/U$3 ( \30103 , RIe1d99b8_3853, \8414 );
nor \g451372/U$1 ( \30104 , \30102 , \30103 );
and \g445060/U$2 ( \30105 , \30098 , \30101 , \30104 );
nor \g445060/U$1 ( \30106 , \30105 , \8477 );
and \g445883/U$2 ( \30107 , RIf149870_5296, \8409 );
and \g445883/U$3 ( \30108 , RIfe96318_8053, \8378 );
and \g448727/U$2 ( \30109 , RIe1b8790_3476, \8373 );
and \g448727/U$3 ( \30110 , \8383 , RIf14ad88_5311);
and \g448727/U$4 ( \30111 , RIfc58d78_6033, \8486 );
nor \g448727/U$1 ( \30112 , \30109 , \30110 , \30111 );
and \g451383/U$2 ( \30113 , \8335 , RIfe96fc0_8062);
and \g451383/U$3 ( \30114 , RIf146cd8_5265, \8340 );
nor \g451383/U$1 ( \30115 , \30113 , \30114 );
and \g451382/U$2 ( \30116 , \8404 , RIfe96480_8054);
and \g451382/U$3 ( \30117 , RIf14c138_5325, \8351 );
nor \g451382/U$1 ( \30118 , \30116 , \30117 );
and \g454497/U$2 ( \30119 , \8313 , RIfe961b0_8052);
and \g454497/U$3 ( \30120 , RIfc591b0_6036, \8323 );
nor \g454497/U$1 ( \30121 , \30119 , \30120 );
not \g454496/U$1 ( \30122 , \30121 );
and \g449759/U$2 ( \30123 , \30122 , \8316 );
and \g449759/U$3 ( \30124 , RIf148628_5283, \8359 );
nor \g449759/U$1 ( \30125 , \30123 , \30124 );
nand \g448158/U$1 ( \30126 , \30112 , \30115 , \30118 , \30125 );
nor \g445883/U$1 ( \30127 , \30107 , \30108 , \30126 );
and \g451379/U$2 ( \30128 , \8356 , RIe1b04c8_3383);
and \g451379/U$3 ( \30129 , RIf14a0e0_5302, \8417 );
nor \g451379/U$1 ( \30130 , \30128 , \30129 );
and \g451377/U$2 ( \30131 , \8531 , RIe1b20e8_3403);
and \g451377/U$3 ( \30132 , RIfe97128_8063, \8414 );
nor \g451377/U$1 ( \30133 , \30131 , \30132 );
and \g445061/U$2 ( \30134 , \30127 , \30130 , \30133 );
nor \g445061/U$1 ( \30135 , \30134 , \8481 );
or \g444198/U$1 ( \30136 , \30077 , \30106 , \30135 );
_DC \g50c1/U$1 ( \30137 , \30136 , \8654 );
and \g448834/U$2 ( \30138 , RIdf08098_1468, \16485 );
and \g448834/U$3 ( \30139 , \16356 , RIdf0ad98_1500);
and \g448834/U$4 ( \30140 , RIdeeeb98_1180, \16398 );
nor \g448834/U$1 ( \30141 , \30138 , \30139 , \30140 );
and \g454726/U$2 ( \30142 , \16317 , RIdf13498_1596);
and \g454726/U$3 ( \30143 , RIdf16198_1628, \16325 );
nor \g454726/U$1 ( \30144 , \30142 , \30143 );
not \g449859/U$3 ( \30145 , \30144 );
not \g449859/U$4 ( \30146 , \16311 );
and \g449859/U$2 ( \30147 , \30145 , \30146 );
and \g449859/U$5 ( \30148 , \16339 , RIdef1898_1212);
nor \g449859/U$1 ( \30149 , \30147 , \30148 );
and \g452208/U$2 ( \30150 , \16377 , RIdf0da98_1532);
and \g452208/U$3 ( \30151 , RIdf10798_1564, \16313 );
nor \g452208/U$1 ( \30152 , \30150 , \30151 );
and \g451725/U$2 ( \30153 , \16334 , RIdf02698_1404);
and \g451725/U$3 ( \30154 , RIdf05398_1436, \16380 );
nor \g451725/U$1 ( \30155 , \30153 , \30154 );
nand \g447305/U$1 ( \30156 , \30141 , \30149 , \30152 , \30155 );
and \g444715/U$2 ( \30157 , \30156 , \16750 );
and \g445966/U$2 ( \30158 , RIee29c98_4934, \16321 );
and \g445966/U$3 ( \30159 , RIee28780_4919, \16313 );
and \g448835/U$2 ( \30160 , RIdf1ee38_1728, \16337 );
and \g448835/U$3 ( \30161 , \16341 , RIfc83d20_6522);
and \g448835/U$4 ( \30162 , RIdf276a0_1825, \16485 );
nor \g448835/U$1 ( \30163 , \30160 , \30161 , \30162 );
and \g454636/U$2 ( \30164 , \16317 , RIfcb73c8_7107);
and \g454636/U$3 ( \30165 , RIfc83ff0_6524, \16325 );
nor \g454636/U$1 ( \30166 , \30164 , \30165 );
not \g449846/U$3 ( \30167 , \30166 );
not \g449846/U$4 ( \30168 , \16351 );
and \g449846/U$2 ( \30169 , \30167 , \30168 );
and \g449846/U$5 ( \30170 , \16356 , RIdf299c8_1850);
nor \g449846/U$1 ( \30171 , \30169 , \30170 );
and \g451733/U$2 ( \30172 , \16361 , RIdf18a60_1657);
and \g451733/U$3 ( \30173 , RIfc51b90_5952, \16364 );
nor \g451733/U$1 ( \30174 , \30172 , \30173 );
and \g451732/U$2 ( \30175 , \16368 , RIfcdaa80_7510);
and \g451732/U$3 ( \30176 , RIfc51320_5946, \16371 );
nor \g451732/U$1 ( \30177 , \30175 , \30176 );
nand \g447636/U$1 ( \30178 , \30163 , \30171 , \30174 , \30177 );
nor \g445966/U$1 ( \30179 , \30158 , \30159 , \30178 );
and \g451730/U$2 ( \30180 , \16377 , RIee27538_4906);
and \g451730/U$3 ( \30181 , RIdf25918_1804, \16380 );
nor \g451730/U$1 ( \30182 , \30180 , \30181 );
and \g451729/U$2 ( \30183 , \16334 , RIdf23cf8_1784);
and \g451729/U$3 ( \30184 , RIee2b318_4950, \16328 );
nor \g451729/U$1 ( \30185 , \30183 , \30184 );
and \g445123/U$2 ( \30186 , \30179 , \30182 , \30185 );
nor \g445123/U$1 ( \30187 , \30186 , \16480 );
nor \g444715/U$1 ( \30188 , \30157 , \30187 );
and \g446755/U$2 ( \30189 , \19208 , RIdee9198_1116);
and \g446755/U$3 ( \30190 , RIdef7298_1276, \19210 );
nor \g446755/U$1 ( \30191 , \30189 , \30190 );
and \g446756/U$2 ( \30192 , \19213 , RIdeebe98_1148);
and \g446756/U$3 ( \30193 , RIdef4598_1244, \19215 );
nor \g446756/U$1 ( \30194 , \30192 , \30193 );
and \g446754/U$2 ( \30195 , \19218 , RIdef9f98_1308);
and \g446754/U$3 ( \30196 , RIdefcc98_1340, \19220 );
nor \g446754/U$1 ( \30197 , \30195 , \30196 );
nand \g444591/U$1 ( \30198 , \30188 , \30191 , \30194 , \30197 );
and \g451740/U$2 ( \30199 , \16398 , RIdee6498_1084);
and \g451740/U$3 ( \30200 , RIdec72c8_730, \16377 );
nor \g451740/U$1 ( \30201 , \30199 , \30200 );
and \g445968/U$2 ( \30202 , RIdec9fc8_762, \16313 );
and \g445968/U$3 ( \30203 , RIde7a798_187, \16361 );
and \g448839/U$2 ( \30204 , RIdecccc8_794, \16321 );
and \g448839/U$3 ( \30205 , \16485 , RIde94850_314);
and \g448839/U$4 ( \30206 , RIdeb37c8_506, \16356 );
nor \g448839/U$1 ( \30207 , \30204 , \30205 , \30206 );
and \g451743/U$2 ( \30208 , \16368 , RIdf1c2a0_1697);
and \g451743/U$3 ( \30209 , RIdf2ba20_1873, \16371 );
nor \g451743/U$1 ( \30210 , \30208 , \30209 );
and \g455164/U$2 ( \30211 , \16317 , RIdf373c0_2005);
and \g455164/U$3 ( \30212 , RIe1429c8_2135, \16325 );
nor \g455164/U$1 ( \30213 , \30211 , \30212 );
not \g449864/U$3 ( \30214 , \30213 );
not \g449864/U$4 ( \30215 , \16351 );
and \g449864/U$2 ( \30216 , \30214 , \30215 );
and \g449864/U$5 ( \30217 , \16328 , RIdecf9c8_826);
nor \g449864/U$1 ( \30218 , \30216 , \30217 );
and \g450716/U$2 ( \30219 , \16334 , RIe1591c8_2391);
and \g450716/U$3 ( \30220 , RIe16d3d0_2620, \16380 );
nor \g450716/U$1 ( \30221 , \30219 , \30220 );
nand \g447637/U$1 ( \30222 , \30207 , \30210 , \30218 , \30221 );
nor \g445968/U$1 ( \30223 , \30202 , \30203 , \30222 );
and \g451741/U$2 ( \30224 , \16364 , RIdedb200_957);
and \g451741/U$3 ( \30225 , RIdeff998_1372, \16341 );
nor \g451741/U$1 ( \30226 , \30224 , \30225 );
nand \g445571/U$1 ( \30227 , \30201 , \30223 , \30226 );
and \g444889/U$2 ( \30228 , \30227 , \16752 );
and \g448837/U$2 ( \30229 , RIdee2118_1036, \16485 );
and \g448837/U$3 ( \30230 , \16356 , RIfe8cca0_7946);
and \g448837/U$4 ( \30231 , RIded6778_904, \16337 );
nor \g448837/U$1 ( \30232 , \30229 , \30230 , \30231 );
and \g454730/U$2 ( \30233 , \16317 , RIee24400_4871);
and \g454730/U$3 ( \30234 , RIee25210_4881, \16325 );
nor \g454730/U$1 ( \30235 , \30233 , \30234 );
not \g449861/U$3 ( \30236 , \30235 );
not \g449861/U$4 ( \30237 , \16311 );
and \g449861/U$2 ( \30238 , \30236 , \30237 );
and \g449861/U$5 ( \30239 , \16341 , RIded8c08_930);
nor \g449861/U$1 ( \30240 , \30238 , \30239 );
and \g451737/U$2 ( \30241 , \16377 , RIee22ee8_4856);
and \g451737/U$3 ( \30242 , RIee238c0_4863, \16313 );
nor \g451737/U$1 ( \30243 , \30241 , \30242 );
and \g451738/U$2 ( \30244 , \16334 , RIdeddf00_989);
and \g451738/U$3 ( \30245 , RIfe8cb38_7945, \16380 );
nor \g451738/U$1 ( \30246 , \30244 , \30245 );
nand \g447306/U$1 ( \30247 , \30232 , \30240 , \30243 , \30246 );
and \g444889/U$3 ( \30248 , \16477 , \30247 );
nor \g444889/U$1 ( \30249 , \30228 , \30248 );
and \g446758/U$2 ( \30250 , \17463 , RIded23f8_856);
and \g446758/U$3 ( \30251 , RIee21f70_4845, \17465 );
nor \g446758/U$1 ( \30252 , \30250 , \30251 );
and \g446757/U$2 ( \30253 , \17468 , RIded4720_881);
and \g446757/U$3 ( \30254 , RIfcc5a68_7271, \17470 );
nor \g446757/U$1 ( \30255 , \30253 , \30254 );
and \g446759/U$2 ( \30256 , \17473 , RIee20e90_4833);
and \g446759/U$3 ( \30257 , RIfcb6cc0_7102, \17475 );
nor \g446759/U$1 ( \30258 , \30256 , \30257 );
nand \g444592/U$1 ( \30259 , \30249 , \30252 , \30255 , \30258 );
and \g445962/U$2 ( \30260 , RIfc85d78_6545, \16448 );
and \g445962/U$3 ( \30261 , RIde9b150_346, \16361 );
and \g448830/U$2 ( \30262 , RIdec18c8_666, \16321 );
and \g448830/U$3 ( \30263 , \16328 , RIdec45c8_698);
and \g448830/U$4 ( \30264 , RIdea8350_410, \16398 );
nor \g448830/U$1 ( \30265 , \30262 , \30263 , \30264 );
and \g454710/U$2 ( \30266 , \16317 , RIdebbec8_602);
and \g454710/U$3 ( \30267 , RIfcb8bb0_7124, \16325 );
nor \g454710/U$1 ( \30268 , \30266 , \30267 );
not \g450268/U$3 ( \30269 , \30268 );
not \g450268/U$4 ( \30270 , \16330 );
and \g450268/U$2 ( \30271 , \30269 , \30270 );
and \g450268/U$5 ( \30272 , \16341 , RIfc4d3d8_5901);
nor \g450268/U$1 ( \30273 , \30271 , \30272 );
and \g451716/U$2 ( \30274 , \16377 , RIdebebc8_634);
and \g451716/U$3 ( \30275 , RIfce85e0_7666, \16313 );
nor \g451716/U$1 ( \30276 , \30274 , \30275 );
and \g451717/U$2 ( \30277 , \16334 , RIdeb64c8_538);
and \g451717/U$3 ( \30278 , RIdeb91c8_570, \16380 );
nor \g451717/U$1 ( \30279 , \30277 , \30278 );
nand \g447303/U$1 ( \30280 , \30265 , \30273 , \30276 , \30279 );
nor \g445962/U$1 ( \30281 , \30260 , \30261 , \30280 );
and \g451713/U$2 ( \30282 , \16364 , RIdea1a50_378);
and \g451713/U$3 ( \30283 , RIdeaddc8_442, \16368 );
nor \g451713/U$1 ( \30284 , \30282 , \30283 );
and \g453528/U$2 ( \30285 , \16371 , RIfc85aa8_6543);
and \g453528/U$3 ( \30286 , RIdeb0ac8_474, \16427 );
nor \g453528/U$1 ( \30287 , \30285 , \30286 );
and \g445119/U$2 ( \30288 , \30281 , \30284 , \30287 );
nor \g445119/U$1 ( \30289 , \30288 , \16618 );
and \g445963/U$2 ( \30290 , RIee2ef90_4993, \16427 );
and \g445963/U$3 ( \30291 , RIee2cdd0_4969, \16368 );
and \g448831/U$2 ( \30292 , RIfe8ce08_7947, \16344 );
and \g448831/U$3 ( \30293 , \16356 , RIfe8cf70_7948);
and \g448831/U$4 ( \30294 , RIfe8d678_7953, \16398 );
nor \g448831/U$1 ( \30295 , \30292 , \30293 , \30294 );
and \g454908/U$2 ( \30296 , \16317 , RIee32c08_5036);
and \g454908/U$3 ( \30297 , RIee33e50_5049, \16325 );
nor \g454908/U$1 ( \30298 , \30296 , \30297 );
not \g449858/U$3 ( \30299 , \30298 );
not \g449858/U$4 ( \30300 , \16311 );
and \g449858/U$2 ( \30301 , \30299 , \30300 );
and \g449858/U$5 ( \30302 , \16341 , RIdf34af8_1976);
nor \g449858/U$1 ( \30303 , \30301 , \30302 );
and \g451720/U$2 ( \30304 , \16377 , RIee30d18_5014);
and \g451720/U$3 ( \30305 , RIee319c0_5023, \16313 );
nor \g451720/U$1 ( \30306 , \30304 , \30305 );
and \g451721/U$2 ( \30307 , \16334 , RIfe8d0d8_7949);
and \g451721/U$3 ( \30308 , RIfe8d240_7950, \16380 );
nor \g451721/U$1 ( \30309 , \30307 , \30308 );
nand \g447304/U$1 ( \30310 , \30295 , \30303 , \30306 , \30309 );
nor \g445963/U$1 ( \30311 , \30290 , \30291 , \30310 );
and \g451719/U$2 ( \30312 , \16361 , RIdf2e720_1905);
and \g451719/U$3 ( \30313 , RIfce9dc8_7683, \16448 );
nor \g451719/U$1 ( \30314 , \30312 , \30313 );
and \g451718/U$2 ( \30315 , \16364 , RIdf30610_1927);
and \g451718/U$3 ( \30316 , RIfce51d8_7629, \16371 );
nor \g451718/U$1 ( \30317 , \30315 , \30316 );
and \g445120/U$2 ( \30318 , \30311 , \30314 , \30317 );
nor \g445120/U$1 ( \30319 , \30318 , \16393 );
or \g444390/U$1 ( \30320 , \30198 , \30259 , \30289 , \30319 );
and \g445958/U$2 ( \30321 , RIe1618c8_2487, \16321 );
and \g445958/U$3 ( \30322 , RIee36b50_5081, \16313 );
and \g448827/U$2 ( \30323 , RIe14b0c8_2231, \16337 );
and \g448827/U$3 ( \30324 , \16341 , RIfce0fc0_7582);
and \g448827/U$4 ( \30325 , RIe15bec8_2423, \16344 );
nor \g448827/U$1 ( \30326 , \30323 , \30324 , \30325 );
and \g454144/U$2 ( \30327 , \16317 , RIe150ac8_2295);
and \g454144/U$3 ( \30328 , RIfc3ef90_5742, \16325 );
nor \g454144/U$1 ( \30329 , \30327 , \30328 );
not \g449854/U$3 ( \30330 , \30329 );
not \g449854/U$4 ( \30331 , \16351 );
and \g449854/U$2 ( \30332 , \30330 , \30331 );
and \g449854/U$5 ( \30333 , \16354 , RIee35d40_5071);
nor \g449854/U$1 ( \30334 , \30332 , \30333 );
and \g451701/U$2 ( \30335 , \16361 , RIe1456c8_2167);
and \g451701/U$3 ( \30336 , RIe1483c8_2199, \16364 );
nor \g451701/U$1 ( \30337 , \30335 , \30336 );
and \g450681/U$2 ( \30338 , \16368 , RIe14ddc8_2263);
and \g450681/U$3 ( \30339 , RIfe8d7e0_7954, \16371 );
nor \g450681/U$1 ( \30340 , \30338 , \30339 );
nand \g447634/U$1 ( \30341 , \30326 , \30334 , \30337 , \30340 );
nor \g445958/U$1 ( \30342 , \30321 , \30322 , \30341 );
and \g451698/U$2 ( \30343 , \16377 , RIe15ebc8_2455);
and \g451698/U$3 ( \30344 , RIe1564c8_2359, \16380 );
nor \g451698/U$1 ( \30345 , \30343 , \30344 );
and \g451697/U$2 ( \30346 , \16334 , RIe1537c8_2327);
and \g451697/U$3 ( \30347 , RIe1645c8_2519, \16326 );
nor \g451697/U$1 ( \30348 , \30346 , \30347 );
and \g445115/U$2 ( \30349 , \30342 , \30345 , \30348 );
nor \g445115/U$1 ( \30350 , \30349 , \16389 );
and \g445960/U$2 ( \30351 , RIde806c0_216, \16448 );
and \g445960/U$3 ( \30352 , RIe167160_2550, \16361 );
and \g448828/U$2 ( \30353 , RIfe8d3a8_7951, \16485 );
and \g448828/U$3 ( \30354 , \16354 , RIfe8d510_7952);
and \g448828/U$4 ( \30355 , RIe16ac70_2592, \16398 );
nor \g448828/U$1 ( \30356 , \30353 , \30354 , \30355 );
and \g454646/U$2 ( \30357 , \16317 , RIfc9c9b0_6804);
and \g454646/U$3 ( \30358 , RIfc85ee0_6546, \16325 );
nor \g454646/U$1 ( \30359 , \30357 , \30358 );
not \g449855/U$3 ( \30360 , \30359 );
not \g449855/U$4 ( \30361 , \16311 );
and \g449855/U$2 ( \30362 , \30360 , \30361 );
and \g449855/U$5 ( \30363 , \16339 , RIee38d10_5105);
nor \g449855/U$1 ( \30364 , \30362 , \30363 );
and \g451707/U$2 ( \30365 , \16377 , RIfcb8778_7121);
and \g451707/U$3 ( \30366 , RIfce13f8_7585, \16313 );
nor \g451707/U$1 ( \30367 , \30365 , \30366 );
and \g451708/U$2 ( \30368 , \16334 , RIde841d0_234);
and \g451708/U$3 ( \30369 , RIde886b8_255, \16380 );
nor \g451708/U$1 ( \30370 , \30368 , \30369 );
nand \g447301/U$1 ( \30371 , \30356 , \30364 , \30367 , \30370 );
nor \g445960/U$1 ( \30372 , \30351 , \30352 , \30371 );
and \g451705/U$2 ( \30373 , \16364 , RIfc850d0_6536);
and \g451705/U$3 ( \30374 , RIfc9c140_6798, \16368 );
nor \g451705/U$1 ( \30375 , \30373 , \30374 );
and \g451704/U$2 ( \30376 , \16371 , RIfce1128_7583);
and \g451704/U$3 ( \30377 , RIfcb8070_7116, \16427 );
nor \g451704/U$1 ( \30378 , \30376 , \30377 );
and \g445117/U$2 ( \30379 , \30372 , \30375 , \30378 );
nor \g445117/U$1 ( \30380 , \30379 , \16649 );
or \g444210/U$1 ( \30381 , \30320 , \30350 , \30380 );
_DC \g5146/U$1 ( \30382 , \30381 , \16652 );
and \g448848/U$2 ( \30383 , RIee396e8_5112, \8531 );
and \g448848/U$3 ( \30384 , \8486 , RIee3aa98_5126);
and \g448848/U$4 ( \30385 , RIf140798_5193, \8330 );
nor \g448848/U$1 ( \30386 , \30383 , \30384 , \30385 );
and \g451773/U$2 ( \30387 , \8356 , RIe172c68_2683);
and \g451773/U$3 ( \30388 , RIee3bb78_5138, \8359 );
nor \g451773/U$1 ( \30389 , \30387 , \30388 );
and \g454658/U$2 ( \30390 , \8313 , RIee3e008_5164);
and \g454658/U$3 ( \30391 , RIf13eb78_5173, \8323 );
nor \g454658/U$1 ( \30392 , \30390 , \30391 );
not \g449872/U$3 ( \30393 , \30392 );
not \g449872/U$4 ( \30394 , \8376 );
and \g449872/U$2 ( \30395 , \30393 , \30394 );
and \g449872/U$5 ( \30396 , \8351 , RIf141cb0_5208);
nor \g449872/U$1 ( \30397 , \30395 , \30396 );
and \g451772/U$2 ( \30398 , \8378 , RIee3cdc0_5151);
and \g451772/U$3 ( \30399 , RIfceb880_7702, \8417 );
nor \g451772/U$1 ( \30400 , \30398 , \30399 );
nand \g447646/U$1 ( \30401 , \30386 , \30389 , \30397 , \30400 );
and \g444682/U$2 ( \30402 , \30401 , \9700 );
and \g445978/U$2 ( \30403 , RIf142ac0_5218, \8340 );
and \g445978/U$3 ( \30404 , RIe196e60_3094, \8404 );
and \g448849/U$2 ( \30405 , RIf1431c8_5223, \8523 );
and \g448849/U$3 ( \30406 , \8486 , RIe186060_2902);
and \g448849/U$4 ( \30407 , RIe199b60_3126, \8330 );
nor \g448849/U$1 ( \30408 , \30405 , \30406 , \30407 );
and \g453180/U$2 ( \30409 , \8356 , RIe183360_2870);
and \g453180/U$3 ( \30410 , RIe188d60_2934, \8359 );
nor \g453180/U$1 ( \30411 , \30409 , \30410 );
and \g454684/U$2 ( \30412 , \8313 , RIe191460_3030);
and \g454684/U$3 ( \30413 , RIe194160_3062, \8323 );
nor \g454684/U$1 ( \30414 , \30412 , \30413 );
not \g449873/U$3 ( \30415 , \30414 );
not \g449873/U$4 ( \30416 , \8376 );
and \g449873/U$2 ( \30417 , \30415 , \30416 );
and \g449873/U$5 ( \30418 , \8351 , RIe19c860_3158);
nor \g449873/U$1 ( \30419 , \30417 , \30418 );
and \g453179/U$2 ( \30420 , \8378 , RIe18e760_2998);
and \g453179/U$3 ( \30421 , RIf144140_5234, \8417 );
nor \g453179/U$1 ( \30422 , \30420 , \30421 );
nand \g447647/U$1 ( \30423 , \30408 , \30411 , \30419 , \30422 );
nor \g445978/U$1 ( \30424 , \30403 , \30404 , \30423 );
and \g451776/U$2 ( \30425 , \8335 , RIe17ac60_2774);
and \g451776/U$3 ( \30426 , RIf145220_5246, \8373 );
nor \g451776/U$1 ( \30427 , \30425 , \30426 );
and \g451777/U$2 ( \30428 , \8319 , RIe17d960_2806);
and \g451777/U$3 ( \30429 , RIe180660_2838, \8326 );
nor \g451777/U$1 ( \30430 , \30428 , \30429 );
and \g445134/U$2 ( \30431 , \30424 , \30427 , \30430 );
nor \g445134/U$1 ( \30432 , \30431 , \8589 );
nor \g444682/U$1 ( \30433 , \30402 , \30432 );
and \g446760/U$2 ( \30434 , \10034 , RIf16ef80_5722);
and \g446760/U$3 ( \30435 , RIf16fac0_5730, \10036 );
nor \g446760/U$1 ( \30436 , \30434 , \30435 );
and \g446761/U$2 ( \30437 , \10039 , RIfe8be90_7936);
and \g446761/U$3 ( \30438 , RIf13ff28_5187, \10041 );
nor \g446761/U$1 ( \30439 , \30437 , \30438 );
and \g446762/U$2 ( \30440 , \10044 , RIfcc4af0_7260);
and \g446762/U$3 ( \30441 , RIf16dbd0_5708, \10046 );
nor \g446762/U$1 ( \30442 , \30440 , \30441 );
nand \g444480/U$1 ( \30443 , \30433 , \30436 , \30439 , \30442 );
and \g451784/U$2 ( \30444 , \8414 , RIfec1e00_8326);
and \g451784/U$3 ( \30445 , RIfc4ebc0_5918, \8407 );
nor \g451784/U$1 ( \30446 , \30444 , \30445 );
and \g445980/U$2 ( \30447 , RIfcd4db0_7444, \8417 );
and \g445980/U$3 ( \30448 , RIfec1b30_8324, \8356 );
and \g448853/U$2 ( \30449 , RIe1b88f8_3477, \8373 );
and \g448853/U$3 ( \30450 , \8383 , RIf14aef0_5312);
and \g448853/U$4 ( \30451 , RIf1476b0_5272, \8488 );
nor \g448853/U$1 ( \30452 , \30449 , \30450 , \30451 );
and \g451787/U$2 ( \30453 , \8335 , RIfec1c98_8325);
and \g451787/U$3 ( \30454 , RIfc4e788_5915, \8340 );
nor \g451787/U$1 ( \30455 , \30453 , \30454 );
and \g451786/U$2 ( \30456 , \8404 , RIe1b68a0_3454);
and \g451786/U$3 ( \30457 , RIf14c2a0_5326, \8351 );
nor \g451786/U$1 ( \30458 , \30456 , \30457 );
and \g455029/U$2 ( \30459 , \8313 , RIfe8bbc0_7934);
and \g455029/U$3 ( \30460 , RIfcb8e80_7126, \8323 );
nor \g455029/U$1 ( \30461 , \30459 , \30460 );
not \g455028/U$1 ( \30462 , \30461 );
and \g449877/U$2 ( \30463 , \30462 , \8316 );
and \g449877/U$3 ( \30464 , RIf148790_5284, \8359 );
nor \g449877/U$1 ( \30465 , \30463 , \30464 );
nand \g448172/U$1 ( \30466 , \30452 , \30455 , \30458 , \30465 );
nor \g445980/U$1 ( \30467 , \30447 , \30448 , \30466 );
and \g451785/U$2 ( \30468 , \8378 , RIfe8bd28_7935);
and \g451785/U$3 ( \30469 , RIfe8ba58_7933, \8531 );
nor \g451785/U$1 ( \30470 , \30468 , \30469 );
nand \g445572/U$1 ( \30471 , \30446 , \30467 , \30470 );
and \g444901/U$2 ( \30472 , \30471 , \8482 );
and \g448850/U$2 ( \30473 , RIe1e4f20_3982, \8373 );
and \g448850/U$3 ( \30474 , \8383 , RIe1e7c20_4014);
and \g448850/U$4 ( \30475 , RIe1ce720_3726, \8488 );
nor \g448850/U$1 ( \30476 , \30473 , \30474 , \30475 );
and \g451781/U$2 ( \30477 , \8335 , RIe1bd920_3534);
and \g451781/U$3 ( \30478 , RIe1c6020_3630, \8340 );
nor \g451781/U$1 ( \30479 , \30477 , \30478 );
and \g453033/U$2 ( \30480 , \8404 , RIe1e2220_3950);
and \g453033/U$3 ( \30481 , RIe1ea920_4046, \8351 );
nor \g453033/U$1 ( \30482 , \30480 , \30481 );
and \g454942/U$2 ( \30483 , \8313 , RIe1c0620_3566);
and \g454942/U$3 ( \30484 , RIe1c3320_3598, \8323 );
nor \g454942/U$1 ( \30485 , \30483 , \30484 );
not \g454941/U$1 ( \30486 , \30485 );
and \g449875/U$2 ( \30487 , \30486 , \8316 );
and \g449875/U$3 ( \30488 , RIe1d1420_3758, \8359 );
nor \g449875/U$1 ( \30489 , \30487 , \30488 );
nand \g448171/U$1 ( \30490 , \30476 , \30479 , \30482 , \30489 );
and \g444901/U$3 ( \30491 , \8478 , \30490 );
nor \g444901/U$1 ( \30492 , \30472 , \30491 );
and \g446765/U$2 ( \30493 , \10534 , RIe1dc820_3886);
and \g446765/U$3 ( \30494 , RIe1df520_3918, \10536 );
nor \g446765/U$1 ( \30495 , \30493 , \30494 );
and \g446766/U$2 ( \30496 , \10539 , RIe1d6e20_3822);
and \g446766/U$3 ( \30497 , RIe1d9b20_3854, \10541 );
nor \g446766/U$1 ( \30498 , \30496 , \30497 );
and \g446767/U$2 ( \30499 , \8775 , RIe1c8d20_3662);
and \g446767/U$3 ( \30500 , RIe1cba20_3694, \8777 );
nor \g446767/U$1 ( \30501 , \30499 , \30500 );
nand \g444593/U$1 ( \30502 , \30492 , \30495 , \30498 , \30501 );
and \g445974/U$2 ( \30503 , RIf15c3f8_5509, \8340 );
and \g445974/U$3 ( \30504 , RIfe8c700_7942, \8404 );
and \g448843/U$2 ( \30505 , RIfe8c598_7941, \8523 );
and \g448843/U$3 ( \30506 , \8488 , RIf15d910_5524);
and \g448843/U$4 ( \30507 , RIf165908_5615, \8330 );
nor \g448843/U$1 ( \30508 , \30505 , \30506 , \30507 );
and \g451765/U$2 ( \30509 , \8356 , RIfe8c868_7943);
and \g451765/U$3 ( \30510 , RIf15f698_5545, \8359 );
nor \g451765/U$1 ( \30511 , \30509 , \30510 );
and \g455141/U$2 ( \30512 , \8313 , RIf162d70_5584);
and \g455141/U$3 ( \30513 , RIf163ce8_5595, \8323 );
nor \g455141/U$1 ( \30514 , \30512 , \30513 );
not \g450411/U$3 ( \30515 , \30514 );
not \g450411/U$4 ( \30516 , \8376 );
and \g450411/U$2 ( \30517 , \30515 , \30516 );
and \g450411/U$5 ( \30518 , \8351 , RIf1669e8_5627);
nor \g450411/U$1 ( \30519 , \30517 , \30518 );
and \g451764/U$2 ( \30520 , \8378 , RIf161588_5567);
and \g451764/U$3 ( \30521 , RIfc9c578_6801, \8417 );
nor \g451764/U$1 ( \30522 , \30520 , \30521 );
nand \g447643/U$1 ( \30523 , \30508 , \30511 , \30519 , \30522 );
nor \g445974/U$1 ( \30524 , \30503 , \30504 , \30523 );
and \g451761/U$2 ( \30525 , \8335 , RIf1596f8_5477);
and \g451761/U$3 ( \30526 , RIfe8c9d0_7944, \8371 );
nor \g451761/U$1 ( \30527 , \30525 , \30526 );
and \g451762/U$2 ( \30528 , \8319 , RIf15a0d0_5484);
and \g451762/U$3 ( \30529 , RIf15aee0_5494, \8326 );
nor \g451762/U$1 ( \30530 , \30528 , \30529 );
and \g445129/U$2 ( \30531 , \30524 , \30527 , \30530 );
nor \g445129/U$1 ( \30532 , \30531 , \8422 );
and \g445975/U$2 ( \30533 , RIe21d1b8_4621, \8409 );
and \g445975/U$3 ( \30534 , RIe214ab8_4525, \8378 );
and \g448845/U$2 ( \30535 , RIe2096b8_4397, \8319 );
and \g448845/U$3 ( \30536 , \8324 , RIe20c3b8_4429);
and \g448845/U$4 ( \30537 , RIe211db8_4493, \8488 );
nor \g448845/U$1 ( \30538 , \30535 , \30536 , \30537 );
and \g451771/U$2 ( \30539 , \8335 , RIe2069b8_4365);
and \g451771/U$3 ( \30540 , RIf167960_5638, \8340 );
nor \g451771/U$1 ( \30541 , \30539 , \30540 );
and \g453533/U$2 ( \30542 , \8404 , RIe21feb8_4653);
and \g453533/U$3 ( \30543 , RIf16c820_5694, \8351 );
nor \g453533/U$1 ( \30544 , \30542 , \30543 );
and \g455074/U$2 ( \30545 , \8313 , RIf16b740_5682);
and \g455074/U$3 ( \30546 , RIe222bb8_4685, \8323 );
nor \g455074/U$1 ( \30547 , \30545 , \30546 );
not \g449871/U$3 ( \30548 , \30547 );
not \g449871/U$4 ( \30549 , \8328 );
and \g449871/U$2 ( \30550 , \30548 , \30549 );
and \g449871/U$5 ( \30551 , \8359 , RIfe8c430_7940);
nor \g449871/U$1 ( \30552 , \30550 , \30551 );
nand \g447645/U$1 ( \30553 , \30538 , \30541 , \30544 , \30552 );
nor \g445975/U$1 ( \30554 , \30533 , \30534 , \30553 );
and \g451769/U$2 ( \30555 , \8356 , RIe20f0b8_4461);
and \g451769/U$3 ( \30556 , RIf16a7c8_5671, \8417 );
nor \g451769/U$1 ( \30557 , \30555 , \30556 );
and \g453580/U$2 ( \30558 , \8531 , RIf1688d8_5649);
and \g453580/U$3 ( \30559 , RIe2177b8_4557, \8412 );
nor \g453580/U$1 ( \30560 , \30558 , \30559 );
and \g445130/U$2 ( \30561 , \30554 , \30557 , \30560 );
nor \g445130/U$1 ( \30562 , \30561 , \8368 );
or \g444365/U$1 ( \30563 , \30443 , \30502 , \30532 , \30562 );
and \g445971/U$2 ( \30564 , RIe177f60_2742, \8409 );
and \g445971/U$3 ( \30565 , RIe21a4b8_4589, \8378 );
and \g448842/U$2 ( \30566 , RIe1bac20_3502, \8326 );
and \g448842/U$3 ( \30567 , \8531 , RIe1f70d0_4188);
and \g448842/U$4 ( \30568 , RIe1fdd18_4265, \8488 );
nor \g448842/U$1 ( \30569 , \30566 , \30567 , \30568 );
and \g455340/U$2 ( \30570 , \8313 , RIe1a2260_3222);
and \g455340/U$3 ( \30571 , RIe1a4f60_3254, \8323 );
nor \g455340/U$1 ( \30572 , \30570 , \30571 );
not \g449868/U$3 ( \30573 , \30572 );
not \g449868/U$4 ( \30574 , \8328 );
and \g449868/U$2 ( \30575 , \30573 , \30574 );
and \g449868/U$5 ( \30576 , \8340 , RIe1d4120_3790);
nor \g449868/U$1 ( \30577 , \30575 , \30576 );
and \g451755/U$2 ( \30578 , \8404 , RIe19f560_3190);
and \g451755/U$3 ( \30579 , RIe1a7c60_3286, \8351 );
nor \g451755/U$1 ( \30580 , \30578 , \30579 );
and \g451756/U$2 ( \30581 , \8356 , RIe1efc18_4105);
and \g451756/U$3 ( \30582 , RIe203cb8_4333, \8359 );
nor \g451756/U$1 ( \30583 , \30581 , \30582 );
nand \g447641/U$1 ( \30584 , \30569 , \30577 , \30580 , \30583 );
nor \g445971/U$1 ( \30585 , \30564 , \30565 , \30584 );
and \g451754/U$2 ( \30586 , \8335 , RIe1700d0_2652);
and \g451754/U$3 ( \30587 , RIe18ba60_2966, \8417 );
nor \g451754/U$1 ( \30588 , \30586 , \30587 );
and \g451753/U$2 ( \30589 , \8319 , RIe1ada98_3353);
and \g451753/U$3 ( \30590 , RIe2258b8_4717, \8414 );
nor \g451753/U$1 ( \30591 , \30589 , \30590 );
and \g445127/U$2 ( \30592 , \30585 , \30588 , \30591 );
nor \g445127/U$1 ( \30593 , \30592 , \8651 );
and \g445970/U$2 ( \30594 , RIf14f270_5360, \8340 );
and \g445970/U$3 ( \30595 , RIfec1f68_8327, \8404 );
and \g448840/U$2 ( \30596 , RIf153fc8_5415, \8414 );
and \g448840/U$3 ( \30597 , \8409 , RIf155378_5429);
and \g448840/U$4 ( \30598 , RIf1573d0_5452, \8383 );
nor \g448840/U$1 ( \30599 , \30596 , \30597 , \30598 );
and \g451750/U$2 ( \30600 , \8356 , RIfe8c2c8_7939);
and \g451750/U$3 ( \30601 , RIf152948_5399, \8359 );
nor \g451750/U$1 ( \30602 , \30600 , \30601 );
and \g455399/U$2 ( \30603 , \8313 , RIf150080_5370);
and \g455399/U$3 ( \30604 , RIf151598_5385, \8323 );
nor \g455399/U$1 ( \30605 , \30603 , \30604 );
not \g449866/U$3 ( \30606 , \30605 );
not \g449866/U$4 ( \30607 , \8347 );
and \g449866/U$2 ( \30608 , \30606 , \30607 );
and \g449866/U$5 ( \30609 , \8351 , RIf158618_5465);
nor \g449866/U$1 ( \30610 , \30608 , \30609 );
and \g451749/U$2 ( \30611 , \8378 , RIfe8bff8_7937);
and \g451749/U$3 ( \30612 , RIf155eb8_5437, \8417 );
nor \g451749/U$1 ( \30613 , \30611 , \30612 );
nand \g447639/U$1 ( \30614 , \30599 , \30602 , \30610 , \30613 );
nor \g445970/U$1 ( \30615 , \30594 , \30595 , \30614 );
and \g451746/U$2 ( \30616 , \8335 , RIfe8c160_7938);
and \g451746/U$3 ( \30617 , RIf156b60_5446, \8373 );
nor \g451746/U$1 ( \30618 , \30616 , \30617 );
and \g451748/U$2 ( \30619 , \8319 , RIf14d650_5340);
and \g451748/U$3 ( \30620 , RIfc503a8_5935, \8326 );
nor \g451748/U$1 ( \30621 , \30619 , \30620 );
and \g445126/U$2 ( \30622 , \30615 , \30618 , \30621 );
nor \g445126/U$1 ( \30623 , \30622 , \8621 );
or \g444188/U$1 ( \30624 , \30563 , \30593 , \30623 );
_DC \g51ca/U$1 ( \30625 , \30624 , \8654 );
and \g448860/U$2 ( \30626 , RIdeeed00_1181, \16398 );
and \g448860/U$3 ( \30627 , \16341 , RIdef1a00_1213);
and \g448860/U$4 ( \30628 , RIdf08200_1469, \16485 );
nor \g448860/U$1 ( \30629 , \30626 , \30627 , \30628 );
and \g454676/U$2 ( \30630 , \16317 , RIdefa100_1309);
and \g454676/U$3 ( \30631 , RIdefce00_1341, \16325 );
nor \g454676/U$1 ( \30632 , \30630 , \30631 );
not \g449885/U$3 ( \30633 , \30632 );
not \g449885/U$4 ( \30634 , \16351 );
and \g449885/U$2 ( \30635 , \30633 , \30634 );
and \g449885/U$5 ( \30636 , \16356 , RIdf0af00_1501);
nor \g449885/U$1 ( \30637 , \30635 , \30636 );
and \g451814/U$2 ( \30638 , \16361 , RIdee9300_1117);
and \g451814/U$3 ( \30639 , RIdeec000_1149, \16364 );
nor \g451814/U$1 ( \30640 , \30638 , \30639 );
and \g452042/U$2 ( \30641 , \16368 , RIdef4700_1245);
and \g452042/U$3 ( \30642 , RIdef7400_1277, \16371 );
nor \g452042/U$1 ( \30643 , \30641 , \30642 );
nand \g447652/U$1 ( \30644 , \30629 , \30637 , \30640 , \30643 );
and \g444716/U$2 ( \30645 , \30644 , \16750 );
and \g445987/U$2 ( \30646 , RIfcd9f40_7502, \16427 );
and \g445987/U$3 ( \30647 , RIfc54cc8_5987, \16368 );
and \g448861/U$2 ( \30648 , RIdf27808_1826, \16344 );
and \g448861/U$3 ( \30649 , \16356 , RIdf29b30_1851);
and \g448861/U$4 ( \30650 , RIdf1efa0_1729, \16398 );
nor \g448861/U$1 ( \30651 , \30648 , \30649 , \30650 );
and \g454666/U$2 ( \30652 , \16317 , RIfec23a0_8330);
and \g454666/U$3 ( \30653 , RIee2b480_4951, \16325 );
nor \g454666/U$1 ( \30654 , \30652 , \30653 );
not \g449911/U$3 ( \30655 , \30654 );
not \g449911/U$4 ( \30656 , \16311 );
and \g449911/U$2 ( \30657 , \30655 , \30656 );
and \g449911/U$5 ( \30658 , \16339 , RIfc4b218_5877);
nor \g449911/U$1 ( \30659 , \30657 , \30658 );
and \g451896/U$2 ( \30660 , \16377 , RIfec2238_8329);
and \g451896/U$3 ( \30661 , RIee288e8_4920, \16313 );
nor \g451896/U$1 ( \30662 , \30660 , \30661 );
and \g451818/U$2 ( \30663 , \16334 , RIdf23e60_1785);
and \g451818/U$3 ( \30664 , RIdf25a80_1805, \16380 );
nor \g451818/U$1 ( \30665 , \30663 , \30664 );
nand \g447310/U$1 ( \30666 , \30651 , \30659 , \30662 , \30665 );
nor \g445987/U$1 ( \30667 , \30646 , \30647 , \30666 );
and \g451816/U$2 ( \30668 , \16361 , RIdf18bc8_1658);
and \g451816/U$3 ( \30669 , RIfc55100_5990, \16448 );
nor \g451816/U$1 ( \30670 , \30668 , \30669 );
and \g451815/U$2 ( \30671 , \16364 , RIfcc69e0_7282);
and \g451815/U$3 ( \30672 , RIfc54f98_5989, \16371 );
nor \g451815/U$1 ( \30673 , \30671 , \30672 );
and \g445141/U$2 ( \30674 , \30667 , \30670 , \30673 );
nor \g445141/U$1 ( \30675 , \30674 , \16480 );
nor \g444716/U$1 ( \30676 , \30645 , \30675 );
and \g446771/U$2 ( \30677 , \19457 , RIdf13600_1597);
and \g446771/U$3 ( \30678 , RIdf16300_1629, \19459 );
nor \g446771/U$1 ( \30679 , \30677 , \30678 );
and \g446773/U$2 ( \30680 , \19462 , RIdf02800_1405);
and \g446773/U$3 ( \30681 , RIdf05500_1437, \19464 );
nor \g446773/U$1 ( \30682 , \30680 , \30681 );
and \g446772/U$2 ( \30683 , \19467 , RIdf0dc00_1533);
and \g446772/U$3 ( \30684 , RIdf10900_1565, \19469 );
nor \g446772/U$1 ( \30685 , \30683 , \30684 );
nand \g444595/U$1 ( \30686 , \30676 , \30679 , \30682 , \30685 );
and \g451825/U$2 ( \30687 , \16364 , RIdedb368_958);
and \g451825/U$3 ( \30688 , RIdf2bb88_1874, \16371 );
nor \g451825/U$1 ( \30689 , \30687 , \30688 );
and \g445989/U$2 ( \30690 , RIdf37528_2006, \16427 );
and \g445989/U$3 ( \30691 , RIdf1c408_1698, \16368 );
and \g448863/U$2 ( \30692 , RIde94b98_315, \16344 );
and \g448863/U$3 ( \30693 , \16354 , RIdeb3930_507);
and \g448863/U$4 ( \30694 , RIdee6600_1085, \16398 );
nor \g448863/U$1 ( \30695 , \30692 , \30693 , \30694 );
and \g455169/U$2 ( \30696 , \16317 , RIdecce30_795);
and \g455169/U$3 ( \30697 , RIdecfb30_827, \16325 );
nor \g455169/U$1 ( \30698 , \30696 , \30697 );
not \g449889/U$3 ( \30699 , \30698 );
not \g449889/U$4 ( \30700 , \16311 );
and \g449889/U$2 ( \30701 , \30699 , \30700 );
and \g449889/U$5 ( \30702 , \16341 , RIdeffb00_1373);
nor \g449889/U$1 ( \30703 , \30701 , \30702 );
and \g451653/U$2 ( \30704 , \16377 , RIdec7430_731);
and \g451653/U$3 ( \30705 , RIdeca130_763, \16313 );
nor \g451653/U$1 ( \30706 , \30704 , \30705 );
and \g451827/U$2 ( \30707 , \16334 , RIe159330_2392);
and \g451827/U$3 ( \30708 , RIe16d538_2621, \16380 );
nor \g451827/U$1 ( \30709 , \30707 , \30708 );
nand \g447313/U$1 ( \30710 , \30695 , \30703 , \30706 , \30709 );
nor \g445989/U$1 ( \30711 , \30690 , \30691 , \30710 );
and \g451826/U$2 ( \30712 , \16361 , RIde7aae0_188);
and \g451826/U$3 ( \30713 , RIe142b30_2136, \16432 );
nor \g451826/U$1 ( \30714 , \30712 , \30713 );
nand \g445574/U$1 ( \30715 , \30689 , \30711 , \30714 );
and \g444890/U$2 ( \30716 , \30715 , \16752 );
and \g448862/U$2 ( \30717 , RIfc9e8a0_6826, \16321 );
and \g448862/U$3 ( \30718 , \16328 , RIfce4ad0_7624);
and \g448862/U$4 ( \30719 , RIded68e0_905, \16398 );
nor \g448862/U$1 ( \30720 , \30717 , \30718 , \30719 );
and \g455134/U$2 ( \30721 , \16317 , RIdee2280_1037);
and \g455134/U$3 ( \30722 , RIdee4440_1061, \16325 );
nor \g455134/U$1 ( \30723 , \30721 , \30722 );
not \g449863/U$3 ( \30724 , \30723 );
not \g449863/U$4 ( \30725 , \16330 );
and \g449863/U$2 ( \30726 , \30724 , \30725 );
and \g449863/U$5 ( \30727 , \16341 , RIded8d70_931);
nor \g449863/U$1 ( \30728 , \30726 , \30727 );
and \g451820/U$2 ( \30729 , \16377 , RIfcd4108_7435);
and \g451820/U$3 ( \30730 , RIfcc46b8_7257, \16313 );
nor \g451820/U$1 ( \30731 , \30729 , \30730 );
and \g451766/U$2 ( \30732 , \16334 , RIdede068_990);
and \g451766/U$3 ( \30733 , RIdee0390_1015, \16380 );
nor \g451766/U$1 ( \30734 , \30732 , \30733 );
nand \g447312/U$1 ( \30735 , \30720 , \30728 , \30731 , \30734 );
and \g444890/U$3 ( \30736 , \16477 , \30735 );
nor \g444890/U$1 ( \30737 , \30716 , \30736 );
and \g446778/U$2 ( \30738 , \17463 , RIded2560_857);
and \g446778/U$3 ( \30739 , RIfce54a8_7631, \17465 );
nor \g446778/U$1 ( \30740 , \30738 , \30739 );
and \g446777/U$2 ( \30741 , \17468 , RIded4888_882);
and \g446777/U$3 ( \30742 , RIfcda0a8_7503, \17470 );
nor \g446777/U$1 ( \30743 , \30741 , \30742 );
and \g446779/U$2 ( \30744 , \17473 , RIfc50ee8_5943);
and \g446779/U$3 ( \30745 , RIfca0790_6848, \17475 );
nor \g446779/U$1 ( \30746 , \30744 , \30745 );
nand \g444596/U$1 ( \30747 , \30737 , \30740 , \30743 , \30746 );
and \g445985/U$2 ( \30748 , RIdec1a30_667, \16321 );
and \g445985/U$3 ( \30749 , RIfce3f90_7616, \16313 );
and \g449015/U$2 ( \30750 , RIdeb0c30_475, \16427 );
and \g449015/U$3 ( \30751 , \16448 , RIfc8c588_6619);
and \g449015/U$4 ( \30752 , RIdebc030_603, \16485 );
nor \g449015/U$1 ( \30753 , \30750 , \30751 , \30752 );
and \g454341/U$2 ( \30754 , \16317 , RIdea8698_411);
and \g454341/U$3 ( \30755 , RIfc99b48_6771, \16325 );
nor \g454341/U$1 ( \30756 , \30754 , \30755 );
not \g454340/U$1 ( \30757 , \30756 );
and \g449881/U$2 ( \30758 , \30757 , \16336 );
and \g449881/U$3 ( \30759 , RIfcc3308_7243, \16356 );
nor \g449881/U$1 ( \30760 , \30758 , \30759 );
and \g451806/U$2 ( \30761 , \16361 , RIde9b498_347);
and \g451806/U$3 ( \30762 , RIdea1d98_379, \16364 );
nor \g451806/U$1 ( \30763 , \30761 , \30762 );
and \g452343/U$2 ( \30764 , \16368 , RIdeadf30_443);
and \g452343/U$3 ( \30765 , RIfc5a998_6053, \16371 );
nor \g452343/U$1 ( \30766 , \30764 , \30765 );
nand \g448056/U$1 ( \30767 , \30753 , \30760 , \30763 , \30766 );
nor \g445985/U$1 ( \30768 , \30748 , \30749 , \30767 );
and \g451803/U$2 ( \30769 , \16377 , RIdebed30_635);
and \g451803/U$3 ( \30770 , RIdeb9330_571, \16380 );
nor \g451803/U$1 ( \30771 , \30769 , \30770 );
and \g451801/U$2 ( \30772 , \16334 , RIdeb6630_539);
and \g451801/U$3 ( \30773 , RIdec4730_699, \16328 );
nor \g451801/U$1 ( \30774 , \30772 , \30773 );
and \g445138/U$2 ( \30775 , \30768 , \30771 , \30774 );
nor \g445138/U$1 ( \30776 , \30775 , \16618 );
and \g445986/U$2 ( \30777 , RIfc56bb8_6009, \16321 );
and \g445986/U$3 ( \30778 , RIfca1ca8_6863, \16313 );
and \g448858/U$2 ( \30779 , RIee2f0f8_4994, \16427 );
and \g448858/U$3 ( \30780 , \16432 , RIfc9a958_6781);
and \g448858/U$4 ( \30781 , RIdf3e440_2085, \16485 );
nor \g448858/U$1 ( \30782 , \30779 , \30780 , \30781 );
and \g454722/U$2 ( \30783 , \16317 , RIfec2940_8334);
and \g454722/U$3 ( \30784 , RIdf34c60_1977, \16325 );
nor \g454722/U$1 ( \30785 , \30783 , \30784 );
not \g454721/U$1 ( \30786 , \30785 );
and \g449883/U$2 ( \30787 , \30786 , \16336 );
and \g449883/U$3 ( \30788 , RIe1406a0_2110, \16356 );
nor \g449883/U$1 ( \30789 , \30787 , \30788 );
and \g451811/U$2 ( \30790 , \16361 , RIdf2e888_1906);
and \g451811/U$3 ( \30791 , RIdf30778_1928, \16364 );
nor \g451811/U$1 ( \30792 , \30790 , \30791 );
and \g451810/U$2 ( \30793 , \16368 , RIee2cf38_4970);
and \g451810/U$3 ( \30794 , RIfcdb458_7517, \16371 );
nor \g451810/U$1 ( \30795 , \30793 , \30794 );
nand \g448057/U$1 ( \30796 , \30782 , \30789 , \30792 , \30795 );
nor \g445986/U$1 ( \30797 , \30777 , \30778 , \30796 );
and \g451809/U$2 ( \30798 , \16377 , RIfcec960_7714);
and \g451809/U$3 ( \30799 , RIdf3c280_2061, \16380 );
nor \g451809/U$1 ( \30800 , \30798 , \30799 );
and \g451808/U$2 ( \30801 , \16334 , RIdf39f58_2036);
and \g451808/U$3 ( \30802 , RIfc9aac0_6782, \16328 );
nor \g451808/U$1 ( \30803 , \30801 , \30802 );
and \g445140/U$2 ( \30804 , \30797 , \30800 , \30803 );
nor \g445140/U$1 ( \30805 , \30804 , \16393 );
or \g444391/U$1 ( \30806 , \30686 , \30747 , \30776 , \30805 );
and \g445982/U$2 ( \30807 , RIe161a30_2488, \16321 );
and \g445982/U$3 ( \30808 , RIee36cb8_5082, \16313 );
and \g448855/U$2 ( \30809 , RIe150c30_2296, \16427 );
and \g448855/U$3 ( \30810 , \16448 , RIfcc7688_7291);
and \g448855/U$4 ( \30811 , RIe15c030_2424, \16485 );
nor \g448855/U$1 ( \30812 , \30809 , \30810 , \30811 );
and \g455387/U$2 ( \30813 , \16317 , RIe14b230_2232);
and \g455387/U$3 ( \30814 , RIfc9a250_6776, \16325 );
nor \g455387/U$1 ( \30815 , \30813 , \30814 );
not \g455386/U$1 ( \30816 , \30815 );
and \g449878/U$2 ( \30817 , \30816 , \16336 );
and \g449878/U$3 ( \30818 , RIfcc7250_7288, \16354 );
nor \g449878/U$1 ( \30819 , \30817 , \30818 );
and \g451792/U$2 ( \30820 , \16361 , RIe145830_2168);
and \g451792/U$3 ( \30821 , RIe148530_2200, \16364 );
nor \g451792/U$1 ( \30822 , \30820 , \30821 );
and \g452689/U$2 ( \30823 , \16368 , RIe14df30_2264);
and \g452689/U$3 ( \30824 , RIfc8af08_6603, \16371 );
nor \g452689/U$1 ( \30825 , \30823 , \30824 );
nand \g448054/U$1 ( \30826 , \30812 , \30819 , \30822 , \30825 );
nor \g445982/U$1 ( \30827 , \30807 , \30808 , \30826 );
and \g451790/U$2 ( \30828 , \16377 , RIe15ed30_2456);
and \g451790/U$3 ( \30829 , RIe156630_2360, \16380 );
nor \g451790/U$1 ( \30830 , \30828 , \30829 );
and \g451789/U$2 ( \30831 , \16334 , RIe153930_2328);
and \g451789/U$3 ( \30832 , RIe164730_2520, \16328 );
nor \g451789/U$1 ( \30833 , \30831 , \30832 );
and \g445135/U$2 ( \30834 , \30827 , \30830 , \30833 );
nor \g445135/U$1 ( \30835 , \30834 , \16389 );
and \g445983/U$2 ( \30836 , RIfcb57a8_7087, \16427 );
and \g445983/U$3 ( \30837 , RIfca3058_6877, \16368 );
and \g448856/U$2 ( \30838 , RIfec2508_8331, \16344 );
and \g448856/U$3 ( \30839 , \16354 , RIfec2670_8332);
and \g448856/U$4 ( \30840 , RIfec27d8_8333, \16398 );
nor \g448856/U$1 ( \30841 , \30838 , \30839 , \30840 );
and \g454661/U$2 ( \30842 , \16317 , RIfcbc558_7165);
and \g454661/U$3 ( \30843 , RIfc78bf0_6396, \16325 );
nor \g454661/U$1 ( \30844 , \30842 , \30843 );
not \g449879/U$3 ( \30845 , \30844 );
not \g449879/U$4 ( \30846 , \16311 );
and \g449879/U$2 ( \30847 , \30845 , \30846 );
and \g449879/U$5 ( \30848 , \16341 , RIee38e78_5106);
nor \g449879/U$1 ( \30849 , \30847 , \30848 );
and \g451798/U$2 ( \30850 , \16377 , RIfca3fd0_6888);
and \g451798/U$3 ( \30851 , RIfca12d0_6856, \16313 );
nor \g451798/U$1 ( \30852 , \30850 , \30851 );
and \g451799/U$2 ( \30853 , \16334 , RIde84518_235);
and \g451799/U$3 ( \30854 , RIde88a00_256, \16380 );
nor \g451799/U$1 ( \30855 , \30853 , \30854 );
nand \g447308/U$1 ( \30856 , \30841 , \30849 , \30852 , \30855 );
nor \g445983/U$1 ( \30857 , \30836 , \30837 , \30856 );
and \g451797/U$2 ( \30858 , \16361 , RIe1672c8_2551);
and \g451797/U$3 ( \30859 , RIfcc35d8_7245, \16432 );
nor \g451797/U$1 ( \30860 , \30858 , \30859 );
and \g451796/U$2 ( \30861 , \16364 , RIfca3328_6879);
and \g451796/U$3 ( \30862 , RIfc5a290_6048, \16371 );
nor \g451796/U$1 ( \30863 , \30861 , \30862 );
and \g445136/U$2 ( \30864 , \30857 , \30860 , \30863 );
nor \g445136/U$1 ( \30865 , \30864 , \16649 );
or \g444211/U$1 ( \30866 , \30806 , \30835 , \30865 );
_DC \g524f/U$1 ( \30867 , \30866 , \16652 );
and \g450773/U$2 ( \30868 , \8326 , RIf16f0e8_5723);
and \g450773/U$3 ( \30869 , RIe1753c8_2711, \8404 );
nor \g450773/U$1 ( \30870 , \30868 , \30869 );
and \g445998/U$2 ( \30871 , RIf140090_5188, \8373 );
and \g445998/U$3 ( \30872 , RIf16dd38_5709, \8317 );
and \g448876/U$2 ( \30873 , RIee39850_5113, \8531 );
and \g448876/U$3 ( \30874 , \8488 , RIee3ac00_5127);
and \g448876/U$4 ( \30875 , RIf140900_5194, \8383 );
nor \g448876/U$1 ( \30876 , \30873 , \30874 , \30875 );
and \g451855/U$2 ( \30877 , \8356 , RIe172dd0_2684);
and \g451855/U$3 ( \30878 , RIee3bce0_5139, \8359 );
nor \g451855/U$1 ( \30879 , \30877 , \30878 );
and \g454440/U$2 ( \30880 , \8313 , RIee3e170_5165);
and \g454440/U$3 ( \30881 , RIf13ece0_5174, \8323 );
nor \g454440/U$1 ( \30882 , \30880 , \30881 );
not \g449557/U$3 ( \30883 , \30882 );
not \g449557/U$4 ( \30884 , \8376 );
and \g449557/U$2 ( \30885 , \30883 , \30884 );
and \g449557/U$5 ( \30886 , \8351 , RIf141e18_5209);
nor \g449557/U$1 ( \30887 , \30885 , \30886 );
and \g450741/U$2 ( \30888 , \8378 , RIee3cf28_5152);
and \g450741/U$3 ( \30889 , RIf13f988_5183, \8417 );
nor \g450741/U$1 ( \30890 , \30888 , \30889 );
nand \g447657/U$1 ( \30891 , \30876 , \30879 , \30887 , \30890 );
nor \g445998/U$1 ( \30892 , \30871 , \30872 , \30891 );
and \g451854/U$2 ( \30893 , \8335 , RIfce9120_7674);
and \g451854/U$3 ( \30894 , RIf16fc28_5731, \8340 );
nor \g451854/U$1 ( \30895 , \30893 , \30894 );
nand \g445575/U$1 ( \30896 , \30870 , \30892 , \30895 );
and \g444695/U$2 ( \30897 , \30896 , \9700 );
and \g448874/U$2 ( \30898 , RIfc68228_6207, \8531 );
and \g448874/U$3 ( \30899 , \8488 , RIe1861c8_2903);
and \g448874/U$4 ( \30900 , RIe199cc8_3127, \8330 );
nor \g448874/U$1 ( \30901 , \30898 , \30899 , \30900 );
and \g451852/U$2 ( \30902 , \8356 , RIe1834c8_2871);
and \g451852/U$3 ( \30903 , RIe188ec8_2935, \8359 );
nor \g451852/U$1 ( \30904 , \30902 , \30903 );
and \g454757/U$2 ( \30905 , \8313 , RIe1915c8_3031);
and \g454757/U$3 ( \30906 , RIe1942c8_3063, \8323 );
nor \g454757/U$1 ( \30907 , \30905 , \30906 );
not \g449897/U$3 ( \30908 , \30907 );
not \g449897/U$4 ( \30909 , \8376 );
and \g449897/U$2 ( \30910 , \30908 , \30909 );
and \g449897/U$5 ( \30911 , \8351 , RIe19c9c8_3159);
nor \g449897/U$1 ( \30912 , \30910 , \30911 );
and \g451851/U$2 ( \30913 , \8378 , RIe18e8c8_2999);
and \g451851/U$3 ( \30914 , RIfec20d0_8328, \8417 );
nor \g451851/U$1 ( \30915 , \30913 , \30914 );
nand \g447656/U$1 ( \30916 , \30901 , \30904 , \30912 , \30915 );
and \g444695/U$3 ( \30917 , \9702 , \30916 );
nor \g444695/U$1 ( \30918 , \30897 , \30917 );
and \g446784/U$2 ( \30919 , \9724 , RIe196fc8_3095);
and \g446784/U$3 ( \30920 , RIfe8ea28_7967, \9726 );
nor \g446784/U$1 ( \30921 , \30919 , \30920 );
and \g446783/U$2 ( \30922 , \9729 , RIe17adc8_2775);
and \g446783/U$3 ( \30923 , RIe17dac8_2807, \9731 );
nor \g446783/U$1 ( \30924 , \30922 , \30923 );
and \g446782/U$2 ( \30925 , \9734 , RIe1807c8_2839);
and \g446782/U$3 ( \30926 , RIfccb5d0_7336, \9736 );
nor \g446782/U$1 ( \30927 , \30925 , \30926 );
nand \g444482/U$1 ( \30928 , \30918 , \30921 , \30924 , \30927 );
and \g451861/U$2 ( \30929 , \8326 , RIf146030_5256);
and \g451861/U$3 ( \30930 , RIe1b6a08_3455, \8404 );
nor \g451861/U$1 ( \30931 , \30929 , \30930 );
and \g446000/U$2 ( \30932 , RIe1b8a60_3478, \8371 );
and \g446000/U$3 ( \30933 , RIfe8dee8_7959, \8317 );
and \g448879/U$2 ( \30934 , RIfe8e050_7960, \8531 );
and \g448879/U$3 ( \30935 , \8488 , RIf147818_5273);
and \g448879/U$4 ( \30936 , RIfc5ea48_6099, \8383 );
nor \g448879/U$1 ( \30937 , \30934 , \30935 , \30936 );
and \g453969/U$2 ( \30938 , \8356 , RIfe8e488_7963);
and \g453969/U$3 ( \30939 , RIf1488f8_5285, \8359 );
nor \g453969/U$1 ( \30940 , \30938 , \30939 );
and \g454679/U$2 ( \30941 , \8313 , RIfe8e5f0_7964);
and \g454679/U$3 ( \30942 , RIfc44fa8_5807, \8323 );
nor \g454679/U$1 ( \30943 , \30941 , \30942 );
not \g449901/U$3 ( \30944 , \30943 );
not \g449901/U$4 ( \30945 , \8376 );
and \g449901/U$2 ( \30946 , \30944 , \30945 );
and \g449901/U$5 ( \30947 , \8351 , RIfca4de0_6898);
nor \g449901/U$1 ( \30948 , \30946 , \30947 );
and \g451863/U$2 ( \30949 , \8378 , RIfe8e1b8_7961);
and \g451863/U$3 ( \30950 , RIfcbd638_7177, \8417 );
nor \g451863/U$1 ( \30951 , \30949 , \30950 );
nand \g447659/U$1 ( \30952 , \30937 , \30940 , \30948 , \30951 );
nor \g446000/U$1 ( \30953 , \30932 , \30933 , \30952 );
and \g451862/U$2 ( \30954 , \8335 , RIfe8e320_7962);
and \g451862/U$3 ( \30955 , RIf146e40_5266, \8340 );
nor \g451862/U$1 ( \30956 , \30954 , \30955 );
nand \g445577/U$1 ( \30957 , \30931 , \30953 , \30956 );
and \g444828/U$2 ( \30958 , \30957 , \8482 );
and \g448877/U$2 ( \30959 , RIe1c0788_3567, \8319 );
and \g448877/U$3 ( \30960 , \8326 , RIe1c3488_3599);
and \g448877/U$4 ( \30961 , RIe1ce888_3727, \8486 );
nor \g448877/U$1 ( \30962 , \30959 , \30960 , \30961 );
and \g451857/U$2 ( \30963 , \8335 , RIe1bda88_3535);
and \g451857/U$3 ( \30964 , RIe1c6188_3631, \8340 );
nor \g451857/U$1 ( \30965 , \30963 , \30964 );
and \g450579/U$2 ( \30966 , \8404 , RIe1e2388_3951);
and \g450579/U$3 ( \30967 , RIe1eaa88_4047, \8351 );
nor \g450579/U$1 ( \30968 , \30966 , \30967 );
and \g454157/U$2 ( \30969 , \8313 , RIe1e5088_3983);
and \g454157/U$3 ( \30970 , RIe1e7d88_4015, \8323 );
nor \g454157/U$1 ( \30971 , \30969 , \30970 );
not \g449899/U$3 ( \30972 , \30971 );
not \g449899/U$4 ( \30973 , \8328 );
and \g449899/U$2 ( \30974 , \30972 , \30973 );
and \g449899/U$5 ( \30975 , \8359 , RIe1d1588_3759);
nor \g449899/U$1 ( \30976 , \30974 , \30975 );
nand \g447658/U$1 ( \30977 , \30962 , \30965 , \30968 , \30976 );
and \g444828/U$3 ( \30978 , \8478 , \30977 );
nor \g444828/U$1 ( \30979 , \30958 , \30978 );
and \g446788/U$2 ( \30980 , \10534 , RIe1dc988_3887);
and \g446788/U$3 ( \30981 , RIe1df688_3919, \10536 );
nor \g446788/U$1 ( \30982 , \30980 , \30981 );
and \g446789/U$2 ( \30983 , \10539 , RIe1d6f88_3823);
and \g446789/U$3 ( \30984 , RIe1d9c88_3855, \10541 );
nor \g446789/U$1 ( \30985 , \30983 , \30984 );
and \g446791/U$2 ( \30986 , \8775 , RIe1c8e88_3663);
and \g446791/U$3 ( \30987 , RIe1cbb88_3695, \8777 );
nor \g446791/U$1 ( \30988 , \30986 , \30987 );
nand \g444599/U$1 ( \30989 , \30979 , \30982 , \30985 , \30988 );
and \g445995/U$2 ( \30990 , RIe21d320_4622, \8407 );
and \g445995/U$3 ( \30991 , RIe214c20_4526, \8378 );
and \g448871/U$2 ( \30992 , RIf16b8a8_5683, \8373 );
and \g448871/U$3 ( \30993 , \8383 , RIe222d20_4686);
and \g448871/U$4 ( \30994 , RIe211f20_4494, \8488 );
nor \g448871/U$1 ( \30995 , \30992 , \30993 , \30994 );
and \g451843/U$2 ( \30996 , \8335 , RIe206b20_4366);
and \g451843/U$3 ( \30997 , RIfe8e758_7965, \8340 );
nor \g451843/U$1 ( \30998 , \30996 , \30997 );
and \g451842/U$2 ( \30999 , \8404 , RIe220020_4654);
and \g451842/U$3 ( \31000 , RIfc404a8_5757, \8351 );
nor \g451842/U$1 ( \31001 , \30999 , \31000 );
and \g454253/U$2 ( \31002 , \8313 , RIe209820_4398);
and \g454253/U$3 ( \31003 , RIe20c520_4430, \8323 );
nor \g454253/U$1 ( \31004 , \31002 , \31003 );
not \g454252/U$1 ( \31005 , \31004 );
and \g449894/U$2 ( \31006 , \31005 , \8316 );
and \g449894/U$3 ( \31007 , RIfc5b910_6064, \8359 );
nor \g449894/U$1 ( \31008 , \31006 , \31007 );
nand \g448175/U$1 ( \31009 , \30995 , \30998 , \31001 , \31008 );
nor \g445995/U$1 ( \31010 , \30990 , \30991 , \31009 );
and \g451841/U$2 ( \31011 , \8356 , RIe20f220_4462);
and \g451841/U$3 ( \31012 , RIf16a930_5672, \8417 );
nor \g451841/U$1 ( \31013 , \31011 , \31012 );
and \g451840/U$2 ( \31014 , \8523 , RIfe8e8c0_7966);
and \g451840/U$3 ( \31015 , RIe217920_4558, \8414 );
nor \g451840/U$1 ( \31016 , \31014 , \31015 );
and \g445147/U$2 ( \31017 , \31010 , \31013 , \31016 );
nor \g445147/U$1 ( \31018 , \31017 , \8368 );
and \g445996/U$2 ( \31019 , RIf162ed8_5585, \8414 );
and \g445996/U$3 ( \31020 , RIf164c60_5606, \8417 );
and \g448872/U$2 ( \31021 , RIfe8dd80_7958, \8373 );
and \g448872/U$3 ( \31022 , \8383 , RIf165a70_5616);
and \g448872/U$4 ( \31023 , RIf15da78_5525, \8488 );
nor \g448872/U$1 ( \31024 , \31021 , \31022 , \31023 );
and \g451848/U$2 ( \31025 , \8335 , RIf159860_5478);
and \g451848/U$3 ( \31026 , RIf15c560_5510, \8340 );
nor \g451848/U$1 ( \31027 , \31025 , \31026 );
and \g451058/U$2 ( \31028 , \8404 , RIfe8dab0_7956);
and \g451058/U$3 ( \31029 , RIf166b50_5628, \8351 );
nor \g451058/U$1 ( \31030 , \31028 , \31029 );
and \g455255/U$2 ( \31031 , \8313 , RIfc62828_6143);
and \g455255/U$3 ( \31032 , RIf15b048_5495, \8323 );
nor \g455255/U$1 ( \31033 , \31031 , \31032 );
not \g455254/U$1 ( \31034 , \31033 );
and \g449896/U$2 ( \31035 , \31034 , \8316 );
and \g449896/U$3 ( \31036 , RIf15f800_5546, \8359 );
nor \g449896/U$1 ( \31037 , \31035 , \31036 );
nand \g448176/U$1 ( \31038 , \31024 , \31027 , \31030 , \31037 );
nor \g445996/U$1 ( \31039 , \31019 , \31020 , \31038 );
and \g451844/U$2 ( \31040 , \8378 , RIf1616f0_5568);
and \g451844/U$3 ( \31041 , RIfe8d948_7955, \8523 );
nor \g451844/U$1 ( \31042 , \31040 , \31041 );
and \g451845/U$2 ( \31043 , \8356 , RIfe8dc18_7957);
and \g451845/U$3 ( \31044 , RIf163e50_5596, \8409 );
nor \g451845/U$1 ( \31045 , \31043 , \31044 );
and \g445148/U$2 ( \31046 , \31039 , \31042 , \31045 );
nor \g445148/U$1 ( \31047 , \31046 , \8422 );
or \g444366/U$1 ( \31048 , \30928 , \30989 , \31018 , \31047 );
and \g445990/U$2 ( \31049 , RIfc61748_6131, \8409 );
and \g445990/U$3 ( \31050 , RIe1f4ad8_4161, \8378 );
and \g448866/U$2 ( \31051 , RIfca6e38_6921, \8373 );
and \g448866/U$3 ( \31052 , \8383 , RIf157538_5453);
and \g448866/U$4 ( \31053 , RIf151700_5386, \8486 );
nor \g448866/U$1 ( \31054 , \31051 , \31052 , \31053 );
and \g451505/U$2 ( \31055 , \8335 , RIe1ed4b8_4077);
and \g451505/U$3 ( \31056 , RIfc60ed8_6125, \8340 );
nor \g451505/U$1 ( \31057 , \31055 , \31056 );
and \g451830/U$2 ( \31058 , \8404 , RIe1f9b00_4218);
and \g451830/U$3 ( \31059 , RIf158780_5466, \8351 );
nor \g451830/U$1 ( \31060 , \31058 , \31059 );
and \g454599/U$2 ( \31061 , \8313 , RIf14d7b8_5341);
and \g454599/U$3 ( \31062 , RIfc7b620_6426, \8323 );
nor \g454599/U$1 ( \31063 , \31061 , \31062 );
not \g454598/U$1 ( \31064 , \31063 );
and \g449890/U$2 ( \31065 , \31064 , \8316 );
and \g449890/U$3 ( \31066 , RIf152ab0_5400, \8359 );
nor \g449890/U$1 ( \31067 , \31065 , \31066 );
nand \g448173/U$1 ( \31068 , \31054 , \31057 , \31060 , \31067 );
nor \g445990/U$1 ( \31069 , \31049 , \31050 , \31068 );
and \g451829/U$2 ( \31070 , \8356 , RIe1f27b0_4136);
and \g451829/U$3 ( \31071 , RIfc61e50_6136, \8417 );
nor \g451829/U$1 ( \31072 , \31070 , \31071 );
and \g451828/U$2 ( \31073 , \8523 , RIf1501e8_5371);
and \g451828/U$3 ( \31074 , RIf154130_5416, \8414 );
nor \g451828/U$1 ( \31075 , \31073 , \31074 );
and \g445142/U$2 ( \31076 , \31069 , \31072 , \31075 );
nor \g445142/U$1 ( \31077 , \31076 , \8621 );
and \g445993/U$2 ( \31078 , RIe1a23c8_3223, \8371 );
and \g445993/U$3 ( \31079 , RIe225a20_4718, \8412 );
and \g448869/U$2 ( \31080 , RIe1f7238_4189, \8523 );
and \g448869/U$3 ( \31081 , \8488 , RIe1fde80_4266);
and \g448869/U$4 ( \31082 , RIe1a50c8_3255, \8383 );
nor \g448869/U$1 ( \31083 , \31080 , \31081 , \31082 );
and \g451837/U$2 ( \31084 , \8335 , RIe170238_2653);
and \g451837/U$3 ( \31085 , RIe1d4288_3791, \8340 );
nor \g451837/U$1 ( \31086 , \31084 , \31085 );
and \g455156/U$2 ( \31087 , \8313 , RIe1adc00_3354);
and \g455156/U$3 ( \31088 , RIe1bad88_3503, \8323 );
nor \g455156/U$1 ( \31089 , \31087 , \31088 );
not \g455155/U$1 ( \31090 , \31089 );
and \g449891/U$2 ( \31091 , \31090 , \8316 );
and \g449891/U$3 ( \31092 , RIe1a7dc8_3287, \8351 );
nor \g449891/U$1 ( \31093 , \31091 , \31092 );
and \g451367/U$2 ( \31094 , \8356 , RIe1efd80_4106);
and \g451367/U$3 ( \31095 , RIe203e20_4334, \8359 );
nor \g451367/U$1 ( \31096 , \31094 , \31095 );
nand \g448174/U$1 ( \31097 , \31083 , \31086 , \31093 , \31096 );
nor \g445993/U$1 ( \31098 , \31078 , \31079 , \31097 );
and \g451834/U$2 ( \31099 , \8404 , RIe19f6c8_3191);
and \g451834/U$3 ( \31100 , RIe18bbc8_2967, \8417 );
nor \g451834/U$1 ( \31101 , \31099 , \31100 );
and \g451835/U$2 ( \31102 , \8378 , RIe21a620_4590);
and \g451835/U$3 ( \31103 , RIe1780c8_2743, \8409 );
nor \g451835/U$1 ( \31104 , \31102 , \31103 );
and \g445145/U$2 ( \31105 , \31098 , \31101 , \31104 );
nor \g445145/U$1 ( \31106 , \31105 , \8651 );
or \g444189/U$1 ( \31107 , \31048 , \31077 , \31106 );
_DC \g52d3/U$1 ( \31108 , \31107 , \8654 );
and \g452127/U$2 ( \31109 , \16398 , RIdee6768_1086);
and \g452127/U$3 ( \31110 , RIdec7598_732, \16377 );
nor \g452127/U$1 ( \31111 , \31109 , \31110 );
and \g446072/U$2 ( \31112 , RIdeca298_764, \16313 );
and \g446072/U$3 ( \31113 , RIde7ae28_189, \16361 );
and \g448968/U$2 ( \31114 , RIdeccf98_796, \16321 );
and \g448968/U$3 ( \31115 , \16485 , RIde94ee0_316);
and \g448968/U$4 ( \31116 , RIdeb3a98_508, \16356 );
nor \g448968/U$1 ( \31117 , \31114 , \31115 , \31116 );
and \g452130/U$2 ( \31118 , \16368 , RIdf1c570_1699);
and \g452130/U$3 ( \31119 , RIdf2bcf0_1875, \16371 );
nor \g452130/U$1 ( \31120 , \31118 , \31119 );
and \g454733/U$2 ( \31121 , \16317 , RIdf37690_2007);
and \g454733/U$3 ( \31122 , RIe142c98_2137, \16325 );
nor \g454733/U$1 ( \31123 , \31121 , \31122 );
not \g449982/U$3 ( \31124 , \31123 );
not \g449982/U$4 ( \31125 , \16351 );
and \g449982/U$2 ( \31126 , \31124 , \31125 );
and \g449982/U$5 ( \31127 , \16328 , RIdecfc98_828);
nor \g449982/U$1 ( \31128 , \31126 , \31127 );
and \g452129/U$2 ( \31129 , \16334 , RIe159498_2393);
and \g452129/U$3 ( \31130 , RIe16d6a0_2622, \16380 );
nor \g452129/U$1 ( \31131 , \31129 , \31130 );
nand \g447711/U$1 ( \31132 , \31117 , \31120 , \31128 , \31131 );
nor \g446072/U$1 ( \31133 , \31112 , \31113 , \31132 );
and \g452128/U$2 ( \31134 , \16364 , RIdedb4d0_959);
and \g452128/U$3 ( \31135 , RIdeffc68_1374, \16341 );
nor \g452128/U$1 ( \31136 , \31134 , \31135 );
nand \g445592/U$1 ( \31137 , \31111 , \31133 , \31136 );
and \g444891/U$2 ( \31138 , \31137 , \16752 );
and \g448967/U$2 ( \31139 , RIee24568_4872, \16321 );
and \g448967/U$3 ( \31140 , \16328 , RIee25378_4882);
and \g448967/U$4 ( \31141 , RIee220d8_4846, \16427 );
nor \g448967/U$1 ( \31142 , \31139 , \31140 , \31141 );
and \g452124/U$2 ( \31143 , \16361 , RIfe8b080_7926);
and \g452124/U$3 ( \31144 , RIded49f0_883, \16364 );
nor \g452124/U$1 ( \31145 , \31143 , \31144 );
and \g452123/U$2 ( \31146 , \16377 , RIee23050_4857);
and \g452123/U$3 ( \31147 , RIee23a28_4864, \16313 );
nor \g452123/U$1 ( \31148 , \31146 , \31147 );
and \g454386/U$2 ( \31149 , \16317 , RIfe8af18_7925);
and \g454386/U$3 ( \31150 , RIded8ed8_932, \16325 );
nor \g454386/U$1 ( \31151 , \31149 , \31150 );
not \g454385/U$1 ( \31152 , \31151 );
and \g449981/U$2 ( \31153 , \31152 , \16336 );
and \g449981/U$3 ( \31154 , RIfca5650_6904, \16448 );
nor \g449981/U$1 ( \31155 , \31153 , \31154 );
nand \g448003/U$1 ( \31156 , \31142 , \31145 , \31148 , \31155 );
and \g444891/U$3 ( \31157 , \16477 , \31156 );
nor \g444891/U$1 ( \31158 , \31138 , \31157 );
and \g446846/U$2 ( \31159 , \17473 , RIee20ff8_4834);
and \g446846/U$3 ( \31160 , RIfceeb20_7738, \17475 );
nor \g446846/U$1 ( \31161 , \31159 , \31160 );
and \g446845/U$2 ( \31162 , \22390 , RIdee23e8_1038);
and \g446845/U$3 ( \31163 , RIfe8adb0_7924, \22392 );
nor \g446845/U$1 ( \31164 , \31162 , \31163 );
and \g446847/U$2 ( \31165 , \18278 , RIdede1d0_991);
and \g446847/U$3 ( \31166 , RIfe8ac48_7923, \18280 );
nor \g446847/U$1 ( \31167 , \31165 , \31166 );
nand \g444605/U$1 ( \31168 , \31158 , \31161 , \31164 , \31167 );
and \g452119/U$2 ( \31169 , \16337 , RIdeeee68_1182);
and \g452119/U$3 ( \31170 , RIdf02968_1406, \16334 );
nor \g452119/U$1 ( \31171 , \31169 , \31170 );
and \g446068/U$2 ( \31172 , RIdf05668_1438, \16380 );
and \g446068/U$3 ( \31173 , RIdee9468_1118, \16361 );
and \g448965/U$2 ( \31174 , RIdefa268_1310, \16427 );
and \g448965/U$3 ( \31175 , \16448 , RIdefcf68_1342);
and \g448965/U$4 ( \31176 , RIdf08368_1470, \16485 );
nor \g448965/U$1 ( \31177 , \31174 , \31175 , \31176 );
and \g454729/U$2 ( \31178 , \16317 , RIdf13768_1598);
and \g454729/U$3 ( \31179 , RIdf16468_1630, \16325 );
nor \g454729/U$1 ( \31180 , \31178 , \31179 );
not \g449980/U$3 ( \31181 , \31180 );
not \g449980/U$4 ( \31182 , \16311 );
and \g449980/U$2 ( \31183 , \31181 , \31182 );
and \g449980/U$5 ( \31184 , \16356 , RIdf0b068_1502);
nor \g449980/U$1 ( \31185 , \31183 , \31184 );
and \g451269/U$2 ( \31186 , \16377 , RIdf0dd68_1534);
and \g451269/U$3 ( \31187 , RIdf10a68_1566, \16313 );
nor \g451269/U$1 ( \31188 , \31186 , \31187 );
and \g452121/U$2 ( \31189 , \16368 , RIdef4868_1246);
and \g452121/U$3 ( \31190 , RIdef7568_1278, \16371 );
nor \g452121/U$1 ( \31191 , \31189 , \31190 );
nand \g447710/U$1 ( \31192 , \31177 , \31185 , \31188 , \31191 );
nor \g446068/U$1 ( \31193 , \31172 , \31173 , \31192 );
and \g452893/U$2 ( \31194 , \16364 , RIdeec168_1150);
and \g452893/U$3 ( \31195 , RIdef1b68_1214, \16341 );
nor \g452893/U$1 ( \31196 , \31194 , \31195 );
nand \g445590/U$1 ( \31197 , \31171 , \31193 , \31196 );
and \g444774/U$2 ( \31198 , \31197 , \16750 );
and \g448964/U$2 ( \31199 , RIfc6ac58_6237, \16427 );
and \g448964/U$3 ( \31200 , \16337 , RIdf1f108_1730);
and \g448964/U$4 ( \31201 , RIdf21160_1753, \16341 );
nor \g448964/U$1 ( \31202 , \31199 , \31200 , \31201 );
and \g452116/U$2 ( \31203 , \16361 , RIfeaa7f0_8256);
and \g452116/U$3 ( \31204 , RIdf1ac20_1681, \16364 );
nor \g452116/U$1 ( \31205 , \31203 , \31204 );
and \g451591/U$2 ( \31206 , \16377 , RIee276a0_4907);
and \g451591/U$3 ( \31207 , RIee28a50_4921, \16313 );
nor \g451591/U$1 ( \31208 , \31206 , \31207 );
and \g454641/U$2 ( \31209 , \16317 , RIee29e00_4935);
and \g454641/U$3 ( \31210 , RIee2b5e8_4952, \16325 );
nor \g454641/U$1 ( \31211 , \31209 , \31210 );
not \g450313/U$3 ( \31212 , \31211 );
not \g450313/U$4 ( \31213 , \16311 );
and \g450313/U$2 ( \31214 , \31212 , \31213 );
and \g450313/U$5 ( \31215 , \16448 , RIfc6aaf0_6236);
nor \g450313/U$1 ( \31216 , \31214 , \31215 );
nand \g447709/U$1 ( \31217 , \31202 , \31205 , \31208 , \31216 );
and \g444774/U$3 ( \31218 , \16481 , \31217 );
nor \g444774/U$1 ( \31219 , \31198 , \31218 );
and \g446842/U$2 ( \31220 , \16511 , RIdf23fc8_1786);
and \g446842/U$3 ( \31221 , RIdf25be8_1806, \16514 );
nor \g446842/U$1 ( \31222 , \31220 , \31221 );
and \g446841/U$2 ( \31223 , \24165 , RIdf27970_1827);
and \g446841/U$3 ( \31224 , RIdf29c98_1852, \24167 );
nor \g446841/U$1 ( \31225 , \31223 , \31224 );
and \g446840/U$2 ( \31226 , \17279 , RIfcdd4b0_7540);
and \g446840/U$3 ( \31227 , RIdf22678_1768, \17281 );
nor \g446840/U$1 ( \31228 , \31226 , \31227 );
nand \g444493/U$1 ( \31229 , \31219 , \31222 , \31225 , \31228 );
and \g446064/U$2 ( \31230 , RIfce6b28_7647, \16356 );
and \g446064/U$3 ( \31231 , RIdeae098_444, \16368 );
and \g448961/U$2 ( \31232 , RIdeb0d98_476, \16427 );
and \g448961/U$3 ( \31233 , \16398 , RIdea89e0_412);
and \g448961/U$4 ( \31234 , RIfcaa510_6960, \16339 );
nor \g448961/U$1 ( \31235 , \31232 , \31233 , \31234 );
and \g452109/U$2 ( \31236 , \16361 , RIde9b7e0_348);
and \g452109/U$3 ( \31237 , RIdea20e0_380, \16364 );
nor \g452109/U$1 ( \31238 , \31236 , \31237 );
and \g452107/U$2 ( \31239 , \16377 , RIdebee98_636);
and \g452107/U$3 ( \31240 , RIfc661d0_6184, \16313 );
nor \g452107/U$1 ( \31241 , \31239 , \31240 );
and \g454720/U$2 ( \31242 , \16317 , RIdec1b98_668);
and \g454720/U$3 ( \31243 , RIdec4898_700, \16325 );
nor \g454720/U$1 ( \31244 , \31242 , \31243 );
not \g449977/U$3 ( \31245 , \31244 );
not \g449977/U$4 ( \31246 , \16311 );
and \g449977/U$2 ( \31247 , \31245 , \31246 );
and \g449977/U$5 ( \31248 , \16448 , RIfc40d18_5763);
nor \g449977/U$1 ( \31249 , \31247 , \31248 );
nand \g447706/U$1 ( \31250 , \31235 , \31238 , \31241 , \31249 );
nor \g446064/U$1 ( \31251 , \31230 , \31231 , \31250 );
and \g452105/U$2 ( \31252 , \16334 , RIdeb6798_540);
and \g452105/U$3 ( \31253 , RIfcad648_6995, \16371 );
nor \g452105/U$1 ( \31254 , \31252 , \31253 );
and \g452104/U$2 ( \31255 , \16380 , RIdeb9498_572);
and \g452104/U$3 ( \31256 , RIdebc198_604, \16485 );
nor \g452104/U$1 ( \31257 , \31255 , \31256 );
and \g445200/U$2 ( \31258 , \31251 , \31254 , \31257 );
nor \g445200/U$1 ( \31259 , \31258 , \16618 );
and \g446066/U$2 ( \31260 , RIee31b28_5024, \16313 );
and \g446066/U$3 ( \31261 , RIdf2e9f0_1907, \16361 );
and \g448963/U$2 ( \31262 , RIee2f260_4995, \16427 );
and \g448963/U$3 ( \31263 , \16448 , RIfc6b1f8_6241);
and \g448963/U$4 ( \31264 , RIfe8a6a8_7919, \16319 );
nor \g448963/U$1 ( \31265 , \31262 , \31263 , \31264 );
and \g452113/U$2 ( \31266 , \16368 , RIee2d0a0_4971);
and \g452113/U$3 ( \31267 , RIfc70d60_6306, \16371 );
nor \g452113/U$1 ( \31268 , \31266 , \31267 );
and \g454605/U$2 ( \31269 , \16317 , RIfe8a540_7918);
and \g454605/U$3 ( \31270 , RIe140808_2111, \16325 );
nor \g454605/U$1 ( \31271 , \31269 , \31270 );
not \g449609/U$3 ( \31272 , \31271 );
not \g449609/U$4 ( \31273 , \16330 );
and \g449609/U$2 ( \31274 , \31272 , \31273 );
and \g449609/U$5 ( \31275 , \16328 , RIfe8a810_7920);
nor \g449609/U$1 ( \31276 , \31274 , \31275 );
and \g452112/U$2 ( \31277 , \16334 , RIdf3a0c0_2037);
and \g452112/U$3 ( \31278 , RIdf3c3e8_2062, \16380 );
nor \g452112/U$1 ( \31279 , \31277 , \31278 );
nand \g447707/U$1 ( \31280 , \31265 , \31268 , \31276 , \31279 );
nor \g446066/U$1 ( \31281 , \31260 , \31261 , \31280 );
and \g452111/U$2 ( \31282 , \16364 , RIdf308e0_1929);
and \g452111/U$3 ( \31283 , RIfe8a978_7921, \16339 );
nor \g452111/U$1 ( \31284 , \31282 , \31283 );
and \g451515/U$2 ( \31285 , \16398 , RIdf32c08_1954);
and \g451515/U$3 ( \31286 , RIee30e80_5015, \16377 );
nor \g451515/U$1 ( \31287 , \31285 , \31286 );
and \g445201/U$2 ( \31288 , \31281 , \31284 , \31287 );
nor \g445201/U$1 ( \31289 , \31288 , \16393 );
or \g444395/U$1 ( \31290 , \31168 , \31229 , \31259 , \31289 );
and \g446061/U$2 ( \31291 , RIfe8a270_7916, \16356 );
and \g446061/U$3 ( \31292 , RIe153a98_2329, \16334 );
and \g448958/U$2 ( \31293 , RIe161b98_2489, \16319 );
and \g448958/U$3 ( \31294 , \16328 , RIe164898_2521);
and \g448958/U$4 ( \31295 , RIe150d98_2297, \16427 );
nor \g448958/U$1 ( \31296 , \31293 , \31294 , \31295 );
and \g452096/U$2 ( \31297 , \16361 , RIe145998_2169);
and \g452096/U$3 ( \31298 , RIe148698_2201, \16364 );
nor \g452096/U$1 ( \31299 , \31297 , \31298 );
and \g452095/U$2 ( \31300 , \16377 , RIe15ee98_2457);
and \g452095/U$3 ( \31301 , RIfe8a3d8_7917, \16313 );
nor \g452095/U$1 ( \31302 , \31300 , \31301 );
and \g454717/U$2 ( \31303 , \16317 , RIe14b398_2233);
and \g454717/U$3 ( \31304 , RIfcca658_7325, \16325 );
nor \g454717/U$1 ( \31305 , \31303 , \31304 );
not \g454716/U$1 ( \31306 , \31305 );
and \g449975/U$2 ( \31307 , \31306 , \16336 );
and \g449975/U$3 ( \31308 , RIfc3f0f8_5743, \16432 );
nor \g449975/U$1 ( \31309 , \31307 , \31308 );
nand \g448064/U$1 ( \31310 , \31296 , \31299 , \31302 , \31309 );
nor \g446061/U$1 ( \31311 , \31291 , \31292 , \31310 );
and \g452092/U$2 ( \31312 , \16371 , RIfcab050_6968);
and \g452092/U$3 ( \31313 , RIe156798_2361, \16380 );
nor \g452092/U$1 ( \31314 , \31312 , \31313 );
and \g452093/U$2 ( \31315 , \16368 , RIe14e098_2265);
and \g452093/U$3 ( \31316 , RIe15c198_2425, \16344 );
nor \g452093/U$1 ( \31317 , \31315 , \31316 );
and \g445196/U$2 ( \31318 , \31311 , \31314 , \31317 );
nor \g445196/U$1 ( \31319 , \31318 , \16389 );
and \g446062/U$2 ( \31320 , RIfc6f6e0_6290, \16313 );
and \g446062/U$3 ( \31321 , RIe1695f0_2576, \16364 );
and \g448960/U$2 ( \31322 , RIfca8350_6936, \16321 );
and \g448960/U$3 ( \31323 , \16485 , RIfe8aae0_7922);
and \g448960/U$4 ( \31324 , RIde8fcd8_291, \16356 );
nor \g448960/U$1 ( \31325 , \31322 , \31323 , \31324 );
and \g452101/U$2 ( \31326 , \16368 , RIfcadeb8_7001);
and \g452101/U$3 ( \31327 , RIfcae020_7002, \16371 );
nor \g452101/U$1 ( \31328 , \31326 , \31327 );
and \g455087/U$2 ( \31329 , \16317 , RIfc64718_6165);
and \g455087/U$3 ( \31330 , RIde80a08_217, \16325 );
nor \g455087/U$1 ( \31331 , \31329 , \31330 );
not \g450226/U$3 ( \31332 , \31331 );
not \g450226/U$4 ( \31333 , \16351 );
and \g450226/U$2 ( \31334 , \31332 , \31333 );
and \g450226/U$5 ( \31335 , \16328 , RIfcab320_6970);
nor \g450226/U$1 ( \31336 , \31334 , \31335 );
and \g453348/U$2 ( \31337 , \16334 , RIde84860_236);
and \g453348/U$3 ( \31338 , RIde88d48_257, \16380 );
nor \g453348/U$1 ( \31339 , \31337 , \31338 );
nand \g447705/U$1 ( \31340 , \31325 , \31328 , \31336 , \31339 );
nor \g446062/U$1 ( \31341 , \31320 , \31321 , \31340 );
and \g453685/U$2 ( \31342 , \16341 , RIee38fe0_5107);
and \g453685/U$3 ( \31343 , RIfcaa240_6958, \16377 );
nor \g453685/U$1 ( \31344 , \31342 , \31343 );
and \g452100/U$2 ( \31345 , \16361 , RIe167430_2552);
and \g452100/U$3 ( \31346 , RIe16add8_2593, \16337 );
nor \g452100/U$1 ( \31347 , \31345 , \31346 );
and \g445197/U$2 ( \31348 , \31341 , \31344 , \31347 );
nor \g445197/U$1 ( \31349 , \31348 , \16649 );
or \g444216/U$1 ( \31350 , \31290 , \31319 , \31349 );
_DC \g5358/U$1 ( \31351 , \31350 , \16652 );
and \g448976/U$2 ( \31352 , RIfc6c440_6254, \8319 );
and \g448976/U$3 ( \31353 , \8324 , RIf16f250_5724);
and \g448976/U$4 ( \31354 , RIfcabb90_6976, \8486 );
nor \g448976/U$1 ( \31355 , \31352 , \31353 , \31354 );
and \g452155/U$2 ( \31356 , \8335 , RIfcaba28_6975);
and \g452155/U$3 ( \31357 , RIf16fd90_5732, \8340 );
nor \g452155/U$1 ( \31358 , \31356 , \31357 );
and \g453144/U$2 ( \31359 , \8404 , RIfea7af0_8224);
and \g453144/U$3 ( \31360 , RIfcccc50_7352, \8351 );
nor \g453144/U$1 ( \31361 , \31359 , \31360 );
and \g455077/U$2 ( \31362 , \8313 , RIe176d18_2729);
and \g455077/U$3 ( \31363 , RIfcccdb8_7353, \8323 );
nor \g455077/U$1 ( \31364 , \31362 , \31363 );
not \g449991/U$3 ( \31365 , \31364 );
not \g449991/U$4 ( \31366 , \8328 );
and \g449991/U$2 ( \31367 , \31365 , \31366 );
and \g449991/U$5 ( \31368 , \8359 , RIfca9868_6951);
nor \g449991/U$1 ( \31369 , \31367 , \31368 );
nand \g447810/U$1 ( \31370 , \31355 , \31358 , \31361 , \31369 );
and \g444686/U$2 ( \31371 , \31370 , \9700 );
and \g446080/U$2 ( \31372 , RIfcabcf8_6977, \8340 );
and \g446080/U$3 ( \31373 , RIe197130_3096, \8404 );
and \g448978/U$2 ( \31374 , RIfc6c878_6257, \8531 );
and \g448978/U$3 ( \31375 , \8488 , RIe186330_2904);
and \g448978/U$4 ( \31376 , RIe199e30_3128, \8383 );
nor \g448978/U$1 ( \31377 , \31374 , \31375 , \31376 );
and \g452162/U$2 ( \31378 , \8356 , RIe183630_2872);
and \g452162/U$3 ( \31379 , RIe189030_2936, \8359 );
nor \g452162/U$1 ( \31380 , \31378 , \31379 );
and \g454742/U$2 ( \31381 , \8313 , RIe191730_3032);
and \g454742/U$3 ( \31382 , RIe194430_3064, \8323 );
nor \g454742/U$1 ( \31383 , \31381 , \31382 );
not \g449756/U$3 ( \31384 , \31383 );
not \g449756/U$4 ( \31385 , \8376 );
and \g449756/U$2 ( \31386 , \31384 , \31385 );
and \g449756/U$5 ( \31387 , \8351 , RIe19cb30_3160);
nor \g449756/U$1 ( \31388 , \31386 , \31387 );
and \g452160/U$2 ( \31389 , \8378 , RIe18ea30_3000);
and \g452160/U$3 ( \31390 , RIfe8a108_7915, \8417 );
nor \g452160/U$1 ( \31391 , \31389 , \31390 );
nand \g447717/U$1 ( \31392 , \31377 , \31380 , \31388 , \31391 );
nor \g446080/U$1 ( \31393 , \31372 , \31373 , \31392 );
and \g452158/U$2 ( \31394 , \8335 , RIe17af30_2776);
and \g452158/U$3 ( \31395 , RIf145388_5247, \8373 );
nor \g452158/U$1 ( \31396 , \31394 , \31395 );
and \g452159/U$2 ( \31397 , \8319 , RIe17dc30_2808);
and \g452159/U$3 ( \31398 , RIe180930_2840, \8326 );
nor \g452159/U$1 ( \31399 , \31397 , \31398 );
and \g445209/U$2 ( \31400 , \31393 , \31396 , \31399 );
nor \g445209/U$1 ( \31401 , \31400 , \8589 );
nor \g444686/U$1 ( \31402 , \31371 , \31401 );
and \g446852/U$2 ( \31403 , \12254 , RIfccb738_7337);
and \g446852/U$3 ( \31404 , RIfcdd078_7537, \12256 );
nor \g446852/U$1 ( \31405 , \31403 , \31404 );
and \g446851/U$2 ( \31406 , \26544 , RIfe89e38_7913);
and \g446851/U$3 ( \31407 , RIfe89fa0_7914, \26546 );
nor \g446851/U$1 ( \31408 , \31406 , \31407 );
and \g446853/U$2 ( \31409 , \12264 , RIe172f38_2685);
and \g446853/U$3 ( \31410 , RIfca99d0_6952, \12266 );
nor \g446853/U$1 ( \31411 , \31409 , \31410 );
nand \g444494/U$1 ( \31412 , \31402 , \31405 , \31408 , \31411 );
and \g452170/U$2 ( \31413 , \8317 , RIe1add68_3355);
and \g452170/U$3 ( \31414 , RIe1baef0_3504, \8326 );
nor \g452170/U$1 ( \31415 , \31413 , \31414 );
and \g446081/U$2 ( \31416 , RIe1d43f0_3792, \8340 );
and \g446081/U$3 ( \31417 , RIe19f830_3192, \8404 );
and \g448981/U$2 ( \31418 , RIe1f73a0_4190, \8523 );
and \g448981/U$3 ( \31419 , \8488 , RIe1fdfe8_4267);
and \g448981/U$4 ( \31420 , RIe1a5230_3256, \8383 );
nor \g448981/U$1 ( \31421 , \31418 , \31419 , \31420 );
and \g452171/U$2 ( \31422 , \8356 , RIe1efee8_4107);
and \g452171/U$3 ( \31423 , RIe203f88_4335, \8359 );
nor \g452171/U$1 ( \31424 , \31422 , \31423 );
and \g454926/U$2 ( \31425 , \8313 , RIe225b88_4719);
and \g454926/U$3 ( \31426 , RIe178230_2744, \8323 );
nor \g454926/U$1 ( \31427 , \31425 , \31426 );
not \g449993/U$3 ( \31428 , \31427 );
not \g449993/U$4 ( \31429 , \8376 );
and \g449993/U$2 ( \31430 , \31428 , \31429 );
and \g449993/U$5 ( \31431 , \8351 , RIe1a7f30_3288);
nor \g449993/U$1 ( \31432 , \31430 , \31431 );
and \g452812/U$2 ( \31433 , \8378 , RIe21a788_4591);
and \g452812/U$3 ( \31434 , RIe18bd30_2968, \8417 );
nor \g452812/U$1 ( \31435 , \31433 , \31434 );
nand \g447942/U$1 ( \31436 , \31421 , \31424 , \31432 , \31435 );
nor \g446081/U$1 ( \31437 , \31416 , \31417 , \31436 );
and \g452169/U$2 ( \31438 , \8335 , RIe1703a0_2654);
and \g452169/U$3 ( \31439 , RIe1a2530_3224, \8371 );
nor \g452169/U$1 ( \31440 , \31438 , \31439 );
nand \g445594/U$1 ( \31441 , \31415 , \31437 , \31440 );
and \g444876/U$2 ( \31442 , \31441 , \9010 );
and \g448980/U$2 ( \31443 , RIe1b2250_3404, \8531 );
and \g448980/U$3 ( \31444 , \8486 , RIfccdd30_7364);
and \g448980/U$4 ( \31445 , RIf14b058_5313, \8383 );
nor \g448980/U$1 ( \31446 , \31443 , \31444 , \31445 );
and \g452167/U$2 ( \31447 , \8356 , RIfec1860_8322);
and \g452167/U$3 ( \31448 , RIf148a60_5286, \8359 );
nor \g452167/U$1 ( \31449 , \31447 , \31448 );
and \g454432/U$2 ( \31450 , \8313 , RIfe89190_7904);
and \g454432/U$3 ( \31451 , RIf1499d8_5297, \8323 );
nor \g454432/U$1 ( \31452 , \31450 , \31451 );
not \g449992/U$3 ( \31453 , \31452 );
not \g449992/U$4 ( \31454 , \8376 );
and \g449992/U$2 ( \31455 , \31453 , \31454 );
and \g449992/U$5 ( \31456 , \8351 , RIfc680c0_6206);
nor \g449992/U$1 ( \31457 , \31455 , \31456 );
and \g452166/U$2 ( \31458 , \8378 , RIfec19c8_8323);
and \g452166/U$3 ( \31459 , RIfcac298_6981, \8417 );
nor \g452166/U$1 ( \31460 , \31458 , \31459 );
nand \g447719/U$1 ( \31461 , \31446 , \31449 , \31457 , \31460 );
and \g444876/U$3 ( \31462 , \8482 , \31461 );
nor \g444876/U$1 ( \31463 , \31442 , \31462 );
and \g446857/U$2 ( \31464 , \8509 , RIe1aa528_3315);
and \g446857/U$3 ( \31465 , RIe1abfe0_3334, \8511 );
nor \g446857/U$1 ( \31466 , \31464 , \31465 );
and \g446856/U$2 ( \31467 , \8514 , RIfc54728_5983);
and \g446856/U$3 ( \31468 , RIfc6e768_6279, \8517 );
nor \g446856/U$1 ( \31469 , \31467 , \31468 );
and \g446858/U$2 ( \31470 , \8969 , RIe1b6b70_3456);
and \g446858/U$3 ( \31471 , RIe1b8bc8_3479, \8971 );
nor \g446858/U$1 ( \31472 , \31470 , \31471 );
nand \g444607/U$1 ( \31473 , \31463 , \31466 , \31469 , \31472 );
and \g446077/U$2 ( \31474 , RIe201f30_4312, \8373 );
and \g446077/U$3 ( \31475 , RIf15a238_5485, \8317 );
and \g448972/U$2 ( \31476 , RIfe89460_7906, \8523 );
and \g448972/U$3 ( \31477 , \8488 , RIfe89898_7909);
and \g448972/U$4 ( \31478 , RIfceec88_7739, \8383 );
nor \g448972/U$1 ( \31479 , \31476 , \31477 , \31478 );
and \g452146/U$2 ( \31480 , \8356 , RIe1fb5b8_4237);
and \g452146/U$3 ( \31481 , RIf15f968_5547, \8359 );
nor \g452146/U$1 ( \31482 , \31480 , \31481 );
and \g454154/U$2 ( \31483 , \8313 , RIf163040_5586);
and \g454154/U$3 ( \31484 , RIf163fb8_5597, \8323 );
nor \g454154/U$1 ( \31485 , \31483 , \31484 );
not \g449986/U$3 ( \31486 , \31485 );
not \g449986/U$4 ( \31487 , \8376 );
and \g449986/U$2 ( \31488 , \31486 , \31487 );
and \g449986/U$5 ( \31489 , \8351 , RIfc6c2d8_6253);
nor \g449986/U$1 ( \31490 , \31488 , \31489 );
and \g452145/U$2 ( \31491 , \8378 , RIfe895c8_7907);
and \g452145/U$3 ( \31492 , RIf164dc8_5607, \8417 );
nor \g452145/U$1 ( \31493 , \31491 , \31492 );
nand \g447715/U$1 ( \31494 , \31479 , \31482 , \31490 , \31493 );
nor \g446077/U$1 ( \31495 , \31474 , \31475 , \31494 );
and \g452143/U$2 ( \31496 , \8335 , RIf1599c8_5479);
and \g452143/U$3 ( \31497 , RIf15c6c8_5511, \8340 );
nor \g452143/U$1 ( \31498 , \31496 , \31497 );
and \g451177/U$2 ( \31499 , \8326 , RIfe89730_7908);
and \g451177/U$3 ( \31500 , RIe200748_4295, \8404 );
nor \g451177/U$1 ( \31501 , \31499 , \31500 );
and \g445206/U$2 ( \31502 , \31495 , \31498 , \31501 );
nor \g445206/U$1 ( \31503 , \31502 , \8422 );
and \g446078/U$2 ( \31504 , RIe21d488_4623, \8407 );
and \g446078/U$3 ( \31505 , RIe214d88_4527, \8378 );
and \g448974/U$2 ( \31506 , RIe209988_4399, \8317 );
and \g448974/U$3 ( \31507 , \8326 , RIe20c688_4431);
and \g448974/U$4 ( \31508 , RIe212088_4495, \8486 );
nor \g448974/U$1 ( \31509 , \31506 , \31507 , \31508 );
and \g452152/U$2 ( \31510 , \8335 , RIe206c88_4367);
and \g452152/U$3 ( \31511 , RIf167ac8_5639, \8340 );
nor \g452152/U$1 ( \31512 , \31510 , \31511 );
and \g452151/U$2 ( \31513 , \8404 , RIe220188_4655);
and \g452151/U$3 ( \31514 , RIfc40610_5758, \8351 );
nor \g452151/U$1 ( \31515 , \31513 , \31514 );
and \g454739/U$2 ( \31516 , \8313 , RIfc5d260_6082);
and \g454739/U$3 ( \31517 , RIe222e88_4687, \8323 );
nor \g454739/U$1 ( \31518 , \31516 , \31517 );
not \g449989/U$3 ( \31519 , \31518 );
not \g449989/U$4 ( \31520 , \8328 );
and \g449989/U$2 ( \31521 , \31519 , \31520 );
and \g449989/U$5 ( \31522 , \8359 , RIfe892f8_7905);
nor \g449989/U$1 ( \31523 , \31521 , \31522 );
nand \g447716/U$1 ( \31524 , \31509 , \31512 , \31515 , \31523 );
nor \g446078/U$1 ( \31525 , \31504 , \31505 , \31524 );
and \g452150/U$2 ( \31526 , \8356 , RIe20f388_4463);
and \g452150/U$3 ( \31527 , RIfcab758_6973, \8417 );
nor \g452150/U$1 ( \31528 , \31526 , \31527 );
and \g452149/U$2 ( \31529 , \8531 , RIf168a40_5650);
and \g452149/U$3 ( \31530 , RIe217a88_4559, \8414 );
nor \g452149/U$1 ( \31531 , \31529 , \31530 );
and \g445208/U$2 ( \31532 , \31525 , \31528 , \31531 );
nor \g445208/U$1 ( \31533 , \31532 , \8368 );
or \g444368/U$1 ( \31534 , \31412 , \31473 , \31503 , \31533 );
and \g446075/U$2 ( \31535 , RIf1554e0_5430, \8409 );
and \g446075/U$3 ( \31536 , RIe1f4c40_4162, \8378 );
and \g448969/U$2 ( \31537 , RIfc5ba78_6065, \8373 );
and \g448969/U$3 ( \31538 , \8383 , RIfe89cd0_7912);
and \g448969/U$4 ( \31539 , RIfe89a00_7910, \8488 );
nor \g448969/U$1 ( \31540 , \31537 , \31538 , \31539 );
and \g452137/U$2 ( \31541 , \8335 , RIe1ed620_4078);
and \g452137/U$3 ( \31542 , RIf14f3d8_5361, \8340 );
nor \g452137/U$1 ( \31543 , \31541 , \31542 );
and \g452683/U$2 ( \31544 , \8404 , RIe1f9c68_4219);
and \g452683/U$3 ( \31545 , RIf1588e8_5467, \8351 );
nor \g452683/U$1 ( \31546 , \31544 , \31545 );
and \g454836/U$2 ( \31547 , \8313 , RIf14d920_5342);
and \g454836/U$3 ( \31548 , RIfccc818_7349, \8323 );
nor \g454836/U$1 ( \31549 , \31547 , \31548 );
not \g454835/U$1 ( \31550 , \31549 );
and \g449984/U$2 ( \31551 , \31550 , \8316 );
and \g449984/U$3 ( \31552 , RIfe89b68_7911, \8359 );
nor \g449984/U$1 ( \31553 , \31551 , \31552 );
nand \g448186/U$1 ( \31554 , \31540 , \31543 , \31546 , \31553 );
nor \g446075/U$1 ( \31555 , \31535 , \31536 , \31554 );
and \g452135/U$2 ( \31556 , \8356 , RIe1f2918_4137);
and \g452135/U$3 ( \31557 , RIfc5bd48_6067, \8417 );
nor \g452135/U$1 ( \31558 , \31556 , \31557 );
and \g452439/U$2 ( \31559 , \8531 , RIf150350_5372);
and \g452439/U$3 ( \31560 , RIf154298_5417, \8412 );
nor \g452439/U$1 ( \31561 , \31559 , \31560 );
and \g445204/U$2 ( \31562 , \31555 , \31558 , \31561 );
nor \g445204/U$1 ( \31563 , \31562 , \8621 );
and \g446076/U$2 ( \31564 , RIe1df7f0_3920, \8417 );
and \g446076/U$3 ( \31565 , RIe1c8ff0_3664, \8356 );
and \g448971/U$2 ( \31566 , RIe1c08f0_3568, \8319 );
and \g448971/U$3 ( \31567 , \8326 , RIe1c35f0_3600);
and \g448971/U$4 ( \31568 , RIe1ce9f0_3728, \8488 );
nor \g448971/U$1 ( \31569 , \31566 , \31567 , \31568 );
and \g452141/U$2 ( \31570 , \8335 , RIe1bdbf0_3536);
and \g452141/U$3 ( \31571 , RIe1c62f0_3632, \8340 );
nor \g452141/U$1 ( \31572 , \31570 , \31571 );
and \g452140/U$2 ( \31573 , \8404 , RIe1e24f0_3952);
and \g452140/U$3 ( \31574 , RIe1eabf0_4048, \8351 );
nor \g452140/U$1 ( \31575 , \31573 , \31574 );
and \g454734/U$2 ( \31576 , \8313 , RIe1e51f0_3984);
and \g454734/U$3 ( \31577 , RIe1e7ef0_4016, \8323 );
nor \g454734/U$1 ( \31578 , \31576 , \31577 );
not \g450190/U$3 ( \31579 , \31578 );
not \g450190/U$4 ( \31580 , \8328 );
and \g450190/U$2 ( \31581 , \31579 , \31580 );
and \g450190/U$5 ( \31582 , \8359 , RIe1d16f0_3760);
nor \g450190/U$1 ( \31583 , \31581 , \31582 );
nand \g447713/U$1 ( \31584 , \31569 , \31572 , \31575 , \31583 );
nor \g446076/U$1 ( \31585 , \31564 , \31565 , \31584 );
and \g452139/U$2 ( \31586 , \8378 , RIe1d70f0_3824);
and \g452139/U$3 ( \31587 , RIe1cbcf0_3696, \8531 );
nor \g452139/U$1 ( \31588 , \31586 , \31587 );
and \g452138/U$2 ( \31589 , \8414 , RIe1d9df0_3856);
and \g452138/U$3 ( \31590 , RIe1dcaf0_3888, \8409 );
nor \g452138/U$1 ( \31591 , \31589 , \31590 );
and \g445205/U$2 ( \31592 , \31585 , \31588 , \31591 );
nor \g445205/U$1 ( \31593 , \31592 , \8477 );
or \g444253/U$1 ( \31594 , \31534 , \31563 , \31593 );
_DC \g53dc/U$1 ( \31595 , \31594 , \8654 );
and \g451768/U$2 ( \31596 , \16377 , RIfccd4c0_7358);
and \g451768/U$3 ( \31597 , RIdee04f8_1016, \16380 );
nor \g451768/U$1 ( \31598 , \31596 , \31597 );
and \g446067/U$2 ( \31599 , RIfc67c88_6203, \16321 );
and \g446067/U$3 ( \31600 , RIfccb300_7334, \16313 );
and \g449014/U$2 ( \31601 , RIded6a48_906, \16398 );
and \g449014/U$3 ( \31602 , \16341 , RIded9040_933);
and \g449014/U$4 ( \31603 , RIfea8360_8230, \16485 );
nor \g449014/U$1 ( \31604 , \31601 , \31602 , \31603 );
and \g454375/U$2 ( \31605 , \16317 , RIfcac130_6980);
and \g454375/U$3 ( \31606 , RIfc6def8_6273, \16325 );
nor \g454375/U$1 ( \31607 , \31605 , \31606 );
not \g449998/U$3 ( \31608 , \31607 );
not \g449998/U$4 ( \31609 , \16351 );
and \g449998/U$2 ( \31610 , \31608 , \31609 );
and \g449998/U$5 ( \31611 , \16354 , RIfea81f8_8229);
nor \g449998/U$1 ( \31612 , \31610 , \31611 );
and \g452084/U$2 ( \31613 , \16361 , RIded26c8_858);
and \g452084/U$3 ( \31614 , RIded4b58_884, \16364 );
nor \g452084/U$1 ( \31615 , \31613 , \31614 );
and \g452062/U$2 ( \31616 , \16368 , RIfc67df0_6204);
and \g452062/U$3 ( \31617 , RIfc67b20_6202, \16371 );
nor \g452062/U$1 ( \31618 , \31616 , \31617 );
nand \g447673/U$1 ( \31619 , \31604 , \31612 , \31615 , \31618 );
nor \g446067/U$1 ( \31620 , \31599 , \31600 , \31619 );
and \g451686/U$2 ( \31621 , \16334 , RIdede338_992);
and \g451686/U$3 ( \31622 , RIfc6dc28_6271, \16326 );
nor \g451686/U$1 ( \31623 , \31621 , \31622 );
nand \g445564/U$1 ( \31624 , \31598 , \31620 , \31623 );
and \g444906/U$2 ( \31625 , \31624 , \16477 );
and \g448753/U$2 ( \31626 , RIfccde98_7365, \16427 );
and \g448753/U$3 ( \31627 , \16448 , RIfc66608_6187);
and \g448753/U$4 ( \31628 , RIdf27ad8_1828, \16485 );
nor \g448753/U$1 ( \31629 , \31626 , \31627 , \31628 );
and \g454255/U$2 ( \31630 , \16317 , RIfeaaef8_8261);
and \g454255/U$3 ( \31631 , RIfcacf40_6990, \16325 );
nor \g454255/U$1 ( \31632 , \31630 , \31631 );
not \g454254/U$1 ( \31633 , \31632 );
and \g449703/U$2 ( \31634 , \31633 , \16336 );
and \g449703/U$3 ( \31635 , RIfe8b788_7931, \16356 );
nor \g449703/U$1 ( \31636 , \31634 , \31635 );
and \g451055/U$2 ( \31637 , \16361 , RIdf18d30_1659);
and \g451055/U$3 ( \31638 , RIfc6e8d0_6280, \16364 );
nor \g451055/U$1 ( \31639 , \31637 , \31638 );
and \g451014/U$2 ( \31640 , \16368 , RIfc668d8_6189);
and \g451014/U$3 ( \31641 , RIfc66a40_6190, \16371 );
nor \g451014/U$1 ( \31642 , \31640 , \31641 );
nand \g448016/U$1 ( \31643 , \31629 , \31636 , \31639 , \31642 );
and \g444906/U$3 ( \31644 , \16481 , \31643 );
nor \g444906/U$1 ( \31645 , \31625 , \31644 );
and \g447206/U$2 ( \31646 , \16505 , RIfc6ee70_6284);
and \g447206/U$3 ( \31647 , RIee2b750_4953, \16507 );
nor \g447206/U$1 ( \31648 , \31646 , \31647 );
and \g446555/U$2 ( \31649 , \16511 , RIdf24130_1787);
and \g446555/U$3 ( \31650 , RIdf25d50_1807, \16514 );
nor \g446555/U$1 ( \31651 , \31649 , \31650 );
and \g446511/U$2 ( \31652 , \16518 , RIee27808_4908);
and \g446511/U$3 ( \31653 , RIfc6efd8_6285, \16521 );
nor \g446511/U$1 ( \31654 , \31652 , \31653 );
nand \g444655/U$1 ( \31655 , \31645 , \31648 , \31651 , \31654 );
and \g453121/U$2 ( \31656 , \16377 , RIdec7700_733);
and \g453121/U$3 ( \31657 , RIe16d808_2623, \16380 );
nor \g453121/U$1 ( \31658 , \31656 , \31657 );
and \g446288/U$2 ( \31659 , RIdecd100_797, \16319 );
and \g446288/U$3 ( \31660 , RIdeca400_765, \16313 );
and \g449364/U$2 ( \31661 , RIdf377f8_2008, \16427 );
and \g449364/U$3 ( \31662 , \16448 , RIe142e00_2138);
and \g449364/U$4 ( \31663 , RIde95228_317, \16344 );
nor \g449364/U$1 ( \31664 , \31661 , \31662 , \31663 );
and \g455334/U$2 ( \31665 , \16317 , RIdee68d0_1087);
and \g455334/U$3 ( \31666 , RIdeffdd0_1375, \16325 );
nor \g455334/U$1 ( \31667 , \31665 , \31666 );
not \g455333/U$1 ( \31668 , \31667 );
and \g450325/U$2 ( \31669 , \31668 , \16336 );
and \g450325/U$3 ( \31670 , RIdeb3c00_509, \16356 );
nor \g450325/U$1 ( \31671 , \31669 , \31670 );
and \g453333/U$2 ( \31672 , \16361 , RIde7b170_190);
and \g453333/U$3 ( \31673 , RIdedb638_960, \16364 );
nor \g453333/U$1 ( \31674 , \31672 , \31673 );
and \g453291/U$2 ( \31675 , \16368 , RIdf1c6d8_1700);
and \g453291/U$3 ( \31676 , RIdf2be58_1876, \16371 );
nor \g453291/U$1 ( \31677 , \31675 , \31676 );
nand \g448100/U$1 ( \31678 , \31664 , \31671 , \31674 , \31677 );
nor \g446288/U$1 ( \31679 , \31659 , \31660 , \31678 );
and \g453083/U$2 ( \31680 , \16334 , RIe159600_2394);
and \g453083/U$3 ( \31681 , RIdecfe00_829, \16328 );
nor \g453083/U$1 ( \31682 , \31680 , \31681 );
nand \g445643/U$1 ( \31683 , \31658 , \31679 , \31682 );
and \g444866/U$2 ( \31684 , \31683 , \16752 );
and \g449215/U$2 ( \31685 , RIdefa3d0_1311, \16427 );
and \g449215/U$3 ( \31686 , \16448 , RIdefd0d0_1343);
and \g449215/U$4 ( \31687 , RIdf084d0_1471, \16344 );
nor \g449215/U$1 ( \31688 , \31685 , \31686 , \31687 );
and \g455064/U$2 ( \31689 , \16317 , RIdeeefd0_1183);
and \g455064/U$3 ( \31690 , RIdef1cd0_1215, \16325 );
nor \g455064/U$1 ( \31691 , \31689 , \31690 );
not \g455063/U$1 ( \31692 , \31691 );
and \g450177/U$2 ( \31693 , \31692 , \16336 );
and \g450177/U$3 ( \31694 , RIdf0b1d0_1503, \16356 );
nor \g450177/U$1 ( \31695 , \31693 , \31694 );
and \g452715/U$2 ( \31696 , \16361 , RIdee95d0_1119);
and \g452715/U$3 ( \31697 , RIdeec2d0_1151, \16364 );
nor \g452715/U$1 ( \31698 , \31696 , \31697 );
and \g452693/U$2 ( \31699 , \16368 , RIdef49d0_1247);
and \g452693/U$3 ( \31700 , RIdef76d0_1279, \16371 );
nor \g452693/U$1 ( \31701 , \31699 , \31700 );
nand \g448086/U$1 ( \31702 , \31688 , \31695 , \31698 , \31701 );
and \g444866/U$3 ( \31703 , \16750 , \31702 );
nor \g444866/U$1 ( \31704 , \31684 , \31703 );
and \g446909/U$2 ( \31705 , \19457 , RIdf138d0_1599);
and \g446909/U$3 ( \31706 , RIdf165d0_1631, \19459 );
nor \g446909/U$1 ( \31707 , \31705 , \31706 );
and \g446935/U$2 ( \31708 , \19462 , RIdf02ad0_1407);
and \g446935/U$3 ( \31709 , RIdf057d0_1439, \19464 );
nor \g446935/U$1 ( \31710 , \31708 , \31709 );
and \g446925/U$2 ( \31711 , \19467 , RIdf0ded0_1535);
and \g446925/U$3 ( \31712 , RIdf10bd0_1567, \19469 );
nor \g446925/U$1 ( \31713 , \31711 , \31712 );
nand \g444617/U$1 ( \31714 , \31704 , \31707 , \31710 , \31713 );
and \g446070/U$2 ( \31715 , RIfc6fc80_6294, \16326 );
and \g446070/U$3 ( \31716 , RIfe8b8f0_7932, \16377 );
and \g449092/U$2 ( \31717 , RIfcad210_6992, \16427 );
and \g449092/U$3 ( \31718 , \16448 , RIfc65ac8_6179);
and \g449092/U$4 ( \31719 , RIde8c510_274, \16344 );
nor \g449092/U$1 ( \31720 , \31717 , \31718 , \31719 );
and \g454232/U$2 ( \31721 , \16317 , RIe16af40_2594);
and \g454232/U$3 ( \31722 , RIfc51488_5947, \16325 );
nor \g454232/U$1 ( \31723 , \31721 , \31722 );
not \g454231/U$1 ( \31724 , \31723 );
and \g450059/U$2 ( \31725 , \31724 , \16336 );
and \g450059/U$3 ( \31726 , RIde90020_292, \16356 );
nor \g450059/U$1 ( \31727 , \31725 , \31726 );
and \g452300/U$2 ( \31728 , \16361 , RIe167598_2553);
and \g452300/U$3 ( \31729 , RIfc65c30_6180, \16364 );
nor \g452300/U$1 ( \31730 , \31728 , \31729 );
and \g452185/U$2 ( \31731 , \16368 , RIfcce2d0_7368);
and \g452185/U$3 ( \31732 , RIfcce168_7367, \16371 );
nor \g452185/U$1 ( \31733 , \31731 , \31732 );
nand \g448062/U$1 ( \31734 , \31720 , \31727 , \31730 , \31733 );
nor \g446070/U$1 ( \31735 , \31715 , \31716 , \31734 );
and \g451595/U$2 ( \31736 , \16334 , RIde84ba8_237);
and \g451595/U$3 ( \31737 , RIfca8080_6934, \16313 );
nor \g451595/U$1 ( \31738 , \31736 , \31737 );
and \g451552/U$2 ( \31739 , \16380 , RIde89090_258);
and \g451552/U$3 ( \31740 , RIee1b760_4771, \16321 );
nor \g451552/U$1 ( \31741 , \31739 , \31740 );
and \g445084/U$2 ( \31742 , \31735 , \31738 , \31741 );
nor \g445084/U$1 ( \31743 , \31742 , \16649 );
and \g446283/U$2 ( \31744 , RIdec4a00_701, \16326 );
and \g446283/U$3 ( \31745 , RIdebf000_637, \16377 );
and \g449378/U$2 ( \31746 , RIdea8d28_413, \16398 );
and \g449378/U$3 ( \31747 , \16341 , RIfce69c0_7646);
and \g449378/U$4 ( \31748 , RIdebc300_605, \16485 );
nor \g449378/U$1 ( \31749 , \31746 , \31747 , \31748 );
and \g455153/U$2 ( \31750 , \16317 , RIdeb0f00_477);
and \g455153/U$3 ( \31751 , RIfc6f9b0_6292, \16325 );
nor \g455153/U$1 ( \31752 , \31750 , \31751 );
not \g450373/U$3 ( \31753 , \31752 );
not \g450373/U$4 ( \31754 , \16351 );
and \g450373/U$2 ( \31755 , \31753 , \31754 );
and \g450373/U$5 ( \31756 , \16356 , RIfc64cb8_6169);
nor \g450373/U$1 ( \31757 , \31755 , \31756 );
and \g453395/U$2 ( \31758 , \16361 , RIde9bb28_349);
and \g453395/U$3 ( \31759 , RIdea2428_381, \16364 );
nor \g453395/U$1 ( \31760 , \31758 , \31759 );
and \g453312/U$2 ( \31761 , \16368 , RIdeae200_445);
and \g453312/U$3 ( \31762 , RIfc657f8_6177, \16371 );
nor \g453312/U$1 ( \31763 , \31761 , \31762 );
nand \g447880/U$1 ( \31764 , \31749 , \31757 , \31760 , \31763 );
nor \g446283/U$1 ( \31765 , \31744 , \31745 , \31764 );
and \g453029/U$2 ( \31766 , \16334 , RIdeb6900_541);
and \g453029/U$3 ( \31767 , RIfcad7b0_6996, \16313 );
nor \g453029/U$1 ( \31768 , \31766 , \31767 );
and \g452881/U$2 ( \31769 , \16380 , RIdeb9600_573);
and \g452881/U$3 ( \31770 , RIdec1d00_669, \16321 );
nor \g452881/U$1 ( \31771 , \31769 , \31770 );
and \g445296/U$2 ( \31772 , \31765 , \31768 , \31771 );
nor \g445296/U$1 ( \31773 , \31772 , \16618 );
or \g444382/U$1 ( \31774 , \31655 , \31714 , \31743 , \31773 );
and \g446157/U$2 ( \31775 , RIee33fb8_5050, \16328 );
and \g446157/U$3 ( \31776 , RIee30fe8_5016, \16377 );
and \g448895/U$2 ( \31777 , RIfcac6d0_6984, \16427 );
and \g448895/U$3 ( \31778 , \16432 , RIfc6e060_6274);
and \g448895/U$4 ( \31779 , RIdf3e5a8_2086, \16485 );
nor \g448895/U$1 ( \31780 , \31777 , \31778 , \31779 );
and \g454673/U$2 ( \31781 , \16317 , RIdf32d70_1955);
and \g454673/U$3 ( \31782 , RIdf34dc8_1978, \16325 );
nor \g454673/U$1 ( \31783 , \31781 , \31782 );
not \g454672/U$1 ( \31784 , \31783 );
and \g449697/U$2 ( \31785 , \31784 , \16336 );
and \g449697/U$3 ( \31786 , RIfea8630_8232, \16356 );
nor \g449697/U$1 ( \31787 , \31785 , \31786 );
and \g453498/U$2 ( \31788 , \16361 , RIdf2eb58_1908);
and \g453498/U$3 ( \31789 , RIfea84c8_8231, \16364 );
nor \g453498/U$1 ( \31790 , \31788 , \31789 );
and \g453165/U$2 ( \31791 , \16368 , RIfc6e600_6278);
and \g453165/U$3 ( \31792 , RIfc56078_6001, \16371 );
nor \g453165/U$1 ( \31793 , \31791 , \31792 );
nand \g448102/U$1 ( \31794 , \31780 , \31787 , \31790 , \31793 );
nor \g446157/U$1 ( \31795 , \31775 , \31776 , \31794 );
and \g450961/U$2 ( \31796 , \16334 , RIfea8798_8233);
and \g450961/U$3 ( \31797 , RIee31c90_5025, \16313 );
nor \g450961/U$1 ( \31798 , \31796 , \31797 );
and \g450855/U$2 ( \31799 , \16380 , RIdf3c550_2063);
and \g450855/U$3 ( \31800 , RIee32d70_5037, \16321 );
nor \g450855/U$1 ( \31801 , \31799 , \31800 );
and \g445453/U$2 ( \31802 , \31795 , \31798 , \31801 );
nor \g445453/U$1 ( \31803 , \31802 , \16393 );
and \g446185/U$2 ( \31804 , RIe161d00_2490, \16321 );
and \g446185/U$3 ( \31805 , RIfc66e78_6193, \16313 );
and \g448503/U$2 ( \31806 , RIe14b500_2234, \16398 );
and \g448503/U$3 ( \31807 , \16341 , RIfc6e1c8_6275);
and \g448503/U$4 ( \31808 , RIe15c300_2426, \16485 );
nor \g448503/U$1 ( \31809 , \31806 , \31807 , \31808 );
and \g454152/U$2 ( \31810 , \16317 , RIe150f00_2298);
and \g454152/U$3 ( \31811 , RIfc6e330_6276, \16325 );
nor \g454152/U$1 ( \31812 , \31810 , \31811 );
not \g450486/U$3 ( \31813 , \31812 );
not \g450486/U$4 ( \31814 , \16351 );
and \g450486/U$2 ( \31815 , \31813 , \31814 );
and \g450486/U$5 ( \31816 , \16356 , RIfc6e498_6277);
nor \g450486/U$1 ( \31817 , \31815 , \31816 );
and \g453602/U$2 ( \31818 , \16361 , RIe145b00_2170);
and \g453602/U$3 ( \31819 , RIe148800_2202, \16364 );
nor \g453602/U$1 ( \31820 , \31818 , \31819 );
and \g453535/U$2 ( \31821 , \16368 , RIe14e200_2266);
and \g453535/U$3 ( \31822 , RIfccda60_7362, \16371 );
nor \g453535/U$1 ( \31823 , \31821 , \31822 );
nand \g447969/U$1 ( \31824 , \31809 , \31817 , \31820 , \31823 );
nor \g446185/U$1 ( \31825 , \31804 , \31805 , \31824 );
and \g452946/U$2 ( \31826 , \16377 , RIe15f000_2458);
and \g452946/U$3 ( \31827 , RIe156900_2362, \16380 );
nor \g452946/U$1 ( \31828 , \31826 , \31827 );
and \g452772/U$2 ( \31829 , \16334 , RIe153c00_2330);
and \g452772/U$3 ( \31830 , RIe164a00_2522, \16328 );
nor \g452772/U$1 ( \31831 , \31829 , \31830 );
and \g445277/U$2 ( \31832 , \31825 , \31828 , \31831 );
nor \g445277/U$1 ( \31833 , \31832 , \16389 );
or \g444219/U$1 ( \31834 , \31774 , \31803 , \31833 );
_DC \g5461/U$1 ( \31835 , \31834 , \16652 );
and \g449105/U$2 ( \31836 , RIfcc9b18_7317, \8373 );
and \g449105/U$3 ( \31837 , \8383 , RIfca6a00_6918);
and \g449105/U$4 ( \31838 , RIee3ad68_5128, \8488 );
nor \g449105/U$1 ( \31839 , \31836 , \31837 , \31838 );
and \g454920/U$2 ( \31840 , \8313 , RIfccf7e8_7383);
and \g454920/U$3 ( \31841 , RIfc726b0_6324, \8323 );
nor \g454920/U$1 ( \31842 , \31840 , \31841 );
not \g450107/U$3 ( \31843 , \31842 );
not \g450107/U$4 ( \31844 , \8376 );
and \g450107/U$2 ( \31845 , \31843 , \31844 );
and \g450107/U$5 ( \31846 , \8359 , RIee3be48_5140);
nor \g450107/U$1 ( \31847 , \31845 , \31846 );
and \g452522/U$2 ( \31848 , \8404 , RIe175530_2712);
and \g452522/U$3 ( \31849 , RIfcaf268_7015, \8351 );
nor \g452522/U$1 ( \31850 , \31848 , \31849 );
and \g452540/U$2 ( \31851 , \8378 , RIfc72548_6323);
and \g452540/U$3 ( \31852 , RIfc72818_6325, \8417 );
nor \g452540/U$1 ( \31853 , \31851 , \31852 );
nand \g447769/U$1 ( \31854 , \31839 , \31847 , \31850 , \31853 );
and \g444687/U$2 ( \31855 , \31854 , \9700 );
and \g446225/U$2 ( \31856 , RIfc72278_6321, \8531 );
and \g446225/U$3 ( \31857 , RIe17dd98_2809, \8319 );
and \g449190/U$2 ( \31858 , RIfc73088_6331, \8371 );
and \g449190/U$3 ( \31859 , \8383 , RIe199f98_3129);
and \g449190/U$4 ( \31860 , RIe186498_2905, \8486 );
nor \g449190/U$1 ( \31861 , \31858 , \31859 , \31860 );
and \g455090/U$2 ( \31862 , \8313 , RIe191898_3033);
and \g455090/U$3 ( \31863 , RIe194598_3065, \8323 );
nor \g455090/U$1 ( \31864 , \31862 , \31863 );
not \g450195/U$3 ( \31865 , \31864 );
not \g450195/U$4 ( \31866 , \8376 );
and \g450195/U$2 ( \31867 , \31865 , \31866 );
and \g450195/U$5 ( \31868 , \8359 , RIe189198_2937);
nor \g450195/U$1 ( \31869 , \31867 , \31868 );
and \g452822/U$2 ( \31870 , \8404 , RIe197298_3097);
and \g452822/U$3 ( \31871 , RIe19cc98_3161, \8351 );
nor \g452822/U$1 ( \31872 , \31870 , \31871 );
and \g452846/U$2 ( \31873 , \8378 , RIe18eb98_3001);
and \g452846/U$3 ( \31874 , RIf1442a8_5235, \8417 );
nor \g452846/U$1 ( \31875 , \31873 , \31874 );
nand \g447803/U$1 ( \31876 , \31861 , \31869 , \31872 , \31875 );
nor \g446225/U$1 ( \31877 , \31856 , \31857 , \31876 );
and \g452716/U$2 ( \31878 , \8335 , RIe17b098_2777);
and \g452716/U$3 ( \31879 , RIfc61ce8_6135, \8340 );
nor \g452716/U$1 ( \31880 , \31878 , \31879 );
and \g452699/U$2 ( \31881 , \8326 , RIe180a98_2841);
and \g452699/U$3 ( \31882 , RIe183798_2873, \8356 );
nor \g452699/U$1 ( \31883 , \31881 , \31882 );
and \g445284/U$2 ( \31884 , \31877 , \31880 , \31883 );
nor \g445284/U$1 ( \31885 , \31884 , \8589 );
nor \g444687/U$1 ( \31886 , \31855 , \31885 );
and \g446910/U$2 ( \31887 , \10044 , RIfc62120_6138);
and \g446910/U$3 ( \31888 , RIfc71e40_6318, \10046 );
nor \g446910/U$1 ( \31889 , \31887 , \31888 );
and \g446903/U$2 ( \31890 , \10034 , RIfccf518_7381);
and \g446903/U$3 ( \31891 , RIfcaef98_7013, \10036 );
nor \g446903/U$1 ( \31892 , \31890 , \31891 );
and \g446918/U$2 ( \31893 , \12264 , RIe1730a0_2686);
and \g446918/U$3 ( \31894 , RIfc71fa8_6319, \12266 );
nor \g446918/U$1 ( \31895 , \31893 , \31894 );
nand \g444500/U$1 ( \31896 , \31886 , \31889 , \31892 , \31895 );
and \g453346/U$2 ( \31897 , \8404 , RIe19f998_3193);
and \g453346/U$3 ( \31898 , RIe178398_2745, \8409 );
nor \g453346/U$1 ( \31899 , \31897 , \31898 );
and \g446323/U$2 ( \31900 , RIe1a2698_3225, \8373 );
and \g446323/U$3 ( \31901 , RIe21a8f0_4592, \8378 );
and \g449342/U$2 ( \31902 , RIe1aded0_3356, \8319 );
and \g449342/U$3 ( \31903 , \8326 , RIe1bb058_3505);
and \g449342/U$4 ( \31904 , RIe1a5398_3257, \8383 );
nor \g449342/U$1 ( \31905 , \31902 , \31903 , \31904 );
and \g453486/U$2 ( \31906 , \8335 , RIe170508_2655);
and \g453486/U$3 ( \31907 , RIe1d4558_3793, \8340 );
nor \g453486/U$1 ( \31908 , \31906 , \31907 );
and \g454162/U$2 ( \31909 , \8313 , RIe1f7508_4191);
and \g454162/U$3 ( \31910 , RIe1fe150_4268, \8323 );
nor \g454162/U$1 ( \31911 , \31909 , \31910 );
not \g450358/U$3 ( \31912 , \31911 );
not \g450358/U$4 ( \31913 , \8347 );
and \g450358/U$2 ( \31914 , \31912 , \31913 );
and \g450358/U$5 ( \31915 , \8351 , RIe1a8098_3289);
nor \g450358/U$1 ( \31916 , \31914 , \31915 );
and \g453418/U$2 ( \31917 , \8356 , RIe1f0050_4108);
and \g453418/U$3 ( \31918 , RIe2040f0_4336, \8359 );
nor \g453418/U$1 ( \31919 , \31917 , \31918 );
nand \g447924/U$1 ( \31920 , \31905 , \31908 , \31916 , \31919 );
nor \g446323/U$1 ( \31921 , \31900 , \31901 , \31920 );
and \g453320/U$2 ( \31922 , \8412 , RIe225cf0_4720);
and \g453320/U$3 ( \31923 , RIe18be98_2969, \8417 );
nor \g453320/U$1 ( \31924 , \31922 , \31923 );
nand \g445657/U$1 ( \31925 , \31899 , \31921 , \31924 );
and \g444882/U$2 ( \31926 , \31925 , \9010 );
and \g449277/U$2 ( \31927 , RIfeaac28_8259, \8317 );
and \g449277/U$3 ( \31928 , \8326 , RIfc700b8_6297);
and \g449277/U$4 ( \31929 , RIf14b1c0_5314, \8383 );
nor \g449277/U$1 ( \31930 , \31927 , \31928 , \31929 );
and \g453182/U$2 ( \31931 , \8335 , RIe1aa690_3316);
and \g453182/U$3 ( \31932 , RIfc645b0_6164, \8340 );
nor \g453182/U$1 ( \31933 , \31931 , \31932 );
and \g454529/U$2 ( \31934 , \8313 , RIe1b23b8_3405);
and \g454529/U$3 ( \31935 , RIfcce870_7372, \8323 );
nor \g454529/U$1 ( \31936 , \31934 , \31935 );
not \g450282/U$3 ( \31937 , \31936 );
not \g450282/U$4 ( \31938 , \8347 );
and \g450282/U$2 ( \31939 , \31937 , \31938 );
and \g450282/U$5 ( \31940 , \8351 , RIf14c408_5327);
nor \g450282/U$1 ( \31941 , \31939 , \31940 );
and \g453155/U$2 ( \31942 , \8356 , RIe1b0630_3384);
and \g453155/U$3 ( \31943 , RIfc70220_6298, \8359 );
nor \g453155/U$1 ( \31944 , \31942 , \31943 );
nand \g447856/U$1 ( \31945 , \31930 , \31933 , \31941 , \31944 );
and \g444882/U$3 ( \31946 , \8482 , \31945 );
nor \g444882/U$1 ( \31947 , \31926 , \31946 );
and \g447023/U$2 ( \31948 , \8964 , RIfca7c48_6931);
and \g447023/U$3 ( \31949 , RIfc707c0_6302, \8966 );
nor \g447023/U$1 ( \31950 , \31948 , \31949 );
and \g447039/U$2 ( \31951 , \8969 , RIe1b6cd8_3457);
and \g447039/U$3 ( \31952 , RIe1b8d30_3480, \8971 );
nor \g447039/U$1 ( \31953 , \31951 , \31952 );
and \g447047/U$2 ( \31954 , \8974 , RIe1b3a38_3421);
and \g447047/U$3 ( \31955 , RIe1b4de8_3435, \8976 );
nor \g447047/U$1 ( \31956 , \31954 , \31955 );
nand \g444628/U$1 ( \31957 , \31947 , \31950 , \31953 , \31956 );
and \g445947/U$2 ( \31958 , RIfcc9f50_7320, \8373 );
and \g445947/U$3 ( \31959 , RIe214ef0_4528, \8378 );
and \g448917/U$2 ( \31960 , RIf168ba8_5651, \8531 );
and \g448917/U$3 ( \31961 , \8488 , RIe2121f0_4496);
and \g448917/U$4 ( \31962 , RIe222ff0_4688, \8383 );
nor \g448917/U$1 ( \31963 , \31960 , \31961 , \31962 );
and \g451833/U$2 ( \31964 , \8335 , RIe206df0_4368);
and \g451833/U$3 ( \31965 , RIfc71300_6310, \8340 );
nor \g451833/U$1 ( \31966 , \31964 , \31965 );
and \g454492/U$2 ( \31967 , \8313 , RIe209af0_4400);
and \g454492/U$3 ( \31968 , RIe20c7f0_4432, \8323 );
nor \g454492/U$1 ( \31969 , \31967 , \31968 );
not \g454491/U$1 ( \31970 , \31969 );
and \g449906/U$2 ( \31971 , \31970 , \8316 );
and \g449906/U$3 ( \31972 , RIfe8b350_7928, \8351 );
nor \g449906/U$1 ( \31973 , \31971 , \31972 );
and \g451791/U$2 ( \31974 , \8356 , RIe20f4f0_4464);
and \g451791/U$3 ( \31975 , RIfccf3b0_7380, \8359 );
nor \g451791/U$1 ( \31976 , \31974 , \31975 );
nand \g448170/U$1 ( \31977 , \31963 , \31966 , \31973 , \31976 );
nor \g445947/U$1 ( \31978 , \31958 , \31959 , \31977 );
and \g451650/U$2 ( \31979 , \8404 , RIe2202f0_4656);
and \g451650/U$3 ( \31980 , RIe21d5f0_4624, \8409 );
nor \g451650/U$1 ( \31981 , \31979 , \31980 );
and \g451601/U$2 ( \31982 , \8414 , RIe217bf0_4560);
and \g451601/U$3 ( \31983 , RIfc4a570_5868, \8417 );
nor \g451601/U$1 ( \31984 , \31982 , \31983 );
and \g445089/U$2 ( \31985 , \31978 , \31981 , \31984 );
nor \g445089/U$1 ( \31986 , \31985 , \8368 );
and \g446102/U$2 ( \31987 , RIe1fc698_4249, \8531 );
and \g446102/U$3 ( \31988 , RIfc63200_6150, \8319 );
and \g449030/U$2 ( \31989 , RIe202098_4313, \8373 );
and \g449030/U$3 ( \31990 , \8383 , RIfc71a08_6315);
and \g449030/U$4 ( \31991 , RIf15dbe0_5526, \8488 );
nor \g449030/U$1 ( \31992 , \31989 , \31990 , \31991 );
and \g454339/U$2 ( \31993 , \8313 , RIfc62c60_6146);
and \g454339/U$3 ( \31994 , RIfce6588_7643, \8323 );
nor \g454339/U$1 ( \31995 , \31993 , \31994 );
not \g450030/U$3 ( \31996 , \31995 );
not \g450030/U$4 ( \31997 , \8376 );
and \g450030/U$2 ( \31998 , \31996 , \31997 );
and \g450030/U$5 ( \31999 , \8359 , RIf15fad0_5548);
nor \g450030/U$1 ( \32000 , \31998 , \31999 );
and \g452240/U$2 ( \32001 , \8404 , RIfe8b1e8_7927);
and \g452240/U$3 ( \32002 , RIfc718a0_6314, \8351 );
nor \g452240/U$1 ( \32003 , \32001 , \32002 );
and \g452287/U$2 ( \32004 , \8378 , RIf161858_5569);
and \g452287/U$3 ( \32005 , RIfc715d0_6312, \8417 );
nor \g452287/U$1 ( \32006 , \32004 , \32005 );
nand \g447724/U$1 ( \32007 , \31992 , \32000 , \32003 , \32006 );
nor \g446102/U$1 ( \32008 , \31987 , \31988 , \32007 );
and \g452118/U$2 ( \32009 , \8335 , RIfc71198_6309);
and \g452118/U$3 ( \32010 , RIfcae5c0_7006, \8340 );
nor \g452118/U$1 ( \32011 , \32009 , \32010 );
and \g452094/U$2 ( \32012 , \8326 , RIfc63098_6149);
and \g452094/U$3 ( \32013 , RIfe8b4b8_7929, \8356 );
nor \g452094/U$1 ( \32014 , \32012 , \32013 );
and \g445198/U$2 ( \32015 , \32008 , \32011 , \32014 );
nor \g445198/U$1 ( \32016 , \32015 , \8422 );
or \g444370/U$1 ( \32017 , \31896 , \31957 , \31986 , \32016 );
and \g446486/U$2 ( \32018 , RIfc4d108_5899, \8531 );
and \g446486/U$3 ( \32019 , RIfca7810_6928, \8319 );
and \g448581/U$2 ( \32020 , RIf154400_5418, \8414 );
and \g448581/U$3 ( \32021 , \8409 , RIfcceb40_7374);
and \g448581/U$4 ( \32022 , RIf151868_5387, \8486 );
nor \g448581/U$1 ( \32023 , \32020 , \32021 , \32022 );
and \g454264/U$2 ( \32024 , \8313 , RIfcdc808_7531);
and \g454264/U$3 ( \32025 , RIf1576a0_5454, \8323 );
nor \g454264/U$1 ( \32026 , \32024 , \32025 );
not \g449576/U$3 ( \32027 , \32026 );
not \g449576/U$4 ( \32028 , \8328 );
and \g449576/U$2 ( \32029 , \32027 , \32028 );
and \g449576/U$5 ( \32030 , \8359 , RIf152c18_5401);
nor \g449576/U$1 ( \32031 , \32029 , \32030 );
and \g450591/U$2 ( \32032 , \8404 , RIfe8b620_7930);
and \g450591/U$3 ( \32033 , RIf158a50_5468, \8351 );
nor \g450591/U$1 ( \32034 , \32032 , \32033 );
and \g450675/U$2 ( \32035 , \8378 , RIe1f4da8_4163);
and \g450675/U$3 ( \32036 , RIfc634d0_6152, \8417 );
nor \g450675/U$1 ( \32037 , \32035 , \32036 );
nand \g447456/U$1 ( \32038 , \32023 , \32031 , \32034 , \32037 );
nor \g446486/U$1 ( \32039 , \32018 , \32019 , \32038 );
and \g453963/U$2 ( \32040 , \8335 , RIe1ed788_4079);
and \g453963/U$3 ( \32041 , RIfc70a90_6304, \8340 );
nor \g453963/U$1 ( \32042 , \32040 , \32041 );
and \g453800/U$2 ( \32043 , \8326 , RIfc63bd8_6157);
and \g453800/U$3 ( \32044 , RIe1f2a80_4138, \8356 );
nor \g453800/U$1 ( \32045 , \32043 , \32044 );
and \g445422/U$2 ( \32046 , \32039 , \32042 , \32045 );
nor \g445422/U$1 ( \32047 , \32046 , \8621 );
and \g445816/U$2 ( \32048 , RIe1c9158_3665, \8356 );
and \g445816/U$3 ( \32049 , RIe1d1858_3761, \8359 );
and \g448746/U$2 ( \32050 , RIe1d9f58_3857, \8412 );
and \g448746/U$3 ( \32051 , \8409 , RIe1dcc58_3889);
and \g448746/U$4 ( \32052 , RIe1c3758_3601, \8324 );
nor \g448746/U$1 ( \32053 , \32050 , \32051 , \32052 );
and \g454647/U$2 ( \32054 , \8313 , RIe1e5358_3985);
and \g454647/U$3 ( \32055 , RIe1e8058_4017, \8323 );
nor \g454647/U$1 ( \32056 , \32054 , \32055 );
not \g449748/U$3 ( \32057 , \32056 );
not \g449748/U$4 ( \32058 , \8328 );
and \g449748/U$2 ( \32059 , \32057 , \32058 );
and \g449748/U$5 ( \32060 , \8340 , RIe1c6458_3633);
nor \g449748/U$1 ( \32061 , \32059 , \32060 );
and \g451217/U$2 ( \32062 , \8404 , RIe1e2658_3953);
and \g451217/U$3 ( \32063 , RIe1ead58_4049, \8351 );
nor \g451217/U$1 ( \32064 , \32062 , \32063 );
and \g451296/U$2 ( \32065 , \8378 , RIe1d7258_3825);
and \g451296/U$3 ( \32066 , RIe1df958_3921, \8417 );
nor \g451296/U$1 ( \32067 , \32065 , \32066 );
nand \g447553/U$1 ( \32068 , \32053 , \32061 , \32064 , \32067 );
nor \g445816/U$1 ( \32069 , \32048 , \32049 , \32068 );
and \g451082/U$2 ( \32070 , \8335 , RIe1bdd58_3537);
and \g451082/U$3 ( \32071 , RIe1ceb58_3729, \8486 );
nor \g451082/U$1 ( \32072 , \32070 , \32071 );
and \g451037/U$2 ( \32073 , \8319 , RIe1c0a58_3569);
and \g451037/U$3 ( \32074 , RIe1cbe58_3697, \8531 );
nor \g451037/U$1 ( \32075 , \32073 , \32074 );
and \g444991/U$2 ( \32076 , \32069 , \32072 , \32075 );
nor \g444991/U$1 ( \32077 , \32076 , \8477 );
or \g444255/U$1 ( \32078 , \32017 , \32047 , \32077 );
_DC \g54e5/U$1 ( \32079 , \32078 , \8654 );
and \g452897/U$2 ( \32080 , \16380 , RIdee0660_1017);
and \g452897/U$3 ( \32081 , RIfccfd88_7387, \16321 );
nor \g452897/U$1 ( \32082 , \32080 , \32081 );
and \g446235/U$2 ( \32083 , RIfcc96e0_7314, \16328 );
and \g446235/U$3 ( \32084 , RIfca5ec0_6910, \16377 );
and \g449195/U$2 ( \32085 , RIded6bb0_907, \16398 );
and \g449195/U$3 ( \32086 , \16339 , RIfe82980_7830);
and \g449195/U$4 ( \32087 , RIdee2550_1039, \16485 );
nor \g449195/U$1 ( \32088 , \32085 , \32086 , \32087 );
and \g454991/U$2 ( \32089 , \16317 , RIfc73bc8_6339);
and \g454991/U$3 ( \32090 , RIfcdeb30_7556, \16325 );
nor \g454991/U$1 ( \32091 , \32089 , \32090 );
not \g450205/U$3 ( \32092 , \32091 );
not \g450205/U$4 ( \32093 , \16351 );
and \g450205/U$2 ( \32094 , \32092 , \32093 );
and \g450205/U$5 ( \32095 , \16354 , RIdee45a8_1062);
nor \g450205/U$1 ( \32096 , \32094 , \32095 );
and \g452928/U$2 ( \32097 , \16361 , RIded2830_859);
and \g452928/U$3 ( \32098 , RIded4cc0_885, \16364 );
nor \g452928/U$1 ( \32099 , \32097 , \32098 );
and \g452915/U$2 ( \32100 , \16368 , RIfc73a60_6338);
and \g452915/U$3 ( \32101 , RIfca5bf0_6908, \16371 );
nor \g452915/U$1 ( \32102 , \32100 , \32101 );
nand \g447818/U$1 ( \32103 , \32088 , \32096 , \32099 , \32102 );
nor \g446235/U$1 ( \32104 , \32083 , \32084 , \32103 );
and \g452903/U$2 ( \32105 , \16334 , RIfe826b0_7828);
and \g452903/U$3 ( \32106 , RIfc60aa0_6122, \16313 );
nor \g452903/U$1 ( \32107 , \32105 , \32106 );
nand \g445637/U$1 ( \32108 , \32082 , \32104 , \32107 );
and \g444920/U$2 ( \32109 , \32108 , \16477 );
and \g449180/U$2 ( \32110 , RIde95570_318, \16344 );
and \g449180/U$3 ( \32111 , \16356 , RIdeb3d68_510);
and \g449180/U$4 ( \32112 , RIdee6a38_1088, \16337 );
nor \g449180/U$1 ( \32113 , \32110 , \32111 , \32112 );
and \g455073/U$2 ( \32114 , \16317 , RIdecd268_798);
and \g455073/U$3 ( \32115 , RIdecff68_830, \16325 );
nor \g455073/U$1 ( \32116 , \32114 , \32115 );
not \g450189/U$3 ( \32117 , \32116 );
not \g450189/U$4 ( \32118 , \16311 );
and \g450189/U$2 ( \32119 , \32117 , \32118 );
and \g450189/U$5 ( \32120 , \16341 , RIdefff38_1376);
nor \g450189/U$1 ( \32121 , \32119 , \32120 );
and \g452871/U$2 ( \32122 , \16377 , RIdec7868_734);
and \g452871/U$3 ( \32123 , RIdeca568_766, \16313 );
nor \g452871/U$1 ( \32124 , \32122 , \32123 );
and \g452878/U$2 ( \32125 , \16334 , RIe159768_2395);
and \g452878/U$3 ( \32126 , RIe16d970_2624, \16380 );
nor \g452878/U$1 ( \32127 , \32125 , \32126 );
nand \g447387/U$1 ( \32128 , \32113 , \32121 , \32124 , \32127 );
and \g444920/U$3 ( \32129 , \16752 , \32128 );
nor \g444920/U$1 ( \32130 , \32109 , \32129 );
and \g446999/U$2 ( \32131 , \16774 , RIde7b4b8_191);
and \g446999/U$3 ( \32132 , RIdedb7a0_961, \16776 );
nor \g446999/U$1 ( \32133 , \32131 , \32132 );
and \g446998/U$2 ( \32134 , \16779 , RIdf1c840_1701);
and \g446998/U$3 ( \32135 , RIdf2bfc0_1877, \16781 );
nor \g446998/U$1 ( \32136 , \32134 , \32135 );
and \g446997/U$2 ( \32137 , \16784 , RIdf37960_2009);
and \g446997/U$3 ( \32138 , RIe142f68_2139, \16786 );
nor \g446997/U$1 ( \32139 , \32137 , \32138 );
nand \g444635/U$1 ( \32140 , \32130 , \32133 , \32136 , \32139 );
and \g452788/U$2 ( \32141 , \16361 , RIe167700_2554);
and \g452788/U$3 ( \32142 , RIfc95a98_6725, \16427 );
nor \g452788/U$1 ( \32143 , \32141 , \32142 );
and \g446212/U$2 ( \32144 , RIde80d50_218, \16448 );
and \g446212/U$3 ( \32145 , RIfced068_7719, \16371 );
and \g449163/U$2 ( \32146 , RIfcc1418_7221, \16321 );
and \g449163/U$3 ( \32147 , \16326 , RIfced4a0_7722);
and \g449163/U$4 ( \32148 , RIe16b0a8_2595, \16337 );
nor \g449163/U$1 ( \32149 , \32146 , \32147 , \32148 );
and \g455037/U$2 ( \32150 , \16317 , RIde8c858_275);
and \g455037/U$3 ( \32151 , RIde90368_293, \16325 );
nor \g455037/U$1 ( \32152 , \32150 , \32151 );
not \g450173/U$3 ( \32153 , \32152 );
not \g450173/U$4 ( \32154 , \16330 );
and \g450173/U$2 ( \32155 , \32153 , \32154 );
and \g450173/U$5 ( \32156 , \16341 , RIfcedfe0_7730);
nor \g450173/U$1 ( \32157 , \32155 , \32156 );
and \g452806/U$2 ( \32158 , \16377 , RIfcec0f0_7708);
and \g452806/U$3 ( \32159 , RIfc95930_6724, \16313 );
nor \g452806/U$1 ( \32160 , \32158 , \32159 );
and \g452809/U$2 ( \32161 , \16334 , RIde84ef0_238);
and \g452809/U$3 ( \32162 , RIde893d8_259, \16380 );
nor \g452809/U$1 ( \32163 , \32161 , \32162 );
nand \g447379/U$1 ( \32164 , \32149 , \32157 , \32160 , \32163 );
nor \g446212/U$1 ( \32165 , \32144 , \32145 , \32164 );
and \g452785/U$2 ( \32166 , \16364 , RIe169758_2577);
and \g452785/U$3 ( \32167 , RIfced1d0_7720, \16368 );
nor \g452785/U$1 ( \32168 , \32166 , \32167 );
nand \g445627/U$1 ( \32169 , \32143 , \32165 , \32168 );
and \g444785/U$2 ( \32170 , \32169 , \17998 );
and \g449149/U$2 ( \32171 , RIe151068_2299, \16427 );
and \g449149/U$3 ( \32172 , \16448 , RIfe82818_7829);
and \g449149/U$4 ( \32173 , RIe15c468_2427, \16485 );
nor \g449149/U$1 ( \32174 , \32171 , \32172 , \32173 );
and \g455002/U$2 ( \32175 , \16317 , RIe14b668_2235);
and \g455002/U$3 ( \32176 , RIfc5f9c0_6110, \16325 );
nor \g455002/U$1 ( \32177 , \32175 , \32176 );
not \g455001/U$1 ( \32178 , \32177 );
and \g450157/U$2 ( \32179 , \32178 , \16336 );
and \g450157/U$3 ( \32180 , RIfc426e0_5778, \16356 );
nor \g450157/U$1 ( \32181 , \32179 , \32180 );
and \g452756/U$2 ( \32182 , \16361 , RIe145c68_2171);
and \g452756/U$3 ( \32183 , RIe148968_2203, \16364 );
nor \g452756/U$1 ( \32184 , \32182 , \32183 );
and \g452751/U$2 ( \32185 , \16368 , RIe14e368_2267);
and \g452751/U$3 ( \32186 , RIee34c60_5059, \16371 );
nor \g452751/U$1 ( \32187 , \32185 , \32186 );
nand \g448088/U$1 ( \32188 , \32174 , \32181 , \32184 , \32187 );
and \g444785/U$3 ( \32189 , \16390 , \32188 );
nor \g444785/U$1 ( \32190 , \32170 , \32189 );
and \g446972/U$2 ( \32191 , \18020 , RIe161e68_2491);
and \g446972/U$3 ( \32192 , RIe164b68_2523, \18022 );
nor \g446972/U$1 ( \32193 , \32191 , \32192 );
and \g446973/U$2 ( \32194 , \18025 , RIe15f168_2459);
and \g446973/U$3 ( \32195 , RIee36e20_5083, \18027 );
nor \g446973/U$1 ( \32196 , \32194 , \32195 );
and \g446976/U$2 ( \32197 , \18030 , RIe153d68_2331);
and \g446976/U$3 ( \32198 , RIe156a68_2363, \18032 );
nor \g446976/U$1 ( \32199 , \32197 , \32198 );
nand \g444509/U$1 ( \32200 , \32190 , \32193 , \32196 , \32199 );
and \g446177/U$2 ( \32201 , RIdeb1068_478, \16427 );
and \g446177/U$3 ( \32202 , RIdeae368_446, \16368 );
and \g449115/U$2 ( \32203 , RIdebc468_606, \16485 );
and \g449115/U$3 ( \32204 , \16354 , RIfce6df8_7649);
and \g449115/U$4 ( \32205 , RIdea9070_414, \16398 );
nor \g449115/U$1 ( \32206 , \32203 , \32204 , \32205 );
and \g454949/U$2 ( \32207 , \16317 , RIdec1e68_670);
and \g454949/U$3 ( \32208 , RIdec4b68_702, \16325 );
nor \g454949/U$1 ( \32209 , \32207 , \32208 );
not \g450127/U$3 ( \32210 , \32209 );
not \g450127/U$4 ( \32211 , \16311 );
and \g450127/U$2 ( \32212 , \32210 , \32211 );
and \g450127/U$5 ( \32213 , \16341 , RIfc5e340_6094);
nor \g450127/U$1 ( \32214 , \32212 , \32213 );
and \g452629/U$2 ( \32215 , \16377 , RIdebf168_638);
and \g452629/U$3 ( \32216 , RIfc5df08_6091, \16313 );
nor \g452629/U$1 ( \32217 , \32215 , \32216 );
and \g452635/U$2 ( \32218 , \16334 , RIdeb6a68_542);
and \g452635/U$3 ( \32219 , RIdeb9768_574, \16380 );
nor \g452635/U$1 ( \32220 , \32218 , \32219 );
nand \g447363/U$1 ( \32221 , \32206 , \32214 , \32217 , \32220 );
nor \g446177/U$1 ( \32222 , \32201 , \32202 , \32221 );
and \g452620/U$2 ( \32223 , \16361 , RIde9be70_350);
and \g452620/U$3 ( \32224 , RIfc75ef0_6364, \16448 );
nor \g452620/U$1 ( \32225 , \32223 , \32224 );
and \g452611/U$2 ( \32226 , \16364 , RIdea2770_382);
and \g452611/U$3 ( \32227 , RIfcc12b0_7220, \16371 );
nor \g452611/U$1 ( \32228 , \32226 , \32227 );
and \g445274/U$2 ( \32229 , \32222 , \32225 , \32228 );
nor \g445274/U$1 ( \32230 , \32229 , \16618 );
and \g446187/U$2 ( \32231 , RIfccfef0_7388, \16328 );
and \g446187/U$3 ( \32232 , RIfcafda8_7023, \16377 );
and \g449128/U$2 ( \32233 , RIfebf100_8294, \16398 );
and \g449128/U$3 ( \32234 , \16339 , RIdf34f30_1979);
and \g449128/U$4 ( \32235 , RIdf3e710_2087, \16485 );
nor \g449128/U$1 ( \32236 , \32233 , \32234 , \32235 );
and \g455346/U$2 ( \32237 , \16317 , RIee2f3c8_4996);
and \g455346/U$3 ( \32238 , RIfc5fc90_6112, \16325 );
nor \g455346/U$1 ( \32239 , \32237 , \32238 );
not \g450140/U$3 ( \32240 , \32239 );
not \g450140/U$4 ( \32241 , \16351 );
and \g450140/U$2 ( \32242 , \32240 , \32241 );
and \g450140/U$5 ( \32243 , \16356 , RIe140970_2112);
nor \g450140/U$1 ( \32244 , \32242 , \32243 );
and \g452688/U$2 ( \32245 , \16361 , RIdf2ecc0_1909);
and \g452688/U$3 ( \32246 , RIdf30a48_1930, \16364 );
nor \g452688/U$1 ( \32247 , \32245 , \32246 );
and \g452680/U$2 ( \32248 , \16368 , RIee2d208_4972);
and \g452680/U$3 ( \32249 , RIfc742d0_6344, \16371 );
nor \g452680/U$1 ( \32250 , \32248 , \32249 );
nand \g447787/U$1 ( \32251 , \32236 , \32244 , \32247 , \32250 );
nor \g446187/U$1 ( \32252 , \32231 , \32232 , \32251 );
and \g452664/U$2 ( \32253 , \16334 , RIdf3a228_2038);
and \g452664/U$3 ( \32254 , RIfc600c8_6115, \16313 );
nor \g452664/U$1 ( \32255 , \32253 , \32254 );
and \g452661/U$2 ( \32256 , \16380 , RIdf3c6b8_2064);
and \g452661/U$3 ( \32257 , RIfca57b8_6905, \16319 );
nor \g452661/U$1 ( \32258 , \32256 , \32257 );
and \g445286/U$2 ( \32259 , \32252 , \32255 , \32258 );
nor \g445286/U$1 ( \32260 , \32259 , \16393 );
or \g444402/U$1 ( \32261 , \32140 , \32200 , \32230 , \32260 );
and \g446158/U$2 ( \32262 , RIfcb08e8_7031, \16326 );
and \g446158/U$3 ( \32263 , RIfcdef68_7559, \16377 );
and \g449088/U$2 ( \32264 , RIfcee850_7736, \16427 );
and \g449088/U$3 ( \32265 , \16432 , RIfc5ed18_6101);
and \g449088/U$4 ( \32266 , RIdf27c40_1829, \16485 );
nor \g449088/U$1 ( \32267 , \32264 , \32265 , \32266 );
and \g454165/U$2 ( \32268 , \16317 , RIfeaa520_8254);
and \g454165/U$3 ( \32269 , RIdf212c8_1754, \16325 );
nor \g454165/U$1 ( \32270 , \32268 , \32269 );
not \g454164/U$1 ( \32271 , \32270 );
and \g450103/U$2 ( \32272 , \32271 , \16336 );
and \g450103/U$3 ( \32273 , RIdf29e00_1853, \16354 );
nor \g450103/U$1 ( \32274 , \32272 , \32273 );
and \g452556/U$2 ( \32275 , \16361 , RIdf18e98_1660);
and \g452556/U$3 ( \32276 , RIdf1ad88_1682, \16364 );
nor \g452556/U$1 ( \32277 , \32275 , \32276 );
and \g452549/U$2 ( \32278 , \16368 , RIfc5efe8_6103);
and \g452549/U$3 ( \32279 , RIdf227e0_1769, \16371 );
nor \g452549/U$1 ( \32280 , \32278 , \32279 );
nand \g448076/U$1 ( \32281 , \32267 , \32274 , \32277 , \32280 );
nor \g446158/U$1 ( \32282 , \32262 , \32263 , \32281 );
and \g452537/U$2 ( \32283 , \16334 , RIdf24298_1788);
and \g452537/U$3 ( \32284 , RIfc95ed0_6728, \16313 );
nor \g452537/U$1 ( \32285 , \32283 , \32284 );
and \g452530/U$2 ( \32286 , \16380 , RIdf25eb8_1808);
and \g452530/U$3 ( \32287 , RIfcee418_7733, \16321 );
nor \g452530/U$1 ( \32288 , \32286 , \32287 );
and \g445261/U$2 ( \32289 , \32282 , \32285 , \32288 );
nor \g445261/U$1 ( \32290 , \32289 , \16480 );
and \g446167/U$2 ( \32291 , RIdf13a38_1600, \16321 );
and \g446167/U$3 ( \32292 , RIdf10d38_1568, \16313 );
and \g449100/U$2 ( \32293 , RIdefa538_1312, \16427 );
and \g449100/U$3 ( \32294 , \16448 , RIdefd238_1344);
and \g449100/U$4 ( \32295 , RIdf08638_1472, \16485 );
nor \g449100/U$1 ( \32296 , \32293 , \32294 , \32295 );
and \g454925/U$2 ( \32297 , \16317 , RIdeef138_1184);
and \g454925/U$3 ( \32298 , RIdef1e38_1216, \16325 );
nor \g454925/U$1 ( \32299 , \32297 , \32298 );
not \g454924/U$1 ( \32300 , \32299 );
and \g450115/U$2 ( \32301 , \32300 , \16336 );
and \g450115/U$3 ( \32302 , RIdf0b338_1504, \16356 );
nor \g450115/U$1 ( \32303 , \32301 , \32302 );
and \g452588/U$2 ( \32304 , \16361 , RIdee9738_1120);
and \g452588/U$3 ( \32305 , RIdeec438_1152, \16364 );
nor \g452588/U$1 ( \32306 , \32304 , \32305 );
and \g452583/U$2 ( \32307 , \16368 , RIdef4b38_1248);
and \g452583/U$3 ( \32308 , RIdef7838_1280, \16371 );
nor \g452583/U$1 ( \32309 , \32307 , \32308 );
nand \g448080/U$1 ( \32310 , \32296 , \32303 , \32306 , \32309 );
nor \g446167/U$1 ( \32311 , \32291 , \32292 , \32310 );
and \g452576/U$2 ( \32312 , \16377 , RIdf0e038_1536);
and \g452576/U$3 ( \32313 , RIdf05938_1440, \16380 );
nor \g452576/U$1 ( \32314 , \32312 , \32313 );
and \g452570/U$2 ( \32315 , \16334 , RIdf02c38_1408);
and \g452570/U$3 ( \32316 , RIdf16738_1632, \16326 );
nor \g452570/U$1 ( \32317 , \32315 , \32316 );
and \g445269/U$2 ( \32318 , \32311 , \32314 , \32317 );
nor \g445269/U$1 ( \32319 , \32318 , \16555 );
or \g444259/U$1 ( \32320 , \32261 , \32290 , \32319 );
_DC \g556a/U$1 ( \32321 , \32320 , \16652 );
and \g453215/U$2 ( \32322 , \8404 , RIfe82548_7827);
and \g453215/U$3 ( \32323 , RIfcbff00_7206, \8409 );
nor \g453215/U$1 ( \32324 , \32322 , \32323 );
and \g446300/U$2 ( \32325 , RIfcb1e00_7046, \8373 );
and \g446300/U$3 ( \32326 , RIee3d090_5153, \8378 );
and \g449271/U$2 ( \32327 , RIfc5c450_6072, \8317 );
and \g449271/U$3 ( \32328 , \8326 , RIfebecc8_8291);
and \g449271/U$4 ( \32329 , RIfce7398_7653, \8383 );
nor \g449271/U$1 ( \32330 , \32327 , \32328 , \32329 );
and \g453230/U$2 ( \32331 , \8335 , RIfce9288_7675);
and \g453230/U$3 ( \32332 , RIf16fef8_5733, \8340 );
nor \g453230/U$1 ( \32333 , \32331 , \32332 );
and \g455276/U$2 ( \32334 , \8313 , RIee399b8_5114);
and \g455276/U$3 ( \32335 , RIfce35b8_7609, \8323 );
nor \g455276/U$1 ( \32336 , \32334 , \32335 );
not \g450287/U$3 ( \32337 , \32336 );
not \g450287/U$4 ( \32338 , \8347 );
and \g450287/U$2 ( \32339 , \32337 , \32338 );
and \g450287/U$5 ( \32340 , \8351 , RIf141f80_5210);
nor \g450287/U$1 ( \32341 , \32339 , \32340 );
and \g453228/U$2 ( \32342 , \8356 , RIfea8a68_8235);
and \g453228/U$3 ( \32343 , RIfc5c180_6070, \8359 );
nor \g453228/U$1 ( \32344 , \32342 , \32343 );
nand \g447867/U$1 ( \32345 , \32330 , \32333 , \32341 , \32344 );
nor \g446300/U$1 ( \32346 , \32325 , \32326 , \32345 );
and \g453212/U$2 ( \32347 , \8414 , RIfcaaee8_6967);
and \g453212/U$3 ( \32348 , RIfca42a0_6890, \8417 );
nor \g453212/U$1 ( \32349 , \32347 , \32348 );
nand \g445650/U$1 ( \32350 , \32324 , \32346 , \32349 );
and \g444697/U$2 ( \32351 , \32350 , \9700 );
and \g449260/U$2 ( \32352 , RIe191a00_3034, \8414 );
and \g449260/U$3 ( \32353 , \8409 , RIe194700_3066);
and \g449260/U$4 ( \32354 , RIe186600_2906, \8488 );
nor \g449260/U$1 ( \32355 , \32352 , \32353 , \32354 );
and \g455290/U$2 ( \32356 , \8313 , RIfce96c0_7678);
and \g455290/U$3 ( \32357 , RIe19a100_3130, \8323 );
nor \g455290/U$1 ( \32358 , \32356 , \32357 );
not \g450276/U$3 ( \32359 , \32358 );
not \g450276/U$4 ( \32360 , \8328 );
and \g450276/U$2 ( \32361 , \32359 , \32360 );
and \g450276/U$5 ( \32362 , \8359 , RIe189300_2938);
nor \g450276/U$1 ( \32363 , \32361 , \32362 );
and \g453186/U$2 ( \32364 , \8404 , RIe197400_3098);
and \g453186/U$3 ( \32365 , RIe19ce00_3162, \8351 );
nor \g453186/U$1 ( \32366 , \32364 , \32365 );
and \g453194/U$2 ( \32367 , \8378 , RIe18ed00_3002);
and \g453194/U$3 ( \32368 , RIf144410_5236, \8417 );
nor \g453194/U$1 ( \32369 , \32367 , \32368 );
nand \g447861/U$1 ( \32370 , \32355 , \32363 , \32366 , \32369 );
and \g444697/U$3 ( \32371 , \9702 , \32370 );
nor \g444697/U$1 ( \32372 , \32351 , \32371 );
and \g447063/U$2 ( \32373 , \9729 , RIe17b200_2778);
and \g447063/U$3 ( \32374 , RIe17df00_2810, \9731 );
nor \g447063/U$1 ( \32375 , \32373 , \32374 );
and \g447058/U$2 ( \32376 , \9230 , RIe183900_2874);
and \g447058/U$3 ( \32377 , RIfebee30_8292, \9232 );
nor \g447058/U$1 ( \32378 , \32376 , \32377 );
and \g447059/U$2 ( \32379 , \9734 , RIe180c00_2842);
and \g447059/U$3 ( \32380 , RIfcdbcc8_7523, \9736 );
nor \g447059/U$1 ( \32381 , \32379 , \32380 );
nand \g444523/U$1 ( \32382 , \32372 , \32375 , \32378 , \32381 );
and \g453298/U$2 ( \32383 , \8404 , RIfebef98_8293);
and \g453298/U$3 ( \32384 , RIfcd7ab0_7476, \8407 );
nor \g453298/U$1 ( \32385 , \32383 , \32384 );
and \g446316/U$2 ( \32386 , RIfc5d0f8_6081, \8371 );
and \g446316/U$3 ( \32387 , RIfeaa0e8_8251, \8378 );
and \g449294/U$2 ( \32388 , RIfcec258_7709, \8319 );
and \g449294/U$3 ( \32389 , \8326 , RIfc772a0_6378);
and \g449294/U$4 ( \32390 , RIf157808_5455, \8383 );
nor \g449294/U$1 ( \32391 , \32388 , \32389 , \32390 );
and \g453313/U$2 ( \32392 , \8335 , RIe1ed8f0_4080);
and \g453313/U$3 ( \32393 , RIf14f540_5362, \8340 );
nor \g453313/U$1 ( \32394 , \32392 , \32393 );
and \g454344/U$2 ( \32395 , \8313 , RIf1504b8_5373);
and \g454344/U$3 ( \32396 , RIfce3450_7608, \8323 );
nor \g454344/U$1 ( \32397 , \32395 , \32396 );
not \g450310/U$3 ( \32398 , \32397 );
not \g450310/U$4 ( \32399 , \8347 );
and \g450310/U$2 ( \32400 , \32398 , \32399 );
and \g450310/U$5 ( \32401 , \8351 , RIf158bb8_5469);
nor \g450310/U$1 ( \32402 , \32400 , \32401 );
and \g453309/U$2 ( \32403 , \8356 , RIe1f2be8_4139);
and \g453309/U$3 ( \32404 , RIfccc548_7347, \8359 );
nor \g453309/U$1 ( \32405 , \32403 , \32404 );
nand \g447881/U$1 ( \32406 , \32391 , \32394 , \32402 , \32405 );
nor \g446316/U$1 ( \32407 , \32386 , \32387 , \32406 );
and \g453293/U$2 ( \32408 , \8414 , RIfcb1428_7039);
and \g453293/U$3 ( \32409 , RIfcc8a38_7305, \8417 );
nor \g453293/U$1 ( \32410 , \32408 , \32409 );
nand \g445658/U$1 ( \32411 , \32385 , \32407 , \32410 );
and \g444729/U$2 ( \32412 , \32411 , \8752 );
and \g449284/U$2 ( \32413 , RIe1e54c0_3986, \8373 );
and \g449284/U$3 ( \32414 , \8383 , RIe1e81c0_4018);
and \g449284/U$4 ( \32415 , RIe1cecc0_3730, \8488 );
nor \g449284/U$1 ( \32416 , \32413 , \32414 , \32415 );
and \g454426/U$2 ( \32417 , \8313 , RIe1da0c0_3858);
and \g454426/U$3 ( \32418 , RIe1dcdc0_3890, \8323 );
nor \g454426/U$1 ( \32419 , \32417 , \32418 );
not \g450301/U$3 ( \32420 , \32419 );
not \g450301/U$4 ( \32421 , \8376 );
and \g450301/U$2 ( \32422 , \32420 , \32421 );
and \g450301/U$5 ( \32423 , \8359 , RIe1d19c0_3762);
nor \g450301/U$1 ( \32424 , \32422 , \32423 );
and \g453268/U$2 ( \32425 , \8404 , RIe1e27c0_3954);
and \g453268/U$3 ( \32426 , RIe1eaec0_4050, \8351 );
nor \g453268/U$1 ( \32427 , \32425 , \32426 );
and \g453274/U$2 ( \32428 , \8378 , RIe1d73c0_3826);
and \g453274/U$3 ( \32429 , RIe1dfac0_3922, \8417 );
nor \g453274/U$1 ( \32430 , \32428 , \32429 );
nand \g447874/U$1 ( \32431 , \32416 , \32424 , \32427 , \32430 );
and \g444729/U$3 ( \32432 , \8478 , \32431 );
nor \g444729/U$1 ( \32433 , \32412 , \32432 );
and \g447079/U$2 ( \32434 , \8775 , RIe1c92c0_3666);
and \g447079/U$3 ( \32435 , RIe1cbfc0_3698, \8777 );
nor \g447079/U$1 ( \32436 , \32434 , \32435 );
and \g447080/U$2 ( \32437 , \8780 , RIe1c38c0_3602);
and \g447080/U$3 ( \32438 , RIe1c65c0_3634, \8782 );
nor \g447080/U$1 ( \32439 , \32437 , \32438 );
and \g447083/U$2 ( \32440 , \8785 , RIe1bdec0_3538);
and \g447083/U$3 ( \32441 , RIe1c0bc0_3570, \8787 );
nor \g447083/U$1 ( \32442 , \32440 , \32441 );
nand \g444651/U$1 ( \32443 , \32433 , \32436 , \32439 , \32442 );
and \g446266/U$2 ( \32444 , RIe1a2800_3226, \8371 );
and \g446266/U$3 ( \32445 , RIe21aa58_4593, \8378 );
and \g449232/U$2 ( \32446 , RIe1ae038_3357, \8319 );
and \g449232/U$3 ( \32447 , \8326 , RIe1bb1c0_3506);
and \g449232/U$4 ( \32448 , RIe1a5500_3258, \8383 );
nor \g449232/U$1 ( \32449 , \32446 , \32447 , \32448 );
and \g453075/U$2 ( \32450 , \8335 , RIe170670_2656);
and \g453075/U$3 ( \32451 , RIe1d46c0_3794, \8340 );
nor \g453075/U$1 ( \32452 , \32450 , \32451 );
and \g455210/U$2 ( \32453 , \8313 , RIe1f7670_4192);
and \g455210/U$3 ( \32454 , RIe1fe2b8_4269, \8323 );
nor \g455210/U$1 ( \32455 , \32453 , \32454 );
not \g450246/U$3 ( \32456 , \32455 );
not \g450246/U$4 ( \32457 , \8347 );
and \g450246/U$2 ( \32458 , \32456 , \32457 );
and \g450246/U$5 ( \32459 , \8351 , RIe1a8200_3290);
nor \g450246/U$1 ( \32460 , \32458 , \32459 );
and \g453072/U$2 ( \32461 , \8356 , RIe1f01b8_4109);
and \g453072/U$3 ( \32462 , RIe204258_4337, \8359 );
nor \g453072/U$1 ( \32463 , \32461 , \32462 );
nand \g447846/U$1 ( \32464 , \32449 , \32452 , \32460 , \32463 );
nor \g446266/U$1 ( \32465 , \32444 , \32445 , \32464 );
and \g453056/U$2 ( \32466 , \8404 , RIe19fb00_3194);
and \g453056/U$3 ( \32467 , RIe178500_2746, \8409 );
nor \g453056/U$1 ( \32468 , \32466 , \32467 );
and \g453053/U$2 ( \32469 , \8414 , RIe225e58_4721);
and \g453053/U$3 ( \32470 , RIe18c000_2970, \8417 );
nor \g453053/U$1 ( \32471 , \32469 , \32470 );
and \g445339/U$2 ( \32472 , \32465 , \32468 , \32471 );
nor \g445339/U$1 ( \32473 , \32472 , \8651 );
and \g446276/U$2 ( \32474 , RIfe823e0_7826, \8523 );
and \g446276/U$3 ( \32475 , RIfe82278_7825, \8319 );
and \g449247/U$2 ( \32476 , RIe1b4f50_3436, \8414 );
and \g449247/U$3 ( \32477 , \8409 , RIfc94b20_6714);
and \g449247/U$4 ( \32478 , RIfceb010_7696, \8488 );
nor \g449247/U$1 ( \32479 , \32476 , \32477 , \32478 );
and \g454690/U$2 ( \32480 , \8313 , RIe1b8e98_3481);
and \g454690/U$3 ( \32481 , RIf14b328_5315, \8323 );
nor \g454690/U$1 ( \32482 , \32480 , \32481 );
not \g450261/U$3 ( \32483 , \32482 );
not \g450261/U$4 ( \32484 , \8328 );
and \g450261/U$2 ( \32485 , \32483 , \32484 );
and \g450261/U$5 ( \32486 , \8359 , RIfcec3c0_7710);
nor \g450261/U$1 ( \32487 , \32485 , \32486 );
and \g453123/U$2 ( \32488 , \8404 , RIe1b6e40_3458);
and \g453123/U$3 ( \32489 , RIf14c570_5328, \8351 );
nor \g453123/U$1 ( \32490 , \32488 , \32489 );
and \g453135/U$2 ( \32491 , \8378 , RIe1b3ba0_3422);
and \g453135/U$3 ( \32492 , RIfc76760_6370, \8417 );
nor \g453135/U$1 ( \32493 , \32491 , \32492 );
nand \g447851/U$1 ( \32494 , \32479 , \32487 , \32490 , \32493 );
nor \g446276/U$1 ( \32495 , \32474 , \32475 , \32494 );
and \g453107/U$2 ( \32496 , \8335 , RIe1aa7f8_3317);
and \g453107/U$3 ( \32497 , RIfcdd8e8_7543, \8340 );
nor \g453107/U$1 ( \32498 , \32496 , \32497 );
and \g453102/U$2 ( \32499 , \8326 , RIfcc0ba8_7215);
and \g453102/U$3 ( \32500 , RIfe82110_7824, \8356 );
nor \g453102/U$1 ( \32501 , \32499 , \32500 );
and \g445341/U$2 ( \32502 , \32495 , \32498 , \32501 );
nor \g445341/U$1 ( \32503 , \32502 , \8481 );
or \g444324/U$1 ( \32504 , \32382 , \32443 , \32473 , \32503 );
and \g446247/U$2 ( \32505 , RIfce1998_7589, \8531 );
and \g446247/U$3 ( \32506 , RIe209c58_4401, \8319 );
and \g449206/U$2 ( \32507 , RIfce77d0_7656, \8373 );
and \g449206/U$3 ( \32508 , \8383 , RIe223158_4689);
and \g449206/U$4 ( \32509 , RIe212358_4497, \8488 );
nor \g449206/U$1 ( \32510 , \32507 , \32508 , \32509 );
and \g455142/U$2 ( \32511 , \8313 , RIe217d58_4561);
and \g455142/U$3 ( \32512 , RIe21d758_4625, \8323 );
nor \g455142/U$1 ( \32513 , \32511 , \32512 );
not \g450219/U$3 ( \32514 , \32513 );
not \g450219/U$4 ( \32515 , \8376 );
and \g450219/U$2 ( \32516 , \32514 , \32515 );
and \g450219/U$5 ( \32517 , \8359 , RIfce8a18_7669);
nor \g450219/U$1 ( \32518 , \32516 , \32517 );
and \g452974/U$2 ( \32519 , \8404 , RIe220458_4657);
and \g452974/U$3 ( \32520 , RIfc40778_5759, \8351 );
nor \g452974/U$1 ( \32521 , \32519 , \32520 );
and \g452977/U$2 ( \32522 , \8378 , RIe215058_4529);
and \g452977/U$3 ( \32523 , RIfce24d8_7597, \8417 );
nor \g452977/U$1 ( \32524 , \32522 , \32523 );
nand \g447829/U$1 ( \32525 , \32510 , \32518 , \32521 , \32524 );
nor \g446247/U$1 ( \32526 , \32505 , \32506 , \32525 );
and \g452959/U$2 ( \32527 , \8335 , RIe206f58_4369);
and \g452959/U$3 ( \32528 , RIfc77840_6382, \8340 );
nor \g452959/U$1 ( \32529 , \32527 , \32528 );
and \g452956/U$2 ( \32530 , \8324 , RIe20c958_4433);
and \g452956/U$3 ( \32531 , RIe20f658_4465, \8356 );
nor \g452956/U$1 ( \32532 , \32530 , \32531 );
and \g445324/U$2 ( \32533 , \32526 , \32529 , \32532 );
nor \g445324/U$1 ( \32534 , \32533 , \8368 );
and \g446257/U$2 ( \32535 , RIfe81fa8_7823, \8373 );
and \g446257/U$3 ( \32536 , RIf1619c0_5570, \8378 );
and \g449220/U$2 ( \32537 , RIfcd0fd0_7400, \8317 );
and \g449220/U$3 ( \32538 , \8326 , RIf15b1b0_5496);
and \g449220/U$4 ( \32539 , RIf165bd8_5617, \8383 );
nor \g449220/U$1 ( \32540 , \32537 , \32538 , \32539 );
and \g453019/U$2 ( \32541 , \8335 , RIfccc6b0_7348);
and \g453019/U$3 ( \32542 , RIf15c830_5512, \8340 );
nor \g453019/U$1 ( \32543 , \32541 , \32542 );
and \g454329/U$2 ( \32544 , \8313 , RIe1fc800_4250);
and \g454329/U$3 ( \32545 , RIfc77570_6380, \8323 );
nor \g454329/U$1 ( \32546 , \32544 , \32545 );
not \g450234/U$3 ( \32547 , \32546 );
not \g450234/U$4 ( \32548 , \8347 );
and \g450234/U$2 ( \32549 , \32547 , \32548 );
and \g450234/U$5 ( \32550 , \8351 , RIf166cb8_5629);
nor \g450234/U$1 ( \32551 , \32549 , \32550 );
and \g453016/U$2 ( \32552 , \8356 , RIe1fb720_4238);
and \g453016/U$3 ( \32553 , RIfccf248_7379, \8359 );
nor \g453016/U$1 ( \32554 , \32552 , \32553 );
nand \g447835/U$1 ( \32555 , \32540 , \32543 , \32551 , \32554 );
nor \g446257/U$1 ( \32556 , \32535 , \32536 , \32555 );
and \g453007/U$2 ( \32557 , \8404 , RIfe81e40_7822);
and \g453007/U$3 ( \32558 , RIfceb178_7697, \8407 );
nor \g453007/U$1 ( \32559 , \32557 , \32558 );
and \g453001/U$2 ( \32560 , \8414 , RIf1631a8_5587);
and \g453001/U$3 ( \32561 , RIfc5c888_6075, \8417 );
nor \g453001/U$1 ( \32562 , \32560 , \32561 );
and \g445325/U$2 ( \32563 , \32556 , \32559 , \32562 );
nor \g445325/U$1 ( \32564 , \32563 , \8422 );
or \g444245/U$1 ( \32565 , \32504 , \32534 , \32564 );
_DC \g55ee/U$1 ( \32566 , \32565 , \8654 );
and \g453594/U$2 ( \32567 , \16364 , RIfc43220_5786);
and \g453594/U$3 ( \32568 , RIfcc2390_7232, \16371 );
nor \g453594/U$1 ( \32569 , \32567 , \32568 );
and \g446382/U$2 ( \32570 , RIfe831f0_7836, \16427 );
and \g446382/U$3 ( \32571 , RIee195a0_4747, \16368 );
and \g449376/U$2 ( \32572 , RIde8cba0_276, \16485 );
and \g449376/U$3 ( \32573 , \16356 , RIde906b0_294);
and \g449376/U$4 ( \32574 , RIfea9e18_8249, \16398 );
nor \g449376/U$1 ( \32575 , \32572 , \32573 , \32574 );
and \g455378/U$2 ( \32576 , \16317 , RIfc7af18_6421);
and \g455378/U$3 ( \32577 , RIfc90ea8_6671, \16325 );
nor \g455378/U$1 ( \32578 , \32576 , \32577 );
not \g450394/U$3 ( \32579 , \32578 );
not \g450394/U$4 ( \32580 , \16311 );
and \g450394/U$2 ( \32581 , \32579 , \32580 );
and \g450394/U$5 ( \32582 , \16341 , RIfcbe718_7189);
nor \g450394/U$1 ( \32583 , \32581 , \32582 );
and \g453609/U$2 ( \32584 , \16377 , RIee1a950_4761);
and \g453609/U$3 ( \32585 , RIfe83088_7835, \16313 );
nor \g453609/U$1 ( \32586 , \32584 , \32585 );
and \g453612/U$2 ( \32587 , \16334 , RIfe82db8_7833);
and \g453612/U$3 ( \32588 , RIfe82f20_7834, \16380 );
nor \g453612/U$1 ( \32589 , \32587 , \32588 );
nand \g447419/U$1 ( \32590 , \32575 , \32583 , \32586 , \32589 );
nor \g446382/U$1 ( \32591 , \32570 , \32571 , \32590 );
and \g453596/U$2 ( \32592 , \16361 , RIe167868_2555);
and \g453596/U$3 ( \32593 , RIee1a248_4756, \16448 );
nor \g453596/U$1 ( \32594 , \32592 , \32593 );
nand \g445675/U$1 ( \32595 , \32569 , \32591 , \32594 );
and \g444712/U$2 ( \32596 , \32595 , \17998 );
and \g449365/U$2 ( \32597 , RIdea93b8_415, \16337 );
and \g449365/U$3 ( \32598 , \16341 , RIfc437c0_5790);
and \g449365/U$4 ( \32599 , RIdebc5d0_607, \16485 );
nor \g449365/U$1 ( \32600 , \32597 , \32598 , \32599 );
and \g454549/U$2 ( \32601 , \16317 , RIdeb11d0_479);
and \g454549/U$3 ( \32602 , RIfe83358_7837, \16325 );
nor \g454549/U$1 ( \32603 , \32601 , \32602 );
not \g450384/U$3 ( \32604 , \32603 );
not \g450384/U$4 ( \32605 , \16351 );
and \g450384/U$2 ( \32606 , \32604 , \32605 );
and \g450384/U$5 ( \32607 , \16356 , RIfc7b1e8_6423);
nor \g450384/U$1 ( \32608 , \32606 , \32607 );
and \g453570/U$2 ( \32609 , \16361 , RIde9c1b8_351);
and \g453570/U$3 ( \32610 , RIdea2ab8_383, \16364 );
nor \g453570/U$1 ( \32611 , \32609 , \32610 );
and \g453561/U$2 ( \32612 , \16368 , RIdeae4d0_447);
and \g453561/U$3 ( \32613 , RIee1e5c8_4804, \16371 );
nor \g453561/U$1 ( \32614 , \32612 , \32613 );
nand \g447922/U$1 ( \32615 , \32600 , \32608 , \32611 , \32614 );
and \g444712/U$3 ( \32616 , \17938 , \32615 );
nor \g444712/U$1 ( \32617 , \32596 , \32616 );
and \g447126/U$2 ( \32618 , \18960 , RIdeb6bd0_543);
and \g447126/U$3 ( \32619 , RIdeb98d0_575, \18962 );
nor \g447126/U$1 ( \32620 , \32618 , \32619 );
and \g447123/U$2 ( \32621 , \18965 , RIdec1fd0_671);
and \g447123/U$3 ( \32622 , RIdec4cd0_703, \18967 );
nor \g447123/U$1 ( \32623 , \32621 , \32622 );
and \g447131/U$2 ( \32624 , \18776 , RIdebf2d0_639);
and \g447131/U$3 ( \32625 , RIfc7b4b8_6425, \18778 );
nor \g447131/U$1 ( \32626 , \32624 , \32625 );
nand \g444531/U$1 ( \32627 , \32617 , \32620 , \32623 , \32626 );
and \g453672/U$2 ( \32628 , \16364 , RIe148ad0_2204);
and \g453672/U$3 ( \32629 , RIfebfda8_8303, \16371 );
nor \g453672/U$1 ( \32630 , \32628 , \32629 );
and \g446399/U$2 ( \32631 , RIe1511d0_2300, \16427 );
and \g446399/U$3 ( \32632 , RIe14e4d0_2268, \16368 );
and \g449401/U$2 ( \32633 , RIe15c5d0_2428, \16344 );
and \g449401/U$3 ( \32634 , \16356 , RIee35ea8_5072);
and \g449401/U$4 ( \32635 , RIe14b7d0_2236, \16398 );
nor \g449401/U$1 ( \32636 , \32633 , \32634 , \32635 );
and \g455120/U$2 ( \32637 , \16317 , RIe161fd0_2492);
and \g455120/U$3 ( \32638 , RIe164cd0_2524, \16325 );
nor \g455120/U$1 ( \32639 , \32637 , \32638 );
not \g450418/U$3 ( \32640 , \32639 );
not \g450418/U$4 ( \32641 , \16311 );
and \g450418/U$2 ( \32642 , \32640 , \32641 );
and \g450418/U$5 ( \32643 , \16339 , RIfebfc40_8302);
nor \g450418/U$1 ( \32644 , \32642 , \32643 );
and \g453689/U$2 ( \32645 , \16377 , RIe15f2d0_2460);
and \g453689/U$3 ( \32646 , RIee36f88_5084, \16313 );
nor \g453689/U$1 ( \32647 , \32645 , \32646 );
and \g453704/U$2 ( \32648 , \16334 , RIe153ed0_2332);
and \g453704/U$3 ( \32649 , RIe156bd0_2364, \16380 );
nor \g453704/U$1 ( \32650 , \32648 , \32649 );
nand \g447422/U$1 ( \32651 , \32636 , \32644 , \32647 , \32650 );
nor \g446399/U$1 ( \32652 , \32631 , \32632 , \32651 );
and \g453682/U$2 ( \32653 , \16361 , RIe145dd0_2172);
and \g453682/U$3 ( \32654 , RIfe83628_7839, \16448 );
nor \g453682/U$1 ( \32655 , \32653 , \32654 );
nand \g445678/U$1 ( \32656 , \32630 , \32652 , \32655 );
and \g444863/U$2 ( \32657 , \32656 , \16390 );
and \g449390/U$2 ( \32658 , RIee32ed8_5038, \16321 );
and \g449390/U$3 ( \32659 , \16328 , RIee34120_5051);
and \g449390/U$4 ( \32660 , RIfeab600_8266, \16398 );
nor \g449390/U$1 ( \32661 , \32658 , \32659 , \32660 );
and \g455286/U$2 ( \32662 , \16317 , RIdf3e878_2088);
and \g455286/U$3 ( \32663 , RIe140ad8_2113, \16325 );
nor \g455286/U$1 ( \32664 , \32662 , \32663 );
not \g450405/U$3 ( \32665 , \32664 );
not \g450405/U$4 ( \32666 , \16330 );
and \g450405/U$2 ( \32667 , \32665 , \32666 );
and \g450405/U$5 ( \32668 , \16339 , RIdf35098_1980);
nor \g450405/U$1 ( \32669 , \32667 , \32668 );
and \g453654/U$2 ( \32670 , \16377 , RIfcc1f58_7229);
and \g453654/U$3 ( \32671 , RIee31df8_5026, \16313 );
nor \g453654/U$1 ( \32672 , \32670 , \32671 );
and \g453656/U$2 ( \32673 , \16334 , RIdf3a390_2039);
and \g453656/U$3 ( \32674 , RIfe834c0_7838, \16380 );
nor \g453656/U$1 ( \32675 , \32673 , \32674 );
nand \g447421/U$1 ( \32676 , \32661 , \32669 , \32672 , \32675 );
and \g444863/U$3 ( \32677 , \16394 , \32676 );
nor \g444863/U$1 ( \32678 , \32657 , \32677 );
and \g447146/U$2 ( \32679 , \16419 , RIfeab768_8267);
and \g447146/U$3 ( \32680 , RIdf30bb0_1931, \16422 );
nor \g447146/U$1 ( \32681 , \32679 , \32680 );
and \g447144/U$2 ( \32682 , \16429 , RIfc91e20_6682);
and \g447144/U$3 ( \32683 , RIfc5a6c8_6051, \16434 );
nor \g447144/U$1 ( \32684 , \32682 , \32683 );
and \g447145/U$2 ( \32685 , \16438 , RIfc96a10_6736);
and \g447145/U$3 ( \32686 , RIee2e888_4988, \16441 );
nor \g447145/U$1 ( \32687 , \32685 , \32686 );
nand \g444659/U$1 ( \32688 , \32678 , \32681 , \32684 , \32687 );
and \g446349/U$2 ( \32689 , RIdefd3a0_1345, \16448 );
and \g446349/U$3 ( \32690 , RIdef79a0_1281, \16371 );
and \g449333/U$2 ( \32691 , RIdf13ba0_1601, \16321 );
and \g449333/U$3 ( \32692 , \16326 , RIdf168a0_1633);
and \g449333/U$4 ( \32693 , RIdeef2a0_1185, \16398 );
nor \g449333/U$1 ( \32694 , \32691 , \32692 , \32693 );
and \g455199/U$2 ( \32695 , \16317 , RIdf087a0_1473);
and \g455199/U$3 ( \32696 , RIdf0b4a0_1505, \16325 );
nor \g455199/U$1 ( \32697 , \32695 , \32696 );
not \g450352/U$3 ( \32698 , \32697 );
not \g450352/U$4 ( \32699 , \16330 );
and \g450352/U$2 ( \32700 , \32698 , \32699 );
and \g450352/U$5 ( \32701 , \16341 , RIdef1fa0_1217);
nor \g450352/U$1 ( \32702 , \32700 , \32701 );
and \g453455/U$2 ( \32703 , \16377 , RIdf0e1a0_1537);
and \g453455/U$3 ( \32704 , RIdf10ea0_1569, \16313 );
nor \g453455/U$1 ( \32705 , \32703 , \32704 );
and \g453463/U$2 ( \32706 , \16334 , RIdf02da0_1409);
and \g453463/U$3 ( \32707 , RIdf05aa0_1441, \16380 );
nor \g453463/U$1 ( \32708 , \32706 , \32707 );
nand \g447416/U$1 ( \32709 , \32694 , \32702 , \32705 , \32708 );
nor \g446349/U$1 ( \32710 , \32689 , \32690 , \32709 );
and \g453437/U$2 ( \32711 , \16364 , RIdeec5a0_1153);
and \g453437/U$3 ( \32712 , RIdef4ca0_1249, \16368 );
nor \g453437/U$1 ( \32713 , \32711 , \32712 );
and \g453443/U$2 ( \32714 , \16361 , RIdee98a0_1121);
and \g453443/U$3 ( \32715 , RIdefa6a0_1313, \16427 );
nor \g453443/U$1 ( \32716 , \32714 , \32715 );
and \g445396/U$2 ( \32717 , \32710 , \32713 , \32716 );
nor \g445396/U$1 ( \32718 , \32717 , \16555 );
and \g446359/U$2 ( \32719 , RIdecd3d0_799, \16321 );
and \g446359/U$3 ( \32720 , RIdeca6d0_767, \16313 );
and \g449348/U$2 ( \32721 , RIdee6ba0_1089, \16398 );
and \g449348/U$3 ( \32722 , \16341 , RIdf000a0_1377);
and \g449348/U$4 ( \32723 , RIde958b8_319, \16485 );
nor \g449348/U$1 ( \32724 , \32721 , \32722 , \32723 );
and \g455191/U$2 ( \32725 , \16317 , RIdf37ac8_2010);
and \g455191/U$3 ( \32726 , RIe1430d0_2140, \16325 );
nor \g455191/U$1 ( \32727 , \32725 , \32726 );
not \g450366/U$3 ( \32728 , \32727 );
not \g450366/U$4 ( \32729 , \16351 );
and \g450366/U$2 ( \32730 , \32728 , \32729 );
and \g450366/U$5 ( \32731 , \16356 , RIdeb3ed0_511);
nor \g450366/U$1 ( \32732 , \32730 , \32731 );
and \g453507/U$2 ( \32733 , \16361 , RIde7b800_192);
and \g453507/U$3 ( \32734 , RIdedb908_962, \16364 );
nor \g453507/U$1 ( \32735 , \32733 , \32734 );
and \g453502/U$2 ( \32736 , \16368 , RIdf1c9a8_1702);
and \g453502/U$3 ( \32737 , RIdf2c128_1878, \16371 );
nor \g453502/U$1 ( \32738 , \32736 , \32737 );
nand \g447919/U$1 ( \32739 , \32724 , \32732 , \32735 , \32738 );
nor \g446359/U$1 ( \32740 , \32719 , \32720 , \32739 );
and \g453487/U$2 ( \32741 , \16377 , RIdec79d0_735);
and \g453487/U$3 ( \32742 , RIe16dad8_2625, \16380 );
nor \g453487/U$1 ( \32743 , \32741 , \32742 );
and \g453482/U$2 ( \32744 , \16334 , RIe1598d0_2396);
and \g453482/U$3 ( \32745 , RIded00d0_831, \16328 );
nor \g453482/U$1 ( \32746 , \32744 , \32745 );
and \g445401/U$2 ( \32747 , \32740 , \32743 , \32746 );
nor \g445401/U$1 ( \32748 , \32747 , \16586 );
or \g444356/U$1 ( \32749 , \32627 , \32688 , \32718 , \32748 );
and \g446326/U$2 ( \32750 , RIfc5add0_6056, \16427 );
and \g446326/U$3 ( \32751 , RIfc92690_6688, \16368 );
and \g449308/U$2 ( \32752 , RIfea95a8_8243, \16344 );
and \g449308/U$3 ( \32753 , \16356 , RIfea7118_8217);
and \g449308/U$4 ( \32754 , RIdf1f270_1731, \16337 );
nor \g449308/U$1 ( \32755 , \32752 , \32753 , \32754 );
and \g455320/U$2 ( \32756 , \16317 , RIfc79fa0_6410);
and \g455320/U$3 ( \32757 , RIfcbe9e8_7191, \16325 );
nor \g455320/U$1 ( \32758 , \32756 , \32757 );
not \g450323/U$3 ( \32759 , \32758 );
not \g450323/U$4 ( \32760 , \16311 );
and \g450323/U$2 ( \32761 , \32759 , \32760 );
and \g450323/U$5 ( \32762 , \16341 , RIfce3018_7605);
nor \g450323/U$1 ( \32763 , \32761 , \32762 );
and \g453356/U$2 ( \32764 , \16377 , RIfc92258_6685);
and \g453356/U$3 ( \32765 , RIfc96740_6734, \16313 );
nor \g453356/U$1 ( \32766 , \32764 , \32765 );
and \g453366/U$2 ( \32767 , \16334 , RIdf24400_1789);
and \g453366/U$3 ( \32768 , RIdf26020_1809, \16380 );
nor \g453366/U$1 ( \32769 , \32767 , \32768 );
nand \g447412/U$1 ( \32770 , \32755 , \32763 , \32766 , \32769 );
nor \g446326/U$1 ( \32771 , \32750 , \32751 , \32770 );
and \g453342/U$2 ( \32772 , \16361 , RIdf19000_1661);
and \g453342/U$3 ( \32773 , RIfc79a00_6406, \16448 );
nor \g453342/U$1 ( \32774 , \32772 , \32773 );
and \g453338/U$2 ( \32775 , \16364 , RIfc79730_6404);
and \g453338/U$3 ( \32776 , RIfce5d18_7637, \16371 );
nor \g453338/U$1 ( \32777 , \32775 , \32776 );
and \g445381/U$2 ( \32778 , \32771 , \32774 , \32777 );
nor \g445381/U$1 ( \32779 , \32778 , \16480 );
and \g446338/U$2 ( \32780 , RIfcbf528_7199, \16427 );
and \g446338/U$3 ( \32781 , RIfc93068_6695, \16368 );
and \g449323/U$2 ( \32782 , RIdee26b8_1040, \16344 );
and \g449323/U$3 ( \32783 , \16356 , RIdee4710_1063);
and \g449323/U$4 ( \32784 , RIded6d18_908, \16337 );
nor \g449323/U$1 ( \32785 , \32782 , \32783 , \32784 );
and \g455218/U$2 ( \32786 , \16317 , RIfc5b640_6062);
and \g455218/U$3 ( \32787 , RIfc5b7a8_6063, \16325 );
nor \g455218/U$1 ( \32788 , \32786 , \32787 );
not \g450337/U$3 ( \32789 , \32788 );
not \g450337/U$4 ( \32790 , \16311 );
and \g450337/U$2 ( \32791 , \32789 , \32790 );
and \g450337/U$5 ( \32792 , \16341 , RIded91a8_934);
nor \g450337/U$1 ( \32793 , \32791 , \32792 );
and \g453402/U$2 ( \32794 , \16377 , RIfcecac8_7715);
and \g453402/U$3 ( \32795 , RIfc931d0_6696, \16313 );
nor \g453402/U$1 ( \32796 , \32794 , \32795 );
and \g453409/U$2 ( \32797 , \16334 , RIdede4a0_993);
and \g453409/U$3 ( \32798 , RIdee07c8_1018, \16380 );
nor \g453409/U$1 ( \32799 , \32797 , \32798 );
nand \g447415/U$1 ( \32800 , \32785 , \32793 , \32796 , \32799 );
nor \g446338/U$1 ( \32801 , \32780 , \32781 , \32800 );
and \g453384/U$2 ( \32802 , \16361 , RIded2998_860);
and \g453384/U$3 ( \32803 , RIfcbf0f0_7196, \16448 );
nor \g453384/U$1 ( \32804 , \32802 , \32803 );
and \g453381/U$2 ( \32805 , \16364 , RIded4e28_886);
and \g453381/U$3 ( \32806 , RIfc792f8_6401, \16371 );
nor \g453381/U$1 ( \32807 , \32805 , \32806 );
and \g445386/U$2 ( \32808 , \32801 , \32804 , \32807 );
nor \g445386/U$1 ( \32809 , \32808 , \16909 );
or \g444179/U$1 ( \32810 , \32749 , \32779 , \32809 );
_DC \g5673/U$1 ( \32811 , \32810 , \16652 );
and \g447196/U$2 ( \32812 , \11521 , RIe1f4f10_4164);
and \g447196/U$3 ( \32813 , RIfc8f288_6651, \11523 );
nor \g447196/U$1 ( \32814 , \32812 , \32813 );
and \g446456/U$2 ( \32815 , RIfc8f828_6655, \8488 );
and \g446456/U$3 ( \32816 , RIf152d80_5402, \8359 );
and \g449470/U$2 ( \32817 , RIf14da88_5343, \8319 );
and \g449470/U$3 ( \32818 , \8326 , RIfc8faf8_6657);
and \g449470/U$4 ( \32819 , RIf155648_5431, \8409 );
nor \g449470/U$1 ( \32820 , \32817 , \32818 , \32819 );
and \g453953/U$2 ( \32821 , \8335 , RIe1eda58_4081);
and \g453953/U$3 ( \32822 , RIfc445d0_5800, \8340 );
nor \g453953/U$1 ( \32823 , \32821 , \32822 );
and \g453952/U$2 ( \32824 , \8404 , RIe1f9dd0_4220);
and \g453952/U$3 ( \32825 , RIfebfad8_8301, \8351 );
nor \g453952/U$1 ( \32826 , \32824 , \32825 );
and \g454322/U$2 ( \32827 , \8313 , RIfc7cca0_6442);
and \g454322/U$3 ( \32828 , RIfebf970_8300, \8323 );
nor \g454322/U$1 ( \32829 , \32827 , \32828 );
not \g450489/U$3 ( \32830 , \32829 );
not \g450489/U$4 ( \32831 , \8328 );
and \g450489/U$2 ( \32832 , \32830 , \32831 );
and \g450489/U$5 ( \32833 , \8417 , RIfe82c50_7832);
nor \g450489/U$1 ( \32834 , \32832 , \32833 );
nand \g447983/U$1 ( \32835 , \32820 , \32823 , \32826 , \32834 );
nor \g446456/U$1 ( \32836 , \32815 , \32816 , \32835 );
not \g444887/U$3 ( \32837 , \32836 );
not \g444887/U$4 ( \32838 , \8621 );
and \g444887/U$2 ( \32839 , \32837 , \32838 );
and \g446463/U$2 ( \32840 , RIe1a2968_3227, \8373 );
and \g446463/U$3 ( \32841 , RIe1a5668_3259, \8383 );
and \g449481/U$2 ( \32842 , RIe1bb328_3507, \8326 );
and \g449481/U$3 ( \32843 , \8531 , RIe1f77d8_4193);
and \g449481/U$4 ( \32844 , RIe1fe420_4270, \8488 );
nor \g449481/U$1 ( \32845 , \32842 , \32843 , \32844 );
and \g454003/U$2 ( \32846 , \8356 , RIe1f0320_4110);
and \g454003/U$3 ( \32847 , RIe2043c0_4338, \8359 );
nor \g454003/U$1 ( \32848 , \32846 , \32847 );
and \g455062/U$2 ( \32849 , \8313 , RIe225fc0_4722);
and \g455062/U$3 ( \32850 , RIe178668_2747, \8323 );
nor \g455062/U$1 ( \32851 , \32849 , \32850 );
not \g450500/U$3 ( \32852 , \32851 );
not \g450500/U$4 ( \32853 , \8376 );
and \g450500/U$2 ( \32854 , \32852 , \32853 );
and \g450500/U$5 ( \32855 , \8340 , RIe1d4828_3795);
nor \g450500/U$1 ( \32856 , \32854 , \32855 );
and \g453995/U$2 ( \32857 , \8378 , RIe21abc0_4594);
and \g453995/U$3 ( \32858 , RIe18c168_2971, \8417 );
nor \g453995/U$1 ( \32859 , \32857 , \32858 );
nand \g447986/U$1 ( \32860 , \32845 , \32848 , \32856 , \32859 );
nor \g446463/U$1 ( \32861 , \32840 , \32841 , \32860 );
and \g453975/U$2 ( \32862 , \8335 , RIe1707d8_2657);
and \g453975/U$3 ( \32863 , RIe1a8368_3291, \8351 );
nor \g453975/U$1 ( \32864 , \32862 , \32863 );
and \g453989/U$2 ( \32865 , \8317 , RIe1ae1a0_3358);
and \g453989/U$3 ( \32866 , RIe19fc68_3195, \8404 );
nor \g453989/U$1 ( \32867 , \32865 , \32866 );
and \g445484/U$2 ( \32868 , \32861 , \32864 , \32867 );
nor \g445484/U$1 ( \32869 , \32868 , \8651 );
nor \g444887/U$1 ( \32870 , \32839 , \32869 );
and \g447192/U$2 ( \32871 , \13486 , RIe1f2d50_4140);
and \g447192/U$3 ( \32872 , RIfcb3b88_7067, \13488 );
nor \g447192/U$1 ( \32873 , \32871 , \32872 );
nand \g444440/U$1 ( \32874 , \32814 , \32870 , \32873 );
and \g454079/U$2 ( \32875 , \8531 , RIe1cc128_3699);
and \g454079/U$3 ( \32876 , RIe1cee28_3731, \8488 );
nor \g454079/U$1 ( \32877 , \32875 , \32876 );
and \g446489/U$2 ( \32878 , RIe1da228_3859, \8414 );
and \g446489/U$3 ( \32879 , RIe1c9428_3667, \8356 );
and \g449510/U$2 ( \32880 , RIe1dcf28_3891, \8409 );
and \g449510/U$3 ( \32881 , \8373 , RIe1e5628_3987);
and \g449510/U$4 ( \32882 , RIe1e8328_4019, \8383 );
nor \g449510/U$1 ( \32883 , \32880 , \32881 , \32882 );
and \g454099/U$2 ( \32884 , \8335 , RIe1be028_3539);
and \g454099/U$3 ( \32885 , RIe1c6728_3635, \8340 );
nor \g454099/U$1 ( \32886 , \32884 , \32885 );
and \g454095/U$2 ( \32887 , \8404 , RIe1e2928_3955);
and \g454095/U$3 ( \32888 , RIe1eb028_4051, \8351 );
nor \g454095/U$1 ( \32889 , \32887 , \32888 );
and \g454810/U$2 ( \32890 , \8313 , RIe1c0d28_3571);
and \g454810/U$3 ( \32891 , RIe1c3a28_3603, \8323 );
nor \g454810/U$1 ( \32892 , \32890 , \32891 );
not \g454809/U$1 ( \32893 , \32892 );
and \g450528/U$2 ( \32894 , \32893 , \8316 );
and \g450528/U$3 ( \32895 , RIe1dfc28_3923, \8417 );
nor \g450528/U$1 ( \32896 , \32894 , \32895 );
nand \g448252/U$1 ( \32897 , \32883 , \32886 , \32889 , \32896 );
nor \g446489/U$1 ( \32898 , \32878 , \32879 , \32897 );
and \g454080/U$2 ( \32899 , \8378 , RIe1d7528_3827);
and \g454080/U$3 ( \32900 , RIe1d1b28_3763, \8359 );
nor \g454080/U$1 ( \32901 , \32899 , \32900 );
nand \g445698/U$1 ( \32902 , \32877 , \32898 , \32901 );
and \g444810/U$2 ( \32903 , \32902 , \8478 );
and \g449498/U$2 ( \32904 , RIe1ac148_3335, \8317 );
and \g449498/U$3 ( \32905 , \8326 , RIfc7ba58_6429);
and \g449498/U$4 ( \32906 , RIfc8ff30_6660, \8409 );
nor \g449498/U$1 ( \32907 , \32904 , \32905 , \32906 );
and \g454053/U$2 ( \32908 , \8335 , RIe1aa960_3318);
and \g454053/U$3 ( \32909 , RIfcdb5c0_7518, \8340 );
nor \g454053/U$1 ( \32910 , \32908 , \32909 );
and \g454049/U$2 ( \32911 , \8404 , RIe1b6fa8_3459);
and \g454049/U$3 ( \32912 , RIfc7bff8_6433, \8351 );
nor \g454049/U$1 ( \32913 , \32911 , \32912 );
and \g455400/U$2 ( \32914 , \8313 , RIe1b9000_3482);
and \g455400/U$3 ( \32915 , RIfc44030_5796, \8323 );
nor \g455400/U$1 ( \32916 , \32914 , \32915 );
not \g450515/U$3 ( \32917 , \32916 );
not \g450515/U$4 ( \32918 , \8328 );
and \g450515/U$2 ( \32919 , \32917 , \32918 );
and \g450515/U$5 ( \32920 , \8417 , RIfcbdd40_7182);
nor \g450515/U$1 ( \32921 , \32919 , \32920 );
nand \g447994/U$1 ( \32922 , \32907 , \32910 , \32913 , \32921 );
and \g444810/U$3 ( \32923 , \8482 , \32922 );
nor \g444810/U$1 ( \32924 , \32903 , \32923 );
and \g447219/U$2 ( \32925 , \8521 , RIe1b0798_3385);
and \g447219/U$3 ( \32926 , RIe1b2520_3406, \8525 );
nor \g447219/U$1 ( \32927 , \32925 , \32926 );
and \g447218/U$2 ( \32928 , \10290 , RIfc43d60_5794);
and \g447218/U$3 ( \32929 , RIfcbe178_7185, \10293 );
nor \g447218/U$1 ( \32930 , \32928 , \32929 );
and \g447220/U$2 ( \32931 , \8974 , RIe1b3d08_3423);
and \g447220/U$3 ( \32932 , RIe1b50b8_3437, \8976 );
nor \g447220/U$1 ( \32933 , \32931 , \32932 );
nand \g444547/U$1 ( \32934 , \32924 , \32927 , \32930 , \32933 );
and \g446431/U$2 ( \32935 , RIe191b68_3035, \8412 );
and \g446431/U$3 ( \32936 , RIe183a68_2875, \8356 );
and \g449440/U$2 ( \32937 , RIe17e068_2811, \8319 );
and \g449440/U$3 ( \32938 , \8326 , RIe180d68_2843);
and \g449440/U$4 ( \32939 , RIe194868_3067, \8409 );
nor \g449440/U$1 ( \32940 , \32937 , \32938 , \32939 );
and \g453845/U$2 ( \32941 , \8335 , RIe17b368_2779);
and \g453845/U$3 ( \32942 , RIfc7d948_6451, \8340 );
nor \g453845/U$1 ( \32943 , \32941 , \32942 );
and \g453842/U$2 ( \32944 , \8404 , RIe197568_3099);
and \g453842/U$3 ( \32945 , RIe19cf68_3163, \8351 );
nor \g453842/U$1 ( \32946 , \32944 , \32945 );
and \g455111/U$2 ( \32947 , \8313 , RIfc8d7d0_6632);
and \g455111/U$3 ( \32948 , RIe19a268_3131, \8323 );
nor \g455111/U$1 ( \32949 , \32947 , \32948 );
not \g450457/U$3 ( \32950 , \32949 );
not \g450457/U$4 ( \32951 , \8328 );
and \g450457/U$2 ( \32952 , \32950 , \32951 );
and \g450457/U$5 ( \32953 , \8417 , RIfc561e0_6002);
nor \g450457/U$1 ( \32954 , \32952 , \32953 );
nand \g447966/U$1 ( \32955 , \32940 , \32943 , \32946 , \32954 );
nor \g446431/U$1 ( \32956 , \32935 , \32936 , \32955 );
and \g453821/U$2 ( \32957 , \8378 , RIe18ee68_3003);
and \g453821/U$3 ( \32958 , RIe189468_2939, \8359 );
nor \g453821/U$1 ( \32959 , \32957 , \32958 );
and \g453829/U$2 ( \32960 , \8531 , RIf143330_5224);
and \g453829/U$3 ( \32961 , RIe186768_2907, \8488 );
nor \g453829/U$1 ( \32962 , \32960 , \32961 );
and \g445451/U$2 ( \32963 , \32956 , \32959 , \32962 );
nor \g445451/U$1 ( \32964 , \32963 , \8589 );
and \g446440/U$2 ( \32965 , RIfc7dc18_6453, \8414 );
and \g446440/U$3 ( \32966 , RIe173208_2687, \8356 );
and \g449454/U$2 ( \32967 , RIfc8e8b0_6644, \8319 );
and \g449454/U$3 ( \32968 , \8324 , RIfc45ae8_5815);
and \g449454/U$4 ( \32969 , RIfc45f20_5818, \8409 );
nor \g449454/U$1 ( \32970 , \32967 , \32968 , \32969 );
and \g453897/U$2 ( \32971 , \8335 , RIfc45980_5814);
and \g453897/U$3 ( \32972 , RIfc8e478_6641, \8340 );
nor \g453897/U$1 ( \32973 , \32971 , \32972 );
and \g453890/U$2 ( \32974 , \8404 , RIe175698_2713);
and \g453890/U$3 ( \32975 , RIfc564b0_6004, \8351 );
nor \g453890/U$1 ( \32976 , \32974 , \32975 );
and \g454550/U$2 ( \32977 , \8313 , RIfc461f0_5820);
and \g454550/U$3 ( \32978 , RIfcd6700_7462, \8323 );
nor \g454550/U$1 ( \32979 , \32977 , \32978 );
not \g450472/U$3 ( \32980 , \32979 );
not \g450472/U$4 ( \32981 , \8328 );
and \g450472/U$2 ( \32982 , \32980 , \32981 );
and \g450472/U$5 ( \32983 , \8417 , RIfc46088_5819);
nor \g450472/U$1 ( \32984 , \32982 , \32983 );
nand \g447973/U$1 ( \32985 , \32970 , \32973 , \32976 , \32984 );
nor \g446440/U$1 ( \32986 , \32965 , \32966 , \32985 );
and \g453874/U$2 ( \32987 , \8378 , RIfcd69d0_7464);
and \g453874/U$3 ( \32988 , RIfc98630_6756, \8359 );
nor \g453874/U$1 ( \32989 , \32987 , \32988 );
and \g453868/U$2 ( \32990 , \8531 , RIfc7d510_6448);
and \g453868/U$3 ( \32991 , RIfcc2a98_7237, \8488 );
nor \g453868/U$1 ( \32992 , \32990 , \32991 );
and \g445459/U$2 ( \32993 , \32986 , \32989 , \32992 );
nor \g445459/U$1 ( \32994 , \32993 , \8558 );
or \g444313/U$1 ( \32995 , \32874 , \32934 , \32964 , \32994 );
and \g446411/U$2 ( \32996 , RIe217ec0_4562, \8412 );
and \g446411/U$3 ( \32997 , RIe20f7c0_4466, \8356 );
and \g449413/U$2 ( \32998 , RIe209dc0_4402, \8319 );
and \g449413/U$3 ( \32999 , \8326 , RIe20cac0_4434);
and \g449413/U$4 ( \33000 , RIe21d8c0_4626, \8409 );
nor \g449413/U$1 ( \33001 , \32998 , \32999 , \33000 );
and \g453746/U$2 ( \33002 , \8335 , RIe2070c0_4370);
and \g453746/U$3 ( \33003 , RIfc7d240_6446, \8340 );
nor \g453746/U$1 ( \33004 , \33002 , \33003 );
and \g453752/U$2 ( \33005 , \8404 , RIe2205c0_4658);
and \g453752/U$3 ( \33006 , RIfe82ae8_7831, \8351 );
nor \g453752/U$1 ( \33007 , \33005 , \33006 );
and \g454438/U$2 ( \33008 , \8313 , RIf16ba10_5684);
and \g454438/U$3 ( \33009 , RIe2232c0_4690, \8323 );
nor \g454438/U$1 ( \33010 , \33008 , \33009 );
not \g450430/U$3 ( \33011 , \33010 );
not \g450430/U$4 ( \33012 , \8328 );
and \g450430/U$2 ( \33013 , \33011 , \33012 );
and \g450430/U$5 ( \33014 , \8417 , RIfcd24e8_7415);
nor \g450430/U$1 ( \33015 , \33013 , \33014 );
nand \g447953/U$1 ( \33016 , \33001 , \33004 , \33007 , \33015 );
nor \g446411/U$1 ( \33017 , \32996 , \32997 , \33016 );
and \g453736/U$2 ( \33018 , \8378 , RIe2151c0_4530);
and \g453736/U$3 ( \33019 , RIfebf268_8295, \8359 );
nor \g453736/U$1 ( \33020 , \33018 , \33019 );
and \g453730/U$2 ( \33021 , \8531 , RIf168d10_5652);
and \g453730/U$3 ( \33022 , RIe2124c0_4498, \8488 );
nor \g453730/U$1 ( \33023 , \33021 , \33022 );
and \g445439/U$2 ( \33024 , \33017 , \33020 , \33023 );
nor \g445439/U$1 ( \33025 , \33024 , \8368 );
and \g446420/U$2 ( \33026 , RIfc453e0_5810, \8412 );
and \g446420/U$3 ( \33027 , RIe1fb888_4239, \8356 );
and \g449424/U$2 ( \33028 , RIfca2518_6869, \8319 );
and \g449424/U$3 ( \33029 , \8324 , RIf15b318_5497);
and \g449424/U$4 ( \33030 , RIf164120_5598, \8409 );
nor \g449424/U$1 ( \33031 , \33028 , \33029 , \33030 );
and \g453797/U$2 ( \33032 , \8335 , RIfc8f120_6650);
and \g453797/U$3 ( \33033 , RIfebf3d0_8296, \8340 );
nor \g453797/U$1 ( \33034 , \33032 , \33033 );
and \g453793/U$2 ( \33035 , \8404 , RIfebf538_8297);
and \g453793/U$3 ( \33036 , RIf166e20_5630, \8351 );
nor \g453793/U$1 ( \33037 , \33035 , \33036 );
and \g455080/U$2 ( \33038 , \8313 , RIfebf808_8299);
and \g455080/U$3 ( \33039 , RIfebf6a0_8298, \8323 );
nor \g455080/U$1 ( \33040 , \33038 , \33039 );
not \g450443/U$3 ( \33041 , \33040 );
not \g450443/U$4 ( \33042 , \8328 );
and \g450443/U$2 ( \33043 , \33041 , \33042 );
and \g450443/U$5 ( \33044 , \8417 , RIfc8eb80_6646);
nor \g450443/U$1 ( \33045 , \33043 , \33044 );
nand \g447960/U$1 ( \33046 , \33031 , \33034 , \33037 , \33045 );
nor \g446420/U$1 ( \33047 , \33026 , \33027 , \33046 );
and \g453781/U$2 ( \33048 , \8378 , RIf161b28_5571);
and \g453781/U$3 ( \33049 , RIf15fc38_5549, \8359 );
nor \g453781/U$1 ( \33050 , \33048 , \33049 );
and \g453775/U$2 ( \33051 , \8531 , RIe1fc968_4251);
and \g453775/U$3 ( \33052 , RIf15dd48_5527, \8488 );
nor \g453775/U$1 ( \33053 , \33051 , \33052 );
and \g445442/U$2 ( \33054 , \33047 , \33050 , \33053 );
nor \g445442/U$1 ( \33055 , \33054 , \8422 );
or \g444237/U$1 ( \33056 , \32995 , \33025 , \33055 );
_DC \g56f7/U$1 ( \33057 , \33056 , \8654 );
and \g452760/U$2 ( \33058 , \16371 , RIfc48518_5845);
and \g452760/U$3 ( \33059 , RIe151338_2301, \16427 );
nor \g452760/U$1 ( \33060 , \33058 , \33059 );
and \g446205/U$2 ( \33061 , RIfc3f260_5744, \16432 );
and \g446205/U$3 ( \33062 , RIe145f38_2173, \16361 );
and \g449147/U$2 ( \33063 , RIe162138_2493, \16321 );
and \g449147/U$3 ( \33064 , \16326 , RIe164e38_2525);
and \g449147/U$4 ( \33065 , RIe14b938_2237, \16398 );
nor \g449147/U$1 ( \33066 , \33063 , \33064 , \33065 );
and \g455227/U$2 ( \33067 , \16317 , RIe15c738_2429);
and \g455227/U$3 ( \33068 , RIfc999e0_6770, \16325 );
nor \g455227/U$1 ( \33069 , \33067 , \33068 );
not \g450162/U$3 ( \33070 , \33069 );
not \g450162/U$4 ( \33071 , \16330 );
and \g450162/U$2 ( \33072 , \33070 , \33071 );
and \g450162/U$5 ( \33073 , \16339 , RIfc99e18_6773);
nor \g450162/U$1 ( \33074 , \33072 , \33073 );
and \g452771/U$2 ( \33075 , \16377 , RIe15f438_2461);
and \g452771/U$3 ( \33076 , RIee370f0_5085, \16313 );
nor \g452771/U$1 ( \33077 , \33075 , \33076 );
and \g452773/U$2 ( \33078 , \16334 , RIe154038_2333);
and \g452773/U$3 ( \33079 , RIe156d38_2365, \16380 );
nor \g452773/U$1 ( \33080 , \33078 , \33079 );
nand \g447378/U$1 ( \33081 , \33066 , \33074 , \33077 , \33080 );
nor \g446205/U$1 ( \33082 , \33061 , \33062 , \33081 );
and \g452766/U$2 ( \33083 , \16364 , RIe148c38_2205);
and \g452766/U$3 ( \33084 , RIe14e638_2269, \16368 );
nor \g452766/U$1 ( \33085 , \33083 , \33084 );
nand \g445625/U$1 ( \33086 , \33060 , \33082 , \33085 );
and \g444861/U$2 ( \33087 , \33086 , \16390 );
and \g449140/U$2 ( \33088 , RIee33040_5039, \16321 );
and \g449140/U$3 ( \33089 , \16328 , RIee34288_5052);
and \g449140/U$4 ( \33090 , RIfec0ff0_8316, \16337 );
nor \g449140/U$1 ( \33091 , \33088 , \33089 , \33090 );
and \g454989/U$2 ( \33092 , \16317 , RIdf3e9e0_2089);
and \g454989/U$3 ( \33093 , RIfe86b98_7877, \16325 );
nor \g454989/U$1 ( \33094 , \33092 , \33093 );
not \g450154/U$3 ( \33095 , \33094 );
not \g450154/U$4 ( \33096 , \16330 );
and \g450154/U$2 ( \33097 , \33095 , \33096 );
and \g450154/U$5 ( \33098 , \16341 , RIdf35200_1981);
nor \g450154/U$1 ( \33099 , \33097 , \33098 );
and \g452742/U$2 ( \33100 , \16377 , RIfcd99a0_7498);
and \g452742/U$3 ( \33101 , RIee31f60_5027, \16313 );
nor \g452742/U$1 ( \33102 , \33100 , \33101 );
and \g452745/U$2 ( \33103 , \16334 , RIdf3a4f8_2040);
and \g452745/U$3 ( \33104 , RIfe86a30_7876, \16380 );
nor \g452745/U$1 ( \33105 , \33103 , \33104 );
nand \g447376/U$1 ( \33106 , \33091 , \33099 , \33102 , \33105 );
and \g444861/U$3 ( \33107 , \16394 , \33106 );
nor \g444861/U$1 ( \33108 , \33087 , \33107 );
and \g446977/U$2 ( \33109 , \16419 , RIfec0e88_8315);
and \g446977/U$3 ( \33110 , RIdf30d18_1932, \16422 );
nor \g446977/U$1 ( \33111 , \33109 , \33110 );
and \g446974/U$2 ( \33112 , \16429 , RIee2f530_4997);
and \g446974/U$3 ( \33113 , RIfcc3470_7244, \16434 );
nor \g446974/U$1 ( \33114 , \33112 , \33113 );
and \g446975/U$2 ( \33115 , \16438 , RIee2d370_4973);
and \g446975/U$3 ( \33116 , RIfc7fdd8_6477, \16441 );
nor \g446975/U$1 ( \33117 , \33115 , \33116 );
nand \g444630/U$1 ( \33118 , \33108 , \33111 , \33114 , \33117 );
and \g452817/U$2 ( \33119 , \16371 , RIdf2c290_1879);
and \g452817/U$3 ( \33120 , RIdf37c30_2011, \16427 );
nor \g452817/U$1 ( \33121 , \33119 , \33120 );
and \g446216/U$2 ( \33122 , RIe143238_2141, \16448 );
and \g446216/U$3 ( \33123 , RIde7bb48_193, \16361 );
and \g449165/U$2 ( \33124 , RIdecd538_800, \16319 );
and \g449165/U$3 ( \33125 , \16328 , RIded0238_832);
and \g449165/U$4 ( \33126 , RIdee6d08_1090, \16398 );
nor \g449165/U$1 ( \33127 , \33124 , \33125 , \33126 );
and \g455044/U$2 ( \33128 , \16317 , RIde95c00_320);
and \g455044/U$3 ( \33129 , RIdeb4038_512, \16325 );
nor \g455044/U$1 ( \33130 , \33128 , \33129 );
not \g450179/U$3 ( \33131 , \33130 );
not \g450179/U$4 ( \33132 , \16330 );
and \g450179/U$2 ( \33133 , \33131 , \33132 );
and \g450179/U$5 ( \33134 , \16341 , RIdf00208_1378);
nor \g450179/U$1 ( \33135 , \33133 , \33134 );
and \g452828/U$2 ( \33136 , \16377 , RIdec7b38_736);
and \g452828/U$3 ( \33137 , RIdeca838_768, \16313 );
nor \g452828/U$1 ( \33138 , \33136 , \33137 );
and \g452831/U$2 ( \33139 , \16334 , RIe159a38_2397);
and \g452831/U$3 ( \33140 , RIe16dc40_2626, \16380 );
nor \g452831/U$1 ( \33141 , \33139 , \33140 );
nand \g447384/U$1 ( \33142 , \33127 , \33135 , \33138 , \33141 );
nor \g446216/U$1 ( \33143 , \33122 , \33123 , \33142 );
and \g452821/U$2 ( \33144 , \16364 , RIdedba70_963);
and \g452821/U$3 ( \33145 , RIdf1cb10_1703, \16368 );
nor \g452821/U$1 ( \33146 , \33144 , \33145 );
nand \g445633/U$1 ( \33147 , \33121 , \33143 , \33146 );
and \g444786/U$2 ( \33148 , \33147 , \16752 );
and \g449156/U$2 ( \33149 , RIdf08908_1474, \16485 );
and \g449156/U$3 ( \33150 , \16356 , RIdf0b608_1506);
and \g449156/U$4 ( \33151 , RIdeef408_1186, \16398 );
nor \g449156/U$1 ( \33152 , \33149 , \33150 , \33151 );
and \g455025/U$2 ( \33153 , \16317 , RIdf13d08_1602);
and \g455025/U$3 ( \33154 , RIdf16a08_1634, \16325 );
nor \g455025/U$1 ( \33155 , \33153 , \33154 );
not \g450170/U$3 ( \33156 , \33155 );
not \g450170/U$4 ( \33157 , \16311 );
and \g450170/U$2 ( \33158 , \33156 , \33157 );
and \g450170/U$5 ( \33159 , \16339 , RIdef2108_1218);
nor \g450170/U$1 ( \33160 , \33158 , \33159 );
and \g452800/U$2 ( \33161 , \16377 , RIdf0e308_1538);
and \g452800/U$3 ( \33162 , RIdf11008_1570, \16313 );
nor \g452800/U$1 ( \33163 , \33161 , \33162 );
and \g452802/U$2 ( \33164 , \16334 , RIdf02f08_1410);
and \g452802/U$3 ( \33165 , RIdf05c08_1442, \16380 );
nor \g452802/U$1 ( \33166 , \33164 , \33165 );
nand \g447380/U$1 ( \33167 , \33152 , \33160 , \33163 , \33166 );
and \g444786/U$3 ( \33168 , \16750 , \33167 );
nor \g444786/U$1 ( \33169 , \33148 , \33168 );
and \g446988/U$2 ( \33170 , \19208 , RIdee9a08_1122);
and \g446988/U$3 ( \33171 , RIdef7b08_1282, \19210 );
nor \g446988/U$1 ( \33172 , \33170 , \33171 );
and \g446989/U$2 ( \33173 , \19213 , RIdeec708_1154);
and \g446989/U$3 ( \33174 , RIdef4e08_1250, \19215 );
nor \g446989/U$1 ( \33175 , \33173 , \33174 );
and \g446987/U$2 ( \33176 , \19218 , RIdefa808_1314);
and \g446987/U$3 ( \33177 , RIdefd508_1346, \19220 );
nor \g446987/U$1 ( \33178 , \33176 , \33177 );
nand \g444633/U$1 ( \33179 , \33169 , \33172 , \33175 , \33178 );
and \g446193/U$2 ( \33180 , RIee254e0_4883, \16326 );
and \g446193/U$3 ( \33181 , RIee231b8_4858, \16377 );
and \g449125/U$2 ( \33182 , RIded6e80_909, \16337 );
and \g449125/U$3 ( \33183 , \16341 , RIded9310_935);
and \g449125/U$4 ( \33184 , RIdee2820_1041, \16485 );
nor \g449125/U$1 ( \33185 , \33182 , \33183 , \33184 );
and \g455359/U$2 ( \33186 , \16331 , RIfc464c0_5822);
and \g455359/U$3 ( \33187 , RIfcc3038_7241, \20087 );
nor \g455359/U$1 ( \33188 , \33186 , \33187 );
not \g450139/U$3 ( \33189 , \33188 );
not \g450139/U$4 ( \33190 , \16351 );
and \g450139/U$2 ( \33191 , \33189 , \33190 );
and \g450139/U$5 ( \33192 , \16356 , RIfe86fd0_7880);
nor \g450139/U$1 ( \33193 , \33191 , \33192 );
and \g452691/U$2 ( \33194 , \16361 , RIded2b00_861);
and \g452691/U$3 ( \33195 , RIded4f90_887, \16364 );
nor \g452691/U$1 ( \33196 , \33194 , \33195 );
and \g452685/U$2 ( \33197 , \16427 , RIfc98a68_6759);
and \g452685/U$3 ( \33198 , RIfc55da8_5999, \16448 );
nor \g452685/U$1 ( \33199 , \33197 , \33198 );
nand \g447788/U$1 ( \33200 , \33185 , \33193 , \33196 , \33199 );
nor \g446193/U$1 ( \33201 , \33180 , \33181 , \33200 );
and \g452672/U$2 ( \33202 , \16334 , RIdede608_994);
and \g452672/U$3 ( \33203 , RIee23b90_4865, \16313 );
nor \g452672/U$1 ( \33204 , \33202 , \33203 );
and \g452671/U$2 ( \33205 , \16380 , RIdee0930_1019);
and \g452671/U$3 ( \33206 , RIee246d0_4873, \16321 );
nor \g452671/U$1 ( \33207 , \33205 , \33206 );
and \g445287/U$2 ( \33208 , \33201 , \33204 , \33207 );
nor \g445287/U$1 ( \33209 , \33208 , \16909 );
and \g446194/U$2 ( \33210 , RIfc8cb28_6623, \16448 );
and \g446194/U$3 ( \33211 , RIdf22948_1770, \16371 );
and \g449133/U$2 ( \33212 , RIdf27da8_1830, \16485 );
and \g449133/U$3 ( \33213 , \16354 , RIdf29f68_1854);
and \g449133/U$4 ( \33214 , RIdf1f3d8_1732, \16398 );
nor \g449133/U$1 ( \33215 , \33212 , \33213 , \33214 );
and \g454974/U$2 ( \33216 , \16317 , RIfc8c858_6621);
and \g454974/U$3 ( \33217 , RIfcd2a88_7419, \16325 );
nor \g454974/U$1 ( \33218 , \33216 , \33217 );
not \g450147/U$3 ( \33219 , \33218 );
not \g450147/U$4 ( \33220 , \16311 );
and \g450147/U$2 ( \33221 , \33219 , \33220 );
and \g450147/U$5 ( \33222 , \16339 , RIdf21430_1755);
nor \g450147/U$1 ( \33223 , \33221 , \33222 );
and \g452714/U$2 ( \33224 , \16377 , RIfcd6430_7460);
and \g452714/U$3 ( \33225 , RIfc47ca8_5839, \16313 );
nor \g452714/U$1 ( \33226 , \33224 , \33225 );
and \g452717/U$2 ( \33227 , \16334 , RIdf24568_1790);
and \g452717/U$3 ( \33228 , RIdf26188_1810, \16380 );
nor \g452717/U$1 ( \33229 , \33227 , \33228 );
nand \g447373/U$1 ( \33230 , \33215 , \33223 , \33226 , \33229 );
nor \g446194/U$1 ( \33231 , \33210 , \33211 , \33230 );
and \g452704/U$2 ( \33232 , \16364 , RIfec0bb8_8313);
and \g452704/U$3 ( \33233 , RIfc475a0_5834, \16368 );
nor \g452704/U$1 ( \33234 , \33232 , \33233 );
and \g452709/U$2 ( \33235 , \16361 , RIfe868c8_7875);
and \g452709/U$3 ( \33236 , RIfcdb188_7515, \16427 );
nor \g452709/U$1 ( \33237 , \33235 , \33236 );
and \g445289/U$2 ( \33238 , \33231 , \33234 , \33237 );
nor \g445289/U$1 ( \33239 , \33238 , \16480 );
or \g444331/U$1 ( \33240 , \33118 , \33179 , \33209 , \33239 );
and \g446178/U$2 ( \33241 , RIdeb1338_480, \16427 );
and \g446178/U$3 ( \33242 , RIdeae638_448, \16368 );
and \g449112/U$2 ( \33243 , RIdec2138_672, \16321 );
and \g449112/U$3 ( \33244 , \16328 , RIdec4e38_704);
and \g449112/U$4 ( \33245 , RIdea9700_416, \16337 );
nor \g449112/U$1 ( \33246 , \33243 , \33244 , \33245 );
and \g454947/U$2 ( \33247 , \16317 , RIdebc738_608);
and \g454947/U$3 ( \33248 , RIfc49490_5856, \16325 );
nor \g454947/U$1 ( \33249 , \33247 , \33248 );
not \g450125/U$3 ( \33250 , \33249 );
not \g450125/U$4 ( \33251 , \16330 );
and \g450125/U$2 ( \33252 , \33250 , \33251 );
and \g450125/U$5 ( \33253 , \16341 , RIfc8b610_6608);
nor \g450125/U$1 ( \33254 , \33252 , \33253 );
and \g452632/U$2 ( \33255 , \16377 , RIdebf438_640);
and \g452632/U$3 ( \33256 , RIee1fc48_4820, \16313 );
nor \g452632/U$1 ( \33257 , \33255 , \33256 );
and \g452634/U$2 ( \33258 , \16334 , RIdeb6d38_544);
and \g452634/U$3 ( \33259 , RIdeb9a38_576, \16380 );
nor \g452634/U$1 ( \33260 , \33258 , \33259 );
nand \g447364/U$1 ( \33261 , \33246 , \33254 , \33257 , \33260 );
nor \g446178/U$1 ( \33262 , \33241 , \33242 , \33261 );
and \g452624/U$2 ( \33263 , \16361 , RIde9c500_352);
and \g452624/U$3 ( \33264 , RIfc48ef0_5852, \16448 );
nor \g452624/U$1 ( \33265 , \33263 , \33264 );
and \g452622/U$2 ( \33266 , \16364 , RIdea2e00_384);
and \g452622/U$3 ( \33267 , RIfcd9b08_7499, \16371 );
nor \g452622/U$1 ( \33268 , \33266 , \33267 );
and \g445278/U$2 ( \33269 , \33262 , \33265 , \33268 );
nor \g445278/U$1 ( \33270 , \33269 , \16618 );
and \g446183/U$2 ( \33271 , RIfc8b8e0_6610, \16427 );
and \g446183/U$3 ( \33272 , RIfce4530_7620, \16368 );
and \g449118/U$2 ( \33273 , RIee1b8c8_4772, \16321 );
and \g449118/U$3 ( \33274 , \16328 , RIee1c9a8_4784);
and \g449118/U$4 ( \33275 , RIe16b210_2596, \16398 );
nor \g449118/U$1 ( \33276 , \33273 , \33274 , \33275 );
and \g454959/U$2 ( \33277 , \16317 , RIde8cee8_277);
and \g454959/U$3 ( \33278 , RIfe86e68_7879, \16325 );
nor \g454959/U$1 ( \33279 , \33277 , \33278 );
not \g450132/U$3 ( \33280 , \33279 );
not \g450132/U$4 ( \33281 , \16330 );
and \g450132/U$2 ( \33282 , \33280 , \33281 );
and \g450132/U$5 ( \33283 , \16341 , RIfc8ba48_6611);
nor \g450132/U$1 ( \33284 , \33282 , \33283 );
and \g452657/U$2 ( \33285 , \16377 , RIfcdad50_7512);
and \g452657/U$3 ( \33286 , RIfc80918_6485, \16313 );
nor \g452657/U$1 ( \33287 , \33285 , \33286 );
and \g452658/U$2 ( \33288 , \16334 , RIfec0d20_8314);
and \g452658/U$3 ( \33289 , RIfe86d00_7878, \16380 );
nor \g452658/U$1 ( \33290 , \33288 , \33289 );
nand \g447368/U$1 ( \33291 , \33276 , \33284 , \33287 , \33290 );
nor \g446183/U$1 ( \33292 , \33271 , \33272 , \33291 );
and \g452651/U$2 ( \33293 , \16361 , RIe1679d0_2556);
and \g452651/U$3 ( \33294 , RIde81098_219, \16448 );
nor \g452651/U$1 ( \33295 , \33293 , \33294 );
and \g452647/U$2 ( \33296 , \16364 , RIe1698c0_2578);
and \g452647/U$3 ( \33297 , RIfcd2d58_7421, \16371 );
nor \g452647/U$1 ( \33298 , \33296 , \33297 );
and \g445281/U$2 ( \33299 , \33292 , \33295 , \33298 );
nor \g445281/U$1 ( \33300 , \33299 , \16649 );
or \g444277/U$1 ( \33301 , \33240 , \33270 , \33300 );
_DC \g577c/U$1 ( \33302 , \33301 , \16652 );
and \g449203/U$2 ( \33303 , RIe218028_4563, \8412 );
and \g449203/U$3 ( \33304 , \8409 , RIe21da28_4627);
and \g449203/U$4 ( \33305 , RIe212628_4499, \8486 );
nor \g449203/U$1 ( \33306 , \33303 , \33304 , \33305 );
and \g455131/U$2 ( \33307 , \8313 , RIf16bb78_5685);
and \g455131/U$3 ( \33308 , RIe223428_4691, \8323 );
nor \g455131/U$1 ( \33309 , \33307 , \33308 );
not \g450216/U$3 ( \33310 , \33309 );
not \g450216/U$4 ( \33311 , \8328 );
and \g450216/U$2 ( \33312 , \33310 , \33311 );
and \g450216/U$5 ( \33313 , \8359 , RIf16a0c0_5666);
nor \g450216/U$1 ( \33314 , \33312 , \33313 );
and \g452966/U$2 ( \33315 , \8404 , RIe220728_4659);
and \g452966/U$3 ( \33316 , RIf16c988_5695, \8351 );
nor \g452966/U$1 ( \33317 , \33315 , \33316 );
and \g452970/U$2 ( \33318 , \8378 , RIe215328_4531);
and \g452970/U$3 ( \33319 , RIf16aa98_5673, \8417 );
nor \g452970/U$1 ( \33320 , \33318 , \33319 );
nand \g447827/U$1 ( \33321 , \33306 , \33314 , \33317 , \33320 );
and \g444791/U$2 ( \33322 , \33321 , \8369 );
and \g446253/U$2 ( \33323 , RIfe85d88_7867, \8356 );
and \g446253/U$3 ( \33324 , RIf15c998_5513, \8340 );
and \g449209/U$2 ( \33325 , RIfec0618_8309, \8371 );
and \g449209/U$3 ( \33326 , \8383 , RIf165d40_5618);
and \g449209/U$4 ( \33327 , RIf15deb0_5528, \8488 );
nor \g449209/U$1 ( \33328 , \33325 , \33326 , \33327 );
and \g454227/U$2 ( \33329 , \8313 , RIf163310_5588);
and \g454227/U$3 ( \33330 , RIf164288_5599, \8323 );
nor \g454227/U$1 ( \33331 , \33329 , \33330 );
not \g450223/U$3 ( \33332 , \33331 );
not \g450223/U$4 ( \33333 , \8376 );
and \g450223/U$2 ( \33334 , \33332 , \33333 );
and \g450223/U$5 ( \33335 , \8359 , RIf15fda0_5550);
nor \g450223/U$1 ( \33336 , \33334 , \33335 );
and \g452988/U$2 ( \33337 , \8404 , RIfe86760_7874);
and \g452988/U$3 ( \33338 , RIf166f88_5631, \8351 );
nor \g452988/U$1 ( \33339 , \33337 , \33338 );
and \g452991/U$2 ( \33340 , \8378 , RIf161c90_5572);
and \g452991/U$3 ( \33341 , RIfc52b08_5963, \8417 );
nor \g452991/U$1 ( \33342 , \33340 , \33341 );
nand \g447832/U$1 ( \33343 , \33328 , \33336 , \33339 , \33342 );
nor \g446253/U$1 ( \33344 , \33323 , \33324 , \33343 );
and \g452985/U$2 ( \33345 , \8335 , RIf159b30_5480);
and \g452985/U$3 ( \33346 , RIfe865f8_7873, \8531 );
nor \g452985/U$1 ( \33347 , \33345 , \33346 );
and \g452982/U$2 ( \33348 , \8319 , RIf15a3a0_5486);
and \g452982/U$3 ( \33349 , RIf15b480_5498, \8324 );
nor \g452982/U$1 ( \33350 , \33348 , \33349 );
and \g445329/U$2 ( \33351 , \33344 , \33347 , \33350 );
nor \g445329/U$1 ( \33352 , \33351 , \8422 );
nor \g444791/U$1 ( \33353 , \33322 , \33352 );
and \g447015/U$2 ( \33354 , \8707 , RIe207228_4371);
and \g447015/U$3 ( \33355 , RIe209f28_4403, \8709 );
nor \g447015/U$1 ( \33356 , \33354 , \33355 );
and \g447014/U$2 ( \33357 , \8712 , RIe20cc28_4435);
and \g447014/U$3 ( \33358 , RIf167c30_5640, \8714 );
nor \g447014/U$1 ( \33359 , \33357 , \33358 );
and \g447019/U$2 ( \33360 , \8717 , RIe20f928_4467);
and \g447019/U$3 ( \33361 , RIf168e78_5653, \8719 );
nor \g447019/U$1 ( \33362 , \33360 , \33361 );
nand \g444517/U$1 ( \33363 , \33353 , \33356 , \33359 , \33362 );
and \g453027/U$2 ( \33364 , \8414 , RIfec0a50_8312);
and \g453027/U$3 ( \33365 , RIfc819f8_6497, \8409 );
nor \g453027/U$1 ( \33366 , \33364 , \33365 );
and \g446262/U$2 ( \33367 , RIf14a248_5303, \8417 );
and \g446262/U$3 ( \33368 , RIfe86490_7872, \8404 );
and \g449223/U$2 ( \33369 , RIfe86058_7869, \8319 );
and \g449223/U$3 ( \33370 , \8326 , RIf146198_5257);
and \g449223/U$4 ( \33371 , RIf14b490_5316, \8383 );
nor \g449223/U$1 ( \33372 , \33369 , \33370 , \33371 );
and \g453042/U$2 ( \33373 , \8335 , RIfec08e8_8311);
and \g453042/U$3 ( \33374 , RIfcbb478_7153, \8340 );
nor \g453042/U$1 ( \33375 , \33373 , \33374 );
and \g454364/U$2 ( \33376 , \8313 , RIfe86328_7871);
and \g454364/U$3 ( \33377 , RIf147980_5274, \8323 );
nor \g454364/U$1 ( \33378 , \33376 , \33377 );
not \g450238/U$3 ( \33379 , \33378 );
not \g450238/U$4 ( \33380 , \8347 );
and \g450238/U$2 ( \33381 , \33379 , \33380 );
and \g450238/U$5 ( \33382 , \8351 , RIf14c6d8_5329);
nor \g450238/U$1 ( \33383 , \33381 , \33382 );
and \g453038/U$2 ( \33384 , \8356 , RIfec0780_8310);
and \g453038/U$3 ( \33385 , RIf148bc8_5287, \8359 );
nor \g453038/U$1 ( \33386 , \33384 , \33385 );
nand \g447839/U$1 ( \33387 , \33372 , \33375 , \33383 , \33386 );
nor \g446262/U$1 ( \33388 , \33367 , \33368 , \33387 );
and \g453031/U$2 ( \33389 , \8378 , RIfe861c0_7870);
and \g453031/U$3 ( \33390 , RIfe85ef0_7868, \8371 );
nor \g453031/U$1 ( \33391 , \33389 , \33390 );
nand \g445642/U$1 ( \33392 , \33366 , \33388 , \33391 );
and \g444902/U$2 ( \33393 , \33392 , \8482 );
and \g449216/U$2 ( \33394 , RIe1cc290_3700, \8531 );
and \g449216/U$3 ( \33395 , \8486 , RIe1cef90_3732);
and \g449216/U$4 ( \33396 , RIe1e8490_4020, \8383 );
nor \g449216/U$1 ( \33397 , \33394 , \33395 , \33396 );
and \g453015/U$2 ( \33398 , \8335 , RIe1be190_3540);
and \g453015/U$3 ( \33399 , RIe1c6890_3636, \8340 );
nor \g453015/U$1 ( \33400 , \33398 , \33399 );
and \g455173/U$2 ( \33401 , \8313 , RIe1c0e90_3572);
and \g455173/U$3 ( \33402 , RIe1c3b90_3604, \8323 );
nor \g455173/U$1 ( \33403 , \33401 , \33402 );
not \g455172/U$1 ( \33404 , \33403 );
and \g450231/U$2 ( \33405 , \33404 , \8316 );
and \g450231/U$3 ( \33406 , RIe1eb190_4052, \8351 );
nor \g450231/U$1 ( \33407 , \33405 , \33406 );
and \g453014/U$2 ( \33408 , \8356 , RIe1c9590_3668);
and \g453014/U$3 ( \33409 , RIe1d1c90_3764, \8359 );
nor \g453014/U$1 ( \33410 , \33408 , \33409 );
nand \g448212/U$1 ( \33411 , \33397 , \33400 , \33407 , \33410 );
and \g444902/U$3 ( \33412 , \8478 , \33411 );
nor \g444902/U$1 ( \33413 , \33393 , \33412 );
and \g447029/U$2 ( \33414 , \9480 , RIe1e2a90_3956);
and \g447029/U$3 ( \33415 , RIe1e5790_3988, \9482 );
nor \g447029/U$1 ( \33416 , \33414 , \33415 );
and \g447030/U$2 ( \33417 , \10539 , RIe1d7690_3828);
and \g447030/U$3 ( \33418 , RIe1da390_3860, \10541 );
nor \g447030/U$1 ( \33419 , \33417 , \33418 );
and \g447025/U$2 ( \33420 , \10534 , RIe1dd090_3892);
and \g447025/U$3 ( \33421 , RIe1dfd90_3924, \10536 );
nor \g447025/U$1 ( \33422 , \33420 , \33421 );
nand \g444638/U$1 ( \33423 , \33413 , \33416 , \33419 , \33422 );
and \g446233/U$2 ( \33424 , RIe183bd0_2876, \8356 );
and \g446233/U$3 ( \33425 , RIfc51758_5949, \8340 );
and \g449184/U$2 ( \33426 , RIf1454f0_5248, \8373 );
and \g449184/U$3 ( \33427 , \8383 , RIe19a3d0_3132);
and \g449184/U$4 ( \33428 , RIe1868d0_2908, \8488 );
nor \g449184/U$1 ( \33429 , \33426 , \33427 , \33428 );
and \g455042/U$2 ( \33430 , \8313 , RIe191cd0_3036);
and \g455042/U$3 ( \33431 , RIe1949d0_3068, \8323 );
nor \g455042/U$1 ( \33432 , \33430 , \33431 );
not \g450199/U$3 ( \33433 , \33432 );
not \g450199/U$4 ( \33434 , \8376 );
and \g450199/U$2 ( \33435 , \33433 , \33434 );
and \g450199/U$5 ( \33436 , \8359 , RIe1895d0_2940);
nor \g450199/U$1 ( \33437 , \33435 , \33436 );
and \g452906/U$2 ( \33438 , \8404 , RIe1976d0_3100);
and \g452906/U$3 ( \33439 , RIe19d0d0_3164, \8351 );
nor \g452906/U$1 ( \33440 , \33438 , \33439 );
and \g452908/U$2 ( \33441 , \8378 , RIe18efd0_3004);
and \g452908/U$3 ( \33442 , RIf144578_5237, \8417 );
nor \g452908/U$1 ( \33443 , \33441 , \33442 );
nand \g447816/U$1 ( \33444 , \33429 , \33437 , \33440 , \33443 );
nor \g446233/U$1 ( \33445 , \33424 , \33425 , \33444 );
and \g452899/U$2 ( \33446 , \8335 , RIe17b4d0_2780);
and \g452899/U$3 ( \33447 , RIf143498_5225, \8531 );
nor \g452899/U$1 ( \33448 , \33446 , \33447 );
and \g452895/U$2 ( \33449 , \8319 , RIe17e1d0_2812);
and \g452895/U$3 ( \33450 , RIe180ed0_2844, \8326 );
nor \g452895/U$1 ( \33451 , \33449 , \33450 );
and \g445315/U$2 ( \33452 , \33445 , \33448 , \33451 );
nor \g445315/U$1 ( \33453 , \33452 , \8589 );
and \g446241/U$2 ( \33454 , RIee39b20_5115, \8531 );
and \g446241/U$3 ( \33455 , RIf16d4c8_5703, \8335 );
and \g449192/U$2 ( \33456 , RIe176e80_2730, \8373 );
and \g449192/U$3 ( \33457 , \8383 , RIfc9ee40_6830);
and \g449192/U$4 ( \33458 , RIee3aed0_5129, \8488 );
nor \g449192/U$1 ( \33459 , \33456 , \33457 , \33458 );
and \g455175/U$2 ( \33460 , \8313 , RIfcc4280_7254);
and \g455175/U$3 ( \33461 , RIfce0cf0_7580, \8323 );
nor \g455175/U$1 ( \33462 , \33460 , \33461 );
not \g450208/U$3 ( \33463 , \33462 );
not \g450208/U$4 ( \33464 , \8376 );
and \g450208/U$2 ( \33465 , \33463 , \33464 );
and \g450208/U$5 ( \33466 , \8359 , RIee3bfb0_5141);
nor \g450208/U$1 ( \33467 , \33465 , \33466 );
and \g452934/U$2 ( \33468 , \8404 , RIe175800_2714);
and \g452934/U$3 ( \33469 , RIfc9b060_6786, \8351 );
nor \g452934/U$1 ( \33470 , \33468 , \33469 );
and \g452935/U$2 ( \33471 , \8378 , RIfcba7d0_7144);
and \g452935/U$3 ( \33472 , RIfcb70f8_7105, \8417 );
nor \g452935/U$1 ( \33473 , \33471 , \33472 );
nand \g447821/U$1 ( \33474 , \33459 , \33467 , \33470 , \33473 );
nor \g446241/U$1 ( \33475 , \33454 , \33455 , \33474 );
and \g452925/U$2 ( \33476 , \8356 , RIe173370_2688);
and \g452925/U$3 ( \33477 , RIf170060_5734, \8340 );
nor \g452925/U$1 ( \33478 , \33476 , \33477 );
and \g452923/U$2 ( \33479 , \8319 , RIf16dea0_5710);
and \g452923/U$3 ( \33480 , RIf16f3b8_5725, \8326 );
nor \g452923/U$1 ( \33481 , \33479 , \33480 );
and \g445316/U$2 ( \33482 , \33475 , \33478 , \33481 );
nor \g445316/U$1 ( \33483 , \33482 , \8558 );
or \g444405/U$1 ( \33484 , \33363 , \33423 , \33453 , \33483 );
and \g446223/U$2 ( \33485 , RIfc4ac78_5873, \8417 );
and \g446223/U$3 ( \33486 , RIe1f9f38_4221, \8404 );
and \g449170/U$2 ( \33487 , RIf150620_5374, \8531 );
and \g449170/U$3 ( \33488 , \8488 , RIfc899f0_6588);
and \g449170/U$4 ( \33489 , RIfc4ade0_5874, \8383 );
nor \g449170/U$1 ( \33490 , \33487 , \33488 , \33489 );
and \g452857/U$2 ( \33491 , \8335 , RIe1edbc0_4082);
and \g452857/U$3 ( \33492 , RIf14f6a8_5363, \8340 );
nor \g452857/U$1 ( \33493 , \33491 , \33492 );
and \g455056/U$2 ( \33494 , \8313 , RIf14dbf0_5344);
and \g455056/U$3 ( \33495 , RIf14ea00_5354, \8323 );
nor \g455056/U$1 ( \33496 , \33494 , \33495 );
not \g455055/U$1 ( \33497 , \33496 );
and \g450185/U$2 ( \33498 , \33497 , \8316 );
and \g450185/U$3 ( \33499 , RIfc83348_6515, \8351 );
nor \g450185/U$1 ( \33500 , \33498 , \33499 );
and \g452856/U$2 ( \33501 , \8356 , RIe1f2eb8_4141);
and \g452856/U$3 ( \33502 , RIf152ee8_5403, \8359 );
nor \g452856/U$1 ( \33503 , \33501 , \33502 );
nand \g448205/U$1 ( \33504 , \33490 , \33493 , \33500 , \33503 );
nor \g446223/U$1 ( \33505 , \33485 , \33486 , \33504 );
and \g452849/U$2 ( \33506 , \8378 , RIe1f5078_4165);
and \g452849/U$3 ( \33507 , RIfc89720_6586, \8373 );
nor \g452849/U$1 ( \33508 , \33506 , \33507 );
and \g452847/U$2 ( \33509 , \8414 , RIfc4ab10_5872);
and \g452847/U$3 ( \33510 , RIfc9f110_6832, \8409 );
nor \g452847/U$1 ( \33511 , \33509 , \33510 );
and \g445306/U$2 ( \33512 , \33505 , \33508 , \33511 );
nor \g445306/U$1 ( \33513 , \33512 , \8621 );
and \g446230/U$2 ( \33514 , RIe18c2d0_2972, \8417 );
and \g446230/U$3 ( \33515 , RIe19fdd0_3196, \8404 );
and \g449176/U$2 ( \33516 , RIe1ae308_3359, \8319 );
and \g449176/U$3 ( \33517 , \8326 , RIe1bb490_3508);
and \g449176/U$4 ( \33518 , RIe1a57d0_3260, \8383 );
nor \g449176/U$1 ( \33519 , \33516 , \33517 , \33518 );
and \g452885/U$2 ( \33520 , \8335 , RIe170940_2658);
and \g452885/U$3 ( \33521 , RIe1d4990_3796, \8340 );
nor \g452885/U$1 ( \33522 , \33520 , \33521 );
and \g455117/U$2 ( \33523 , \8313 , RIe1f7940_4194);
and \g455117/U$3 ( \33524 , RIe1fe588_4271, \8323 );
nor \g455117/U$1 ( \33525 , \33523 , \33524 );
not \g450193/U$3 ( \33526 , \33525 );
not \g450193/U$4 ( \33527 , \8347 );
and \g450193/U$2 ( \33528 , \33526 , \33527 );
and \g450193/U$5 ( \33529 , \8351 , RIe1a84d0_3292);
nor \g450193/U$1 ( \33530 , \33528 , \33529 );
and \g452883/U$2 ( \33531 , \8356 , RIe1f0488_4111);
and \g452883/U$3 ( \33532 , RIe204528_4339, \8359 );
nor \g452883/U$1 ( \33533 , \33531 , \33532 );
nand \g447812/U$1 ( \33534 , \33519 , \33522 , \33530 , \33533 );
nor \g446230/U$1 ( \33535 , \33514 , \33515 , \33534 );
and \g452877/U$2 ( \33536 , \8378 , RIe21ad28_4595);
and \g452877/U$3 ( \33537 , RIe1a2ad0_3228, \8373 );
nor \g452877/U$1 ( \33538 , \33536 , \33537 );
and \g452873/U$2 ( \33539 , \8412 , RIe226128_4723);
and \g452873/U$3 ( \33540 , RIe1787d0_2748, \8409 );
nor \g452873/U$1 ( \33541 , \33539 , \33540 );
and \g445313/U$2 ( \33542 , \33535 , \33538 , \33541 );
nor \g445313/U$1 ( \33543 , \33542 , \8651 );
or \g444192/U$1 ( \33544 , \33484 , \33513 , \33543 );
_DC \g5800/U$1 ( \33545 , \33544 , \8654 );
and \g453233/U$2 ( \33546 , \16361 , RIde7be90_194);
and \g453233/U$3 ( \33547 , RIdf37d98_2012, \16427 );
nor \g453233/U$1 ( \33548 , \33546 , \33547 );
and \g446303/U$2 ( \33549 , RIe1433a0_2142, \16432 );
and \g446303/U$3 ( \33550 , RIdf2c3f8_1880, \16371 );
and \g449273/U$2 ( \33551 , RIde95f48_321, \16485 );
and \g449273/U$3 ( \33552 , \16356 , RIdeb41a0_513);
and \g449273/U$4 ( \33553 , RIdee6e70_1091, \16398 );
nor \g449273/U$1 ( \33554 , \33551 , \33552 , \33553 );
and \g455299/U$2 ( \33555 , \16317 , RIdecd6a0_801);
and \g455299/U$3 ( \33556 , RIded03a0_833, \16325 );
nor \g455299/U$1 ( \33557 , \33555 , \33556 );
not \g450290/U$3 ( \33558 , \33557 );
not \g450290/U$4 ( \33559 , \16311 );
and \g450290/U$2 ( \33560 , \33558 , \33559 );
and \g450290/U$5 ( \33561 , \16339 , RIdf00370_1379);
nor \g450290/U$1 ( \33562 , \33560 , \33561 );
and \g453241/U$2 ( \33563 , \16377 , RIdec7ca0_737);
and \g453241/U$3 ( \33564 , RIdeca9a0_769, \16313 );
nor \g453241/U$1 ( \33565 , \33563 , \33564 );
and \g453242/U$2 ( \33566 , \16334 , RIe159ba0_2398);
and \g453242/U$3 ( \33567 , RIe16dda8_2627, \16380 );
nor \g453242/U$1 ( \33568 , \33566 , \33567 );
nand \g447406/U$1 ( \33569 , \33554 , \33562 , \33565 , \33568 );
nor \g446303/U$1 ( \33570 , \33549 , \33550 , \33569 );
and \g453231/U$2 ( \33571 , \16364 , RIdedbbd8_964);
and \g453231/U$3 ( \33572 , RIdf1cc78_1704, \16368 );
nor \g453231/U$1 ( \33573 , \33571 , \33572 );
nand \g445653/U$1 ( \33574 , \33548 , \33570 , \33573 );
and \g444895/U$2 ( \33575 , \33574 , \16752 );
and \g449268/U$2 ( \33576 , RIfcd43d8_7437, \16427 );
and \g449268/U$3 ( \33577 , \16448 , RIfcd7ee8_7479);
and \g449268/U$4 ( \33578 , RIdee2988_1042, \16344 );
nor \g449268/U$1 ( \33579 , \33576 , \33577 , \33578 );
and \g454576/U$2 ( \33580 , \16317 , RIded6fe8_910);
and \g454576/U$3 ( \33581 , RIded9478_936, \16325 );
nor \g454576/U$1 ( \33582 , \33580 , \33581 );
not \g454575/U$1 ( \33583 , \33582 );
and \g450284/U$2 ( \33584 , \33583 , \16336 );
and \g450284/U$3 ( \33585 , RIfec0078_8305, \16356 );
nor \g450284/U$1 ( \33586 , \33584 , \33585 );
and \g453219/U$2 ( \33587 , \16361 , RIfeab330_8264);
and \g453219/U$3 ( \33588 , RIded50f8_888, \16364 );
nor \g453219/U$1 ( \33589 , \33587 , \33588 );
and \g453217/U$2 ( \33590 , \16368 , RIfc9e5d0_6824);
and \g453217/U$3 ( \33591 , RIfc88eb0_6580, \16371 );
nor \g453217/U$1 ( \33592 , \33590 , \33591 );
nand \g448099/U$1 ( \33593 , \33579 , \33586 , \33589 , \33592 );
and \g444895/U$3 ( \33594 , \16477 , \33593 );
nor \g444895/U$1 ( \33595 , \33575 , \33594 );
and \g447067/U$2 ( \33596 , \18268 , RIfcb54d8_7085);
and \g447067/U$3 ( \33597 , RIfec0348_8307, \18270 );
nor \g447067/U$1 ( \33598 , \33596 , \33597 );
and \g447068/U$2 ( \33599 , \18273 , RIfc54e30_5988);
and \g447068/U$3 ( \33600 , RIee23cf8_4866, \18275 );
nor \g447068/U$1 ( \33601 , \33599 , \33600 );
and \g447071/U$2 ( \33602 , \18278 , RIdede770_995);
and \g447071/U$3 ( \33603 , RIfec01e0_8306, \18280 );
nor \g447071/U$1 ( \33604 , \33602 , \33603 );
nand \g444645/U$1 ( \33605 , \33595 , \33598 , \33601 , \33604 );
and \g449256/U$2 ( \33606 , RIdf08a70_1475, \16485 );
and \g449256/U$3 ( \33607 , \16356 , RIdf0b770_1507);
and \g449256/U$4 ( \33608 , RIdeef570_1187, \16398 );
nor \g449256/U$1 ( \33609 , \33606 , \33607 , \33608 );
and \g454655/U$2 ( \33610 , \16317 , RIdf13e70_1603);
and \g454655/U$3 ( \33611 , RIdf16b70_1635, \16325 );
nor \g454655/U$1 ( \33612 , \33610 , \33611 );
not \g450272/U$3 ( \33613 , \33612 );
not \g450272/U$4 ( \33614 , \16311 );
and \g450272/U$2 ( \33615 , \33613 , \33614 );
and \g450272/U$5 ( \33616 , \16341 , RIdef2270_1219);
nor \g450272/U$1 ( \33617 , \33615 , \33616 );
and \g453170/U$2 ( \33618 , \16377 , RIdf0e470_1539);
and \g453170/U$3 ( \33619 , RIdf11170_1571, \16313 );
nor \g453170/U$1 ( \33620 , \33618 , \33619 );
and \g453173/U$2 ( \33621 , \16334 , RIdf03070_1411);
and \g453173/U$3 ( \33622 , RIdf05d70_1443, \16380 );
nor \g453173/U$1 ( \33623 , \33621 , \33622 );
nand \g447399/U$1 ( \33624 , \33609 , \33617 , \33620 , \33623 );
and \g444718/U$2 ( \33625 , \33624 , \16750 );
and \g446295/U$2 ( \33626 , RIee29f68_4936, \16321 );
and \g446295/U$3 ( \33627 , RIee28bb8_4922, \16313 );
and \g449263/U$2 ( \33628 , RIee26b60_4899, \16427 );
and \g449263/U$3 ( \33629 , \16448 , RIee27100_4903);
and \g449263/U$4 ( \33630 , RIfe84e10_7856, \16344 );
nor \g449263/U$1 ( \33631 , \33628 , \33629 , \33630 );
and \g454624/U$2 ( \33632 , \16317 , RIdf1f540_1733);
and \g454624/U$3 ( \33633 , RIfc9e300_6822, \16325 );
nor \g454624/U$1 ( \33634 , \33632 , \33633 );
not \g454623/U$1 ( \33635 , \33634 );
and \g450278/U$2 ( \33636 , \33635 , \16336 );
and \g450278/U$3 ( \33637 , RIdf2a0d0_1855, \16356 );
nor \g450278/U$1 ( \33638 , \33636 , \33637 );
and \g453201/U$2 ( \33639 , \16361 , RIfe84b40_7854);
and \g453201/U$3 ( \33640 , RIee25eb8_4890, \16364 );
nor \g453201/U$1 ( \33641 , \33639 , \33640 );
and \g453198/U$2 ( \33642 , \16368 , RIee265c0_4895);
and \g453198/U$3 ( \33643 , RIfcd32f8_7425, \16371 );
nor \g453198/U$1 ( \33644 , \33642 , \33643 );
nand \g448098/U$1 ( \33645 , \33631 , \33638 , \33641 , \33644 );
nor \g446295/U$1 ( \33646 , \33626 , \33627 , \33645 );
and \g453190/U$2 ( \33647 , \16377 , RIee27970_4909);
and \g453190/U$3 ( \33648 , RIdf262f0_1811, \16380 );
nor \g453190/U$1 ( \33649 , \33647 , \33648 );
and \g453188/U$2 ( \33650 , \16334 , RIfe84ca8_7855);
and \g453188/U$3 ( \33651 , RIee2b8b8_4954, \16328 );
nor \g453188/U$1 ( \33652 , \33650 , \33651 );
and \g445360/U$2 ( \33653 , \33646 , \33649 , \33652 );
nor \g445360/U$1 ( \33654 , \33653 , \16480 );
nor \g444718/U$1 ( \33655 , \33625 , \33654 );
and \g447061/U$2 ( \33656 , \19208 , RIdee9b70_1123);
and \g447061/U$3 ( \33657 , RIdef7c70_1283, \19210 );
nor \g447061/U$1 ( \33658 , \33656 , \33657 );
and \g447062/U$2 ( \33659 , \19213 , RIdeec870_1155);
and \g447062/U$3 ( \33660 , RIdef4f70_1251, \19215 );
nor \g447062/U$1 ( \33661 , \33659 , \33660 );
and \g447060/U$2 ( \33662 , \19218 , RIdefa970_1315);
and \g447060/U$3 ( \33663 , RIdefd670_1347, \19220 );
nor \g447060/U$1 ( \33664 , \33662 , \33663 );
nand \g444644/U$1 ( \33665 , \33655 , \33658 , \33661 , \33664 );
and \g446278/U$2 ( \33666 , RIee1cb10_4785, \16328 );
and \g446278/U$3 ( \33667 , RIfe84f78_7857, \16334 );
and \g449242/U$2 ( \33668 , RIfe853b0_7860, \16427 );
and \g449242/U$3 ( \33669 , \16448 , RIee1a3b0_4757);
and \g449242/U$4 ( \33670 , RIde8d230_278, \16485 );
nor \g449242/U$1 ( \33671 , \33668 , \33669 , \33670 );
and \g454542/U$2 ( \33672 , \16317 , RIe16b378_2597);
and \g454542/U$3 ( \33673 , RIee39148_5108, \16325 );
nor \g454542/U$1 ( \33674 , \33672 , \33673 );
not \g454541/U$1 ( \33675 , \33674 );
and \g450257/U$2 ( \33676 , \33675 , \16336 );
and \g450257/U$3 ( \33677 , RIfe850e0_7858, \16356 );
nor \g450257/U$1 ( \33678 , \33676 , \33677 );
and \g453120/U$2 ( \33679 , \16361 , RIe167b38_2557);
and \g453120/U$3 ( \33680 , RIee38608_5100, \16364 );
nor \g453120/U$1 ( \33681 , \33679 , \33680 );
and \g453119/U$2 ( \33682 , \16368 , RIfe85248_7859);
and \g453119/U$3 ( \33683 , RIee199d8_4750, \16371 );
nor \g453119/U$1 ( \33684 , \33682 , \33683 );
nand \g448097/U$1 ( \33685 , \33671 , \33678 , \33681 , \33684 );
nor \g446278/U$1 ( \33686 , \33666 , \33667 , \33685 );
and \g453111/U$2 ( \33687 , \16377 , RIfec04b0_8308);
and \g453111/U$3 ( \33688 , RIfea9cb0_8248, \16380 );
nor \g453111/U$1 ( \33689 , \33687 , \33688 );
and \g453110/U$2 ( \33690 , \16313 , RIee1b1c0_4767);
and \g453110/U$3 ( \33691 , RIee1ba30_4773, \16321 );
nor \g453110/U$1 ( \33692 , \33690 , \33691 );
and \g445349/U$2 ( \33693 , \33686 , \33689 , \33692 );
nor \g445349/U$1 ( \33694 , \33693 , \16649 );
and \g446285/U$2 ( \33695 , RIfe85c20_7866, \16432 );
and \g446285/U$3 ( \33696 , RIee34dc8_5060, \16371 );
and \g449251/U$2 ( \33697 , RIe15c8a0_2430, \16485 );
and \g449251/U$3 ( \33698 , \16356 , RIee36010_5073);
and \g449251/U$4 ( \33699 , RIe14baa0_2238, \16337 );
nor \g449251/U$1 ( \33700 , \33697 , \33698 , \33699 );
and \g455263/U$2 ( \33701 , \16317 , RIe1622a0_2494);
and \g455263/U$3 ( \33702 , RIe164fa0_2526, \16325 );
nor \g455263/U$1 ( \33703 , \33701 , \33702 );
not \g450265/U$3 ( \33704 , \33703 );
not \g450265/U$4 ( \33705 , \16311 );
and \g450265/U$2 ( \33706 , \33704 , \33705 );
and \g450265/U$5 ( \33707 , \16341 , RIfc861b0_6548);
nor \g450265/U$1 ( \33708 , \33706 , \33707 );
and \g453147/U$2 ( \33709 , \16377 , RIe15f5a0_2462);
and \g453147/U$3 ( \33710 , RIfe85950_7864, \16313 );
nor \g453147/U$1 ( \33711 , \33709 , \33710 );
and \g453150/U$2 ( \33712 , \16334 , RIe1541a0_2334);
and \g453150/U$3 ( \33713 , RIe156ea0_2366, \16380 );
nor \g453150/U$1 ( \33714 , \33712 , \33713 );
nand \g447398/U$1 ( \33715 , \33700 , \33708 , \33711 , \33714 );
nor \g446285/U$1 ( \33716 , \33695 , \33696 , \33715 );
and \g453137/U$2 ( \33717 , \16364 , RIe148da0_2206);
and \g453137/U$3 ( \33718 , RIe14e7a0_2270, \16368 );
nor \g453137/U$1 ( \33719 , \33717 , \33718 );
and \g453140/U$2 ( \33720 , \16361 , RIe1460a0_2174);
and \g453140/U$3 ( \33721 , RIe1514a0_2302, \16427 );
nor \g453140/U$1 ( \33722 , \33720 , \33721 );
and \g445353/U$2 ( \33723 , \33716 , \33719 , \33722 );
nor \g445353/U$1 ( \33724 , \33723 , \16389 );
or \g444345/U$1 ( \33725 , \33605 , \33665 , \33694 , \33724 );
and \g446267/U$2 ( \33726 , RIdeb14a0_481, \16427 );
and \g446267/U$3 ( \33727 , RIdeae7a0_449, \16368 );
and \g449229/U$2 ( \33728 , RIdec22a0_673, \16321 );
and \g449229/U$3 ( \33729 , \16328 , RIdec4fa0_705);
and \g449229/U$4 ( \33730 , RIdea9a48_417, \16398 );
nor \g449229/U$1 ( \33731 , \33728 , \33729 , \33730 );
and \g455201/U$2 ( \33732 , \16317 , RIdebc8a0_609);
and \g455201/U$3 ( \33733 , RIee1f270_4813, \16325 );
nor \g455201/U$1 ( \33734 , \33732 , \33733 );
not \g450243/U$3 ( \33735 , \33734 );
not \g450243/U$4 ( \33736 , \16330 );
and \g450243/U$2 ( \33737 , \33735 , \33736 );
and \g450243/U$5 ( \33738 , \16339 , RIee1d920_4795);
nor \g450243/U$1 ( \33739 , \33737 , \33738 );
and \g453067/U$2 ( \33740 , \16377 , RIdebf5a0_641);
and \g453067/U$3 ( \33741 , RIee1fdb0_4821, \16313 );
nor \g453067/U$1 ( \33742 , \33740 , \33741 );
and \g453069/U$2 ( \33743 , \16334 , RIdeb6ea0_545);
and \g453069/U$3 ( \33744 , RIdeb9ba0_577, \16380 );
nor \g453069/U$1 ( \33745 , \33743 , \33744 );
nand \g447396/U$1 ( \33746 , \33731 , \33739 , \33742 , \33745 );
nor \g446267/U$1 ( \33747 , \33726 , \33727 , \33746 );
and \g453057/U$2 ( \33748 , \16361 , RIde9c848_353);
and \g453057/U$3 ( \33749 , RIee1ecd0_4809, \16432 );
nor \g453057/U$1 ( \33750 , \33748 , \33749 );
and \g453054/U$2 ( \33751 , \16364 , RIdea3148_385);
and \g453054/U$3 ( \33752 , RIee1e730_4805, \16371 );
nor \g453054/U$1 ( \33753 , \33751 , \33752 );
and \g445342/U$2 ( \33754 , \33747 , \33750 , \33753 );
nor \g445342/U$1 ( \33755 , \33754 , \16618 );
and \g446273/U$2 ( \33756 , RIee343f0_5053, \16328 );
and \g446273/U$3 ( \33757 , RIfe85680_7862, \16377 );
and \g449235/U$2 ( \33758 , RIee2f698_4998, \16427 );
and \g449235/U$3 ( \33759 , \16448 , RIfc9d4f0_6812);
and \g449235/U$4 ( \33760 , RIdf3eb48_2090, \16485 );
nor \g449235/U$1 ( \33761 , \33758 , \33759 , \33760 );
and \g454487/U$2 ( \33762 , \16317 , RIdf32ed8_1956);
and \g454487/U$3 ( \33763 , RIdf35368_1982, \16325 );
nor \g454487/U$1 ( \33764 , \33762 , \33763 );
not \g454486/U$1 ( \33765 , \33764 );
and \g450250/U$2 ( \33766 , \33765 , \16336 );
and \g450250/U$3 ( \33767 , RIe140c40_2114, \16356 );
nor \g450250/U$1 ( \33768 , \33766 , \33767 );
and \g453095/U$2 ( \33769 , \16361 , RIfe85ab8_7865);
and \g453095/U$3 ( \33770 , RIdf30e80_1933, \16364 );
nor \g453095/U$1 ( \33771 , \33769 , \33770 );
and \g453093/U$2 ( \33772 , \16368 , RIee2d4d8_4974);
and \g453093/U$3 ( \33773 , RIfc52298_5957, \16371 );
nor \g453093/U$1 ( \33774 , \33772 , \33773 );
nand \g448096/U$1 ( \33775 , \33761 , \33768 , \33771 , \33774 );
nor \g446273/U$1 ( \33776 , \33756 , \33757 , \33775 );
and \g453084/U$2 ( \33777 , \16334 , RIdf3a660_2041);
and \g453084/U$3 ( \33778 , RIfe857e8_7863, \16313 );
nor \g453084/U$1 ( \33779 , \33777 , \33778 );
and \g453082/U$2 ( \33780 , \16380 , RIdf3c820_2065);
and \g453082/U$3 ( \33781 , RIfe85518_7861, \16319 );
nor \g453082/U$1 ( \33782 , \33780 , \33781 );
and \g445348/U$2 ( \33783 , \33776 , \33779 , \33782 );
nor \g445348/U$1 ( \33784 , \33783 , \16393 );
or \g444281/U$1 ( \33785 , \33725 , \33755 , \33784 );
_DC \g5885/U$1 ( \33786 , \33785 , \16652 );
and \g449381/U$2 ( \33787 , RIee3e2d8_5166, \8414 );
and \g449381/U$3 ( \33788 , \8409 , RIf13ee48_5175);
and \g449381/U$4 ( \33789 , RIf140a68_5195, \8383 );
nor \g449381/U$1 ( \33790 , \33787 , \33788 , \33789 );
and \g453633/U$2 ( \33791 , \8356 , RIfe838f8_7841);
and \g453633/U$3 ( \33792 , RIee3c118_5142, \8359 );
nor \g453633/U$1 ( \33793 , \33791 , \33792 );
and \g455353/U$2 ( \33794 , \8313 , RIee39c88_5116);
and \g455353/U$3 ( \33795 , RIee3b038_5130, \8323 );
nor \g455353/U$1 ( \33796 , \33794 , \33795 );
not \g450400/U$3 ( \33797 , \33796 );
not \g450400/U$4 ( \33798 , \8347 );
and \g450400/U$2 ( \33799 , \33797 , \33798 );
and \g450400/U$5 ( \33800 , \8351 , RIf1420e8_5211);
nor \g450400/U$1 ( \33801 , \33799 , \33800 );
and \g453631/U$2 ( \33802 , \8378 , RIee3d1f8_5154);
and \g453631/U$3 ( \33803 , RIf13faf0_5184, \8417 );
nor \g453631/U$1 ( \33804 , \33802 , \33803 );
nand \g447935/U$1 ( \33805 , \33790 , \33793 , \33801 , \33804 );
and \g444689/U$2 ( \33806 , \33805 , \9700 );
and \g446394/U$2 ( \33807 , RIe194b38_3069, \8409 );
and \g446394/U$3 ( \33808 , RIe18f138_3005, \8378 );
and \g449386/U$2 ( \33809 , RIf145658_5249, \8373 );
and \g449386/U$3 ( \33810 , \8383 , RIe19a538_3133);
and \g449386/U$4 ( \33811 , RIe186a38_2909, \8488 );
nor \g449386/U$1 ( \33812 , \33809 , \33810 , \33811 );
and \g453660/U$2 ( \33813 , \8335 , RIe17b638_2781);
and \g453660/U$3 ( \33814 , RIf142c28_5219, \8340 );
nor \g453660/U$1 ( \33815 , \33813 , \33814 );
and \g453658/U$2 ( \33816 , \8404 , RIe197838_3101);
and \g453658/U$3 ( \33817 , RIe19d238_3165, \8351 );
nor \g453658/U$1 ( \33818 , \33816 , \33817 );
and \g455279/U$2 ( \33819 , \8313 , RIe17e338_2813);
and \g455279/U$3 ( \33820 , RIe181038_2845, \8323 );
nor \g455279/U$1 ( \33821 , \33819 , \33820 );
not \g455278/U$1 ( \33822 , \33821 );
and \g450407/U$2 ( \33823 , \33822 , \8316 );
and \g450407/U$3 ( \33824 , RIe189738_2941, \8359 );
nor \g450407/U$1 ( \33825 , \33823 , \33824 );
nand \g448234/U$1 ( \33826 , \33812 , \33815 , \33818 , \33825 );
nor \g446394/U$1 ( \33827 , \33807 , \33808 , \33826 );
and \g453652/U$2 ( \33828 , \8356 , RIe183d38_2877);
and \g453652/U$3 ( \33829 , RIf1446e0_5238, \8417 );
nor \g453652/U$1 ( \33830 , \33828 , \33829 );
and \g453650/U$2 ( \33831 , \8523 , RIf143600_5226);
and \g453650/U$3 ( \33832 , RIe191e38_3037, \8414 );
nor \g453650/U$1 ( \33833 , \33831 , \33832 );
and \g445426/U$2 ( \33834 , \33827 , \33830 , \33833 );
nor \g445426/U$1 ( \33835 , \33834 , \8589 );
nor \g444689/U$1 ( \33836 , \33806 , \33835 );
and \g447142/U$2 ( \33837 , \10034 , RIfc5ab00_6054);
and \g447142/U$3 ( \33838 , RIf1701c8_5735, \10036 );
nor \g447142/U$1 ( \33839 , \33837 , \33838 );
and \g447138/U$2 ( \33840 , \10039 , RIfebff10_8304);
and \g447138/U$3 ( \33841 , RIf1401f8_5189, \10041 );
nor \g447138/U$1 ( \33842 , \33840 , \33841 );
and \g447143/U$2 ( \33843 , \10044 , RIfcb0e88_7035);
and \g447143/U$3 ( \33844 , RIf16e008_5711, \10046 );
nor \g447143/U$1 ( \33845 , \33843 , \33844 );
nand \g444536/U$1 ( \33846 , \33836 , \33839 , \33842 , \33845 );
and \g453690/U$2 ( \33847 , \8319 , RIe1c0ff8_3573);
and \g453690/U$3 ( \33848 , RIe1c3cf8_3605, \8326 );
nor \g453690/U$1 ( \33849 , \33847 , \33848 );
and \g446401/U$2 ( \33850 , RIe1c69f8_3637, \8340 );
and \g446401/U$3 ( \33851 , RIe1e2bf8_3957, \8404 );
and \g449398/U$2 ( \33852 , RIe1da4f8_3861, \8414 );
and \g449398/U$3 ( \33853 , \8409 , RIe1dd1f8_3893);
and \g449398/U$4 ( \33854 , RIe1e85f8_4021, \8383 );
nor \g449398/U$1 ( \33855 , \33852 , \33853 , \33854 );
and \g453700/U$2 ( \33856 , \8356 , RIe1c96f8_3669);
and \g453700/U$3 ( \33857 , RIe1d1df8_3765, \8359 );
nor \g453700/U$1 ( \33858 , \33856 , \33857 );
and \g455364/U$2 ( \33859 , \8313 , RIe1cc3f8_3701);
and \g455364/U$3 ( \33860 , RIe1cf0f8_3733, \8323 );
nor \g455364/U$1 ( \33861 , \33859 , \33860 );
not \g450419/U$3 ( \33862 , \33861 );
not \g450419/U$4 ( \33863 , \8347 );
and \g450419/U$2 ( \33864 , \33862 , \33863 );
and \g450419/U$5 ( \33865 , \8351 , RIe1eb2f8_4053);
nor \g450419/U$1 ( \33866 , \33864 , \33865 );
and \g453697/U$2 ( \33867 , \8378 , RIe1d77f8_3829);
and \g453697/U$3 ( \33868 , RIe1dfef8_3925, \8417 );
nor \g453697/U$1 ( \33869 , \33867 , \33868 );
nand \g447944/U$1 ( \33870 , \33855 , \33858 , \33866 , \33869 );
nor \g446401/U$1 ( \33871 , \33850 , \33851 , \33870 );
and \g453688/U$2 ( \33872 , \8335 , RIe1be2f8_3541);
and \g453688/U$3 ( \33873 , RIe1e58f8_3989, \8373 );
nor \g453688/U$1 ( \33874 , \33872 , \33873 );
nand \g445681/U$1 ( \33875 , \33849 , \33871 , \33874 );
and \g444804/U$2 ( \33876 , \33875 , \8478 );
and \g449393/U$2 ( \33877 , RIfe83a60_7842, \8373 );
and \g449393/U$3 ( \33878 , \8383 , RIf14b5f8_5317);
and \g449393/U$4 ( \33879 , RIf147ae8_5275, \8486 );
nor \g449393/U$1 ( \33880 , \33877 , \33878 , \33879 );
and \g453678/U$2 ( \33881 , \8335 , RIfe83790_7840);
and \g453678/U$3 ( \33882 , RIf146fa8_5267, \8340 );
nor \g453678/U$1 ( \33883 , \33881 , \33882 );
and \g453673/U$2 ( \33884 , \8404 , RIfe849d8_7853);
and \g453673/U$3 ( \33885 , RIf14c840_5330, \8351 );
nor \g453673/U$1 ( \33886 , \33884 , \33885 );
and \g455163/U$2 ( \33887 , \8313 , RIfe845a0_7850);
and \g455163/U$3 ( \33888 , RIf146300_5258, \8323 );
nor \g455163/U$1 ( \33889 , \33887 , \33888 );
not \g455162/U$1 ( \33890 , \33889 );
and \g450414/U$2 ( \33891 , \33890 , \8316 );
and \g450414/U$3 ( \33892 , RIf148d30_5288, \8359 );
nor \g450414/U$1 ( \33893 , \33891 , \33892 );
nand \g448235/U$1 ( \33894 , \33880 , \33883 , \33886 , \33893 );
and \g444804/U$3 ( \33895 , \8482 , \33894 );
nor \g444804/U$1 ( \33896 , \33876 , \33895 );
and \g447152/U$2 ( \33897 , \8964 , RIf149b40_5298);
and \g447152/U$3 ( \33898 , RIfc74168_6343, \8966 );
nor \g447152/U$1 ( \33899 , \33897 , \33898 );
and \g447153/U$2 ( \33900 , \8521 , RIe1b0900_3386);
and \g447153/U$3 ( \33901 , RIfe84870_7852, \8525 );
nor \g447153/U$1 ( \33902 , \33900 , \33901 );
and \g447154/U$2 ( \33903 , \8974 , RIfe84708_7851);
and \g447154/U$3 ( \33904 , RIfe83bc8_7843, \8976 );
nor \g447154/U$1 ( \33905 , \33903 , \33904 );
nand \g444537/U$1 ( \33906 , \33896 , \33899 , \33902 , \33905 );
and \g446379/U$2 ( \33907 , RIf16bce0_5686, \8373 );
and \g446379/U$3 ( \33908 , RIe20a090_4404, \8319 );
and \g449369/U$2 ( \33909 , RIf168fe0_5654, \8523 );
and \g449369/U$3 ( \33910 , \8488 , RIe212790_4500);
and \g449369/U$4 ( \33911 , RIe223590_4692, \8383 );
nor \g449369/U$1 ( \33912 , \33909 , \33910 , \33911 );
and \g453591/U$2 ( \33913 , \8356 , RIe20fa90_4468);
and \g453591/U$3 ( \33914 , RIf16a228_5667, \8359 );
nor \g453591/U$1 ( \33915 , \33913 , \33914 );
and \g455160/U$2 ( \33916 , \8313 , RIe218190_4564);
and \g455160/U$3 ( \33917 , RIe21db90_4628, \8323 );
nor \g455160/U$1 ( \33918 , \33916 , \33917 );
not \g450389/U$3 ( \33919 , \33918 );
not \g450389/U$4 ( \33920 , \8376 );
and \g450389/U$2 ( \33921 , \33919 , \33920 );
and \g450389/U$5 ( \33922 , \8351 , RIf16caf0_5696);
nor \g450389/U$1 ( \33923 , \33921 , \33922 );
and \g453588/U$2 ( \33924 , \8378 , RIe215490_4532);
and \g453588/U$3 ( \33925 , RIf16ac00_5674, \8417 );
nor \g453588/U$1 ( \33926 , \33924 , \33925 );
nand \g447925/U$1 ( \33927 , \33912 , \33915 , \33923 , \33926 );
nor \g446379/U$1 ( \33928 , \33907 , \33908 , \33927 );
and \g453582/U$2 ( \33929 , \8335 , RIe207390_4372);
and \g453582/U$3 ( \33930 , RIf167d98_5641, \8340 );
nor \g453582/U$1 ( \33931 , \33929 , \33930 );
and \g453579/U$2 ( \33932 , \8326 , RIe20cd90_4436);
and \g453579/U$3 ( \33933 , RIe220890_4660, \8404 );
nor \g453579/U$1 ( \33934 , \33932 , \33933 );
and \g445414/U$2 ( \33935 , \33928 , \33931 , \33934 );
nor \g445414/U$1 ( \33936 , \33935 , \8368 );
and \g446384/U$2 ( \33937 , RIe202200_4314, \8371 );
and \g446384/U$3 ( \33938 , RIf15a508_5487, \8317 );
and \g449374/U$2 ( \33939 , RIfe83d30_7844, \8523 );
and \g449374/U$3 ( \33940 , \8488 , RIf15e018_5529);
and \g449374/U$4 ( \33941 , RIf165ea8_5619, \8383 );
nor \g449374/U$1 ( \33942 , \33939 , \33940 , \33941 );
and \g453615/U$2 ( \33943 , \8356 , RIfe84000_7846);
and \g453615/U$3 ( \33944 , RIf15ff08_5551, \8359 );
nor \g453615/U$1 ( \33945 , \33943 , \33944 );
and \g455348/U$2 ( \33946 , \8313 , RIfce8310_7664);
and \g455348/U$3 ( \33947 , RIf1643f0_5600, \8323 );
nor \g455348/U$1 ( \33948 , \33946 , \33947 );
not \g450393/U$3 ( \33949 , \33948 );
not \g450393/U$4 ( \33950 , \8376 );
and \g450393/U$2 ( \33951 , \33949 , \33950 );
and \g450393/U$5 ( \33952 , \8351 , RIf1670f0_5632);
nor \g450393/U$1 ( \33953 , \33951 , \33952 );
and \g453614/U$2 ( \33954 , \8378 , RIf161df8_5573);
and \g453614/U$3 ( \33955 , RIf164f30_5608, \8417 );
nor \g453614/U$1 ( \33956 , \33954 , \33955 );
nand \g447929/U$1 ( \33957 , \33942 , \33945 , \33953 , \33956 );
nor \g446384/U$1 ( \33958 , \33937 , \33938 , \33957 );
and \g453606/U$2 ( \33959 , \8335 , RIfc887a8_6575);
and \g453606/U$3 ( \33960 , RIf15cb00_5514, \8340 );
nor \g453606/U$1 ( \33961 , \33959 , \33960 );
and \g453604/U$2 ( \33962 , \8326 , RIf15b5e8_5499);
and \g453604/U$3 ( \33963 , RIfe83e98_7845, \8404 );
nor \g453604/U$1 ( \33964 , \33962 , \33963 );
and \g445418/U$2 ( \33965 , \33958 , \33961 , \33964 );
nor \g445418/U$1 ( \33966 , \33965 , \8422 );
or \g444374/U$1 ( \33967 , \33846 , \33906 , \33936 , \33966 );
and \g446369/U$2 ( \33968 , RIfc51fc8_5955, \8409 );
and \g446369/U$3 ( \33969 , RIe1f51e0_4166, \8378 );
and \g449355/U$2 ( \33970 , RIf156cc8_5447, \8373 );
and \g449355/U$3 ( \33971 , \8383 , RIf157970_5456);
and \g449355/U$4 ( \33972 , RIf1519d0_5388, \8488 );
nor \g449355/U$1 ( \33973 , \33970 , \33971 , \33972 );
and \g453541/U$2 ( \33974 , \8335 , RIfe84168_7847);
and \g453541/U$3 ( \33975 , RIf14f810_5364, \8340 );
nor \g453541/U$1 ( \33976 , \33974 , \33975 );
and \g453539/U$2 ( \33977 , \8404 , RIfe84438_7849);
and \g453539/U$3 ( \33978 , RIf158d20_5470, \8351 );
nor \g453539/U$1 ( \33979 , \33977 , \33978 );
and \g454697/U$2 ( \33980 , \8313 , RIf14dd58_5345);
and \g454697/U$3 ( \33981 , RIf14eb68_5355, \8323 );
nor \g454697/U$1 ( \33982 , \33980 , \33981 );
not \g454696/U$1 ( \33983 , \33982 );
and \g450375/U$2 ( \33984 , \33983 , \8316 );
and \g450375/U$3 ( \33985 , RIf153050_5404, \8359 );
nor \g450375/U$1 ( \33986 , \33984 , \33985 );
nand \g448228/U$1 ( \33987 , \33973 , \33976 , \33979 , \33986 );
nor \g446369/U$1 ( \33988 , \33968 , \33969 , \33987 );
and \g453532/U$2 ( \33989 , \8356 , RIfe842d0_7848);
and \g453532/U$3 ( \33990 , RIf156020_5438, \8417 );
nor \g453532/U$1 ( \33991 , \33989 , \33990 );
and \g453529/U$2 ( \33992 , \8523 , RIf150788_5375);
and \g453529/U$3 ( \33993 , RIf154568_5419, \8414 );
nor \g453529/U$1 ( \33994 , \33992 , \33993 );
and \g445406/U$2 ( \33995 , \33988 , \33991 , \33994 );
nor \g445406/U$1 ( \33996 , \33995 , \8621 );
and \g446372/U$2 ( \33997 , RIe226290_4724, \8414 );
and \g446372/U$3 ( \33998 , RIe18c438_2973, \8417 );
and \g449362/U$2 ( \33999 , RIe1a2c38_3229, \8373 );
and \g449362/U$3 ( \34000 , \8383 , RIe1a5938_3261);
and \g449362/U$4 ( \34001 , RIe1fe6f0_4272, \8488 );
nor \g449362/U$1 ( \34002 , \33999 , \34000 , \34001 );
and \g453569/U$2 ( \34003 , \8335 , RIe170aa8_2659);
and \g453569/U$3 ( \34004 , RIe1d4af8_3797, \8340 );
nor \g453569/U$1 ( \34005 , \34003 , \34004 );
and \g453564/U$2 ( \34006 , \8404 , RIe19ff38_3197);
and \g453564/U$3 ( \34007 , RIe1a8638_3293, \8351 );
nor \g453564/U$1 ( \34008 , \34006 , \34007 );
and \g454587/U$2 ( \34009 , \8313 , RIe1ae470_3360);
and \g454587/U$3 ( \34010 , RIe1bb5f8_3509, \8323 );
nor \g454587/U$1 ( \34011 , \34009 , \34010 );
not \g454586/U$1 ( \34012 , \34011 );
and \g450383/U$2 ( \34013 , \34012 , \8316 );
and \g450383/U$3 ( \34014 , RIe204690_4340, \8359 );
nor \g450383/U$1 ( \34015 , \34013 , \34014 );
nand \g448231/U$1 ( \34016 , \34002 , \34005 , \34008 , \34015 );
nor \g446372/U$1 ( \34017 , \33997 , \33998 , \34016 );
and \g453554/U$2 ( \34018 , \8378 , RIe21ae90_4596);
and \g453554/U$3 ( \34019 , RIe1f7aa8_4195, \8531 );
nor \g453554/U$1 ( \34020 , \34018 , \34019 );
and \g453558/U$2 ( \34021 , \8356 , RIe1f05f0_4112);
and \g453558/U$3 ( \34022 , RIe178938_2749, \8409 );
nor \g453558/U$1 ( \34023 , \34021 , \34022 );
and \g445408/U$2 ( \34024 , \34017 , \34020 , \34023 );
nor \g445408/U$1 ( \34025 , \34024 , \8651 );
or \g444193/U$1 ( \34026 , \33967 , \33996 , \34025 );
_DC \g5909/U$1 ( \34027 , \34026 , \8654 );
and \g451322/U$2 ( \34028 , \16364 , RIe169a28_2579);
and \g451322/U$3 ( \34029 , RIfc82100_6502, \16371 );
nor \g451322/U$1 ( \34030 , \34028 , \34029 );
and \g445869/U$2 ( \34031 , RIfc52f40_5966, \16427 );
and \g445869/U$3 ( \34032 , RIfca7108_6923, \16368 );
and \g448714/U$2 ( \34033 , RIfe7f9b0_7796, \16485 );
and \g448714/U$3 ( \34034 , \16356 , RIde90d40_296);
and \g448714/U$4 ( \34035 , RIe16b648_2599, \16398 );
nor \g448714/U$1 ( \34036 , \34033 , \34034 , \34035 );
and \g455252/U$2 ( \34037 , \16317 , RIfcce438_7369);
and \g455252/U$3 ( \34038 , RIfcdc3d0_7528, \16325 );
nor \g455252/U$1 ( \34039 , \34037 , \34038 );
not \g449743/U$3 ( \34040 , \34039 );
not \g449743/U$4 ( \34041 , \16311 );
and \g449743/U$2 ( \34042 , \34040 , \34041 );
and \g449743/U$5 ( \34043 , \16341 , RIfe7fb18_7797);
nor \g449743/U$1 ( \34044 , \34042 , \34043 );
and \g451331/U$2 ( \34045 , \16377 , RIfc75680_6358);
and \g451331/U$3 ( \34046 , RIfcb0a50_7032, \16313 );
nor \g451331/U$1 ( \34047 , \34045 , \34046 );
and \g451336/U$2 ( \34048 , \16334 , RIde85580_240);
and \g451336/U$3 ( \34049 , RIde89720_260, \16380 );
nor \g451336/U$1 ( \34050 , \34048 , \34049 );
nand \g447278/U$1 ( \34051 , \34036 , \34044 , \34047 , \34050 );
nor \g445869/U$1 ( \34052 , \34031 , \34032 , \34051 );
and \g451323/U$2 ( \34053 , \16361 , RIe167ca0_2558);
and \g451323/U$3 ( \34054 , RIde81728_221, \16448 );
nor \g451323/U$1 ( \34055 , \34053 , \34054 );
nand \g445544/U$1 ( \34056 , \34030 , \34052 , \34055 );
and \g444704/U$2 ( \34057 , \34056 , \17998 );
and \g448706/U$2 ( \34058 , RIdeaa0d8_419, \16337 );
and \g448706/U$3 ( \34059 , \16341 , RIfcaf808_7019);
and \g448706/U$4 ( \34060 , RIdebcb70_611, \16485 );
nor \g448706/U$1 ( \34061 , \34058 , \34059 , \34060 );
and \g454992/U$2 ( \34062 , \16317 , RIdeb1770_483);
and \g454992/U$3 ( \34063 , RIfe7fc80_7798, \16325 );
nor \g454992/U$1 ( \34064 , \34062 , \34063 );
not \g449737/U$3 ( \34065 , \34064 );
not \g449737/U$4 ( \34066 , \16351 );
and \g449737/U$2 ( \34067 , \34065 , \34066 );
and \g449737/U$5 ( \34068 , \16356 , RIfe7f848_7795);
nor \g449737/U$1 ( \34069 , \34067 , \34068 );
and \g451313/U$2 ( \34070 , \16361 , RIde9ced8_355);
and \g451313/U$3 ( \34071 , RIdea37d8_387, \16364 );
nor \g451313/U$1 ( \34072 , \34070 , \34071 );
and \g454077/U$2 ( \34073 , \16368 , RIdeaea70_451);
and \g454077/U$3 ( \34074 , RIfca5d58_6909, \16371 );
nor \g454077/U$1 ( \34075 , \34073 , \34074 );
nand \g447572/U$1 ( \34076 , \34061 , \34069 , \34072 , \34075 );
and \g444704/U$3 ( \34077 , \17938 , \34076 );
nor \g444704/U$1 ( \34078 , \34057 , \34077 );
and \g446650/U$2 ( \34079 , \18960 , RIdeb7170_547);
and \g446650/U$3 ( \34080 , RIdeb9e70_579, \18962 );
nor \g446650/U$1 ( \34081 , \34079 , \34080 );
and \g446649/U$2 ( \34082 , \18965 , RIdec2570_675);
and \g446649/U$3 ( \34083 , RIdec5270_707, \18967 );
nor \g446649/U$1 ( \34084 , \34082 , \34083 );
and \g446653/U$2 ( \34085 , \18776 , RIdebf870_643);
and \g446653/U$3 ( \34086 , RIee1ff18_4822, \18778 );
nor \g446653/U$1 ( \34087 , \34085 , \34086 );
nand \g444466/U$1 ( \34088 , \34078 , \34081 , \34084 , \34087 );
and \g451371/U$2 ( \34089 , \16377 , RIee23320_4859);
and \g451371/U$3 ( \34090 , RIfe80220_7802, \16380 );
nor \g451371/U$1 ( \34091 , \34089 , \34090 );
and \g445880/U$2 ( \34092 , RIee24838_4874, \16321 );
and \g445880/U$3 ( \34093 , RIfc4cb68_5895, \16313 );
and \g448729/U$2 ( \34094 , RIee223a8_4848, \16427 );
and \g448729/U$3 ( \34095 , \16432 , RIfc98900_6758);
and \g448729/U$4 ( \34096 , RIdee2c58_1044, \16485 );
nor \g448729/U$1 ( \34097 , \34094 , \34095 , \34096 );
and \g454592/U$2 ( \34098 , \16317 , RIfe804f0_7804);
and \g454592/U$3 ( \34099 , RIded9748_938, \16325 );
nor \g454592/U$1 ( \34100 , \34098 , \34099 );
not \g454591/U$1 ( \34101 , \34100 );
and \g449760/U$2 ( \34102 , \34101 , \16336 );
and \g449760/U$3 ( \34103 , RIfe80388_7803, \16356 );
nor \g449760/U$1 ( \34104 , \34102 , \34103 );
and \g451381/U$2 ( \34105 , \16361 , RIded2c68_862);
and \g451381/U$3 ( \34106 , RIded53c8_890, \16364 );
nor \g451381/U$1 ( \34107 , \34105 , \34106 );
and \g451376/U$2 ( \34108 , \16368 , RIee212c8_4836);
and \g451376/U$3 ( \34109 , RIfcc8600_7302, \16371 );
nor \g451376/U$1 ( \34110 , \34108 , \34109 );
nand \g448037/U$1 ( \34111 , \34097 , \34104 , \34107 , \34110 );
nor \g445880/U$1 ( \34112 , \34092 , \34093 , \34111 );
and \g452258/U$2 ( \34113 , \16334 , RIdedea40_997);
and \g452258/U$3 ( \34114 , RIfcb7800_7110, \16326 );
nor \g452258/U$1 ( \34115 , \34113 , \34114 );
nand \g445547/U$1 ( \34116 , \34091 , \34112 , \34115 );
and \g444909/U$2 ( \34117 , \34116 , \16477 );
and \g448723/U$2 ( \34118 , RIee2a0d0_4937, \16321 );
and \g448723/U$3 ( \34119 , \16328 , RIee2bb88_4956);
and \g448723/U$4 ( \34120 , RIdf1f810_1735, \16398 );
nor \g448723/U$1 ( \34121 , \34118 , \34119 , \34120 );
and \g454273/U$2 ( \34122 , \16317 , RIdf27f10_1831);
and \g454273/U$3 ( \34123 , RIdf2a238_1856, \16325 );
nor \g454273/U$1 ( \34124 , \34122 , \34123 );
not \g449752/U$3 ( \34125 , \34124 );
not \g449752/U$4 ( \34126 , \16330 );
and \g449752/U$2 ( \34127 , \34125 , \34126 );
and \g449752/U$5 ( \34128 , \16341 , RIdf21700_1757);
nor \g449752/U$1 ( \34129 , \34127 , \34128 );
and \g451351/U$2 ( \34130 , \16377 , RIfe7f578_7793);
and \g451351/U$3 ( \34131 , RIee28d20_4923, \16313 );
nor \g451351/U$1 ( \34132 , \34130 , \34131 );
and \g451355/U$2 ( \34133 , \16334 , RIdf246d0_1791);
and \g451355/U$3 ( \34134 , RIfe7f6e0_7794, \16380 );
nor \g451355/U$1 ( \34135 , \34133 , \34134 );
nand \g447283/U$1 ( \34136 , \34121 , \34129 , \34132 , \34135 );
and \g444909/U$3 ( \34137 , \16481 , \34136 );
nor \g444909/U$1 ( \34138 , \34117 , \34137 );
and \g446665/U$2 ( \34139 , \17274 , RIfc63638_6153);
and \g446665/U$3 ( \34140 , RIfcce9d8_7373, \17276 );
nor \g446665/U$1 ( \34141 , \34139 , \34140 );
and \g446666/U$2 ( \34142 , \17279 , RIfc62990_6144);
and \g446666/U$3 ( \34143 , RIdf22c18_1772, \17281 );
nor \g446666/U$1 ( \34144 , \34142 , \34143 );
and \g446669/U$2 ( \34145 , \17284 , RIdf19168_1662);
and \g446669/U$3 ( \34146 , RIfeaa958_8257, \17286 );
nor \g446669/U$1 ( \34147 , \34145 , \34146 );
nand \g444574/U$1 ( \34148 , \34138 , \34141 , \34144 , \34147 );
and \g445854/U$2 ( \34149 , RIee331a8_5040, \16321 );
and \g445854/U$3 ( \34150 , RIee320c8_5028, \16313 );
and \g448691/U$2 ( \34151 , RIee2f800_4999, \16427 );
and \g448691/U$3 ( \34152 , \16448 , RIfcc8330_7300);
and \g448691/U$4 ( \34153 , RIfe7ff50_7800, \16485 );
nor \g448691/U$1 ( \34154 , \34151 , \34152 , \34153 );
and \g455102/U$2 ( \34155 , \16317 , RIdf331a8_1958);
and \g455102/U$3 ( \34156 , RIdf35638_1984, \16325 );
nor \g455102/U$1 ( \34157 , \34155 , \34156 );
not \g455101/U$1 ( \34158 , \34157 );
and \g449720/U$2 ( \34159 , \34158 , \16336 );
and \g449720/U$3 ( \34160 , RIfe800b8_7801, \16356 );
nor \g449720/U$1 ( \34161 , \34159 , \34160 );
and \g451266/U$2 ( \34162 , \16361 , RIdf2ef90_1911);
and \g451266/U$3 ( \34163 , RIdf31150_1935, \16364 );
nor \g451266/U$1 ( \34164 , \34162 , \34163 );
and \g451262/U$2 ( \34165 , \16368 , RIee2d640_4975);
and \g451262/U$3 ( \34166 , RIfca0d30_6852, \16371 );
nor \g451262/U$1 ( \34167 , \34165 , \34166 );
nand \g448028/U$1 ( \34168 , \34154 , \34161 , \34164 , \34167 );
nor \g445854/U$1 ( \34169 , \34149 , \34150 , \34168 );
and \g451257/U$2 ( \34170 , \16377 , RIee31150_5017);
and \g451257/U$3 ( \34171 , RIdf3caf0_2067, \16380 );
nor \g451257/U$1 ( \34172 , \34170 , \34171 );
and \g451256/U$2 ( \34173 , \16334 , RIfe7fde8_7799);
and \g451256/U$3 ( \34174 , RIee34558_5054, \16328 );
nor \g451256/U$1 ( \34175 , \34173 , \34174 );
and \g445041/U$2 ( \34176 , \34169 , \34172 , \34175 );
nor \g445041/U$1 ( \34177 , \34176 , \16393 );
and \g445860/U$2 ( \34178 , RIe162570_2496, \16321 );
and \g445860/U$3 ( \34179 , RIee37258_5086, \16313 );
and \g448698/U$2 ( \34180 , RIe14bd70_2240, \16398 );
and \g448698/U$3 ( \34181 , \16339 , RIfce1290_7584);
and \g448698/U$4 ( \34182 , RIe15cb70_2432, \16485 );
nor \g448698/U$1 ( \34183 , \34180 , \34181 , \34182 );
and \g454229/U$2 ( \34184 , \16317 , RIe151770_2304);
and \g454229/U$3 ( \34185 , RIfc86fc0_6558, \16325 );
nor \g454229/U$1 ( \34186 , \34184 , \34185 );
not \g449728/U$3 ( \34187 , \34186 );
not \g449728/U$4 ( \34188 , \16351 );
and \g449728/U$2 ( \34189 , \34187 , \34188 );
and \g449728/U$5 ( \34190 , \16354 , RIee36178_5074);
nor \g449728/U$1 ( \34191 , \34189 , \34190 );
and \g450811/U$2 ( \34192 , \16361 , RIe146370_2176);
and \g450811/U$3 ( \34193 , RIe149070_2208, \16364 );
nor \g450811/U$1 ( \34194 , \34192 , \34193 );
and \g451287/U$2 ( \34195 , \16368 , RIe14ea70_2272);
and \g451287/U$3 ( \34196 , RIfc4eff8_5921, \16371 );
nor \g451287/U$1 ( \34197 , \34195 , \34196 );
nand \g447568/U$1 ( \34198 , \34183 , \34191 , \34194 , \34197 );
nor \g445860/U$1 ( \34199 , \34178 , \34179 , \34198 );
and \g451281/U$2 ( \34200 , \16377 , RIe15f870_2464);
and \g451281/U$3 ( \34201 , RIe157170_2368, \16380 );
nor \g451281/U$1 ( \34202 , \34200 , \34201 );
and \g450952/U$2 ( \34203 , \16334 , RIe154470_2336);
and \g450952/U$3 ( \34204 , RIe165270_2528, \16328 );
nor \g450952/U$1 ( \34205 , \34203 , \34204 );
and \g445043/U$2 ( \34206 , \34199 , \34202 , \34205 );
nor \g445043/U$1 ( \34207 , \34206 , \16389 );
or \g444340/U$1 ( \34208 , \34088 , \34148 , \34177 , \34207 );
and \g445842/U$2 ( \34209 , RIdefac40_1317, \16427 );
and \g445842/U$3 ( \34210 , RIdef5240_1253, \16368 );
and \g448675/U$2 ( \34211 , RIdf14140_1605, \16321 );
and \g448675/U$3 ( \34212 , \16328 , RIdf16e40_1637);
and \g448675/U$4 ( \34213 , RIdeef840_1189, \16398 );
nor \g448675/U$1 ( \34214 , \34211 , \34212 , \34213 );
and \g454418/U$2 ( \34215 , \16317 , RIdf08d40_1477);
and \g454418/U$3 ( \34216 , RIdf0ba40_1509, \16325 );
nor \g454418/U$1 ( \34217 , \34215 , \34216 );
not \g449706/U$3 ( \34218 , \34217 );
not \g449706/U$4 ( \34219 , \16330 );
and \g449706/U$2 ( \34220 , \34218 , \34219 );
and \g449706/U$5 ( \34221 , \16339 , RIdef2540_1221);
nor \g449706/U$1 ( \34222 , \34220 , \34221 );
and \g451209/U$2 ( \34223 , \16377 , RIdf0e740_1541);
and \g451209/U$3 ( \34224 , RIdf11440_1573, \16313 );
nor \g451209/U$1 ( \34225 , \34223 , \34224 );
and \g451212/U$2 ( \34226 , \16334 , RIdf03340_1413);
and \g451212/U$3 ( \34227 , RIdf06040_1445, \16380 );
nor \g451212/U$1 ( \34228 , \34226 , \34227 );
nand \g447268/U$1 ( \34229 , \34214 , \34222 , \34225 , \34228 );
nor \g445842/U$1 ( \34230 , \34209 , \34210 , \34229 );
and \g451206/U$2 ( \34231 , \16361 , RIdee9e40_1125);
and \g451206/U$3 ( \34232 , RIdefd940_1349, \16448 );
nor \g451206/U$1 ( \34233 , \34231 , \34232 );
and \g451201/U$2 ( \34234 , \16364 , RIdeecb40_1157);
and \g451201/U$3 ( \34235 , RIdef7f40_1285, \16371 );
nor \g451201/U$1 ( \34236 , \34234 , \34235 );
and \g445033/U$2 ( \34237 , \34230 , \34233 , \34236 );
nor \g445033/U$1 ( \34238 , \34237 , \16555 );
and \g445846/U$2 ( \34239 , RIdf38068_2014, \16427 );
and \g445846/U$3 ( \34240 , RIdf1cf48_1706, \16368 );
and \g448684/U$2 ( \34241 , RIdecd970_803, \16319 );
and \g448684/U$3 ( \34242 , \16328 , RIded0670_835);
and \g448684/U$4 ( \34243 , RIdee7140_1093, \16398 );
nor \g448684/U$1 ( \34244 , \34241 , \34242 , \34243 );
and \g454506/U$2 ( \34245 , \16317 , RIde965d8_323);
and \g454506/U$3 ( \34246 , RIdeb4470_515, \16325 );
nor \g454506/U$1 ( \34247 , \34245 , \34246 );
not \g449712/U$3 ( \34248 , \34247 );
not \g449712/U$4 ( \34249 , \16330 );
and \g449712/U$2 ( \34250 , \34248 , \34249 );
and \g449712/U$5 ( \34251 , \16339 , RIdf00640_1381);
nor \g449712/U$1 ( \34252 , \34250 , \34251 );
and \g451236/U$2 ( \34253 , \16377 , RIdec7f70_739);
and \g451236/U$3 ( \34254 , RIdecac70_771, \16313 );
nor \g451236/U$1 ( \34255 , \34253 , \34254 );
and \g451243/U$2 ( \34256 , \16334 , RIe159e70_2400);
and \g451243/U$3 ( \34257 , RIe16e078_2629, \16380 );
nor \g451243/U$1 ( \34258 , \34256 , \34257 );
nand \g447270/U$1 ( \34259 , \34244 , \34252 , \34255 , \34258 );
nor \g445846/U$1 ( \34260 , \34239 , \34240 , \34259 );
and \g451227/U$2 ( \34261 , \16361 , RIde7c520_196);
and \g451227/U$3 ( \34262 , RIe143670_2144, \16448 );
nor \g451227/U$1 ( \34263 , \34261 , \34262 );
and \g451226/U$2 ( \34264 , \16364 , RIdedbea8_966);
and \g451226/U$3 ( \34265 , RIdf2c6c8_1882, \16371 );
nor \g451226/U$1 ( \34266 , \34264 , \34265 );
and \g445038/U$2 ( \34267 , \34260 , \34263 , \34266 );
nor \g445038/U$1 ( \34268 , \34267 , \16586 );
or \g444222/U$1 ( \34269 , \34208 , \34238 , \34268 );
_DC \g598e/U$1 ( \34270 , \34269 , \16652 );
and \g448763/U$2 ( \34271 , RIe176fe8_2731, \8373 );
and \g448763/U$3 ( \34272 , \8383 , RIf140d38_5197);
and \g448763/U$4 ( \34273 , RIee3b1a0_5131, \8488 );
nor \g448763/U$1 ( \34274 , \34271 , \34272 , \34273 );
and \g455304/U$2 ( \34275 , \8313 , RIee3e440_5167);
and \g455304/U$3 ( \34276 , RIf13f118_5177, \8323 );
nor \g455304/U$1 ( \34277 , \34275 , \34276 );
not \g449791/U$3 ( \34278 , \34277 );
not \g449791/U$4 ( \34279 , \8376 );
and \g449791/U$2 ( \34280 , \34278 , \34279 );
and \g449791/U$5 ( \34281 , \8359 , RIee3c280_5143);
nor \g449791/U$1 ( \34282 , \34280 , \34281 );
and \g451484/U$2 ( \34283 , \8404 , RIe175ad0_2716);
and \g451484/U$3 ( \34284 , RIfe7f410_7792, \8351 );
nor \g451484/U$1 ( \34285 , \34283 , \34284 );
and \g451486/U$2 ( \34286 , \8378 , RIee3d360_5155);
and \g451486/U$3 ( \34287 , RIfe7f2a8_7791, \8417 );
nor \g451486/U$1 ( \34288 , \34286 , \34287 );
nand \g447602/U$1 ( \34289 , \34274 , \34282 , \34285 , \34288 );
and \g444680/U$2 ( \34290 , \34289 , \9700 );
and \g445913/U$2 ( \34291 , RIf143768_5227, \8531 );
and \g445913/U$3 ( \34292 , RIe17e608_2815, \8319 );
and \g448768/U$2 ( \34293 , RIfe7ee70_7788, \8373 );
and \g448768/U$3 ( \34294 , \8383 , RIe19a808_3135);
and \g448768/U$4 ( \34295 , RIe186d08_2911, \8488 );
nor \g448768/U$1 ( \34296 , \34293 , \34294 , \34295 );
and \g454518/U$2 ( \34297 , \8313 , RIe192108_3039);
and \g454518/U$3 ( \34298 , RIe194e08_3071, \8323 );
nor \g454518/U$1 ( \34299 , \34297 , \34298 );
not \g449797/U$3 ( \34300 , \34299 );
not \g449797/U$4 ( \34301 , \8376 );
and \g449797/U$2 ( \34302 , \34300 , \34301 );
and \g449797/U$5 ( \34303 , \8359 , RIe189a08_2943);
nor \g449797/U$1 ( \34304 , \34302 , \34303 );
and \g451509/U$2 ( \34305 , \8404 , RIe197b08_3103);
and \g451509/U$3 ( \34306 , RIe19d508_3167, \8351 );
nor \g451509/U$1 ( \34307 , \34305 , \34306 );
and \g451512/U$2 ( \34308 , \8378 , RIe18f408_3007);
and \g451512/U$3 ( \34309 , RIfe7efd8_7789, \8417 );
nor \g451512/U$1 ( \34310 , \34308 , \34309 );
nand \g447605/U$1 ( \34311 , \34296 , \34304 , \34307 , \34310 );
nor \g445913/U$1 ( \34312 , \34291 , \34292 , \34311 );
and \g451502/U$2 ( \34313 , \8335 , RIe17b908_2783);
and \g451502/U$3 ( \34314 , RIfc4bbf0_5884, \8340 );
nor \g451502/U$1 ( \34315 , \34313 , \34314 );
and \g451499/U$2 ( \34316 , \8326 , RIe181308_2847);
and \g451499/U$3 ( \34317 , RIe184008_2879, \8356 );
nor \g451499/U$1 ( \34318 , \34316 , \34317 );
and \g445085/U$2 ( \34319 , \34312 , \34315 , \34318 );
nor \g445085/U$1 ( \34320 , \34319 , \8589 );
nor \g444680/U$1 ( \34321 , \34290 , \34320 );
and \g446697/U$2 ( \34322 , \10044 , RIf16d630_5704);
and \g446697/U$3 ( \34323 , RIf16e2d8_5713, \10046 );
nor \g446697/U$1 ( \34324 , \34322 , \34323 );
and \g446696/U$2 ( \34325 , \10034 , RIf16f520_5726);
and \g446696/U$3 ( \34326 , RIf170330_5736, \10036 );
nor \g446696/U$1 ( \34327 , \34325 , \34326 );
and \g446699/U$2 ( \34328 , \12264 , RIe173640_2690);
and \g446699/U$3 ( \34329 , RIfe7f140_7790, \12266 );
nor \g446699/U$1 ( \34330 , \34328 , \34329 );
nand \g444473/U$1 ( \34331 , \34321 , \34324 , \34327 , \34330 );
and \g451549/U$2 ( \34332 , \8404 , RIfe7e600_7782);
and \g451549/U$3 ( \34333 , RIfca1f78_6865, \8409 );
nor \g451549/U$1 ( \34334 , \34332 , \34333 );
and \g445924/U$2 ( \34335 , RIfe7ed08_7787, \8373 );
and \g445924/U$3 ( \34336 , RIfe7e498_7781, \8378 );
and \g448781/U$2 ( \34337 , RIe1ac418_3337, \8317 );
and \g448781/U$3 ( \34338 , \8326 , RIf1465d0_5260);
and \g448781/U$4 ( \34339 , RIf14b760_5318, \8383 );
nor \g448781/U$1 ( \34340 , \34337 , \34338 , \34339 );
and \g451556/U$2 ( \34341 , \8335 , RIe1aac30_3320);
and \g451556/U$3 ( \34342 , RIf147278_5269, \8340 );
nor \g451556/U$1 ( \34343 , \34341 , \34342 );
and \g454581/U$2 ( \34344 , \8313 , RIfe7e330_7780);
and \g454581/U$3 ( \34345 , RIf147c50_5276, \8323 );
nor \g454581/U$1 ( \34346 , \34344 , \34345 );
not \g449808/U$3 ( \34347 , \34346 );
not \g449808/U$4 ( \34348 , \8347 );
and \g449808/U$2 ( \34349 , \34347 , \34348 );
and \g449808/U$5 ( \34350 , \8351 , RIf14c9a8_5331);
nor \g449808/U$1 ( \34351 , \34349 , \34350 );
and \g451555/U$2 ( \34352 , \8356 , RIe1b0a68_3387);
and \g451555/U$3 ( \34353 , RIf148e98_5289, \8359 );
nor \g451555/U$1 ( \34354 , \34352 , \34353 );
nand \g447613/U$1 ( \34355 , \34340 , \34343 , \34351 , \34354 );
nor \g445924/U$1 ( \34356 , \34335 , \34336 , \34355 );
and \g451546/U$2 ( \34357 , \8414 , RIfe7eba0_7786);
and \g451546/U$3 ( \34358 , RIf14a518_5305, \8417 );
nor \g451546/U$1 ( \34359 , \34357 , \34358 );
nand \g445558/U$1 ( \34360 , \34334 , \34356 , \34359 );
and \g444900/U$2 ( \34361 , \34360 , \8482 );
and \g448775/U$2 ( \34362 , RIe1cc6c8_3703, \8531 );
and \g448775/U$3 ( \34363 , \8488 , RIe1cf3c8_3735);
and \g448775/U$4 ( \34364 , RIe1e88c8_4023, \8383 );
nor \g448775/U$1 ( \34365 , \34362 , \34363 , \34364 );
and \g451533/U$2 ( \34366 , \8335 , RIe1be5c8_3543);
and \g451533/U$3 ( \34367 , RIe1c6cc8_3639, \8340 );
nor \g451533/U$1 ( \34368 , \34366 , \34367 );
and \g454412/U$2 ( \34369 , \8313 , RIe1c12c8_3575);
and \g454412/U$3 ( \34370 , RIe1c3fc8_3607, \8323 );
nor \g454412/U$1 ( \34371 , \34369 , \34370 );
not \g454411/U$1 ( \34372 , \34371 );
and \g449802/U$2 ( \34373 , \34372 , \8316 );
and \g449802/U$3 ( \34374 , RIe1eb5c8_4055, \8351 );
nor \g449802/U$1 ( \34375 , \34373 , \34374 );
and \g451530/U$2 ( \34376 , \8356 , RIe1c99c8_3671);
and \g451530/U$3 ( \34377 , RIe1d20c8_3767, \8359 );
nor \g451530/U$1 ( \34378 , \34376 , \34377 );
nand \g448163/U$1 ( \34379 , \34365 , \34368 , \34375 , \34378 );
and \g444900/U$3 ( \34380 , \8478 , \34379 );
nor \g444900/U$1 ( \34381 , \34361 , \34380 );
and \g446707/U$2 ( \34382 , \9480 , RIe1e2ec8_3959);
and \g446707/U$3 ( \34383 , RIe1e5bc8_3991, \9482 );
nor \g446707/U$1 ( \34384 , \34382 , \34383 );
and \g446708/U$2 ( \34385 , \10539 , RIe1d7ac8_3831);
and \g446708/U$3 ( \34386 , RIe1da7c8_3863, \10541 );
nor \g446708/U$1 ( \34387 , \34385 , \34386 );
and \g446706/U$2 ( \34388 , \10534 , RIe1dd4c8_3895);
and \g446706/U$3 ( \34389 , RIe1e01c8_3927, \10536 );
nor \g446706/U$1 ( \34390 , \34388 , \34389 );
nand \g444581/U$1 ( \34391 , \34381 , \34384 , \34387 , \34390 );
and \g445899/U$2 ( \34392 , RIe202368_4315, \8373 );
and \g445899/U$3 ( \34393 , RIf161f60_5574, \8378 );
and \g448751/U$2 ( \34394 , RIe1fcc38_4253, \8531 );
and \g448751/U$3 ( \34395 , \8486 , RIf15e180_5530);
and \g448751/U$4 ( \34396 , RIfc4e4b8_5913, \8383 );
nor \g448751/U$1 ( \34397 , \34394 , \34395 , \34396 );
and \g451454/U$2 ( \34398 , \8335 , RIf159c98_5481);
and \g451454/U$3 ( \34399 , RIf15cc68_5515, \8340 );
nor \g451454/U$1 ( \34400 , \34398 , \34399 );
and \g454579/U$2 ( \34401 , \8313 , RIf15a670_5488);
and \g454579/U$3 ( \34402 , RIf15b750_5500, \8323 );
nor \g454579/U$1 ( \34403 , \34401 , \34402 );
not \g454578/U$1 ( \34404 , \34403 );
and \g449780/U$2 ( \34405 , \34404 , \8316 );
and \g449780/U$3 ( \34406 , RIfc86750_6552, \8351 );
nor \g449780/U$1 ( \34407 , \34405 , \34406 );
and \g451451/U$2 ( \34408 , \8356 , RIe1fb9f0_4240);
and \g451451/U$3 ( \34409 , RIf160070_5552, \8359 );
nor \g451451/U$1 ( \34410 , \34408 , \34409 );
nand \g448161/U$1 ( \34411 , \34397 , \34400 , \34407 , \34410 );
nor \g445899/U$1 ( \34412 , \34392 , \34393 , \34411 );
and \g451445/U$2 ( \34413 , \8404 , RIe200a18_4297);
and \g451445/U$3 ( \34414 , RIf164558_5601, \8409 );
nor \g451445/U$1 ( \34415 , \34413 , \34414 );
and \g451443/U$2 ( \34416 , \8414 , RIf163478_5589);
and \g451443/U$3 ( \34417 , RIf165200_5610, \8417 );
nor \g451443/U$1 ( \34418 , \34416 , \34417 );
and \g445073/U$2 ( \34419 , \34412 , \34415 , \34418 );
nor \g445073/U$1 ( \34420 , \34419 , \8422 );
and \g445905/U$2 ( \34421 , RIfc4ddb0_5908, \8531 );
and \g445905/U$3 ( \34422 , RIe20a360_4406, \8319 );
and \g448758/U$2 ( \34423 , RIfc9c410_6800, \8373 );
and \g448758/U$3 ( \34424 , \8383 , RIe223860_4694);
and \g448758/U$4 ( \34425 , RIe212a60_4502, \8486 );
nor \g448758/U$1 ( \34426 , \34423 , \34424 , \34425 );
and \g454382/U$2 ( \34427 , \8313 , RIe218460_4566);
and \g454382/U$3 ( \34428 , RIe21de60_4630, \8323 );
nor \g454382/U$1 ( \34429 , \34427 , \34428 );
not \g449785/U$3 ( \34430 , \34429 );
not \g449785/U$4 ( \34431 , \8376 );
and \g449785/U$2 ( \34432 , \34430 , \34431 );
and \g449785/U$5 ( \34433 , \8359 , RIfc9cc80_6806);
nor \g449785/U$1 ( \34434 , \34432 , \34433 );
and \g453830/U$2 ( \34435 , \8404 , RIe220b60_4662);
and \g453830/U$3 ( \34436 , RIfe7ea38_7785, \8351 );
nor \g453830/U$1 ( \34437 , \34435 , \34436 );
and \g451468/U$2 ( \34438 , \8378 , RIe215760_4534);
and \g451468/U$3 ( \34439 , RIfcb8340_7118, \8417 );
nor \g451468/U$1 ( \34440 , \34438 , \34439 );
nand \g447597/U$1 ( \34441 , \34426 , \34434 , \34437 , \34440 );
nor \g445905/U$1 ( \34442 , \34421 , \34422 , \34441 );
and \g451467/U$2 ( \34443 , \8335 , RIe207660_4374);
and \g451467/U$3 ( \34444 , RIfc873f8_6561, \8340 );
nor \g451467/U$1 ( \34445 , \34443 , \34444 );
and \g451463/U$2 ( \34446 , \8326 , RIe20d060_4438);
and \g451463/U$3 ( \34447 , RIe20fd60_4470, \8356 );
nor \g451463/U$1 ( \34448 , \34446 , \34447 );
and \g445078/U$2 ( \34449 , \34442 , \34445 , \34448 );
nor \g445078/U$1 ( \34450 , \34449 , \8368 );
or \g444363/U$1 ( \34451 , \34331 , \34391 , \34420 , \34450 );
and \g445887/U$2 ( \34452 , RIf150a58_5377, \8531 );
and \g445887/U$3 ( \34453 , RIf14dec0_5346, \8319 );
and \g448736/U$2 ( \34454 , RIf154838_5421, \8414 );
and \g448736/U$3 ( \34455 , \8409 , RIf1557b0_5432);
and \g448736/U$4 ( \34456 , RIfc52400_5958, \8488 );
nor \g448736/U$1 ( \34457 , \34454 , \34455 , \34456 );
and \g454439/U$2 ( \34458 , \8313 , RIf156e30_5448);
and \g454439/U$3 ( \34459 , RIf157ad8_5457, \8323 );
nor \g454439/U$1 ( \34460 , \34458 , \34459 );
not \g449766/U$3 ( \34461 , \34460 );
not \g449766/U$4 ( \34462 , \8328 );
and \g449766/U$2 ( \34463 , \34461 , \34462 );
and \g449766/U$5 ( \34464 , \8359 , RIf1531b8_5405);
nor \g449766/U$1 ( \34465 , \34463 , \34464 );
and \g451397/U$2 ( \34466 , \8404 , RIfe7e768_7783);
and \g451397/U$3 ( \34467 , RIf158e88_5471, \8351 );
nor \g451397/U$1 ( \34468 , \34466 , \34467 );
and \g451402/U$2 ( \34469 , \8378 , RIfe7e8d0_7784);
and \g451402/U$3 ( \34470 , RIf1562f0_5440, \8417 );
nor \g451402/U$1 ( \34471 , \34469 , \34470 );
nand \g447582/U$1 ( \34472 , \34457 , \34465 , \34468 , \34471 );
nor \g445887/U$1 ( \34473 , \34452 , \34453 , \34472 );
and \g451395/U$2 ( \34474 , \8335 , RIe1ede90_4084);
and \g451395/U$3 ( \34475 , RIf14f978_5365, \8340 );
nor \g451395/U$1 ( \34476 , \34474 , \34475 );
and \g451656/U$2 ( \34477 , \8326 , RIf14ecd0_5356);
and \g451656/U$3 ( \34478 , RIe1f3188_4143, \8356 );
nor \g451656/U$1 ( \34479 , \34477 , \34478 );
and \g445065/U$2 ( \34480 , \34473 , \34476 , \34479 );
nor \g445065/U$1 ( \34481 , \34480 , \8621 );
and \g445893/U$2 ( \34482 , RIe18c708_2975, \8417 );
and \g445893/U$3 ( \34483 , RIe1a0208_3199, \8404 );
and \g448743/U$2 ( \34484 , RIe1ae740_3362, \8319 );
and \g448743/U$3 ( \34485 , \8326 , RIe1bb8c8_3511);
and \g448743/U$4 ( \34486 , RIe1a5c08_3263, \8383 );
nor \g448743/U$1 ( \34487 , \34484 , \34485 , \34486 );
and \g451427/U$2 ( \34488 , \8335 , RIe170d78_2661);
and \g451427/U$3 ( \34489 , RIe1d4dc8_3799, \8340 );
nor \g451427/U$1 ( \34490 , \34488 , \34489 );
and \g454642/U$2 ( \34491 , \8313 , RIe1f7d78_4197);
and \g454642/U$3 ( \34492 , RIe1fe9c0_4274, \8323 );
nor \g454642/U$1 ( \34493 , \34491 , \34492 );
not \g449772/U$3 ( \34494 , \34493 );
not \g449772/U$4 ( \34495 , \8347 );
and \g449772/U$2 ( \34496 , \34494 , \34495 );
and \g449772/U$5 ( \34497 , \8351 , RIe1a8908_3295);
nor \g449772/U$1 ( \34498 , \34496 , \34497 );
and \g451425/U$2 ( \34499 , \8356 , RIe1f08c0_4114);
and \g451425/U$3 ( \34500 , RIe204960_4342, \8359 );
nor \g451425/U$1 ( \34501 , \34499 , \34500 );
nand \g447588/U$1 ( \34502 , \34487 , \34490 , \34498 , \34501 );
nor \g445893/U$1 ( \34503 , \34482 , \34483 , \34502 );
and \g451419/U$2 ( \34504 , \8378 , RIe21b160_4598);
and \g451419/U$3 ( \34505 , RIe1a2f08_3231, \8373 );
nor \g451419/U$1 ( \34506 , \34504 , \34505 );
and \g451039/U$2 ( \34507 , \8412 , RIe226560_4726);
and \g451039/U$3 ( \34508 , RIe178c08_2751, \8409 );
nor \g451039/U$1 ( \34509 , \34507 , \34508 );
and \g445068/U$2 ( \34510 , \34503 , \34506 , \34509 );
nor \g445068/U$1 ( \34511 , \34510 , \8651 );
or \g444185/U$1 ( \34512 , \34451 , \34481 , \34511 );
_DC \g5a12/U$1 ( \34513 , \34512 , \8654 );
and \g451669/U$2 ( \34514 , \16313 , RIee32230_5029);
and \g451669/U$3 ( \34515 , RIfe7d688_7771, \16321 );
nor \g451669/U$1 ( \34516 , \34514 , \34515 );
and \g445953/U$2 ( \34517 , RIfe7d7f0_7772, \16328 );
and \g445953/U$3 ( \34518 , RIfe7d3b8_7769, \16334 );
and \g448819/U$2 ( \34519 , RIee2f968_5000, \16427 );
and \g448819/U$3 ( \34520 , \16448 , RIfc734c0_6334);
and \g448819/U$4 ( \34521 , RIfe7d520_7770, \16344 );
nor \g448819/U$1 ( \34522 , \34519 , \34520 , \34521 );
and \g455122/U$2 ( \34523 , \16317 , RIdf33310_1959);
and \g455122/U$3 ( \34524 , RIdf357a0_1985, \16325 );
nor \g455122/U$1 ( \34525 , \34523 , \34524 );
not \g455121/U$1 ( \34526 , \34525 );
and \g449844/U$2 ( \34527 , \34526 , \16336 );
and \g449844/U$3 ( \34528 , RIfebdd50_8280, \16356 );
nor \g449844/U$1 ( \34529 , \34527 , \34528 );
and \g451678/U$2 ( \34530 , \16361 , RIdf2f0f8_1912);
and \g451678/U$3 ( \34531 , RIdf312b8_1936, \16364 );
nor \g451678/U$1 ( \34532 , \34530 , \34531 );
and \g451676/U$2 ( \34533 , \16368 , RIee2d7a8_4976);
and \g451676/U$3 ( \34534 , RIfccfab8_7385, \16371 );
nor \g451676/U$1 ( \34535 , \34533 , \34534 );
nand \g448049/U$1 ( \34536 , \34522 , \34529 , \34532 , \34535 );
nor \g445953/U$1 ( \34537 , \34517 , \34518 , \34536 );
and \g451670/U$2 ( \34538 , \16377 , RIfceb9e8_7703);
and \g451670/U$3 ( \34539 , RIfebdbe8_8279, \16380 );
nor \g451670/U$1 ( \34540 , \34538 , \34539 );
nand \g445565/U$1 ( \34541 , \34516 , \34537 , \34540 );
and \g444767/U$2 ( \34542 , \34541 , \16394 );
and \g448814/U$2 ( \34543 , RIe14bed8_2241, \16398 );
and \g448814/U$3 ( \34544 , \16339 , RIfc649e8_6167);
and \g448814/U$4 ( \34545 , RIe15ccd8_2433, \16344 );
nor \g448814/U$1 ( \34546 , \34543 , \34544 , \34545 );
and \g454700/U$2 ( \34547 , \16317 , RIe1518d8_2305);
and \g454700/U$3 ( \34548 , RIfe7def8_7777, \16325 );
nor \g454700/U$1 ( \34549 , \34547 , \34548 );
not \g449839/U$3 ( \34550 , \34549 );
not \g449839/U$4 ( \34551 , \16351 );
and \g449839/U$2 ( \34552 , \34550 , \34551 );
and \g449839/U$5 ( \34553 , \16354 , RIee362e0_5075);
nor \g449839/U$1 ( \34554 , \34552 , \34553 );
and \g451659/U$2 ( \34555 , \16361 , RIe1464d8_2177);
and \g451659/U$3 ( \34556 , RIe1491d8_2209, \16364 );
nor \g451659/U$1 ( \34557 , \34555 , \34556 );
and \g451657/U$2 ( \34558 , \16368 , RIe14ebd8_2273);
and \g451657/U$3 ( \34559 , RIfebdeb8_8281, \16371 );
nor \g451657/U$1 ( \34560 , \34558 , \34559 );
nand \g447629/U$1 ( \34561 , \34546 , \34554 , \34557 , \34560 );
and \g444767/U$3 ( \34562 , \16390 , \34561 );
nor \g444767/U$1 ( \34563 , \34542 , \34562 );
and \g446733/U$2 ( \34564 , \18020 , RIe1626d8_2497);
and \g446733/U$3 ( \34565 , RIe1653d8_2529, \18022 );
nor \g446733/U$1 ( \34566 , \34564 , \34565 );
and \g446734/U$2 ( \34567 , \18025 , RIe15f9d8_2465);
and \g446734/U$3 ( \34568 , RIee373c0_5087, \18027 );
nor \g446734/U$1 ( \34569 , \34567 , \34568 );
and \g446736/U$2 ( \34570 , \18030 , RIe1545d8_2337);
and \g446736/U$3 ( \34571 , RIe1572d8_2369, \18032 );
nor \g446736/U$1 ( \34572 , \34570 , \34571 );
nand \g444479/U$1 ( \34573 , \34563 , \34566 , \34569 , \34572 );
and \g451699/U$2 ( \34574 , \16371 , RIfc787b8_6393);
and \g451699/U$3 ( \34575 , RIfc7aae0_6418, \16427 );
nor \g451699/U$1 ( \34576 , \34574 , \34575 );
and \g445959/U$2 ( \34577 , RIfcbf7f8_7201, \16448 );
and \g445959/U$3 ( \34578 , RIded2dd0_863, \16361 );
and \g448832/U$2 ( \34579 , RIee249a0_4875, \16319 );
and \g448832/U$3 ( \34580 , \16328 , RIee25648_4884);
and \g448832/U$4 ( \34581 , RIded72b8_912, \16398 );
nor \g448832/U$1 ( \34582 , \34579 , \34580 , \34581 );
and \g455149/U$2 ( \34583 , \16317 , RIfebe188_8283);
and \g455149/U$3 ( \34584 , RIfebe2f0_8284, \16325 );
nor \g455149/U$1 ( \34585 , \34583 , \34584 );
not \g449856/U$3 ( \34586 , \34585 );
not \g449856/U$4 ( \34587 , \16330 );
and \g449856/U$2 ( \34588 , \34586 , \34587 );
and \g449856/U$5 ( \34589 , \16341 , RIded98b0_939);
nor \g449856/U$1 ( \34590 , \34588 , \34589 );
and \g451709/U$2 ( \34591 , \16377 , RIee23488_4860);
and \g451709/U$3 ( \34592 , RIfebe020_8282, \16313 );
nor \g451709/U$1 ( \34593 , \34591 , \34592 );
and \g451712/U$2 ( \34594 , \16334 , RIfe7e060_7778);
and \g451712/U$3 ( \34595 , RIfe7e1c8_7779, \16380 );
nor \g451712/U$1 ( \34596 , \34594 , \34595 );
nand \g447302/U$1 ( \34597 , \34582 , \34590 , \34593 , \34596 );
nor \g445959/U$1 ( \34598 , \34577 , \34578 , \34597 );
and \g451702/U$2 ( \34599 , \16364 , RIded5530_891);
and \g451702/U$3 ( \34600 , RIfc618b0_6132, \16368 );
nor \g451702/U$1 ( \34601 , \34599 , \34600 );
nand \g445570/U$1 ( \34602 , \34576 , \34598 , \34601 );
and \g444911/U$2 ( \34603 , \34602 , \16477 );
and \g448824/U$2 ( \34604 , RIfe7ccb0_7764, \16485 );
and \g448824/U$3 ( \34605 , \16356 , RIfe7ce18_7765);
and \g448824/U$4 ( \34606 , RIfe7d250_7768, \16398 );
nor \g448824/U$1 ( \34607 , \34604 , \34605 , \34606 );
and \g454265/U$2 ( \34608 , \16317 , RIee2a238_4938);
and \g454265/U$3 ( \34609 , RIee2bcf0_4957, \16325 );
nor \g454265/U$1 ( \34610 , \34608 , \34609 );
not \g449850/U$3 ( \34611 , \34610 );
not \g449850/U$4 ( \34612 , \16311 );
and \g449850/U$2 ( \34613 , \34611 , \34612 );
and \g449850/U$5 ( \34614 , \16341 , RIee262f0_4893);
nor \g449850/U$1 ( \34615 , \34613 , \34614 );
and \g451688/U$2 ( \34616 , \16377 , RIee27c40_4911);
and \g451688/U$3 ( \34617 , RIee28e88_4924, \16313 );
nor \g451688/U$1 ( \34618 , \34616 , \34617 );
and \g451690/U$2 ( \34619 , \16334 , RIfe7cb48_7763);
and \g451690/U$3 ( \34620 , RIfe7cf80_7766, \16380 );
nor \g451690/U$1 ( \34621 , \34619 , \34620 );
nand \g447299/U$1 ( \34622 , \34607 , \34615 , \34618 , \34621 );
and \g444911/U$3 ( \34623 , \16481 , \34622 );
nor \g444911/U$1 ( \34624 , \34603 , \34623 );
and \g446747/U$2 ( \34625 , \17274 , RIee26e30_4901);
and \g446747/U$3 ( \34626 , RIee27268_4904, \17276 );
nor \g446747/U$1 ( \34627 , \34625 , \34626 );
and \g446749/U$2 ( \34628 , \17279 , RIfcaa0d8_6957);
and \g446749/U$3 ( \34629 , RIee26890_4897, \17281 );
nor \g446749/U$1 ( \34630 , \34628 , \34629 );
and \g446748/U$2 ( \34631 , \17284 , RIfe7d0e8_7767);
and \g446748/U$3 ( \34632 , RIee26020_4891, \17286 );
nor \g446748/U$1 ( \34633 , \34631 , \34632 );
nand \g444587/U$1 ( \34634 , \34624 , \34627 , \34630 , \34633 );
and \g445938/U$2 ( \34635 , RIdf16fa8_1638, \16328 );
and \g445938/U$3 ( \34636 , RIdf034a8_1414, \16334 );
and \g448801/U$2 ( \34637 , RIdeef9a8_1190, \16337 );
and \g448801/U$3 ( \34638 , \16341 , RIdef26a8_1222);
and \g448801/U$4 ( \34639 , RIdf08ea8_1478, \16485 );
nor \g448801/U$1 ( \34640 , \34637 , \34638 , \34639 );
and \g454421/U$2 ( \34641 , \16317 , RIdefada8_1318);
and \g454421/U$3 ( \34642 , RIdefdaa8_1350, \16325 );
nor \g454421/U$1 ( \34643 , \34641 , \34642 );
not \g449826/U$3 ( \34644 , \34643 );
not \g449826/U$4 ( \34645 , \16351 );
and \g449826/U$2 ( \34646 , \34644 , \34645 );
and \g449826/U$5 ( \34647 , \16356 , RIdf0bba8_1510);
nor \g449826/U$1 ( \34648 , \34646 , \34647 );
and \g451618/U$2 ( \34649 , \16361 , RIdee9fa8_1126);
and \g451618/U$3 ( \34650 , RIdeecca8_1158, \16364 );
nor \g451618/U$1 ( \34651 , \34649 , \34650 );
and \g451617/U$2 ( \34652 , \16368 , RIdef53a8_1254);
and \g451617/U$3 ( \34653 , RIdef80a8_1286, \16371 );
nor \g451617/U$1 ( \34654 , \34652 , \34653 );
nand \g447626/U$1 ( \34655 , \34640 , \34648 , \34651 , \34654 );
nor \g445938/U$1 ( \34656 , \34635 , \34636 , \34655 );
and \g451611/U$2 ( \34657 , \16377 , RIdf0e8a8_1542);
and \g451611/U$3 ( \34658 , RIdf061a8_1446, \16380 );
nor \g451611/U$1 ( \34659 , \34657 , \34658 );
and \g451607/U$2 ( \34660 , \16313 , RIdf115a8_1574);
and \g451607/U$3 ( \34661 , RIdf142a8_1606, \16321 );
nor \g451607/U$1 ( \34662 , \34660 , \34661 );
and \g445102/U$2 ( \34663 , \34656 , \34659 , \34662 );
nor \g445102/U$1 ( \34664 , \34663 , \16555 );
and \g445944/U$2 ( \34665 , RIe1437d8_2145, \16432 );
and \g445944/U$3 ( \34666 , RIde7c868_197, \16361 );
and \g448807/U$2 ( \34667 , RIdecdad8_804, \16321 );
and \g448807/U$3 ( \34668 , \16328 , RIded07d8_836);
and \g448807/U$4 ( \34669 , RIdee72a8_1094, \16398 );
nor \g448807/U$1 ( \34670 , \34667 , \34668 , \34669 );
and \g454620/U$2 ( \34671 , \16317 , RIde96920_324);
and \g454620/U$3 ( \34672 , RIdeb45d8_516, \16325 );
nor \g454620/U$1 ( \34673 , \34671 , \34672 );
not \g449834/U$3 ( \34674 , \34673 );
not \g449834/U$4 ( \34675 , \16330 );
and \g449834/U$2 ( \34676 , \34674 , \34675 );
and \g449834/U$5 ( \34677 , \16341 , RIdf007a8_1382);
nor \g449834/U$1 ( \34678 , \34676 , \34677 );
and \g451637/U$2 ( \34679 , \16377 , RIdec80d8_740);
and \g451637/U$3 ( \34680 , RIdecadd8_772, \16313 );
nor \g451637/U$1 ( \34681 , \34679 , \34680 );
and \g451639/U$2 ( \34682 , \16334 , RIe159fd8_2401);
and \g451639/U$3 ( \34683 , RIe16e1e0_2630, \16380 );
nor \g451639/U$1 ( \34684 , \34682 , \34683 );
nand \g447292/U$1 ( \34685 , \34670 , \34678 , \34681 , \34684 );
nor \g445944/U$1 ( \34686 , \34665 , \34666 , \34685 );
and \g451631/U$2 ( \34687 , \16364 , RIdedc010_967);
and \g451631/U$3 ( \34688 , RIdf1d0b0_1707, \16368 );
nor \g451631/U$1 ( \34689 , \34687 , \34688 );
and \g451630/U$2 ( \34690 , \16371 , RIdf2c830_1883);
and \g451630/U$3 ( \34691 , RIdf381d0_2015, \16427 );
nor \g451630/U$1 ( \34692 , \34690 , \34691 );
and \g445106/U$2 ( \34693 , \34686 , \34689 , \34692 );
nor \g445106/U$1 ( \34694 , \34693 , \16586 );
or \g444352/U$1 ( \34695 , \34573 , \34634 , \34664 , \34694 );
and \g445930/U$2 ( \34696 , RIee1cde0_4787, \16328 );
and \g445930/U$3 ( \34697 , RIfe7d958_7773, \16334 );
and \g448786/U$2 ( \34698 , RIee19e10_4753, \16427 );
and \g448786/U$3 ( \34699 , \16448 , RIee1a518_4758);
and \g448786/U$4 ( \34700 , RIde8d8c0_280, \16344 );
nor \g448786/U$1 ( \34701 , \34698 , \34699 , \34700 );
and \g455313/U$2 ( \34702 , \16317 , RIfe7dd90_7776);
and \g455313/U$3 ( \34703 , RIfcd05f8_7393, \16325 );
nor \g455313/U$1 ( \34704 , \34702 , \34703 );
not \g455312/U$1 ( \34705 , \34704 );
and \g449816/U$2 ( \34706 , \34705 , \16336 );
and \g449816/U$3 ( \34707 , RIde91088_297, \16354 );
nor \g449816/U$1 ( \34708 , \34706 , \34707 );
and \g451576/U$2 ( \34709 , \16361 , RIfe7dc28_7775);
and \g451576/U$3 ( \34710 , RIee38770_5101, \16364 );
nor \g451576/U$1 ( \34711 , \34709 , \34710 );
and \g451575/U$2 ( \34712 , \16368 , RIfc768c8_6371);
and \g451575/U$3 ( \34713 , RIee19b40_4751, \16371 );
nor \g451575/U$1 ( \34714 , \34712 , \34713 );
nand \g448043/U$1 ( \34715 , \34701 , \34708 , \34711 , \34714 );
nor \g445930/U$1 ( \34716 , \34696 , \34697 , \34715 );
and \g451571/U$2 ( \34717 , \16377 , RIfcd8a28_7487);
and \g451571/U$3 ( \34718 , RIfe7dac0_7774, \16380 );
nor \g451571/U$1 ( \34719 , \34717 , \34718 );
and \g451570/U$2 ( \34720 , \16313 , RIee1b490_4769);
and \g451570/U$3 ( \34721 , RIee1bd00_4775, \16319 );
nor \g451570/U$1 ( \34722 , \34720 , \34721 );
and \g445094/U$2 ( \34723 , \34716 , \34719 , \34722 );
nor \g445094/U$1 ( \34724 , \34723 , \16649 );
and \g445932/U$2 ( \34725 , RIee1ee38_4810, \16448 );
and \g445932/U$3 ( \34726 , RIde9d220_356, \16361 );
and \g448795/U$2 ( \34727 , RIdebccd8_612, \16344 );
and \g448795/U$3 ( \34728 , \16356 , RIee1f3d8_4814);
and \g448795/U$4 ( \34729 , RIdeaa420_420, \16398 );
nor \g448795/U$1 ( \34730 , \34727 , \34728 , \34729 );
and \g454601/U$2 ( \34731 , \16317 , RIdec26d8_676);
and \g454601/U$3 ( \34732 , RIdec53d8_708, \16325 );
nor \g454601/U$1 ( \34733 , \34731 , \34732 );
not \g449821/U$3 ( \34734 , \34733 );
not \g449821/U$4 ( \34735 , \16311 );
and \g449821/U$2 ( \34736 , \34734 , \34735 );
and \g449821/U$5 ( \34737 , \16341 , RIee1da88_4796);
nor \g449821/U$1 ( \34738 , \34736 , \34737 );
and \g451593/U$2 ( \34739 , \16377 , RIdebf9d8_644);
and \g451593/U$3 ( \34740 , RIee20080_4823, \16313 );
nor \g451593/U$1 ( \34741 , \34739 , \34740 );
and \g451596/U$2 ( \34742 , \16334 , RIdeb72d8_548);
and \g451596/U$3 ( \34743 , RIdeb9fd8_580, \16380 );
nor \g451596/U$1 ( \34744 , \34742 , \34743 );
nand \g447288/U$1 ( \34745 , \34730 , \34738 , \34741 , \34744 );
nor \g445932/U$1 ( \34746 , \34725 , \34726 , \34745 );
and \g451589/U$2 ( \34747 , \16364 , RIdea3b20_388);
and \g451589/U$3 ( \34748 , RIdeaebd8_452, \16368 );
nor \g451589/U$1 ( \34749 , \34747 , \34748 );
and \g451587/U$2 ( \34750 , \16371 , RIee1e898_4806);
and \g451587/U$3 ( \34751 , RIdeb18d8_484, \16427 );
nor \g451587/U$1 ( \34752 , \34750 , \34751 );
and \g445098/U$2 ( \34753 , \34746 , \34749 , \34752 );
nor \g445098/U$1 ( \34754 , \34753 , \16618 );
or \g444275/U$1 ( \34755 , \34695 , \34724 , \34754 );
_DC \g5a97/U$1 ( \34756 , \34755 , \16652 );
and \g446813/U$2 ( \34757 , \9724 , RIe197c70_3104);
and \g446813/U$3 ( \34758 , RIfe7b630_7748, \9726 );
nor \g446813/U$1 ( \34759 , \34757 , \34758 );
and \g446031/U$2 ( \34760 , RIe19d670_3168, \8351 );
and \g446031/U$3 ( \34761 , RIe19a970_3136, \8383 );
and \g448923/U$2 ( \34762 , RIe181470_2848, \8326 );
and \g448923/U$3 ( \34763 , \8531 , RIfe7b360_7746);
and \g448923/U$4 ( \34764 , RIe186e70_2912, \8488 );
nor \g448923/U$1 ( \34765 , \34762 , \34763 , \34764 );
and \g451979/U$2 ( \34766 , \8356 , RIe184170_2880);
and \g451979/U$3 ( \34767 , RIe189b70_2944, \8359 );
nor \g451979/U$1 ( \34768 , \34766 , \34767 );
and \g454795/U$2 ( \34769 , \8313 , RIe192270_3040);
and \g454795/U$3 ( \34770 , RIe194f70_3072, \8323 );
nor \g454795/U$1 ( \34771 , \34769 , \34770 );
not \g449936/U$3 ( \34772 , \34771 );
not \g449936/U$4 ( \34773 , \8376 );
and \g449936/U$2 ( \34774 , \34772 , \34773 );
and \g449936/U$5 ( \34775 , \8340 , RIfe7b1f8_7745);
nor \g449936/U$1 ( \34776 , \34774 , \34775 );
and \g451978/U$2 ( \34777 , \8378 , RIe18f570_3008);
and \g451978/U$3 ( \34778 , RIfe7b4c8_7747, \8417 );
nor \g451978/U$1 ( \34779 , \34777 , \34778 );
nand \g447681/U$1 ( \34780 , \34765 , \34768 , \34776 , \34779 );
nor \g446031/U$1 ( \34781 , \34760 , \34761 , \34780 );
not \g444817/U$3 ( \34782 , \34781 );
not \g444817/U$4 ( \34783 , \8589 );
and \g444817/U$2 ( \34784 , \34782 , \34783 );
and \g446034/U$2 ( \34785 , RIf140360_5190, \8371 );
and \g446034/U$3 ( \34786 , RIf140ea0_5198, \8383 );
and \g448928/U$2 ( \34787 , RIfe7ac58_7741, \8326 );
and \g448928/U$3 ( \34788 , \8531 , RIee39df0_5117);
and \g448928/U$4 ( \34789 , RIfe7af28_7743, \8488 );
nor \g448928/U$1 ( \34790 , \34787 , \34788 , \34789 );
and \g451999/U$2 ( \34791 , \8356 , RIe1737a8_2691);
and \g451999/U$3 ( \34792 , RIfe7b090_7744, \8359 );
nor \g451999/U$1 ( \34793 , \34791 , \34792 );
and \g455341/U$2 ( \34794 , \8313 , RIfc79460_6402);
and \g455341/U$3 ( \34795 , RIf13f280_5178, \8323 );
nor \g455341/U$1 ( \34796 , \34794 , \34795 );
not \g449942/U$3 ( \34797 , \34796 );
not \g449942/U$4 ( \34798 , \8376 );
and \g449942/U$2 ( \34799 , \34797 , \34798 );
and \g449942/U$5 ( \34800 , \8340 , RIfe7adc0_7742);
nor \g449942/U$1 ( \34801 , \34799 , \34800 );
and \g451998/U$2 ( \34802 , \8378 , RIee3d4c8_5156);
and \g451998/U$3 ( \34803 , RIf13fc58_5185, \8417 );
nor \g451998/U$1 ( \34804 , \34802 , \34803 );
nand \g447685/U$1 ( \34805 , \34790 , \34793 , \34801 , \34804 );
nor \g446034/U$1 ( \34806 , \34785 , \34786 , \34805 );
and \g453937/U$2 ( \34807 , \8335 , RIfcb20d0_7048);
and \g453937/U$3 ( \34808 , RIf1423b8_5213, \8351 );
nor \g453937/U$1 ( \34809 , \34807 , \34808 );
and \g451990/U$2 ( \34810 , \8319 , RIf16e440_5714);
and \g451990/U$3 ( \34811 , RIfe7b798_7749, \8404 );
nor \g451990/U$1 ( \34812 , \34810 , \34811 );
and \g445177/U$2 ( \34813 , \34806 , \34809 , \34812 );
nor \g445177/U$1 ( \34814 , \34813 , \8558 );
nor \g444817/U$1 ( \34815 , \34784 , \34814 );
and \g446812/U$2 ( \34816 , \9729 , RIe17ba70_2784);
and \g446812/U$3 ( \34817 , RIe17e770_2816, \9731 );
nor \g446812/U$1 ( \34818 , \34816 , \34817 );
nand \g444426/U$1 ( \34819 , \34759 , \34815 , \34818 );
and \g448934/U$2 ( \34820 , RIe2185c8_4567, \8414 );
and \g448934/U$3 ( \34821 , \8409 , RIe21dfc8_4631);
and \g448934/U$4 ( \34822 , RIe20d1c8_4439, \8326 );
nor \g448934/U$1 ( \34823 , \34820 , \34821 , \34822 );
and \g452019/U$2 ( \34824 , \8356 , RIe20fec8_4471);
and \g452019/U$3 ( \34825 , RIfebd7b0_8276, \8359 );
nor \g452019/U$1 ( \34826 , \34824 , \34825 );
and \g455139/U$2 ( \34827 , \8313 , RIfebd648_8275);
and \g455139/U$3 ( \34828 , RIe212bc8_4503, \8323 );
nor \g455139/U$1 ( \34829 , \34827 , \34828 );
not \g449948/U$3 ( \34830 , \34829 );
not \g449948/U$4 ( \34831 , \8347 );
and \g449948/U$2 ( \34832 , \34830 , \34831 );
and \g449948/U$5 ( \34833 , \8340 , RIfe7b900_7750);
nor \g449948/U$1 ( \34834 , \34832 , \34833 );
and \g452015/U$2 ( \34835 , \8378 , RIe2158c8_4535);
and \g452015/U$3 ( \34836 , RIf16aed0_5676, \8417 );
nor \g452015/U$1 ( \34837 , \34835 , \34836 );
nand \g447690/U$1 ( \34838 , \34823 , \34826 , \34834 , \34837 );
and \g444771/U$2 ( \34839 , \34838 , \8369 );
and \g446045/U$2 ( \34840 , RIe2024d0_4316, \8373 );
and \g446045/U$3 ( \34841 , RIf166178_5621, \8383 );
and \g448941/U$2 ( \34842 , RIf15b8b8_5501, \8326 );
and \g448941/U$3 ( \34843 , \8523 , RIfe7ba68_7751);
and \g448941/U$4 ( \34844 , RIf15e2e8_5531, \8488 );
nor \g448941/U$1 ( \34845 , \34842 , \34843 , \34844 );
and \g451434/U$2 ( \34846 , \8356 , RIfe7bea0_7754);
and \g451434/U$3 ( \34847 , RIf1601d8_5553, \8359 );
nor \g451434/U$1 ( \34848 , \34846 , \34847 );
and \g454728/U$2 ( \34849 , \8313 , RIfcd0a30_7396);
and \g454728/U$3 ( \34850 , RIf1646c0_5602, \8323 );
nor \g454728/U$1 ( \34851 , \34849 , \34850 );
not \g449955/U$3 ( \34852 , \34851 );
not \g449955/U$4 ( \34853 , \8376 );
and \g449955/U$2 ( \34854 , \34852 , \34853 );
and \g449955/U$5 ( \34855 , \8340 , RIf15cdd0_5516);
nor \g449955/U$1 ( \34856 , \34854 , \34855 );
and \g452032/U$2 ( \34857 , \8378 , RIf1620c8_5575);
and \g452032/U$3 ( \34858 , RIf165368_5611, \8417 );
nor \g452032/U$1 ( \34859 , \34857 , \34858 );
nand \g447695/U$1 ( \34860 , \34845 , \34848 , \34856 , \34859 );
nor \g446045/U$1 ( \34861 , \34840 , \34841 , \34860 );
and \g452028/U$2 ( \34862 , \8335 , RIfca4840_6894);
and \g452028/U$3 ( \34863 , RIf167258_5633, \8351 );
nor \g452028/U$1 ( \34864 , \34862 , \34863 );
and \g452064/U$2 ( \34865 , \8319 , RIf15a7d8_5489);
and \g452064/U$3 ( \34866 , RIfe7bbd0_7752, \8404 );
nor \g452064/U$1 ( \34867 , \34865 , \34866 );
and \g445183/U$2 ( \34868 , \34861 , \34864 , \34867 );
nor \g445183/U$1 ( \34869 , \34868 , \8422 );
nor \g444771/U$1 ( \34870 , \34839 , \34869 );
and \g446824/U$2 ( \34871 , \8426 , RIe220cc8_4663);
and \g446824/U$3 ( \34872 , RIf16be48_5687, \8428 );
nor \g446824/U$1 ( \34873 , \34871 , \34872 );
and \g446823/U$2 ( \34874 , \13735 , RIe2239c8_4695);
and \g446823/U$3 ( \34875 , RIfe7bd38_7753, \13737 );
nor \g446823/U$1 ( \34876 , \34874 , \34875 );
and \g446825/U$2 ( \34877 , \8707 , RIe2077c8_4375);
and \g446825/U$3 ( \34878 , RIe20a4c8_4407, \8709 );
nor \g446825/U$1 ( \34879 , \34877 , \34878 );
nand \g444488/U$1 ( \34880 , \34870 , \34873 , \34876 , \34879 );
and \g446021/U$2 ( \34881 , RIfebda80_8278, \8373 );
and \g446021/U$3 ( \34882 , RIf14b8c8_5319, \8383 );
and \g448910/U$2 ( \34883 , RIfe7c9e0_7762, \8414 );
and \g448910/U$3 ( \34884 , \8407 , RIfe7c2d8_7757);
and \g448910/U$4 ( \34885 , RIf146738_5261, \8324 );
nor \g448910/U$1 ( \34886 , \34883 , \34884 , \34885 );
and \g451938/U$2 ( \34887 , \8356 , RIfebd918_8277);
and \g451938/U$3 ( \34888 , RIf149000_5290, \8359 );
nor \g451938/U$1 ( \34889 , \34887 , \34888 );
and \g454333/U$2 ( \34890 , \8313 , RIe1b2688_3407);
and \g454333/U$3 ( \34891 , RIf147db8_5277, \8323 );
nor \g454333/U$1 ( \34892 , \34890 , \34891 );
not \g449928/U$3 ( \34893 , \34892 );
not \g449928/U$4 ( \34894 , \8347 );
and \g449928/U$2 ( \34895 , \34893 , \34894 );
and \g449928/U$5 ( \34896 , \8340 , RIfe7c5a8_7759);
nor \g449928/U$1 ( \34897 , \34895 , \34896 );
and \g451700/U$2 ( \34898 , \8378 , RIfe7c440_7758);
and \g451700/U$3 ( \34899 , RIf14a680_5306, \8417 );
nor \g451700/U$1 ( \34900 , \34898 , \34899 );
nand \g447671/U$1 ( \34901 , \34886 , \34889 , \34897 , \34900 );
nor \g446021/U$1 ( \34902 , \34881 , \34882 , \34901 );
and \g451931/U$2 ( \34903 , \8335 , RIe1aad98_3321);
and \g451931/U$3 ( \34904 , RIf14cb10_5332, \8351 );
nor \g451931/U$1 ( \34905 , \34903 , \34904 );
and \g451934/U$2 ( \34906 , \8319 , RIfe7c710_7760);
and \g451934/U$3 ( \34907 , RIfe7c878_7761, \8404 );
nor \g451934/U$1 ( \34908 , \34906 , \34907 );
and \g445165/U$2 ( \34909 , \34902 , \34905 , \34908 );
nor \g445165/U$1 ( \34910 , \34909 , \8481 );
and \g446025/U$2 ( \34911 , RIe1d7c30_3832, \8378 );
and \g446025/U$3 ( \34912 , RIe1d2230_3768, \8359 );
and \g448915/U$2 ( \34913 , RIe1c1430_3576, \8319 );
and \g448915/U$3 ( \34914 , \8326 , RIe1c4130_3608);
and \g448915/U$4 ( \34915 , RIe1dd630_3896, \8409 );
nor \g448915/U$1 ( \34916 , \34913 , \34914 , \34915 );
and \g451960/U$2 ( \34917 , \8335 , RIe1be730_3544);
and \g451960/U$3 ( \34918 , RIe1c6e30_3640, \8340 );
nor \g451960/U$1 ( \34919 , \34917 , \34918 );
and \g451959/U$2 ( \34920 , \8404 , RIe1e3030_3960);
and \g451959/U$3 ( \34921 , RIe1eb730_4056, \8351 );
nor \g451959/U$1 ( \34922 , \34920 , \34921 );
and \g454311/U$2 ( \34923 , \8313 , RIe1e5d30_3992);
and \g454311/U$3 ( \34924 , RIe1e8a30_4024, \8323 );
nor \g454311/U$1 ( \34925 , \34923 , \34924 );
not \g449932/U$3 ( \34926 , \34925 );
not \g449932/U$4 ( \34927 , \8328 );
and \g449932/U$2 ( \34928 , \34926 , \34927 );
and \g449932/U$5 ( \34929 , \8417 , RIe1e0330_3928);
nor \g449932/U$1 ( \34930 , \34928 , \34929 );
nand \g447677/U$1 ( \34931 , \34916 , \34919 , \34922 , \34930 );
nor \g446025/U$1 ( \34932 , \34911 , \34912 , \34931 );
and \g451953/U$2 ( \34933 , \8356 , RIe1c9b30_3672);
and \g451953/U$3 ( \34934 , RIe1da930_3864, \8414 );
nor \g451953/U$1 ( \34935 , \34933 , \34934 );
and \g451951/U$2 ( \34936 , \8531 , RIe1cc830_3704);
and \g451951/U$3 ( \34937 , RIe1cf530_3736, \8488 );
nor \g451951/U$1 ( \34938 , \34936 , \34937 );
and \g445168/U$2 ( \34939 , \34932 , \34935 , \34938 );
nor \g445168/U$1 ( \34940 , \34939 , \8477 );
or \g444295/U$1 ( \34941 , \34819 , \34880 , \34910 , \34940 );
and \g446018/U$2 ( \34942 , RIe1a3070_3232, \8373 );
and \g446018/U$3 ( \34943 , RIe1a5d70_3264, \8383 );
and \g448902/U$2 ( \34944 , RIe1bba30_3512, \8326 );
and \g448902/U$3 ( \34945 , \8531 , RIe1f7ee0_4198);
and \g448902/U$4 ( \34946 , RIe1feb28_4275, \8488 );
nor \g448902/U$1 ( \34947 , \34944 , \34945 , \34946 );
and \g451922/U$2 ( \34948 , \8356 , RIe1f0a28_4115);
and \g451922/U$3 ( \34949 , RIe204ac8_4343, \8359 );
nor \g451922/U$1 ( \34950 , \34948 , \34949 );
and \g454691/U$2 ( \34951 , \8313 , RIe2266c8_4727);
and \g454691/U$3 ( \34952 , RIe178d70_2752, \8323 );
nor \g454691/U$1 ( \34953 , \34951 , \34952 );
not \g449920/U$3 ( \34954 , \34953 );
not \g449920/U$4 ( \34955 , \8376 );
and \g449920/U$2 ( \34956 , \34954 , \34955 );
and \g449920/U$5 ( \34957 , \8340 , RIe1d4f30_3800);
nor \g449920/U$1 ( \34958 , \34956 , \34957 );
and \g452276/U$2 ( \34959 , \8378 , RIe21b2c8_4599);
and \g452276/U$3 ( \34960 , RIe18c870_2976, \8417 );
nor \g452276/U$1 ( \34961 , \34959 , \34960 );
nand \g447668/U$1 ( \34962 , \34947 , \34950 , \34958 , \34961 );
nor \g446018/U$1 ( \34963 , \34942 , \34943 , \34962 );
and \g451911/U$2 ( \34964 , \8335 , RIe170ee0_2662);
and \g451911/U$3 ( \34965 , RIe1a8a70_3296, \8351 );
nor \g451911/U$1 ( \34966 , \34964 , \34965 );
and \g451915/U$2 ( \34967 , \8319 , RIe1ae8a8_3363);
and \g451915/U$3 ( \34968 , RIe1a0370_3200, \8404 );
nor \g451915/U$1 ( \34969 , \34967 , \34968 );
and \g445163/U$2 ( \34970 , \34963 , \34966 , \34969 );
nor \g445163/U$1 ( \34971 , \34970 , \8651 );
and \g446009/U$2 ( \34972 , RIf156f98_5449, \8371 );
and \g446009/U$3 ( \34973 , RIf157c40_5458, \8330 );
and \g448894/U$2 ( \34974 , RIf1549a0_5422, \8414 );
and \g448894/U$3 ( \34975 , \8409 , RIf155918_5433);
and \g448894/U$4 ( \34976 , RIf14ee38_5357, \8326 );
nor \g448894/U$1 ( \34977 , \34974 , \34975 , \34976 );
and \g451900/U$2 ( \34978 , \8356 , RIe1f32f0_4144);
and \g451900/U$3 ( \34979 , RIfe7c008_7755, \8359 );
nor \g451900/U$1 ( \34980 , \34978 , \34979 );
and \g455197/U$2 ( \34981 , \8313 , RIf150bc0_5378);
and \g455197/U$3 ( \34982 , RIf151b38_5389, \8323 );
nor \g455197/U$1 ( \34983 , \34981 , \34982 );
not \g449915/U$3 ( \34984 , \34983 );
not \g449915/U$4 ( \34985 , \8347 );
and \g449915/U$2 ( \34986 , \34984 , \34985 );
and \g449915/U$5 ( \34987 , \8340 , RIf14fae0_5366);
nor \g449915/U$1 ( \34988 , \34986 , \34987 );
and \g452947/U$2 ( \34989 , \8378 , RIe1f54b0_4168);
and \g452947/U$3 ( \34990 , RIf156458_5441, \8417 );
nor \g452947/U$1 ( \34991 , \34989 , \34990 );
nand \g447833/U$1 ( \34992 , \34977 , \34980 , \34988 , \34991 );
nor \g446009/U$1 ( \34993 , \34972 , \34973 , \34992 );
and \g453174/U$2 ( \34994 , \8335 , RIe1edff8_4085);
and \g453174/U$3 ( \34995 , RIf158ff0_5472, \8351 );
nor \g453174/U$1 ( \34996 , \34994 , \34995 );
and \g453059/U$2 ( \34997 , \8319 , RIf14e028_5347);
and \g453059/U$3 ( \34998 , RIfe7c170_7756, \8404 );
nor \g453059/U$1 ( \34999 , \34997 , \34998 );
and \g445156/U$2 ( \35000 , \34993 , \34996 , \34999 );
nor \g445156/U$1 ( \35001 , \35000 , \8621 );
or \g444162/U$1 ( \35002 , \34941 , \34971 , \35001 );
_DC \g5b1b/U$1 ( \35003 , \35002 , \8654 );
and \g452674/U$2 ( \35004 , \16313 , RIfc7dab0_6452);
and \g452674/U$3 ( \35005 , RIfca19d8_6861, \16321 );
nor \g452674/U$1 ( \35006 , \35004 , \35005 );
and \g446191/U$2 ( \35007 , RIfc7e1b8_6457, \16328 );
and \g446191/U$3 ( \35008 , RIfe80bf8_7809, \16334 );
and \g449123/U$2 ( \35009 , RIded7420_913, \16398 );
and \g449123/U$3 ( \35010 , \16339 , RIfe81030_7812);
and \g449123/U$4 ( \35011 , RIfe80d60_7810, \16485 );
nor \g449123/U$1 ( \35012 , \35009 , \35010 , \35011 );
and \g455363/U$2 ( \35013 , \16317 , RIfce9f30_7684);
and \g455363/U$3 ( \35014 , RIfcb3750_7064, \16325 );
nor \g455363/U$1 ( \35015 , \35013 , \35014 );
not \g450137/U$3 ( \35016 , \35015 );
not \g450137/U$4 ( \35017 , \16351 );
and \g450137/U$2 ( \35018 , \35016 , \35017 );
and \g450137/U$5 ( \35019 , \16354 , RIdee49e0_1065);
nor \g450137/U$1 ( \35020 , \35018 , \35019 );
and \g452682/U$2 ( \35021 , \16361 , RIded2f38_864);
and \g452682/U$3 ( \35022 , RIfe80ec8_7811, \16364 );
nor \g452682/U$1 ( \35023 , \35021 , \35022 );
and \g452681/U$2 ( \35024 , \16368 , RIfc56a50_6008);
and \g452681/U$3 ( \35025 , RIfc7e5f0_6460, \16371 );
nor \g452681/U$1 ( \35026 , \35024 , \35025 );
nand \g447786/U$1 ( \35027 , \35012 , \35020 , \35023 , \35026 );
nor \g446191/U$1 ( \35028 , \35007 , \35008 , \35027 );
and \g452677/U$2 ( \35029 , \16377 , RIfc7e488_6459);
and \g452677/U$3 ( \35030 , RIfeabba0_8270, \16380 );
nor \g452677/U$1 ( \35031 , \35029 , \35030 );
nand \g445621/U$1 ( \35032 , \35006 , \35028 , \35031 );
and \g444918/U$2 ( \35033 , \35032 , \16477 );
and \g449120/U$2 ( \35034 , RIfce7ed8_7661, \16427 );
and \g449120/U$3 ( \35035 , \16448 , RIfc84428_6527);
and \g449120/U$4 ( \35036 , RIdf28078_1832, \16485 );
nor \g449120/U$1 ( \35037 , \35034 , \35035 , \35036 );
and \g455100/U$2 ( \35038 , \16317 , RIdf1f978_1736);
and \g455100/U$3 ( \35039 , RIdf21868_1758, \16325 );
nor \g455100/U$1 ( \35040 , \35038 , \35039 );
not \g455099/U$1 ( \35041 , \35040 );
and \g450134/U$2 ( \35042 , \35041 , \16336 );
and \g450134/U$3 ( \35043 , RIdf2a3a0_1857, \16356 );
nor \g450134/U$1 ( \35044 , \35042 , \35043 );
and \g452666/U$2 ( \35045 , \16361 , RIdf192d0_1663);
and \g452666/U$3 ( \35046 , RIdf1b058_1684, \16364 );
nor \g452666/U$1 ( \35047 , \35045 , \35046 );
and \g452665/U$2 ( \35048 , \16368 , RIfc515f0_5948);
and \g452665/U$3 ( \35049 , RIdf22d80_1773, \16371 );
nor \g452665/U$1 ( \35050 , \35048 , \35049 );
nand \g448084/U$1 ( \35051 , \35037 , \35044 , \35047 , \35050 );
and \g444918/U$3 ( \35052 , \16481 , \35051 );
nor \g444918/U$1 ( \35053 , \35033 , \35052 );
and \g446957/U$2 ( \35054 , \16505 , RIee2a3a0_4939);
and \g446957/U$3 ( \35055 , RIfcb7968_7111, \16507 );
nor \g446957/U$1 ( \35056 , \35054 , \35055 );
and \g446959/U$2 ( \35057 , \16511 , RIdf24838_1792);
and \g446959/U$3 ( \35058 , RIfe81198_7813, \16514 );
nor \g446959/U$1 ( \35059 , \35057 , \35058 );
and \g446958/U$2 ( \35060 , \16518 , RIfcd3fa0_7434);
and \g446958/U$3 ( \35061 , RIfc51050_5944, \16521 );
nor \g446958/U$1 ( \35062 , \35060 , \35061 );
nand \g444626/U$1 ( \35063 , \35053 , \35056 , \35059 , \35062 );
and \g452705/U$2 ( \35064 , \16371 , RIdf2c998_1884);
and \g452705/U$3 ( \35065 , RIdf38338_2016, \16427 );
nor \g452705/U$1 ( \35066 , \35064 , \35065 );
and \g446195/U$2 ( \35067 , RIe143940_2146, \16448 );
and \g446195/U$3 ( \35068 , RIde7cbb0_198, \16361 );
and \g449131/U$2 ( \35069 , RIdecdc40_805, \16321 );
and \g449131/U$3 ( \35070 , \16328 , RIded0940_837);
and \g449131/U$4 ( \35071 , RIdee7410_1095, \16337 );
nor \g449131/U$1 ( \35072 , \35069 , \35070 , \35071 );
and \g455349/U$2 ( \35073 , \16317 , RIde96c68_325);
and \g455349/U$3 ( \35074 , RIdeb4740_517, \16325 );
nor \g455349/U$1 ( \35075 , \35073 , \35074 );
not \g450145/U$3 ( \35076 , \35075 );
not \g450145/U$4 ( \35077 , \16330 );
and \g450145/U$2 ( \35078 , \35076 , \35077 );
and \g450145/U$5 ( \35079 , \16339 , RIdf00910_1383);
nor \g450145/U$1 ( \35080 , \35078 , \35079 );
and \g452712/U$2 ( \35081 , \16377 , RIdec8240_741);
and \g452712/U$3 ( \35082 , RIdecaf40_773, \16313 );
nor \g452712/U$1 ( \35083 , \35081 , \35082 );
and \g452713/U$2 ( \35084 , \16334 , RIe15a140_2402);
and \g452713/U$3 ( \35085 , RIe16e348_2631, \16380 );
nor \g452713/U$1 ( \35086 , \35084 , \35085 );
nand \g447372/U$1 ( \35087 , \35072 , \35080 , \35083 , \35086 );
nor \g446195/U$1 ( \35088 , \35067 , \35068 , \35087 );
and \g452706/U$2 ( \35089 , \16364 , RIdedc178_968);
and \g452706/U$3 ( \35090 , RIdf1d218_1708, \16368 );
nor \g452706/U$1 ( \35091 , \35089 , \35090 );
nand \g445622/U$1 ( \35092 , \35066 , \35088 , \35091 );
and \g444784/U$2 ( \35093 , \35092 , \16752 );
and \g449127/U$2 ( \35094 , RIdeefb10_1191, \16398 );
and \g449127/U$3 ( \35095 , \16341 , RIdef2810_1223);
and \g449127/U$4 ( \35096 , RIdf09010_1479, \16344 );
nor \g449127/U$1 ( \35097 , \35094 , \35095 , \35096 );
and \g454970/U$2 ( \35098 , \16317 , RIdefaf10_1319);
and \g454970/U$3 ( \35099 , RIdefdc10_1351, \16325 );
nor \g454970/U$1 ( \35100 , \35098 , \35099 );
not \g450142/U$3 ( \35101 , \35100 );
not \g450142/U$4 ( \35102 , \16351 );
and \g450142/U$2 ( \35103 , \35101 , \35102 );
and \g450142/U$5 ( \35104 , \16356 , RIdf0bd10_1511);
nor \g450142/U$1 ( \35105 , \35103 , \35104 );
and \g452700/U$2 ( \35106 , \16361 , RIdeea110_1127);
and \g452700/U$3 ( \35107 , RIdeece10_1159, \16364 );
nor \g452700/U$1 ( \35108 , \35106 , \35107 );
and \g452698/U$2 ( \35109 , \16368 , RIdef5510_1255);
and \g452698/U$3 ( \35110 , RIdef8210_1287, \16371 );
nor \g452698/U$1 ( \35111 , \35109 , \35110 );
nand \g447790/U$1 ( \35112 , \35097 , \35105 , \35108 , \35111 );
and \g444784/U$3 ( \35113 , \16750 , \35112 );
nor \g444784/U$1 ( \35114 , \35093 , \35113 );
and \g446962/U$2 ( \35115 , \19457 , RIdf14410_1607);
and \g446962/U$3 ( \35116 , RIdf17110_1639, \19459 );
nor \g446962/U$1 ( \35117 , \35115 , \35116 );
and \g446964/U$2 ( \35118 , \19462 , RIdf03610_1415);
and \g446964/U$3 ( \35119 , RIdf06310_1447, \19464 );
nor \g446964/U$1 ( \35120 , \35118 , \35119 );
and \g446963/U$2 ( \35121 , \19467 , RIdf0ea10_1543);
and \g446963/U$3 ( \35122 , RIdf11710_1575, \19469 );
nor \g446963/U$1 ( \35123 , \35121 , \35122 );
nand \g444627/U$1 ( \35124 , \35114 , \35117 , \35120 , \35123 );
and \g446181/U$2 ( \35125 , RIe165540_2530, \16328 );
and \g446181/U$3 ( \35126 , RIe154740_2338, \16334 );
and \g449113/U$2 ( \35127 , RIe151a40_2306, \16427 );
and \g449113/U$3 ( \35128 , \16448 , RIfcd35c8_7427);
and \g449113/U$4 ( \35129 , RIe15ce40_2434, \16485 );
nor \g449113/U$1 ( \35130 , \35127 , \35128 , \35129 );
and \g454951/U$2 ( \35131 , \16317 , RIe14c040_2242);
and \g454951/U$3 ( \35132 , RIfcc6170_7276, \16325 );
nor \g454951/U$1 ( \35133 , \35131 , \35132 );
not \g454950/U$1 ( \35134 , \35133 );
and \g450128/U$2 ( \35135 , \35134 , \16336 );
and \g450128/U$3 ( \35136 , RIfcb5be0_7090, \16356 );
nor \g450128/U$1 ( \35137 , \35135 , \35136 );
and \g452644/U$2 ( \35138 , \16361 , RIe146640_2178);
and \g452644/U$3 ( \35139 , RIe149340_2210, \16364 );
nor \g452644/U$1 ( \35140 , \35138 , \35139 );
and \g452642/U$2 ( \35141 , \16368 , RIe14ed40_2274);
and \g452642/U$3 ( \35142 , RIfc53a80_5974, \16371 );
nor \g452642/U$1 ( \35143 , \35141 , \35142 );
nand \g448083/U$1 ( \35144 , \35130 , \35137 , \35140 , \35143 );
nor \g446181/U$1 ( \35145 , \35125 , \35126 , \35144 );
and \g452639/U$2 ( \35146 , \16377 , RIe15fb40_2466);
and \g452639/U$3 ( \35147 , RIe157440_2370, \16380 );
nor \g452639/U$1 ( \35148 , \35146 , \35147 );
and \g452638/U$2 ( \35149 , \16313 , RIee37528_5088);
and \g452638/U$3 ( \35150 , RIe162840_2498, \16321 );
nor \g452638/U$1 ( \35151 , \35149 , \35150 );
and \g445282/U$2 ( \35152 , \35145 , \35148 , \35151 );
nor \g445282/U$1 ( \35153 , \35152 , \16389 );
and \g446184/U$2 ( \35154 , RIfc7fc70_6476, \16448 );
and \g446184/U$3 ( \35155 , RIdf2f260_1913, \16361 );
and \g449117/U$2 ( \35156 , RIee33310_5041, \16319 );
and \g449117/U$3 ( \35157 , \16326 , RIfc7f130_6468);
and \g449117/U$4 ( \35158 , RIdf33478_1960, \16398 );
nor \g449117/U$1 ( \35159 , \35156 , \35157 , \35158 );
and \g455071/U$2 ( \35160 , \16317 , RIdf3ee18_2092);
and \g455071/U$3 ( \35161 , RIe140f10_2116, \16325 );
nor \g455071/U$1 ( \35162 , \35160 , \35161 );
not \g450131/U$3 ( \35163 , \35162 );
not \g450131/U$4 ( \35164 , \16330 );
and \g450131/U$2 ( \35165 , \35163 , \35164 );
and \g450131/U$5 ( \35166 , \16341 , RIdf35908_1986);
nor \g450131/U$1 ( \35167 , \35165 , \35166 );
and \g452654/U$2 ( \35168 , \16377 , RIfc47f78_5841);
and \g452654/U$3 ( \35169 , RIfcb4f38_7081, \16313 );
nor \g452654/U$1 ( \35170 , \35168 , \35169 );
and \g452656/U$2 ( \35171 , \16334 , RIdf3a7c8_2042);
and \g452656/U$3 ( \35172 , RIdf3cc58_2068, \16380 );
nor \g452656/U$1 ( \35173 , \35171 , \35172 );
nand \g447366/U$1 ( \35174 , \35159 , \35167 , \35170 , \35173 );
nor \g446184/U$1 ( \35175 , \35154 , \35155 , \35174 );
and \g452650/U$2 ( \35176 , \16364 , RIfebe9f8_8289);
and \g452650/U$3 ( \35177 , RIfcc6b48_7283, \16368 );
nor \g452650/U$1 ( \35178 , \35176 , \35177 );
and \g452649/U$2 ( \35179 , \16371 , RIfca1000_6854);
and \g452649/U$3 ( \35180 , RIfcd27b8_7417, \16427 );
nor \g452649/U$1 ( \35181 , \35179 , \35180 );
and \g445283/U$2 ( \35182 , \35175 , \35178 , \35181 );
nor \g445283/U$1 ( \35183 , \35182 , \16393 );
or \g444343/U$1 ( \35184 , \35063 , \35124 , \35153 , \35183 );
and \g446175/U$2 ( \35185 , RIdec5540_709, \16326 );
and \g446175/U$3 ( \35186 , RIdeb7440_549, \16334 );
and \g449107/U$2 ( \35187 , RIdeb1a40_485, \16427 );
and \g449107/U$3 ( \35188 , \16448 , RIfc4d978_5905);
and \g449107/U$4 ( \35189 , RIdebce40_613, \16344 );
nor \g449107/U$1 ( \35190 , \35187 , \35188 , \35189 );
and \g454940/U$2 ( \35191 , \16317 , RIdeaa768_421);
and \g454940/U$3 ( \35192 , RIfcb8610_7120, \16325 );
nor \g454940/U$1 ( \35193 , \35191 , \35192 );
not \g454939/U$1 ( \35194 , \35193 );
and \g450121/U$2 ( \35195 , \35194 , \16336 );
and \g450121/U$3 ( \35196 , RIfc9d7c0_6814, \16356 );
nor \g450121/U$1 ( \35197 , \35195 , \35196 );
and \g452618/U$2 ( \35198 , \16361 , RIde9d568_357);
and \g452618/U$3 ( \35199 , RIdea3e68_389, \16364 );
nor \g452618/U$1 ( \35200 , \35198 , \35199 );
and \g452616/U$2 ( \35201 , \16368 , RIdeaed40_453);
and \g452616/U$3 ( \35202 , RIfc9dbf8_6817, \16371 );
nor \g452616/U$1 ( \35203 , \35201 , \35202 );
nand \g448081/U$1 ( \35204 , \35190 , \35197 , \35200 , \35203 );
nor \g446175/U$1 ( \35205 , \35185 , \35186 , \35204 );
and \g452613/U$2 ( \35206 , \16377 , RIdebfb40_645);
and \g452613/U$3 ( \35207 , RIdeba140_581, \16380 );
nor \g452613/U$1 ( \35208 , \35206 , \35207 );
and \g452612/U$2 ( \35209 , \16313 , RIfcc4dc0_7262);
and \g452612/U$3 ( \35210 , RIdec2840_677, \16321 );
nor \g452612/U$1 ( \35211 , \35209 , \35210 );
and \g445275/U$2 ( \35212 , \35205 , \35208 , \35211 );
nor \g445275/U$1 ( \35213 , \35212 , \16618 );
and \g446180/U$2 ( \35214 , RIfc50678_5937, \16328 );
and \g446180/U$3 ( \35215 , RIde858c8_241, \16334 );
and \g449110/U$2 ( \35216 , RIe16b7b0_2600, \16337 );
and \g449110/U$3 ( \35217 , \16339 , RIfcb7da0_7114);
and \g449110/U$4 ( \35218 , RIde8dc08_281, \16485 );
nor \g449110/U$1 ( \35219 , \35216 , \35217 , \35218 );
and \g454945/U$2 ( \35220 , \16317 , RIfc84860_6530);
and \g454945/U$3 ( \35221 , RIde81a70_222, \16325 );
nor \g454945/U$1 ( \35222 , \35220 , \35221 );
not \g450124/U$3 ( \35223 , \35222 );
not \g450124/U$4 ( \35224 , \16351 );
and \g450124/U$2 ( \35225 , \35223 , \35224 );
and \g450124/U$5 ( \35226 , \16356 , RIde913d0_298);
nor \g450124/U$1 ( \35227 , \35225 , \35226 );
and \g452631/U$2 ( \35228 , \16361 , RIe167e08_2559);
and \g452631/U$3 ( \35229 , RIe169b90_2580, \16364 );
nor \g452631/U$1 ( \35230 , \35228 , \35229 );
and \g452630/U$2 ( \35231 , \16368 , RIfc84c98_6533);
and \g452630/U$3 ( \35232 , RIfc50948_5939, \16371 );
nor \g452630/U$1 ( \35233 , \35231 , \35232 );
nand \g447784/U$1 ( \35234 , \35219 , \35227 , \35230 , \35233 );
nor \g446180/U$1 ( \35235 , \35214 , \35215 , \35234 );
and \g452627/U$2 ( \35236 , \16377 , RIfc853a0_6538);
and \g452627/U$3 ( \35237 , RIde89a68_261, \16380 );
nor \g452627/U$1 ( \35238 , \35236 , \35237 );
and \g452625/U$2 ( \35239 , \16313 , RIfc9dec8_6819);
and \g452625/U$3 ( \35240 , RIfc507e0_5938, \16319 );
nor \g452625/U$1 ( \35241 , \35239 , \35240 );
and \g445280/U$2 ( \35242 , \35235 , \35238 , \35241 );
nor \g445280/U$1 ( \35243 , \35242 , \16649 );
or \g444278/U$1 ( \35244 , \35184 , \35213 , \35243 );
_DC \g5ba0/U$1 ( \35245 , \35244 , \16652 );
and \g452816/U$2 ( \35246 , \8324 , RIfcb7f08_7115);
and \g452816/U$3 ( \35247 , RIfebe458_8285, \8356 );
nor \g452816/U$1 ( \35248 , \35246 , \35247 );
and \g446217/U$2 ( \35249 , RIf150d28_5379, \8531 );
and \g446217/U$3 ( \35250 , RIf14e190_5348, \8319 );
and \g449161/U$2 ( \35251 , RIfcb9f60_7138, \8373 );
and \g449161/U$3 ( \35252 , \8330 , RIf157da8_5459);
and \g449161/U$4 ( \35253 , RIfcc4988_7259, \8488 );
nor \g449161/U$1 ( \35254 , \35251 , \35252 , \35253 );
and \g455039/U$2 ( \35255 , \8313 , RIfc9f6b0_6836);
and \g455039/U$3 ( \35256 , RIfc529a0_5962, \8323 );
nor \g455039/U$1 ( \35257 , \35255 , \35256 );
not \g450176/U$3 ( \35258 , \35257 );
not \g450176/U$4 ( \35259 , \8376 );
and \g450176/U$2 ( \35260 , \35258 , \35259 );
and \g450176/U$5 ( \35261 , \8359 , RIf153320_5406);
nor \g450176/U$1 ( \35262 , \35260 , \35261 );
and \g452825/U$2 ( \35263 , \8404 , RIe1fa208_4223);
and \g452825/U$3 ( \35264 , RIfc9e468_6823, \8351 );
nor \g452825/U$1 ( \35265 , \35263 , \35264 );
and \g452826/U$2 ( \35266 , \8378 , RIe1f5618_4169);
and \g452826/U$3 ( \35267 , RIfc849c8_6531, \8417 );
nor \g452826/U$1 ( \35268 , \35266 , \35267 );
nand \g447807/U$1 ( \35269 , \35254 , \35262 , \35265 , \35268 );
nor \g446217/U$1 ( \35270 , \35249 , \35250 , \35269 );
and \g452818/U$2 ( \35271 , \8335 , RIfe80658_7805);
and \g452818/U$3 ( \35272 , RIfc87f38_6569, \8340 );
nor \g452818/U$1 ( \35273 , \35271 , \35272 );
nand \g445634/U$1 ( \35274 , \35248 , \35270 , \35273 );
and \g444726/U$2 ( \35275 , \35274 , \8752 );
and \g449157/U$2 ( \35276 , RIe1daa98_3865, \8414 );
and \g449157/U$3 ( \35277 , \8409 , RIe1dd798_3897);
and \g449157/U$4 ( \35278 , RIe1cf698_3737, \8486 );
nor \g449157/U$1 ( \35279 , \35276 , \35277 , \35278 );
and \g455031/U$2 ( \35280 , \8313 , RIe1e5e98_3993);
and \g455031/U$3 ( \35281 , RIe1e8b98_4025, \8323 );
nor \g455031/U$1 ( \35282 , \35280 , \35281 );
not \g450172/U$3 ( \35283 , \35282 );
not \g450172/U$4 ( \35284 , \8328 );
and \g450172/U$2 ( \35285 , \35283 , \35284 );
and \g450172/U$5 ( \35286 , \8359 , RIe1d2398_3769);
nor \g450172/U$1 ( \35287 , \35285 , \35286 );
and \g452810/U$2 ( \35288 , \8404 , RIe1e3198_3961);
and \g452810/U$3 ( \35289 , RIe1eb898_4057, \8351 );
nor \g452810/U$1 ( \35290 , \35288 , \35289 );
and \g452811/U$2 ( \35291 , \8378 , RIe1d7d98_3833);
and \g452811/U$3 ( \35292 , RIe1e0498_3929, \8417 );
nor \g452811/U$1 ( \35293 , \35291 , \35292 );
nand \g447806/U$1 ( \35294 , \35279 , \35287 , \35290 , \35293 );
and \g444726/U$3 ( \35295 , \8478 , \35294 );
nor \g444726/U$1 ( \35296 , \35275 , \35295 );
and \g446991/U$2 ( \35297 , \8775 , RIe1c9c98_3673);
and \g446991/U$3 ( \35298 , RIe1cc998_3705, \8777 );
nor \g446991/U$1 ( \35299 , \35297 , \35298 );
and \g446990/U$2 ( \35300 , \8780 , RIe1c4298_3609);
and \g446990/U$3 ( \35301 , RIe1c6f98_3641, \8782 );
nor \g446990/U$1 ( \35302 , \35300 , \35301 );
and \g446992/U$2 ( \35303 , \8785 , RIe1be898_3545);
and \g446992/U$3 ( \35304 , RIe1c1598_3577, \8787 );
nor \g446992/U$1 ( \35305 , \35303 , \35304 );
nand \g444634/U$1 ( \35306 , \35296 , \35299 , \35302 , \35305 );
and \g452789/U$2 ( \35307 , \8414 , RIfc8ada0_6602);
and \g452789/U$3 ( \35308 , RIfc59b88_6043, \8407 );
nor \g452789/U$1 ( \35309 , \35307 , \35308 );
and \g446210/U$2 ( \35310 , RIfcdb890_7520, \8417 );
and \g446210/U$3 ( \35311 , RIe175c38_2717, \8404 );
and \g449153/U$2 ( \35312 , RIfc57428_6015, \8319 );
and \g449153/U$3 ( \35313 , \8324 , RIfc8a968_6599);
and \g449153/U$4 ( \35314 , RIfc59480_6038, \8330 );
nor \g449153/U$1 ( \35315 , \35312 , \35313 , \35314 );
and \g452796/U$2 ( \35316 , \8335 , RIfc56d20_6010);
and \g452796/U$3 ( \35317 , RIfcc62d8_7277, \8340 );
nor \g452796/U$1 ( \35318 , \35316 , \35317 );
and \g455266/U$2 ( \35319 , \8313 , RIfc58aa8_6031);
and \g455266/U$3 ( \35320 , RIfc57158_6013, \8323 );
nor \g455266/U$1 ( \35321 , \35319 , \35320 );
not \g450168/U$3 ( \35322 , \35321 );
not \g450168/U$4 ( \35323 , \8347 );
and \g450168/U$2 ( \35324 , \35322 , \35323 );
and \g450168/U$5 ( \35325 , \8351 , RIfcbb748_7155);
nor \g450168/U$1 ( \35326 , \35324 , \35325 );
and \g452795/U$2 ( \35327 , \8356 , RIe173910_2692);
and \g452795/U$3 ( \35328 , RIfc57c98_6021, \8359 );
nor \g452795/U$1 ( \35329 , \35327 , \35328 );
nand \g447804/U$1 ( \35330 , \35315 , \35318 , \35326 , \35329 );
nor \g446210/U$1 ( \35331 , \35310 , \35311 , \35330 );
and \g452791/U$2 ( \35332 , \8378 , RIfcb5eb0_7092);
and \g452791/U$3 ( \35333 , RIfcbbce8_7159, \8373 );
nor \g452791/U$1 ( \35334 , \35332 , \35333 );
nand \g445629/U$1 ( \35335 , \35309 , \35331 , \35334 );
and \g444696/U$2 ( \35336 , \35335 , \9700 );
and \g449150/U$2 ( \35337 , RIe1923d8_3041, \8414 );
and \g449150/U$3 ( \35338 , \8409 , RIe1950d8_3073);
and \g449150/U$4 ( \35339 , RIe186fd8_2913, \8486 );
nor \g449150/U$1 ( \35340 , \35337 , \35338 , \35339 );
and \g455011/U$2 ( \35341 , \8313 , RIfcc2d68_7239);
and \g455011/U$3 ( \35342 , RIe19aad8_3137, \8323 );
nor \g455011/U$1 ( \35343 , \35341 , \35342 );
not \g450164/U$3 ( \35344 , \35343 );
not \g450164/U$4 ( \35345 , \8328 );
and \g450164/U$2 ( \35346 , \35344 , \35345 );
and \g450164/U$5 ( \35347 , \8359 , RIe189cd8_2945);
nor \g450164/U$1 ( \35348 , \35346 , \35347 );
and \g452781/U$2 ( \35349 , \8404 , RIe197dd8_3105);
and \g452781/U$3 ( \35350 , RIe19d7d8_3169, \8351 );
nor \g452781/U$1 ( \35351 , \35349 , \35350 );
and \g452782/U$2 ( \35352 , \8378 , RIe18f6d8_3009);
and \g452782/U$3 ( \35353 , RIfc5c5b8_6073, \8417 );
nor \g452782/U$1 ( \35354 , \35352 , \35353 );
nand \g447801/U$1 ( \35355 , \35340 , \35348 , \35351 , \35354 );
and \g444696/U$3 ( \35356 , \9702 , \35355 );
nor \g444696/U$1 ( \35357 , \35336 , \35356 );
and \g446986/U$2 ( \35358 , \9729 , RIe17bbd8_2785);
and \g446986/U$3 ( \35359 , RIe17e8d8_2817, \9731 );
nor \g446986/U$1 ( \35360 , \35358 , \35359 );
and \g446984/U$2 ( \35361 , \9230 , RIe1842d8_2881);
and \g446984/U$3 ( \35362 , RIf1438d0_5228, \9232 );
nor \g446984/U$1 ( \35363 , \35361 , \35362 );
and \g446985/U$2 ( \35364 , \9734 , RIe1815d8_2849);
and \g446985/U$3 ( \35365 , RIfc5b370_6060, \9736 );
nor \g446985/U$1 ( \35366 , \35364 , \35365 );
nand \g444512/U$1 ( \35367 , \35357 , \35360 , \35363 , \35366 );
and \g446203/U$2 ( \35368 , RIe202638_4317, \8373 );
and \g446203/U$3 ( \35369 , RIfcba398_7141, \8378 );
and \g449143/U$2 ( \35370 , RIe1fcda0_4254, \8523 );
and \g449143/U$3 ( \35371 , \8486 , RIfcba0c8_7139);
and \g449143/U$4 ( \35372 , RIfc4bec0_5886, \8383 );
nor \g449143/U$1 ( \35373 , \35370 , \35371 , \35372 );
and \g452755/U$2 ( \35374 , \8335 , RIfc4c5c8_5891);
and \g452755/U$3 ( \35375 , RIfc53d50_5976, \8340 );
nor \g452755/U$1 ( \35376 , \35374 , \35375 );
and \g455336/U$2 ( \35377 , \8313 , RIfc537b0_5972);
and \g455336/U$3 ( \35378 , RIfc9b768_6791, \8323 );
nor \g455336/U$1 ( \35379 , \35377 , \35378 );
not \g455335/U$1 ( \35380 , \35379 );
and \g450156/U$2 ( \35381 , \35380 , \8316 );
and \g450156/U$3 ( \35382 , RIfc88d48_6579, \8351 );
nor \g450156/U$1 ( \35383 , \35381 , \35382 );
and \g452754/U$2 ( \35384 , \8356 , RIe1fbb58_4241);
and \g452754/U$3 ( \35385 , RIfcd4270_7436, \8359 );
nor \g452754/U$1 ( \35386 , \35384 , \35385 );
nand \g448204/U$1 ( \35387 , \35373 , \35376 , \35383 , \35386 );
nor \g446203/U$1 ( \35388 , \35368 , \35369 , \35387 );
and \g452750/U$2 ( \35389 , \8404 , RIe200b80_4298);
and \g452750/U$3 ( \35390 , RIfc4c190_5888, \8409 );
nor \g452750/U$1 ( \35391 , \35389 , \35390 );
and \g452747/U$2 ( \35392 , \8414 , RIfc4c2f8_5889);
and \g452747/U$3 ( \35393 , RIfc88910_6576, \8417 );
nor \g452747/U$1 ( \35394 , \35392 , \35393 );
and \g445298/U$2 ( \35395 , \35388 , \35391 , \35394 );
nor \g445298/U$1 ( \35396 , \35395 , \8422 );
and \g446206/U$2 ( \35397 , RIf169148_5655, \8531 );
and \g446206/U$3 ( \35398 , RIe207930_4376, \8335 );
and \g449145/U$2 ( \35399 , RIe218730_4568, \8414 );
and \g449145/U$3 ( \35400 , \8407 , RIe21e130_4632);
and \g449145/U$4 ( \35401 , RIe212d30_4504, \8488 );
nor \g449145/U$1 ( \35402 , \35399 , \35400 , \35401 );
and \g455318/U$2 ( \35403 , \8313 , RIfc82970_6508);
and \g455318/U$3 ( \35404 , RIe223b30_4696, \8323 );
nor \g455318/U$1 ( \35405 , \35403 , \35404 );
not \g450160/U$3 ( \35406 , \35405 );
not \g450160/U$4 ( \35407 , \8328 );
and \g450160/U$2 ( \35408 , \35406 , \35407 );
and \g450160/U$5 ( \35409 , \8359 , RIfc3fad0_5750);
nor \g450160/U$1 ( \35410 , \35408 , \35409 );
and \g452769/U$2 ( \35411 , \8404 , RIe220e30_4664);
and \g452769/U$3 ( \35412 , RIfc408e0_5760, \8351 );
nor \g452769/U$1 ( \35413 , \35411 , \35412 );
and \g452770/U$2 ( \35414 , \8378 , RIe215a30_4536);
and \g452770/U$3 ( \35415 , RIfcecc30_7716, \8417 );
nor \g452770/U$1 ( \35416 , \35414 , \35415 );
nand \g447798/U$1 ( \35417 , \35402 , \35410 , \35413 , \35416 );
nor \g446206/U$1 ( \35418 , \35397 , \35398 , \35417 );
and \g452762/U$2 ( \35419 , \8356 , RIe210030_4472);
and \g452762/U$3 ( \35420 , RIfc545c0_5982, \8340 );
nor \g452762/U$1 ( \35421 , \35419 , \35420 );
and \g452764/U$2 ( \35422 , \8319 , RIe20a630_4408);
and \g452764/U$3 ( \35423 , RIe20d330_4440, \8324 );
nor \g452764/U$1 ( \35424 , \35422 , \35423 );
and \g445300/U$2 ( \35425 , \35418 , \35421 , \35424 );
nor \g445300/U$1 ( \35426 , \35425 , \8368 );
or \g444371/U$1 ( \35427 , \35306 , \35367 , \35396 , \35426 );
and \g446198/U$2 ( \35428 , RIe18c9d8_2977, \8417 );
and \g446198/U$3 ( \35429 , RIe1a04d8_3201, \8404 );
and \g449135/U$2 ( \35430 , RIe1aea10_3364, \8319 );
and \g449135/U$3 ( \35431 , \8326 , RIe1bbb98_3513);
and \g449135/U$4 ( \35432 , RIe1a5ed8_3265, \8330 );
nor \g449135/U$1 ( \35433 , \35430 , \35431 , \35432 );
and \g452727/U$2 ( \35434 , \8335 , RIe171048_2663);
and \g452727/U$3 ( \35435 , RIe1d5098_3801, \8340 );
nor \g452727/U$1 ( \35436 , \35434 , \35435 );
and \g455174/U$2 ( \35437 , \8313 , RIe1f8048_4199);
and \g455174/U$3 ( \35438 , RIe1fec90_4276, \8323 );
nor \g455174/U$1 ( \35439 , \35437 , \35438 );
not \g450149/U$3 ( \35440 , \35439 );
not \g450149/U$4 ( \35441 , \8347 );
and \g450149/U$2 ( \35442 , \35440 , \35441 );
and \g450149/U$5 ( \35443 , \8351 , RIe1a8bd8_3297);
nor \g450149/U$1 ( \35444 , \35442 , \35443 );
and \g452726/U$2 ( \35445 , \8356 , RIe1f0b90_4116);
and \g452726/U$3 ( \35446 , RIe204c30_4344, \8359 );
nor \g452726/U$1 ( \35447 , \35445 , \35446 );
nand \g447792/U$1 ( \35448 , \35433 , \35436 , \35444 , \35447 );
nor \g446198/U$1 ( \35449 , \35428 , \35429 , \35448 );
and \g452723/U$2 ( \35450 , \8378 , RIe21b430_4600);
and \g452723/U$3 ( \35451 , RIe1a31d8_3233, \8373 );
nor \g452723/U$1 ( \35452 , \35450 , \35451 );
and \g452720/U$2 ( \35453 , \8412 , RIe226830_4728);
and \g452720/U$3 ( \35454 , RIe178ed8_2753, \8407 );
nor \g452720/U$1 ( \35455 , \35453 , \35454 );
and \g445292/U$2 ( \35456 , \35449 , \35452 , \35455 );
nor \g445292/U$1 ( \35457 , \35456 , \8651 );
and \g446200/U$2 ( \35458 , RIfebe890_8288, \8356 );
and \g446200/U$3 ( \35459 , RIfc9cde8_6807, \8340 );
and \g449138/U$2 ( \35460 , RIfebe5c0_8286, \8414 );
and \g449138/U$3 ( \35461 , \8407 , RIf149ca8_5299);
and \g449138/U$4 ( \35462 , RIfce4f08_7627, \8486 );
nor \g449138/U$1 ( \35463 , \35460 , \35461 , \35462 );
and \g455338/U$2 ( \35464 , \8313 , RIe1b92d0_3484);
and \g455338/U$3 ( \35465 , RIf14ba30_5320, \8323 );
nor \g455338/U$1 ( \35466 , \35464 , \35465 );
not \g450152/U$3 ( \35467 , \35466 );
not \g450152/U$4 ( \35468 , \8328 );
and \g450152/U$2 ( \35469 , \35467 , \35468 );
and \g450152/U$5 ( \35470 , \8359 , RIfc50510_5936);
nor \g450152/U$1 ( \35471 , \35469 , \35470 );
and \g452739/U$2 ( \35472 , \8404 , RIe1b7278_3461);
and \g452739/U$3 ( \35473 , RIf14cc78_5333, \8351 );
nor \g452739/U$1 ( \35474 , \35472 , \35473 );
and \g452740/U$2 ( \35475 , \8378 , RIfe807c0_7806);
and \g452740/U$3 ( \35476 , RIf14a7e8_5307, \8417 );
nor \g452740/U$1 ( \35477 , \35475 , \35476 );
nand \g447794/U$1 ( \35478 , \35463 , \35471 , \35474 , \35477 );
nor \g446200/U$1 ( \35479 , \35458 , \35459 , \35478 );
and \g452735/U$2 ( \35480 , \8335 , RIfebe728_8287);
and \g452735/U$3 ( \35481 , RIfe80a90_7808, \8523 );
nor \g452735/U$1 ( \35482 , \35480 , \35481 );
and \g452733/U$2 ( \35483 , \8317 , RIfe80928_7807);
and \g452733/U$3 ( \35484 , RIfc87560_6562, \8326 );
nor \g452733/U$1 ( \35485 , \35483 , \35484 );
and \g445294/U$2 ( \35486 , \35479 , \35482 , \35485 );
nor \g445294/U$1 ( \35487 , \35486 , \8481 );
or \g444172/U$1 ( \35488 , \35427 , \35457 , \35487 );
_DC \g5c24/U$1 ( \35489 , \35488 , \8654 );
and \g452998/U$2 ( \35490 , \16380 , RIdeba2a8_582);
and \g452998/U$3 ( \35491 , RIdec29a8_678, \16321 );
nor \g452998/U$1 ( \35492 , \35490 , \35491 );
and \g446256/U$2 ( \35493 , RIdec56a8_710, \16328 );
and \g446256/U$3 ( \35494 , RIdebfca8_646, \16377 );
and \g449211/U$2 ( \35495 , RIdeaaab0_422, \16398 );
and \g449211/U$3 ( \35496 , \16341 , RIfc6a118_6229);
and \g449211/U$4 ( \35497 , RIdebcfa8_614, \16485 );
nor \g449211/U$1 ( \35498 , \35495 , \35496 , \35497 );
and \g455154/U$2 ( \35499 , \16317 , RIdeb1ba8_486);
and \g455154/U$3 ( \35500 , RIfc4fe08_5931, \16325 );
nor \g455154/U$1 ( \35501 , \35499 , \35500 );
not \g450227/U$3 ( \35502 , \35501 );
not \g450227/U$4 ( \35503 , \16351 );
and \g450227/U$2 ( \35504 , \35502 , \35503 );
and \g450227/U$5 ( \35505 , \16356 , RIee1f540_4815);
nor \g450227/U$1 ( \35506 , \35504 , \35505 );
and \g453004/U$2 ( \35507 , \16361 , RIde9d8b0_358);
and \g453004/U$3 ( \35508 , RIdea41b0_390, \16364 );
nor \g453004/U$1 ( \35509 , \35507 , \35508 );
and \g453003/U$2 ( \35510 , \16368 , RIdeaeea8_454);
and \g453003/U$3 ( \35511 , RIfc6b630_6244, \16371 );
nor \g453003/U$1 ( \35512 , \35510 , \35511 );
nand \g447834/U$1 ( \35513 , \35498 , \35506 , \35509 , \35512 );
nor \g446256/U$1 ( \35514 , \35493 , \35494 , \35513 );
and \g453000/U$2 ( \35515 , \16334 , RIdeb75a8_550);
and \g453000/U$3 ( \35516 , RIfc54020_5978, \16313 );
nor \g453000/U$1 ( \35517 , \35515 , \35516 );
nand \g445640/U$1 ( \35518 , \35492 , \35514 , \35517 );
and \g444735/U$2 ( \35519 , \35518 , \17938 );
and \g449208/U$2 ( \35520 , RIfc687c8_6211, \16321 );
and \g449208/U$3 ( \35521 , \16326 , RIfcde2c0_7550);
and \g449208/U$4 ( \35522 , RIdf335e0_1961, \16398 );
nor \g449208/U$1 ( \35523 , \35520 , \35521 , \35522 );
and \g454876/U$2 ( \35524 , \16317 , RIdf3ef80_2093);
and \g454876/U$3 ( \35525 , RIe141078_2117, \16325 );
nor \g454876/U$1 ( \35526 , \35524 , \35525 );
not \g450224/U$3 ( \35527 , \35526 );
not \g450224/U$4 ( \35528 , \16330 );
and \g450224/U$2 ( \35529 , \35527 , \35528 );
and \g450224/U$5 ( \35530 , \16341 , RIdf35a70_1987);
nor \g450224/U$1 ( \35531 , \35529 , \35530 );
and \g452993/U$2 ( \35532 , \16377 , RIfcb1590_7040);
and \g452993/U$3 ( \35533 , RIfca9160_6946, \16313 );
nor \g452993/U$1 ( \35534 , \35532 , \35533 );
and \g452994/U$2 ( \35535 , \16334 , RIfebeb60_8290);
and \g452994/U$3 ( \35536 , RIdf3cdc0_2069, \16380 );
nor \g452994/U$1 ( \35537 , \35535 , \35536 );
nand \g447394/U$1 ( \35538 , \35523 , \35531 , \35534 , \35537 );
and \g444735/U$3 ( \35539 , \16394 , \35538 );
nor \g444735/U$1 ( \35540 , \35519 , \35539 );
and \g447022/U$2 ( \35541 , \16419 , RIdf2f3c8_1914);
and \g447022/U$3 ( \35542 , RIdf31420_1937, \16422 );
nor \g447022/U$1 ( \35543 , \35541 , \35542 );
and \g447020/U$2 ( \35544 , \16429 , RIee2fad0_5001);
and \g447020/U$3 ( \35545 , RIfc64448_6163, \16434 );
nor \g447020/U$1 ( \35546 , \35544 , \35545 );
and \g447021/U$2 ( \35547 , \16438 , RIfc676e8_6199);
and \g447021/U$3 ( \35548 , RIfca7978_6929, \16441 );
nor \g447021/U$1 ( \35549 , \35547 , \35548 );
nand \g444519/U$1 ( \35550 , \35540 , \35543 , \35546 , \35549 );
and \g449214/U$2 ( \35551 , RIdf09178_1480, \16344 );
and \g449214/U$3 ( \35552 , \16356 , RIdf0be78_1512);
and \g449214/U$4 ( \35553 , RIdeefc78_1192, \16398 );
nor \g449214/U$1 ( \35554 , \35551 , \35552 , \35553 );
and \g455166/U$2 ( \35555 , \16317 , RIdf14578_1608);
and \g455166/U$3 ( \35556 , RIdf17278_1640, \16325 );
nor \g455166/U$1 ( \35557 , \35555 , \35556 );
not \g450229/U$3 ( \35558 , \35557 );
not \g450229/U$4 ( \35559 , \16311 );
and \g450229/U$2 ( \35560 , \35558 , \35559 );
and \g450229/U$5 ( \35561 , \16341 , RIdef2978_1224);
nor \g450229/U$1 ( \35562 , \35560 , \35561 );
and \g453010/U$2 ( \35563 , \16377 , RIdf0eb78_1544);
and \g453010/U$3 ( \35564 , RIdf11878_1576, \16313 );
nor \g453010/U$1 ( \35565 , \35563 , \35564 );
and \g453012/U$2 ( \35566 , \16334 , RIdf03778_1416);
and \g453012/U$3 ( \35567 , RIdf06478_1448, \16380 );
nor \g453012/U$1 ( \35568 , \35566 , \35567 );
nand \g447395/U$1 ( \35569 , \35554 , \35562 , \35565 , \35568 );
and \g444717/U$2 ( \35570 , \35569 , \16750 );
and \g446259/U$2 ( \35571 , RIfccef78_7377, \16328 );
and \g446259/U$3 ( \35572 , RIfc61fb8_6137, \16377 );
and \g449218/U$2 ( \35573 , RIfcafc40_7022, \16427 );
and \g449218/U$3 ( \35574 , \16432 , RIfc44300_5798);
and \g449218/U$4 ( \35575 , RIdf281e0_1833, \16485 );
nor \g449218/U$1 ( \35576 , \35573 , \35574 , \35575 );
and \g454675/U$2 ( \35577 , \16317 , RIdf1fae0_1737);
and \g454675/U$3 ( \35578 , RIdf219d0_1759, \16325 );
nor \g454675/U$1 ( \35579 , \35577 , \35578 );
not \g454674/U$1 ( \35580 , \35579 );
and \g450233/U$2 ( \35581 , \35580 , \16336 );
and \g450233/U$3 ( \35582 , RIfe81b70_7820, \16356 );
nor \g450233/U$1 ( \35583 , \35581 , \35582 );
and \g453023/U$2 ( \35584 , \16361 , RIdf19438_1664);
and \g453023/U$3 ( \35585 , RIdf1b1c0_1685, \16364 );
nor \g453023/U$1 ( \35586 , \35584 , \35585 );
and \g453022/U$2 ( \35587 , \16368 , RIfcaac18_6965);
and \g453022/U$3 ( \35588 , RIdf22ee8_1774, \16371 );
nor \g453022/U$1 ( \35589 , \35587 , \35588 );
nand \g448095/U$1 ( \35590 , \35576 , \35583 , \35586 , \35589 );
nor \g446259/U$1 ( \35591 , \35571 , \35572 , \35590 );
and \g453018/U$2 ( \35592 , \16334 , RIdf249a0_1793);
and \g453018/U$3 ( \35593 , RIfc62558_6141, \16313 );
nor \g453018/U$1 ( \35594 , \35592 , \35593 );
and \g453017/U$2 ( \35595 , \16380 , RIfe81cd8_7821);
and \g453017/U$3 ( \35596 , RIfca6fa0_6922, \16321 );
nor \g453017/U$1 ( \35597 , \35595 , \35596 );
and \g445335/U$2 ( \35598 , \35591 , \35594 , \35597 );
nor \g445335/U$1 ( \35599 , \35598 , \16480 );
nor \g444717/U$1 ( \35600 , \35570 , \35599 );
and \g447032/U$2 ( \35601 , \19208 , RIdeea278_1128);
and \g447032/U$3 ( \35602 , RIdef8378_1288, \19210 );
nor \g447032/U$1 ( \35603 , \35601 , \35602 );
and \g447033/U$2 ( \35604 , \19213 , RIdeecf78_1160);
and \g447033/U$3 ( \35605 , RIdef5678_1256, \19215 );
nor \g447033/U$1 ( \35606 , \35604 , \35605 );
and \g447031/U$2 ( \35607 , \19218 , RIdefb078_1320);
and \g447031/U$3 ( \35608 , RIdefdd78_1352, \19220 );
nor \g447031/U$1 ( \35609 , \35607 , \35608 );
nand \g444639/U$1 ( \35610 , \35600 , \35603 , \35606 , \35609 );
and \g446249/U$2 ( \35611 , RIfc611a8_6127, \16328 );
and \g446249/U$3 ( \35612 , RIfca6b68_6919, \16377 );
and \g449201/U$2 ( \35613 , RIfc738f8_6337, \16427 );
and \g449201/U$3 ( \35614 , \16432 , RIfc626c0_6142);
and \g449201/U$4 ( \35615 , RIdee2dc0_1045, \16485 );
nor \g449201/U$1 ( \35616 , \35613 , \35614 , \35615 );
and \g454916/U$2 ( \35617 , \16317 , RIded7588_914);
and \g454916/U$3 ( \35618 , RIded9a18_940, \16325 );
nor \g454916/U$1 ( \35619 , \35617 , \35618 );
not \g454915/U$1 ( \35620 , \35619 );
and \g450217/U$2 ( \35621 , \35620 , \16336 );
and \g450217/U$3 ( \35622 , RIdee4b48_1066, \16356 );
nor \g450217/U$1 ( \35623 , \35621 , \35622 );
and \g452968/U$2 ( \35624 , \16361 , RIded30a0_865);
and \g452968/U$3 ( \35625 , RIded5698_892, \16364 );
nor \g452968/U$1 ( \35626 , \35624 , \35625 );
and \g452967/U$2 ( \35627 , \16368 , RIee21430_4837);
and \g452967/U$3 ( \35628 , RIfcb31b0_7060, \16371 );
nor \g452967/U$1 ( \35629 , \35627 , \35628 );
nand \g448094/U$1 ( \35630 , \35616 , \35623 , \35626 , \35629 );
nor \g446249/U$1 ( \35631 , \35611 , \35612 , \35630 );
and \g452963/U$2 ( \35632 , \16334 , RIdedeba8_998);
and \g452963/U$3 ( \35633 , RIfca65c8_6915, \16313 );
nor \g452963/U$1 ( \35634 , \35632 , \35633 );
and \g452962/U$2 ( \35635 , \16380 , RIdee0c00_1021);
and \g452962/U$3 ( \35636 , RIfc61a18_6133, \16319 );
nor \g452962/U$1 ( \35637 , \35635 , \35636 );
and \g445326/U$2 ( \35638 , \35631 , \35634 , \35637 );
nor \g445326/U$1 ( \35639 , \35638 , \16909 );
and \g446251/U$2 ( \35640 , RIe143aa8_2147, \16448 );
and \g446251/U$3 ( \35641 , RIde7cef8_199, \16361 );
and \g449204/U$2 ( \35642 , RIde96fb0_326, \16485 );
and \g449204/U$3 ( \35643 , \16356 , RIdeb48a8_518);
and \g449204/U$4 ( \35644 , RIdee7578_1096, \16398 );
nor \g449204/U$1 ( \35645 , \35642 , \35643 , \35644 );
and \g455137/U$2 ( \35646 , \16317 , RIdecdda8_806);
and \g455137/U$3 ( \35647 , RIded0aa8_838, \16325 );
nor \g455137/U$1 ( \35648 , \35646 , \35647 );
not \g450220/U$3 ( \35649 , \35648 );
not \g450220/U$4 ( \35650 , \16311 );
and \g450220/U$2 ( \35651 , \35649 , \35650 );
and \g450220/U$5 ( \35652 , \16341 , RIdf00a78_1384);
nor \g450220/U$1 ( \35653 , \35651 , \35652 );
and \g452980/U$2 ( \35654 , \16377 , RIdec83a8_742);
and \g452980/U$3 ( \35655 , RIdecb0a8_774, \16313 );
nor \g452980/U$1 ( \35656 , \35654 , \35655 );
and \g452981/U$2 ( \35657 , \16334 , RIe15a2a8_2403);
and \g452981/U$3 ( \35658 , RIe16e4b0_2632, \16380 );
nor \g452981/U$1 ( \35659 , \35657 , \35658 );
nand \g447393/U$1 ( \35660 , \35645 , \35653 , \35656 , \35659 );
nor \g446251/U$1 ( \35661 , \35640 , \35641 , \35660 );
and \g452976/U$2 ( \35662 , \16364 , RIdedc2e0_969);
and \g452976/U$3 ( \35663 , RIdf1d380_1709, \16368 );
nor \g452976/U$1 ( \35664 , \35662 , \35663 );
and \g452975/U$2 ( \35665 , \16371 , RIdf2cb00_1885);
and \g452975/U$3 ( \35666 , RIdf384a0_2017, \16427 );
nor \g452975/U$1 ( \35667 , \35665 , \35666 );
and \g445330/U$2 ( \35668 , \35661 , \35664 , \35667 );
nor \g445330/U$1 ( \35669 , \35668 , \16586 );
or \g444319/U$1 ( \35670 , \35550 , \35610 , \35639 , \35669 );
and \g446243/U$2 ( \35671 , RIee1be68_4776, \16321 );
and \g446243/U$3 ( \35672 , RIfc653c0_6174, \16313 );
and \g449193/U$2 ( \35673 , RIe16b918_2601, \16398 );
and \g449193/U$3 ( \35674 , \16341 , RIfc6b360_6242);
and \g449193/U$4 ( \35675 , RIde8df50_282, \16485 );
nor \g449193/U$1 ( \35676 , \35673 , \35674 , \35675 );
and \g454971/U$2 ( \35677 , \16317 , RIfca76a8_6927);
and \g454971/U$3 ( \35678 , RIde81db8_223, \16325 );
nor \g454971/U$1 ( \35679 , \35677 , \35678 );
not \g450210/U$3 ( \35680 , \35679 );
not \g450210/U$4 ( \35681 , \16351 );
and \g450210/U$2 ( \35682 , \35680 , \35681 );
and \g450210/U$5 ( \35683 , \16356 , RIde91718_299);
nor \g450210/U$1 ( \35684 , \35682 , \35683 );
and \g452943/U$2 ( \35685 , \16361 , RIe167f70_2560);
and \g452943/U$3 ( \35686 , RIe169cf8_2581, \16364 );
nor \g452943/U$1 ( \35687 , \35685 , \35686 );
and \g452942/U$2 ( \35688 , \16368 , RIfc4ce38_5897);
and \g452942/U$3 ( \35689 , RIfcca4f0_7324, \16371 );
nor \g452942/U$1 ( \35690 , \35688 , \35689 );
nand \g447824/U$1 ( \35691 , \35676 , \35684 , \35687 , \35690 );
nor \g446243/U$1 ( \35692 , \35671 , \35672 , \35691 );
and \g452939/U$2 ( \35693 , \16377 , RIee1ac20_4763);
and \g452939/U$3 ( \35694 , RIde89db0_262, \16380 );
nor \g452939/U$1 ( \35695 , \35693 , \35694 );
and \g452937/U$2 ( \35696 , \16334 , RIde85c10_242);
and \g452937/U$3 ( \35697 , RIfc69ce0_6226, \16328 );
nor \g452937/U$1 ( \35698 , \35696 , \35697 );
and \g445320/U$2 ( \35699 , \35692 , \35695 , \35698 );
nor \g445320/U$1 ( \35700 , \35699 , \16649 );
and \g446246/U$2 ( \35701 , RIee35908_5068, \16448 );
and \g446246/U$3 ( \35702 , RIe1467a8_2179, \16361 );
and \g449197/U$2 ( \35703 , RIe15cfa8_2435, \16485 );
and \g449197/U$3 ( \35704 , \16354 , RIfce93f0_7676);
and \g449197/U$4 ( \35705 , RIe14c1a8_2243, \16398 );
nor \g449197/U$1 ( \35706 , \35703 , \35704 , \35705 );
and \g455126/U$2 ( \35707 , \16317 , RIe1629a8_2499);
and \g455126/U$3 ( \35708 , RIe1656a8_2531, \16325 );
nor \g455126/U$1 ( \35709 , \35707 , \35708 );
not \g450213/U$3 ( \35710 , \35709 );
not \g450213/U$4 ( \35711 , \16311 );
and \g450213/U$2 ( \35712 , \35710 , \35711 );
and \g450213/U$5 ( \35713 , \16341 , RIfce32e8_7607);
nor \g450213/U$1 ( \35714 , \35712 , \35713 );
and \g452954/U$2 ( \35715 , \16377 , RIe15fca8_2467);
and \g452954/U$3 ( \35716 , RIee37690_5089, \16313 );
nor \g452954/U$1 ( \35717 , \35715 , \35716 );
and \g452955/U$2 ( \35718 , \16334 , RIe1548a8_2339);
and \g452955/U$3 ( \35719 , RIe1575a8_2371, \16380 );
nor \g452955/U$1 ( \35720 , \35718 , \35719 );
nand \g447392/U$1 ( \35721 , \35706 , \35714 , \35717 , \35720 );
nor \g446246/U$1 ( \35722 , \35701 , \35702 , \35721 );
and \g452951/U$2 ( \35723 , \16364 , RIe1494a8_2211);
and \g452951/U$3 ( \35724 , RIe14eea8_2275, \16368 );
nor \g452951/U$1 ( \35725 , \35723 , \35724 );
and \g452949/U$2 ( \35726 , \16371 , RIee34f30_5061);
and \g452949/U$3 ( \35727 , RIe151ba8_2307, \16427 );
nor \g452949/U$1 ( \35728 , \35726 , \35727 );
and \g445322/U$2 ( \35729 , \35722 , \35725 , \35728 );
nor \g445322/U$1 ( \35730 , \35729 , \16389 );
or \g444218/U$1 ( \35731 , \35670 , \35700 , \35730 );
_DC \g5ca9/U$1 ( \35732 , \35731 , \16652 );
and \g453098/U$2 ( \35733 , \8412 , RIfca81e8_6935);
and \g453098/U$3 ( \35734 , RIf13f3e8_5179, \8407 );
nor \g453098/U$1 ( \35735 , \35733 , \35734 );
and \g446275/U$2 ( \35736 , RIfccabf8_7329, \8417 );
and \g446275/U$3 ( \35737 , RIfe81738_7817, \8404 );
and \g449237/U$2 ( \35738 , RIfcdde88_7547, \8523 );
and \g449237/U$3 ( \35739 , \8488 , RIfc6ed08_6283);
and \g449237/U$4 ( \35740 , RIf141008_5199, \8383 );
nor \g449237/U$1 ( \35741 , \35738 , \35739 , \35740 );
and \g453105/U$2 ( \35742 , \8335 , RIfcacdd8_6989);
and \g453105/U$3 ( \35743 , RIfc66338_6185, \8340 );
nor \g453105/U$1 ( \35744 , \35742 , \35743 );
and \g454706/U$2 ( \35745 , \8313 , RIfc664a0_6186);
and \g454706/U$3 ( \35746 , RIfc6eba0_6282, \8323 );
nor \g454706/U$1 ( \35747 , \35745 , \35746 );
not \g454705/U$1 ( \35748 , \35747 );
and \g450252/U$2 ( \35749 , \35748 , \8316 );
and \g450252/U$3 ( \35750 , RIfc64f88_6171, \8351 );
nor \g450252/U$1 ( \35751 , \35749 , \35750 );
and \g453103/U$2 ( \35752 , \8356 , RIe173a78_2693);
and \g453103/U$3 ( \35753 , RIfc66068_6183, \8359 );
nor \g453103/U$1 ( \35754 , \35752 , \35753 );
nand \g448215/U$1 ( \35755 , \35741 , \35744 , \35751 , \35754 );
nor \g446275/U$1 ( \35756 , \35736 , \35737 , \35755 );
and \g453100/U$2 ( \35757 , \8378 , RIee3d630_5157);
and \g453100/U$3 ( \35758 , RIe177150_2732, \8373 );
nor \g453100/U$1 ( \35759 , \35757 , \35758 );
nand \g445644/U$1 ( \35760 , \35735 , \35756 , \35759 );
and \g444746/U$2 ( \35761 , \35760 , \9700 );
and \g449234/U$2 ( \35762 , RIf143a38_5229, \8531 );
and \g449234/U$3 ( \35763 , \8486 , RIe187140_2914);
and \g449234/U$4 ( \35764 , RIe19ac40_3138, \8383 );
nor \g449234/U$1 ( \35765 , \35762 , \35763 , \35764 );
and \g453094/U$2 ( \35766 , \8335 , RIe17bd40_2786);
and \g453094/U$3 ( \35767 , RIfc6f140_6286, \8340 );
nor \g453094/U$1 ( \35768 , \35766 , \35767 );
and \g455220/U$2 ( \35769 , \8313 , RIe17ea40_2818);
and \g455220/U$3 ( \35770 , RIe181740_2850, \8323 );
nor \g455220/U$1 ( \35771 , \35769 , \35770 );
not \g455219/U$1 ( \35772 , \35771 );
and \g450249/U$2 ( \35773 , \35772 , \8316 );
and \g450249/U$3 ( \35774 , RIe19d940_3170, \8351 );
nor \g450249/U$1 ( \35775 , \35773 , \35774 );
and \g453092/U$2 ( \35776 , \8356 , RIe184440_2882);
and \g453092/U$3 ( \35777 , RIe189e40_2946, \8359 );
nor \g453092/U$1 ( \35778 , \35776 , \35777 );
nand \g448214/U$1 ( \35779 , \35765 , \35768 , \35775 , \35778 );
and \g444746/U$3 ( \35780 , \9702 , \35779 );
nor \g444746/U$1 ( \35781 , \35761 , \35780 );
and \g447042/U$2 ( \35782 , \11700 , RIe195240_3074);
and \g447042/U$3 ( \35783 , RIf144848_5239, \11702 );
nor \g447042/U$1 ( \35784 , \35782 , \35783 );
and \g447044/U$2 ( \35785 , \9724 , RIe197f40_3106);
and \g447044/U$3 ( \35786 , RIfc64880_6166, \9726 );
nor \g447044/U$1 ( \35787 , \35785 , \35786 );
and \g447043/U$2 ( \35788 , \9170 , RIe18f840_3010);
and \g447043/U$3 ( \35789 , RIe192540_3042, \9172 );
nor \g447043/U$1 ( \35790 , \35788 , \35789 );
nand \g444522/U$1 ( \35791 , \35781 , \35784 , \35787 , \35790 );
and \g453128/U$2 ( \35792 , \8378 , RIe1f5780_4170);
and \g453128/U$3 ( \35793 , RIfcabe60_6978, \8409 );
nor \g453128/U$1 ( \35794 , \35792 , \35793 );
and \g446281/U$2 ( \35795 , RIfc6d3b8_6265, \8373 );
and \g446281/U$3 ( \35796 , RIfc6d0e8_6263, \8414 );
and \g449244/U$2 ( \35797 , RIfc68c00_6214, \8531 );
and \g449244/U$3 ( \35798 , \8488 , RIfc68d68_6215);
and \g449244/U$4 ( \35799 , RIfc6cf80_6262, \8383 );
nor \g449244/U$1 ( \35800 , \35797 , \35798 , \35799 );
and \g453132/U$2 ( \35801 , \8335 , RIe1ee160_4086);
and \g453132/U$3 ( \35802 , RIfc68a98_6213, \8340 );
nor \g453132/U$1 ( \35803 , \35801 , \35802 );
and \g454689/U$2 ( \35804 , \8313 , RIfca9b38_6953);
and \g454689/U$3 ( \35805 , RIfccb8a0_7338, \8323 );
nor \g454689/U$1 ( \35806 , \35804 , \35805 );
not \g454688/U$1 ( \35807 , \35806 );
and \g450259/U$2 ( \35808 , \35807 , \8316 );
and \g450259/U$3 ( \35809 , RIfc587d8_6029, \8351 );
nor \g450259/U$1 ( \35810 , \35808 , \35809 );
and \g453131/U$2 ( \35811 , \8356 , RIe1f3458_4145);
and \g453131/U$3 ( \35812 , RIfc6c5a8_6255, \8359 );
nor \g453131/U$1 ( \35813 , \35811 , \35812 );
nand \g448219/U$1 ( \35814 , \35800 , \35803 , \35810 , \35813 );
nor \g446281/U$1 ( \35815 , \35795 , \35796 , \35814 );
and \g453127/U$2 ( \35816 , \8404 , RIfe815d0_7816);
and \g453127/U$3 ( \35817 , RIfc6d520_6266, \8417 );
nor \g453127/U$1 ( \35818 , \35816 , \35817 );
nand \g445646/U$1 ( \35819 , \35794 , \35815 , \35818 );
and \g444727/U$2 ( \35820 , \35819 , \8752 );
and \g449240/U$2 ( \35821 , RIe1dac00_3866, \8414 );
and \g449240/U$3 ( \35822 , \8407 , RIe1dd900_3898);
and \g449240/U$4 ( \35823 , RIe1cf800_3738, \8488 );
nor \g449240/U$1 ( \35824 , \35821 , \35822 , \35823 );
and \g454695/U$2 ( \35825 , \8313 , RIe1e6000_3994);
and \g454695/U$3 ( \35826 , RIe1e8d00_4026, \8323 );
nor \g454695/U$1 ( \35827 , \35825 , \35826 );
not \g450256/U$3 ( \35828 , \35827 );
not \g450256/U$4 ( \35829 , \8328 );
and \g450256/U$2 ( \35830 , \35828 , \35829 );
and \g450256/U$5 ( \35831 , \8359 , RIe1d2500_3770);
nor \g450256/U$1 ( \35832 , \35830 , \35831 );
and \g453115/U$2 ( \35833 , \8404 , RIe1e3300_3962);
and \g453115/U$3 ( \35834 , RIe1eba00_4058, \8351 );
nor \g453115/U$1 ( \35835 , \35833 , \35834 );
and \g453117/U$2 ( \35836 , \8378 , RIe1d7f00_3834);
and \g453117/U$3 ( \35837 , RIe1e0600_3930, \8417 );
nor \g453117/U$1 ( \35838 , \35836 , \35837 );
nand \g447852/U$1 ( \35839 , \35824 , \35832 , \35835 , \35838 );
and \g444727/U$3 ( \35840 , \8478 , \35839 );
nor \g444727/U$1 ( \35841 , \35820 , \35840 );
and \g447049/U$2 ( \35842 , \8775 , RIe1c9e00_3674);
and \g447049/U$3 ( \35843 , RIe1ccb00_3706, \8777 );
nor \g447049/U$1 ( \35844 , \35842 , \35843 );
and \g447050/U$2 ( \35845 , \8780 , RIe1c4400_3610);
and \g447050/U$3 ( \35846 , RIe1c7100_3642, \8782 );
nor \g447050/U$1 ( \35847 , \35845 , \35846 );
and \g447051/U$2 ( \35848 , \8785 , RIe1bea00_3546);
and \g447051/U$3 ( \35849 , RIe1c1700_3578, \8787 );
nor \g447051/U$1 ( \35850 , \35848 , \35849 );
nand \g444641/U$1 ( \35851 , \35841 , \35844 , \35847 , \35850 );
and \g446269/U$2 ( \35852 , RIe1b0bd0_3388, \8356 );
and \g446269/U$3 ( \35853 , RIfc6ce18_6261, \8340 );
and \g449227/U$2 ( \35854 , RIe1b9438_3485, \8373 );
and \g449227/U$3 ( \35855 , \8383 , RIfcdd348_7539);
and \g449227/U$4 ( \35856 , RIfcab488_6971, \8488 );
nor \g449227/U$1 ( \35857 , \35854 , \35855 , \35856 );
and \g454415/U$2 ( \35858 , \8313 , RIe1b5220_3438);
and \g454415/U$3 ( \35859 , RIfccbb70_7340, \8323 );
nor \g454415/U$1 ( \35860 , \35858 , \35859 );
not \g450242/U$3 ( \35861 , \35860 );
not \g450242/U$4 ( \35862 , \8376 );
and \g450242/U$2 ( \35863 , \35861 , \35862 );
and \g450242/U$5 ( \35864 , \8359 , RIfc6c9e0_6258);
nor \g450242/U$1 ( \35865 , \35863 , \35864 );
and \g453064/U$2 ( \35866 , \8404 , RIe1b73e0_3462);
and \g453064/U$3 ( \35867 , RIfc6bbd0_6248, \8351 );
nor \g453064/U$1 ( \35868 , \35866 , \35867 );
and \g453065/U$2 ( \35869 , \8378 , RIe1b3e70_3424);
and \g453065/U$3 ( \35870 , RIfcab5f0_6972, \8417 );
nor \g453065/U$1 ( \35871 , \35869 , \35870 );
nand \g447845/U$1 ( \35872 , \35857 , \35865 , \35868 , \35871 );
nor \g446269/U$1 ( \35873 , \35852 , \35853 , \35872 );
and \g453061/U$2 ( \35874 , \8335 , RIe1aaf00_3322);
and \g453061/U$3 ( \35875 , RIfea7dc0_8226, \8531 );
nor \g453061/U$1 ( \35876 , \35874 , \35875 );
and \g453060/U$2 ( \35877 , \8319 , RIe1ac580_3338);
and \g453060/U$3 ( \35878 , RIfcabfc8_6979, \8324 );
nor \g453060/U$1 ( \35879 , \35877 , \35878 );
and \g445344/U$2 ( \35880 , \35873 , \35876 , \35879 );
nor \g445344/U$1 ( \35881 , \35880 , \8481 );
and \g446271/U$2 ( \35882 , RIe1f81b0_4200, \8531 );
and \g446271/U$3 ( \35883 , RIe1aeb78_3365, \8319 );
and \g449230/U$2 ( \35884 , RIe1a3340_3234, \8371 );
and \g449230/U$3 ( \35885 , \8330 , RIe1a6040_3266);
and \g449230/U$4 ( \35886 , RIe1fedf8_4277, \8488 );
nor \g449230/U$1 ( \35887 , \35884 , \35885 , \35886 );
and \g454732/U$2 ( \35888 , \8313 , RIe226998_4729);
and \g454732/U$3 ( \35889 , RIe179040_2754, \8323 );
nor \g454732/U$1 ( \35890 , \35888 , \35889 );
not \g450245/U$3 ( \35891 , \35890 );
not \g450245/U$4 ( \35892 , \8376 );
and \g450245/U$2 ( \35893 , \35891 , \35892 );
and \g450245/U$5 ( \35894 , \8359 , RIe204d98_4345);
nor \g450245/U$1 ( \35895 , \35893 , \35894 );
and \g453076/U$2 ( \35896 , \8404 , RIe1a0640_3202);
and \g453076/U$3 ( \35897 , RIe1a8d40_3298, \8351 );
nor \g453076/U$1 ( \35898 , \35896 , \35897 );
and \g453078/U$2 ( \35899 , \8378 , RIe21b598_4601);
and \g453078/U$3 ( \35900 , RIe18cb40_2978, \8417 );
nor \g453078/U$1 ( \35901 , \35899 , \35900 );
nand \g447848/U$1 ( \35902 , \35887 , \35895 , \35898 , \35901 );
nor \g446271/U$1 ( \35903 , \35882 , \35883 , \35902 );
and \g453074/U$2 ( \35904 , \8335 , RIe1711b0_2664);
and \g453074/U$3 ( \35905 , RIe1d5200_3802, \8340 );
nor \g453074/U$1 ( \35906 , \35904 , \35905 );
and \g453073/U$2 ( \35907 , \8326 , RIe1bbd00_3514);
and \g453073/U$3 ( \35908 , RIe1f0cf8_4117, \8356 );
nor \g453073/U$1 ( \35909 , \35907 , \35908 );
and \g445346/U$2 ( \35910 , \35903 , \35906 , \35909 );
nor \g445346/U$1 ( \35911 , \35910 , \8651 );
or \g444326/U$1 ( \35912 , \35791 , \35851 , \35881 , \35911 );
and \g446261/U$2 ( \35913 , RIfc67850_6200, \8531 );
and \g446261/U$3 ( \35914 , RIe20a798_4409, \8317 );
and \g449221/U$2 ( \35915 , RIfc66d10_6192, \8373 );
and \g449221/U$3 ( \35916 , \8383 , RIe223c98_4697);
and \g449221/U$4 ( \35917 , RIe212e98_4505, \8488 );
nor \g449221/U$1 ( \35918 , \35915 , \35916 , \35917 );
and \g454786/U$2 ( \35919 , \8313 , RIe218898_4569);
and \g454786/U$3 ( \35920 , RIe21e298_4633, \8323 );
nor \g454786/U$1 ( \35921 , \35919 , \35920 );
not \g450236/U$3 ( \35922 , \35921 );
not \g450236/U$4 ( \35923 , \8376 );
and \g450236/U$2 ( \35924 , \35922 , \35923 );
and \g450236/U$5 ( \35925 , \8359 , RIfc3fc38_5751);
nor \g450236/U$1 ( \35926 , \35924 , \35925 );
and \g453037/U$2 ( \35927 , \8404 , RIe220f98_4665);
and \g453037/U$3 ( \35928 , RIfe81468_7815, \8351 );
nor \g453037/U$1 ( \35929 , \35927 , \35928 );
and \g453040/U$2 ( \35930 , \8378 , RIe215b98_4537);
and \g453040/U$3 ( \35931 , RIf16b038_5677, \8417 );
nor \g453040/U$1 ( \35932 , \35930 , \35931 );
nand \g447840/U$1 ( \35933 , \35918 , \35926 , \35929 , \35932 );
nor \g446261/U$1 ( \35934 , \35913 , \35914 , \35933 );
and \g453035/U$2 ( \35935 , \8335 , RIe207a98_4377);
and \g453035/U$3 ( \35936 , RIf167f00_5642, \8340 );
nor \g453035/U$1 ( \35937 , \35935 , \35936 );
and \g453034/U$2 ( \35938 , \8326 , RIe20d498_4441);
and \g453034/U$3 ( \35939 , RIe210198_4473, \8356 );
nor \g453034/U$1 ( \35940 , \35938 , \35939 );
and \g445336/U$2 ( \35941 , \35934 , \35937 , \35940 );
nor \g445336/U$1 ( \35942 , \35941 , \8368 );
and \g446264/U$2 ( \35943 , RIfe81300_7814, \8356 );
and \g446264/U$3 ( \35944 , RIfc6dac0_6270, \8340 );
and \g449225/U$2 ( \35945 , RIfea8900_8234, \8371 );
and \g449225/U$3 ( \35946 , \8383 , RIfcac9a0_6986);
and \g449225/U$4 ( \35947 , RIf15e450_5532, \8486 );
nor \g449225/U$1 ( \35948 , \35945 , \35946 , \35947 );
and \g455196/U$2 ( \35949 , \8313 , RIfcac838_6985);
and \g455196/U$3 ( \35950 , RIfccad60_7330, \8323 );
nor \g455196/U$1 ( \35951 , \35949 , \35950 );
not \g450240/U$3 ( \35952 , \35951 );
not \g450240/U$4 ( \35953 , \8376 );
and \g450240/U$2 ( \35954 , \35952 , \35953 );
and \g450240/U$5 ( \35955 , \8359 , RIf160340_5554);
nor \g450240/U$1 ( \35956 , \35954 , \35955 );
and \g453049/U$2 ( \35957 , \8404 , RIfe818a0_7818);
and \g453049/U$3 ( \35958 , RIfcacb08_6987, \8351 );
nor \g453049/U$1 ( \35959 , \35957 , \35958 );
and \g453052/U$2 ( \35960 , \8378 , RIfc67418_6197);
and \g453052/U$3 ( \35961 , RIfca8a58_6941, \8417 );
nor \g453052/U$1 ( \35962 , \35960 , \35961 );
nand \g447842/U$1 ( \35963 , \35948 , \35956 , \35959 , \35962 );
nor \g446264/U$1 ( \35964 , \35943 , \35944 , \35963 );
and \g453046/U$2 ( \35965 , \8335 , RIfc6d7f0_6268);
and \g453046/U$3 ( \35966 , RIfe81a08_7819, \8523 );
nor \g453046/U$1 ( \35967 , \35965 , \35966 );
and \g453045/U$2 ( \35968 , \8317 , RIfc6d958_6269);
and \g453045/U$3 ( \35969 , RIf15ba20_5502, \8326 );
nor \g453045/U$1 ( \35970 , \35968 , \35969 );
and \g445338/U$2 ( \35971 , \35964 , \35967 , \35970 );
nor \g445338/U$1 ( \35972 , \35971 , \8422 );
or \g444246/U$1 ( \35973 , \35912 , \35942 , \35972 );
_DC \g5d2d/U$1 ( \35974 , \35973 , \8654 );
and \g453774/U$2 ( \35975 , \16334 , RIdeded10_999);
and \g453774/U$3 ( \35976 , RIfce6858_7645, \16427 );
nor \g453774/U$1 ( \35977 , \35975 , \35976 );
and \g446417/U$2 ( \35978 , RIdee0d68_1022, \16380 );
and \g446417/U$3 ( \35979 , RIfcdc970_7532, \16368 );
and \g449418/U$2 ( \35980 , RIfeaaac0_8258, \16398 );
and \g449418/U$3 ( \35981 , \16341 , RIded9b80_941);
and \g449418/U$4 ( \35982 , RIdee2f28_1046, \16485 );
nor \g449418/U$1 ( \35983 , \35980 , \35981 , \35982 );
and \g453780/U$2 ( \35984 , \16361 , RIded3208_866);
and \g453780/U$3 ( \35985 , RIded5800_893, \16364 );
nor \g453780/U$1 ( \35986 , \35984 , \35985 );
and \g453778/U$2 ( \35987 , \16377 , RIfce66f0_7644);
and \g453778/U$3 ( \35988 , RIee23e60_4867, \16313 );
nor \g453778/U$1 ( \35989 , \35987 , \35988 );
and \g455098/U$2 ( \35990 , \16317 , RIfca73d8_6925);
and \g455098/U$3 ( \35991 , RIee257b0_4885, \16325 );
nor \g455098/U$1 ( \35992 , \35990 , \35991 );
not \g450439/U$3 ( \35993 , \35992 );
not \g450439/U$4 ( \35994 , \16311 );
and \g450439/U$2 ( \35995 , \35993 , \35994 );
and \g450439/U$5 ( \35996 , \16356 , RIdee4cb0_1067);
nor \g450439/U$1 ( \35997 , \35995 , \35996 );
nand \g447958/U$1 ( \35998 , \35983 , \35986 , \35989 , \35997 );
nor \g446417/U$1 ( \35999 , \35978 , \35979 , \35998 );
and \g453771/U$2 ( \36000 , \16371 , RIfcceca8_7375);
and \g453771/U$3 ( \36001 , RIfcca388_7323, \16448 );
nor \g453771/U$1 ( \36002 , \36000 , \36001 );
nand \g445686/U$1 ( \36003 , \35977 , \35999 , \36002 );
and \g444924/U$2 ( \36004 , \36003 , \16477 );
and \g449414/U$2 ( \36005 , RIde972f8_327, \16344 );
and \g449414/U$3 ( \36006 , \16356 , RIdeb4a10_519);
and \g449414/U$4 ( \36007 , RIdee76e0_1097, \16398 );
nor \g449414/U$1 ( \36008 , \36005 , \36006 , \36007 );
and \g455103/U$2 ( \36009 , \16317 , RIdecdf10_807);
and \g455103/U$3 ( \36010 , RIded0c10_839, \16325 );
nor \g455103/U$1 ( \36011 , \36009 , \36010 );
not \g450434/U$3 ( \36012 , \36011 );
not \g450434/U$4 ( \36013 , \16311 );
and \g450434/U$2 ( \36014 , \36012 , \36013 );
and \g450434/U$5 ( \36015 , \16341 , RIdf00be0_1385);
nor \g450434/U$1 ( \36016 , \36014 , \36015 );
and \g453764/U$2 ( \36017 , \16377 , RIdec8510_743);
and \g453764/U$3 ( \36018 , RIdecb210_775, \16313 );
nor \g453764/U$1 ( \36019 , \36017 , \36018 );
and \g453765/U$2 ( \36020 , \16334 , RIe15a410_2404);
and \g453765/U$3 ( \36021 , RIe16e618_2633, \16380 );
nor \g453765/U$1 ( \36022 , \36020 , \36021 );
nand \g447425/U$1 ( \36023 , \36008 , \36016 , \36019 , \36022 );
and \g444924/U$3 ( \36024 , \16752 , \36023 );
nor \g444924/U$1 ( \36025 , \36004 , \36024 );
and \g447169/U$2 ( \36026 , \16774 , RIde7d240_200);
and \g447169/U$3 ( \36027 , RIdedc448_970, \16776 );
nor \g447169/U$1 ( \36028 , \36026 , \36027 );
and \g447168/U$2 ( \36029 , \16779 , RIdf1d4e8_1710);
and \g447168/U$3 ( \36030 , RIdf2cc68_1886, \16781 );
nor \g447168/U$1 ( \36031 , \36029 , \36030 );
and \g447167/U$2 ( \36032 , \16784 , RIdf38608_2018);
and \g447167/U$3 ( \36033 , RIe143c10_2148, \16786 );
nor \g447167/U$1 ( \36034 , \36032 , \36033 );
nand \g444660/U$1 ( \36035 , \36025 , \36028 , \36031 , \36034 );
and \g453749/U$2 ( \36036 , \16377 , RIdf0ece0_1545);
and \g453749/U$3 ( \36037 , RIdf065e0_1449, \16380 );
nor \g453749/U$1 ( \36038 , \36036 , \36037 );
and \g446413/U$2 ( \36039 , RIdf146e0_1609, \16319 );
and \g446413/U$3 ( \36040 , RIdf119e0_1577, \16313 );
and \g449411/U$2 ( \36041 , RIdefb1e0_1321, \16427 );
and \g449411/U$3 ( \36042 , \16448 , RIdefdee0_1353);
and \g449411/U$4 ( \36043 , RIdf092e0_1481, \16344 );
nor \g449411/U$1 ( \36044 , \36041 , \36042 , \36043 );
and \g455108/U$2 ( \36045 , \16317 , RIdeefde0_1193);
and \g455108/U$3 ( \36046 , RIdef2ae0_1225, \16325 );
nor \g455108/U$1 ( \36047 , \36045 , \36046 );
not \g455107/U$1 ( \36048 , \36047 );
and \g450432/U$2 ( \36049 , \36048 , \16336 );
and \g450432/U$3 ( \36050 , RIdf0bfe0_1513, \16354 );
nor \g450432/U$1 ( \36051 , \36049 , \36050 );
and \g453754/U$2 ( \36052 , \16361 , RIdeea3e0_1129);
and \g453754/U$3 ( \36053 , RIdeed0e0_1161, \16364 );
nor \g453754/U$1 ( \36054 , \36052 , \36053 );
and \g453753/U$2 ( \36055 , \16368 , RIdef57e0_1257);
and \g453753/U$3 ( \36056 , RIdef84e0_1289, \16371 );
nor \g453753/U$1 ( \36057 , \36055 , \36056 );
nand \g448120/U$1 ( \36058 , \36044 , \36051 , \36054 , \36057 );
nor \g446413/U$1 ( \36059 , \36039 , \36040 , \36058 );
and \g453747/U$2 ( \36060 , \16334 , RIdf038e0_1417);
and \g453747/U$3 ( \36061 , RIdf173e0_1641, \16328 );
nor \g453747/U$1 ( \36062 , \36060 , \36061 );
nand \g445683/U$1 ( \36063 , \36038 , \36059 , \36062 );
and \g444805/U$2 ( \36064 , \36063 , \16750 );
and \g449409/U$2 ( \36065 , RIdf28348_1834, \16485 );
and \g449409/U$3 ( \36066 , \16356 , RIdf2a508_1858);
and \g449409/U$4 ( \36067 , RIdf1fc48_1738, \16398 );
nor \g449409/U$1 ( \36068 , \36065 , \36066 , \36067 );
and \g454573/U$2 ( \36069 , \16317 , RIee2a508_4940);
and \g454573/U$3 ( \36070 , RIee2be58_4958, \16325 );
nor \g454573/U$1 ( \36071 , \36069 , \36070 );
not \g450429/U$3 ( \36072 , \36071 );
not \g450429/U$4 ( \36073 , \16311 );
and \g450429/U$2 ( \36074 , \36072 , \36073 );
and \g450429/U$5 ( \36075 , \16341 , RIfcb0078_7025);
nor \g450429/U$1 ( \36076 , \36074 , \36075 );
and \g453743/U$2 ( \36077 , \16377 , RIee27da8_4912);
and \g453743/U$3 ( \36078 , RIee28ff0_4925, \16313 );
nor \g453743/U$1 ( \36079 , \36077 , \36078 );
and \g453745/U$2 ( \36080 , \16334 , RIdf24b08_1794);
and \g453745/U$3 ( \36081 , RIdf265c0_1813, \16380 );
nor \g453745/U$1 ( \36082 , \36080 , \36081 );
nand \g447424/U$1 ( \36083 , \36068 , \36076 , \36079 , \36082 );
and \g444805/U$3 ( \36084 , \16481 , \36083 );
nor \g444805/U$1 ( \36085 , \36064 , \36084 );
and \g447161/U$2 ( \36086 , \17274 , RIfc42578_5777);
and \g447161/U$3 ( \36087 , RIfc74708_6347, \17276 );
nor \g447161/U$1 ( \36088 , \36086 , \36087 );
and \g447163/U$2 ( \36089 , \17279 , RIfc745a0_6346);
and \g447163/U$3 ( \36090 , RIfc43388_5787, \17281 );
nor \g447163/U$1 ( \36091 , \36089 , \36090 );
and \g447162/U$2 ( \36092 , \17284 , RIdf195a0_1665);
and \g447162/U$3 ( \36093 , RIfcaff10_7024, \17286 );
nor \g447162/U$1 ( \36094 , \36092 , \36093 );
nand \g444538/U$1 ( \36095 , \36085 , \36088 , \36091 , \36094 );
and \g446406/U$2 ( \36096 , RIdeb1d10_487, \16427 );
and \g446406/U$3 ( \36097 , RIdeaf010_455, \16368 );
and \g449403/U$2 ( \36098 , RIdec2b10_679, \16319 );
and \g449403/U$3 ( \36099 , \16326 , RIdec5810_711);
and \g449403/U$4 ( \36100 , RIdeaadf8_423, \16398 );
nor \g449403/U$1 ( \36101 , \36098 , \36099 , \36100 );
and \g455118/U$2 ( \36102 , \16317 , RIdebd110_615);
and \g455118/U$3 ( \36103 , RIfc95228_6719, \16325 );
nor \g455118/U$1 ( \36104 , \36102 , \36103 );
not \g450423/U$3 ( \36105 , \36104 );
not \g450423/U$4 ( \36106 , \16330 );
and \g450423/U$2 ( \36107 , \36105 , \36106 );
and \g450423/U$5 ( \36108 , \16341 , RIfca4f48_6899);
nor \g450423/U$1 ( \36109 , \36107 , \36108 );
and \g453717/U$2 ( \36110 , \16377 , RIdebfe10_647);
and \g453717/U$3 ( \36111 , RIfce6f60_7650, \16313 );
nor \g453717/U$1 ( \36112 , \36110 , \36111 );
and \g453718/U$2 ( \36113 , \16334 , RIdeb7710_551);
and \g453718/U$3 ( \36114 , RIdeba410_583, \16380 );
nor \g453718/U$1 ( \36115 , \36113 , \36114 );
nand \g447423/U$1 ( \36116 , \36101 , \36109 , \36112 , \36115 );
nor \g446406/U$1 ( \36117 , \36096 , \36097 , \36116 );
and \g453714/U$2 ( \36118 , \16361 , RIde9dbf8_359);
and \g453714/U$3 ( \36119 , RIfe879a8_7887, \16448 );
nor \g453714/U$1 ( \36120 , \36118 , \36119 );
and \g453712/U$2 ( \36121 , \16364 , RIdea44f8_391);
and \g453712/U$3 ( \36122 , RIfcc16e8_7223, \16371 );
nor \g453712/U$1 ( \36123 , \36121 , \36122 );
and \g445436/U$2 ( \36124 , \36117 , \36120 , \36123 );
nor \g445436/U$1 ( \36125 , \36124 , \16618 );
and \g446410/U$2 ( \36126 , RIee33478_5042, \16319 );
and \g446410/U$3 ( \36127 , RIfc71b70_6316, \16313 );
and \g449405/U$2 ( \36128 , RIdf33748_1962, \16398 );
and \g449405/U$3 ( \36129 , \16341 , RIdf35bd8_1988);
and \g449405/U$4 ( \36130 , RIfe87570_7884, \16485 );
nor \g449405/U$1 ( \36131 , \36128 , \36129 , \36130 );
and \g455367/U$2 ( \36132 , \16317 , RIfccf0e0_7378);
and \g455367/U$3 ( \36133 , RIfcc99b0_7316, \16325 );
nor \g455367/U$1 ( \36134 , \36132 , \36133 );
not \g450425/U$3 ( \36135 , \36134 );
not \g450425/U$4 ( \36136 , \16351 );
and \g450425/U$2 ( \36137 , \36135 , \36136 );
and \g450425/U$5 ( \36138 , \16354 , RIe1411e0_2118);
nor \g450425/U$1 ( \36139 , \36137 , \36138 );
and \g453734/U$2 ( \36140 , \16361 , RIdf2f530_1915);
and \g453734/U$3 ( \36141 , RIdf31588_1938, \16364 );
nor \g453734/U$1 ( \36142 , \36140 , \36141 );
and \g453732/U$2 ( \36143 , \16368 , RIfcca220_7322);
and \g453732/U$3 ( \36144 , RIfcaeb60_7010, \16371 );
nor \g453732/U$1 ( \36145 , \36143 , \36144 );
nand \g447951/U$1 ( \36146 , \36131 , \36139 , \36142 , \36145 );
nor \g446410/U$1 ( \36147 , \36126 , \36127 , \36146 );
and \g453728/U$2 ( \36148 , \16377 , RIee312b8_5018);
and \g453728/U$3 ( \36149 , RIdf3cf28_2070, \16380 );
nor \g453728/U$1 ( \36150 , \36148 , \36149 );
and \g453726/U$2 ( \36151 , \16334 , RIfe87408_7883);
and \g453726/U$3 ( \36152 , RIfc62288_6139, \16328 );
nor \g453726/U$1 ( \36153 , \36151 , \36152 );
and \g445438/U$2 ( \36154 , \36147 , \36150 , \36153 );
nor \g445438/U$1 ( \36155 , \36154 , \16393 );
or \g444411/U$1 ( \36156 , \36035 , \36095 , \36125 , \36155 );
and \g446400/U$2 ( \36157 , RIe162b10_2500, \16321 );
and \g446400/U$3 ( \36158 , RIee377f8_5090, \16313 );
and \g449396/U$2 ( \36159 , RIe151d10_2308, \16427 );
and \g449396/U$3 ( \36160 , \16448 , RIfc3f3c8_5745);
and \g449396/U$4 ( \36161 , RIe15d110_2436, \16344 );
nor \g449396/U$1 ( \36162 , \36159 , \36160 , \36161 );
and \g454850/U$2 ( \36163 , \16317 , RIe14c310_2244);
and \g454850/U$3 ( \36164 , RIfc4a2a0_5866, \16325 );
nor \g454850/U$1 ( \36165 , \36163 , \36164 );
not \g454849/U$1 ( \36166 , \36165 );
and \g450416/U$2 ( \36167 , \36166 , \16336 );
and \g450416/U$3 ( \36168 , RIee36448_5076, \16356 );
nor \g450416/U$1 ( \36169 , \36167 , \36168 );
and \g453694/U$2 ( \36170 , \16361 , RIe146910_2180);
and \g453694/U$3 ( \36171 , RIe149610_2212, \16364 );
nor \g453694/U$1 ( \36172 , \36170 , \36171 );
and \g453692/U$2 ( \36173 , \16368 , RIe14f010_2276);
and \g453692/U$3 ( \36174 , RIfcde9c8_7555, \16371 );
nor \g453692/U$1 ( \36175 , \36173 , \36174 );
nand \g448119/U$1 ( \36176 , \36162 , \36169 , \36172 , \36175 );
nor \g446400/U$1 ( \36177 , \36157 , \36158 , \36176 );
and \g453687/U$2 ( \36178 , \16377 , RIe15fe10_2468);
and \g453687/U$3 ( \36179 , RIe157710_2372, \16380 );
nor \g453687/U$1 ( \36180 , \36178 , \36179 );
and \g453686/U$2 ( \36181 , \16334 , RIe154a10_2340);
and \g453686/U$3 ( \36182 , RIe165810_2532, \16328 );
nor \g453686/U$1 ( \36183 , \36181 , \36182 );
and \g445429/U$2 ( \36184 , \36177 , \36180 , \36183 );
nor \g445429/U$1 ( \36185 , \36184 , \16389 );
and \g446403/U$2 ( \36186 , RIee1bfd0_4777, \16321 );
and \g446403/U$3 ( \36187 , RIfc95660_6722, \16313 );
and \g449400/U$2 ( \36188 , RIe16ba80_2602, \16398 );
and \g449400/U$3 ( \36189 , \16341 , RIfcd8050_7480);
and \g449400/U$4 ( \36190 , RIfe876d8_7885, \16485 );
nor \g449400/U$1 ( \36191 , \36188 , \36189 , \36190 );
and \g455119/U$2 ( \36192 , \16317 , RIfcee9b8_7737);
and \g455119/U$3 ( \36193 , RIfcb0780_7030, \16325 );
nor \g455119/U$1 ( \36194 , \36192 , \36193 );
not \g450421/U$3 ( \36195 , \36194 );
not \g450421/U$4 ( \36196 , \16351 );
and \g450421/U$2 ( \36197 , \36195 , \36196 );
and \g450421/U$5 ( \36198 , \16356 , RIfe87840_7886);
nor \g450421/U$1 ( \36199 , \36197 , \36198 );
and \g453707/U$2 ( \36200 , \16361 , RIe1680d8_2561);
and \g453707/U$3 ( \36201 , RIfca5380_6902, \16364 );
nor \g453707/U$1 ( \36202 , \36200 , \36201 );
and \g453706/U$2 ( \36203 , \16368 , RIfcdee00_7558);
and \g453706/U$3 ( \36204 , RIfc5f150_6104, \16371 );
nor \g453706/U$1 ( \36205 , \36203 , \36204 );
nand \g447946/U$1 ( \36206 , \36191 , \36199 , \36202 , \36205 );
nor \g446403/U$1 ( \36207 , \36186 , \36187 , \36206 );
and \g453701/U$2 ( \36208 , \16377 , RIfcee148_7731);
and \g453701/U$3 ( \36209 , RIde8a0f8_263, \16380 );
nor \g453701/U$1 ( \36210 , \36208 , \36209 );
and \g453699/U$2 ( \36211 , \16334 , RIde85f58_243);
and \g453699/U$3 ( \36212 , RIee1cf48_4788, \16328 );
nor \g453699/U$1 ( \36213 , \36211 , \36212 );
and \g445432/U$2 ( \36214 , \36207 , \36210 , \36213 );
nor \g445432/U$1 ( \36215 , \36214 , \16649 );
or \g444220/U$1 ( \36216 , \36156 , \36185 , \36215 );
_DC \g5db2/U$1 ( \36217 , \36216 , \16652 );
and \g447174/U$2 ( \36218 , \13244 , RIe171318_2665);
and \g447174/U$3 ( \36219 , RIe1aece0_3366, \13246 );
nor \g447174/U$1 ( \36220 , \36218 , \36219 );
and \g446432/U$2 ( \36221 , RIe1fef60_4278, \8488 );
and \g446432/U$3 ( \36222 , RIe204f00_4346, \8359 );
and \g449433/U$2 ( \36223 , RIe226b00_4730, \8414 );
and \g449433/U$3 ( \36224 , \8409 , RIe1791a8_2755);
and \g449433/U$4 ( \36225 , RIe1bbe68_3515, \8326 );
nor \g449433/U$1 ( \36226 , \36223 , \36224 , \36225 );
and \g455068/U$2 ( \36227 , \8313 , RIe1a34a8_3235);
and \g455068/U$3 ( \36228 , RIe1a61a8_3267, \8323 );
nor \g455068/U$1 ( \36229 , \36227 , \36228 );
not \g450454/U$3 ( \36230 , \36229 );
not \g450454/U$4 ( \36231 , \8328 );
and \g450454/U$2 ( \36232 , \36230 , \36231 );
and \g450454/U$5 ( \36233 , \8340 , RIe1d5368_3803);
nor \g450454/U$1 ( \36234 , \36232 , \36233 );
and \g453838/U$2 ( \36235 , \8404 , RIe1a07a8_3203);
and \g453838/U$3 ( \36236 , RIe1a8ea8_3299, \8351 );
nor \g453838/U$1 ( \36237 , \36235 , \36236 );
and \g453839/U$2 ( \36238 , \8378 , RIe21b700_4602);
and \g453839/U$3 ( \36239 , RIe18cca8_2979, \8417 );
nor \g453839/U$1 ( \36240 , \36238 , \36239 );
nand \g447968/U$1 ( \36241 , \36226 , \36234 , \36237 , \36240 );
nor \g446432/U$1 ( \36242 , \36221 , \36222 , \36241 );
not \g444848/U$3 ( \36243 , \36242 );
not \g444848/U$4 ( \36244 , \8651 );
and \g444848/U$2 ( \36245 , \36243 , \36244 );
and \g446435/U$2 ( \36246 , RIfcb23a0_7050, \8351 );
and \g446435/U$3 ( \36247 , RIe1f58e8_4171, \8378 );
and \g449437/U$2 ( \36248 , RIfce1dd0_7592, \8409 );
and \g449437/U$3 ( \36249 , \8531 , RIfc93770_6700);
and \g449437/U$4 ( \36250 , RIfc78380_6390, \8488 );
nor \g449437/U$1 ( \36251 , \36248 , \36249 , \36250 );
and \g455125/U$2 ( \36252 , \8313 , RIfc93a40_6702);
and \g455125/U$3 ( \36253 , RIfce1b00_7590, \8323 );
nor \g455125/U$1 ( \36254 , \36252 , \36253 );
not \g455124/U$1 ( \36255 , \36254 );
and \g450459/U$2 ( \36256 , \36255 , \8316 );
and \g450459/U$3 ( \36257 , RIfcd4c48_7443, \8417 );
nor \g450459/U$1 ( \36258 , \36256 , \36257 );
and \g453853/U$2 ( \36259 , \8335 , RIe1ee2c8_4087);
and \g453853/U$3 ( \36260 , RIfcb1f68_7047, \8340 );
nor \g453853/U$1 ( \36261 , \36259 , \36260 );
and \g453852/U$2 ( \36262 , \8356 , RIe1f35c0_4146);
and \g453852/U$3 ( \36263 , RIfcbfc30_7204, \8359 );
nor \g453852/U$1 ( \36264 , \36262 , \36263 );
nand \g448241/U$1 ( \36265 , \36251 , \36258 , \36261 , \36264 );
nor \g446435/U$1 ( \36266 , \36246 , \36247 , \36265 );
and \g453847/U$2 ( \36267 , \8404 , RIe1fa370_4224);
and \g453847/U$3 ( \36268 , RIfcbf960_7202, \8414 );
nor \g453847/U$1 ( \36269 , \36267 , \36268 );
and \g453846/U$2 ( \36270 , \8373 , RIfcede78_7729);
and \g453846/U$3 ( \36271 , RIfc5bbe0_6066, \8330 );
nor \g453846/U$1 ( \36272 , \36270 , \36271 );
and \g445456/U$2 ( \36273 , \36266 , \36269 , \36272 );
nor \g445456/U$1 ( \36274 , \36273 , \8621 );
nor \g444848/U$1 ( \36275 , \36245 , \36274 );
and \g447175/U$2 ( \36276 , \11213 , RIe1f0e60_4118);
and \g447175/U$3 ( \36277 , RIe1f8318_4201, \11215 );
nor \g447175/U$1 ( \36278 , \36276 , \36277 );
nand \g444438/U$1 ( \36279 , \36220 , \36275 , \36278 );
and \g453869/U$2 ( \36280 , \8531 , RIfcbee20_7194);
and \g453869/U$3 ( \36281 , RIe213000_4506, \8488 );
nor \g453869/U$1 ( \36282 , \36280 , \36281 );
and \g446441/U$2 ( \36283 , RIe215d00_4538, \8378 );
and \g446441/U$3 ( \36284 , RIfc79e38_6409, \8359 );
and \g449445/U$2 ( \36285 , RIe21e400_4634, \8407 );
and \g449445/U$3 ( \36286 , \8373 , RIfcd8488_7483);
and \g449445/U$4 ( \36287 , RIe223e00_4698, \8383 );
nor \g449445/U$1 ( \36288 , \36285 , \36286 , \36287 );
and \g453877/U$2 ( \36289 , \8335 , RIe207c00_4378);
and \g453877/U$3 ( \36290 , RIf168068_5643, \8340 );
nor \g453877/U$1 ( \36291 , \36289 , \36290 );
and \g453876/U$2 ( \36292 , \8404 , RIe221100_4666);
and \g453876/U$3 ( \36293 , RIfea9710_8244, \8351 );
nor \g453876/U$1 ( \36294 , \36292 , \36293 );
and \g454843/U$2 ( \36295 , \8313 , RIe20a900_4410);
and \g454843/U$3 ( \36296 , RIe20d600_4442, \8323 );
nor \g454843/U$1 ( \36297 , \36295 , \36296 );
not \g454842/U$1 ( \36298 , \36297 );
and \g450465/U$2 ( \36299 , \36298 , \8316 );
and \g450465/U$3 ( \36300 , RIfc920f0_6684, \8417 );
nor \g450465/U$1 ( \36301 , \36299 , \36300 );
nand \g448242/U$1 ( \36302 , \36288 , \36291 , \36294 , \36301 );
nor \g446441/U$1 ( \36303 , \36283 , \36284 , \36302 );
and \g453873/U$2 ( \36304 , \8356 , RIe210300_4474);
and \g453873/U$3 ( \36305 , RIe218a00_4570, \8414 );
nor \g453873/U$1 ( \36306 , \36304 , \36305 );
nand \g445690/U$1 ( \36307 , \36282 , \36303 , \36306 );
and \g444855/U$2 ( \36308 , \36307 , \8369 );
and \g449442/U$2 ( \36309 , RIfc93338_6697, \8319 );
and \g449442/U$3 ( \36310 , \8324 , RIfec1158_8317);
and \g449442/U$4 ( \36311 , RIfcdf940_7566, \8407 );
nor \g449442/U$1 ( \36312 , \36309 , \36310 , \36311 );
and \g454930/U$2 ( \36313 , \8313 , RIfe872a0_7882);
and \g454930/U$3 ( \36314 , RIf15e5b8_5533, \8323 );
nor \g454930/U$1 ( \36315 , \36313 , \36314 );
not \g450462/U$3 ( \36316 , \36315 );
not \g450462/U$4 ( \36317 , \8347 );
and \g450462/U$2 ( \36318 , \36316 , \36317 );
and \g450462/U$5 ( \36319 , \8417 , RIfcb2670_7052);
nor \g450462/U$1 ( \36320 , \36318 , \36319 );
and \g453864/U$2 ( \36321 , \8335 , RIfcea368_7687);
and \g453864/U$3 ( \36322 , RIfc78920_6394, \8340 );
nor \g453864/U$1 ( \36323 , \36321 , \36322 );
and \g453862/U$2 ( \36324 , \8356 , RIfe87138_7881);
and \g453862/U$3 ( \36325 , RIf1604a8_5555, \8359 );
nor \g453862/U$1 ( \36326 , \36324 , \36325 );
nand \g447971/U$1 ( \36327 , \36312 , \36320 , \36323 , \36326 );
and \g444855/U$3 ( \36328 , \9266 , \36327 );
nor \g444855/U$1 ( \36329 , \36308 , \36328 );
and \g447181/U$2 ( \36330 , \14165 , RIfcbf3c0_7198);
and \g447181/U$3 ( \36331 , RIfc5b208_6059, \14167 );
nor \g447181/U$1 ( \36332 , \36330 , \36331 );
and \g447178/U$2 ( \36333 , \9293 , RIfcd73a8_7471);
and \g447178/U$3 ( \36334 , RIfc5af38_6057, \9296 );
nor \g447178/U$1 ( \36335 , \36333 , \36334 );
and \g447183/U$2 ( \36336 , \9288 , RIe200ce8_4299);
and \g447183/U$3 ( \36337 , RIe2027a0_4318, \9290 );
nor \g447183/U$1 ( \36338 , \36336 , \36337 );
nand \g444662/U$1 ( \36339 , \36329 , \36332 , \36335 , \36338 );
and \g446426/U$2 ( \36340 , RIe1ebb68_4059, \8351 );
and \g446426/U$3 ( \36341 , RIe1d8068_3835, \8378 );
and \g449427/U$2 ( \36342 , RIe1dda68_3899, \8409 );
and \g449427/U$3 ( \36343 , \8531 , RIe1ccc68_3707);
and \g449427/U$4 ( \36344 , RIe1cf968_3739, \8488 );
nor \g449427/U$1 ( \36345 , \36342 , \36343 , \36344 );
and \g455079/U$2 ( \36346 , \8313 , RIe1c1868_3579);
and \g455079/U$3 ( \36347 , RIe1c4568_3611, \8323 );
nor \g455079/U$1 ( \36348 , \36346 , \36347 );
not \g455078/U$1 ( \36349 , \36348 );
and \g450449/U$2 ( \36350 , \36349 , \8316 );
and \g450449/U$3 ( \36351 , RIe1e0768_3931, \8417 );
nor \g450449/U$1 ( \36352 , \36350 , \36351 );
and \g453815/U$2 ( \36353 , \8335 , RIe1beb68_3547);
and \g453815/U$3 ( \36354 , RIe1c7268_3643, \8340 );
nor \g453815/U$1 ( \36355 , \36353 , \36354 );
and \g453814/U$2 ( \36356 , \8356 , RIe1c9f68_3675);
and \g453814/U$3 ( \36357 , RIe1d2668_3771, \8359 );
nor \g453814/U$1 ( \36358 , \36356 , \36357 );
nand \g448239/U$1 ( \36359 , \36345 , \36352 , \36355 , \36358 );
nor \g446426/U$1 ( \36360 , \36340 , \36341 , \36359 );
and \g453811/U$2 ( \36361 , \8404 , RIe1e3468_3963);
and \g453811/U$3 ( \36362 , RIe1dad68_3867, \8414 );
nor \g453811/U$1 ( \36363 , \36361 , \36362 );
and \g453810/U$2 ( \36364 , \8373 , RIe1e6168_3995);
and \g453810/U$3 ( \36365 , RIe1e8e68_4027, \8330 );
nor \g453810/U$1 ( \36366 , \36364 , \36365 );
and \g445447/U$2 ( \36367 , \36360 , \36363 , \36366 );
nor \g445447/U$1 ( \36368 , \36367 , \8477 );
and \g446428/U$2 ( \36369 , RIfcdec98_7557, \8351 );
and \g446428/U$3 ( \36370 , RIe1b3fd8_3425, \8378 );
and \g449430/U$2 ( \36371 , RIfceabd8_7693, \8409 );
and \g449430/U$3 ( \36372 , \8531 , RIe1b27f0_3408);
and \g449430/U$4 ( \36373 , RIfcd7c18_7477, \8488 );
nor \g449430/U$1 ( \36374 , \36371 , \36372 , \36373 );
and \g455177/U$2 ( \36375 , \8313 , RIe1ac6e8_3339);
and \g455177/U$3 ( \36376 , RIfce2640_7598, \8323 );
nor \g455177/U$1 ( \36377 , \36375 , \36376 );
not \g455176/U$1 ( \36378 , \36377 );
and \g450451/U$2 ( \36379 , \36378 , \8316 );
and \g450451/U$3 ( \36380 , RIfcd12a0_7402, \8417 );
nor \g450451/U$1 ( \36381 , \36379 , \36380 );
and \g453826/U$2 ( \36382 , \8335 , RIe1ab068_3323);
and \g453826/U$3 ( \36383 , RIfc76a30_6372, \8340 );
nor \g453826/U$1 ( \36384 , \36382 , \36383 );
and \g453823/U$2 ( \36385 , \8356 , RIe1b0d38_3389);
and \g453823/U$3 ( \36386 , RIfc94850_6712, \8359 );
nor \g453823/U$1 ( \36387 , \36385 , \36386 );
nand \g448240/U$1 ( \36388 , \36374 , \36381 , \36384 , \36387 );
nor \g446428/U$1 ( \36389 , \36369 , \36370 , \36388 );
and \g453819/U$2 ( \36390 , \8404 , RIe1b7548_3463);
and \g453819/U$3 ( \36391 , RIe1b5388_3439, \8414 );
nor \g453819/U$1 ( \36392 , \36390 , \36391 );
and \g453818/U$2 ( \36393 , \8373 , RIe1b95a0_3486);
and \g453818/U$3 ( \36394 , RIfc94148_6707, \8330 );
nor \g453818/U$1 ( \36395 , \36393 , \36394 );
and \g445452/U$2 ( \36396 , \36389 , \36392 , \36395 );
nor \g445452/U$1 ( \36397 , \36396 , \8481 );
or \g444296/U$1 ( \36398 , \36279 , \36339 , \36368 , \36397 );
and \g446421/U$2 ( \36399 , RIe19daa8_3171, \8351 );
and \g446421/U$3 ( \36400 , RIe1980a8_3107, \8404 );
and \g449420/U$2 ( \36401 , RIe1953a8_3075, \8409 );
and \g449420/U$3 ( \36402 , \8523 , RIf143ba0_5230);
and \g449420/U$4 ( \36403 , RIe1872a8_2915, \8486 );
nor \g449420/U$1 ( \36404 , \36401 , \36402 , \36403 );
and \g454160/U$2 ( \36405 , \8313 , RIe17eba8_2819);
and \g454160/U$3 ( \36406 , RIe1818a8_2851, \8323 );
nor \g454160/U$1 ( \36407 , \36405 , \36406 );
not \g454159/U$1 ( \36408 , \36407 );
and \g450441/U$2 ( \36409 , \36408 , \8316 );
and \g450441/U$3 ( \36410 , RIf1449b0_5240, \8417 );
nor \g450441/U$1 ( \36411 , \36409 , \36410 );
and \g453790/U$2 ( \36412 , \8335 , RIe17bea8_2787);
and \g453790/U$3 ( \36413 , RIfc912e0_6674, \8340 );
nor \g453790/U$1 ( \36414 , \36412 , \36413 );
and \g453789/U$2 ( \36415 , \8356 , RIe1845a8_2883);
and \g453789/U$3 ( \36416 , RIe189fa8_2947, \8359 );
nor \g453789/U$1 ( \36417 , \36415 , \36416 );
nand \g448238/U$1 ( \36418 , \36404 , \36411 , \36414 , \36417 );
nor \g446421/U$1 ( \36419 , \36399 , \36400 , \36418 );
and \g453787/U$2 ( \36420 , \8378 , RIe18f9a8_3011);
and \g453787/U$3 ( \36421 , RIe19ada8_3139, \8383 );
nor \g453787/U$1 ( \36422 , \36420 , \36421 );
and \g453785/U$2 ( \36423 , \8412 , RIe1926a8_3043);
and \g453785/U$3 ( \36424 , RIf1457c0_5250, \8373 );
nor \g453785/U$1 ( \36425 , \36423 , \36424 );
and \g445445/U$2 ( \36426 , \36419 , \36422 , \36425 );
nor \g445445/U$1 ( \36427 , \36426 , \8589 );
and \g446424/U$2 ( \36428 , RIfc7a810_6416, \8359 );
and \g446424/U$3 ( \36429 , RIfc429b0_5780, \8335 );
and \g449422/U$2 ( \36430 , RIfc7a540_6414, \8326 );
and \g449422/U$3 ( \36431 , \8373 , RIfce3b58_7613);
and \g449422/U$4 ( \36432 , RIfcbe5b0_7188, \8383 );
nor \g449422/U$1 ( \36433 , \36430 , \36431 , \36432 );
and \g455030/U$2 ( \36434 , \8313 , RIfc42de8_5783);
and \g455030/U$3 ( \36435 , RIfcc7958_7293, \8323 );
nor \g455030/U$1 ( \36436 , \36434 , \36435 );
not \g450445/U$3 ( \36437 , \36436 );
not \g450445/U$4 ( \36438 , \8376 );
and \g450445/U$2 ( \36439 , \36437 , \36438 );
and \g450445/U$5 ( \36440 , \8340 , RIfce39f0_7612);
nor \g450445/U$1 ( \36441 , \36439 , \36440 );
and \g453803/U$2 ( \36442 , \8404 , RIe175da0_2718);
and \g453803/U$3 ( \36443 , RIfc915b0_6676, \8351 );
nor \g453803/U$1 ( \36444 , \36442 , \36443 );
and \g453805/U$2 ( \36445 , \8378 , RIfc96e48_6739);
and \g453805/U$3 ( \36446 , RIfceb448_7699, \8417 );
nor \g453805/U$1 ( \36447 , \36445 , \36446 );
nand \g447962/U$1 ( \36448 , \36433 , \36441 , \36444 , \36447 );
nor \g446424/U$1 ( \36449 , \36428 , \36429 , \36448 );
and \g453799/U$2 ( \36450 , \8319 , RIfc91b50_6680);
and \g453799/U$3 ( \36451 , RIe173be0_2694, \8356 );
nor \g453799/U$1 ( \36452 , \36450 , \36451 );
and \g453798/U$2 ( \36453 , \8531 , RIfcc7ac0_7294);
and \g453798/U$3 ( \36454 , RIfc96ce0_6738, \8486 );
nor \g453798/U$1 ( \36455 , \36453 , \36454 );
and \g445446/U$2 ( \36456 , \36449 , \36452 , \36455 );
nor \g445446/U$1 ( \36457 , \36456 , \8558 );
or \g444203/U$1 ( \36458 , \36398 , \36427 , \36457 );
_DC \g5e36/U$1 ( \36459 , \36458 , \8654 );
and \g447224/U$2 ( \36460 , \17779 , RIdec8678_744);
and \g447224/U$3 ( \36461 , RIdecb378_776, \17781 );
nor \g447224/U$1 ( \36462 , \36460 , \36461 );
and \g446490/U$2 ( \36463 , RIded0d78_840, \16328 );
and \g446490/U$3 ( \36464 , RIdece078_808, \16321 );
and \g449500/U$2 ( \36465 , RIdee7848_1098, \16398 );
and \g449500/U$3 ( \36466 , \16341 , RIdf00d48_1386);
and \g449500/U$4 ( \36467 , RIde97640_328, \16485 );
nor \g449500/U$1 ( \36468 , \36465 , \36466 , \36467 );
and \g455110/U$2 ( \36469 , \16317 , RIdf38770_2019);
and \g455110/U$3 ( \36470 , RIe143d78_2149, \16325 );
nor \g455110/U$1 ( \36471 , \36469 , \36470 );
not \g450522/U$3 ( \36472 , \36471 );
not \g450522/U$4 ( \36473 , \16351 );
and \g450522/U$2 ( \36474 , \36472 , \36473 );
and \g450522/U$5 ( \36475 , \16356 , RIdeb4b78_520);
nor \g450522/U$1 ( \36476 , \36474 , \36475 );
and \g454082/U$2 ( \36477 , \16361 , RIde7d588_201);
and \g454082/U$3 ( \36478 , RIdedc5b0_971, \16364 );
nor \g454082/U$1 ( \36479 , \36477 , \36478 );
and \g454081/U$2 ( \36480 , \16368 , RIdf1d650_1711);
and \g454081/U$3 ( \36481 , RIdf2cdd0_1887, \16371 );
nor \g454081/U$1 ( \36482 , \36480 , \36481 );
nand \g447998/U$1 ( \36483 , \36468 , \36476 , \36479 , \36482 );
nor \g446490/U$1 ( \36484 , \36463 , \36464 , \36483 );
not \g444928/U$3 ( \36485 , \36484 );
not \g444928/U$4 ( \36486 , \16586 );
and \g444928/U$2 ( \36487 , \36485 , \36486 );
and \g446491/U$2 ( \36488 , RIfc7cb38_6441, \16321 );
and \g446491/U$3 ( \36489 , RIfc97af0_6748, \16313 );
and \g449503/U$2 ( \36490 , RIfcc2930_7236, \16427 );
and \g449503/U$3 ( \36491 , \16448 , RIfc97dc0_6750);
and \g449503/U$4 ( \36492 , RIdee3090_1047, \16344 );
nor \g449503/U$1 ( \36493 , \36490 , \36491 , \36492 );
and \g455311/U$2 ( \36494 , \16317 , RIded76f0_915);
and \g455311/U$3 ( \36495 , RIded9ce8_942, \16325 );
nor \g455311/U$1 ( \36496 , \36494 , \36495 );
not \g455310/U$1 ( \36497 , \36496 );
and \g450527/U$2 ( \36498 , \36497 , \16336 );
and \g450527/U$3 ( \36499 , RIdee4e18_1068, \16354 );
nor \g450527/U$1 ( \36500 , \36498 , \36499 );
and \g454097/U$2 ( \36501 , \16361 , RIded3370_867);
and \g454097/U$3 ( \36502 , RIded5968_894, \16364 );
nor \g454097/U$1 ( \36503 , \36501 , \36502 );
and \g454093/U$2 ( \36504 , \16368 , RIfc7c868_6439);
and \g454093/U$3 ( \36505 , RIfcd9298_7493, \16371 );
nor \g454093/U$1 ( \36506 , \36504 , \36505 );
nand \g448129/U$1 ( \36507 , \36493 , \36500 , \36503 , \36506 );
nor \g446491/U$1 ( \36508 , \36488 , \36489 , \36507 );
and \g454090/U$2 ( \36509 , \16377 , RIfcb3e58_7069);
and \g454090/U$3 ( \36510 , RIdee0ed0_1023, \16380 );
nor \g454090/U$1 ( \36511 , \36509 , \36510 );
and \g454089/U$2 ( \36512 , \16334 , RIfe88380_7894);
and \g454089/U$3 ( \36513 , RIfcd9130_7492, \16326 );
nor \g454089/U$1 ( \36514 , \36512 , \36513 );
and \g445494/U$2 ( \36515 , \36508 , \36511 , \36514 );
nor \g445494/U$1 ( \36516 , \36515 , \16909 );
nor \g444928/U$1 ( \36517 , \36487 , \36516 );
and \g447223/U$2 ( \36518 , \17032 , RIe15a578_2405);
and \g447223/U$3 ( \36519 , RIe16e780_2634, \17029 );
nor \g447223/U$1 ( \36520 , \36518 , \36519 );
nand \g444443/U$1 ( \36521 , \36462 , \36517 , \36520 );
and \g449507/U$2 ( \36522 , RIdf14848_1610, \16321 );
and \g449507/U$3 ( \36523 , \16328 , RIdf17548_1642);
and \g449507/U$4 ( \36524 , RIdeeff48_1194, \16398 );
nor \g449507/U$1 ( \36525 , \36522 , \36523 , \36524 );
and \g454948/U$2 ( \36526 , \16317 , RIdf09448_1482);
and \g454948/U$3 ( \36527 , RIdf0c148_1514, \16325 );
nor \g454948/U$1 ( \36528 , \36526 , \36527 );
not \g450530/U$3 ( \36529 , \36528 );
not \g450530/U$4 ( \36530 , \16330 );
and \g450530/U$2 ( \36531 , \36529 , \36530 );
and \g450530/U$5 ( \36532 , \16339 , RIdef2c48_1226);
nor \g450530/U$1 ( \36533 , \36531 , \36532 );
and \g454104/U$2 ( \36534 , \16377 , RIdf0ee48_1546);
and \g454104/U$3 ( \36535 , RIdf11b48_1578, \16313 );
nor \g454104/U$1 ( \36536 , \36534 , \36535 );
and \g454105/U$2 ( \36537 , \16334 , RIdf03a48_1418);
and \g454105/U$3 ( \36538 , RIdf06748_1450, \16380 );
nor \g454105/U$1 ( \36539 , \36537 , \36538 );
nand \g447449/U$1 ( \36540 , \36525 , \36533 , \36536 , \36539 );
and \g444720/U$2 ( \36541 , \36540 , \16750 );
and \g446496/U$2 ( \36542 , RIfc7ecf8_6465, \16448 );
and \g446496/U$3 ( \36543 , RIfc99008_6763, \16371 );
and \g449511/U$2 ( \36544 , RIfce4260_7618, \16319 );
and \g449511/U$3 ( \36545 , \16328 , RIfc7f9a0_6474);
and \g449511/U$4 ( \36546 , RIdf1fdb0_1739, \16398 );
nor \g449511/U$1 ( \36547 , \36544 , \36545 , \36546 );
and \g454982/U$2 ( \36548 , \16317 , RIdf284b0_1835);
and \g454982/U$3 ( \36549 , RIdf2a670_1859, \16325 );
nor \g454982/U$1 ( \36550 , \36548 , \36549 );
not \g450532/U$3 ( \36551 , \36550 );
not \g450532/U$4 ( \36552 , \16330 );
and \g450532/U$2 ( \36553 , \36551 , \36552 );
and \g450532/U$5 ( \36554 , \16341 , RIfce2a78_7601);
nor \g450532/U$1 ( \36555 , \36553 , \36554 );
and \g454114/U$2 ( \36556 , \16377 , RIfce9990_7680);
and \g454114/U$3 ( \36557 , RIfcd62c8_7459, \16313 );
nor \g454114/U$1 ( \36558 , \36556 , \36557 );
and \g454115/U$2 ( \36559 , \16334 , RIdf24c70_1795);
and \g454115/U$3 ( \36560 , RIdf26728_1814, \16380 );
nor \g454115/U$1 ( \36561 , \36559 , \36560 );
nand \g447451/U$1 ( \36562 , \36547 , \36555 , \36558 , \36561 );
nor \g446496/U$1 ( \36563 , \36542 , \36543 , \36562 );
and \g454112/U$2 ( \36564 , \16364 , RIfcc6e18_7285);
and \g454112/U$3 ( \36565 , RIfc46e98_5829, \16368 );
nor \g454112/U$1 ( \36566 , \36564 , \36565 );
and \g454113/U$2 ( \36567 , \16361 , RIdf19708_1666);
and \g454113/U$3 ( \36568 , RIfcc31a0_7242, \16427 );
nor \g454113/U$1 ( \36569 , \36567 , \36568 );
and \g445498/U$2 ( \36570 , \36563 , \36566 , \36569 );
nor \g445498/U$1 ( \36571 , \36570 , \16480 );
nor \g444720/U$1 ( \36572 , \36541 , \36571 );
and \g447229/U$2 ( \36573 , \19208 , RIdeea548_1130);
and \g447229/U$3 ( \36574 , RIdef8648_1290, \19210 );
nor \g447229/U$1 ( \36575 , \36573 , \36574 );
and \g447230/U$2 ( \36576 , \19213 , RIdeed248_1162);
and \g447230/U$3 ( \36577 , RIdef5948_1258, \19215 );
nor \g447230/U$1 ( \36578 , \36576 , \36577 );
and \g447228/U$2 ( \36579 , \19218 , RIdefb348_1322);
and \g447228/U$3 ( \36580 , RIdefe048_1354, \19220 );
nor \g447228/U$1 ( \36581 , \36579 , \36580 );
nand \g444667/U$1 ( \36582 , \36572 , \36575 , \36578 , \36581 );
and \g446483/U$2 ( \36583 , RIdec2c78_680, \16321 );
and \g446483/U$3 ( \36584 , RIfc8aad0_6600, \16313 );
and \g449493/U$2 ( \36585 , RIdeb1e78_488, \16427 );
and \g449493/U$3 ( \36586 , \16448 , RIfc40e80_5764);
and \g449493/U$4 ( \36587 , RIdebd278_616, \16485 );
nor \g449493/U$1 ( \36588 , \36585 , \36586 , \36587 );
and \g455296/U$2 ( \36589 , \16317 , RIdeab140_424);
and \g455296/U$3 ( \36590 , RIee1dbf0_4797, \16325 );
nor \g455296/U$1 ( \36591 , \36589 , \36590 );
not \g455295/U$1 ( \36592 , \36591 );
and \g450517/U$2 ( \36593 , \36592 , \16336 );
and \g450517/U$3 ( \36594 , RIfc8ac38_6601, \16356 );
nor \g450517/U$1 ( \36595 , \36593 , \36594 );
and \g454061/U$2 ( \36596 , \16361 , RIde9df40_360);
and \g454061/U$3 ( \36597 , RIdea4840_392, \16364 );
nor \g454061/U$1 ( \36598 , \36596 , \36597 );
and \g454060/U$2 ( \36599 , \16368 , RIdeaf178_456);
and \g454060/U$3 ( \36600 , RIfcdaeb8_7513, \16371 );
nor \g454060/U$1 ( \36601 , \36599 , \36600 );
nand \g448128/U$1 ( \36602 , \36588 , \36595 , \36598 , \36601 );
nor \g446483/U$1 ( \36603 , \36583 , \36584 , \36602 );
and \g454057/U$2 ( \36604 , \16377 , RIdebff78_648);
and \g454057/U$3 ( \36605 , RIdeba578_584, \16380 );
nor \g454057/U$1 ( \36606 , \36604 , \36605 );
and \g454056/U$2 ( \36607 , \16334 , RIdeb7878_552);
and \g454056/U$3 ( \36608 , RIdec5978_712, \16328 );
nor \g454056/U$1 ( \36609 , \36607 , \36608 );
and \g445489/U$2 ( \36610 , \36603 , \36606 , \36609 );
nor \g445489/U$1 ( \36611 , \36610 , \16618 );
and \g446484/U$2 ( \36612 , RIfc56780_6006, \16427 );
and \g446484/U$3 ( \36613 , RIfce2eb0_7604, \16368 );
and \g449497/U$2 ( \36614 , RIee335e0_5043, \16321 );
and \g449497/U$3 ( \36615 , \16328 , RIee346c0_5055);
and \g449497/U$4 ( \36616 , RIfe88218_7893, \16398 );
nor \g449497/U$1 ( \36617 , \36614 , \36615 , \36616 );
and \g454999/U$2 ( \36618 , \16317 , RIe13f020_2094);
and \g454999/U$3 ( \36619 , RIe141348_2119, \16325 );
nor \g454999/U$1 ( \36620 , \36618 , \36619 );
not \g450520/U$3 ( \36621 , \36620 );
not \g450520/U$4 ( \36622 , \16330 );
and \g450520/U$2 ( \36623 , \36621 , \36622 );
and \g450520/U$5 ( \36624 , \16341 , RIdf35d40_1989);
nor \g450520/U$1 ( \36625 , \36623 , \36624 );
and \g454068/U$2 ( \36626 , \16377 , RIee31420_5019);
and \g454068/U$3 ( \36627 , RIee32398_5030, \16313 );
nor \g454068/U$1 ( \36628 , \36626 , \36627 );
and \g454071/U$2 ( \36629 , \16334 , RIdf3a930_2043);
and \g454071/U$3 ( \36630 , RIfec16f8_8321, \16380 );
nor \g454071/U$1 ( \36631 , \36629 , \36630 );
nand \g447448/U$1 ( \36632 , \36617 , \36625 , \36628 , \36631 );
nor \g446484/U$1 ( \36633 , \36612 , \36613 , \36632 );
and \g454067/U$2 ( \36634 , \16361 , RIdf2f698_1916);
and \g454067/U$3 ( \36635 , RIfce3e28_7615, \16448 );
nor \g454067/U$1 ( \36636 , \36634 , \36635 );
and \g454066/U$2 ( \36637 , \16364 , RIdf316f0_1939);
and \g454066/U$3 ( \36638 , RIfcb4128_7071, \16371 );
nor \g454066/U$1 ( \36639 , \36637 , \36638 );
and \g445491/U$2 ( \36640 , \36633 , \36636 , \36639 );
nor \g445491/U$1 ( \36641 , \36640 , \16393 );
or \g444314/U$1 ( \36642 , \36521 , \36582 , \36611 , \36641 );
and \g446476/U$2 ( \36643 , RIe162c78_2501, \16321 );
and \g446476/U$3 ( \36644 , RIee37960_5091, \16313 );
and \g449488/U$2 ( \36645 , RIe151e78_2309, \16427 );
and \g449488/U$3 ( \36646 , \16432 , RIfc8e5e0_6642);
and \g449488/U$4 ( \36647 , RIe15d278_2437, \16485 );
nor \g449488/U$1 ( \36648 , \36645 , \36646 , \36647 );
and \g455010/U$2 ( \36649 , \16317 , RIe14c478_2245);
and \g455010/U$3 ( \36650 , RIfc56ff0_6012, \16325 );
nor \g455010/U$1 ( \36651 , \36649 , \36650 );
not \g455009/U$1 ( \36652 , \36651 );
and \g450509/U$2 ( \36653 , \36652 , \16336 );
and \g450509/U$3 ( \36654 , RIfcd6b38_7465, \16354 );
nor \g450509/U$1 ( \36655 , \36653 , \36654 );
and \g454035/U$2 ( \36656 , \16361 , RIe146a78_2181);
and \g454035/U$3 ( \36657 , RIe149778_2213, \16364 );
nor \g454035/U$1 ( \36658 , \36656 , \36657 );
and \g454034/U$2 ( \36659 , \16368 , RIe14f178_2277);
and \g454034/U$3 ( \36660 , RIfcb4290_7072, \16371 );
nor \g454034/U$1 ( \36661 , \36659 , \36660 );
nand \g448126/U$1 ( \36662 , \36648 , \36655 , \36658 , \36661 );
nor \g446476/U$1 ( \36663 , \36643 , \36644 , \36662 );
and \g454030/U$2 ( \36664 , \16377 , RIe15ff78_2469);
and \g454030/U$3 ( \36665 , RIe157878_2373, \16380 );
nor \g454030/U$1 ( \36666 , \36664 , \36665 );
and \g454029/U$2 ( \36667 , \16334 , RIe154b78_2341);
and \g454029/U$3 ( \36668 , RIe165978_2533, \16328 );
nor \g454029/U$1 ( \36669 , \36667 , \36668 );
and \g445481/U$2 ( \36670 , \36663 , \36666 , \36669 );
nor \g445481/U$1 ( \36671 , \36670 , \16389 );
and \g446478/U$2 ( \36672 , RIfcbbb80_7158, \16427 );
and \g446478/U$3 ( \36673 , RIfcbbfb8_7161, \16368 );
and \g449491/U$2 ( \36674 , RIde8e298_283, \16485 );
and \g449491/U$3 ( \36675 , \16356 , RIde91a60_300);
and \g449491/U$4 ( \36676 , RIe16bbe8_2603, \16398 );
nor \g449491/U$1 ( \36677 , \36674 , \36675 , \36676 );
and \g454257/U$2 ( \36678 , \16317 , RIfcc38a8_7247);
and \g454257/U$3 ( \36679 , RIfc8b070_6604, \16325 );
nor \g454257/U$1 ( \36680 , \36678 , \36679 );
not \g450512/U$3 ( \36681 , \36680 );
not \g450512/U$4 ( \36682 , \16311 );
and \g450512/U$2 ( \36683 , \36681 , \36682 );
and \g450512/U$5 ( \36684 , \16341 , RIfc54458_5981);
nor \g450512/U$1 ( \36685 , \36683 , \36684 );
and \g454047/U$2 ( \36686 , \16377 , RIfcbb8b0_7156);
and \g454047/U$3 ( \36687 , RIfc807b0_6484, \16313 );
nor \g454047/U$1 ( \36688 , \36686 , \36687 );
and \g454048/U$2 ( \36689 , \16334 , RIde862a0_244);
and \g454048/U$3 ( \36690 , RIde8a440_264, \16380 );
nor \g454048/U$1 ( \36691 , \36689 , \36690 );
nand \g447446/U$1 ( \36692 , \36677 , \36685 , \36688 , \36691 );
nor \g446478/U$1 ( \36693 , \36672 , \36673 , \36692 );
and \g454044/U$2 ( \36694 , \16361 , RIe168240_2562);
and \g454044/U$3 ( \36695 , RIde82100_224, \16448 );
nor \g454044/U$1 ( \36696 , \36694 , \36695 );
and \g454040/U$2 ( \36697 , \16364 , RIfc8c2b8_6617);
and \g454040/U$3 ( \36698 , RIfc8c150_6616, \16371 );
nor \g454040/U$1 ( \36699 , \36697 , \36698 );
and \g445486/U$2 ( \36700 , \36693 , \36696 , \36699 );
nor \g445486/U$1 ( \36701 , \36700 , \16649 );
or \g444204/U$1 ( \36702 , \36642 , \36671 , \36701 );
_DC \g5ebb/U$1 ( \36703 , \36702 , \16652 );
and \g450610/U$2 ( \36704 , \8317 , RIe1ac850_3340);
and \g450610/U$3 ( \36705 , RIe1b9708_3487, \8371 );
nor \g450610/U$1 ( \36706 , \36704 , \36705 );
and \g445715/U$2 ( \36707 , RIfce0b88_7579, \8351 );
and \g445715/U$3 ( \36708 , RIe1b76b0_3464, \8404 );
and \g448511/U$2 ( \36709 , RIfc8a260_6594, \8324 );
and \g448511/U$3 ( \36710 , \8531 , RIe1b2958_3409);
and \g448511/U$4 ( \36711 , RIfce9af8_7681, \8488 );
nor \g448511/U$1 ( \36712 , \36709 , \36710 , \36711 );
and \g450616/U$2 ( \36713 , \8356 , RIe1b0ea0_3390);
and \g450616/U$3 ( \36714 , RIfc89f90_6592, \8359 );
nor \g450616/U$1 ( \36715 , \36713 , \36714 );
and \g454532/U$2 ( \36716 , \8313 , RIe1b54f0_3440);
and \g454532/U$3 ( \36717 , RIfcb69f0_7100, \8323 );
nor \g454532/U$1 ( \36718 , \36716 , \36717 );
not \g449532/U$3 ( \36719 , \36718 );
not \g449532/U$4 ( \36720 , \8376 );
and \g449532/U$2 ( \36721 , \36719 , \36720 );
and \g449532/U$5 ( \36722 , \8340 , RIfc4a138_5865);
nor \g449532/U$1 ( \36723 , \36721 , \36722 );
and \g450615/U$2 ( \36724 , \8378 , RIe1b4140_3426);
and \g450615/U$3 ( \36725 , RIfcd5bc0_7454, \8417 );
nor \g450615/U$1 ( \36726 , \36724 , \36725 );
nand \g447466/U$1 ( \36727 , \36712 , \36715 , \36723 , \36726 );
nor \g445715/U$1 ( \36728 , \36707 , \36708 , \36727 );
and \g450613/U$2 ( \36729 , \8335 , RIe1ab1d0_3324);
and \g450613/U$3 ( \36730 , RIfc82808_6507, \8383 );
nor \g450613/U$1 ( \36731 , \36729 , \36730 );
nand \g445509/U$1 ( \36732 , \36706 , \36728 , \36731 );
and \g444903/U$2 ( \36733 , \36732 , \8482 );
and \g448509/U$2 ( \36734 , RIe226c68_4731, \8414 );
and \g448509/U$3 ( \36735 , \8409 , RIe179310_2756);
and \g448509/U$4 ( \36736 , RIe1bbfd0_3516, \8324 );
nor \g448509/U$1 ( \36737 , \36734 , \36735 , \36736 );
and \g450607/U$2 ( \36738 , \8356 , RIe1f0fc8_4119);
and \g450607/U$3 ( \36739 , RIe205068_4347, \8359 );
nor \g450607/U$1 ( \36740 , \36738 , \36739 );
and \g454174/U$2 ( \36741 , \8313 , RIe1f8480_4202);
and \g454174/U$3 ( \36742 , RIe1ff0c8_4279, \8323 );
nor \g454174/U$1 ( \36743 , \36741 , \36742 );
not \g449530/U$3 ( \36744 , \36743 );
not \g449530/U$4 ( \36745 , \8347 );
and \g449530/U$2 ( \36746 , \36744 , \36745 );
and \g449530/U$5 ( \36747 , \8340 , RIe1d54d0_3804);
nor \g449530/U$1 ( \36748 , \36746 , \36747 );
and \g450606/U$2 ( \36749 , \8378 , RIe21b868_4603);
and \g450606/U$3 ( \36750 , RIe18ce10_2980, \8417 );
nor \g450606/U$1 ( \36751 , \36749 , \36750 );
nand \g447464/U$1 ( \36752 , \36737 , \36740 , \36748 , \36751 );
and \g444903/U$3 ( \36753 , \9010 , \36752 );
nor \g444903/U$1 ( \36754 , \36733 , \36753 );
and \g446516/U$2 ( \36755 , \9041 , RIe1a0910_3204);
and \g446516/U$3 ( \36756 , RIe1a3610_3236, \9043 );
nor \g446516/U$1 ( \36757 , \36755 , \36756 );
and \g446515/U$2 ( \36758 , \14956 , RIe1a6310_3268);
and \g446515/U$3 ( \36759 , RIe1a9010_3300, \14958 );
nor \g446515/U$1 ( \36760 , \36758 , \36759 );
and \g446517/U$2 ( \36761 , \13244 , RIe171480_2666);
and \g446517/U$3 ( \36762 , RIe1aee48_3367, \13246 );
nor \g446517/U$1 ( \36763 , \36761 , \36762 );
nand \g444550/U$1 ( \36764 , \36754 , \36757 , \36760 , \36763 );
and \g446510/U$2 ( \36765 , \8775 , RIe1ca0d0_3676);
and \g446510/U$3 ( \36766 , RIe1ccdd0_3708, \8777 );
nor \g446510/U$1 ( \36767 , \36765 , \36766 );
and \g445707/U$2 ( \36768 , RIe1cfad0_3740, \8488 );
and \g445707/U$3 ( \36769 , RIe1d27d0_3772, \8359 );
and \g448502/U$2 ( \36770 , RIe1c19d0_3580, \8317 );
and \g448502/U$3 ( \36771 , \8326 , RIe1c46d0_3612);
and \g448502/U$4 ( \36772 , RIe1ddbd0_3900, \8407 );
nor \g448502/U$1 ( \36773 , \36770 , \36771 , \36772 );
and \g450581/U$2 ( \36774 , \8335 , RIe1becd0_3548);
and \g450581/U$3 ( \36775 , RIe1c73d0_3644, \8340 );
nor \g450581/U$1 ( \36776 , \36774 , \36775 );
and \g450580/U$2 ( \36777 , \8404 , RIe1e35d0_3964);
and \g450580/U$3 ( \36778 , RIe1ebcd0_4060, \8351 );
nor \g450580/U$1 ( \36779 , \36777 , \36778 );
and \g454593/U$2 ( \36780 , \8313 , RIe1e62d0_3996);
and \g454593/U$3 ( \36781 , RIe1e8fd0_4028, \8323 );
nor \g454593/U$1 ( \36782 , \36780 , \36781 );
not \g449524/U$3 ( \36783 , \36782 );
not \g449524/U$4 ( \36784 , \8328 );
and \g449524/U$2 ( \36785 , \36783 , \36784 );
and \g449524/U$5 ( \36786 , \8417 , RIe1e08d0_3932);
nor \g449524/U$1 ( \36787 , \36785 , \36786 );
nand \g447459/U$1 ( \36788 , \36773 , \36776 , \36779 , \36787 );
nor \g445707/U$1 ( \36789 , \36768 , \36769 , \36788 );
not \g444846/U$3 ( \36790 , \36789 );
not \g444846/U$4 ( \36791 , \8477 );
and \g444846/U$2 ( \36792 , \36790 , \36791 );
and \g445710/U$2 ( \36793 , RIfc47b40_5838, \8351 );
and \g445710/U$3 ( \36794 , RIe1ee430_4088, \8335 );
and \g448505/U$2 ( \36795 , RIfcd58f0_7452, \8412 );
and \g448505/U$3 ( \36796 , \8407 , RIfcb7530_7108);
and \g448505/U$4 ( \36797 , RIfcbaaa0_7146, \8324 );
nor \g448505/U$1 ( \36798 , \36795 , \36796 , \36797 );
and \g450595/U$2 ( \36799 , \8356 , RIe1f3728_4147);
and \g450595/U$3 ( \36800 , RIf153488_5407, \8359 );
nor \g450595/U$1 ( \36801 , \36799 , \36800 );
and \g454166/U$2 ( \36802 , \8313 , RIfc51e60_5954);
and \g454166/U$3 ( \36803 , RIf151ca0_5390, \8323 );
nor \g454166/U$1 ( \36804 , \36802 , \36803 );
not \g449526/U$3 ( \36805 , \36804 );
not \g449526/U$4 ( \36806 , \8347 );
and \g449526/U$2 ( \36807 , \36805 , \36806 );
and \g449526/U$5 ( \36808 , \8340 , RIfc9aef8_6785);
nor \g449526/U$1 ( \36809 , \36807 , \36808 );
and \g450593/U$2 ( \36810 , \8378 , RIe1f5a50_4172);
and \g450593/U$3 ( \36811 , RIfc4ba88_5883, \8417 );
nor \g450593/U$1 ( \36812 , \36810 , \36811 );
nand \g447461/U$1 ( \36813 , \36798 , \36801 , \36809 , \36812 );
nor \g445710/U$1 ( \36814 , \36793 , \36794 , \36813 );
and \g450590/U$2 ( \36815 , \8319 , RIfc52130_5956);
and \g450590/U$3 ( \36816 , RIe1fa4d8_4225, \8404 );
nor \g450590/U$1 ( \36817 , \36815 , \36816 );
and \g450589/U$2 ( \36818 , \8371 , RIfc4b920_5882);
and \g450589/U$3 ( \36819 , RIfc84158_6525, \8330 );
nor \g450589/U$1 ( \36820 , \36818 , \36819 );
and \g444935/U$2 ( \36821 , \36814 , \36817 , \36820 );
nor \g444935/U$1 ( \36822 , \36821 , \8621 );
nor \g444846/U$1 ( \36823 , \36792 , \36822 );
and \g446512/U$2 ( \36824 , \10539 , RIe1d81d0_3836);
and \g446512/U$3 ( \36825 , RIe1daed0_3868, \10541 );
nor \g446512/U$1 ( \36826 , \36824 , \36825 );
nand \g444415/U$1 ( \36827 , \36767 , \36823 , \36826 );
and \g445703/U$2 ( \36828 , RIfc42140_5774, \8378 );
and \g445703/U$3 ( \36829 , RIfca3b98_6885, \8359 );
and \g448495/U$2 ( \36830 , RIfcc6008_7275, \8409 );
and \g448495/U$3 ( \36831 , \8373 , RIfca88f0_6940);
and \g448495/U$4 ( \36832 , RIfc5f858_6109, \8383 );
nor \g448495/U$1 ( \36833 , \36830 , \36831 , \36832 );
and \g450561/U$2 ( \36834 , \8335 , RIfc5f588_6107);
and \g450561/U$3 ( \36835 , RIfc9b330_6788, \8340 );
nor \g450561/U$1 ( \36836 , \36834 , \36835 );
and \g450560/U$2 ( \36837 , \8404 , RIe175f08_2719);
and \g450560/U$3 ( \36838 , RIfc6ccb0_6260, \8351 );
nor \g450560/U$1 ( \36839 , \36837 , \36838 );
and \g454149/U$2 ( \36840 , \8313 , RIfc42410_5776);
and \g454149/U$3 ( \36841 , RIf16f688_5727, \8323 );
nor \g454149/U$1 ( \36842 , \36840 , \36841 );
not \g454148/U$1 ( \36843 , \36842 );
and \g449517/U$2 ( \36844 , \36843 , \8316 );
and \g449517/U$3 ( \36845 , RIfc81020_6490, \8417 );
nor \g449517/U$1 ( \36846 , \36844 , \36845 );
nand \g448130/U$1 ( \36847 , \36833 , \36836 , \36839 , \36846 );
nor \g445703/U$1 ( \36848 , \36828 , \36829 , \36847 );
and \g450557/U$2 ( \36849 , \8356 , RIe173d48_2695);
and \g450557/U$3 ( \36850 , RIfc4ea58_5917, \8412 );
nor \g450557/U$1 ( \36851 , \36849 , \36850 );
and \g450556/U$2 ( \36852 , \8523 , RIfc984c8_6755);
and \g450556/U$3 ( \36853 , RIfc5ac68_6055, \8486 );
nor \g450556/U$1 ( \36854 , \36852 , \36853 );
and \g444931/U$2 ( \36855 , \36848 , \36851 , \36854 );
nor \g444931/U$1 ( \36856 , \36855 , \8558 );
and \g445704/U$2 ( \36857 , RIe19dc10_3172, \8351 );
and \g445704/U$3 ( \36858 , RIe17c010_2788, \8335 );
and \g448498/U$2 ( \36859 , RIe192810_3044, \8414 );
and \g448498/U$3 ( \36860 , \8409 , RIe195510_3076);
and \g448498/U$4 ( \36861 , RIe181a10_2852, \8326 );
nor \g448498/U$1 ( \36862 , \36859 , \36860 , \36861 );
and \g450573/U$2 ( \36863 , \8356 , RIe184710_2884);
and \g450573/U$3 ( \36864 , RIe18a110_2948, \8359 );
nor \g450573/U$1 ( \36865 , \36863 , \36864 );
and \g454153/U$2 ( \36866 , \8313 , RIfec12c0_8318);
and \g454153/U$3 ( \36867 , RIe187410_2916, \8323 );
nor \g454153/U$1 ( \36868 , \36866 , \36867 );
not \g449522/U$3 ( \36869 , \36868 );
not \g449522/U$4 ( \36870 , \8347 );
and \g449522/U$2 ( \36871 , \36869 , \36870 );
and \g449522/U$5 ( \36872 , \8340 , RIfc88370_6572);
nor \g449522/U$1 ( \36873 , \36871 , \36872 );
and \g450572/U$2 ( \36874 , \8378 , RIe18fb10_3012);
and \g450572/U$3 ( \36875 , RIfec1428_8319, \8417 );
nor \g450572/U$1 ( \36876 , \36874 , \36875 );
nand \g447457/U$1 ( \36877 , \36862 , \36865 , \36873 , \36876 );
nor \g445704/U$1 ( \36878 , \36857 , \36858 , \36877 );
and \g450567/U$2 ( \36879 , \8317 , RIe17ed10_2820);
and \g450567/U$3 ( \36880 , RIe198210_3108, \8404 );
nor \g450567/U$1 ( \36881 , \36879 , \36880 );
and \g450570/U$2 ( \36882 , \8373 , RIfec1590_8320);
and \g450570/U$3 ( \36883 , RIe19af10_3140, \8383 );
nor \g450570/U$1 ( \36884 , \36882 , \36883 );
and \g444932/U$2 ( \36885 , \36878 , \36881 , \36884 );
nor \g444932/U$1 ( \36886 , \36885 , \8589 );
or \g444307/U$1 ( \36887 , \36764 , \36827 , \36856 , \36886 );
and \g446498/U$2 ( \36888 , RIe215e68_4539, \8378 );
and \g446498/U$3 ( \36889 , RIfe87de0_7890, \8359 );
and \g448490/U$2 ( \36890 , RIe21e568_4635, \8409 );
and \g448490/U$3 ( \36891 , \8373 , RIf16bfb0_5688);
and \g448490/U$4 ( \36892 , RIe223f68_4699, \8383 );
nor \g448490/U$1 ( \36893 , \36890 , \36891 , \36892 );
and \g454129/U$2 ( \36894 , \8335 , RIe207d68_4379);
and \g454129/U$3 ( \36895 , RIfcdf670_7564, \8340 );
nor \g454129/U$1 ( \36896 , \36894 , \36895 );
and \g454127/U$2 ( \36897 , \8404 , RIe221268_4667);
and \g454127/U$3 ( \36898 , RIfe880b0_7892, \8351 );
nor \g454127/U$1 ( \36899 , \36897 , \36898 );
and \g454137/U$2 ( \36900 , \8313 , RIe20aa68_4411);
and \g454137/U$3 ( \36901 , RIe20d768_4443, \8323 );
nor \g454137/U$1 ( \36902 , \36900 , \36901 );
not \g454136/U$1 ( \36903 , \36902 );
and \g450535/U$2 ( \36904 , \36903 , \8316 );
and \g450535/U$3 ( \36905 , RIfc86cf0_6556, \8417 );
nor \g450535/U$1 ( \36906 , \36904 , \36905 );
nand \g448254/U$1 ( \36907 , \36893 , \36896 , \36899 , \36906 );
nor \g446498/U$1 ( \36908 , \36888 , \36889 , \36907 );
and \g454124/U$2 ( \36909 , \8356 , RIe210468_4475);
and \g454124/U$3 ( \36910 , RIe218b68_4571, \8414 );
nor \g454124/U$1 ( \36911 , \36909 , \36910 );
and \g454122/U$2 ( \36912 , \8531 , RIf1692b0_5656);
and \g454122/U$3 ( \36913 , RIe213168_4507, \8488 );
nor \g454122/U$1 ( \36914 , \36912 , \36913 );
and \g445501/U$2 ( \36915 , \36908 , \36911 , \36914 );
nor \g445501/U$1 ( \36916 , \36915 , \8368 );
and \g445700/U$2 ( \36917 , RIe202908_4319, \8373 );
and \g445700/U$3 ( \36918 , RIf1662e0_5622, \8383 );
and \g448493/U$2 ( \36919 , RIfccd790_7360, \8414 );
and \g448493/U$3 ( \36920 , \8409 , RIfc50ab0_5940);
and \g448493/U$4 ( \36921 , RIfc86480_6550, \8326 );
nor \g448493/U$1 ( \36922 , \36919 , \36920 , \36921 );
and \g450551/U$2 ( \36923 , \8356 , RIfe87f48_7891);
and \g450551/U$3 ( \36924 , RIf160610_5556, \8359 );
nor \g450551/U$1 ( \36925 , \36923 , \36924 );
and \g454145/U$2 ( \36926 , \8313 , RIfe87c78_7889);
and \g454145/U$3 ( \36927 , RIf15e720_5534, \8323 );
nor \g454145/U$1 ( \36928 , \36926 , \36927 );
not \g449514/U$3 ( \36929 , \36928 );
not \g449514/U$4 ( \36930 , \8347 );
and \g449514/U$2 ( \36931 , \36929 , \36930 );
and \g449514/U$5 ( \36932 , \8340 , RIfce7668_7655);
nor \g449514/U$1 ( \36933 , \36931 , \36932 );
and \g450550/U$2 ( \36934 , \8378 , RIfccd1f0_7356);
and \g450550/U$3 ( \36935 , RIfc58c10_6032, \8417 );
nor \g450550/U$1 ( \36936 , \36934 , \36935 );
nand \g447453/U$1 ( \36937 , \36922 , \36925 , \36933 , \36936 );
nor \g445700/U$1 ( \36938 , \36917 , \36918 , \36937 );
and \g450546/U$2 ( \36939 , \8335 , RIfcb01e0_7026);
and \g450546/U$3 ( \36940 , RIfca6460_6914, \8351 );
nor \g450546/U$1 ( \36941 , \36939 , \36940 );
and \g450547/U$2 ( \36942 , \8319 , RIfcd2218_7413);
and \g450547/U$3 ( \36943 , RIfe87b10_7888, \8404 );
nor \g450547/U$1 ( \36944 , \36942 , \36943 );
and \g444930/U$2 ( \36945 , \36938 , \36941 , \36944 );
nor \g444930/U$1 ( \36946 , \36945 , \8422 );
or \g444238/U$1 ( \36947 , \36887 , \36916 , \36946 );
_DC \g5f3f/U$1 ( \36948 , \36947 , \8654 );
and \g448697/U$2 ( \36949 , RIdec2de0_681, \16319 );
and \g448697/U$3 ( \36950 , \16328 , RIdec5ae0_713);
and \g448697/U$4 ( \36951 , RIdeab488_425, \16398 );
nor \g448697/U$1 ( \36952 , \36949 , \36950 , \36951 );
and \g454446/U$2 ( \36953 , \16317 , RIdebd3e0_617);
and \g454446/U$3 ( \36954 , RIfcb8d18_7125, \16325 );
nor \g454446/U$1 ( \36955 , \36953 , \36954 );
not \g449726/U$3 ( \36956 , \36955 );
not \g449726/U$4 ( \36957 , \16330 );
and \g449726/U$2 ( \36958 , \36956 , \36957 );
and \g449726/U$5 ( \36959 , \16341 , RIfce0750_7576);
nor \g449726/U$1 ( \36960 , \36958 , \36959 );
and \g451289/U$2 ( \36961 , \16377 , RIdec00e0_649);
and \g451289/U$3 ( \36962 , RIfc82268_6503, \16313 );
nor \g451289/U$1 ( \36963 , \36961 , \36962 );
and \g451290/U$2 ( \36964 , \16334 , RIdeb79e0_553);
and \g451290/U$3 ( \36965 , RIdeba6e0_585, \16380 );
nor \g451290/U$1 ( \36966 , \36964 , \36965 );
nand \g447276/U$1 ( \36967 , \36952 , \36960 , \36963 , \36966 );
and \g444703/U$2 ( \36968 , \36967 , \17938 );
and \g445864/U$2 ( \36969 , RIfc85670_6540, \16319 );
and \g445864/U$3 ( \36970 , RIfc81f98_6501, \16313 );
and \g448700/U$2 ( \36971 , RIfc7d7e0_6450, \16427 );
and \g448700/U$3 ( \36972 , \16448 , RIfcd2920_7418);
and \g448700/U$4 ( \36973 , RIe13f188_2095, \16485 );
nor \g448700/U$1 ( \36974 , \36971 , \36972 , \36973 );
and \g454184/U$2 ( \36975 , \16317 , RIdf338b0_1963);
and \g454184/U$3 ( \36976 , RIdf35ea8_1990, \16325 );
nor \g454184/U$1 ( \36977 , \36975 , \36976 );
not \g454183/U$1 ( \36978 , \36977 );
and \g449732/U$2 ( \36979 , \36978 , \16336 );
and \g449732/U$3 ( \36980 , RIe1414b0_2120, \16356 );
nor \g449732/U$1 ( \36981 , \36979 , \36980 );
and \g451304/U$2 ( \36982 , \16361 , RIdf2f800_1917);
and \g451304/U$3 ( \36983 , RIfe88920_7898, \16364 );
nor \g451304/U$1 ( \36984 , \36982 , \36983 );
and \g451301/U$2 ( \36985 , \16368 , RIfce5a48_7635);
and \g451301/U$3 ( \36986 , RIfc49760_5858, \16371 );
nor \g451301/U$1 ( \36987 , \36985 , \36986 );
nand \g448031/U$1 ( \36988 , \36974 , \36981 , \36984 , \36987 );
nor \g445864/U$1 ( \36989 , \36969 , \36970 , \36988 );
and \g451299/U$2 ( \36990 , \16377 , RIfcc4f28_7263);
and \g451299/U$3 ( \36991 , RIdf3d090_2071, \16380 );
nor \g451299/U$1 ( \36992 , \36990 , \36991 );
and \g451297/U$2 ( \36993 , \16334 , RIdf3aa98_2044);
and \g451297/U$3 ( \36994 , RIfc88208_6571, \16326 );
nor \g451297/U$1 ( \36995 , \36993 , \36994 );
and \g445049/U$2 ( \36996 , \36989 , \36992 , \36995 );
nor \g445049/U$1 ( \36997 , \36996 , \16393 );
nor \g444703/U$1 ( \36998 , \36968 , \36997 );
and \g446646/U$2 ( \36999 , \18457 , RIdeb1fe0_489);
and \g446646/U$3 ( \37000 , RIfcb9858_7133, \18459 );
nor \g446646/U$1 ( \37001 , \36999 , \37000 );
and \g446647/U$2 ( \37002 , \18462 , RIdeaf2e0_457);
and \g446647/U$3 ( \37003 , RIfc9efa8_6831, \18464 );
nor \g446647/U$1 ( \37004 , \37002 , \37003 );
and \g446648/U$2 ( \37005 , \18467 , RIde9e288_361);
and \g446648/U$3 ( \37006 , RIdea4b88_393, \18469 );
nor \g446648/U$1 ( \37007 , \37005 , \37006 );
nand \g444465/U$1 ( \37008 , \36998 , \37001 , \37004 , \37007 );
and \g453859/U$2 ( \37009 , \16313 , RIfe88a88_7899);
and \g453859/U$3 ( \37010 , RIe162de0_2502, \16321 );
nor \g453859/U$1 ( \37011 , \37009 , \37010 );
and \g445867/U$2 ( \37012 , RIe165ae0_2534, \16328 );
and \g445867/U$3 ( \37013 , RIe154ce0_2342, \16334 );
and \g448710/U$2 ( \37014 , RIe151fe0_2310, \16427 );
and \g448710/U$3 ( \37015 , \16448 , RIfc698a8_6223);
and \g448710/U$4 ( \37016 , RIe15d3e0_2438, \16485 );
nor \g448710/U$1 ( \37017 , \37014 , \37015 , \37016 );
and \g455408/U$2 ( \37018 , \16317 , RIe14c5e0_2246);
and \g455408/U$3 ( \37019 , RIfcc0338_7209, \16325 );
nor \g455408/U$1 ( \37020 , \37018 , \37019 );
not \g455407/U$1 ( \37021 , \37020 );
and \g449738/U$2 ( \37022 , \37021 , \16336 );
and \g449738/U$3 ( \37023 , RIfcc9140_7310, \16354 );
nor \g449738/U$1 ( \37024 , \37022 , \37023 );
and \g451320/U$2 ( \37025 , \16361 , RIe146be0_2182);
and \g451320/U$3 ( \37026 , RIe1498e0_2214, \16364 );
nor \g451320/U$1 ( \37027 , \37025 , \37026 );
and \g451318/U$2 ( \37028 , \16368 , RIe14f2e0_2278);
and \g451318/U$3 ( \37029 , RIee35098_5062, \16371 );
nor \g451318/U$1 ( \37030 , \37028 , \37029 );
nand \g448032/U$1 ( \37031 , \37017 , \37024 , \37027 , \37030 );
nor \g445867/U$1 ( \37032 , \37012 , \37013 , \37031 );
and \g451314/U$2 ( \37033 , \16377 , RIe1600e0_2470);
and \g451314/U$3 ( \37034 , RIe1579e0_2374, \16380 );
nor \g451314/U$1 ( \37035 , \37033 , \37034 );
nand \g445543/U$1 ( \37036 , \37011 , \37032 , \37035 );
and \g444738/U$2 ( \37037 , \37036 , \16390 );
and \g448704/U$2 ( \37038 , RIfe88d58_7901, \16344 );
and \g448704/U$3 ( \37039 , \16354 , RIfe89028_7903);
and \g448704/U$4 ( \37040 , RIe16bd50_2604, \16398 );
nor \g448704/U$1 ( \37041 , \37038 , \37039 , \37040 );
and \g455035/U$2 ( \37042 , \16317 , RIee1c138_4778);
and \g455035/U$3 ( \37043 , RIee1d0b0_4789, \16325 );
nor \g455035/U$1 ( \37044 , \37042 , \37043 );
not \g449734/U$3 ( \37045 , \37044 );
not \g449734/U$4 ( \37046 , \16311 );
and \g449734/U$2 ( \37047 , \37045 , \37046 );
and \g449734/U$5 ( \37048 , \16341 , RIfc4f868_5927);
nor \g449734/U$1 ( \37049 , \37047 , \37048 );
and \g451307/U$2 ( \37050 , \16377 , RIfc76d00_6374);
and \g451307/U$3 ( \37051 , RIfcd0e68_7399, \16313 );
nor \g451307/U$1 ( \37052 , \37050 , \37051 );
and \g451310/U$2 ( \37053 , \16334 , RIfe88bf0_7900);
and \g451310/U$3 ( \37054 , RIfe88ec0_7902, \16380 );
nor \g451310/U$1 ( \37055 , \37053 , \37054 );
nand \g447277/U$1 ( \37056 , \37041 , \37049 , \37052 , \37055 );
and \g444738/U$3 ( \37057 , \17998 , \37056 );
nor \g444738/U$1 ( \37058 , \37037 , \37057 );
and \g446656/U$2 ( \37059 , \18523 , RIfcde590_7552);
and \g446656/U$3 ( \37060 , RIfcda7b0_7508, \18525 );
nor \g446656/U$1 ( \37061 , \37059 , \37060 );
and \g446654/U$2 ( \37062 , \18528 , RIfc52dd8_5965);
and \g446654/U$3 ( \37063 , RIfc4d810_5904, \18530 );
nor \g446654/U$1 ( \37064 , \37062 , \37063 );
and \g446657/U$2 ( \37065 , \18533 , RIe1683a8_2563);
and \g446657/U$3 ( \37066 , RIfc68930_6212, \18535 );
nor \g446657/U$1 ( \37067 , \37065 , \37066 );
nand \g444573/U$1 ( \37068 , \37058 , \37061 , \37064 , \37067 );
and \g445855/U$2 ( \37069 , RIfcad918_6997, \16448 );
and \g445855/U$3 ( \37070 , RIdf19870_1667, \16361 );
and \g448639/U$2 ( \37071 , RIee2a670_4941, \16321 );
and \g448639/U$3 ( \37072 , \16328 , RIee2bfc0_4959);
and \g448639/U$4 ( \37073 , RIdf1ff18_1740, \16337 );
nor \g448639/U$1 ( \37074 , \37071 , \37072 , \37073 );
and \g454996/U$2 ( \37075 , \16317 , RIdf28618_1836);
and \g454996/U$3 ( \37076 , RIdf2a7d8_1860, \16325 );
nor \g454996/U$1 ( \37077 , \37075 , \37076 );
not \g449718/U$3 ( \37078 , \37077 );
not \g449718/U$4 ( \37079 , \16330 );
and \g449718/U$2 ( \37080 , \37078 , \37079 );
and \g449718/U$5 ( \37081 , \16341 , RIfc60938_6121);
nor \g449718/U$1 ( \37082 , \37080 , \37081 );
and \g451263/U$2 ( \37083 , \16377 , RIee27f10_4913);
and \g451263/U$3 ( \37084 , RIee29158_4926, \16313 );
nor \g451263/U$1 ( \37085 , \37083 , \37084 );
and \g451264/U$2 ( \37086 , \16334 , RIdf24dd8_1796);
and \g451264/U$3 ( \37087 , RIdf26890_1815, \16380 );
nor \g451264/U$1 ( \37088 , \37086 , \37087 );
nand \g447273/U$1 ( \37089 , \37074 , \37082 , \37085 , \37088 );
nor \g445855/U$1 ( \37090 , \37069 , \37070 , \37089 );
and \g451261/U$2 ( \37091 , \16364 , RIfcba500_7142);
and \g451261/U$3 ( \37092 , RIfc623f0_6140, \16368 );
nor \g451261/U$1 ( \37093 , \37091 , \37092 );
and \g451204/U$2 ( \37094 , \16371 , RIfc63368_6151);
and \g451204/U$3 ( \37095 , RIfc69fb0_6228, \16427 );
nor \g451204/U$1 ( \37096 , \37094 , \37095 );
and \g445044/U$2 ( \37097 , \37090 , \37093 , \37096 );
nor \g445044/U$1 ( \37098 , \37097 , \16480 );
and \g445857/U$2 ( \37099 , RIdefe1b0_1355, \16448 );
and \g445857/U$3 ( \37100 , RIdeea6b0_1131, \16361 );
and \g448694/U$2 ( \37101 , RIdf095b0_1483, \16485 );
and \g448694/U$3 ( \37102 , \16356 , RIdf0c2b0_1515);
and \g448694/U$4 ( \37103 , RIdef00b0_1195, \16398 );
nor \g448694/U$1 ( \37104 , \37101 , \37102 , \37103 );
and \g454993/U$2 ( \37105 , \16317 , RIdf149b0_1611);
and \g454993/U$3 ( \37106 , RIdf176b0_1643, \16325 );
nor \g454993/U$1 ( \37107 , \37105 , \37106 );
not \g449723/U$3 ( \37108 , \37107 );
not \g449723/U$4 ( \37109 , \16311 );
and \g449723/U$2 ( \37110 , \37108 , \37109 );
and \g449723/U$5 ( \37111 , \16339 , RIdef2db0_1227);
nor \g449723/U$1 ( \37112 , \37110 , \37111 );
and \g451275/U$2 ( \37113 , \16377 , RIdf0efb0_1547);
and \g451275/U$3 ( \37114 , RIdf11cb0_1579, \16313 );
nor \g451275/U$1 ( \37115 , \37113 , \37114 );
and \g451278/U$2 ( \37116 , \16334 , RIdf03bb0_1419);
and \g451278/U$3 ( \37117 , RIdf068b0_1451, \16380 );
nor \g451278/U$1 ( \37118 , \37116 , \37117 );
nand \g447275/U$1 ( \37119 , \37104 , \37112 , \37115 , \37118 );
nor \g445857/U$1 ( \37120 , \37099 , \37100 , \37119 );
and \g451272/U$2 ( \37121 , \16364 , RIdeed3b0_1163);
and \g451272/U$3 ( \37122 , RIdef5ab0_1259, \16368 );
nor \g451272/U$1 ( \37123 , \37121 , \37122 );
and \g451270/U$2 ( \37124 , \16371 , RIdef87b0_1291);
and \g451270/U$3 ( \37125 , RIdefb4b0_1323, \16427 );
nor \g451270/U$1 ( \37126 , \37124 , \37125 );
and \g445046/U$2 ( \37127 , \37120 , \37123 , \37126 );
nor \g445046/U$1 ( \37128 , \37127 , \16555 );
or \g444379/U$1 ( \37129 , \37008 , \37068 , \37098 , \37128 );
and \g445848/U$2 ( \37130 , RIfc84590_6528, \16448 );
and \g445848/U$3 ( \37131 , RIded34d8_868, \16361 );
and \g448682/U$2 ( \37132 , RIdee31f8_1048, \16485 );
and \g448682/U$3 ( \37133 , \16356 , RIdee4f80_1069);
and \g448682/U$4 ( \37134 , RIded7858_916, \16398 );
nor \g448682/U$1 ( \37135 , \37132 , \37133 , \37134 );
and \g454526/U$2 ( \37136 , \16317 , RIfc69a10_6224);
and \g454526/U$3 ( \37137 , RIfcc9848_7315, \16325 );
nor \g454526/U$1 ( \37138 , \37136 , \37137 );
not \g449710/U$3 ( \37139 , \37138 );
not \g449710/U$4 ( \37140 , \16311 );
and \g449710/U$2 ( \37141 , \37139 , \37140 );
and \g449710/U$5 ( \37142 , \16341 , RIded9e50_943);
nor \g449710/U$1 ( \37143 , \37141 , \37142 );
and \g451238/U$2 ( \37144 , \16377 , RIfccbfa8_7343);
and \g451238/U$3 ( \37145 , RIfcacc70_6988, \16313 );
nor \g451238/U$1 ( \37146 , \37144 , \37145 );
and \g451239/U$2 ( \37147 , \16334 , RIdedee78_1000);
and \g451239/U$3 ( \37148 , RIdee1038_1024, \16380 );
nor \g451239/U$1 ( \37149 , \37147 , \37148 );
nand \g447271/U$1 ( \37150 , \37135 , \37143 , \37146 , \37149 );
nor \g445848/U$1 ( \37151 , \37130 , \37131 , \37150 );
and \g451235/U$2 ( \37152 , \16364 , RIfe887b8_7897);
and \g451235/U$3 ( \37153 , RIfc47168_5831, \16368 );
nor \g451235/U$1 ( \37154 , \37152 , \37153 );
and \g451231/U$2 ( \37155 , \16371 , RIee21b38_4842);
and \g451231/U$3 ( \37156 , RIfc9bba0_6794, \16427 );
nor \g451231/U$1 ( \37157 , \37155 , \37156 );
and \g445036/U$2 ( \37158 , \37151 , \37154 , \37157 );
nor \g445036/U$1 ( \37159 , \37158 , \16909 );
and \g445851/U$2 ( \37160 , RIe143ee0_2150, \16448 );
and \g445851/U$3 ( \37161 , RIde7d8d0_202, \16361 );
and \g448687/U$2 ( \37162 , RIde97988_329, \16344 );
and \g448687/U$3 ( \37163 , \16354 , RIdeb4ce0_521);
and \g448687/U$4 ( \37164 , RIdee79b0_1099, \16398 );
nor \g448687/U$1 ( \37165 , \37162 , \37163 , \37164 );
and \g454455/U$2 ( \37166 , \16317 , RIdece1e0_809);
and \g454455/U$3 ( \37167 , RIded0ee0_841, \16325 );
nor \g454455/U$1 ( \37168 , \37166 , \37167 );
not \g449715/U$3 ( \37169 , \37168 );
not \g449715/U$4 ( \37170 , \16311 );
and \g449715/U$2 ( \37171 , \37169 , \37170 );
and \g449715/U$5 ( \37172 , \16339 , RIdf00eb0_1387);
nor \g449715/U$1 ( \37173 , \37171 , \37172 );
and \g451250/U$2 ( \37174 , \16377 , RIdec87e0_745);
and \g451250/U$3 ( \37175 , RIdecb4e0_777, \16313 );
nor \g451250/U$1 ( \37176 , \37174 , \37175 );
and \g451252/U$2 ( \37177 , \16334 , RIe15a6e0_2406);
and \g451252/U$3 ( \37178 , RIe16e8e8_2635, \16380 );
nor \g451252/U$1 ( \37179 , \37177 , \37178 );
nand \g447272/U$1 ( \37180 , \37165 , \37173 , \37176 , \37179 );
nor \g445851/U$1 ( \37181 , \37160 , \37161 , \37180 );
and \g451247/U$2 ( \37182 , \16364 , RIdedc718_972);
and \g451247/U$3 ( \37183 , RIdf1d7b8_1712, \16368 );
nor \g451247/U$1 ( \37184 , \37182 , \37183 );
and \g451246/U$2 ( \37185 , \16371 , RIdf2cf38_1888);
and \g451246/U$3 ( \37186 , RIdf388d8_2020, \16427 );
nor \g451246/U$1 ( \37187 , \37185 , \37186 );
and \g445039/U$2 ( \37188 , \37181 , \37184 , \37187 );
nor \g445039/U$1 ( \37189 , \37188 , \16586 );
or \g444166/U$1 ( \37190 , \37129 , \37159 , \37189 );
_DC \g5fc4/U$1 ( \37191 , \37190 , \16652 );
and \g446675/U$2 ( \37192 , \8969 , RIe1b7818_3465);
and \g446675/U$3 ( \37193 , RIe1b9870_3488, \8971 );
nor \g446675/U$1 ( \37194 , \37192 , \37193 );
and \g445882/U$2 ( \37195 , RIfcb8a48_7123, \8351 );
and \g445882/U$3 ( \37196 , RIfcb84a8_7119, \8383 );
and \g448728/U$2 ( \37197 , RIfeac140_8274, \8414 );
and \g448728/U$3 ( \37198 , \8409 , RIfc9e198_6821);
and \g448728/U$4 ( \37199 , RIfc82ad8_6509, \8324 );
nor \g448728/U$1 ( \37200 , \37197 , \37198 , \37199 );
and \g451380/U$2 ( \37201 , \8356 , RIe1b1008_3391);
and \g451380/U$3 ( \37202 , RIfc518c0_5950, \8359 );
nor \g451380/U$1 ( \37203 , \37201 , \37202 );
and \g454498/U$2 ( \37204 , \8313 , RIfe884e8_7895);
and \g454498/U$3 ( \37205 , RIfc838e8_6519, \8323 );
nor \g454498/U$1 ( \37206 , \37204 , \37205 );
not \g449758/U$3 ( \37207 , \37206 );
not \g449758/U$4 ( \37208 , \8347 );
and \g449758/U$2 ( \37209 , \37207 , \37208 );
and \g449758/U$5 ( \37210 , \8340 , RIfcc5900_7270);
nor \g449758/U$1 ( \37211 , \37209 , \37210 );
and \g451378/U$2 ( \37212 , \8378 , RIe1b42a8_3427);
and \g451378/U$3 ( \37213 , RIfc85940_6542, \8417 );
nor \g451378/U$1 ( \37214 , \37212 , \37213 );
nand \g447577/U$1 ( \37215 , \37200 , \37203 , \37211 , \37214 );
nor \g445882/U$1 ( \37216 , \37195 , \37196 , \37215 );
not \g444814/U$3 ( \37217 , \37216 );
not \g444814/U$4 ( \37218 , \8481 );
and \g444814/U$2 ( \37219 , \37217 , \37218 );
and \g445885/U$2 ( \37220 , RIe1e6438_3997, \8371 );
and \g445885/U$3 ( \37221 , RIe1e9138_4029, \8383 );
and \g448733/U$2 ( \37222 , RIe1db038_3869, \8414 );
and \g448733/U$3 ( \37223 , \8409 , RIe1ddd38_3901);
and \g448733/U$4 ( \37224 , RIe1c4838_3613, \8326 );
nor \g448733/U$1 ( \37225 , \37222 , \37223 , \37224 );
and \g451393/U$2 ( \37226 , \8356 , RIe1ca238_3677);
and \g451393/U$3 ( \37227 , RIe1d2938_3773, \8359 );
nor \g451393/U$1 ( \37228 , \37226 , \37227 );
and \g454622/U$2 ( \37229 , \8313 , RIe1ccf38_3709);
and \g454622/U$3 ( \37230 , RIe1cfc38_3741, \8323 );
nor \g454622/U$1 ( \37231 , \37229 , \37230 );
not \g449762/U$3 ( \37232 , \37231 );
not \g449762/U$4 ( \37233 , \8347 );
and \g449762/U$2 ( \37234 , \37232 , \37233 );
and \g449762/U$5 ( \37235 , \8340 , RIe1c7538_3645);
nor \g449762/U$1 ( \37236 , \37234 , \37235 );
and \g451390/U$2 ( \37237 , \8378 , RIe1d8338_3837);
and \g451390/U$3 ( \37238 , RIe1e0a38_3933, \8417 );
nor \g451390/U$1 ( \37239 , \37237 , \37238 );
nand \g447579/U$1 ( \37240 , \37225 , \37228 , \37236 , \37239 );
nor \g445885/U$1 ( \37241 , \37220 , \37221 , \37240 );
and \g451386/U$2 ( \37242 , \8335 , RIe1bee38_3549);
and \g451386/U$3 ( \37243 , RIe1ebe38_4061, \8351 );
nor \g451386/U$1 ( \37244 , \37242 , \37243 );
and \g451387/U$2 ( \37245 , \8319 , RIe1c1b38_3581);
and \g451387/U$3 ( \37246 , RIe1e3738_3965, \8404 );
nor \g451387/U$1 ( \37247 , \37245 , \37246 );
and \g445063/U$2 ( \37248 , \37241 , \37244 , \37247 );
nor \g445063/U$1 ( \37249 , \37248 , \8477 );
nor \g444814/U$1 ( \37250 , \37219 , \37249 );
and \g446674/U$2 ( \37251 , \8509 , RIfe88650_7896);
and \g446674/U$3 ( \37252 , RIe1ac9b8_3341, \8511 );
nor \g446674/U$1 ( \37253 , \37251 , \37252 );
nand \g444422/U$1 ( \37254 , \37194 , \37250 , \37253 );
and \g448688/U$2 ( \37255 , RIe20abd0_4412, \8317 );
and \g448688/U$3 ( \37256 , \8324 , RIe20d8d0_4444);
and \g448688/U$4 ( \37257 , RIe21e6d0_4636, \8407 );
nor \g448688/U$1 ( \37258 , \37255 , \37256 , \37257 );
and \g451401/U$2 ( \37259 , \8335 , RIe207ed0_4380);
and \g451401/U$3 ( \37260 , RIfc97988_6747, \8340 );
nor \g451401/U$1 ( \37261 , \37259 , \37260 );
and \g451399/U$2 ( \37262 , \8404 , RIe2213d0_4668);
and \g451399/U$3 ( \37263 , RIfc40a48_5761, \8351 );
nor \g451399/U$1 ( \37264 , \37262 , \37263 );
and \g454185/U$2 ( \37265 , \8313 , RIfc85508_6539);
and \g454185/U$3 ( \37266 , RIe2240d0_4700, \8323 );
nor \g454185/U$1 ( \37267 , \37265 , \37266 );
not \g449765/U$3 ( \37268 , \37267 );
not \g449765/U$4 ( \37269 , \8328 );
and \g449765/U$2 ( \37270 , \37268 , \37269 );
and \g449765/U$5 ( \37271 , \8417 , RIfc9ba38_6793);
nor \g449765/U$1 ( \37272 , \37270 , \37271 );
nand \g447583/U$1 ( \37273 , \37258 , \37261 , \37264 , \37272 );
and \g444764/U$2 ( \37274 , \37273 , \8369 );
and \g445890/U$2 ( \37275 , RIe202a70_4320, \8373 );
and \g445890/U$3 ( \37276 , RIfcddbb8_7545, \8330 );
and \g448739/U$2 ( \37277 , RIfc71468_6311, \8414 );
and \g448739/U$3 ( \37278 , \8409 , RIfcaf100_7014);
and \g448739/U$4 ( \37279 , RIfcdd1e0_7538, \8326 );
nor \g448739/U$1 ( \37280 , \37277 , \37278 , \37279 );
and \g451414/U$2 ( \37281 , \8356 , RIe1fbcc0_4242);
and \g451414/U$3 ( \37282 , RIfcdda50_7544, \8359 );
nor \g451414/U$1 ( \37283 , \37281 , \37282 );
and \g454513/U$2 ( \37284 , \8313 , RIe1fcf08_4255);
and \g454513/U$3 ( \37285 , RIfca8620_6938, \8323 );
nor \g454513/U$1 ( \37286 , \37284 , \37285 );
not \g449768/U$3 ( \37287 , \37286 );
not \g449768/U$4 ( \37288 , \8347 );
and \g449768/U$2 ( \37289 , \37287 , \37288 );
and \g449768/U$5 ( \37290 , \8340 , RIfc6c008_6251);
nor \g449768/U$1 ( \37291 , \37289 , \37290 );
and \g451413/U$2 ( \37292 , \8378 , RIfcdcad8_7533);
and \g451413/U$3 ( \37293 , RIfc73d30_6340, \8417 );
nor \g451413/U$1 ( \37294 , \37292 , \37293 );
nand \g447586/U$1 ( \37295 , \37280 , \37283 , \37291 , \37294 );
nor \g445890/U$1 ( \37296 , \37275 , \37276 , \37295 );
and \g451409/U$2 ( \37297 , \8335 , RIfca92c8_6947);
and \g451409/U$3 ( \37298 , RIfceb5b0_7700, \8351 );
nor \g451409/U$1 ( \37299 , \37297 , \37298 );
and \g451410/U$2 ( \37300 , \8319 , RIfca9700_6950);
and \g451410/U$3 ( \37301 , RIe200e50_4300, \8404 );
nor \g451410/U$1 ( \37302 , \37300 , \37301 );
and \g445067/U$2 ( \37303 , \37296 , \37299 , \37302 );
nor \g445067/U$1 ( \37304 , \37303 , \8422 );
nor \g444764/U$1 ( \37305 , \37274 , \37304 );
and \g446681/U$2 ( \37306 , \8438 , RIe215fd0_4540);
and \g446681/U$3 ( \37307 , RIe218cd0_4572, \8440 );
nor \g446681/U$1 ( \37308 , \37306 , \37307 );
and \g446679/U$2 ( \37309 , \12506 , RIe2132d0_4508);
and \g446679/U$3 ( \37310 , RIfc52c70_5964, \12508 );
nor \g446679/U$1 ( \37311 , \37309 , \37310 );
and \g446682/U$2 ( \37312 , \8717 , RIe2105d0_4476);
and \g446682/U$3 ( \37313 , RIfca3760_6882, \8719 );
nor \g446682/U$1 ( \37314 , \37312 , \37313 );
nand \g444471/U$1 ( \37315 , \37305 , \37308 , \37311 , \37314 );
and \g445876/U$2 ( \37316 , RIfcce708_7371, \8414 );
and \g445876/U$3 ( \37317 , RIe1f3890_4148, \8356 );
and \g448720/U$2 ( \37318 , RIfc53918_5973, \8407 );
and \g448720/U$3 ( \37319 , \8373 , RIfc6f410_6288);
and \g448720/U$4 ( \37320 , RIfc6ba68_6247, \8383 );
nor \g448720/U$1 ( \37321 , \37318 , \37319 , \37320 );
and \g451354/U$2 ( \37322 , \8335 , RIe1ee598_4089);
and \g451354/U$3 ( \37323 , RIf14fc48_5367, \8340 );
nor \g451354/U$1 ( \37324 , \37322 , \37323 );
and \g451352/U$2 ( \37325 , \8404 , RIe1fa640_4226);
and \g451352/U$3 ( \37326 , RIfcce5a0_7370, \8351 );
nor \g451352/U$1 ( \37327 , \37325 , \37326 );
and \g454885/U$2 ( \37328 , \8313 , RIfc73e98_6341);
and \g454885/U$3 ( \37329 , RIfc72c50_6328, \8323 );
nor \g454885/U$1 ( \37330 , \37328 , \37329 );
not \g454884/U$1 ( \37331 , \37330 );
and \g449750/U$2 ( \37332 , \37331 , \8316 );
and \g449750/U$3 ( \37333 , RIfcce000_7366, \8417 );
nor \g449750/U$1 ( \37334 , \37332 , \37333 );
nand \g448155/U$1 ( \37335 , \37321 , \37324 , \37327 , \37334 );
nor \g445876/U$1 ( \37336 , \37316 , \37317 , \37335 );
and \g451349/U$2 ( \37337 , \8378 , RIe1f5bb8_4173);
and \g451349/U$3 ( \37338 , RIf1535f0_5408, \8359 );
nor \g451349/U$1 ( \37339 , \37337 , \37338 );
and \g452757/U$2 ( \37340 , \8531 , RIfc72db8_6329);
and \g452757/U$3 ( \37341 , RIf151e08_5391, \8488 );
nor \g452757/U$1 ( \37342 , \37340 , \37341 );
and \g445058/U$2 ( \37343 , \37336 , \37339 , \37342 );
nor \g445058/U$1 ( \37344 , \37343 , \8621 );
and \g445878/U$2 ( \37345 , RIe1a3778_3237, \8373 );
and \g445878/U$3 ( \37346 , RIe1a6478_3269, \8383 );
and \g448725/U$2 ( \37347 , RIe1bc138_3517, \8324 );
and \g448725/U$3 ( \37348 , \8523 , RIe1f85e8_4203);
and \g448725/U$4 ( \37349 , RIe1ff230_4280, \8488 );
nor \g448725/U$1 ( \37350 , \37347 , \37348 , \37349 );
and \g451368/U$2 ( \37351 , \8356 , RIe1f1130_4120);
and \g451368/U$3 ( \37352 , RIe2051d0_4348, \8359 );
nor \g451368/U$1 ( \37353 , \37351 , \37352 );
and \g454752/U$2 ( \37354 , \8313 , RIe226dd0_4732);
and \g454752/U$3 ( \37355 , RIe179478_2757, \8323 );
nor \g454752/U$1 ( \37356 , \37354 , \37355 );
not \g449754/U$3 ( \37357 , \37356 );
not \g449754/U$4 ( \37358 , \8376 );
and \g449754/U$2 ( \37359 , \37357 , \37358 );
and \g449754/U$5 ( \37360 , \8340 , RIe1d5638_3805);
nor \g449754/U$1 ( \37361 , \37359 , \37360 );
and \g451364/U$2 ( \37362 , \8378 , RIe21b9d0_4604);
and \g451364/U$3 ( \37363 , RIe18cf78_2981, \8417 );
nor \g451364/U$1 ( \37364 , \37362 , \37363 );
nand \g447576/U$1 ( \37365 , \37350 , \37353 , \37361 , \37364 );
nor \g445878/U$1 ( \37366 , \37345 , \37346 , \37365 );
and \g452435/U$2 ( \37367 , \8335 , RIe1715e8_2667);
and \g452435/U$3 ( \37368 , RIe1a9178_3301, \8351 );
nor \g452435/U$1 ( \37369 , \37367 , \37368 );
and \g451360/U$2 ( \37370 , \8317 , RIe1aefb0_3368);
and \g451360/U$3 ( \37371 , RIe1a0a78_3205, \8404 );
nor \g451360/U$1 ( \37372 , \37370 , \37371 );
and \g445059/U$2 ( \37373 , \37366 , \37369 , \37372 );
nor \g445059/U$1 ( \37374 , \37373 , \8651 );
or \g444291/U$1 ( \37375 , \37254 , \37315 , \37344 , \37374 );
and \g445872/U$2 ( \37376 , RIe19dd78_3173, \8351 );
and \g445872/U$3 ( \37377 , RIe198378_3109, \8404 );
and \g448712/U$2 ( \37378 , RIe192978_3045, \8412 );
and \g448712/U$3 ( \37379 , \8407 , RIe195678_3077);
and \g448712/U$4 ( \37380 , RIe181b78_2853, \8324 );
nor \g448712/U$1 ( \37381 , \37378 , \37379 , \37380 );
and \g451335/U$2 ( \37382 , \8356 , RIe184878_2885);
and \g451335/U$3 ( \37383 , RIe18a278_2949, \8359 );
nor \g451335/U$1 ( \37384 , \37382 , \37383 );
and \g454469/U$2 ( \37385 , \8313 , RIfcba230_7140);
and \g454469/U$3 ( \37386 , RIe187578_2917, \8323 );
nor \g454469/U$1 ( \37387 , \37385 , \37386 );
not \g449741/U$3 ( \37388 , \37387 );
not \g449741/U$4 ( \37389 , \8347 );
and \g449741/U$2 ( \37390 , \37388 , \37389 );
and \g449741/U$5 ( \37391 , \8340 , RIf142d90_5220);
nor \g449741/U$1 ( \37392 , \37390 , \37391 );
and \g451332/U$2 ( \37393 , \8378 , RIe18fc78_3013);
and \g451332/U$3 ( \37394 , RIfca35f8_6881, \8417 );
nor \g451332/U$1 ( \37395 , \37393 , \37394 );
nand \g447574/U$1 ( \37396 , \37381 , \37384 , \37392 , \37395 );
nor \g445872/U$1 ( \37397 , \37376 , \37377 , \37396 );
and \g451328/U$2 ( \37398 , \8335 , RIe17c178_2789);
and \g451328/U$3 ( \37399 , RIe19b078_3141, \8383 );
nor \g451328/U$1 ( \37400 , \37398 , \37399 );
and \g451326/U$2 ( \37401 , \8317 , RIe17ee78_2821);
and \g451326/U$3 ( \37402 , RIfca1438_6857, \8373 );
nor \g451326/U$1 ( \37403 , \37401 , \37402 );
and \g445053/U$2 ( \37404 , \37397 , \37400 , \37403 );
nor \g445053/U$1 ( \37405 , \37404 , \8589 );
and \g445874/U$2 ( \37406 , RIfc4ccd0_5896, \8373 );
and \g445874/U$3 ( \37407 , RIfc9bd08_6795, \8383 );
and \g448717/U$2 ( \37408 , RIfcc4c58_7261, \8414 );
and \g448717/U$3 ( \37409 , \8407 , RIfc87b00_6566);
and \g448717/U$4 ( \37410 , RIfc4e080_5910, \8326 );
nor \g448717/U$1 ( \37411 , \37408 , \37409 , \37410 );
and \g451346/U$2 ( \37412 , \8356 , RIe173eb0_2696);
and \g451346/U$3 ( \37413 , RIfc4f598_5925, \8359 );
nor \g451346/U$1 ( \37414 , \37412 , \37413 );
and \g455067/U$2 ( \37415 , \8313 , RIfc4dae0_5906);
and \g455067/U$3 ( \37416 , RIfc876c8_6563, \8323 );
nor \g455067/U$1 ( \37417 , \37415 , \37416 );
not \g449745/U$3 ( \37418 , \37417 );
not \g449745/U$4 ( \37419 , \8347 );
and \g449745/U$2 ( \37420 , \37418 , \37419 );
and \g449745/U$5 ( \37421 , \8340 , RIfcb9420_7130);
nor \g449745/U$1 ( \37422 , \37420 , \37421 );
and \g451344/U$2 ( \37423 , \8378 , RIfc4fca0_5930);
and \g451344/U$3 ( \37424 , RIfc87c68_6567, \8417 );
nor \g451344/U$1 ( \37425 , \37423 , \37424 );
nand \g447575/U$1 ( \37426 , \37411 , \37414 , \37422 , \37425 );
nor \g445874/U$1 ( \37427 , \37406 , \37407 , \37426 );
and \g451340/U$2 ( \37428 , \8335 , RIfc9d388_6811);
and \g451340/U$3 ( \37429 , RIfc9be70_6796, \8351 );
nor \g451340/U$1 ( \37430 , \37428 , \37429 );
and \g451342/U$2 ( \37431 , \8317 , RIfc4e350_5912);
and \g451342/U$3 ( \37432 , RIe176070_2720, \8404 );
nor \g451342/U$1 ( \37433 , \37431 , \37432 );
and \g445055/U$2 ( \37434 , \37427 , \37430 , \37433 );
nor \g445055/U$1 ( \37435 , \37434 , \8558 );
or \g444233/U$1 ( \37436 , \37375 , \37405 , \37435 );
_DC \g6048/U$1 ( \37437 , \37436 , \8654 );
and \g452652/U$2 ( \37438 , \16380 , RIe157b48_2375);
and \g452652/U$3 ( \37439 , RIe15d548_2439, \16485 );
nor \g452652/U$1 ( \37440 , \37438 , \37439 );
and \g445911/U$2 ( \37441 , RIfc4e8f0_5916, \16356 );
and \g445911/U$3 ( \37442 , RIe14f448_2279, \16368 );
and \g448765/U$2 ( \37443 , RIe152148_2311, \16427 );
and \g448765/U$3 ( \37444 , \16398 , RIe14c748_2247);
and \g448765/U$4 ( \37445 , RIfc865e8_6551, \16341 );
nor \g448765/U$1 ( \37446 , \37443 , \37444 , \37445 );
and \g451497/U$2 ( \37447 , \16361 , RIe146d48_2183);
and \g451497/U$3 ( \37448 , RIe149a48_2215, \16364 );
nor \g451497/U$1 ( \37449 , \37447 , \37448 );
and \g451495/U$2 ( \37450 , \16377 , RIe160248_2471);
and \g451495/U$3 ( \37451 , RIfc4f9d0_5928, \16313 );
nor \g451495/U$1 ( \37452 , \37450 , \37451 );
and \g454861/U$2 ( \37453 , \16317 , RIe162f48_2503);
and \g454861/U$3 ( \37454 , RIe165c48_2535, \16325 );
nor \g454861/U$1 ( \37455 , \37453 , \37454 );
not \g449793/U$3 ( \37456 , \37455 );
not \g449793/U$4 ( \37457 , \16311 );
and \g449793/U$2 ( \37458 , \37456 , \37457 );
and \g449793/U$5 ( \37459 , \16448 , RIfc4e1e8_5911);
nor \g449793/U$1 ( \37460 , \37458 , \37459 );
nand \g447604/U$1 ( \37461 , \37446 , \37449 , \37452 , \37460 );
nor \g445911/U$1 ( \37462 , \37441 , \37442 , \37461 );
and \g451492/U$2 ( \37463 , \16334 , RIe154e48_2343);
and \g451492/U$3 ( \37464 , RIfc868b8_6553, \16371 );
nor \g451492/U$1 ( \37465 , \37463 , \37464 );
nand \g445554/U$1 ( \37466 , \37440 , \37462 , \37465 );
and \g444740/U$2 ( \37467 , \37466 , \16390 );
and \g448761/U$2 ( \37468 , RIfcb1b30_7044, \16427 );
and \g448761/U$3 ( \37469 , \16432 , RIfcdf508_7563);
and \g448761/U$4 ( \37470 , RIfc5b0a0_6058, \16321 );
nor \g448761/U$1 ( \37471 , \37468 , \37469 , \37470 );
and \g451487/U$2 ( \37472 , \16368 , RIfcb16f8_7041);
and \g451487/U$3 ( \37473 , RIfc5ccc0_6078, \16371 );
nor \g451487/U$1 ( \37474 , \37472 , \37473 );
and \g455006/U$2 ( \37475 , \16317 , RIde8e5e0_284);
and \g455006/U$3 ( \37476 , RIfea92d8_8241, \16325 );
nor \g455006/U$1 ( \37477 , \37475 , \37476 );
not \g449790/U$3 ( \37478 , \37477 );
not \g449790/U$4 ( \37479 , \16330 );
and \g449790/U$2 ( \37480 , \37478 , \37479 );
and \g449790/U$5 ( \37481 , \16328 , RIfc41e70_5772);
nor \g449790/U$1 ( \37482 , \37480 , \37481 );
and \g451485/U$2 ( \37483 , \16334 , RIfea0bd8_8173);
and \g451485/U$3 ( \37484 , RIfea0d40_8174, \16380 );
nor \g451485/U$1 ( \37485 , \37483 , \37484 );
nand \g447603/U$1 ( \37486 , \37471 , \37474 , \37482 , \37485 );
and \g444740/U$3 ( \37487 , \17998 , \37486 );
nor \g444740/U$1 ( \37488 , \37467 , \37487 );
and \g446700/U$2 ( \37489 , \18711 , RIfc78650_6392);
and \g446700/U$3 ( \37490 , RIfcdbb60_7522, \18713 );
nor \g446700/U$1 ( \37491 , \37489 , \37490 );
and \g446701/U$2 ( \37492 , \18716 , RIe16beb8_2605);
and \g446701/U$3 ( \37493 , RIfc77b10_6384, \18718 );
nor \g446701/U$1 ( \37494 , \37492 , \37493 );
and \g446702/U$2 ( \37495 , \18533 , RIe168510_2564);
and \g446702/U$3 ( \37496 , RIe169e60_2582, \18535 );
nor \g446702/U$1 ( \37497 , \37495 , \37496 );
nand \g444580/U$1 ( \37498 , \37488 , \37491 , \37494 , \37497 );
and \g446690/U$2 ( \37499 , \16779 , RIdf1d920_1713);
and \g446690/U$3 ( \37500 , RIdf2d0a0_1889, \16781 );
nor \g446690/U$1 ( \37501 , \37499 , \37500 );
and \g445906/U$2 ( \37502 , RIdeb4e48_522, \16356 );
and \g445906/U$3 ( \37503 , RIde97cd0_330, \16485 );
and \g448756/U$2 ( \37504 , RIdece348_810, \16321 );
and \g448756/U$3 ( \37505 , \16326 , RIded1048_842);
and \g448756/U$4 ( \37506 , RIdf38a40_2021, \16427 );
nor \g448756/U$1 ( \37507 , \37504 , \37505 , \37506 );
and \g451470/U$2 ( \37508 , \16361 , RIde7dc18_203);
and \g451470/U$3 ( \37509 , RIdedc880_973, \16364 );
nor \g451470/U$1 ( \37510 , \37508 , \37509 );
and \g453733/U$2 ( \37511 , \16377 , RIdec8948_746);
and \g453733/U$3 ( \37512 , RIdecb648_778, \16313 );
nor \g453733/U$1 ( \37513 , \37511 , \37512 );
and \g455185/U$2 ( \37514 , \16317 , RIdee7b18_1100);
and \g455185/U$3 ( \37515 , RIdf01018_1388, \16325 );
nor \g455185/U$1 ( \37516 , \37514 , \37515 );
not \g455184/U$1 ( \37517 , \37516 );
and \g449784/U$2 ( \37518 , \37517 , \16336 );
and \g449784/U$3 ( \37519 , RIe144048_2151, \16448 );
nor \g449784/U$1 ( \37520 , \37518 , \37519 );
nand \g448040/U$1 ( \37521 , \37507 , \37510 , \37513 , \37520 );
nor \g445906/U$1 ( \37522 , \37502 , \37503 , \37521 );
not \g444926/U$3 ( \37523 , \37522 );
not \g444926/U$4 ( \37524 , \16586 );
and \g444926/U$2 ( \37525 , \37523 , \37524 );
and \g445908/U$2 ( \37526 , RIfcdc538_7529, \16313 );
and \g445908/U$3 ( \37527 , RIded5ad0_895, \16364 );
and \g448760/U$2 ( \37528 , RIfcd4978_7441, \16427 );
and \g448760/U$3 ( \37529 , \16448 , RIfcb0d20_7034);
and \g448760/U$4 ( \37530 , RIfca5218_6901, \16321 );
nor \g448760/U$1 ( \37531 , \37528 , \37529 , \37530 );
and \g451479/U$2 ( \37532 , \16368 , RIfca1708_6859);
and \g451479/U$3 ( \37533 , RIfca49a8_6895, \16371 );
nor \g451479/U$1 ( \37534 , \37532 , \37533 );
and \g454384/U$2 ( \37535 , \16317 , RIdee3360_1049);
and \g454384/U$3 ( \37536 , RIdee50e8_1070, \16325 );
nor \g454384/U$1 ( \37537 , \37535 , \37536 );
not \g449788/U$3 ( \37538 , \37537 );
not \g449788/U$4 ( \37539 , \16330 );
and \g449788/U$2 ( \37540 , \37538 , \37539 );
and \g449788/U$5 ( \37541 , \16326 , RIfcdf3a0_7562);
nor \g449788/U$1 ( \37542 , \37540 , \37541 );
and \g451478/U$2 ( \37543 , \16334 , RIdedefe0_1001);
and \g451478/U$3 ( \37544 , RIfea07a0_8170, \16380 );
nor \g451478/U$1 ( \37545 , \37543 , \37544 );
nand \g447601/U$1 ( \37546 , \37531 , \37534 , \37542 , \37545 );
nor \g445908/U$1 ( \37547 , \37526 , \37527 , \37546 );
and \g451473/U$2 ( \37548 , \16341 , RIded9fb8_944);
and \g451473/U$3 ( \37549 , RIfcdc6a0_7530, \16377 );
nor \g451473/U$1 ( \37550 , \37548 , \37549 );
and \g451475/U$2 ( \37551 , \16361 , RIfeab498_8265);
and \g451475/U$3 ( \37552 , RIded79c0_917, \16398 );
nor \g451475/U$1 ( \37553 , \37551 , \37552 );
and \g445080/U$2 ( \37554 , \37547 , \37550 , \37553 );
nor \g445080/U$1 ( \37555 , \37554 , \16909 );
nor \g444926/U$1 ( \37556 , \37525 , \37555 );
and \g446691/U$2 ( \37557 , \17032 , RIe15a848_2407);
and \g446691/U$3 ( \37558 , RIe16ea50_2636, \17029 );
nor \g446691/U$1 ( \37559 , \37557 , \37558 );
nand \g444423/U$1 ( \37560 , \37501 , \37556 , \37559 );
and \g445900/U$2 ( \37561 , RIfc7c160_6434, \16313 );
and \g445900/U$3 ( \37562 , RIde9e5d0_362, \16361 );
and \g448749/U$2 ( \37563 , RIdeb2148_490, \16427 );
and \g448749/U$3 ( \37564 , \16432 , RIfce7c08_7659);
and \g448749/U$4 ( \37565 , RIdec2f48_682, \16319 );
nor \g448749/U$1 ( \37566 , \37563 , \37564 , \37565 );
and \g451455/U$2 ( \37567 , \16368 , RIdeaf448_458);
and \g451455/U$3 ( \37568 , RIfce7aa0_7658, \16371 );
nor \g451455/U$1 ( \37569 , \37567 , \37568 );
and \g454648/U$2 ( \37570 , \16317 , RIdebd548_618);
and \g454648/U$3 ( \37571 , RIfcb38b8_7065, \16325 );
nor \g454648/U$1 ( \37572 , \37570 , \37571 );
not \g449779/U$3 ( \37573 , \37572 );
not \g449779/U$4 ( \37574 , \16330 );
and \g449779/U$2 ( \37575 , \37573 , \37574 );
and \g449779/U$5 ( \37576 , \16328 , RIdec5c48_714);
nor \g449779/U$1 ( \37577 , \37575 , \37576 );
and \g451453/U$2 ( \37578 , \16334 , RIdeb7b48_554);
and \g451453/U$3 ( \37579 , RIdeba848_586, \16380 );
nor \g451453/U$1 ( \37580 , \37578 , \37579 );
nand \g447594/U$1 ( \37581 , \37566 , \37569 , \37577 , \37580 );
nor \g445900/U$1 ( \37582 , \37561 , \37562 , \37581 );
and \g451450/U$2 ( \37583 , \16364 , RIdea4ed0_394);
and \g451450/U$3 ( \37584 , RIfca38c8_6883, \16339 );
nor \g451450/U$1 ( \37585 , \37583 , \37584 );
and \g451448/U$2 ( \37586 , \16398 , RIdeab7d0_426);
and \g451448/U$3 ( \37587 , RIdec0248_650, \16377 );
nor \g451448/U$1 ( \37588 , \37586 , \37587 );
and \g445075/U$2 ( \37589 , \37582 , \37585 , \37588 );
nor \g445075/U$1 ( \37590 , \37589 , \16618 );
and \g445902/U$2 ( \37591 , RIe141618_2121, \16356 );
and \g445902/U$3 ( \37592 , RIdf3ac00_2045, \16334 );
and \g448752/U$2 ( \37593 , RIfc9ecd8_6829, \16321 );
and \g448752/U$3 ( \37594 , \16326 , RIfc9eb70_6828);
and \g448752/U$4 ( \37595 , RIfcd3cd0_7432, \16427 );
nor \g448752/U$1 ( \37596 , \37593 , \37594 , \37595 );
and \g451461/U$2 ( \37597 , \16361 , RIdf2f968_1918);
and \g451461/U$3 ( \37598 , RIdf31858_1940, \16364 );
nor \g451461/U$1 ( \37599 , \37597 , \37598 );
and \g451460/U$2 ( \37600 , \16377 , RIfc83bb8_6521);
and \g451460/U$3 ( \37601 , RIfcc5630_7268, \16313 );
nor \g451460/U$1 ( \37602 , \37600 , \37601 );
and \g454995/U$2 ( \37603 , \16317 , RIdf33a18_1964);
and \g454995/U$3 ( \37604 , RIdf36010_1991, \16325 );
nor \g454995/U$1 ( \37605 , \37603 , \37604 );
not \g454994/U$1 ( \37606 , \37605 );
and \g449782/U$2 ( \37607 , \37606 , \16336 );
and \g449782/U$3 ( \37608 , RIee308e0_5011, \16448 );
nor \g449782/U$1 ( \37609 , \37607 , \37608 );
nand \g448039/U$1 ( \37610 , \37596 , \37599 , \37602 , \37609 );
nor \g445902/U$1 ( \37611 , \37591 , \37592 , \37610 );
and \g451456/U$2 ( \37612 , \16371 , RIfc84e00_6534);
and \g451456/U$3 ( \37613 , RIdf3d1f8_2072, \16380 );
nor \g451456/U$1 ( \37614 , \37612 , \37613 );
and \g451458/U$2 ( \37615 , \16368 , RIfc834b0_6516);
and \g451458/U$3 ( \37616 , RIfea0ea8_8175, \16485 );
nor \g451458/U$1 ( \37617 , \37615 , \37616 );
and \g445077/U$2 ( \37618 , \37611 , \37614 , \37617 );
nor \g445077/U$1 ( \37619 , \37618 , \16393 );
or \g444309/U$1 ( \37620 , \37498 , \37560 , \37590 , \37619 );
and \g445895/U$2 ( \37621 , RIdf0c418_1516, \16356 );
and \g445895/U$3 ( \37622 , RIdf03d18_1420, \16334 );
and \g448741/U$2 ( \37623 , RIdf14b18_1612, \16321 );
and \g448741/U$3 ( \37624 , \16328 , RIdf17818_1644);
and \g448741/U$4 ( \37625 , RIdefb618_1324, \16427 );
nor \g448741/U$1 ( \37626 , \37623 , \37624 , \37625 );
and \g451428/U$2 ( \37627 , \16361 , RIdeea818_1132);
and \g451428/U$3 ( \37628 , RIdeed518_1164, \16364 );
nor \g451428/U$1 ( \37629 , \37627 , \37628 );
and \g451426/U$2 ( \37630 , \16377 , RIdf0f118_1548);
and \g451426/U$3 ( \37631 , RIdf11e18_1580, \16313 );
nor \g451426/U$1 ( \37632 , \37630 , \37631 );
and \g454141/U$2 ( \37633 , \16317 , RIdef0218_1196);
and \g454141/U$3 ( \37634 , RIdef2f18_1228, \16325 );
nor \g454141/U$1 ( \37635 , \37633 , \37634 );
not \g454140/U$1 ( \37636 , \37635 );
and \g449771/U$2 ( \37637 , \37636 , \16336 );
and \g449771/U$3 ( \37638 , RIdefe318_1356, \16432 );
nor \g449771/U$1 ( \37639 , \37637 , \37638 );
nand \g448038/U$1 ( \37640 , \37626 , \37629 , \37632 , \37639 );
nor \g445895/U$1 ( \37641 , \37621 , \37622 , \37640 );
and \g451421/U$2 ( \37642 , \16371 , RIdef8918_1292);
and \g451421/U$3 ( \37643 , RIdf06a18_1452, \16380 );
nor \g451421/U$1 ( \37644 , \37642 , \37643 );
and \g451423/U$2 ( \37645 , \16368 , RIdef5c18_1260);
and \g451423/U$3 ( \37646 , RIdf09718_1484, \16485 );
nor \g451423/U$1 ( \37647 , \37645 , \37646 );
and \g445070/U$2 ( \37648 , \37641 , \37644 , \37647 );
nor \g445070/U$1 ( \37649 , \37648 , \16555 );
and \g445897/U$2 ( \37650 , RIdf21b38_1760, \16341 );
and \g445897/U$3 ( \37651 , RIee28078_4914, \16377 );
and \g448744/U$2 ( \37652 , RIfca0628_6847, \16427 );
and \g448744/U$3 ( \37653 , \16432 , RIfcd4f18_7445);
and \g448744/U$4 ( \37654 , RIee2a7d8_4942, \16319 );
nor \g448744/U$1 ( \37655 , \37652 , \37653 , \37654 );
and \g451442/U$2 ( \37656 , \16368 , RIfcd3190_7424);
and \g451442/U$3 ( \37657 , RIdf23050_1775, \16371 );
nor \g451442/U$1 ( \37658 , \37656 , \37657 );
and \g454627/U$2 ( \37659 , \16317 , RIdf28780_1837);
and \g454627/U$3 ( \37660 , RIdf2a940_1861, \16325 );
nor \g454627/U$1 ( \37661 , \37659 , \37660 );
not \g449774/U$3 ( \37662 , \37661 );
not \g449774/U$4 ( \37663 , \16330 );
and \g449774/U$2 ( \37664 , \37662 , \37663 );
and \g449774/U$5 ( \37665 , \16328 , RIee2c128_4960);
nor \g449774/U$1 ( \37666 , \37664 , \37665 );
and \g451440/U$2 ( \37667 , \16334 , RIfea0908_8171);
and \g451440/U$3 ( \37668 , RIfea0a70_8172, \16380 );
nor \g451440/U$1 ( \37669 , \37667 , \37668 );
nand \g447592/U$1 ( \37670 , \37655 , \37658 , \37666 , \37669 );
nor \g445897/U$1 ( \37671 , \37650 , \37651 , \37670 );
and \g451435/U$2 ( \37672 , \16361 , RIdf199d8_1668);
and \g451435/U$3 ( \37673 , RIee292c0_4927, \16313 );
nor \g451435/U$1 ( \37674 , \37672 , \37673 );
and \g451436/U$2 ( \37675 , \16364 , RIdf1b328_1686);
and \g451436/U$3 ( \37676 , RIdf20080_1741, \16398 );
nor \g451436/U$1 ( \37677 , \37675 , \37676 );
and \g445072/U$2 ( \37678 , \37671 , \37674 , \37677 );
nor \g445072/U$1 ( \37679 , \37678 , \16480 );
or \g444256/U$1 ( \37680 , \37620 , \37649 , \37679 );
_DC \g60cd/U$1 ( \37681 , \37680 , \16652 );
and \g448779/U$2 ( \37682 , RIfca9f70_6956, \8373 );
and \g448779/U$3 ( \37683 , \8330 , RIe224238_4701);
and \g448779/U$4 ( \37684 , RIe213438_4509, \8488 );
nor \g448779/U$1 ( \37685 , \37682 , \37683 , \37684 );
and \g454170/U$2 ( \37686 , \8313 , RIe218e38_4573);
and \g454170/U$3 ( \37687 , RIe21e838_4637, \8323 );
nor \g454170/U$1 ( \37688 , \37686 , \37687 );
not \g449807/U$3 ( \37689 , \37688 );
not \g449807/U$4 ( \37690 , \8376 );
and \g449807/U$2 ( \37691 , \37689 , \37690 );
and \g449807/U$5 ( \37692 , \8359 , RIfc3fda0_5752);
nor \g449807/U$1 ( \37693 , \37691 , \37692 );
and \g451557/U$2 ( \37694 , \8404 , RIe221538_4669);
and \g451557/U$3 ( \37695 , RIfc65528_6175, \8351 );
nor \g451557/U$1 ( \37696 , \37694 , \37695 );
and \g451559/U$2 ( \37697 , \8378 , RIe216138_4541);
and \g451559/U$3 ( \37698 , RIfc6b4c8_6243, \8417 );
nor \g451559/U$1 ( \37699 , \37697 , \37698 );
nand \g447614/U$1 ( \37700 , \37685 , \37693 , \37696 , \37699 );
and \g444766/U$2 ( \37701 , \37700 , \8369 );
and \g445926/U$2 ( \37702 , RIfcadbe8_6999, \8417 );
and \g445926/U$3 ( \37703 , RIe200fb8_4301, \8404 );
and \g448783/U$2 ( \37704 , RIe1fd070_4256, \8531 );
and \g448783/U$3 ( \37705 , \8488 , RIfc73358_6333);
and \g448783/U$4 ( \37706 , RIfccbcd8_7341, \8383 );
nor \g448783/U$1 ( \37707 , \37704 , \37705 , \37706 );
and \g451569/U$2 ( \37708 , \8335 , RIfca7270_6924);
and \g451569/U$3 ( \37709 , RIfcc2660_7234, \8340 );
nor \g451569/U$1 ( \37710 , \37708 , \37709 );
and \g455049/U$2 ( \37711 , \8313 , RIf15a940_5490);
and \g455049/U$3 ( \37712 , RIfc44468_5799, \8323 );
nor \g455049/U$1 ( \37713 , \37711 , \37712 );
not \g455048/U$1 ( \37714 , \37713 );
and \g449811/U$2 ( \37715 , \37714 , \8316 );
and \g449811/U$3 ( \37716 , RIfc66ba8_6191, \8351 );
nor \g449811/U$1 ( \37717 , \37715 , \37716 );
and \g451567/U$2 ( \37718 , \8356 , RIe1fbe28_4243);
and \g451567/U$3 ( \37719 , RIfca6898_6917, \8359 );
nor \g451567/U$1 ( \37720 , \37718 , \37719 );
nand \g448166/U$1 ( \37721 , \37707 , \37710 , \37717 , \37720 );
nor \g445926/U$1 ( \37722 , \37702 , \37703 , \37721 );
and \g451564/U$2 ( \37723 , \8378 , RIfc6a3e8_6231);
and \g451564/U$3 ( \37724 , RIe202bd8_4321, \8373 );
nor \g451564/U$1 ( \37725 , \37723 , \37724 );
and \g451562/U$2 ( \37726 , \8414 , RIfca7540_6926);
and \g451562/U$3 ( \37727 , RIfccbe40_7342, \8409 );
nor \g451562/U$1 ( \37728 , \37726 , \37727 );
and \g445095/U$2 ( \37729 , \37722 , \37725 , \37728 );
nor \g445095/U$1 ( \37730 , \37729 , \8422 );
nor \g444766/U$1 ( \37731 , \37701 , \37730 );
and \g446712/U$2 ( \37732 , \8707 , RIe208038_4381);
and \g446712/U$3 ( \37733 , RIe20ad38_4413, \8709 );
nor \g446712/U$1 ( \37734 , \37732 , \37733 );
and \g446714/U$2 ( \37735 , \8712 , RIe20da38_4445);
and \g446714/U$3 ( \37736 , RIfc60c08_6123, \8714 );
nor \g446714/U$1 ( \37737 , \37735 , \37736 );
and \g446713/U$2 ( \37738 , \8717 , RIe210738_4477);
and \g446713/U$3 ( \37739 , RIfc61310_6128, \8719 );
nor \g446713/U$1 ( \37740 , \37738 , \37739 );
nand \g444474/U$1 ( \37741 , \37731 , \37734 , \37737 , \37740 );
and \g451581/U$2 ( \37742 , \8319 , RIfc5a128_6047);
and \g451581/U$3 ( \37743 , RIfcbc3f0_7164, \8326 );
nor \g451581/U$1 ( \37744 , \37742 , \37743 );
and \g445929/U$2 ( \37745 , RIe1f39f8_4149, \8356 );
and \g445929/U$3 ( \37746 , RIfc99440_6766, \8340 );
and \g448789/U$2 ( \37747 , RIfc7e050_6456, \8373 );
and \g448789/U$3 ( \37748 , \8383 , RIfc5dda0_6090);
and \g448789/U$4 ( \37749 , RIfc8cdf8_6625, \8488 );
nor \g448789/U$1 ( \37750 , \37747 , \37748 , \37749 );
and \g454594/U$2 ( \37751 , \8313 , RIfc8d668_6631);
and \g454594/U$3 ( \37752 , RIfcd9568_7495, \8323 );
nor \g454594/U$1 ( \37753 , \37751 , \37752 );
not \g449818/U$3 ( \37754 , \37753 );
not \g449818/U$4 ( \37755 , \8376 );
and \g449818/U$2 ( \37756 , \37754 , \37755 );
and \g449818/U$5 ( \37757 , \8359 , RIfca4138_6889);
nor \g449818/U$1 ( \37758 , \37756 , \37757 );
and \g451584/U$2 ( \37759 , \8404 , RIe1fa7a8_4227);
and \g451584/U$3 ( \37760 , RIfc5e070_6092, \8351 );
nor \g451584/U$1 ( \37761 , \37759 , \37760 );
and \g451586/U$2 ( \37762 , \8378 , RIe1f5d20_4174);
and \g451586/U$3 ( \37763 , RIfc5d968_6087, \8417 );
nor \g451586/U$1 ( \37764 , \37762 , \37763 );
nand \g447619/U$1 ( \37765 , \37750 , \37758 , \37761 , \37764 );
nor \g445929/U$1 ( \37766 , \37745 , \37746 , \37765 );
and \g451582/U$2 ( \37767 , \8335 , RIe1ee700_4090);
and \g451582/U$3 ( \37768 , RIfcc7c28_7295, \8531 );
nor \g451582/U$1 ( \37769 , \37767 , \37768 );
nand \g445559/U$1 ( \37770 , \37744 , \37766 , \37769 );
and \g444723/U$2 ( \37771 , \37770 , \8752 );
and \g448785/U$2 ( \37772 , RIe1c1ca0_3582, \8317 );
and \g448785/U$3 ( \37773 , \8326 , RIe1c49a0_3614);
and \g448785/U$4 ( \37774 , RIe1e92a0_4030, \8330 );
nor \g448785/U$1 ( \37775 , \37772 , \37773 , \37774 );
and \g451578/U$2 ( \37776 , \8335 , RIe1befa0_3550);
and \g451578/U$3 ( \37777 , RIe1c76a0_3646, \8340 );
nor \g451578/U$1 ( \37778 , \37776 , \37777 );
and \g454735/U$2 ( \37779 , \8313 , RIe1cd0a0_3710);
and \g454735/U$3 ( \37780 , RIe1cfda0_3742, \8323 );
nor \g454735/U$1 ( \37781 , \37779 , \37780 );
not \g449815/U$3 ( \37782 , \37781 );
not \g449815/U$4 ( \37783 , \8347 );
and \g449815/U$2 ( \37784 , \37782 , \37783 );
and \g449815/U$5 ( \37785 , \8351 , RIe1ebfa0_4062);
nor \g449815/U$1 ( \37786 , \37784 , \37785 );
and \g451577/U$2 ( \37787 , \8356 , RIe1ca3a0_3678);
and \g451577/U$3 ( \37788 , RIe1d2aa0_3774, \8359 );
nor \g451577/U$1 ( \37789 , \37787 , \37788 );
nand \g447617/U$1 ( \37790 , \37775 , \37778 , \37786 , \37789 );
and \g444723/U$3 ( \37791 , \8478 , \37790 );
nor \g444723/U$1 ( \37792 , \37771 , \37791 );
and \g446716/U$2 ( \37793 , \9480 , RIe1e38a0_3966);
and \g446716/U$3 ( \37794 , RIe1e65a0_3998, \9482 );
nor \g446716/U$1 ( \37795 , \37793 , \37794 );
and \g446717/U$2 ( \37796 , \10539 , RIe1d84a0_3838);
and \g446717/U$3 ( \37797 , RIe1db1a0_3870, \10541 );
nor \g446717/U$1 ( \37798 , \37796 , \37797 );
and \g446715/U$2 ( \37799 , \10534 , RIe1ddea0_3902);
and \g446715/U$3 ( \37800 , RIe1e0ba0_3934, \10536 );
nor \g446715/U$1 ( \37801 , \37799 , \37800 );
nand \g444584/U$1 ( \37802 , \37792 , \37795 , \37798 , \37801 );
and \g445919/U$2 ( \37803 , RIfc4c460_5890, \8417 );
and \g445919/U$3 ( \37804 , RIe1b7980_3466, \8404 );
and \g448773/U$2 ( \37805 , RIe1b2ac0_3410, \8531 );
and \g448773/U$3 ( \37806 , \8488 , RIf147f20_5278);
and \g448773/U$4 ( \37807 , RIf14bb98_5321, \8330 );
nor \g448773/U$1 ( \37808 , \37805 , \37806 , \37807 );
and \g451535/U$2 ( \37809 , \8335 , RIe1ab338_3325);
and \g451535/U$3 ( \37810 , RIf1473e0_5270, \8340 );
nor \g451535/U$1 ( \37811 , \37809 , \37810 );
and \g454725/U$2 ( \37812 , \8313 , RIe1acb20_3342);
and \g454725/U$3 ( \37813 , RIf1468a0_5262, \8323 );
nor \g454725/U$1 ( \37814 , \37812 , \37813 );
not \g454724/U$1 ( \37815 , \37814 );
and \g449803/U$2 ( \37816 , \37815 , \8316 );
and \g449803/U$3 ( \37817 , RIf14cde0_5334, \8351 );
nor \g449803/U$1 ( \37818 , \37816 , \37817 );
and \g451531/U$2 ( \37819 , \8356 , RIe1b1170_3392);
and \g451531/U$3 ( \37820 , RIf149168_5291, \8359 );
nor \g451531/U$1 ( \37821 , \37819 , \37820 );
nand \g448164/U$1 ( \37822 , \37808 , \37811 , \37818 , \37821 );
nor \g445919/U$1 ( \37823 , \37803 , \37804 , \37822 );
and \g451529/U$2 ( \37824 , \8378 , RIfec54d8_8365);
and \g451529/U$3 ( \37825 , RIe1b99d8_3489, \8373 );
nor \g451529/U$1 ( \37826 , \37824 , \37825 );
and \g451528/U$2 ( \37827 , \8412 , RIe1b5658_3441);
and \g451528/U$3 ( \37828 , RIfc9e738_6825, \8409 );
nor \g451528/U$1 ( \37829 , \37827 , \37828 );
and \g445090/U$2 ( \37830 , \37823 , \37826 , \37829 );
nor \g445090/U$1 ( \37831 , \37830 , \8481 );
and \g445921/U$2 ( \37832 , RIe18d0e0_2982, \8417 );
and \g445921/U$3 ( \37833 , RIe1a0be0_3206, \8404 );
and \g448777/U$2 ( \37834 , RIe1af118_3369, \8319 );
and \g448777/U$3 ( \37835 , \8326 , RIe1bc2a0_3518);
and \g448777/U$4 ( \37836 , RIe1a65e0_3270, \8383 );
nor \g448777/U$1 ( \37837 , \37834 , \37835 , \37836 );
and \g451545/U$2 ( \37838 , \8335 , RIe171750_2668);
and \g451545/U$3 ( \37839 , RIe1d57a0_3806, \8340 );
nor \g451545/U$1 ( \37840 , \37838 , \37839 );
and \g454337/U$2 ( \37841 , \8313 , RIe1f8750_4204);
and \g454337/U$3 ( \37842 , RIe1ff398_4281, \8323 );
nor \g454337/U$1 ( \37843 , \37841 , \37842 );
not \g449805/U$3 ( \37844 , \37843 );
not \g449805/U$4 ( \37845 , \8347 );
and \g449805/U$2 ( \37846 , \37844 , \37845 );
and \g449805/U$5 ( \37847 , \8351 , RIe1a92e0_3302);
nor \g449805/U$1 ( \37848 , \37846 , \37847 );
and \g451544/U$2 ( \37849 , \8356 , RIe1f1298_4121);
and \g451544/U$3 ( \37850 , RIe205338_4349, \8359 );
nor \g451544/U$1 ( \37851 , \37849 , \37850 );
nand \g447610/U$1 ( \37852 , \37837 , \37840 , \37848 , \37851 );
nor \g445921/U$1 ( \37853 , \37832 , \37833 , \37852 );
and \g451541/U$2 ( \37854 , \8378 , RIe21bb38_4605);
and \g451541/U$3 ( \37855 , RIe1a38e0_3238, \8373 );
nor \g451541/U$1 ( \37856 , \37854 , \37855 );
and \g451539/U$2 ( \37857 , \8414 , RIe226f38_4733);
and \g451539/U$3 ( \37858 , RIe1795e0_2758, \8409 );
nor \g451539/U$1 ( \37859 , \37857 , \37858 );
and \g445091/U$2 ( \37860 , \37853 , \37856 , \37859 );
nor \g445091/U$1 ( \37861 , \37860 , \8651 );
or \g444323/U$1 ( \37862 , \37741 , \37802 , \37831 , \37861 );
and \g445915/U$2 ( \37863 , RIfcca928_7327, \8417 );
and \g445915/U$3 ( \37864 , RIfea0638_8169, \8404 );
and \g448767/U$2 ( \37865 , RIf16e5a8_5715, \8317 );
and \g448767/U$3 ( \37866 , \8326 , RIfc650f0_6172);
and \g448767/U$4 ( \37867 , RIfc65690_6176, \8330 );
nor \g448767/U$1 ( \37868 , \37865 , \37866 , \37867 );
and \g451513/U$2 ( \37869 , \8335 , RIfc43a90_5792);
and \g451513/U$3 ( \37870 , RIfcecf00_7718, \8340 );
nor \g451513/U$1 ( \37871 , \37869 , \37870 );
and \g454560/U$2 ( \37872 , \8313 , RIee39f58_5118);
and \g454560/U$3 ( \37873 , RIfca9430_6948, \8323 );
nor \g454560/U$1 ( \37874 , \37872 , \37873 );
not \g449796/U$3 ( \37875 , \37874 );
not \g449796/U$4 ( \37876 , \8347 );
and \g449796/U$2 ( \37877 , \37875 , \37876 );
and \g449796/U$5 ( \37878 , \8351 , RIfc65d98_6181);
nor \g449796/U$1 ( \37879 , \37877 , \37878 );
and \g451511/U$2 ( \37880 , \8356 , RIe174018_2697);
and \g451511/U$3 ( \37881 , RIee3c3e8_5144, \8359 );
nor \g451511/U$1 ( \37882 , \37880 , \37881 );
nand \g447606/U$1 ( \37883 , \37868 , \37871 , \37879 , \37882 );
nor \g445915/U$1 ( \37884 , \37863 , \37864 , \37883 );
and \g451507/U$2 ( \37885 , \8378 , RIee3d798_5158);
and \g451507/U$3 ( \37886 , RIe1772b8_2733, \8373 );
nor \g451507/U$1 ( \37887 , \37885 , \37886 );
and \g451506/U$2 ( \37888 , \8414 , RIfc65258_6173);
and \g451506/U$3 ( \37889 , RIfc607d0_6120, \8409 );
nor \g451506/U$1 ( \37890 , \37888 , \37889 );
and \g445086/U$2 ( \37891 , \37884 , \37887 , \37890 );
nor \g445086/U$1 ( \37892 , \37891 , \8558 );
and \g445917/U$2 ( \37893 , RIe1849e0_2886, \8356 );
and \g445917/U$3 ( \37894 , RIfcaa7e0_6962, \8340 );
and \g448771/U$2 ( \37895 , RIe192ae0_3046, \8414 );
and \g448771/U$3 ( \37896 , \8409 , RIe1957e0_3078);
and \g448771/U$4 ( \37897 , RIe1876e0_2918, \8488 );
nor \g448771/U$1 ( \37898 , \37895 , \37896 , \37897 );
and \g454656/U$2 ( \37899 , \8313 , RIfc67580_6198);
and \g454656/U$3 ( \37900 , RIe19b1e0_3142, \8323 );
nor \g454656/U$1 ( \37901 , \37899 , \37900 );
not \g449799/U$3 ( \37902 , \37901 );
not \g449799/U$4 ( \37903 , \8328 );
and \g449799/U$2 ( \37904 , \37902 , \37903 );
and \g449799/U$5 ( \37905 , \8359 , RIe18a3e0_2950);
nor \g449799/U$1 ( \37906 , \37904 , \37905 );
and \g451519/U$2 ( \37907 , \8404 , RIe1984e0_3110);
and \g451519/U$3 ( \37908 , RIe19dee0_3174, \8351 );
nor \g451519/U$1 ( \37909 , \37907 , \37908 );
and \g451522/U$2 ( \37910 , \8378 , RIe18fde0_3014);
and \g451522/U$3 ( \37911 , RIfccb030_7332, \8417 );
nor \g451522/U$1 ( \37912 , \37910 , \37911 );
nand \g447607/U$1 ( \37913 , \37898 , \37906 , \37909 , \37912 );
nor \g445917/U$1 ( \37914 , \37893 , \37894 , \37913 );
and \g451517/U$2 ( \37915 , \8335 , RIe17c2e0_2790);
and \g451517/U$3 ( \37916 , RIfc6a550_6232, \8531 );
nor \g451517/U$1 ( \37917 , \37915 , \37916 );
and \g451516/U$2 ( \37918 , \8319 , RIe17efe0_2822);
and \g451516/U$3 ( \37919 , RIe181ce0_2854, \8324 );
nor \g451516/U$1 ( \37920 , \37918 , \37919 );
and \g445088/U$2 ( \37921 , \37914 , \37917 , \37920 );
nor \g445088/U$1 ( \37922 , \37921 , \8589 );
or \g444273/U$1 ( \37923 , \37862 , \37892 , \37922 );
_DC \g6151/U$1 ( \37924 , \37923 , \8654 );
and \g452204/U$2 ( \37925 , \16371 , RIfc750e0_6354);
and \g452204/U$3 ( \37926 , RIfea1448_8179, \16427 );
nor \g452204/U$1 ( \37927 , \37925 , \37926 );
and \g446089/U$2 ( \37928 , RIde82448_225, \16432 );
and \g446089/U$3 ( \37929 , RIe168678_2565, \16361 );
and \g448991/U$2 ( \37930 , RIfcedd10_7728, \16321 );
and \g448991/U$3 ( \37931 , \16328 , RIee1d218_4790);
and \g448991/U$4 ( \37932 , RIfec5eb0_8372, \16398 );
nor \g448991/U$1 ( \37933 , \37930 , \37931 , \37932 );
and \g454400/U$2 ( \37934 , \16317 , RIde8e928_285);
and \g454400/U$3 ( \37935 , RIde91da8_301, \16325 );
nor \g454400/U$1 ( \37936 , \37934 , \37935 );
not \g450004/U$3 ( \37937 , \37936 );
not \g450004/U$4 ( \37938 , \16330 );
and \g450004/U$2 ( \37939 , \37937 , \37938 );
and \g450004/U$5 ( \37940 , \16341 , RIfced8d8_7725);
nor \g450004/U$1 ( \37941 , \37939 , \37940 );
and \g452209/U$2 ( \37942 , \16377 , RIfcc92a8_7311);
and \g452209/U$3 ( \37943 , RIfce62b8_7641, \16313 );
nor \g452209/U$1 ( \37944 , \37942 , \37943 );
and \g452210/U$2 ( \37945 , \16334 , RIde865e8_245);
and \g452210/U$3 ( \37946 , RIde8a788_265, \16380 );
nor \g452210/U$1 ( \37947 , \37945 , \37946 );
nand \g447341/U$1 ( \37948 , \37933 , \37941 , \37944 , \37947 );
nor \g446089/U$1 ( \37949 , \37928 , \37929 , \37948 );
and \g452205/U$2 ( \37950 , \16364 , RIe169fc8_2583);
and \g452205/U$3 ( \37951 , RIfcc19b8_7225, \16368 );
nor \g452205/U$1 ( \37952 , \37950 , \37951 );
nand \g445596/U$1 ( \37953 , \37927 , \37949 , \37952 );
and \g444707/U$2 ( \37954 , \37953 , \17998 );
and \g448989/U$2 ( \37955 , RIdebd6b0_619, \16485 );
and \g448989/U$3 ( \37956 , \16356 , RIfcaf538_7017);
and \g448989/U$4 ( \37957 , RIdeabb18_427, \16337 );
nor \g448989/U$1 ( \37958 , \37955 , \37956 , \37957 );
and \g454751/U$2 ( \37959 , \16317 , RIdec30b0_683);
and \g454751/U$3 ( \37960 , RIdec5db0_715, \16325 );
nor \g454751/U$1 ( \37961 , \37959 , \37960 );
not \g450003/U$3 ( \37962 , \37961 );
not \g450003/U$4 ( \37963 , \16311 );
and \g450003/U$2 ( \37964 , \37962 , \37963 );
and \g450003/U$5 ( \37965 , \16341 , RIee1dd58_4798);
nor \g450003/U$1 ( \37966 , \37964 , \37965 );
and \g452201/U$2 ( \37967 , \16377 , RIdec03b0_651);
and \g452201/U$3 ( \37968 , RIee201e8_4824, \16313 );
nor \g452201/U$1 ( \37969 , \37967 , \37968 );
and \g452202/U$2 ( \37970 , \16334 , RIdeb7cb0_555);
and \g452202/U$3 ( \37971 , RIdeba9b0_587, \16380 );
nor \g452202/U$1 ( \37972 , \37970 , \37971 );
nand \g447340/U$1 ( \37973 , \37958 , \37966 , \37969 , \37972 );
and \g444707/U$3 ( \37974 , \17938 , \37973 );
nor \g444707/U$1 ( \37975 , \37954 , \37974 );
and \g446860/U$2 ( \37976 , \18457 , RIdeb22b0_491);
and \g446860/U$3 ( \37977 , RIfc40fe8_5765, \18459 );
nor \g446860/U$1 ( \37978 , \37976 , \37977 );
and \g446861/U$2 ( \37979 , \18462 , RIdeaf5b0_459);
and \g446861/U$3 ( \37980 , RIfcd08c8_7395, \18464 );
nor \g446861/U$1 ( \37981 , \37979 , \37980 );
and \g446862/U$2 ( \37982 , \18467 , RIde9e918_363);
and \g446862/U$3 ( \37983 , RIdea5218_395, \18469 );
nor \g446862/U$1 ( \37984 , \37982 , \37983 );
nand \g444495/U$1 ( \37985 , \37975 , \37978 , \37981 , \37984 );
and \g452217/U$2 ( \37986 , \16380 , RIe157cb0_2376);
and \g452217/U$3 ( \37987 , RIe1630b0_2504, \16321 );
nor \g452217/U$1 ( \37988 , \37986 , \37987 );
and \g446091/U$2 ( \37989 , RIe165db0_2536, \16328 );
and \g446091/U$3 ( \37990 , RIe1603b0_2472, \16377 );
and \g448994/U$2 ( \37991 , RIe1522b0_2312, \16427 );
and \g448994/U$3 ( \37992 , \16448 , RIfea1718_8181);
and \g448994/U$4 ( \37993 , RIe15d6b0_2440, \16485 );
nor \g448994/U$1 ( \37994 , \37991 , \37992 , \37993 );
and \g454759/U$2 ( \37995 , \16317 , RIe14c8b0_2248);
and \g454759/U$3 ( \37996 , RIfcb0348_7027, \16325 );
nor \g454759/U$1 ( \37997 , \37995 , \37996 );
not \g454758/U$1 ( \37998 , \37997 );
and \g450007/U$2 ( \37999 , \37998 , \16336 );
and \g450007/U$3 ( \38000 , RIee365b0_5077, \16356 );
nor \g450007/U$1 ( \38001 , \37999 , \38000 );
and \g452220/U$2 ( \38002 , \16361 , RIe146eb0_2184);
and \g452220/U$3 ( \38003 , RIe149bb0_2216, \16364 );
nor \g452220/U$1 ( \38004 , \38002 , \38003 );
and \g452219/U$2 ( \38005 , \16368 , RIe14f5b0_2280);
and \g452219/U$3 ( \38006 , RIee35200_5063, \16371 );
nor \g452219/U$1 ( \38007 , \38005 , \38006 );
nand \g448066/U$1 ( \38008 , \37994 , \38001 , \38004 , \38007 );
nor \g446091/U$1 ( \38009 , \37989 , \37990 , \38008 );
and \g452216/U$2 ( \38010 , \16334 , RIe154fb0_2344);
and \g452216/U$3 ( \38011 , RIfccfc20_7386, \16313 );
nor \g452216/U$1 ( \38012 , \38010 , \38011 );
nand \g445597/U$1 ( \38013 , \37988 , \38009 , \38012 );
and \g444858/U$2 ( \38014 , \38013 , \16390 );
and \g448992/U$2 ( \38015 , RIdf33b80_1965, \16398 );
and \g448992/U$3 ( \38016 , \16341 , RIdf36178_1992);
and \g448992/U$4 ( \38017 , RIe13f2f0_2096, \16344 );
nor \g448992/U$1 ( \38018 , \38015 , \38016 , \38017 );
and \g454755/U$2 ( \38019 , \16317 , RIfc5fb28_6111);
and \g454755/U$3 ( \38020 , RIfea15b0_8180, \16325 );
nor \g454755/U$1 ( \38021 , \38019 , \38020 );
not \g450005/U$3 ( \38022 , \38021 );
not \g450005/U$4 ( \38023 , \16351 );
and \g450005/U$2 ( \38024 , \38022 , \38023 );
and \g450005/U$5 ( \38025 , \16356 , RIe141780_2122);
nor \g450005/U$1 ( \38026 , \38024 , \38025 );
and \g452215/U$2 ( \38027 , \16361 , RIdf2fad0_1919);
and \g452215/U$3 ( \38028 , RIdf319c0_1941, \16364 );
nor \g452215/U$1 ( \38029 , \38027 , \38028 );
and \g452212/U$2 ( \38030 , \16368 , RIfc74438_6345);
and \g452212/U$3 ( \38031 , RIfcae728_7007, \16371 );
nor \g452212/U$1 ( \38032 , \38030 , \38031 );
nand \g447723/U$1 ( \38033 , \38018 , \38026 , \38029 , \38032 );
and \g444858/U$3 ( \38034 , \16394 , \38033 );
nor \g444858/U$1 ( \38035 , \38014 , \38034 );
and \g446867/U$2 ( \38036 , \16705 , RIdf3ad68_2046);
and \g446867/U$3 ( \38037 , RIfec5be0_8370, \16707 );
nor \g446867/U$1 ( \38038 , \38036 , \38037 );
and \g446866/U$2 ( \38039 , \16710 , RIfcdf238_7561);
and \g446866/U$3 ( \38040 , RIfc73790_6336, \16712 );
nor \g446866/U$1 ( \38041 , \38039 , \38040 );
and \g446868/U$2 ( \38042 , \16715 , RIfc94f58_6717);
and \g446868/U$3 ( \38043 , RIee32500_5031, \16717 );
nor \g446868/U$1 ( \38044 , \38042 , \38043 );
nand \g444610/U$1 ( \38045 , \38035 , \38038 , \38041 , \38044 );
and \g446086/U$2 ( \38046 , RIfccaa90_7328, \16427 );
and \g446086/U$3 ( \38047 , RIfcad4e0_6994, \16368 );
and \g448986/U$2 ( \38048 , RIee2a940_4943, \16321 );
and \g448986/U$3 ( \38049 , \16326 , RIee2c290_4961);
and \g448986/U$4 ( \38050 , RIfeaad90_8260, \16337 );
nor \g448986/U$1 ( \38051 , \38048 , \38049 , \38050 );
and \g454343/U$2 ( \38052 , \16317 , RIdf288e8_1838);
and \g454343/U$3 ( \38053 , RIdf2aaa8_1862, \16325 );
nor \g454343/U$1 ( \38054 , \38052 , \38053 );
not \g449999/U$3 ( \38055 , \38054 );
not \g449999/U$4 ( \38056 , \16330 );
and \g449999/U$2 ( \38057 , \38055 , \38056 );
and \g449999/U$5 ( \38058 , \16341 , RIdf21ca0_1761);
nor \g449999/U$1 ( \38059 , \38057 , \38058 );
and \g452190/U$2 ( \38060 , \16377 , RIfc704f0_6300);
and \g452190/U$3 ( \38061 , RIfc70658_6301, \16313 );
nor \g452190/U$1 ( \38062 , \38060 , \38061 );
and \g452191/U$2 ( \38063 , \16334 , RIdf24f40_1797);
and \g452191/U$3 ( \38064 , RIdf269f8_1816, \16380 );
nor \g452191/U$1 ( \38065 , \38063 , \38064 );
nand \g447337/U$1 ( \38066 , \38051 , \38059 , \38062 , \38065 );
nor \g446086/U$1 ( \38067 , \38046 , \38047 , \38066 );
and \g452188/U$2 ( \38068 , \16361 , RIdf19b40_1669);
and \g452188/U$3 ( \38069 , RIfc64b50_6168, \16448 );
nor \g452188/U$1 ( \38070 , \38068 , \38069 );
and \g452187/U$2 ( \38071 , \16364 , RIdf1b490_1687);
and \g452187/U$3 ( \38072 , RIdf231b8_1776, \16371 );
nor \g452187/U$1 ( \38073 , \38071 , \38072 );
and \g445214/U$2 ( \38074 , \38067 , \38070 , \38073 );
nor \g445214/U$1 ( \38075 , \38074 , \16480 );
and \g446088/U$2 ( \38076 , RIee22510_4849, \16427 );
and \g446088/U$3 ( \38077 , RIfc6cb48_6259, \16368 );
and \g448987/U$2 ( \38078 , RIfea7f28_8227, \16485 );
and \g448987/U$3 ( \38079 , \16356 , RIdee5250_1071);
and \g448987/U$4 ( \38080 , RIded7b28_918, \16398 );
nor \g448987/U$1 ( \38081 , \38078 , \38079 , \38080 );
and \g454410/U$2 ( \38082 , \16317 , RIfcac568_6983);
and \g454410/U$3 ( \38083 , RIfc595e8_6039, \16325 );
nor \g454410/U$1 ( \38084 , \38082 , \38083 );
not \g450001/U$3 ( \38085 , \38084 );
not \g450001/U$4 ( \38086 , \16311 );
and \g450001/U$2 ( \38087 , \38085 , \38086 );
and \g450001/U$5 ( \38088 , \16341 , RIdeda120_945);
nor \g450001/U$1 ( \38089 , \38087 , \38088 );
and \g452198/U$2 ( \38090 , \16377 , RIfccd358_7357);
and \g452198/U$3 ( \38091 , RIfcccf20_7354, \16313 );
nor \g452198/U$1 ( \38092 , \38090 , \38091 );
and \g452199/U$2 ( \38093 , \16334 , RIfea12e0_8178);
and \g452199/U$3 ( \38094 , RIdee11a0_1025, \16380 );
nor \g452199/U$1 ( \38095 , \38093 , \38094 );
nand \g447339/U$1 ( \38096 , \38081 , \38089 , \38092 , \38095 );
nor \g446088/U$1 ( \38097 , \38076 , \38077 , \38096 );
and \g452195/U$2 ( \38098 , \16361 , RIfec5d48_8371);
and \g452195/U$3 ( \38099 , RIfc679b8_6201, \16448 );
nor \g452195/U$1 ( \38100 , \38098 , \38099 );
and \g452194/U$2 ( \38101 , \16364 , RIded5c38_896);
and \g452194/U$3 ( \38102 , RIfc6dd90_6272, \16371 );
nor \g452194/U$1 ( \38103 , \38101 , \38102 );
and \g445215/U$2 ( \38104 , \38097 , \38100 , \38103 );
nor \g445215/U$1 ( \38105 , \38104 , \16909 );
or \g444330/U$1 ( \38106 , \37985 , \38045 , \38075 , \38105 );
and \g446082/U$2 ( \38107 , RIdf38ba8_2022, \16427 );
and \g446082/U$3 ( \38108 , RIdf1da88_1714, \16368 );
and \g448982/U$2 ( \38109 , RIdece4b0_811, \16321 );
and \g448982/U$3 ( \38110 , \16328 , RIded11b0_843);
and \g448982/U$4 ( \38111 , RIdee7c80_1101, \16398 );
nor \g448982/U$1 ( \38112 , \38109 , \38110 , \38111 );
and \g454423/U$2 ( \38113 , \16317 , RIde98018_331);
and \g454423/U$3 ( \38114 , RIdeb4fb0_523, \16325 );
nor \g454423/U$1 ( \38115 , \38113 , \38114 );
not \g449994/U$3 ( \38116 , \38115 );
not \g449994/U$4 ( \38117 , \16330 );
and \g449994/U$2 ( \38118 , \38116 , \38117 );
and \g449994/U$5 ( \38119 , \16341 , RIdf01180_1389);
nor \g449994/U$1 ( \38120 , \38118 , \38119 );
and \g452177/U$2 ( \38121 , \16377 , RIdec8ab0_747);
and \g452177/U$3 ( \38122 , RIdecb7b0_779, \16313 );
nor \g452177/U$1 ( \38123 , \38121 , \38122 );
and \g452176/U$2 ( \38124 , \16334 , RIe15a9b0_2408);
and \g452176/U$3 ( \38125 , RIe16ebb8_2637, \16380 );
nor \g452176/U$1 ( \38126 , \38124 , \38125 );
nand \g447335/U$1 ( \38127 , \38112 , \38120 , \38123 , \38126 );
nor \g446082/U$1 ( \38128 , \38107 , \38108 , \38127 );
and \g452174/U$2 ( \38129 , \16361 , RIde7df60_204);
and \g452174/U$3 ( \38130 , RIe1441b0_2152, \16448 );
nor \g452174/U$1 ( \38131 , \38129 , \38130 );
and \g452172/U$2 ( \38132 , \16364 , RIdedc9e8_974);
and \g452172/U$3 ( \38133 , RIdf2d208_1890, \16371 );
nor \g452172/U$1 ( \38134 , \38132 , \38133 );
and \g445212/U$2 ( \38135 , \38128 , \38131 , \38134 );
nor \g445212/U$1 ( \38136 , \38135 , \16586 );
and \g446083/U$2 ( \38137 , RIdefb780_1325, \16427 );
and \g446083/U$3 ( \38138 , RIdef5d80_1261, \16368 );
and \g448984/U$2 ( \38139 , RIdf09880_1485, \16485 );
and \g448984/U$3 ( \38140 , \16354 , RIdf0c580_1517);
and \g448984/U$4 ( \38141 , RIdef0380_1197, \16337 );
nor \g448984/U$1 ( \38142 , \38139 , \38140 , \38141 );
and \g454747/U$2 ( \38143 , \16317 , RIdf14c80_1613);
and \g454747/U$3 ( \38144 , RIdf17980_1645, \16325 );
nor \g454747/U$1 ( \38145 , \38143 , \38144 );
not \g449997/U$3 ( \38146 , \38145 );
not \g449997/U$4 ( \38147 , \16311 );
and \g449997/U$2 ( \38148 , \38146 , \38147 );
and \g449997/U$5 ( \38149 , \16341 , RIdef3080_1229);
nor \g449997/U$1 ( \38150 , \38148 , \38149 );
and \g452182/U$2 ( \38151 , \16377 , RIdf0f280_1549);
and \g452182/U$3 ( \38152 , RIdf11f80_1581, \16313 );
nor \g452182/U$1 ( \38153 , \38151 , \38152 );
and \g452184/U$2 ( \38154 , \16334 , RIdf03e80_1421);
and \g452184/U$3 ( \38155 , RIdf06b80_1453, \16380 );
nor \g452184/U$1 ( \38156 , \38154 , \38155 );
nand \g447336/U$1 ( \38157 , \38142 , \38150 , \38153 , \38156 );
nor \g446083/U$1 ( \38158 , \38137 , \38138 , \38157 );
and \g452181/U$2 ( \38159 , \16361 , RIdeea980_1133);
and \g452181/U$3 ( \38160 , RIdefe480_1357, \16448 );
nor \g452181/U$1 ( \38161 , \38159 , \38160 );
and \g452180/U$2 ( \38162 , \16364 , RIdeed680_1165);
and \g452180/U$3 ( \38163 , RIdef8a80_1293, \16371 );
nor \g452180/U$1 ( \38164 , \38162 , \38163 );
and \g445213/U$2 ( \38165 , \38158 , \38161 , \38164 );
nor \g445213/U$1 ( \38166 , \38165 , \16555 );
or \g444226/U$1 ( \38167 , \38106 , \38136 , \38166 );
_DC \g61d6/U$1 ( \38168 , \38167 , \16652 );
and \g452266/U$2 ( \38169 , \8317 , RIfec57a8_8367);
and \g452266/U$3 ( \38170 , RIfec5910_8368, \8404 );
nor \g452266/U$1 ( \38171 , \38169 , \38170 );
and \g446103/U$2 ( \38172 , RIe1b9b40_3490, \8373 );
and \g446103/U$3 ( \38173 , RIfc78d58_6397, \8383 );
and \g449007/U$2 ( \38174 , RIf146a08_5263, \8326 );
and \g449007/U$3 ( \38175 , \8531 , RIe1b2c28_3411);
and \g449007/U$4 ( \38176 , RIfec5a78_8369, \8488 );
nor \g449007/U$1 ( \38177 , \38174 , \38175 , \38176 );
and \g452270/U$2 ( \38178 , \8356 , RIe1b12d8_3393);
and \g452270/U$3 ( \38179 , RIf1492d0_5292, \8359 );
nor \g452270/U$1 ( \38180 , \38178 , \38179 );
and \g454776/U$2 ( \38181 , \8313 , RIe1b57c0_3442);
and \g454776/U$3 ( \38182 , RIfcd51e8_7447, \8323 );
nor \g454776/U$1 ( \38183 , \38181 , \38182 );
not \g450021/U$3 ( \38184 , \38183 );
not \g450021/U$4 ( \38185 , \8376 );
and \g450021/U$2 ( \38186 , \38184 , \38185 );
and \g450021/U$5 ( \38187 , \8340 , RIfec5640_8366);
nor \g450021/U$1 ( \38188 , \38186 , \38187 );
and \g452269/U$2 ( \38189 , \8378 , RIfea1010_8176);
and \g452269/U$3 ( \38190 , RIfc78a88_6395, \8417 );
nor \g452269/U$1 ( \38191 , \38189 , \38190 );
nand \g447735/U$1 ( \38192 , \38177 , \38180 , \38188 , \38191 );
nor \g446103/U$1 ( \38193 , \38172 , \38173 , \38192 );
and \g452265/U$2 ( \38194 , \8335 , RIfea1178_8177);
and \g452265/U$3 ( \38195 , RIf14cf48_5335, \8351 );
nor \g452265/U$1 ( \38196 , \38194 , \38195 );
nand \g445599/U$1 ( \38197 , \38171 , \38193 , \38196 );
and \g444916/U$2 ( \38198 , \38197 , \8482 );
and \g449005/U$2 ( \38199 , RIe2270a0_4734, \8414 );
and \g449005/U$3 ( \38200 , \8409 , RIe179748_2759);
and \g449005/U$4 ( \38201 , RIe1bc408_3519, \8326 );
nor \g449005/U$1 ( \38202 , \38199 , \38200 , \38201 );
and \g452262/U$2 ( \38203 , \8356 , RIe1f1400_4122);
and \g452262/U$3 ( \38204 , RIe2054a0_4350, \8359 );
nor \g452262/U$1 ( \38205 , \38203 , \38204 );
and \g454775/U$2 ( \38206 , \8313 , RIe1f88b8_4205);
and \g454775/U$3 ( \38207 , RIe1ff500_4282, \8323 );
nor \g454775/U$1 ( \38208 , \38206 , \38207 );
not \g450019/U$3 ( \38209 , \38208 );
not \g450019/U$4 ( \38210 , \8347 );
and \g450019/U$2 ( \38211 , \38209 , \38210 );
and \g450019/U$5 ( \38212 , \8340 , RIe1d5908_3807);
nor \g450019/U$1 ( \38213 , \38211 , \38212 );
and \g452261/U$2 ( \38214 , \8378 , RIe21bca0_4606);
and \g452261/U$3 ( \38215 , RIe18d248_2983, \8417 );
nor \g452261/U$1 ( \38216 , \38214 , \38215 );
nand \g447733/U$1 ( \38217 , \38202 , \38205 , \38213 , \38216 );
and \g444916/U$3 ( \38218 , \9010 , \38217 );
nor \g444916/U$1 ( \38219 , \38198 , \38218 );
and \g446875/U$2 ( \38220 , \9041 , RIe1a0d48_3207);
and \g446875/U$3 ( \38221 , RIe1a3a48_3239, \9043 );
nor \g446875/U$1 ( \38222 , \38220 , \38221 );
and \g446874/U$2 ( \38223 , \14956 , RIe1a6748_3271);
and \g446874/U$3 ( \38224 , RIe1a9448_3303, \14958 );
nor \g446874/U$1 ( \38225 , \38223 , \38224 );
and \g446876/U$2 ( \38226 , \13244 , RIe1718b8_2669);
and \g446876/U$3 ( \38227 , RIe1af280_3370, \13246 );
nor \g446876/U$1 ( \38228 , \38226 , \38227 );
nand \g444611/U$1 ( \38229 , \38219 , \38222 , \38225 , \38228 );
and \g446869/U$2 ( \38230 , \10230 , RIe1fbf90_4244);
and \g446869/U$3 ( \38231 , RIe1fd1d8_4257, \10232 );
nor \g446869/U$1 ( \38232 , \38230 , \38231 );
and \g446099/U$2 ( \38233 , RIfc44a08_5803, \8488 );
and \g446099/U$3 ( \38234 , RIfca2680_6870, \8359 );
and \g449001/U$2 ( \38235 , RIfc487e8_5847, \8409 );
and \g449001/U$3 ( \38236 , \8371 , RIe202d40_4322);
and \g449001/U$4 ( \38237 , RIfc7f568_6471, \8383 );
nor \g449001/U$1 ( \38238 , \38235 , \38236 , \38237 );
and \g452252/U$2 ( \38239 , \8335 , RIfce01b0_7572);
and \g452252/U$3 ( \38240 , RIfc580d0_6024, \8340 );
nor \g452252/U$1 ( \38241 , \38239 , \38240 );
and \g452251/U$2 ( \38242 , \8404 , RIe201120_4302);
and \g452251/U$3 ( \38243 , RIfc8c9c0_6622, \8351 );
nor \g452251/U$1 ( \38244 , \38242 , \38243 );
and \g454769/U$2 ( \38245 , \8313 , RIfc8dd70_6636);
and \g454769/U$3 ( \38246 , RIfcbdbd8_7181, \8323 );
nor \g454769/U$1 ( \38247 , \38245 , \38246 );
not \g454768/U$1 ( \38248 , \38247 );
and \g450016/U$2 ( \38249 , \38248 , \8316 );
and \g450016/U$3 ( \38250 , RIfce2910_7600, \8417 );
nor \g450016/U$1 ( \38251 , \38249 , \38250 );
nand \g448188/U$1 ( \38252 , \38238 , \38241 , \38244 , \38251 );
nor \g446099/U$1 ( \38253 , \38233 , \38234 , \38252 );
not \g444868/U$3 ( \38254 , \38253 );
not \g444868/U$4 ( \38255 , \8422 );
and \g444868/U$2 ( \38256 , \38254 , \38255 );
and \g446100/U$2 ( \38257 , RIe218fa0_4574, \8414 );
and \g446100/U$3 ( \38258 , RIf169418_5657, \8523 );
and \g449004/U$2 ( \38259 , RIe20aea0_4414, \8319 );
and \g449004/U$3 ( \38260 , \8324 , RIe20dba0_4446);
and \g449004/U$4 ( \38261 , RIe21e9a0_4638, \8407 );
nor \g449004/U$1 ( \38262 , \38259 , \38260 , \38261 );
and \g452257/U$2 ( \38263 , \8335 , RIe2081a0_4382);
and \g452257/U$3 ( \38264 , RIfc8bfe8_6615, \8340 );
nor \g452257/U$1 ( \38265 , \38263 , \38264 );
and \g452256/U$2 ( \38266 , \8404 , RIe2216a0_4670);
and \g452256/U$3 ( \38267 , RIfc48c20_5850, \8351 );
nor \g452256/U$1 ( \38268 , \38266 , \38267 );
and \g454773/U$2 ( \38269 , \8313 , RIfca0358_6845);
and \g454773/U$3 ( \38270 , RIe2243a0_4702, \8323 );
nor \g454773/U$1 ( \38271 , \38269 , \38270 );
not \g450018/U$3 ( \38272 , \38271 );
not \g450018/U$4 ( \38273 , \8328 );
and \g450018/U$2 ( \38274 , \38272 , \38273 );
and \g450018/U$5 ( \38275 , \8417 , RIfc9a688_6779);
nor \g450018/U$1 ( \38276 , \38274 , \38275 );
nand \g447732/U$1 ( \38277 , \38262 , \38265 , \38268 , \38276 );
nor \g446100/U$1 ( \38278 , \38257 , \38258 , \38277 );
and \g452254/U$2 ( \38279 , \8356 , RIe2108a0_4478);
and \g452254/U$3 ( \38280 , RIfc456b0_5812, \8359 );
nor \g452254/U$1 ( \38281 , \38279 , \38280 );
and \g452255/U$2 ( \38282 , \8378 , RIe2162a0_4542);
and \g452255/U$3 ( \38283 , RIe2135a0_4510, \8488 );
nor \g452255/U$1 ( \38284 , \38282 , \38283 );
and \g445222/U$2 ( \38285 , \38278 , \38281 , \38284 );
nor \g445222/U$1 ( \38286 , \38285 , \8368 );
nor \g444868/U$1 ( \38287 , \38256 , \38286 );
and \g446870/U$2 ( \38288 , \14165 , RIfc992d8_6765);
and \g446870/U$3 ( \38289 , RIfc46d30_5828, \14167 );
nor \g446870/U$1 ( \38290 , \38288 , \38289 );
nand \g444427/U$1 ( \38291 , \38232 , \38287 , \38290 );
and \g446096/U$2 ( \38292 , RIe19e048_3175, \8351 );
and \g446096/U$3 ( \38293 , RIe198648_3111, \8404 );
and \g448998/U$2 ( \38294 , RIe181e48_2855, \8326 );
and \g448998/U$3 ( \38295 , \8531 , RIfc46790_5824);
and \g448998/U$4 ( \38296 , RIe187848_2919, \8488 );
nor \g448998/U$1 ( \38297 , \38294 , \38295 , \38296 );
and \g452242/U$2 ( \38298 , \8356 , RIe184b48_2887);
and \g452242/U$3 ( \38299 , RIe18a548_2951, \8359 );
nor \g452242/U$1 ( \38300 , \38298 , \38299 );
and \g454763/U$2 ( \38301 , \8313 , RIe192c48_3047);
and \g454763/U$3 ( \38302 , RIe195948_3079, \8323 );
nor \g454763/U$1 ( \38303 , \38301 , \38302 );
not \g450012/U$3 ( \38304 , \38303 );
not \g450012/U$4 ( \38305 , \8376 );
and \g450012/U$2 ( \38306 , \38304 , \38305 );
and \g450012/U$5 ( \38307 , \8340 , RIfc98d38_6761);
nor \g450012/U$1 ( \38308 , \38306 , \38307 );
and \g452241/U$2 ( \38309 , \8378 , RIe18ff48_3015);
and \g452241/U$3 ( \38310 , RIfc7efc8_6467, \8417 );
nor \g452241/U$1 ( \38311 , \38309 , \38310 );
nand \g447730/U$1 ( \38312 , \38297 , \38300 , \38308 , \38311 );
nor \g446096/U$1 ( \38313 , \38292 , \38293 , \38312 );
and \g452239/U$2 ( \38314 , \8335 , RIe17c448_2791);
and \g452239/U$3 ( \38315 , RIe19b348_3143, \8383 );
nor \g452239/U$1 ( \38316 , \38314 , \38315 );
and \g452238/U$2 ( \38317 , \8319 , RIe17f148_2823);
and \g452238/U$3 ( \38318 , RIfcc3ce0_7250, \8373 );
nor \g452238/U$1 ( \38319 , \38317 , \38318 );
and \g445218/U$2 ( \38320 , \38313 , \38316 , \38319 );
nor \g445218/U$1 ( \38321 , \38320 , \8589 );
and \g446097/U$2 ( \38322 , RIfc8b778_6609, \8414 );
and \g446097/U$3 ( \38323 , RIee3a0c0_5119, \8531 );
and \g448999/U$2 ( \38324 , RIf16e710_5716, \8319 );
and \g448999/U$3 ( \38325 , \8324 , RIfcbc288_7163);
and \g448999/U$4 ( \38326 , RIfcd2bf0_7420, \8409 );
nor \g448999/U$1 ( \38327 , \38324 , \38325 , \38326 );
and \g452248/U$2 ( \38328 , \8335 , RIfc8fdc8_6659);
and \g452248/U$3 ( \38329 , RIfc46628_5823, \8340 );
nor \g452248/U$1 ( \38330 , \38328 , \38329 );
and \g452247/U$2 ( \38331 , \8404 , RIe1761d8_2721);
and \g452247/U$3 ( \38332 , RIfcb5d48_7091, \8351 );
nor \g452247/U$1 ( \38333 , \38331 , \38332 );
and \g454766/U$2 ( \38334 , \8313 , RIfc9a3b8_6777);
and \g454766/U$3 ( \38335 , RIfc995a8_6767, \8323 );
nor \g454766/U$1 ( \38336 , \38334 , \38335 );
not \g450015/U$3 ( \38337 , \38336 );
not \g450015/U$4 ( \38338 , \8328 );
and \g450015/U$2 ( \38339 , \38337 , \38338 );
and \g450015/U$5 ( \38340 , \8417 , RIfc54188_5979);
nor \g450015/U$1 ( \38341 , \38339 , \38340 );
nand \g447731/U$1 ( \38342 , \38327 , \38330 , \38333 , \38341 );
nor \g446097/U$1 ( \38343 , \38322 , \38323 , \38342 );
and \g452245/U$2 ( \38344 , \8356 , RIfeaba38_8269);
and \g452245/U$3 ( \38345 , RIee3c550_5145, \8359 );
nor \g452245/U$1 ( \38346 , \38344 , \38345 );
and \g452244/U$2 ( \38347 , \8378 , RIfc7dee8_6455);
and \g452244/U$3 ( \38348 , RIfc8c420_6618, \8488 );
nor \g452244/U$1 ( \38349 , \38347 , \38348 );
and \g445220/U$2 ( \38350 , \38343 , \38346 , \38349 );
nor \g445220/U$1 ( \38351 , \38350 , \8558 );
or \g444310/U$1 ( \38352 , \38229 , \38291 , \38321 , \38351 );
and \g446094/U$2 ( \38353 , RIfc7b8f0_6428, \8373 );
and \g446094/U$3 ( \38354 , RIfc90368_6663, \8330 );
and \g448995/U$2 ( \38355 , RIfc7b788_6427, \8414 );
and \g448995/U$3 ( \38356 , \8409 , RIfc43ec8_5795);
and \g448995/U$4 ( \38357 , RIfcdb728_7519, \8326 );
nor \g448995/U$1 ( \38358 , \38355 , \38356 , \38357 );
and \g452228/U$2 ( \38359 , \8356 , RIe1f3b60_4150);
and \g452228/U$3 ( \38360 , RIfc7b350_6424, \8359 );
nor \g452228/U$1 ( \38361 , \38359 , \38360 );
and \g454760/U$2 ( \38362 , \8313 , RIfca3490_6880);
and \g454760/U$3 ( \38363 , RIfc90d40_6670, \8323 );
nor \g454760/U$1 ( \38364 , \38362 , \38363 );
not \g450008/U$3 ( \38365 , \38364 );
not \g450008/U$4 ( \38366 , \8347 );
and \g450008/U$2 ( \38367 , \38365 , \38366 );
and \g450008/U$5 ( \38368 , \8340 , RIfc91010_6672);
nor \g450008/U$1 ( \38369 , \38367 , \38368 );
and \g452227/U$2 ( \38370 , \8378 , RIe1f5e88_4175);
and \g452227/U$3 ( \38371 , RIfcd8b90_7488, \8417 );
nor \g452227/U$1 ( \38372 , \38370 , \38371 );
nand \g447727/U$1 ( \38373 , \38358 , \38361 , \38369 , \38372 );
nor \g446094/U$1 ( \38374 , \38353 , \38354 , \38373 );
and \g452223/U$2 ( \38375 , \8335 , RIe1ee868_4091);
and \g452223/U$3 ( \38376 , RIfc7bbc0_6430, \8351 );
nor \g452223/U$1 ( \38377 , \38375 , \38376 );
and \g452224/U$2 ( \38378 , \8319 , RIfcd8758_7485);
and \g452224/U$3 ( \38379 , RIe1fa910_4228, \8404 );
nor \g452224/U$1 ( \38380 , \38378 , \38379 );
and \g445216/U$2 ( \38381 , \38374 , \38377 , \38380 );
nor \g445216/U$1 ( \38382 , \38381 , \8621 );
and \g446095/U$2 ( \38383 , RIe1db308_3871, \8412 );
and \g446095/U$3 ( \38384 , RIe1ca508_3679, \8356 );
and \g448996/U$2 ( \38385 , RIe1c1e08_3583, \8319 );
and \g448996/U$3 ( \38386 , \8326 , RIe1c4b08_3615);
and \g448996/U$4 ( \38387 , RIe1de008_3903, \8409 );
nor \g448996/U$1 ( \38388 , \38385 , \38386 , \38387 );
and \g452235/U$2 ( \38389 , \8335 , RIe1bf108_3551);
and \g452235/U$3 ( \38390 , RIe1c7808_3647, \8340 );
nor \g452235/U$1 ( \38391 , \38389 , \38390 );
and \g452236/U$2 ( \38392 , \8404 , RIe1e3a08_3967);
and \g452236/U$3 ( \38393 , RIe1ec108_4063, \8351 );
nor \g452236/U$1 ( \38394 , \38392 , \38393 );
and \g454387/U$2 ( \38395 , \8313 , RIe1e6708_3999);
and \g454387/U$3 ( \38396 , RIe1e9408_4031, \8323 );
nor \g454387/U$1 ( \38397 , \38395 , \38396 );
not \g450009/U$3 ( \38398 , \38397 );
not \g450009/U$4 ( \38399 , \8328 );
and \g450009/U$2 ( \38400 , \38398 , \38399 );
and \g450009/U$5 ( \38401 , \8417 , RIe1e0d08_3935);
nor \g450009/U$1 ( \38402 , \38400 , \38401 );
nand \g447728/U$1 ( \38403 , \38388 , \38391 , \38394 , \38402 );
nor \g446095/U$1 ( \38404 , \38383 , \38384 , \38403 );
and \g452233/U$2 ( \38405 , \8378 , RIe1d8608_3839);
and \g452233/U$3 ( \38406 , RIe1d2c08_3775, \8359 );
nor \g452233/U$1 ( \38407 , \38405 , \38406 );
and \g452232/U$2 ( \38408 , \8531 , RIe1cd208_3711);
and \g452232/U$3 ( \38409 , RIe1cff08_3743, \8488 );
nor \g452232/U$1 ( \38410 , \38408 , \38409 );
and \g445217/U$2 ( \38411 , \38404 , \38407 , \38410 );
nor \g445217/U$1 ( \38412 , \38411 , \8477 );
or \g444252/U$1 ( \38413 , \38352 , \38382 , \38412 );
_DC \g625a/U$1 ( \38414 , \38413 , \8654 );
and \g452306/U$2 ( \38415 , \16361 , RIdeeaae8_1134);
and \g452306/U$3 ( \38416 , RIdefb8e8_1326, \16427 );
nor \g452306/U$1 ( \38417 , \38415 , \38416 );
and \g446111/U$2 ( \38418 , RIdefe5e8_1358, \16448 );
and \g446111/U$3 ( \38419 , RIdef8be8_1294, \16371 );
and \g449018/U$2 ( \38420 , RIdf099e8_1486, \16485 );
and \g449018/U$3 ( \38421 , \16356 , RIdf0c6e8_1518);
and \g449018/U$4 ( \38422 , RIdef04e8_1198, \16398 );
nor \g449018/U$1 ( \38423 , \38420 , \38421 , \38422 );
and \g454789/U$2 ( \38424 , \16317 , RIdf14de8_1614);
and \g454789/U$3 ( \38425 , RIdf17ae8_1646, \16325 );
nor \g454789/U$1 ( \38426 , \38424 , \38425 );
not \g450033/U$3 ( \38427 , \38426 );
not \g450033/U$4 ( \38428 , \16311 );
and \g450033/U$2 ( \38429 , \38427 , \38428 );
and \g450033/U$5 ( \38430 , \16341 , RIdef31e8_1230);
nor \g450033/U$1 ( \38431 , \38429 , \38430 );
and \g452307/U$2 ( \38432 , \16377 , RIdf0f3e8_1550);
and \g452307/U$3 ( \38433 , RIdf120e8_1582, \16313 );
nor \g452307/U$1 ( \38434 , \38432 , \38433 );
and \g452308/U$2 ( \38435 , \16334 , RIdf03fe8_1422);
and \g452308/U$3 ( \38436 , RIdf06ce8_1454, \16380 );
nor \g452308/U$1 ( \38437 , \38435 , \38436 );
nand \g447346/U$1 ( \38438 , \38423 , \38431 , \38434 , \38437 );
nor \g446111/U$1 ( \38439 , \38418 , \38419 , \38438 );
and \g452304/U$2 ( \38440 , \16364 , RIdeed7e8_1166);
and \g452304/U$3 ( \38441 , RIdef5ee8_1262, \16368 );
nor \g452304/U$1 ( \38442 , \38440 , \38441 );
nand \g445601/U$1 ( \38443 , \38417 , \38439 , \38442 );
and \g444775/U$2 ( \38444 , \38443 , \16750 );
and \g449017/U$2 ( \38445 , RIdf201e8_1742, \16398 );
and \g449017/U$3 ( \38446 , \16341 , RIfeabfd8_8273);
and \g449017/U$4 ( \38447 , RIdf28a50_1839, \16344 );
nor \g449017/U$1 ( \38448 , \38445 , \38446 , \38447 );
and \g454787/U$2 ( \38449 , \16317 , RIfcb9df8_7137);
and \g454787/U$3 ( \38450 , RIfc9b600_6790, \16325 );
nor \g454787/U$1 ( \38451 , \38449 , \38450 );
not \g450031/U$3 ( \38452 , \38451 );
not \g450031/U$4 ( \38453 , \16351 );
and \g450031/U$2 ( \38454 , \38452 , \38453 );
and \g450031/U$5 ( \38455 , \16356 , RIfea3e78_8209);
nor \g450031/U$1 ( \38456 , \38454 , \38455 );
and \g452299/U$2 ( \38457 , \16361 , RIdf19ca8_1670);
and \g452299/U$3 ( \38458 , RIdf1b5f8_1688, \16364 );
nor \g452299/U$1 ( \38459 , \38457 , \38458 );
and \g452298/U$2 ( \38460 , \16368 , RIfc86318_6549);
and \g452298/U$3 ( \38461 , RIdf23320_1777, \16371 );
nor \g452298/U$1 ( \38462 , \38460 , \38461 );
nand \g447737/U$1 ( \38463 , \38448 , \38456 , \38459 , \38462 );
and \g444775/U$3 ( \38464 , \16481 , \38463 );
nor \g444775/U$1 ( \38465 , \38444 , \38464 );
and \g446881/U$2 ( \38466 , \16505 , RIfc4cfa0_5898);
and \g446881/U$3 ( \38467 , RIee2c3f8_4962, \16507 );
nor \g446881/U$1 ( \38468 , \38466 , \38467 );
and \g446882/U$2 ( \38469 , \16511 , RIdf250a8_1798);
and \g446882/U$3 ( \38470 , RIdf26b60_1817, \16514 );
nor \g446882/U$1 ( \38471 , \38469 , \38470 );
and \g446880/U$2 ( \38472 , \16518 , RIfc4f430_5924);
and \g446880/U$3 ( \38473 , RIfc572c0_6014, \16521 );
nor \g446880/U$1 ( \38474 , \38472 , \38473 );
nand \g444498/U$1 ( \38475 , \38465 , \38468 , \38471 , \38474 );
and \g452315/U$2 ( \38476 , \16377 , RIdec8c18_748);
and \g452315/U$3 ( \38477 , RIe16ed20_2638, \16380 );
nor \g452315/U$1 ( \38478 , \38476 , \38477 );
and \g446113/U$2 ( \38479 , RIdece618_812, \16321 );
and \g446113/U$3 ( \38480 , RIdecb918_780, \16313 );
and \g449021/U$2 ( \38481 , RIdf38d10_2023, \16427 );
and \g449021/U$3 ( \38482 , \16448 , RIe144318_2153);
and \g449021/U$4 ( \38483 , RIde98360_332, \16344 );
nor \g449021/U$1 ( \38484 , \38481 , \38482 , \38483 );
and \g454794/U$2 ( \38485 , \16317 , RIdee7de8_1102);
and \g454794/U$3 ( \38486 , RIdf012e8_1390, \16325 );
nor \g454794/U$1 ( \38487 , \38485 , \38486 );
not \g454793/U$1 ( \38488 , \38487 );
and \g450036/U$2 ( \38489 , \38488 , \16336 );
and \g450036/U$3 ( \38490 , RIdeb5118_524, \16356 );
nor \g450036/U$1 ( \38491 , \38489 , \38490 );
and \g452317/U$2 ( \38492 , \16361 , RIde7e2a8_205);
and \g452317/U$3 ( \38493 , RIdedcb50_975, \16364 );
nor \g452317/U$1 ( \38494 , \38492 , \38493 );
and \g452316/U$2 ( \38495 , \16368 , RIdf1dbf0_1715);
and \g452316/U$3 ( \38496 , RIdf2d370_1891, \16371 );
nor \g452316/U$1 ( \38497 , \38495 , \38496 );
nand \g448071/U$1 ( \38498 , \38484 , \38491 , \38494 , \38497 );
nor \g446113/U$1 ( \38499 , \38479 , \38480 , \38498 );
and \g452314/U$2 ( \38500 , \16334 , RIe15ab18_2409);
and \g452314/U$3 ( \38501 , RIded1318_844, \16326 );
nor \g452314/U$1 ( \38502 , \38500 , \38501 );
nand \g445602/U$1 ( \38503 , \38478 , \38499 , \38502 );
and \g444892/U$2 ( \38504 , \38503 , \16752 );
and \g449020/U$2 ( \38505 , RIded7c90_919, \16398 );
and \g449020/U$3 ( \38506 , \16341 , RIdeda288_946);
and \g449020/U$4 ( \38507 , RIdee34c8_1050, \16485 );
nor \g449020/U$1 ( \38508 , \38505 , \38506 , \38507 );
and \g454792/U$2 ( \38509 , \16317 , RIfc4b0b0_5876);
and \g454792/U$3 ( \38510 , RIfcae188_7003, \16325 );
nor \g454792/U$1 ( \38511 , \38509 , \38510 );
not \g450035/U$3 ( \38512 , \38511 );
not \g450035/U$4 ( \38513 , \16351 );
and \g450035/U$2 ( \38514 , \38512 , \38513 );
and \g450035/U$5 ( \38515 , \16356 , RIdee53b8_1072);
nor \g450035/U$1 ( \38516 , \38514 , \38515 );
and \g452312/U$2 ( \38517 , \16361 , RIded3640_869);
and \g452312/U$3 ( \38518 , RIded5da0_897, \16364 );
nor \g452312/U$1 ( \38519 , \38517 , \38518 );
and \g452311/U$2 ( \38520 , \16368 , RIfce4968_7623);
and \g452311/U$3 ( \38521 , RIfc74870_6348, \16371 );
nor \g452311/U$1 ( \38522 , \38520 , \38521 );
nand \g447738/U$1 ( \38523 , \38508 , \38516 , \38519 , \38522 );
and \g444892/U$3 ( \38524 , \16477 , \38523 );
nor \g444892/U$1 ( \38525 , \38504 , \38524 );
and \g446883/U$2 ( \38526 , \18268 , RIfcc54c8_7267);
and \g446883/U$3 ( \38527 , RIfc89018_6581, \18270 );
nor \g446883/U$1 ( \38528 , \38526 , \38527 );
and \g446884/U$2 ( \38529 , \18273 , RIfc4b380_5878);
and \g446884/U$3 ( \38530 , RIfc89180_6582, \18275 );
nor \g446884/U$1 ( \38531 , \38529 , \38530 );
and \g446885/U$2 ( \38532 , \18278 , RIdedf148_1002);
and \g446885/U$3 ( \38533 , RIfea3d10_8208, \18280 );
nor \g446885/U$1 ( \38534 , \38532 , \38533 );
nand \g444612/U$1 ( \38535 , \38525 , \38528 , \38531 , \38534 );
and \g446107/U$2 ( \38536 , RIfce4da0_7626, \16448 );
and \g446107/U$3 ( \38537 , RIfcea908_7691, \16371 );
and \g449012/U$2 ( \38538 , RIdec3218_684, \16321 );
and \g449012/U$3 ( \38539 , \16328 , RIdec5f18_716);
and \g449012/U$4 ( \38540 , RIdeabe60_428, \16398 );
nor \g449012/U$1 ( \38541 , \38538 , \38539 , \38540 );
and \g454783/U$2 ( \38542 , \16317 , RIdebd818_620);
and \g454783/U$3 ( \38543 , RIee1f6a8_4816, \16325 );
nor \g454783/U$1 ( \38544 , \38542 , \38543 );
not \g450028/U$3 ( \38545 , \38544 );
not \g450028/U$4 ( \38546 , \16330 );
and \g450028/U$2 ( \38547 , \38545 , \38546 );
and \g450028/U$5 ( \38548 , \16341 , RIfce20a0_7594);
nor \g450028/U$1 ( \38549 , \38547 , \38548 );
and \g452288/U$2 ( \38550 , \16377 , RIdec0518_652);
and \g452288/U$3 ( \38551 , RIee20350_4825, \16313 );
nor \g452288/U$1 ( \38552 , \38550 , \38551 );
and \g452289/U$2 ( \38553 , \16334 , RIdeb7e18_556);
and \g452289/U$3 ( \38554 , RIdebab18_588, \16380 );
nor \g452289/U$1 ( \38555 , \38553 , \38554 );
nand \g447343/U$1 ( \38556 , \38541 , \38549 , \38552 , \38555 );
nor \g446107/U$1 ( \38557 , \38536 , \38537 , \38556 );
and \g452283/U$2 ( \38558 , \16364 , RIdea5560_396);
and \g452283/U$3 ( \38559 , RIdeaf718_460, \16368 );
nor \g452283/U$1 ( \38560 , \38558 , \38559 );
and \g452284/U$2 ( \38561 , \16361 , RIde9ec60_364);
and \g452284/U$3 ( \38562 , RIdeb2418_492, \16427 );
nor \g452284/U$1 ( \38563 , \38561 , \38562 );
and \g445228/U$2 ( \38564 , \38557 , \38560 , \38563 );
nor \g445228/U$1 ( \38565 , \38564 , \16618 );
and \g446108/U$2 ( \38566 , RIee33748_5044, \16321 );
and \g446108/U$3 ( \38567 , RIee32668_5032, \16313 );
and \g449016/U$2 ( \38568 , RIfc42848_5779, \16427 );
and \g449016/U$3 ( \38569 , \16432 , RIfc526d0_5960);
and \g449016/U$4 ( \38570 , RIe13f458_2097, \16344 );
nor \g449016/U$1 ( \38571 , \38568 , \38569 , \38570 );
and \g454351/U$2 ( \38572 , \16317 , RIdf33ce8_1966);
and \g454351/U$3 ( \38573 , RIfea42b0_8212, \16325 );
nor \g454351/U$1 ( \38574 , \38572 , \38573 );
not \g454350/U$1 ( \38575 , \38574 );
and \g450029/U$2 ( \38576 , \38575 , \16336 );
and \g450029/U$3 ( \38577 , RIe1418e8_2123, \16356 );
nor \g450029/U$1 ( \38578 , \38576 , \38577 );
and \g452294/U$2 ( \38579 , \16361 , RIdf2fc38_1920);
and \g452294/U$3 ( \38580 , RIdf31b28_1942, \16364 );
nor \g452294/U$1 ( \38581 , \38579 , \38580 );
and \g452293/U$2 ( \38582 , \16368 , RIfcb7260_7106);
and \g452293/U$3 ( \38583 , RIfcae9f8_7009, \16371 );
nor \g452293/U$1 ( \38584 , \38582 , \38583 );
nand \g448070/U$1 ( \38585 , \38571 , \38578 , \38581 , \38584 );
nor \g446108/U$1 ( \38586 , \38566 , \38567 , \38585 );
and \g452292/U$2 ( \38587 , \16377 , RIee31588_5020);
and \g452292/U$3 ( \38588 , RIdf3d360_2073, \16380 );
nor \g452292/U$1 ( \38589 , \38587 , \38588 );
and \g452291/U$2 ( \38590 , \16334 , RIdf3aed0_2047);
and \g452291/U$3 ( \38591 , RIee34828_5056, \16326 );
nor \g452291/U$1 ( \38592 , \38590 , \38591 );
and \g445229/U$2 ( \38593 , \38586 , \38589 , \38592 );
nor \g445229/U$1 ( \38594 , \38593 , \16393 );
or \g444396/U$1 ( \38595 , \38475 , \38535 , \38565 , \38594 );
and \g446104/U$2 ( \38596 , RIe165f18_2537, \16328 );
and \g446104/U$3 ( \38597 , RIe160518_2473, \16377 );
and \g449009/U$2 ( \38598 , RIe152418_2313, \16427 );
and \g449009/U$3 ( \38599 , \16448 , RIfc45548_5811);
and \g449009/U$4 ( \38600 , RIe15d818_2441, \16344 );
nor \g449009/U$1 ( \38601 , \38598 , \38599 , \38600 );
and \g454780/U$2 ( \38602 , \16317 , RIe14ca18_2249);
and \g454780/U$3 ( \38603 , RIfcbda70_7180, \16325 );
nor \g454780/U$1 ( \38604 , \38602 , \38603 );
not \g454779/U$1 ( \38605 , \38604 );
and \g450023/U$2 ( \38606 , \38605 , \16336 );
and \g450023/U$3 ( \38607 , RIfc55268_5991, \16356 );
nor \g450023/U$1 ( \38608 , \38606 , \38607 );
and \g452274/U$2 ( \38609 , \16361 , RIe147018_2185);
and \g452274/U$3 ( \38610 , RIe149d18_2217, \16364 );
nor \g452274/U$1 ( \38611 , \38609 , \38610 );
and \g452273/U$2 ( \38612 , \16368 , RIe14f718_2281);
and \g452273/U$3 ( \38613 , RIfc498c8_5859, \16371 );
nor \g452273/U$1 ( \38614 , \38612 , \38613 );
nand \g448068/U$1 ( \38615 , \38601 , \38608 , \38611 , \38614 );
nor \g446104/U$1 ( \38616 , \38596 , \38597 , \38615 );
and \g452272/U$2 ( \38617 , \16334 , RIe155118_2345);
and \g452272/U$3 ( \38618 , RIfcadd50_7000, \16313 );
nor \g452272/U$1 ( \38619 , \38617 , \38618 );
and \g452271/U$2 ( \38620 , \16380 , RIe157e18_2377);
and \g452271/U$3 ( \38621 , RIe163218_2505, \16321 );
nor \g452271/U$1 ( \38622 , \38620 , \38621 );
and \g445224/U$2 ( \38623 , \38616 , \38619 , \38622 );
nor \g445224/U$1 ( \38624 , \38623 , \16389 );
and \g446105/U$2 ( \38625 , RIfc6f848_6291, \16427 );
and \g446105/U$3 ( \38626 , RIfc76b98_6373, \16368 );
and \g449011/U$2 ( \38627 , RIee1c2a0_4779, \16321 );
and \g449011/U$3 ( \38628 , \16328 , RIfce6420_7642);
and \g449011/U$4 ( \38629 , RIe16c020_2606, \16337 );
nor \g449011/U$1 ( \38630 , \38627 , \38628 , \38629 );
and \g454781/U$2 ( \38631 , \16317 , RIfea4148_8211);
and \g454781/U$3 ( \38632 , RIde920f0_302, \16325 );
nor \g454781/U$1 ( \38633 , \38631 , \38632 );
not \g450025/U$3 ( \38634 , \38633 );
not \g450025/U$4 ( \38635 , \16330 );
and \g450025/U$2 ( \38636 , \38634 , \38635 );
and \g450025/U$5 ( \38637 , \16339 , RIfcae2f0_7004);
nor \g450025/U$1 ( \38638 , \38636 , \38637 );
and \g452280/U$2 ( \38639 , \16377 , RIee1ad88_4764);
and \g452280/U$3 ( \38640 , RIfc75950_6360, \16313 );
nor \g452280/U$1 ( \38641 , \38639 , \38640 );
and \g452281/U$2 ( \38642 , \16334 , RIfea3fe0_8210);
and \g452281/U$3 ( \38643 , RIfeaa688_8255, \16380 );
nor \g452281/U$1 ( \38644 , \38642 , \38643 );
nand \g447342/U$1 ( \38645 , \38630 , \38638 , \38641 , \38644 );
nor \g446105/U$1 ( \38646 , \38625 , \38626 , \38645 );
and \g452278/U$2 ( \38647 , \16361 , RIe1687e0_2566);
and \g452278/U$3 ( \38648 , RIde82790_226, \16432 );
nor \g452278/U$1 ( \38649 , \38647 , \38648 );
and \g452277/U$2 ( \38650 , \16364 , RIe16a130_2584);
and \g452277/U$3 ( \38651 , RIfc5dc38_6089, \16371 );
nor \g452277/U$1 ( \38652 , \38650 , \38651 );
and \g445227/U$2 ( \38653 , \38646 , \38649 , \38652 );
nor \g445227/U$1 ( \38654 , \38653 , \16649 );
or \g444217/U$1 ( \38655 , \38595 , \38624 , \38654 );
_DC \g62df/U$1 ( \38656 , \38655 , \16652 );
and \g452347/U$2 ( \38657 , \8523 , RIe1cd370_3712);
and \g452347/U$3 ( \38658 , RIe1d0070_3744, \8486 );
nor \g452347/U$1 ( \38659 , \38657 , \38658 );
and \g446119/U$2 ( \38660 , RIe1db470_3872, \8414 );
and \g446119/U$3 ( \38661 , RIe1ca670_3680, \8356 );
and \g449033/U$2 ( \38662 , RIe1de170_3904, \8409 );
and \g449033/U$3 ( \38663 , \8373 , RIe1e6870_4000);
and \g449033/U$4 ( \38664 , RIe1e9570_4032, \8383 );
nor \g449033/U$1 ( \38665 , \38662 , \38663 , \38664 );
and \g452352/U$2 ( \38666 , \8335 , RIe1bf270_3552);
and \g452352/U$3 ( \38667 , RIe1c7970_3648, \8340 );
nor \g452352/U$1 ( \38668 , \38666 , \38667 );
and \g452350/U$2 ( \38669 , \8404 , RIe1e3b70_3968);
and \g452350/U$3 ( \38670 , RIe1ec270_4064, \8351 );
nor \g452350/U$1 ( \38671 , \38669 , \38670 );
and \g454815/U$2 ( \38672 , \8313 , RIe1c1f70_3584);
and \g454815/U$3 ( \38673 , RIe1c4c70_3616, \8323 );
nor \g454815/U$1 ( \38674 , \38672 , \38673 );
not \g454814/U$1 ( \38675 , \38674 );
and \g450046/U$2 ( \38676 , \38675 , \8316 );
and \g450046/U$3 ( \38677 , RIe1e0e70_3936, \8417 );
nor \g450046/U$1 ( \38678 , \38676 , \38677 );
nand \g448192/U$1 ( \38679 , \38665 , \38668 , \38671 , \38678 );
nor \g446119/U$1 ( \38680 , \38660 , \38661 , \38679 );
and \g452349/U$2 ( \38681 , \8378 , RIe1d8770_3840);
and \g452349/U$3 ( \38682 , RIe1d2d70_3776, \8359 );
nor \g452349/U$1 ( \38683 , \38681 , \38682 );
nand \g445603/U$1 ( \38684 , \38659 , \38680 , \38683 );
and \g444777/U$2 ( \38685 , \38684 , \8478 );
and \g449031/U$2 ( \38686 , RIe1acc88_3343, \8317 );
and \g449031/U$3 ( \38687 , \8326 , RIfcb9588_7131);
and \g449031/U$4 ( \38688 , RIfca6190_6912, \8409 );
nor \g449031/U$1 ( \38689 , \38686 , \38687 , \38688 );
and \g452345/U$2 ( \38690 , \8335 , RIe1ab4a0_3326);
and \g452345/U$3 ( \38691 , RIfcd5350_7448, \8340 );
nor \g452345/U$1 ( \38692 , \38690 , \38691 );
and \g452344/U$2 ( \38693 , \8404 , RIe1b7ae8_3467);
and \g452344/U$3 ( \38694 , RIfc784e8_6391, \8351 );
nor \g452344/U$1 ( \38695 , \38693 , \38694 );
and \g454812/U$2 ( \38696 , \8313 , RIe1b9ca8_3491);
and \g454812/U$3 ( \38697 , RIfcbef88_7195, \8323 );
nor \g454812/U$1 ( \38698 , \38696 , \38697 );
not \g450045/U$3 ( \38699 , \38698 );
not \g450045/U$4 ( \38700 , \8328 );
and \g450045/U$2 ( \38701 , \38699 , \38700 );
and \g450045/U$5 ( \38702 , \8417 , RIfcc20c0_7230);
nor \g450045/U$1 ( \38703 , \38701 , \38702 );
nand \g447743/U$1 ( \38704 , \38689 , \38692 , \38695 , \38703 );
and \g444777/U$3 ( \38705 , \8482 , \38704 );
nor \g444777/U$1 ( \38706 , \38685 , \38705 );
and \g446893/U$2 ( \38707 , \8521 , RIe1b1440_3394);
and \g446893/U$3 ( \38708 , RIe1b2d90_3412, \8525 );
nor \g446893/U$1 ( \38709 , \38707 , \38708 );
and \g446892/U$2 ( \38710 , \10290 , RIfcc5090_7264);
and \g446892/U$3 ( \38711 , RIfcb81d8_7117, \10293 );
nor \g446892/U$1 ( \38712 , \38710 , \38711 );
and \g446894/U$2 ( \38713 , \8974 , RIe1b4410_3428);
and \g446894/U$3 ( \38714 , RIe1b5928_3443, \8976 );
nor \g446894/U$1 ( \38715 , \38713 , \38714 );
nand \g444501/U$1 ( \38716 , \38706 , \38709 , \38712 , \38715 );
and \g452361/U$2 ( \38717 , \8531 , RIfccb468_7335);
and \g452361/U$3 ( \38718 , RIf151f70_5392, \8486 );
nor \g452361/U$1 ( \38719 , \38717 , \38718 );
and \g446121/U$2 ( \38720 , RIfce0e58_7581, \8412 );
and \g446121/U$3 ( \38721 , RIe1f3cc8_4151, \8356 );
and \g449036/U$2 ( \38722 , RIfc4ed28_5919, \8409 );
and \g449036/U$3 ( \38723 , \8373 , RIfcae890_7008);
and \g449036/U$4 ( \38724 , RIf157f10_5460, \8383 );
nor \g449036/U$1 ( \38725 , \38722 , \38723 , \38724 );
and \g452364/U$2 ( \38726 , \8335 , RIe1ee9d0_4092);
and \g452364/U$3 ( \38727 , RIfc68ed0_6216, \8340 );
nor \g452364/U$1 ( \38728 , \38726 , \38727 );
and \g452363/U$2 ( \38729 , \8404 , RIe1faa78_4229);
and \g452363/U$3 ( \38730 , RIf159158_5473, \8351 );
nor \g452363/U$1 ( \38731 , \38729 , \38730 );
and \g454819/U$2 ( \38732 , \8313 , RIfca9ca0_6954);
and \g454819/U$3 ( \38733 , RIfc6d250_6264, \8323 );
nor \g454819/U$1 ( \38734 , \38732 , \38733 );
not \g454818/U$1 ( \38735 , \38734 );
and \g450049/U$2 ( \38736 , \38735 , \8316 );
and \g450049/U$3 ( \38737 , RIfc4a840_5870, \8417 );
nor \g450049/U$1 ( \38738 , \38736 , \38737 );
nand \g448193/U$1 ( \38739 , \38725 , \38728 , \38731 , \38738 );
nor \g446121/U$1 ( \38740 , \38720 , \38721 , \38739 );
and \g452362/U$2 ( \38741 , \8378 , RIe1f5ff0_4176);
and \g452362/U$3 ( \38742 , RIf153758_5409, \8359 );
nor \g452362/U$1 ( \38743 , \38741 , \38742 );
nand \g445606/U$1 ( \38744 , \38719 , \38740 , \38743 );
and \g444844/U$2 ( \38745 , \38744 , \8752 );
and \g449034/U$2 ( \38746 , RIe1bc570_3520, \8324 );
and \g449034/U$3 ( \38747 , \8531 , RIe1f8a20_4206);
and \g449034/U$4 ( \38748 , RIe1ff668_4283, \8488 );
nor \g449034/U$1 ( \38749 , \38746 , \38747 , \38748 );
and \g452357/U$2 ( \38750 , \8356 , RIe1f1568_4123);
and \g452357/U$3 ( \38751 , RIe205608_4351, \8359 );
nor \g452357/U$1 ( \38752 , \38750 , \38751 );
and \g454817/U$2 ( \38753 , \8313 , RIe227208_4735);
and \g454817/U$3 ( \38754 , RIe1798b0_2760, \8323 );
nor \g454817/U$1 ( \38755 , \38753 , \38754 );
not \g450048/U$3 ( \38756 , \38755 );
not \g450048/U$4 ( \38757 , \8376 );
and \g450048/U$2 ( \38758 , \38756 , \38757 );
and \g450048/U$5 ( \38759 , \8340 , RIe1d5a70_3808);
nor \g450048/U$1 ( \38760 , \38758 , \38759 );
and \g452356/U$2 ( \38761 , \8378 , RIe21be08_4607);
and \g452356/U$3 ( \38762 , RIe18d3b0_2984, \8417 );
nor \g452356/U$1 ( \38763 , \38761 , \38762 );
nand \g447745/U$1 ( \38764 , \38749 , \38752 , \38760 , \38763 );
and \g444844/U$3 ( \38765 , \9010 , \38764 );
nor \g444844/U$1 ( \38766 , \38745 , \38765 );
and \g446899/U$2 ( \38767 , \9041 , RIe1a0eb0_3208);
and \g446899/U$3 ( \38768 , RIe1a3bb0_3240, \9043 );
nor \g446899/U$1 ( \38769 , \38767 , \38768 );
and \g446898/U$2 ( \38770 , \14956 , RIe1a68b0_3272);
and \g446898/U$3 ( \38771 , RIe1a95b0_3304, \14958 );
nor \g446898/U$1 ( \38772 , \38770 , \38771 );
and \g446900/U$2 ( \38773 , \13244 , RIe171a20_2670);
and \g446900/U$3 ( \38774 , RIe1af3e8_3371, \13246 );
nor \g446900/U$1 ( \38775 , \38773 , \38774 );
nand \g444614/U$1 ( \38776 , \38766 , \38769 , \38772 , \38775 );
and \g446117/U$2 ( \38777 , RIfce8040_7662, \8378 );
and \g446117/U$3 ( \38778 , RIee3c6b8_5146, \8359 );
and \g449027/U$2 ( \38779 , RIfcc4820_7258, \8409 );
and \g449027/U$3 ( \38780 , \8371 , RIe177420_2734);
and \g449027/U$4 ( \38781 , RIfc9e030_6820, \8383 );
nor \g449027/U$1 ( \38782 , \38779 , \38780 , \38781 );
and \g452333/U$2 ( \38783 , \8335 , RIfc472d0_5832);
and \g452333/U$3 ( \38784 , RIfcd3028_7423, \8340 );
nor \g452333/U$1 ( \38785 , \38783 , \38784 );
and \g452332/U$2 ( \38786 , \8404 , RIe176340_2722);
and \g452332/U$3 ( \38787 , RIfc9d0b8_6809, \8351 );
nor \g452332/U$1 ( \38788 , \38786 , \38787 );
and \g454328/U$2 ( \38789 , \8313 , RIfc46a60_5826);
and \g454328/U$3 ( \38790 , RIfc7f400_6470, \8323 );
nor \g454328/U$1 ( \38791 , \38789 , \38790 );
not \g454327/U$1 ( \38792 , \38791 );
and \g450041/U$2 ( \38793 , \38792 , \8316 );
and \g450041/U$3 ( \38794 , RIfc4f700_5926, \8417 );
nor \g450041/U$1 ( \38795 , \38793 , \38794 );
nand \g448191/U$1 ( \38796 , \38782 , \38785 , \38788 , \38795 );
nor \g446117/U$1 ( \38797 , \38777 , \38778 , \38796 );
and \g452331/U$2 ( \38798 , \8356 , RIe174180_2698);
and \g452331/U$3 ( \38799 , RIfc4fb38_5929, \8414 );
nor \g452331/U$1 ( \38800 , \38798 , \38799 );
and \g452330/U$2 ( \38801 , \8523 , RIfc812f0_6492);
and \g452330/U$3 ( \38802 , RIee3b308_5132, \8488 );
nor \g452330/U$1 ( \38803 , \38801 , \38802 );
and \g445234/U$2 ( \38804 , \38797 , \38800 , \38803 );
nor \g445234/U$1 ( \38805 , \38804 , \8558 );
and \g446118/U$2 ( \38806 , RIe192db0_3048, \8414 );
and \g446118/U$3 ( \38807 , RIe184cb0_2888, \8356 );
and \g449028/U$2 ( \38808 , RIe17f2b0_2824, \8317 );
and \g449028/U$3 ( \38809 , \8326 , RIe181fb0_2856);
and \g449028/U$4 ( \38810 , RIe195ab0_3080, \8407 );
nor \g449028/U$1 ( \38811 , \38808 , \38809 , \38810 );
and \g452342/U$2 ( \38812 , \8335 , RIe17c5b0_2792);
and \g452342/U$3 ( \38813 , RIfc83a50_6520, \8340 );
nor \g452342/U$1 ( \38814 , \38812 , \38813 );
and \g452341/U$2 ( \38815 , \8404 , RIe1987b0_3112);
and \g452341/U$3 ( \38816 , RIe19e1b0_3176, \8351 );
nor \g452341/U$1 ( \38817 , \38815 , \38816 );
and \g454808/U$2 ( \38818 , \8313 , RIfc9cf50_6808);
and \g454808/U$3 ( \38819 , RIe19b4b0_3144, \8323 );
nor \g454808/U$1 ( \38820 , \38818 , \38819 );
not \g450043/U$3 ( \38821 , \38820 );
not \g450043/U$4 ( \38822 , \8328 );
and \g450043/U$2 ( \38823 , \38821 , \38822 );
and \g450043/U$5 ( \38824 , \8417 , RIfc87290_6560);
nor \g450043/U$1 ( \38825 , \38823 , \38824 );
nand \g447742/U$1 ( \38826 , \38811 , \38814 , \38817 , \38825 );
nor \g446118/U$1 ( \38827 , \38806 , \38807 , \38826 );
and \g452339/U$2 ( \38828 , \8378 , RIe1900b0_3016);
and \g452339/U$3 ( \38829 , RIe18a6b0_2952, \8359 );
nor \g452339/U$1 ( \38830 , \38828 , \38829 );
and \g452337/U$2 ( \38831 , \8531 , RIfc842c0_6526);
and \g452337/U$3 ( \38832 , RIe1879b0_2920, \8486 );
nor \g452337/U$1 ( \38833 , \38831 , \38832 );
and \g445235/U$2 ( \38834 , \38827 , \38830 , \38833 );
nor \g445235/U$1 ( \38835 , \38834 , \8589 );
or \g444397/U$1 ( \38836 , \38716 , \38776 , \38805 , \38835 );
and \g446114/U$2 ( \38837 , RIfcc81c8_7299, \8414 );
and \g446114/U$3 ( \38838 , RIfea46e8_8215, \8356 );
and \g449023/U$2 ( \38839 , RIfcd19a8_7407, \8409 );
and \g449023/U$3 ( \38840 , \8371 , RIfea9b48_8247);
and \g449023/U$4 ( \38841 , RIfc59cf0_6044, \8330 );
nor \g449023/U$1 ( \38842 , \38839 , \38840 , \38841 );
and \g452323/U$2 ( \38843 , \8335 , RIfc7c430_6436);
and \g452323/U$3 ( \38844 , RIfc77f48_6387, \8340 );
nor \g452323/U$1 ( \38845 , \38843 , \38844 );
and \g452322/U$2 ( \38846 , \8404 , RIfea4418_8213);
and \g452322/U$3 ( \38847 , RIfc7b080_6422, \8351 );
nor \g452322/U$1 ( \38848 , \38846 , \38847 );
and \g454799/U$2 ( \38849 , \8313 , RIf15aaa8_5491);
and \g454799/U$3 ( \38850 , RIfc41fd8_5773, \8323 );
nor \g454799/U$1 ( \38851 , \38849 , \38850 );
not \g454798/U$1 ( \38852 , \38851 );
and \g450039/U$2 ( \38853 , \38852 , \8316 );
and \g450039/U$3 ( \38854 , RIfc79cd0_6408, \8417 );
nor \g450039/U$1 ( \38855 , \38853 , \38854 );
nand \g448190/U$1 ( \38856 , \38842 , \38845 , \38848 , \38855 );
nor \g446114/U$1 ( \38857 , \38837 , \38838 , \38856 );
and \g452320/U$2 ( \38858 , \8378 , RIf162230_5576);
and \g452320/U$3 ( \38859 , RIf160778_5557, \8359 );
nor \g452320/U$1 ( \38860 , \38858 , \38859 );
and \g452319/U$2 ( \38861 , \8531 , RIfea4580_8214);
and \g452319/U$3 ( \38862 , RIf15e888_5535, \8486 );
nor \g452319/U$1 ( \38863 , \38861 , \38862 );
and \g445231/U$2 ( \38864 , \38857 , \38860 , \38863 );
nor \g445231/U$1 ( \38865 , \38864 , \8422 );
and \g446115/U$2 ( \38866 , RIf16cc58_5697, \8351 );
and \g446115/U$3 ( \38867 , RIe221808_4671, \8404 );
and \g449025/U$2 ( \38868 , RIe219108_4575, \8412 );
and \g449025/U$3 ( \38869 , \8409 , RIe21eb08_4639);
and \g449025/U$4 ( \38870 , RIe20dd08_4447, \8326 );
nor \g449025/U$1 ( \38871 , \38868 , \38869 , \38870 );
and \g452327/U$2 ( \38872 , \8356 , RIe210a08_4479);
and \g452327/U$3 ( \38873 , RIfcdbe30_7524, \8359 );
nor \g452327/U$1 ( \38874 , \38872 , \38873 );
and \g454803/U$2 ( \38875 , \8313 , RIf169580_5658);
and \g454803/U$3 ( \38876 , RIe213708_4511, \8323 );
nor \g454803/U$1 ( \38877 , \38875 , \38876 );
not \g450040/U$3 ( \38878 , \38877 );
not \g450040/U$4 ( \38879 , \8347 );
and \g450040/U$2 ( \38880 , \38878 , \38879 );
and \g450040/U$5 ( \38881 , \8340 , RIfca4570_6892);
nor \g450040/U$1 ( \38882 , \38880 , \38881 );
and \g452326/U$2 ( \38883 , \8378 , RIe216408_4543);
and \g452326/U$3 ( \38884 , RIfc97c58_6749, \8417 );
nor \g452326/U$1 ( \38885 , \38883 , \38884 );
nand \g447739/U$1 ( \38886 , \38871 , \38874 , \38882 , \38885 );
nor \g446115/U$1 ( \38887 , \38866 , \38867 , \38886 );
and \g452325/U$2 ( \38888 , \8335 , RIe208308_4383);
and \g452325/U$3 ( \38889 , RIe224508_4703, \8383 );
nor \g452325/U$1 ( \38890 , \38888 , \38889 );
and \g452324/U$2 ( \38891 , \8317 , RIe20b008_4415);
and \g452324/U$3 ( \38892 , RIfc7d3a8_6447, \8373 );
nor \g452324/U$1 ( \38893 , \38891 , \38892 );
and \g445233/U$2 ( \38894 , \38887 , \38890 , \38893 );
nor \g445233/U$1 ( \38895 , \38894 , \8368 );
or \g444243/U$1 ( \38896 , \38836 , \38865 , \38895 );
_DC \g6363/U$1 ( \38897 , \38896 , \8654 );
and \g452708/U$2 ( \38898 , \16377 , RIdec07e8_654);
and \g452708/U$3 ( \38899 , RIdebade8_590, \16380 );
nor \g452708/U$1 ( \38900 , \38898 , \38899 );
and \g446196/U$2 ( \38901 , RIdec34e8_686, \16321 );
and \g446196/U$3 ( \38902 , RIee20620_4827, \16313 );
and \g449130/U$2 ( \38903 , RIdeac4f0_430, \16398 );
and \g449130/U$3 ( \38904 , \16341 , RIee1dec0_4799);
and \g449130/U$4 ( \38905 , RIdebdae8_622, \16344 );
nor \g449130/U$1 ( \38906 , \38903 , \38904 , \38905 );
and \g455347/U$2 ( \38907 , \16317 , RIdeb26e8_494);
and \g455347/U$3 ( \38908 , RIfc41150_5766, \16325 );
nor \g455347/U$1 ( \38909 , \38907 , \38908 );
not \g450144/U$3 ( \38910 , \38909 );
not \g450144/U$4 ( \38911 , \16351 );
and \g450144/U$2 ( \38912 , \38910 , \38911 );
and \g450144/U$5 ( \38913 , \16356 , RIfc4b7b8_5881);
nor \g450144/U$1 ( \38914 , \38912 , \38913 );
and \g452711/U$2 ( \38915 , \16361 , RIde9f2f0_366);
and \g452711/U$3 ( \38916 , RIdea5bf0_398, \16364 );
nor \g452711/U$1 ( \38917 , \38915 , \38916 );
and \g452710/U$2 ( \38918 , \16368 , RIdeaf9e8_462);
and \g452710/U$3 ( \38919 , RIfc87830_6564, \16371 );
nor \g452710/U$1 ( \38920 , \38918 , \38919 );
nand \g447791/U$1 ( \38921 , \38906 , \38914 , \38917 , \38920 );
nor \g446196/U$1 ( \38922 , \38901 , \38902 , \38921 );
and \g452707/U$2 ( \38923 , \16334 , RIdeb80e8_558);
and \g452707/U$3 ( \38924 , RIdec61e8_718, \16328 );
nor \g452707/U$1 ( \38925 , \38923 , \38924 );
nand \g445623/U$1 ( \38926 , \38900 , \38922 , \38925 );
and \g444734/U$2 ( \38927 , \38926 , \17938 );
and \g449129/U$2 ( \38928 , RIfcb7ad0_7112, \16321 );
and \g449129/U$3 ( \38929 , \16328 , RIfcea4d0_7688);
and \g449129/U$4 ( \38930 , RIdf33fb8_1968, \16398 );
nor \g449129/U$1 ( \38931 , \38928 , \38929 , \38930 );
and \g455352/U$2 ( \38932 , \16317 , RIe13f728_2099);
and \g455352/U$3 ( \38933 , RIe141a50_2124, \16325 );
nor \g455352/U$1 ( \38934 , \38932 , \38933 );
not \g450143/U$3 ( \38935 , \38934 );
not \g450143/U$4 ( \38936 , \16330 );
and \g450143/U$2 ( \38937 , \38935 , \38936 );
and \g450143/U$5 ( \38938 , \16339 , RIdf36448_1994);
nor \g450143/U$1 ( \38939 , \38937 , \38938 );
and \g452702/U$2 ( \38940 , \16377 , RIfc51a28_5951);
and \g452702/U$3 ( \38941 , RIfc695d8_6221, \16313 );
nor \g452702/U$1 ( \38942 , \38940 , \38941 );
and \g452703/U$2 ( \38943 , \16334 , RIdf3b1a0_2049);
and \g452703/U$3 ( \38944 , RIdf3d630_2075, \16380 );
nor \g452703/U$1 ( \38945 , \38943 , \38944 );
nand \g447371/U$1 ( \38946 , \38931 , \38939 , \38942 , \38945 );
and \g444734/U$3 ( \38947 , \16394 , \38946 );
nor \g444734/U$1 ( \38948 , \38927 , \38947 );
and \g446967/U$2 ( \38949 , \16419 , RIfea2258_8189);
and \g446967/U$3 ( \38950 , RIdf31df8_1944, \16422 );
nor \g446967/U$1 ( \38951 , \38949 , \38950 );
and \g446965/U$2 ( \38952 , \16429 , RIee2fda0_5003);
and \g446965/U$3 ( \38953 , RIfca9e08_6955, \16434 );
nor \g446965/U$1 ( \38954 , \38952 , \38953 );
and \g446966/U$2 ( \38955 , \16438 , RIee2da78_4978);
and \g446966/U$3 ( \38956 , RIfc88a78_6577, \16441 );
nor \g446966/U$1 ( \38957 , \38955 , \38956 );
nand \g444510/U$1 ( \38958 , \38948 , \38951 , \38954 , \38957 );
and \g452721/U$2 ( \38959 , \16364 , RIfea23c0_8190);
and \g452721/U$3 ( \38960 , RIfcbd7a0_7178, \16371 );
nor \g452721/U$1 ( \38961 , \38959 , \38960 );
and \g446197/U$2 ( \38962 , RIfcb35e8_7063, \16427 );
and \g446197/U$3 ( \38963 , RIfc91178_6673, \16368 );
and \g449134/U$2 ( \38964 , RIfc57f68_6023, \16319 );
and \g449134/U$3 ( \38965 , \16328 , RIfcd1f48_7411);
and \g449134/U$4 ( \38966 , RIded7df8_920, \16398 );
nor \g449134/U$1 ( \38967 , \38964 , \38965 , \38966 );
and \g454975/U$2 ( \38968 , \16317 , RIfea2690_8192);
and \g454975/U$3 ( \38969 , RIdee5520_1073, \16325 );
nor \g454975/U$1 ( \38970 , \38968 , \38969 );
not \g450148/U$3 ( \38971 , \38970 );
not \g450148/U$4 ( \38972 , \16330 );
and \g450148/U$2 ( \38973 , \38971 , \38972 );
and \g450148/U$5 ( \38974 , \16341 , RIfea2528_8191);
nor \g450148/U$1 ( \38975 , \38973 , \38974 );
and \g452724/U$2 ( \38976 , \16377 , RIfcd8fc8_7491);
and \g452724/U$3 ( \38977 , RIfcbe2e0_7186, \16313 );
nor \g452724/U$1 ( \38978 , \38976 , \38977 );
and \g452725/U$2 ( \38979 , \16334 , RIdedf418_1004);
and \g452725/U$3 ( \38980 , RIdee1470_1027, \16380 );
nor \g452725/U$1 ( \38981 , \38979 , \38980 );
nand \g447375/U$1 ( \38982 , \38967 , \38975 , \38978 , \38981 );
nor \g446197/U$1 ( \38983 , \38962 , \38963 , \38982 );
and \g452722/U$2 ( \38984 , \16361 , RIded3910_871);
and \g452722/U$3 ( \38985 , RIfc57b30_6020, \16432 );
nor \g452722/U$1 ( \38986 , \38984 , \38985 );
nand \g445624/U$1 ( \38987 , \38961 , \38983 , \38986 );
and \g444919/U$2 ( \38988 , \38987 , \16477 );
and \g449132/U$2 ( \38989 , RIde989f0_334, \16485 );
and \g449132/U$3 ( \38990 , \16354 , RIdeb53e8_526);
and \g449132/U$4 ( \38991 , RIdee80b8_1104, \16398 );
nor \g449132/U$1 ( \38992 , \38989 , \38990 , \38991 );
and \g454972/U$2 ( \38993 , \16317 , RIdece8e8_814);
and \g454972/U$3 ( \38994 , RIded15e8_846, \16325 );
nor \g454972/U$1 ( \38995 , \38993 , \38994 );
not \g450146/U$3 ( \38996 , \38995 );
not \g450146/U$4 ( \38997 , \16311 );
and \g450146/U$2 ( \38998 , \38996 , \38997 );
and \g450146/U$5 ( \38999 , \16341 , RIdf015b8_1392);
nor \g450146/U$1 ( \39000 , \38998 , \38999 );
and \g452718/U$2 ( \39001 , \16377 , RIdec8ee8_750);
and \g452718/U$3 ( \39002 , RIdecbbe8_782, \16313 );
nor \g452718/U$1 ( \39003 , \39001 , \39002 );
and \g452719/U$2 ( \39004 , \16334 , RIe15ade8_2411);
and \g452719/U$3 ( \39005 , RIe16eff0_2640, \16380 );
nor \g452719/U$1 ( \39006 , \39004 , \39005 );
nand \g447374/U$1 ( \39007 , \38992 , \39000 , \39003 , \39006 );
and \g444919/U$3 ( \39008 , \16752 , \39007 );
nor \g444919/U$1 ( \39009 , \38988 , \39008 );
and \g446970/U$2 ( \39010 , \16774 , RIde7e938_207);
and \g446970/U$3 ( \39011 , RIdedce20_977, \16776 );
nor \g446970/U$1 ( \39012 , \39010 , \39011 );
and \g446969/U$2 ( \39013 , \16779 , RIdf1dec0_1717);
and \g446969/U$3 ( \39014 , RIdf2d640_1893, \16781 );
nor \g446969/U$1 ( \39015 , \39013 , \39014 );
and \g446968/U$2 ( \39016 , \16784 , RIdf38fe0_2025);
and \g446968/U$3 ( \39017 , RIe1445e8_2155, \16786 );
nor \g446968/U$1 ( \39018 , \39016 , \39017 );
nand \g444629/U$1 ( \39019 , \39009 , \39012 , \39015 , \39018 );
and \g446190/U$2 ( \39020 , RIfc77c78_6385, \16319 );
and \g446190/U$3 ( \39021 , RIfc84f68_6535, \16313 );
and \g449124/U$2 ( \39022 , RIee19f78_4754, \16427 );
and \g449124/U$3 ( \39023 , \16432 , RIee1a680_4759);
and \g449124/U$4 ( \39024 , RIde8efb8_287, \16485 );
nor \g449124/U$1 ( \39025 , \39022 , \39023 , \39024 );
and \g454966/U$2 ( \39026 , \16317 , RIe16c2f0_2608);
and \g454966/U$3 ( \39027 , RIfc76328_6367, \16325 );
nor \g454966/U$1 ( \39028 , \39026 , \39027 );
not \g454965/U$1 ( \39029 , \39028 );
and \g450138/U$2 ( \39030 , \39029 , \16336 );
and \g450138/U$3 ( \39031 , RIde92780_304, \16356 );
nor \g450138/U$1 ( \39032 , \39030 , \39031 );
and \g452692/U$2 ( \39033 , \16361 , RIfea20f0_8188);
and \g452692/U$3 ( \39034 , RIee388d8_5102, \16364 );
nor \g452692/U$1 ( \39035 , \39033 , \39034 );
and \g452690/U$2 ( \39036 , \16368 , RIfcbeb50_7192);
and \g452690/U$3 ( \39037 , RIfcd7240_7470, \16371 );
nor \g452690/U$1 ( \39038 , \39036 , \39037 );
nand \g448087/U$1 ( \39039 , \39025 , \39032 , \39035 , \39038 );
nor \g446190/U$1 ( \39040 , \39020 , \39021 , \39039 );
and \g452686/U$2 ( \39041 , \16377 , RIfc6ff50_6296);
and \g452686/U$3 ( \39042 , RIde8ae18_267, \16380 );
nor \g452686/U$1 ( \39043 , \39041 , \39042 );
and \g452684/U$2 ( \39044 , \16334 , RIde86c78_247);
and \g452684/U$3 ( \39045 , RIee1d380_4791, \16328 );
nor \g452684/U$1 ( \39046 , \39044 , \39045 );
and \g445290/U$2 ( \39047 , \39040 , \39043 , \39046 );
nor \g445290/U$1 ( \39048 , \39047 , \16649 );
and \g446192/U$2 ( \39049 , RIe1634e8_2507, \16321 );
and \g446192/U$3 ( \39050 , RIee37c30_5093, \16313 );
and \g449126/U$2 ( \39051 , RIe14cce8_2251, \16398 );
and \g449126/U$3 ( \39052 , \16341 , RIfc83e88_6523);
and \g449126/U$4 ( \39053 , RIe15dae8_2443, \16485 );
nor \g449126/U$1 ( \39054 , \39051 , \39052 , \39053 );
and \g454968/U$2 ( \39055 , \16317 , RIe1526e8_2315);
and \g454968/U$3 ( \39056 , RIfc3f698_5747, \16325 );
nor \g454968/U$1 ( \39057 , \39055 , \39056 );
not \g450141/U$3 ( \39058 , \39057 );
not \g450141/U$4 ( \39059 , \16351 );
and \g450141/U$2 ( \39060 , \39058 , \39059 );
and \g450141/U$5 ( \39061 , \16356 , RIfce7500_7654);
nor \g450141/U$1 ( \39062 , \39060 , \39061 );
and \g452697/U$2 ( \39063 , \16361 , RIe1472e8_2187);
and \g452697/U$3 ( \39064 , RIe149fe8_2219, \16364 );
nor \g452697/U$1 ( \39065 , \39063 , \39064 );
and \g452696/U$2 ( \39066 , \16368 , RIe14f9e8_2283);
and \g452696/U$3 ( \39067 , RIee354d0_5065, \16371 );
nor \g452696/U$1 ( \39068 , \39066 , \39067 );
nand \g447789/U$1 ( \39069 , \39054 , \39062 , \39065 , \39068 );
nor \g446192/U$1 ( \39070 , \39049 , \39050 , \39069 );
and \g452695/U$2 ( \39071 , \16377 , RIe1607e8_2475);
and \g452695/U$3 ( \39072 , RIe1580e8_2379, \16380 );
nor \g452695/U$1 ( \39073 , \39071 , \39072 );
and \g452694/U$2 ( \39074 , \16334 , RIe1553e8_2347);
and \g452694/U$3 ( \39075 , RIe1661e8_2539, \16328 );
nor \g452694/U$1 ( \39076 , \39074 , \39075 );
and \g445291/U$2 ( \39077 , \39070 , \39073 , \39076 );
nor \g445291/U$1 ( \39078 , \39077 , \16389 );
or \g444344/U$1 ( \39079 , \38958 , \39019 , \39048 , \39078 );
and \g446188/U$2 ( \39080 , RIdf150b8_1616, \16321 );
and \g446188/U$3 ( \39081 , RIdf123b8_1584, \16313 );
and \g449121/U$2 ( \39082 , RIdefbbb8_1328, \16427 );
and \g449121/U$3 ( \39083 , \16448 , RIdefe8b8_1360);
and \g449121/U$4 ( \39084 , RIdf09cb8_1488, \16485 );
nor \g449121/U$1 ( \39085 , \39082 , \39083 , \39084 );
and \g454961/U$2 ( \39086 , \16317 , RIdef07b8_1200);
and \g454961/U$3 ( \39087 , RIdef34b8_1232, \16325 );
nor \g454961/U$1 ( \39088 , \39086 , \39087 );
not \g454960/U$1 ( \39089 , \39088 );
and \g450135/U$2 ( \39090 , \39089 , \16336 );
and \g450135/U$3 ( \39091 , RIdf0c9b8_1520, \16356 );
nor \g450135/U$1 ( \39092 , \39090 , \39091 );
and \g452670/U$2 ( \39093 , \16361 , RIdeeadb8_1136);
and \g452670/U$3 ( \39094 , RIdeedab8_1168, \16364 );
nor \g452670/U$1 ( \39095 , \39093 , \39094 );
and \g452669/U$2 ( \39096 , \16368 , RIdef61b8_1264);
and \g452669/U$3 ( \39097 , RIdef8eb8_1296, \16371 );
nor \g452669/U$1 ( \39098 , \39096 , \39097 );
nand \g448085/U$1 ( \39099 , \39085 , \39092 , \39095 , \39098 );
nor \g446188/U$1 ( \39100 , \39080 , \39081 , \39099 );
and \g452668/U$2 ( \39101 , \16377 , RIdf0f6b8_1552);
and \g452668/U$3 ( \39102 , RIdf06fb8_1456, \16380 );
nor \g452668/U$1 ( \39103 , \39101 , \39102 );
and \g452667/U$2 ( \39104 , \16334 , RIdf042b8_1424);
and \g452667/U$3 ( \39105 , RIdf17db8_1648, \16328 );
nor \g452667/U$1 ( \39106 , \39104 , \39105 );
and \g445285/U$2 ( \39107 , \39100 , \39103 , \39106 );
nor \g445285/U$1 ( \39108 , \39107 , \16555 );
and \g446189/U$2 ( \39109 , RIfca08f8_6849, \16427 );
and \g446189/U$3 ( \39110 , RIfc49058_5853, \16368 );
and \g449122/U$2 ( \39111 , RIdf28d20_1841, \16485 );
and \g449122/U$3 ( \39112 , \16356 , RIdf2ac10_1863);
and \g449122/U$4 ( \39113 , RIdf204b8_1744, \16398 );
nor \g449122/U$1 ( \39114 , \39111 , \39112 , \39113 );
and \g454964/U$2 ( \39115 , \16317 , RIee2aaa8_4944);
and \g454964/U$3 ( \39116 , RIee2c560_4963, \16325 );
nor \g454964/U$1 ( \39117 , \39115 , \39116 );
not \g450136/U$3 ( \39118 , \39117 );
not \g450136/U$4 ( \39119 , \16311 );
and \g450136/U$2 ( \39120 , \39118 , \39119 );
and \g450136/U$5 ( \39121 , \16341 , RIfca0a60_6850);
nor \g450136/U$1 ( \39122 , \39120 , \39121 );
and \g452678/U$2 ( \39123 , \16377 , RIee281e0_4915);
and \g452678/U$3 ( \39124 , RIee29428_4928, \16313 );
nor \g452678/U$1 ( \39125 , \39123 , \39124 );
and \g452679/U$2 ( \39126 , \16334 , RIfea2960_8194);
and \g452679/U$3 ( \39127 , RIfea27f8_8193, \16380 );
nor \g452679/U$1 ( \39128 , \39126 , \39127 );
nand \g447370/U$1 ( \39129 , \39114 , \39122 , \39125 , \39128 );
nor \g446189/U$1 ( \39130 , \39109 , \39110 , \39129 );
and \g452676/U$2 ( \39131 , \16361 , RIdf19f78_1672);
and \g452676/U$3 ( \39132 , RIfcdabe8_7511, \16448 );
nor \g452676/U$1 ( \39133 , \39131 , \39132 );
and \g452675/U$2 ( \39134 , \16364 , RIfc99cb0_6772);
and \g452675/U$3 ( \39135 , RIfc8b1d8_6605, \16371 );
nor \g452675/U$1 ( \39136 , \39134 , \39135 );
and \g445288/U$2 ( \39137 , \39130 , \39133 , \39136 );
nor \g445288/U$1 ( \39138 , \39137 , \16480 );
or \g444262/U$1 ( \39139 , \39079 , \39108 , \39138 );
_DC \g63e8/U$1 ( \39140 , \39139 , \16652 );
and \g452763/U$2 ( \39141 , \8326 , RIe1bc840_3522);
and \g452763/U$3 ( \39142 , RIe1f1838_4125, \8356 );
nor \g452763/U$1 ( \39143 , \39141 , \39142 );
and \g446207/U$2 ( \39144 , RIe1f8cf0_4208, \8523 );
and \g446207/U$3 ( \39145 , RIe1af6b8_3373, \8319 );
and \g449144/U$2 ( \39146 , RIe1a3e80_3242, \8373 );
and \g449144/U$3 ( \39147 , \8383 , RIe1a6b80_3274);
and \g449144/U$4 ( \39148 , RIe1ff938_4285, \8488 );
nor \g449144/U$1 ( \39149 , \39146 , \39147 , \39148 );
and \g455214/U$2 ( \39150 , \8313 , RIe2274d8_4737);
and \g455214/U$3 ( \39151 , RIe179b80_2762, \8323 );
nor \g455214/U$1 ( \39152 , \39150 , \39151 );
not \g450159/U$3 ( \39153 , \39152 );
not \g450159/U$4 ( \39154 , \8376 );
and \g450159/U$2 ( \39155 , \39153 , \39154 );
and \g450159/U$5 ( \39156 , \8359 , RIe2058d8_4353);
nor \g450159/U$1 ( \39157 , \39155 , \39156 );
and \g452767/U$2 ( \39158 , \8404 , RIe1a1180_3210);
and \g452767/U$3 ( \39159 , RIe1a9880_3306, \8351 );
nor \g452767/U$1 ( \39160 , \39158 , \39159 );
and \g452768/U$2 ( \39161 , \8378 , RIe21c0d8_4609);
and \g452768/U$3 ( \39162 , RIe18d680_2986, \8417 );
nor \g452768/U$1 ( \39163 , \39161 , \39162 );
nand \g447797/U$1 ( \39164 , \39149 , \39157 , \39160 , \39163 );
nor \g446207/U$1 ( \39165 , \39144 , \39145 , \39164 );
and \g452765/U$2 ( \39166 , \8335 , RIe171cf0_2672);
and \g452765/U$3 ( \39167 , RIe1d5d40_3810, \8340 );
nor \g452765/U$1 ( \39168 , \39166 , \39167 );
nand \g445626/U$1 ( \39169 , \39143 , \39165 , \39168 );
and \g444880/U$2 ( \39170 , \39169 , \9010 );
and \g449142/U$2 ( \39171 , RIfc65f00_6182, \8319 );
and \g449142/U$3 ( \39172 , \8326 , RIfcad378_6993);
and \g449142/U$4 ( \39173 , RIfc71030_6308, \8383 );
nor \g449142/U$1 ( \39174 , \39171 , \39172 , \39173 );
and \g452761/U$2 ( \39175 , \8335 , RIe1eeca0_4094);
and \g452761/U$3 ( \39176 , RIfcde158_7549, \8340 );
nor \g452761/U$1 ( \39177 , \39175 , \39176 );
and \g454997/U$2 ( \39178 , \8313 , RIfc6f578_6289);
and \g454997/U$3 ( \39179 , RIfc6fde8_6295, \8323 );
nor \g454997/U$1 ( \39180 , \39178 , \39179 );
not \g450158/U$3 ( \39181 , \39180 );
not \g450158/U$4 ( \39182 , \8347 );
and \g450158/U$2 ( \39183 , \39181 , \39182 );
and \g450158/U$5 ( \39184 , \8351 , RIfc4ca00_5894);
nor \g450158/U$1 ( \39185 , \39183 , \39184 );
and \g452759/U$2 ( \39186 , \8356 , RIe1f3f98_4153);
and \g452759/U$3 ( \39187 , RIfcada80_6998, \8359 );
nor \g452759/U$1 ( \39188 , \39186 , \39187 );
nand \g447796/U$1 ( \39189 , \39174 , \39177 , \39185 , \39188 );
and \g444880/U$3 ( \39190 , \8752 , \39189 );
nor \g444880/U$1 ( \39191 , \39170 , \39190 );
and \g446978/U$2 ( \39192 , \11511 , RIe1fad48_4231);
and \g446978/U$3 ( \39193 , RIfcde428_7551, \11513 );
nor \g446978/U$1 ( \39194 , \39192 , \39193 );
and \g446979/U$2 ( \39195 , \11516 , RIfc63a70_6156);
and \g446979/U$3 ( \39196 , RIfc70bf8_6305, \11518 );
nor \g446979/U$1 ( \39197 , \39195 , \39196 );
and \g446980/U$2 ( \39198 , \11521 , RIe1f62c0_4178);
and \g446980/U$3 ( \39199 , RIfca7db0_6932, \11523 );
nor \g446980/U$1 ( \39200 , \39198 , \39199 );
nand \g444631/U$1 ( \39201 , \39191 , \39194 , \39197 , \39200 );
and \g452777/U$2 ( \39202 , \8324 , RIe20dfd8_4449);
and \g452777/U$3 ( \39203 , RIe210cd8_4481, \8356 );
nor \g452777/U$1 ( \39204 , \39202 , \39203 );
and \g446208/U$2 ( \39205 , RIf169850_5660, \8523 );
and \g446208/U$3 ( \39206 , RIe20b2d8_4417, \8317 );
and \g449148/U$2 ( \39207 , RIe2193d8_4577, \8414 );
and \g449148/U$3 ( \39208 , \8409 , RIe21edd8_4641);
and \g449148/U$4 ( \39209 , RIe2139d8_4513, \8486 );
nor \g449148/U$1 ( \39210 , \39207 , \39208 , \39209 );
and \g455008/U$2 ( \39211 , \8313 , RIfc77138_6377);
and \g455008/U$3 ( \39212 , RIe2247d8_4705, \8323 );
nor \g455008/U$1 ( \39213 , \39211 , \39212 );
not \g450163/U$3 ( \39214 , \39213 );
not \g450163/U$4 ( \39215 , \8328 );
and \g450163/U$2 ( \39216 , \39214 , \39215 );
and \g450163/U$5 ( \39217 , \8359 , RIfc40070_5754);
nor \g450163/U$1 ( \39218 , \39216 , \39217 );
and \g452779/U$2 ( \39219 , \8404 , RIe221ad8_4673);
and \g452779/U$3 ( \39220 , RIfc40bb0_5762, \8351 );
nor \g452779/U$1 ( \39221 , \39219 , \39220 );
and \g452780/U$2 ( \39222 , \8378 , RIe2166d8_4545);
and \g452780/U$3 ( \39223 , RIfcd7d80_7478, \8417 );
nor \g452780/U$1 ( \39224 , \39222 , \39223 );
nand \g447800/U$1 ( \39225 , \39210 , \39218 , \39221 , \39224 );
nor \g446208/U$1 ( \39226 , \39205 , \39206 , \39225 );
and \g452778/U$2 ( \39227 , \8335 , RIe2085d8_4385);
and \g452778/U$3 ( \39228 , RIfcc1580_7222, \8340 );
nor \g452778/U$1 ( \39229 , \39227 , \39228 );
nand \g445628/U$1 ( \39230 , \39204 , \39226 , \39229 );
and \g444853/U$2 ( \39231 , \39230 , \8369 );
and \g449146/U$2 ( \39232 , RIe203010_4324, \8373 );
and \g449146/U$3 ( \39233 , \8383 , RIfc749d8_6349);
and \g449146/U$4 ( \39234 , RIf15eb58_5537, \8488 );
nor \g449146/U$1 ( \39235 , \39232 , \39233 , \39234 );
and \g455224/U$2 ( \39236 , \8313 , RIfcaf970_7020);
and \g455224/U$3 ( \39237 , RIfc60668_6119, \8323 );
nor \g455224/U$1 ( \39238 , \39236 , \39237 );
not \g450161/U$3 ( \39239 , \39238 );
not \g450161/U$4 ( \39240 , \8376 );
and \g450161/U$2 ( \39241 , \39239 , \39240 );
and \g450161/U$5 ( \39242 , \8359 , RIf160a48_5559);
nor \g450161/U$1 ( \39243 , \39241 , \39242 );
and \g452774/U$2 ( \39244 , \8404 , RIe2013f0_4304);
and \g452774/U$3 ( \39245 , RIfcd0058_7389, \8351 );
nor \g452774/U$1 ( \39246 , \39244 , \39245 );
and \g452775/U$2 ( \39247 , \8378 , RIfc45818_5813);
and \g452775/U$3 ( \39248 , RIfc60230_6116, \8417 );
nor \g452775/U$1 ( \39249 , \39247 , \39248 );
nand \g447799/U$1 ( \39250 , \39235 , \39243 , \39246 , \39249 );
and \g444853/U$3 ( \39251 , \9266 , \39250 );
nor \g444853/U$1 ( \39252 , \39231 , \39251 );
and \g446981/U$2 ( \39253 , \10230 , RIfea19e8_8183);
and \g446981/U$3 ( \39254 , RIfea1880_8182, \10232 );
nor \g446981/U$1 ( \39255 , \39253 , \39254 );
and \g446982/U$2 ( \39256 , \13424 , RIfc49b98_5861);
and \g446982/U$3 ( \39257 , RIfc72110_6320, \13426 );
nor \g446982/U$1 ( \39258 , \39256 , \39257 );
and \g446983/U$2 ( \39259 , \9299 , RIfc71738_6313);
and \g446983/U$3 ( \39260 , RIfcca0b8_7321, \9301 );
nor \g446983/U$1 ( \39261 , \39259 , \39260 );
nand \g444632/U$1 ( \39262 , \39252 , \39255 , \39258 , \39261 );
and \g446202/U$2 ( \39263 , RIe1e6b40_4002, \8371 );
and \g446202/U$3 ( \39264 , RIe1d8a40_3842, \8378 );
and \g449139/U$2 ( \39265 , RIe1cd640_3714, \8531 );
and \g449139/U$3 ( \39266 , \8488 , RIe1d0340_3746);
and \g449139/U$4 ( \39267 , RIe1e9840_4034, \8383 );
nor \g449139/U$1 ( \39268 , \39265 , \39266 , \39267 );
and \g452746/U$2 ( \39269 , \8335 , RIe1bf540_3554);
and \g452746/U$3 ( \39270 , RIe1c7c40_3650, \8340 );
nor \g452746/U$1 ( \39271 , \39269 , \39270 );
and \g454986/U$2 ( \39272 , \8313 , RIe1c2240_3586);
and \g454986/U$3 ( \39273 , RIe1c4f40_3618, \8323 );
nor \g454986/U$1 ( \39274 , \39272 , \39273 );
not \g454985/U$1 ( \39275 , \39274 );
and \g450153/U$2 ( \39276 , \39275 , \8316 );
and \g450153/U$3 ( \39277 , RIe1ec540_4066, \8351 );
nor \g450153/U$1 ( \39278 , \39276 , \39277 );
and \g452744/U$2 ( \39279 , \8356 , RIe1ca940_3682);
and \g452744/U$3 ( \39280 , RIe1d3040_3778, \8359 );
nor \g452744/U$1 ( \39281 , \39279 , \39280 );
nand \g448203/U$1 ( \39282 , \39268 , \39271 , \39278 , \39281 );
nor \g446202/U$1 ( \39283 , \39263 , \39264 , \39282 );
and \g452743/U$2 ( \39284 , \8404 , RIe1e3e40_3970);
and \g452743/U$3 ( \39285 , RIe1de440_3906, \8409 );
nor \g452743/U$1 ( \39286 , \39284 , \39285 );
and \g452741/U$2 ( \39287 , \8414 , RIe1db740_3874);
and \g452741/U$3 ( \39288 , RIe1e1140_3938, \8417 );
nor \g452741/U$1 ( \39289 , \39287 , \39288 );
and \g445297/U$2 ( \39290 , \39283 , \39286 , \39289 );
nor \g445297/U$1 ( \39291 , \39290 , \8477 );
and \g446204/U$2 ( \39292 , RIe1b3060_3414, \8531 );
and \g446204/U$3 ( \39293 , RIe1acf58_3345, \8317 );
and \g449141/U$2 ( \39294 , RIe1b5bf8_3445, \8414 );
and \g449141/U$3 ( \39295 , \8409 , RIfc69740_6222);
and \g449141/U$4 ( \39296 , RIf148088_5279, \8488 );
nor \g449141/U$1 ( \39297 , \39294 , \39295 , \39296 );
and \g454990/U$2 ( \39298 , \8313 , RIe1b9f78_3493);
and \g454990/U$3 ( \39299 , RIfccba08_7339, \8323 );
nor \g454990/U$1 ( \39300 , \39298 , \39299 );
not \g450155/U$3 ( \39301 , \39300 );
not \g450155/U$4 ( \39302 , \8328 );
and \g450155/U$2 ( \39303 , \39301 , \39302 );
and \g450155/U$5 ( \39304 , \8359 , RIfccf950_7384);
nor \g450155/U$1 ( \39305 , \39303 , \39304 );
and \g452752/U$2 ( \39306 , \8404 , RIe1b7db8_3469);
and \g452752/U$3 ( \39307 , RIfc69308_6219, \8351 );
nor \g452752/U$1 ( \39308 , \39306 , \39307 );
and \g452753/U$2 ( \39309 , \8378 , RIe1b4578_3429);
and \g452753/U$3 ( \39310 , RIfccd628_7359, \8417 );
nor \g452753/U$1 ( \39311 , \39309 , \39310 );
nand \g447795/U$1 ( \39312 , \39297 , \39305 , \39308 , \39311 );
nor \g446204/U$1 ( \39313 , \39292 , \39293 , \39312 );
and \g452749/U$2 ( \39314 , \8335 , RIe1ab770_3328);
and \g452749/U$3 ( \39315 , RIfc9f818_6837, \8340 );
nor \g452749/U$1 ( \39316 , \39314 , \39315 );
and \g452748/U$2 ( \39317 , \8324 , RIfcb9c90_7136);
and \g452748/U$3 ( \39318 , RIe1b1710_3396, \8356 );
nor \g452748/U$1 ( \39319 , \39317 , \39318 );
and \g445299/U$2 ( \39320 , \39313 , \39316 , \39319 );
nor \g445299/U$1 ( \39321 , \39320 , \8481 );
or \g444336/U$1 ( \39322 , \39201 , \39262 , \39291 , \39321 );
and \g446199/U$2 ( \39323 , RIfcc1148_7219, \8417 );
and \g446199/U$3 ( \39324 , RIe198a80_3114, \8404 );
and \g449136/U$2 ( \39325 , RIfcb2ee0_7058, \8531 );
and \g449136/U$3 ( \39326 , \8488 , RIe187c80_2922);
and \g449136/U$4 ( \39327 , RIe19b780_3146, \8330 );
nor \g449136/U$1 ( \39328 , \39325 , \39326 , \39327 );
and \g452731/U$2 ( \39329 , \8335 , RIe17c880_2794);
and \g452731/U$3 ( \39330 , RIfc615e0_6130, \8340 );
nor \g452731/U$1 ( \39331 , \39329 , \39330 );
and \g454979/U$2 ( \39332 , \8313 , RIe17f580_2826);
and \g454979/U$3 ( \39333 , RIe182280_2858, \8323 );
nor \g454979/U$1 ( \39334 , \39332 , \39333 );
not \g454978/U$1 ( \39335 , \39334 );
and \g450150/U$2 ( \39336 , \39335 , \8316 );
and \g450150/U$3 ( \39337 , RIe19e480_3178, \8351 );
nor \g450150/U$1 ( \39338 , \39336 , \39337 );
and \g452730/U$2 ( \39339 , \8356 , RIe184f80_2890);
and \g452730/U$3 ( \39340 , RIe18a980_2954, \8359 );
nor \g452730/U$1 ( \39341 , \39339 , \39340 );
nand \g448202/U$1 ( \39342 , \39328 , \39331 , \39338 , \39341 );
nor \g446199/U$1 ( \39343 , \39323 , \39324 , \39342 );
and \g452729/U$2 ( \39344 , \8378 , RIe190380_3018);
and \g452729/U$3 ( \39345 , RIfccc980_7350, \8373 );
nor \g452729/U$1 ( \39346 , \39344 , \39345 );
and \g452728/U$2 ( \39347 , \8412 , RIe193080_3050);
and \g452728/U$3 ( \39348 , RIe195d80_3082, \8409 );
nor \g452728/U$1 ( \39349 , \39347 , \39348 );
and \g445293/U$2 ( \39350 , \39343 , \39346 , \39349 );
nor \g445293/U$1 ( \39351 , \39350 , \8589 );
and \g446201/U$2 ( \39352 , RIfea1cb8_8185, \8531 );
and \g446201/U$3 ( \39353 , RIfea1e20_8186, \8319 );
and \g449137/U$2 ( \39354 , RIfc6f2a8_6287, \8373 );
and \g449137/U$3 ( \39355 , \8383 , RIfc4c898_5893);
and \g449137/U$4 ( \39356 , RIfc56e88_6011, \8488 );
nor \g449137/U$1 ( \39357 , \39354 , \39355 , \39356 );
and \g454983/U$2 ( \39358 , \8313 , RIfc70388_6299);
and \g454983/U$3 ( \39359 , RIfc6adc0_6238, \8323 );
nor \g454983/U$1 ( \39360 , \39358 , \39359 );
not \g450151/U$3 ( \39361 , \39360 );
not \g450151/U$4 ( \39362 , \8376 );
and \g450151/U$2 ( \39363 , \39361 , \39362 );
and \g450151/U$5 ( \39364 , \8359 , RIfea1f88_8187);
nor \g450151/U$1 ( \39365 , \39363 , \39364 );
and \g452737/U$2 ( \39366 , \8404 , RIe1764a8_2723);
and \g452737/U$3 ( \39367 , RIfc69038_6217, \8351 );
nor \g452737/U$1 ( \39368 , \39366 , \39367 );
and \g452738/U$2 ( \39369 , \8378 , RIfea1b50_8184);
and \g452738/U$3 ( \39370 , RIfcad0a8_6991, \8417 );
nor \g452738/U$1 ( \39371 , \39369 , \39370 );
nand \g447793/U$1 ( \39372 , \39357 , \39365 , \39368 , \39371 );
nor \g446201/U$1 ( \39373 , \39352 , \39353 , \39372 );
and \g452736/U$2 ( \39374 , \8335 , RIf16d798_5705);
and \g452736/U$3 ( \39375 , RIfc60d70_6124, \8340 );
nor \g452736/U$1 ( \39376 , \39374 , \39375 );
and \g452734/U$2 ( \39377 , \8324 , RIfc6a820_6234);
and \g452734/U$3 ( \39378 , RIe174450_2700, \8356 );
nor \g452734/U$1 ( \39379 , \39377 , \39378 );
and \g445295/U$2 ( \39380 , \39373 , \39376 , \39379 );
nor \g445295/U$1 ( \39381 , \39380 , \8558 );
or \g444279/U$1 ( \39382 , \39322 , \39351 , \39381 );
_DC \g646c/U$1 ( \39383 , \39382 , \8654 );
and \g446209/U$2 ( \39384 , RIdec3650_687, \16319 );
and \g446209/U$3 ( \39385 , RIfcaf3d0_7016, \16313 );
and \g449151/U$2 ( \39386 , RIdeac838_431, \16398 );
and \g449151/U$3 ( \39387 , \16341 , RIfc8c6f0_6620);
and \g449151/U$4 ( \39388 , RIdebdc50_623, \16344 );
nor \g449151/U$1 ( \39389 , \39386 , \39387 , \39388 );
and \g455315/U$2 ( \39390 , \16317 , RIdeb2850_495);
and \g455315/U$3 ( \39391 , RIfc42f50_5784, \16325 );
nor \g455315/U$1 ( \39392 , \39390 , \39391 );
not \g450165/U$3 ( \39393 , \39392 );
not \g450165/U$4 ( \39394 , \16351 );
and \g450165/U$2 ( \39395 , \39393 , \39394 );
and \g450165/U$5 ( \39396 , \16356 , RIfc6a280_6230);
nor \g450165/U$1 ( \39397 , \39395 , \39396 );
and \g452787/U$2 ( \39398 , \16361 , RIde9f638_367);
and \g452787/U$3 ( \39399 , RIdea5f38_399, \16364 );
nor \g452787/U$1 ( \39400 , \39398 , \39399 );
and \g452786/U$2 ( \39401 , \16368 , RIdeafb50_463);
and \g452786/U$3 ( \39402 , RIfc981f8_6753, \16371 );
nor \g452786/U$1 ( \39403 , \39401 , \39402 );
nand \g447802/U$1 ( \39404 , \39389 , \39397 , \39400 , \39403 );
nor \g446209/U$1 ( \39405 , \39384 , \39385 , \39404 );
and \g452784/U$2 ( \39406 , \16377 , RIdec0950_655);
and \g452784/U$3 ( \39407 , RIdebaf50_591, \16380 );
nor \g452784/U$1 ( \39408 , \39406 , \39407 );
and \g452783/U$2 ( \39409 , \16334 , RIdeb8250_559);
and \g452783/U$3 ( \39410 , RIdec6350_719, \16326 );
nor \g452783/U$1 ( \39411 , \39409 , \39410 );
and \g445301/U$2 ( \39412 , \39405 , \39408 , \39411 );
nor \g445301/U$1 ( \39413 , \39412 , \16618 );
and \g446211/U$2 ( \39414 , RIfc89888_6587, \16321 );
and \g446211/U$3 ( \39415 , RIfc8f558_6653, \16313 );
and \g449152/U$2 ( \39416 , RIfc568e8_6007, \16427 );
and \g449152/U$3 ( \39417 , \16448 , RIee30a48_5012);
and \g449152/U$4 ( \39418 , RIe13f890_2100, \16485 );
nor \g449152/U$1 ( \39419 , \39416 , \39417 , \39418 );
and \g455022/U$2 ( \39420 , \16317 , RIfea38d8_8205);
and \g455022/U$3 ( \39421 , RIdf365b0_1995, \16325 );
nor \g455022/U$1 ( \39422 , \39420 , \39421 );
not \g455021/U$1 ( \39423 , \39422 );
and \g450166/U$2 ( \39424 , \39423 , \16336 );
and \g450166/U$3 ( \39425 , RIe141bb8_2125, \16354 );
nor \g450166/U$1 ( \39426 , \39424 , \39425 );
and \g452794/U$2 ( \39427 , \16361 , RIdf2ff08_1922);
and \g452794/U$3 ( \39428 , RIfea3a40_8206, \16364 );
nor \g452794/U$1 ( \39429 , \39427 , \39428 );
and \g452793/U$2 ( \39430 , \16368 , RIee2dbe0_4979);
and \g452793/U$3 ( \39431 , RIee2e9f0_4989, \16371 );
nor \g452793/U$1 ( \39432 , \39430 , \39431 );
nand \g448089/U$1 ( \39433 , \39419 , \39426 , \39429 , \39432 );
nor \g446211/U$1 ( \39434 , \39414 , \39415 , \39433 );
and \g452792/U$2 ( \39435 , \16377 , RIfc52838_5961);
and \g452792/U$3 ( \39436 , RIdf3d798_2076, \16380 );
nor \g452792/U$1 ( \39437 , \39435 , \39436 );
and \g452790/U$2 ( \39438 , \16334 , RIdf3b308_2050);
and \g452790/U$3 ( \39439 , RIfc97f28_6751, \16328 );
nor \g452790/U$1 ( \39440 , \39438 , \39439 );
and \g445302/U$2 ( \39441 , \39434 , \39437 , \39440 );
nor \g445302/U$1 ( \39442 , \39441 , \16393 );
nor \g444672/U$1 ( \39443 , \39413 , \39442 );
and \g446993/U$2 ( \39444 , \22457 , RIe14fb50_2284);
and \g446993/U$3 ( \39445 , RIee35638_5066, \22459 );
nor \g446993/U$1 ( \39446 , \39444 , \39445 );
not \g444413/U$2 ( \39447 , \39446 );
and \g452833/U$2 ( \39448 , \16364 , RIdeedc20_1169);
and \g452833/U$3 ( \39449 , RIdef9020_1297, \16371 );
nor \g452833/U$1 ( \39450 , \39448 , \39449 );
and \g446219/U$2 ( \39451 , RIdefbd20_1329, \16427 );
and \g446219/U$3 ( \39452 , RIdef6320_1265, \16368 );
and \g449164/U$2 ( \39453 , RIdf15220_1617, \16319 );
and \g449164/U$3 ( \39454 , \16328 , RIdf17f20_1649);
and \g449164/U$4 ( \39455 , RIdef0920_1201, \16398 );
nor \g449164/U$1 ( \39456 , \39453 , \39454 , \39455 );
and \g455045/U$2 ( \39457 , \16317 , RIdf09e20_1489);
and \g455045/U$3 ( \39458 , RIdf0cb20_1521, \16325 );
nor \g455045/U$1 ( \39459 , \39457 , \39458 );
not \g450180/U$3 ( \39460 , \39459 );
not \g450180/U$4 ( \39461 , \16330 );
and \g450180/U$2 ( \39462 , \39460 , \39461 );
and \g450180/U$5 ( \39463 , \16341 , RIdef3620_1233);
nor \g450180/U$1 ( \39464 , \39462 , \39463 );
and \g452836/U$2 ( \39465 , \16377 , RIdf0f820_1553);
and \g452836/U$3 ( \39466 , RIdf12520_1585, \16313 );
nor \g452836/U$1 ( \39467 , \39465 , \39466 );
and \g452837/U$2 ( \39468 , \16334 , RIdf04420_1425);
and \g452837/U$3 ( \39469 , RIdf07120_1457, \16380 );
nor \g452837/U$1 ( \39470 , \39468 , \39469 );
nand \g447385/U$1 ( \39471 , \39456 , \39464 , \39467 , \39470 );
nor \g446219/U$1 ( \39472 , \39451 , \39452 , \39471 );
and \g452835/U$2 ( \39473 , \16361 , RIdeeaf20_1137);
and \g452835/U$3 ( \39474 , RIdefea20_1361, \16448 );
nor \g452835/U$1 ( \39475 , \39473 , \39474 );
nand \g445635/U$1 ( \39476 , \39450 , \39472 , \39475 );
and \g444787/U$2 ( \39477 , \39476 , \16750 );
and \g449162/U$2 ( \39478 , RIfc75c20_6362, \16427 );
and \g449162/U$3 ( \39479 , \16448 , RIfcc0d10_7216);
and \g449162/U$4 ( \39480 , RIdf28e88_1842, \16485 );
nor \g449162/U$1 ( \39481 , \39478 , \39479 , \39480 );
and \g455041/U$2 ( \39482 , \16317 , RIdf20620_1745);
and \g455041/U$3 ( \39483 , RIfcc9410_7312, \16325 );
nor \g455041/U$1 ( \39484 , \39482 , \39483 );
not \g455040/U$1 ( \39485 , \39484 );
and \g450178/U$2 ( \39486 , \39485 , \16336 );
and \g450178/U$3 ( \39487 , RIdf2ad78_1864, \16356 );
nor \g450178/U$1 ( \39488 , \39486 , \39487 );
and \g452830/U$2 ( \39489 , \16361 , RIdf1a0e0_1673);
and \g452830/U$3 ( \39490 , RIfc73628_6335, \16364 );
nor \g452830/U$1 ( \39491 , \39489 , \39490 );
and \g452829/U$2 ( \39492 , \16368 , RIfc74e10_6352);
and \g452829/U$3 ( \39493 , RIfca50b0_6900, \16371 );
nor \g452829/U$1 ( \39494 , \39492 , \39493 );
nand \g448090/U$1 ( \39495 , \39481 , \39488 , \39491 , \39494 );
and \g444787/U$3 ( \39496 , \16481 , \39495 );
nor \g444787/U$1 ( \39497 , \39477 , \39496 );
and \g446994/U$2 ( \39498 , \16505 , RIee2ac10_4945);
and \g446994/U$3 ( \39499 , RIee2c6c8_4964, \16507 );
nor \g446994/U$1 ( \39500 , \39498 , \39499 );
and \g446996/U$2 ( \39501 , \16511 , RIfea3770_8204);
and \g446996/U$3 ( \39502 , RIfea3608_8203, \16514 );
nor \g446996/U$1 ( \39503 , \39501 , \39502 );
and \g446995/U$2 ( \39504 , \16518 , RIee28348_4916);
and \g446995/U$3 ( \39505 , RIee29590_4929, \16521 );
nor \g446995/U$1 ( \39506 , \39504 , \39505 );
nand \g444513/U$1 ( \39507 , \39497 , \39500 , \39503 , \39506 );
and \g446215/U$2 ( \39508 , RIfea3ba8_8207, \16448 );
and \g446215/U$3 ( \39509 , RIe147450_2188, \16361 );
and \g449159/U$2 ( \39510 , RIe163650_2508, \16321 );
and \g449159/U$3 ( \39511 , \16328 , RIe166350_2540);
and \g449159/U$4 ( \39512 , RIe14ce50_2252, \16337 );
nor \g449159/U$1 ( \39513 , \39510 , \39511 , \39512 );
and \g455033/U$2 ( \39514 , \16317 , RIe15dc50_2444);
and \g455033/U$3 ( \39515 , RIfcaa678_6961, \16325 );
nor \g455033/U$1 ( \39516 , \39514 , \39515 );
not \g450174/U$3 ( \39517 , \39516 );
not \g450174/U$4 ( \39518 , \16330 );
and \g450174/U$2 ( \39519 , \39517 , \39518 );
and \g450174/U$5 ( \39520 , \16341 , RIfc62f30_6148);
nor \g450174/U$1 ( \39521 , \39519 , \39520 );
and \g452814/U$2 ( \39522 , \16377 , RIe160950_2476);
and \g452814/U$3 ( \39523 , RIee37d98_5094, \16313 );
nor \g452814/U$1 ( \39524 , \39522 , \39523 );
and \g452815/U$2 ( \39525 , \16334 , RIe155550_2348);
and \g452815/U$3 ( \39526 , RIe158250_2380, \16380 );
nor \g452815/U$1 ( \39527 , \39525 , \39526 );
nand \g447382/U$1 ( \39528 , \39513 , \39521 , \39524 , \39527 );
nor \g446215/U$1 ( \39529 , \39508 , \39509 , \39528 );
and \g452813/U$2 ( \39530 , \16364 , RIe14a150_2220);
and \g452813/U$3 ( \39531 , RIe152850_2316, \16427 );
nor \g452813/U$1 ( \39532 , \39530 , \39531 );
and \g445505/U$2 ( \39533 , \39529 , \39532 );
nor \g445505/U$1 ( \39534 , \39533 , \16389 );
and \g446218/U$2 ( \39535 , RIfcb6b58_7101, \16448 );
and \g446218/U$3 ( \39536 , RIfc9dd60_6818, \16371 );
and \g449160/U$2 ( \39537 , RIfcda648_7507, \16321 );
and \g449160/U$3 ( \39538 , \16328 , RIee1d4e8_4792);
and \g449160/U$4 ( \39539 , RIe16c458_2609, \16398 );
nor \g449160/U$1 ( \39540 , \39537 , \39538 , \39539 );
and \g455292/U$2 ( \39541 , \16317 , RIfea34a0_8202);
and \g455292/U$3 ( \39542 , RIde92ac8_305, \16325 );
nor \g455292/U$1 ( \39543 , \39541 , \39542 );
not \g450175/U$3 ( \39544 , \39543 );
not \g450175/U$4 ( \39545 , \16330 );
and \g450175/U$2 ( \39546 , \39544 , \39545 );
and \g450175/U$5 ( \39547 , \16341 , RIfc50c18_5941);
nor \g450175/U$1 ( \39548 , \39546 , \39547 );
and \g452823/U$2 ( \39549 , \16377 , RIfcd5620_7450);
and \g452823/U$3 ( \39550 , RIfcc6440_7278, \16313 );
nor \g452823/U$1 ( \39551 , \39549 , \39550 );
and \g452824/U$2 ( \39552 , \16334 , RIfea3338_8201);
and \g452824/U$3 ( \39553 , RIfea31d0_8200, \16380 );
nor \g452824/U$1 ( \39554 , \39552 , \39553 );
nand \g447383/U$1 ( \39555 , \39540 , \39548 , \39551 , \39554 );
nor \g446218/U$1 ( \39556 , \39535 , \39536 , \39555 );
and \g452819/U$2 ( \39557 , \16364 , RIfc80a80_6486);
and \g452819/U$3 ( \39558 , RIee19708_4748, \16368 );
nor \g452819/U$1 ( \39559 , \39557 , \39558 );
and \g452820/U$2 ( \39560 , \16361 , RIfec62e8_8375);
and \g452820/U$3 ( \39561 , RIfcb6888_7099, \16427 );
nor \g452820/U$1 ( \39562 , \39560 , \39561 );
and \g445303/U$2 ( \39563 , \39556 , \39559 , \39562 );
nor \g445303/U$1 ( \39564 , \39563 , \16649 );
nor \g444413/U$1 ( \39565 , \39447 , \39507 , \39534 , \39564 );
and \g452804/U$2 ( \39566 , \16364 , RIdedcf88_978);
and \g452804/U$3 ( \39567 , RIdf2d7a8_1894, \16371 );
nor \g452804/U$1 ( \39568 , \39566 , \39567 );
and \g446214/U$2 ( \39569 , RIdf39148_2026, \16427 );
and \g446214/U$3 ( \39570 , RIdf1e028_1718, \16368 );
and \g449155/U$2 ( \39571 , RIdecea50_815, \16321 );
and \g449155/U$3 ( \39572 , \16328 , RIded1750_847);
and \g449155/U$4 ( \39573 , RIdee8220_1105, \16398 );
nor \g449155/U$1 ( \39574 , \39571 , \39572 , \39573 );
and \g455273/U$2 ( \39575 , \16317 , RIde98d38_335);
and \g455273/U$3 ( \39576 , RIdeb5550_527, \16325 );
nor \g455273/U$1 ( \39577 , \39575 , \39576 );
not \g450171/U$3 ( \39578 , \39577 );
not \g450171/U$4 ( \39579 , \16330 );
and \g450171/U$2 ( \39580 , \39578 , \39579 );
and \g450171/U$5 ( \39581 , \16341 , RIdf01720_1393);
nor \g450171/U$1 ( \39582 , \39580 , \39581 );
and \g452807/U$2 ( \39583 , \16377 , RIdec9050_751);
and \g452807/U$3 ( \39584 , RIdecbd50_783, \16313 );
nor \g452807/U$1 ( \39585 , \39583 , \39584 );
and \g452808/U$2 ( \39586 , \16334 , RIe15af50_2412);
and \g452808/U$3 ( \39587 , RIe16f158_2641, \16380 );
nor \g452808/U$1 ( \39588 , \39586 , \39587 );
nand \g447381/U$1 ( \39589 , \39574 , \39582 , \39585 , \39588 );
nor \g446214/U$1 ( \39590 , \39569 , \39570 , \39589 );
and \g452805/U$2 ( \39591 , \16361 , RIde7ec80_208);
and \g452805/U$3 ( \39592 , RIe144750_2156, \16432 );
nor \g452805/U$1 ( \39593 , \39591 , \39592 );
nand \g445631/U$1 ( \39594 , \39568 , \39590 , \39593 );
and \g444673/U$2 ( \39595 , \39594 , \16752 );
and \g452798/U$2 ( \39596 , \16377 , RIfc58ee0_6034);
and \g452798/U$3 ( \39597 , RIdee15d8_1028, \16380 );
nor \g452798/U$1 ( \39598 , \39596 , \39597 );
and \g446213/U$2 ( \39599 , RIfc7c598_6437, \16321 );
and \g446213/U$3 ( \39600 , RIfc5beb0_6068, \16313 );
and \g449154/U$2 ( \39601 , RIded7f60_921, \16398 );
and \g449154/U$3 ( \39602 , \16339 , RIdeda558_948);
and \g449154/U$4 ( \39603 , RIdee3798_1052, \16344 );
nor \g449154/U$1 ( \39604 , \39601 , \39602 , \39603 );
and \g455023/U$2 ( \39605 , \16317 , RIfc72ae8_6327);
and \g455023/U$3 ( \39606 , RIfcb3048_7059, \16325 );
nor \g455023/U$1 ( \39607 , \39605 , \39606 );
not \g450169/U$3 ( \39608 , \39607 );
not \g450169/U$4 ( \39609 , \16351 );
and \g450169/U$2 ( \39610 , \39608 , \39609 );
and \g450169/U$5 ( \39611 , \16356 , RIdee5688_1074);
nor \g450169/U$1 ( \39612 , \39610 , \39611 );
and \g452801/U$2 ( \39613 , \16361 , RIded3a78_872);
and \g452801/U$3 ( \39614 , RIfea3068_8199, \16364 );
nor \g452801/U$1 ( \39615 , \39613 , \39614 );
and \g452799/U$2 ( \39616 , \16368 , RIfcb6450_7096);
and \g452799/U$3 ( \39617 , RIfca3d00_6886, \16371 );
nor \g452799/U$1 ( \39618 , \39616 , \39617 );
nand \g447805/U$1 ( \39619 , \39604 , \39612 , \39615 , \39618 );
nor \g446213/U$1 ( \39620 , \39599 , \39600 , \39619 );
and \g452797/U$2 ( \39621 , \16334 , RIdedf580_1005);
and \g452797/U$3 ( \39622 , RIfcab8c0_6974, \16328 );
nor \g452797/U$1 ( \39623 , \39621 , \39622 );
nand \g445630/U$1 ( \39624 , \39598 , \39620 , \39623 );
and \g444673/U$3 ( \39625 , \16477 , \39624 );
nor \g444673/U$1 ( \39626 , \39595 , \39625 );
nand \g444286/U$1 ( \39627 , \39443 , \39565 , \39626 );
_DC \g64f1/U$1 ( \39628 , \39627 , \16652 );
and \g449198/U$2 ( \39629 , RIe20b440_4418, \8317 );
and \g449198/U$3 ( \39630 , \8326 , RIe20e140_4450);
and \g449198/U$4 ( \39631 , RIe21ef40_4642, \8409 );
nor \g449198/U$1 ( \39632 , \39629 , \39630 , \39631 );
and \g452958/U$2 ( \39633 , \8335 , RIe208740_4386);
and \g452958/U$3 ( \39634 , RIfcab1b8_6969, \8340 );
nor \g452958/U$1 ( \39635 , \39633 , \39634 );
and \g452957/U$2 ( \39636 , \8404 , RIe221c40_4674);
and \g452957/U$3 ( \39637 , RIfc44cd8_5805, \8351 );
nor \g452957/U$1 ( \39638 , \39636 , \39637 );
and \g454943/U$2 ( \39639 , \8313 , RIfcb6180_7094);
and \g454943/U$3 ( \39640 , RIe224940_4706, \8323 );
nor \g454943/U$1 ( \39641 , \39639 , \39640 );
not \g450214/U$3 ( \39642 , \39641 );
not \g450214/U$4 ( \39643 , \8328 );
and \g450214/U$2 ( \39644 , \39642 , \39643 );
and \g450214/U$5 ( \39645 , \8417 , RIfc55ad8_5997);
nor \g450214/U$1 ( \39646 , \39644 , \39645 );
nand \g447826/U$1 ( \39647 , \39632 , \39635 , \39638 , \39646 );
and \g444790/U$2 ( \39648 , \39647 , \8369 );
and \g446248/U$2 ( \39649 , RIe203178_4325, \8373 );
and \g446248/U$3 ( \39650 , RIfc64178_6161, \8330 );
and \g449199/U$2 ( \39651 , RIfc4f160_5922, \8324 );
and \g449199/U$3 ( \39652 , \8531 , RIfea2ac8_8195);
and \g449199/U$4 ( \39653 , RIfca8bc0_6942, \8488 );
nor \g449199/U$1 ( \39654 , \39651 , \39652 , \39653 );
and \g452965/U$2 ( \39655 , \8356 , RIfea2c30_8196);
and \g452965/U$3 ( \39656 , RIfcc9c80_7318, \8359 );
nor \g452965/U$1 ( \39657 , \39655 , \39656 );
and \g454929/U$2 ( \39658 , \8313 , RIfc7f838_6473);
and \g454929/U$3 ( \39659 , RIf164828_5603, \8323 );
nor \g454929/U$1 ( \39660 , \39658 , \39659 );
not \g450215/U$3 ( \39661 , \39660 );
not \g450215/U$4 ( \39662 , \8376 );
and \g450215/U$2 ( \39663 , \39661 , \39662 );
and \g450215/U$5 ( \39664 , \8340 , RIfc59318_6037);
nor \g450215/U$1 ( \39665 , \39663 , \39664 );
and \g452964/U$2 ( \39666 , \8378 , RIf162398_5577);
and \g452964/U$3 ( \39667 , RIfcd2ec0_7422, \8417 );
nor \g452964/U$1 ( \39668 , \39666 , \39667 );
nand \g447828/U$1 ( \39669 , \39654 , \39657 , \39665 , \39668 );
nor \g446248/U$1 ( \39670 , \39649 , \39650 , \39669 );
and \g452960/U$2 ( \39671 , \8335 , RIfcebf88_7707);
and \g452960/U$3 ( \39672 , RIfce3720_7610, \8351 );
nor \g452960/U$1 ( \39673 , \39671 , \39672 );
and \g452961/U$2 ( \39674 , \8319 , RIf15ac10_5492);
and \g452961/U$3 ( \39675 , RIe201558_4305, \8404 );
nor \g452961/U$1 ( \39676 , \39674 , \39675 );
and \g445327/U$2 ( \39677 , \39670 , \39673 , \39676 );
nor \g445327/U$1 ( \39678 , \39677 , \8422 );
nor \g444790/U$1 ( \39679 , \39648 , \39678 );
and \g447017/U$2 ( \39680 , \8438 , RIe216840_4546);
and \g447017/U$3 ( \39681 , RIe219540_4578, \8440 );
nor \g447017/U$1 ( \39682 , \39680 , \39681 );
and \g447016/U$2 ( \39683 , \12506 , RIe213b40_4514);
and \g447016/U$3 ( \39684 , RIfc4dc48_5907, \12508 );
nor \g447016/U$1 ( \39685 , \39683 , \39684 );
and \g447018/U$2 ( \39686 , \8717 , RIe210e40_4482);
and \g447018/U$3 ( \39687 , RIfcdcf10_7536, \8719 );
nor \g447018/U$1 ( \39688 , \39686 , \39687 );
nand \g444518/U$1 ( \39689 , \39679 , \39682 , \39685 , \39688 );
and \g447013/U$2 ( \39690 , \9170 , RIe1904e8_3019);
and \g447013/U$3 ( \39691 , RIe1931e8_3051, \9172 );
nor \g447013/U$1 ( \39692 , \39690 , \39691 );
and \g446244/U$2 ( \39693 , RIe187de8_2923, \8486 );
and \g446244/U$3 ( \39694 , RIe18aae8_2955, \8359 );
and \g449194/U$2 ( \39695 , RIe195ee8_3083, \8409 );
and \g449194/U$3 ( \39696 , \8373 , RIfca84b8_6937);
and \g449194/U$4 ( \39697 , RIe19b8e8_3147, \8383 );
nor \g449194/U$1 ( \39698 , \39695 , \39696 , \39697 );
and \g452945/U$2 ( \39699 , \8335 , RIe17c9e8_2795);
and \g452945/U$3 ( \39700 , RIfc8e310_6640, \8340 );
nor \g452945/U$1 ( \39701 , \39699 , \39700 );
and \g452944/U$2 ( \39702 , \8404 , RIe198be8_3115);
and \g452944/U$3 ( \39703 , RIe19e5e8_3179, \8351 );
nor \g452944/U$1 ( \39704 , \39702 , \39703 );
and \g455369/U$2 ( \39705 , \8313 , RIe17f6e8_2827);
and \g455369/U$3 ( \39706 , RIe1823e8_2859, \8323 );
nor \g455369/U$1 ( \39707 , \39705 , \39706 );
not \g455368/U$1 ( \39708 , \39707 );
and \g450211/U$2 ( \39709 , \39708 , \8316 );
and \g450211/U$3 ( \39710 , RIfc846f8_6529, \8417 );
nor \g450211/U$1 ( \39711 , \39709 , \39710 );
nand \g448208/U$1 ( \39712 , \39698 , \39701 , \39704 , \39711 );
nor \g446244/U$1 ( \39713 , \39693 , \39694 , \39712 );
not \g444818/U$3 ( \39714 , \39713 );
not \g444818/U$4 ( \39715 , \8589 );
and \g444818/U$2 ( \39716 , \39714 , \39715 );
and \g446245/U$2 ( \39717 , RIf1404c8_5191, \8373 );
and \g446245/U$3 ( \39718 , RIfccc278_7345, \8383 );
and \g449196/U$2 ( \39719 , RIee3e5a8_5168, \8414 );
and \g449196/U$3 ( \39720 , \8409 , RIfc60398_6117);
and \g449196/U$4 ( \39721 , RIfc5c720_6074, \8326 );
nor \g449196/U$1 ( \39722 , \39719 , \39720 , \39721 );
and \g452953/U$2 ( \39723 , \8356 , RIfec6180_8374);
and \g452953/U$3 ( \39724 , RIfc642e0_6162, \8359 );
nor \g452953/U$1 ( \39725 , \39723 , \39724 );
and \g455123/U$2 ( \39726 , \8313 , RIee3a228_5120);
and \g455123/U$3 ( \39727 , RIfca7f18_6933, \8323 );
nor \g455123/U$1 ( \39728 , \39726 , \39727 );
not \g450212/U$3 ( \39729 , \39728 );
not \g450212/U$4 ( \39730 , \8347 );
and \g450212/U$2 ( \39731 , \39729 , \39730 );
and \g450212/U$5 ( \39732 , \8340 , RIfca9598_6949);
nor \g450212/U$1 ( \39733 , \39731 , \39732 );
and \g452952/U$2 ( \39734 , \8378 , RIee3da68_5160);
and \g452952/U$3 ( \39735 , RIfcc1b20_7226, \8417 );
nor \g452952/U$1 ( \39736 , \39734 , \39735 );
nand \g447825/U$1 ( \39737 , \39722 , \39725 , \39733 , \39736 );
nor \g446245/U$1 ( \39738 , \39717 , \39718 , \39737 );
and \g452948/U$2 ( \39739 , \8335 , RIfccaec8_7331);
and \g452948/U$3 ( \39740 , RIfcd1570_7404, \8351 );
nor \g452948/U$1 ( \39741 , \39739 , \39740 );
and \g452950/U$2 ( \39742 , \8319 , RIfc6bea0_6250);
and \g452950/U$3 ( \39743 , RIfea2d98_8197, \8404 );
nor \g452950/U$1 ( \39744 , \39742 , \39743 );
and \g445323/U$2 ( \39745 , \39738 , \39741 , \39744 );
nor \g445323/U$1 ( \39746 , \39745 , \8558 );
nor \g444818/U$1 ( \39747 , \39716 , \39746 );
and \g447012/U$2 ( \39748 , \9230 , RIe1850e8_2891);
and \g447012/U$3 ( \39749 , RIfce2be0_7602, \9232 );
nor \g447012/U$1 ( \39750 , \39748 , \39749 );
nand \g444429/U$1 ( \39751 , \39692 , \39747 , \39750 );
and \g446240/U$2 ( \39752 , RIfc45c50_5816, \8414 );
and \g446240/U$3 ( \39753 , RIfec6018_8373, \8356 );
and \g449189/U$2 ( \39754 , RIfc4c028_5887, \8319 );
and \g449189/U$3 ( \39755 , \8326 , RIfc434f0_5788);
and \g449189/U$4 ( \39756 , RIf155a80_5434, \8407 );
nor \g449189/U$1 ( \39757 , \39754 , \39755 , \39756 );
and \g452933/U$2 ( \39758 , \8335 , RIe1eee08_4095);
and \g452933/U$3 ( \39759 , RIfc64010_6160, \8340 );
nor \g452933/U$1 ( \39760 , \39758 , \39759 );
and \g452932/U$2 ( \39761 , \8404 , RIe1faeb0_4232);
and \g452932/U$3 ( \39762 , RIfcbb040_7150, \8351 );
nor \g452932/U$1 ( \39763 , \39761 , \39762 );
and \g454984/U$2 ( \39764 , \8313 , RIfc93d10_6704);
and \g454984/U$3 ( \39765 , RIfca1870_6860, \8323 );
nor \g454984/U$1 ( \39766 , \39764 , \39765 );
not \g450206/U$3 ( \39767 , \39766 );
not \g450206/U$4 ( \39768 , \8328 );
and \g450206/U$2 ( \39769 , \39767 , \39768 );
and \g450206/U$5 ( \39770 , \8417 , RIf1565c0_5442);
nor \g450206/U$1 ( \39771 , \39769 , \39770 );
nand \g447822/U$1 ( \39772 , \39757 , \39760 , \39763 , \39771 );
nor \g446240/U$1 ( \39773 , \39752 , \39753 , \39772 );
and \g452931/U$2 ( \39774 , \8378 , RIe1f6428_4179);
and \g452931/U$3 ( \39775 , RIfccdbc8_7363, \8359 );
nor \g452931/U$1 ( \39776 , \39774 , \39775 );
and \g452930/U$2 ( \39777 , \8531 , RIfca6cd0_6920);
and \g452930/U$3 ( \39778 , RIfcccae8_7351, \8488 );
nor \g452930/U$1 ( \39779 , \39777 , \39778 );
and \g445319/U$2 ( \39780 , \39773 , \39776 , \39779 );
nor \g445319/U$1 ( \39781 , \39780 , \8621 );
and \g446242/U$2 ( \39782 , RIe1db8a8_3875, \8414 );
and \g446242/U$3 ( \39783 , RIe1cd7a8_3715, \8531 );
and \g449191/U$2 ( \39784 , RIe1c23a8_3587, \8317 );
and \g449191/U$3 ( \39785 , \8326 , RIe1c50a8_3619);
and \g449191/U$4 ( \39786 , RIe1de5a8_3907, \8409 );
nor \g449191/U$1 ( \39787 , \39784 , \39785 , \39786 );
and \g452941/U$2 ( \39788 , \8335 , RIe1bf6a8_3555);
and \g452941/U$3 ( \39789 , RIe1c7da8_3651, \8340 );
nor \g452941/U$1 ( \39790 , \39788 , \39789 );
and \g452940/U$2 ( \39791 , \8404 , RIe1e3fa8_3971);
and \g452940/U$3 ( \39792 , RIe1ec6a8_4067, \8351 );
nor \g452940/U$1 ( \39793 , \39791 , \39792 );
and \g455113/U$2 ( \39794 , \8313 , RIe1e6ca8_4003);
and \g455113/U$3 ( \39795 , RIe1e99a8_4035, \8323 );
nor \g455113/U$1 ( \39796 , \39794 , \39795 );
not \g450209/U$3 ( \39797 , \39796 );
not \g450209/U$4 ( \39798 , \8328 );
and \g450209/U$2 ( \39799 , \39797 , \39798 );
and \g450209/U$5 ( \39800 , \8417 , RIe1e12a8_3939);
nor \g450209/U$1 ( \39801 , \39799 , \39800 );
nand \g447823/U$1 ( \39802 , \39787 , \39790 , \39793 , \39801 );
nor \g446242/U$1 ( \39803 , \39782 , \39783 , \39802 );
and \g452936/U$2 ( \39804 , \8356 , RIe1caaa8_3683);
and \g452936/U$3 ( \39805 , RIe1d31a8_3779, \8359 );
nor \g452936/U$1 ( \39806 , \39804 , \39805 );
and \g452938/U$2 ( \39807 , \8378 , RIe1d8ba8_3843);
and \g452938/U$3 ( \39808 , RIe1d04a8_3747, \8488 );
nor \g452938/U$1 ( \39809 , \39807 , \39808 );
and \g445321/U$2 ( \39810 , \39803 , \39806 , \39809 );
nor \g445321/U$1 ( \39811 , \39810 , \8477 );
or \g444306/U$1 ( \39812 , \39689 , \39751 , \39781 , \39811 );
and \g446237/U$2 ( \39813 , RIfea2f00_8198, \8378 );
and \g446237/U$3 ( \39814 , RIfc9bfd8_6797, \8359 );
and \g449186/U$2 ( \39815 , RIfc92ac8_6691, \8407 );
and \g449186/U$3 ( \39816 , \8373 , RIe1ba0e0_3494);
and \g449186/U$4 ( \39817 , RIfc6bd38_6249, \8330 );
nor \g449186/U$1 ( \39818 , \39815 , \39816 , \39817 );
and \g452917/U$2 ( \39819 , \8335 , RIe1ab8d8_3329);
and \g452917/U$3 ( \39820 , RIfc4df18_5909, \8340 );
nor \g452917/U$1 ( \39821 , \39819 , \39820 );
and \g452916/U$2 ( \39822 , \8404 , RIe1b7f20_3470);
and \g452916/U$3 ( \39823 , RIfc63908_6155, \8351 );
nor \g452916/U$1 ( \39824 , \39822 , \39823 );
and \g455013/U$2 ( \39825 , \8313 , RIe1ad0c0_3346);
and \g455013/U$3 ( \39826 , RIfc9d658_6813, \8323 );
nor \g455013/U$1 ( \39827 , \39825 , \39826 );
not \g455012/U$1 ( \39828 , \39827 );
and \g450202/U$2 ( \39829 , \39828 , \8316 );
and \g450202/U$3 ( \39830 , RIfc66fe0_6194, \8417 );
nor \g450202/U$1 ( \39831 , \39829 , \39830 );
nand \g448207/U$1 ( \39832 , \39818 , \39821 , \39824 , \39831 );
nor \g446237/U$1 ( \39833 , \39813 , \39814 , \39832 );
and \g452913/U$2 ( \39834 , \8356 , RIe1b1878_3397);
and \g452913/U$3 ( \39835 , RIe1b5d60_3446, \8412 );
nor \g452913/U$1 ( \39836 , \39834 , \39835 );
and \g452912/U$2 ( \39837 , \8531 , RIe1b31c8_3415);
and \g452912/U$3 ( \39838 , RIfc50d80_5942, \8488 );
nor \g452912/U$1 ( \39839 , \39837 , \39838 );
and \g445317/U$2 ( \39840 , \39833 , \39836 , \39839 );
nor \g445317/U$1 ( \39841 , \39840 , \8481 );
and \g446238/U$2 ( \39842 , RIe1a3fe8_3243, \8371 );
and \g446238/U$3 ( \39843 , RIe1a6ce8_3275, \8330 );
and \g449187/U$2 ( \39844 , RIe227640_4738, \8414 );
and \g449187/U$3 ( \39845 , \8409 , RIe179ce8_2763);
and \g449187/U$4 ( \39846 , RIe1bc9a8_3523, \8324 );
nor \g449187/U$1 ( \39847 , \39844 , \39845 , \39846 );
and \g452924/U$2 ( \39848 , \8356 , RIe1f19a0_4126);
and \g452924/U$3 ( \39849 , RIe205a40_4354, \8359 );
nor \g452924/U$1 ( \39850 , \39848 , \39849 );
and \g455109/U$2 ( \39851 , \8313 , RIe1f8e58_4209);
and \g455109/U$3 ( \39852 , RIe1ffaa0_4286, \8323 );
nor \g455109/U$1 ( \39853 , \39851 , \39852 );
not \g450203/U$3 ( \39854 , \39853 );
not \g450203/U$4 ( \39855 , \8347 );
and \g450203/U$2 ( \39856 , \39854 , \39855 );
and \g450203/U$5 ( \39857 , \8340 , RIe1d5ea8_3811);
nor \g450203/U$1 ( \39858 , \39856 , \39857 );
and \g452922/U$2 ( \39859 , \8378 , RIe21c240_4610);
and \g452922/U$3 ( \39860 , RIe18d7e8_2987, \8417 );
nor \g452922/U$1 ( \39861 , \39859 , \39860 );
nand \g447819/U$1 ( \39862 , \39847 , \39850 , \39858 , \39861 );
nor \g446238/U$1 ( \39863 , \39842 , \39843 , \39862 );
and \g452918/U$2 ( \39864 , \8335 , RIe171e58_2673);
and \g452918/U$3 ( \39865 , RIe1a99e8_3307, \8351 );
nor \g452918/U$1 ( \39866 , \39864 , \39865 );
and \g452920/U$2 ( \39867 , \8319 , RIe1af820_3374);
and \g452920/U$3 ( \39868 , RIe1a12e8_3211, \8404 );
nor \g452920/U$1 ( \39869 , \39867 , \39868 );
and \g445318/U$2 ( \39870 , \39863 , \39866 , \39869 );
nor \g445318/U$1 ( \39871 , \39870 , \8651 );
or \g444164/U$1 ( \39872 , \39812 , \39841 , \39871 );
_DC \g6575/U$1 ( \39873 , \39872 , \8654 );
_DC \g6577/U$1 ( \39874 , \24539 , \16652 );
_DC \g6578/U$1 ( \39875 , \24783 , \8654 );
_DC \g657a/U$1 ( \39876 , \25025 , \16652 );
_DC \g657b/U$1 ( \39877 , \25270 , \8654 );
_DC \g657d/U$1 ( \39878 , \25513 , \16652 );
_DC \g657e/U$1 ( \39879 , \25758 , \8654 );
_DC \g6580/U$1 ( \39880 , \26001 , \16652 );
_DC \g6581/U$1 ( \39881 , \26243 , \8654 );
_DC \g6583/U$1 ( \39882 , \26489 , \16652 );
_DC \g6584/U$1 ( \39883 , \26735 , \8654 );
_DC \g6586/U$1 ( \39884 , \26978 , \16652 );
_DC \g6587/U$1 ( \39885 , \27219 , \8654 );
_DC \g6589/U$1 ( \39886 , \27463 , \16652 );
_DC \g658a/U$1 ( \39887 , \27706 , \8654 );
_DC \g658c/U$1 ( \39888 , \27951 , \16652 );
_DC \g658d/U$1 ( \39889 , \28196 , \8654 );
_DC \g658f/U$1 ( \39890 , \28438 , \16652 );
_DC \g6590/U$1 ( \39891 , \28681 , \8654 );
_DC \g6592/U$1 ( \39892 , \28924 , \16652 );
_DC \g6593/U$1 ( \39893 , \29169 , \8654 );
_DC \g6595/U$1 ( \39894 , \29410 , \16652 );
_DC \g6596/U$1 ( \39895 , \29652 , \8654 );
_DC \g6598/U$1 ( \39896 , \29893 , \16652 );
_DC \g6599/U$1 ( \39897 , \30136 , \8654 );
_DC \g659b/U$1 ( \39898 , \30381 , \16652 );
_DC \g659c/U$1 ( \39899 , \30624 , \8654 );
_DC \g659e/U$1 ( \39900 , \30866 , \16652 );
_DC \g659f/U$1 ( \39901 , \31107 , \8654 );
_DC \g65a1/U$1 ( \39902 , \31350 , \16652 );
_DC \g65a2/U$1 ( \39903 , \31594 , \8654 );
_DC \g65a4/U$1 ( \39904 , \31834 , \16652 );
_DC \g65a5/U$1 ( \39905 , \32078 , \8654 );
_DC \g65a7/U$1 ( \39906 , \32320 , \16652 );
_DC \g65a8/U$1 ( \39907 , \32565 , \8654 );
_DC \g65aa/U$1 ( \39908 , \32810 , \16652 );
_DC \g65ab/U$1 ( \39909 , \33056 , \8654 );
_DC \g65ad/U$1 ( \39910 , \33301 , \16652 );
_DC \g65ae/U$1 ( \39911 , \33544 , \8654 );
_DC \g65b0/U$1 ( \39912 , \33785 , \16652 );
_DC \g65b1/U$1 ( \39913 , \34026 , \8654 );
_DC \g65b3/U$1 ( \39914 , \34269 , \16652 );
_DC \g65b4/U$1 ( \39915 , \34512 , \8654 );
_DC \g65b6/U$1 ( \39916 , \34755 , \16652 );
_DC \g65b7/U$1 ( \39917 , \35002 , \8654 );
_DC \g65b9/U$1 ( \39918 , \35244 , \16652 );
_DC \g65ba/U$1 ( \39919 , \35488 , \8654 );
_DC \g65bc/U$1 ( \39920 , \35731 , \16652 );
_DC \g65bd/U$1 ( \39921 , \35973 , \8654 );
_DC \g65bf/U$1 ( \39922 , \36216 , \16652 );
_DC \g65c0/U$1 ( \39923 , \36458 , \8654 );
_DC \g65c2/U$1 ( \39924 , \36702 , \16652 );
_DC \g65c3/U$1 ( \39925 , \36947 , \8654 );
_DC \g65c5/U$1 ( \39926 , \37190 , \16652 );
_DC \g65c6/U$1 ( \39927 , \37436 , \8654 );
_DC \g65c8/U$1 ( \39928 , \37680 , \16652 );
_DC \g65c9/U$1 ( \39929 , \37923 , \8654 );
_DC \g65cb/U$1 ( \39930 , \38167 , \16652 );
_DC \g65cc/U$1 ( \39931 , \38413 , \8654 );
_DC \g65ce/U$1 ( \39932 , \38655 , \16652 );
_DC \g65cf/U$1 ( \39933 , \38896 , \8654 );
_DC \g65d1/U$1 ( \39934 , \39139 , \16652 );
_DC \g65d2/U$1 ( \39935 , \39382 , \8654 );
_DC \g65d4/U$1 ( \39936 , \39627 , \16652 );
_DC \g65d5/U$1 ( \39937 , \39872 , \8654 );
xor \g132399/U$1 ( \39938 , \16653 , \8655 );
xor \g132463/U$4 ( \39939 , \16912 , \8913 );
xor \g132520/U$4 ( \39940 , \17162 , \9169 );
xor \g132578/U$4 ( \39941 , \17412 , \9425 );
xor \g132633/U$4 ( \39942 , \17661 , \9670 );
xor \g132693/U$4 ( \39943 , \17908 , \9922 );
xor \g132737/U$4 ( \39944 , \18157 , \10170 );
xor \g132792/U$4 ( \39945 , \18405 , \10422 );
xor \g132835/U$4 ( \39946 , \18659 , \10670 );
xor \g132885/U$4 ( \39947 , \18910 , \10912 );
xor \g132923/U$4 ( \39948 , \19156 , \11157 );
xor \g132971/U$4 ( \39949 , \19406 , \11400 );
xor \g133005/U$4 ( \39950 , \19652 , \11649 );
xor \g133048/U$4 ( \39951 , \19894 , \11898 );
xor \g133086/U$4 ( \39952 , \20139 , \12140 );
xor \g133124/U$4 ( \39953 , \20384 , \12391 );
xor \g133152/U$4 ( \39954 , \20628 , \12636 );
xor \g133202/U$4 ( \39955 , \20875 , \12879 );
xor \g133252/U$4 ( \39956 , \21118 , \13123 );
xor \g133295/U$4 ( \39957 , \21361 , \13370 );
xor \g133353/U$4 ( \39958 , \21605 , \13617 );
xor \g133405/U$4 ( \39959 , \21847 , \13864 );
xor \g133476/U$4 ( \39960 , \22092 , \14107 );
xor \g133539/U$4 ( \39961 , \22336 , \14354 );
xor \g133630/U$4 ( \39962 , \22585 , \14597 );
xor \g133728/U$4 ( \39963 , \22831 , \14840 );
xor \g133847/U$4 ( \39964 , \23076 , \15087 );
xor \g134037/U$4 ( \39965 , \23318 , \15330 );
xor \g134140/U$4 ( \39966 , \23562 , \15573 );
xor \g134673/U$4 ( \39967 , \15818 , \23804 );
xor \g135269/U$4 ( \39968 , \24050 , \16062 );
and \g135396/U$2 ( \39969 , \24296 , \16306 );
and \g135269/U$3 ( \39970 , \39968 , \39969 );
and \g135269/U$5 ( \39971 , \24050 , \16062 );
or \g135269/U$2 ( \39972 , \39970 , \39971 );
and \g134673/U$3 ( \39973 , \39967 , \39972 );
and \g134673/U$5 ( \39974 , \15818 , \23804 );
or \g134673/U$2 ( \39975 , \39973 , \39974 );
and \g134140/U$3 ( \39976 , \39966 , \39975 );
and \g134140/U$5 ( \39977 , \23562 , \15573 );
or \g134140/U$2 ( \39978 , \39976 , \39977 );
and \g134037/U$3 ( \39979 , \39965 , \39978 );
and \g134037/U$5 ( \39980 , \23318 , \15330 );
or \g134037/U$2 ( \39981 , \39979 , \39980 );
and \g133847/U$3 ( \39982 , \39964 , \39981 );
and \g133847/U$5 ( \39983 , \23076 , \15087 );
or \g133847/U$2 ( \39984 , \39982 , \39983 );
and \g133728/U$3 ( \39985 , \39963 , \39984 );
and \g133728/U$5 ( \39986 , \22831 , \14840 );
or \g133728/U$2 ( \39987 , \39985 , \39986 );
and \g133630/U$3 ( \39988 , \39962 , \39987 );
and \g133630/U$5 ( \39989 , \22585 , \14597 );
or \g133630/U$2 ( \39990 , \39988 , \39989 );
and \g133539/U$3 ( \39991 , \39961 , \39990 );
and \g133539/U$5 ( \39992 , \22336 , \14354 );
or \g133539/U$2 ( \39993 , \39991 , \39992 );
and \g133476/U$3 ( \39994 , \39960 , \39993 );
and \g133476/U$5 ( \39995 , \22092 , \14107 );
or \g133476/U$2 ( \39996 , \39994 , \39995 );
and \g133405/U$3 ( \39997 , \39959 , \39996 );
and \g133405/U$5 ( \39998 , \21847 , \13864 );
or \g133405/U$2 ( \39999 , \39997 , \39998 );
and \g133353/U$3 ( \40000 , \39958 , \39999 );
and \g133353/U$5 ( \40001 , \21605 , \13617 );
or \g133353/U$2 ( \40002 , \40000 , \40001 );
and \g133295/U$3 ( \40003 , \39957 , \40002 );
and \g133295/U$5 ( \40004 , \21361 , \13370 );
or \g133295/U$2 ( \40005 , \40003 , \40004 );
and \g133252/U$3 ( \40006 , \39956 , \40005 );
and \g133252/U$5 ( \40007 , \21118 , \13123 );
or \g133252/U$2 ( \40008 , \40006 , \40007 );
and \g133202/U$3 ( \40009 , \39955 , \40008 );
and \g133202/U$5 ( \40010 , \20875 , \12879 );
or \g133202/U$2 ( \40011 , \40009 , \40010 );
and \g133152/U$3 ( \40012 , \39954 , \40011 );
and \g133152/U$5 ( \40013 , \20628 , \12636 );
or \g133152/U$2 ( \40014 , \40012 , \40013 );
and \g133124/U$3 ( \40015 , \39953 , \40014 );
and \g133124/U$5 ( \40016 , \20384 , \12391 );
or \g133124/U$2 ( \40017 , \40015 , \40016 );
and \g133086/U$3 ( \40018 , \39952 , \40017 );
and \g133086/U$5 ( \40019 , \20139 , \12140 );
or \g133086/U$2 ( \40020 , \40018 , \40019 );
and \g133048/U$3 ( \40021 , \39951 , \40020 );
and \g133048/U$5 ( \40022 , \19894 , \11898 );
or \g133048/U$2 ( \40023 , \40021 , \40022 );
and \g133005/U$3 ( \40024 , \39950 , \40023 );
and \g133005/U$5 ( \40025 , \19652 , \11649 );
or \g133005/U$2 ( \40026 , \40024 , \40025 );
and \g132971/U$3 ( \40027 , \39949 , \40026 );
and \g132971/U$5 ( \40028 , \19406 , \11400 );
or \g132971/U$2 ( \40029 , \40027 , \40028 );
and \g132923/U$3 ( \40030 , \39948 , \40029 );
and \g132923/U$5 ( \40031 , \19156 , \11157 );
or \g132923/U$2 ( \40032 , \40030 , \40031 );
and \g132885/U$3 ( \40033 , \39947 , \40032 );
and \g132885/U$5 ( \40034 , \18910 , \10912 );
or \g132885/U$2 ( \40035 , \40033 , \40034 );
and \g132835/U$3 ( \40036 , \39946 , \40035 );
and \g132835/U$5 ( \40037 , \18659 , \10670 );
or \g132835/U$2 ( \40038 , \40036 , \40037 );
and \g132792/U$3 ( \40039 , \39945 , \40038 );
and \g132792/U$5 ( \40040 , \18405 , \10422 );
or \g132792/U$2 ( \40041 , \40039 , \40040 );
and \g132737/U$3 ( \40042 , \39944 , \40041 );
and \g132737/U$5 ( \40043 , \18157 , \10170 );
or \g132737/U$2 ( \40044 , \40042 , \40043 );
and \g132693/U$3 ( \40045 , \39943 , \40044 );
and \g132693/U$5 ( \40046 , \17908 , \9922 );
or \g132693/U$2 ( \40047 , \40045 , \40046 );
and \g132633/U$3 ( \40048 , \39942 , \40047 );
and \g132633/U$5 ( \40049 , \17661 , \9670 );
or \g132633/U$2 ( \40050 , \40048 , \40049 );
and \g132578/U$3 ( \40051 , \39941 , \40050 );
and \g132578/U$5 ( \40052 , \17412 , \9425 );
or \g132578/U$2 ( \40053 , \40051 , \40052 );
and \g132520/U$3 ( \40054 , \39940 , \40053 );
and \g132520/U$5 ( \40055 , \17162 , \9169 );
or \g132520/U$2 ( \40056 , \40054 , \40055 );
and \g132463/U$3 ( \40057 , \39939 , \40056 );
and \g132463/U$5 ( \40058 , \16912 , \8913 );
or \g132463/U$2 ( \40059 , \40057 , \40058 );
xnor \g132399/U$1_r1 ( \40060 , \39938 , \40059 );
not \g132398/U$1 ( \40061 , \40060 );
xnor \g135604/U$1 ( \40062 , \39628 , \39873 );
not \g135572/U$2 ( \40063 , \40062 );
and \g135476/U$1 ( \40064 , \39936 , \39937 );
nand \g135572/U$1 ( \40065 , \40063 , \40064 );
not \g135271/U$3 ( \40066 , \40065 );
and \g135455/U$1 ( \40067 , \39934 , \39935 );
not \g135578/U$2 ( \40068 , \40067 );
nor \g135578/U$1 ( \40069 , \40068 , \40062 );
not \g135271/U$4 ( \40070 , \40069 );
or \g135271/U$2 ( \40071 , \40066 , \40070 );
or \g135271/U$5 ( \40072 , \40069 , \40065 );
nand \g135271/U$1 ( \40073 , \40071 , \40072 );
xnor \g135429/U$1 ( \40074 , \38897 , \38656 );
not \g135253/U$3 ( \40075 , \40074 );
xnor \g135407/U$1 ( \40076 , \39383 , \39140 );
not \g135253/U$4 ( \40077 , \40076 );
and \g135253/U$2 ( \40078 , \40075 , \40077 );
nor \g135253/U$1 ( \40079 , \40078 , \40062 );
not \g135252/U$1 ( \40080 , \40079 );
not \g133664/U$3 ( \40081 , \40080 );
not \g135428/U$1 ( \40082 , \40074 );
and \g135334/U$2 ( \40083 , \40076 , \40082 );
nor \g135388/U$1 ( \40084 , \40076 , \40082 );
nor \g135334/U$1 ( \40085 , \40083 , \40084 );
not \g135345/U$3 ( \40086 , \40062 );
not \g135345/U$4 ( \40087 , \40076 );
and \g135345/U$2 ( \40088 , \40086 , \40087 );
and \g135345/U$5 ( \40089 , \40062 , \40076 );
nor \g135345/U$1 ( \40090 , \40088 , \40089 );
and \g135232/U$1 ( \40091 , \40085 , \40090 );
nand \g135155/U$1 ( \40092 , \40064 , \40091 );
and \g134645/U$2 ( \40093 , \40092 , \40079 );
not \g134645/U$4 ( \40094 , \40092 );
and \g134645/U$3 ( \40095 , \40094 , \40080 );
nor \g134645/U$1 ( \40096 , \40093 , \40095 );
not \g133875/U$3 ( \40097 , \40096 );
not \g133875/U$4 ( \40098 , \40069 );
and \g133875/U$2 ( \40099 , \40097 , \40098 );
and \g133884/U$2 ( \40100 , \40096 , \40069 );
xnor \g135443/U$1 ( \40101 , \37924 , \37681 );
not \g135263/U$3 ( \40102 , \40101 );
xnor \g135408/U$1 ( \40103 , \38414 , \38168 );
not \g135263/U$4 ( \40104 , \40103 );
and \g135263/U$2 ( \40105 , \40102 , \40104 );
nor \g135263/U$1 ( \40106 , \40105 , \40074 );
not \g135262/U$1 ( \40107 , \40106 );
and \g135457/U$1 ( \40108 , \39932 , \39933 );
not \g135579/U$2 ( \40109 , \40108 );
nor \g135579/U$1 ( \40110 , \40109 , \40062 );
xor \g134035/U$4 ( \40111 , \40107 , \40110 );
and \g135119/U$2 ( \40112 , \40091 , \40067 );
not \g135285/U$1 ( \40113 , \40085 );
and \g135119/U$3 ( \40114 , \40064 , \40113 );
nor \g135119/U$1 ( \40115 , \40112 , \40114 );
and \g134598/U$2 ( \40116 , \40115 , \40080 );
not \g134598/U$4 ( \40117 , \40115 );
and \g134598/U$3 ( \40118 , \40117 , \40079 );
nor \g134598/U$1 ( \40119 , \40116 , \40118 );
and \g134035/U$3 ( \40120 , \40111 , \40119 );
and \g134035/U$5 ( \40121 , \40107 , \40110 );
or \g134035/U$2 ( \40122 , \40120 , \40121 );
not \g134034/U$1 ( \40123 , \40122 );
nor \g133884/U$1 ( \40124 , \40100 , \40123 );
nor \g133875/U$1 ( \40125 , \40099 , \40124 );
not \g133664/U$4 ( \40126 , \40125 );
or \g133664/U$2 ( \40127 , \40081 , \40126 );
or \g133664/U$5 ( \40128 , \40125 , \40080 );
nand \g133664/U$1 ( \40129 , \40127 , \40128 );
not \g129493/U$3 ( \40130 , \40129 );
xnor \g135415/U$1 ( \40131 , \36948 , \36703 );
not \g135251/U$3 ( \40132 , \40131 );
xnor \g135439/U$1 ( \40133 , \37437 , \37191 );
not \g135251/U$4 ( \40134 , \40133 );
and \g135251/U$2 ( \40135 , \40132 , \40134 );
nor \g135251/U$1 ( \40136 , \40135 , \40101 );
not \g135250/U$1 ( \40137 , \40136 );
and \g135463/U$1 ( \40138 , \39928 , \39929 );
not \g135582/U$2 ( \40139 , \40138 );
nor \g135582/U$1 ( \40140 , \40139 , \40062 );
xor \g134039/U$1 ( \40141 , \40137 , \40140 );
xnor \g455964/U$1 ( \40142 , \40103 , \40101 );
and \g135339/U$2 ( \40143 , \40103 , \40074 );
not \g135339/U$4 ( \40144 , \40103 );
and \g135339/U$3 ( \40145 , \40144 , \40082 );
nor \g135339/U$1 ( \40146 , \40143 , \40145 );
and \g135235/U$1 ( \40147 , \40142 , \40146 );
and \g134979/U$2 ( \40148 , \40147 , \40067 );
not \g135277/U$1 ( \40149 , \40142 );
and \g134979/U$3 ( \40150 , \40064 , \40149 );
nor \g134979/U$1 ( \40151 , \40148 , \40150 );
and \g134467/U$2 ( \40152 , \40151 , \40107 );
not \g134467/U$4 ( \40153 , \40151 );
and \g134467/U$3 ( \40154 , \40153 , \40106 );
nor \g134467/U$1 ( \40155 , \40152 , \40154 );
xor \g134039/U$1_r1 ( \40156 , \40141 , \40155 );
not \g133646/U$3 ( \40157 , \40156 );
and \g135453/U$1 ( \40158 , \39930 , \39931 );
and \g134872/U$2 ( \40159 , \40091 , \40158 );
and \g134872/U$3 ( \40160 , \40108 , \40113 );
nor \g134872/U$1 ( \40161 , \40159 , \40160 );
and \g134374/U$2 ( \40162 , \40161 , \40080 );
not \g134374/U$4 ( \40163 , \40161 );
and \g134374/U$3 ( \40164 , \40163 , \40079 );
nor \g134374/U$1 ( \40165 , \40162 , \40164 );
not \g135414/U$1 ( \40166 , \40131 );
and \g135321/U$2 ( \40167 , \40133 , \40166 );
nor \g135384/U$1 ( \40168 , \40133 , \40166 );
nor \g135321/U$1 ( \40169 , \40167 , \40168 );
not \g135328/U$3 ( \40170 , \40133 );
not \g135328/U$4 ( \40171 , \40101 );
and \g135328/U$2 ( \40172 , \40170 , \40171 );
and \g135328/U$5 ( \40173 , \40101 , \40133 );
nor \g135328/U$1 ( \40174 , \40172 , \40173 );
and \g135233/U$1 ( \40175 , \40169 , \40174 );
nand \g135143/U$1 ( \40176 , \40064 , \40175 );
and \g134663/U$2 ( \40177 , \40176 , \40137 );
not \g134663/U$4 ( \40178 , \40176 );
and \g134663/U$3 ( \40179 , \40178 , \40136 );
nor \g134663/U$1 ( \40180 , \40177 , \40179 );
xor \g133767/U$1 ( \40181 , \40165 , \40180 );
and \g135082/U$2 ( \40182 , \40147 , \40108 );
and \g135082/U$3 ( \40183 , \40067 , \40149 );
nor \g135082/U$1 ( \40184 , \40182 , \40183 );
and \g134457/U$2 ( \40185 , \40184 , \40107 );
not \g134457/U$4 ( \40186 , \40184 );
and \g134457/U$3 ( \40187 , \40186 , \40106 );
nor \g134457/U$1 ( \40188 , \40185 , \40187 );
and \g135500/U$1 ( \40189 , \39926 , \39927 );
not \g135599/U$2 ( \40190 , \40189 );
nor \g135599/U$1 ( \40191 , \40190 , \40062 );
xor \g133997/U$4 ( \40192 , \40188 , \40191 );
and \g134968/U$2 ( \40193 , \40091 , \40138 );
and \g134968/U$3 ( \40194 , \40158 , \40113 );
nor \g134968/U$1 ( \40195 , \40193 , \40194 );
or \g134154/U$2 ( \40196 , \40195 , \40079 );
nand \g134633/U$1 ( \40197 , \40079 , \40195 );
nand \g134154/U$1 ( \40198 , \40196 , \40197 );
and \g133997/U$3 ( \40199 , \40192 , \40198 );
and \g133997/U$5 ( \40200 , \40188 , \40191 );
or \g133997/U$2 ( \40201 , \40199 , \40200 );
xor \g133767/U$1_r1 ( \40202 , \40181 , \40201 );
not \g133646/U$4 ( \40203 , \40202 );
or \g133646/U$2 ( \40204 , \40157 , \40203 );
or \g133661/U$2 ( \40205 , \40202 , \40156 );
and \g134987/U$2 ( \40206 , \40175 , \40067 );
not \g135282/U$1 ( \40207 , \40169 );
and \g134987/U$3 ( \40208 , \40064 , \40207 );
nor \g134987/U$1 ( \40209 , \40206 , \40208 );
and \g134586/U$2 ( \40210 , \40209 , \40137 );
not \g134586/U$4 ( \40211 , \40209 );
and \g134586/U$3 ( \40212 , \40211 , \40136 );
nor \g134586/U$1 ( \40213 , \40210 , \40212 );
xnor \g135441/U$1 ( \40214 , \35974 , \35732 );
not \g135267/U$3 ( \40215 , \40214 );
xnor \g135398/U$1 ( \40216 , \36459 , \36217 );
not \g135267/U$4 ( \40217 , \40216 );
and \g135267/U$2 ( \40218 , \40215 , \40217 );
nor \g135267/U$1 ( \40219 , \40218 , \40131 );
not \g135266/U$1 ( \40220 , \40219 );
xor \g134015/U$4 ( \40221 , \40213 , \40220 );
and \g135085/U$2 ( \40222 , \40091 , \40189 );
and \g135085/U$3 ( \40223 , \40138 , \40113 );
nor \g135085/U$1 ( \40224 , \40222 , \40223 );
and \g134493/U$2 ( \40225 , \40224 , \40080 );
not \g134493/U$4 ( \40226 , \40224 );
and \g134493/U$3 ( \40227 , \40226 , \40079 );
nor \g134493/U$1 ( \40228 , \40225 , \40227 );
and \g134015/U$3 ( \40229 , \40221 , \40228 );
and \g134015/U$5 ( \40230 , \40213 , \40220 );
or \g134015/U$2 ( \40231 , \40229 , \40230 );
not \g134662/U$1 ( \40232 , \40180 );
xor \g133748/U$4 ( \40233 , \40231 , \40232 );
xor \g133997/U$1 ( \40234 , \40188 , \40191 );
xor \g133997/U$1_r1 ( \40235 , \40234 , \40198 );
and \g133748/U$3 ( \40236 , \40233 , \40235 );
and \g133748/U$5 ( \40237 , \40231 , \40232 );
or \g133748/U$2 ( \40238 , \40236 , \40237 );
nand \g133661/U$1 ( \40239 , \40205 , \40238 );
nand \g133646/U$1 ( \40240 , \40204 , \40239 );
nand \g135148/U$1 ( \40241 , \40064 , \40147 );
and \g134647/U$2 ( \40242 , \40241 , \40106 );
not \g134647/U$4 ( \40243 , \40241 );
and \g134647/U$3 ( \40244 , \40243 , \40107 );
nor \g134647/U$1 ( \40245 , \40242 , \40244 );
not \g135577/U$2 ( \40246 , \40158 );
nor \g135577/U$1 ( \40247 , \40246 , \40062 );
xor \g134006/U$1 ( \40248 , \40245 , \40247 );
and \g135053/U$2 ( \40249 , \40091 , \40108 );
and \g135053/U$3 ( \40250 , \40067 , \40113 );
nor \g135053/U$1 ( \40251 , \40249 , \40250 );
and \g134355/U$2 ( \40252 , \40251 , \40080 );
not \g134355/U$4 ( \40253 , \40251 );
and \g134355/U$3 ( \40254 , \40253 , \40079 );
nor \g134355/U$1 ( \40255 , \40252 , \40254 );
xor \g134006/U$1_r1 ( \40256 , \40248 , \40255 );
xor \g133767/U$4 ( \40257 , \40165 , \40180 );
and \g133767/U$3 ( \40258 , \40257 , \40201 );
and \g133767/U$5 ( \40259 , \40165 , \40180 );
or \g133767/U$2 ( \40260 , \40258 , \40259 );
xor \g456235/U$1 ( \40261 , \40256 , \40260 );
xor \g134039/U$4 ( \40262 , \40137 , \40140 );
and \g134039/U$3 ( \40263 , \40262 , \40155 );
and \g134039/U$5 ( \40264 , \40137 , \40140 );
or \g134039/U$2 ( \40265 , \40263 , \40264 );
xor \g456235/U$1_r1 ( \40266 , \40261 , \40265 );
and \g129735/U$2 ( \40267 , \40240 , \40266 );
xor \g133507/U$1 ( \40268 , \40266 , \40240 );
xor \g133748/U$1 ( \40269 , \40231 , \40232 );
xor \g133748/U$1_r1 ( \40270 , \40269 , \40235 );
and \g134850/U$2 ( \40271 , \40147 , \40158 );
and \g134850/U$3 ( \40272 , \40108 , \40149 );
nor \g134850/U$1 ( \40273 , \40271 , \40272 );
and \g134340/U$2 ( \40274 , \40273 , \40107 );
not \g134340/U$4 ( \40275 , \40273 );
and \g134340/U$3 ( \40276 , \40275 , \40106 );
nor \g134340/U$1 ( \40277 , \40274 , \40276 );
and \g135482/U$1 ( \40278 , \39924 , \39925 );
not \g135591/U$2 ( \40279 , \40278 );
nor \g135591/U$1 ( \40280 , \40279 , \40062 );
xor \g134033/U$4 ( \40281 , \40277 , \40280 );
and \g134867/U$2 ( \40282 , \40175 , \40108 );
and \g134867/U$3 ( \40283 , \40067 , \40207 );
nor \g134867/U$1 ( \40284 , \40282 , \40283 );
and \g134292/U$2 ( \40285 , \40284 , \40136 );
not \g134292/U$4 ( \40286 , \40284 );
and \g134292/U$3 ( \40287 , \40286 , \40137 );
nor \g134292/U$1 ( \40288 , \40285 , \40287 );
not \g134291/U$1 ( \40289 , \40288 );
and \g134033/U$3 ( \40290 , \40281 , \40289 );
and \g134033/U$5 ( \40291 , \40277 , \40280 );
or \g134033/U$2 ( \40292 , \40290 , \40291 );
xor \g456233/U$4 ( \40293 , \40270 , \40292 );
xor \g134015/U$1 ( \40294 , \40213 , \40220 );
xor \g134015/U$1_r1 ( \40295 , \40294 , \40228 );
xnor \g455965/U$1 ( \40296 , \40216 , \40214 );
and \g135338/U$2 ( \40297 , \40216 , \40131 );
not \g135338/U$4 ( \40298 , \40216 );
and \g135338/U$3 ( \40299 , \40298 , \40166 );
nor \g135338/U$1 ( \40300 , \40297 , \40299 );
and \g135227/U$1 ( \40301 , \40296 , \40300 );
nand \g135151/U$1 ( \40302 , \40064 , \40301 );
and \g134667/U$2 ( \40303 , \40302 , \40220 );
not \g134667/U$4 ( \40304 , \40302 );
and \g134667/U$3 ( \40305 , \40304 , \40219 );
nor \g134667/U$1 ( \40306 , \40303 , \40305 );
and \g135473/U$1 ( \40307 , \39922 , \39923 );
not \g135587/U$2 ( \40308 , \40307 );
nor \g135587/U$1 ( \40309 , \40308 , \40062 );
xor \g133971/U$4 ( \40310 , \40306 , \40309 );
and \g134995/U$2 ( \40311 , \40091 , \40278 );
and \g134995/U$3 ( \40312 , \40189 , \40113 );
nor \g134995/U$1 ( \40313 , \40311 , \40312 );
and \g134244/U$2 ( \40314 , \40313 , \40080 );
not \g134244/U$4 ( \40315 , \40313 );
and \g134244/U$3 ( \40316 , \40315 , \40079 );
nor \g134244/U$1 ( \40317 , \40314 , \40316 );
and \g133971/U$3 ( \40318 , \40310 , \40317 );
and \g133971/U$5 ( \40319 , \40306 , \40309 );
or \g133971/U$2 ( \40320 , \40318 , \40319 );
xor \g456208/U$5 ( \40321 , \40295 , \40320 );
xor \g134033/U$1 ( \40322 , \40277 , \40280 );
xor \g134033/U$1_r1 ( \40323 , \40322 , \40289 );
and \g456208/U$4 ( \40324 , \40321 , \40323 );
and \g456208/U$6 ( \40325 , \40295 , \40320 );
or \g456208/U$3 ( \40326 , \40324 , \40325 );
and \g456233/U$3 ( \40327 , \40293 , \40326 );
and \g456233/U$5 ( \40328 , \40270 , \40292 );
nor \g456233/U$2 ( \40329 , \40327 , \40328 );
xnor \g455960/U$1 ( \40330 , \40238 , \40156 );
not \g133614/U$3 ( \40331 , \40330 );
not \g133614/U$4 ( \40332 , \40202 );
and \g133614/U$2 ( \40333 , \40331 , \40332 );
and \g133614/U$5 ( \40334 , \40330 , \40202 );
nor \g133614/U$1 ( \40335 , \40333 , \40334 );
or \g129824/U$2 ( \40336 , \40329 , \40335 );
xnor \g133506/U$1 ( \40337 , \40335 , \40329 );
and \g134706/U$2 ( \40338 , \40147 , \40138 );
and \g134706/U$3 ( \40339 , \40158 , \40149 );
nor \g134706/U$1 ( \40340 , \40338 , \40339 );
and \g134528/U$2 ( \40341 , \40340 , \40107 );
not \g134528/U$4 ( \40342 , \40340 );
and \g134528/U$3 ( \40343 , \40342 , \40106 );
nor \g134528/U$1 ( \40344 , \40341 , \40343 );
xor \g133794/U$4 ( \40345 , \40288 , \40344 );
and \g134745/U$2 ( \40346 , \40091 , \40307 );
and \g134745/U$3 ( \40347 , \40278 , \40113 );
nor \g134745/U$1 ( \40348 , \40346 , \40347 );
and \g134581/U$2 ( \40349 , \40348 , \40080 );
not \g134581/U$4 ( \40350 , \40348 );
and \g134581/U$3 ( \40351 , \40350 , \40079 );
nor \g134581/U$1 ( \40352 , \40349 , \40351 );
and \g135451/U$1 ( \40353 , \39920 , \39921 );
not \g135576/U$2 ( \40354 , \40353 );
nor \g135576/U$1 ( \40355 , \40354 , \40062 );
xor \g133945/U$4 ( \40356 , \40352 , \40355 );
and \g134764/U$2 ( \40357 , \40175 , \40158 );
and \g134764/U$3 ( \40358 , \40108 , \40207 );
nor \g134764/U$1 ( \40359 , \40357 , \40358 );
and \g134593/U$2 ( \40360 , \40359 , \40137 );
not \g134593/U$4 ( \40361 , \40359 );
and \g134593/U$3 ( \40362 , \40361 , \40136 );
nor \g134593/U$1 ( \40363 , \40360 , \40362 );
and \g133945/U$3 ( \40364 , \40356 , \40363 );
and \g133945/U$5 ( \40365 , \40352 , \40355 );
or \g133945/U$2 ( \40366 , \40364 , \40365 );
and \g133794/U$3 ( \40367 , \40345 , \40366 );
and \g133794/U$5 ( \40368 , \40288 , \40344 );
or \g133794/U$2 ( \40369 , \40367 , \40368 );
xor \g456208/U$9 ( \40370 , \40295 , \40320 );
xor \g456208/U$9_r1 ( \40371 , \40370 , \40323 );
and \g456208/U$8 ( \40372 , \40369 , \40371 );
xor \g133971/U$1 ( \40373 , \40306 , \40309 );
xor \g133971/U$1_r1 ( \40374 , \40373 , \40317 );
and \g134949/U$2 ( \40375 , \40147 , \40189 );
and \g134949/U$3 ( \40376 , \40138 , \40149 );
nor \g134949/U$1 ( \40377 , \40375 , \40376 );
and \g134271/U$2 ( \40378 , \40377 , \40107 );
not \g134271/U$4 ( \40379 , \40377 );
and \g134271/U$3 ( \40380 , \40379 , \40106 );
nor \g134271/U$1 ( \40381 , \40378 , \40380 );
xnor \g135412/U$1 ( \40382 , \35003 , \34756 );
not \g135255/U$3 ( \40383 , \40382 );
xnor \g135413/U$1 ( \40384 , \35489 , \35245 );
not \g135255/U$4 ( \40385 , \40384 );
and \g135255/U$2 ( \40386 , \40383 , \40385 );
nor \g135255/U$1 ( \40387 , \40386 , \40214 );
not \g135254/U$1 ( \40388 , \40387 );
xor \g456236/U$5 ( \40389 , \40381 , \40388 );
and \g135021/U$2 ( \40390 , \40301 , \40067 );
not \g135280/U$1 ( \40391 , \40296 );
and \g135021/U$3 ( \40392 , \40064 , \40391 );
nor \g135021/U$1 ( \40393 , \40390 , \40392 );
and \g134402/U$2 ( \40394 , \40393 , \40220 );
not \g134402/U$4 ( \40395 , \40393 );
and \g134402/U$3 ( \40396 , \40395 , \40219 );
nor \g134402/U$1 ( \40397 , \40394 , \40396 );
and \g456236/U$4 ( \40398 , \40389 , \40397 );
and \g456236/U$6 ( \40399 , \40381 , \40388 );
or \g456236/U$3 ( \40400 , \40398 , \40399 );
xor \g456209/U$5 ( \40401 , \40374 , \40400 );
xor \g133794/U$1 ( \40402 , \40288 , \40344 );
xor \g133794/U$1_r1 ( \40403 , \40402 , \40366 );
and \g456209/U$4 ( \40404 , \40401 , \40403 );
and \g456209/U$6 ( \40405 , \40374 , \40400 );
or \g456209/U$3 ( \40406 , \40404 , \40405 );
xor \g456208/U$11 ( \40407 , \40295 , \40320 );
xor \g456208/U$11_r1 ( \40408 , \40407 , \40323 );
and \g456208/U$10 ( \40409 , \40406 , \40408 );
and \g456208/U$12 ( \40410 , \40369 , \40406 );
or \g456208/U$7 ( \40411 , \40372 , \40409 , \40410 );
xor \g456233/U$1 ( \40412 , \40270 , \40292 );
xor \g456233/U$1_r1 ( \40413 , \40412 , \40326 );
and \g129915/U$2 ( \40414 , \40411 , \40413 );
xor \g133467/U$1 ( \40415 , \40413 , \40411 );
and \g134694/U$2 ( \40416 , \40147 , \40278 );
and \g134694/U$3 ( \40417 , \40189 , \40149 );
nor \g134694/U$1 ( \40418 , \40416 , \40417 );
and \g134398/U$2 ( \40419 , \40418 , \40107 );
not \g134398/U$4 ( \40420 , \40418 );
and \g134398/U$3 ( \40421 , \40420 , \40106 );
nor \g134398/U$1 ( \40422 , \40419 , \40421 );
not \g135411/U$1 ( \40423 , \40382 );
and \g135322/U$2 ( \40424 , \40384 , \40423 );
nor \g135390/U$1 ( \40425 , \40384 , \40423 );
nor \g135322/U$1 ( \40426 , \40424 , \40425 );
not \g135326/U$3 ( \40427 , \40384 );
not \g135326/U$4 ( \40428 , \40214 );
and \g135326/U$2 ( \40429 , \40427 , \40428 );
and \g135326/U$5 ( \40430 , \40214 , \40384 );
nor \g135326/U$1 ( \40431 , \40429 , \40430 );
and \g135234/U$1 ( \40432 , \40426 , \40431 );
nand \g135153/U$1 ( \40433 , \40064 , \40432 );
and \g134655/U$2 ( \40434 , \40433 , \40388 );
not \g134655/U$4 ( \40435 , \40433 );
and \g134655/U$3 ( \40436 , \40435 , \40387 );
nor \g134655/U$1 ( \40437 , \40434 , \40436 );
xor \g134013/U$4 ( \40438 , \40422 , \40437 );
and \g134713/U$2 ( \40439 , \40091 , \40353 );
and \g134713/U$3 ( \40440 , \40307 , \40113 );
nor \g134713/U$1 ( \40441 , \40439 , \40440 );
and \g134172/U$2 ( \40442 , \40441 , \40080 );
not \g134172/U$4 ( \40443 , \40441 );
and \g134172/U$3 ( \40444 , \40443 , \40079 );
nor \g134172/U$1 ( \40445 , \40442 , \40444 );
and \g134013/U$3 ( \40446 , \40438 , \40445 );
and \g134013/U$5 ( \40447 , \40422 , \40437 );
or \g134013/U$2 ( \40448 , \40446 , \40447 );
and \g134952/U$2 ( \40449 , \40301 , \40108 );
and \g134952/U$3 ( \40450 , \40067 , \40391 );
nor \g134952/U$1 ( \40451 , \40449 , \40450 );
and \g134167/U$2 ( \40452 , \40451 , \40220 );
not \g134167/U$4 ( \40453 , \40451 );
and \g134167/U$3 ( \40454 , \40453 , \40219 );
nor \g134167/U$1 ( \40455 , \40452 , \40454 );
xor \g133791/U$4 ( \40456 , \40448 , \40455 );
xor \g133945/U$1 ( \40457 , \40352 , \40355 );
xor \g133945/U$1_r1 ( \40458 , \40457 , \40363 );
and \g133791/U$3 ( \40459 , \40456 , \40458 );
and \g133791/U$5 ( \40460 , \40448 , \40455 );
or \g133791/U$2 ( \40461 , \40459 , \40460 );
xor \g456209/U$9 ( \40462 , \40374 , \40400 );
xor \g456209/U$9_r1 ( \40463 , \40462 , \40403 );
and \g456209/U$8 ( \40464 , \40461 , \40463 );
and \g134842/U$2 ( \40465 , \40175 , \40138 );
and \g134842/U$3 ( \40466 , \40158 , \40207 );
nor \g134842/U$1 ( \40467 , \40465 , \40466 );
and \g134212/U$2 ( \40468 , \40467 , \40137 );
not \g134212/U$4 ( \40469 , \40467 );
and \g134212/U$3 ( \40470 , \40469 , \40136 );
nor \g134212/U$1 ( \40471 , \40468 , \40470 );
and \g135465/U$1 ( \40472 , \39918 , \39919 );
not \g135583/U$2 ( \40473 , \40472 );
nor \g135583/U$1 ( \40474 , \40473 , \40062 );
xor \g133963/U$4 ( \40475 , \40471 , \40474 );
not \g134166/U$1 ( \40476 , \40455 );
and \g133963/U$3 ( \40477 , \40475 , \40476 );
and \g133963/U$5 ( \40478 , \40471 , \40474 );
or \g133963/U$2 ( \40479 , \40477 , \40478 );
xor \g456236/U$9 ( \40480 , \40381 , \40388 );
xor \g456236/U$9_r1 ( \40481 , \40480 , \40397 );
and \g456236/U$8 ( \40482 , \40479 , \40481 );
xor \g133791/U$1 ( \40483 , \40448 , \40455 );
xor \g133791/U$1_r1 ( \40484 , \40483 , \40458 );
xor \g456236/U$11 ( \40485 , \40381 , \40388 );
xor \g456236/U$11_r1 ( \40486 , \40485 , \40397 );
and \g456236/U$10 ( \40487 , \40484 , \40486 );
and \g456236/U$12 ( \40488 , \40479 , \40484 );
or \g456236/U$7 ( \40489 , \40482 , \40487 , \40488 );
xor \g456209/U$11 ( \40490 , \40374 , \40400 );
xor \g456209/U$11_r1 ( \40491 , \40490 , \40403 );
and \g456209/U$10 ( \40492 , \40489 , \40491 );
and \g456209/U$12 ( \40493 , \40461 , \40489 );
or \g456209/U$7 ( \40494 , \40464 , \40492 , \40493 );
not \g130012/U$3 ( \40495 , \40494 );
xor \g456208/U$2 ( \40496 , \40295 , \40320 );
xor \g456208/U$1 ( \40497 , \40496 , \40323 );
xor \g456208/U$1_r1 ( \40498 , \40369 , \40406 );
xor \g456208/U$1_r2 ( \40499 , \40497 , \40498 );
not \g130012/U$4 ( \40500 , \40499 );
or \g130012/U$2 ( \40501 , \40495 , \40500 );
xor \g456209/U$2 ( \40502 , \40374 , \40400 );
xor \g456209/U$1 ( \40503 , \40502 , \40403 );
xor \g456209/U$1_r1 ( \40504 , \40461 , \40489 );
xor \g456209/U$1_r2 ( \40505 , \40503 , \40504 );
xnor \g135432/U$1 ( \40506 , \34513 , \34270 );
xnor \g135422/U$1 ( \40507 , \34027 , \33786 );
xnor \g455967/U$1 ( \40508 , \40506 , \40507 );
and \g135347/U$2 ( \40509 , \40506 , \40382 );
not \g135347/U$4 ( \40510 , \40506 );
and \g135347/U$3 ( \40511 , \40510 , \40423 );
nor \g135347/U$1 ( \40512 , \40509 , \40511 );
and \g135231/U$1 ( \40513 , \40508 , \40512 );
nand \g135147/U$1 ( \40514 , \40064 , \40513 );
not \g135257/U$3 ( \40515 , \40507 );
not \g135257/U$4 ( \40516 , \40506 );
and \g135257/U$2 ( \40517 , \40515 , \40516 );
nor \g135257/U$1 ( \40518 , \40517 , \40382 );
and \g134666/U$2 ( \40519 , \40514 , \40518 );
not \g134666/U$4 ( \40520 , \40514 );
not \g135256/U$1 ( \40521 , \40518 );
and \g134666/U$3 ( \40522 , \40520 , \40521 );
nor \g134666/U$1 ( \40523 , \40519 , \40522 );
not \g134665/U$1 ( \40524 , \40523 );
and \g135496/U$1 ( \40525 , \39916 , \39917 );
not \g135597/U$2 ( \40526 , \40525 );
nor \g135597/U$1 ( \40527 , \40526 , \40062 );
xor \g133775/U$4 ( \40528 , \40524 , \40527 );
and \g134753/U$2 ( \40529 , \40432 , \40108 );
not \g135275/U$1 ( \40530 , \40426 );
and \g134753/U$3 ( \40531 , \40067 , \40530 );
nor \g134753/U$1 ( \40532 , \40529 , \40531 );
and \g134370/U$2 ( \40533 , \40532 , \40388 );
not \g134370/U$4 ( \40534 , \40532 );
and \g134370/U$3 ( \40535 , \40534 , \40387 );
nor \g134370/U$1 ( \40536 , \40533 , \40535 );
and \g134956/U$2 ( \40537 , \40175 , \40278 );
and \g134956/U$3 ( \40538 , \40189 , \40207 );
nor \g134956/U$1 ( \40539 , \40537 , \40538 );
and \g134572/U$2 ( \40540 , \40539 , \40137 );
not \g134572/U$4 ( \40541 , \40539 );
and \g134572/U$3 ( \40542 , \40541 , \40136 );
nor \g134572/U$1 ( \40543 , \40540 , \40542 );
xor \g134041/U$4 ( \40544 , \40536 , \40543 );
and \g135134/U$2 ( \40545 , \40147 , \40353 );
and \g135134/U$3 ( \40546 , \40307 , \40149 );
nor \g135134/U$1 ( \40547 , \40545 , \40546 );
and \g134198/U$2 ( \40548 , \40547 , \40107 );
not \g134198/U$4 ( \40549 , \40547 );
and \g134198/U$3 ( \40550 , \40549 , \40106 );
nor \g134198/U$1 ( \40551 , \40548 , \40550 );
and \g134041/U$3 ( \40552 , \40544 , \40551 );
and \g134041/U$5 ( \40553 , \40536 , \40543 );
or \g134041/U$2 ( \40554 , \40552 , \40553 );
and \g133775/U$3 ( \40555 , \40528 , \40554 );
and \g133775/U$5 ( \40556 , \40524 , \40527 );
or \g133775/U$2 ( \40557 , \40555 , \40556 );
xor \g133963/U$1 ( \40558 , \40471 , \40474 );
xor \g133963/U$1_r1 ( \40559 , \40558 , \40476 );
xor \g133588/U$4 ( \40560 , \40557 , \40559 );
and \g134788/U$2 ( \40561 , \40091 , \40525 );
and \g134788/U$3 ( \40562 , \40472 , \40113 );
nor \g134788/U$1 ( \40563 , \40561 , \40562 );
and \g134312/U$2 ( \40564 , \40563 , \40080 );
not \g134312/U$4 ( \40565 , \40563 );
and \g134312/U$3 ( \40566 , \40565 , \40079 );
nor \g134312/U$1 ( \40567 , \40564 , \40566 );
and \g135467/U$1 ( \40568 , \39914 , \39915 );
not \g135584/U$2 ( \40569 , \40568 );
nor \g135584/U$1 ( \40570 , \40569 , \40062 );
xor \g456267/U$5 ( \40571 , \40567 , \40570 );
and \g134771/U$2 ( \40572 , \40301 , \40138 );
and \g134771/U$3 ( \40573 , \40158 , \40391 );
nor \g134771/U$1 ( \40574 , \40572 , \40573 );
and \g134155/U$2 ( \40575 , \40574 , \40220 );
not \g134155/U$4 ( \40576 , \40574 );
and \g134155/U$3 ( \40577 , \40576 , \40219 );
nor \g134155/U$1 ( \40578 , \40575 , \40577 );
and \g456267/U$4 ( \40579 , \40571 , \40578 );
and \g456267/U$6 ( \40580 , \40567 , \40570 );
or \g456267/U$3 ( \40581 , \40579 , \40580 );
and \g134983/U$2 ( \40582 , \40301 , \40158 );
and \g134983/U$3 ( \40583 , \40108 , \40391 );
nor \g134983/U$1 ( \40584 , \40582 , \40583 );
and \g134465/U$2 ( \40585 , \40584 , \40220 );
not \g134465/U$4 ( \40586 , \40584 );
and \g134465/U$3 ( \40587 , \40586 , \40219 );
nor \g134465/U$1 ( \40588 , \40585 , \40587 );
and \g135117/U$2 ( \40589 , \40147 , \40307 );
and \g135117/U$3 ( \40590 , \40278 , \40149 );
nor \g135117/U$1 ( \40591 , \40589 , \40590 );
and \g134184/U$2 ( \40592 , \40591 , \40107 );
not \g134184/U$4 ( \40593 , \40591 );
and \g134184/U$3 ( \40594 , \40593 , \40106 );
nor \g134184/U$1 ( \40595 , \40592 , \40594 );
xor \g456255/U$9 ( \40596 , \40588 , \40595 );
and \g135090/U$2 ( \40597 , \40091 , \40472 );
and \g135090/U$3 ( \40598 , \40353 , \40113 );
nor \g135090/U$1 ( \40599 , \40597 , \40598 );
and \g134481/U$2 ( \40600 , \40599 , \40080 );
not \g134481/U$4 ( \40601 , \40599 );
and \g134481/U$3 ( \40602 , \40601 , \40079 );
nor \g134481/U$1 ( \40603 , \40600 , \40602 );
xor \g456255/U$9_r1 ( \40604 , \40596 , \40603 );
and \g456255/U$8 ( \40605 , \40581 , \40604 );
and \g134915/U$2 ( \40606 , \40432 , \40067 );
and \g134915/U$3 ( \40607 , \40064 , \40530 );
nor \g134915/U$1 ( \40608 , \40606 , \40607 );
and \g134438/U$2 ( \40609 , \40608 , \40388 );
not \g134438/U$4 ( \40610 , \40608 );
and \g134438/U$3 ( \40611 , \40610 , \40387 );
nor \g134438/U$1 ( \40612 , \40609 , \40611 );
xor \g133943/U$1 ( \40613 , \40612 , \40521 );
and \g135000/U$2 ( \40614 , \40175 , \40189 );
and \g135000/U$3 ( \40615 , \40138 , \40207 );
nor \g135000/U$1 ( \40616 , \40614 , \40615 );
and \g134532/U$2 ( \40617 , \40616 , \40137 );
not \g134532/U$4 ( \40618 , \40616 );
and \g134532/U$3 ( \40619 , \40618 , \40136 );
nor \g134532/U$1 ( \40620 , \40617 , \40619 );
xor \g133943/U$1_r1 ( \40621 , \40613 , \40620 );
xor \g456255/U$11 ( \40622 , \40588 , \40595 );
xor \g456255/U$11_r1 ( \40623 , \40622 , \40603 );
and \g456255/U$10 ( \40624 , \40621 , \40623 );
and \g456255/U$12 ( \40625 , \40581 , \40621 );
or \g456255/U$7 ( \40626 , \40605 , \40624 , \40625 );
and \g133588/U$3 ( \40627 , \40560 , \40626 );
and \g133588/U$5 ( \40628 , \40557 , \40559 );
or \g133588/U$2 ( \40629 , \40627 , \40628 );
xor \g456255/U$5 ( \40630 , \40588 , \40595 );
and \g456255/U$4 ( \40631 , \40630 , \40603 );
and \g456255/U$6 ( \40632 , \40588 , \40595 );
or \g456255/U$3 ( \40633 , \40631 , \40632 );
xor \g133943/U$4 ( \40634 , \40612 , \40521 );
and \g133943/U$3 ( \40635 , \40634 , \40620 );
and \g133943/U$5 ( \40636 , \40612 , \40521 );
or \g133943/U$2 ( \40637 , \40635 , \40636 );
xor \g133793/U$4 ( \40638 , \40633 , \40637 );
xor \g134013/U$1 ( \40639 , \40422 , \40437 );
xor \g134013/U$1_r1 ( \40640 , \40639 , \40445 );
and \g133793/U$3 ( \40641 , \40638 , \40640 );
and \g133793/U$5 ( \40642 , \40633 , \40637 );
or \g133793/U$2 ( \40643 , \40641 , \40642 );
xor \g133457/U$4 ( \40644 , \40629 , \40643 );
xor \g456236/U$2 ( \40645 , \40381 , \40388 );
xor \g456236/U$1 ( \40646 , \40645 , \40397 );
xor \g456236/U$1_r1 ( \40647 , \40479 , \40484 );
xor \g456236/U$1_r2 ( \40648 , \40646 , \40647 );
and \g133457/U$3 ( \40649 , \40644 , \40648 );
and \g133457/U$5 ( \40650 , \40629 , \40643 );
or \g133457/U$2 ( \40651 , \40649 , \40650 );
and \g130105/U$2 ( \40652 , \40505 , \40651 );
xor \g133392/U$1 ( \40653 , \40651 , \40505 );
xor \g133457/U$1 ( \40654 , \40629 , \40643 );
xor \g133457/U$1_r1 ( \40655 , \40654 , \40648 );
not \g130180/U$3 ( \40656 , \40655 );
and \g134904/U$2 ( \40657 , \40147 , \40472 );
and \g134904/U$3 ( \40658 , \40353 , \40149 );
nor \g134904/U$1 ( \40659 , \40657 , \40658 );
and \g134609/U$2 ( \40660 , \40659 , \40107 );
not \g134609/U$4 ( \40661 , \40659 );
and \g134609/U$3 ( \40662 , \40661 , \40106 );
nor \g134609/U$1 ( \40663 , \40660 , \40662 );
xnor \g135406/U$1 ( \40664 , \33545 , \33302 );
xnor \g135434/U$1 ( \40665 , \33057 , \32811 );
xnor \g455966/U$1 ( \40666 , \40664 , \40665 );
not \g135336/U$3 ( \40667 , \40664 );
not \g135336/U$4 ( \40668 , \40507 );
and \g135336/U$2 ( \40669 , \40667 , \40668 );
and \g135336/U$5 ( \40670 , \40507 , \40664 );
nor \g135336/U$1 ( \40671 , \40669 , \40670 );
and \g135224/U$1 ( \40672 , \40666 , \40671 );
nand \g135149/U$1 ( \40673 , \40064 , \40672 );
not \g135259/U$3 ( \40674 , \40665 );
not \g135259/U$4 ( \40675 , \40664 );
and \g135259/U$2 ( \40676 , \40674 , \40675 );
nor \g135259/U$1 ( \40677 , \40676 , \40507 );
not \g135258/U$1 ( \40678 , \40677 );
and \g134650/U$2 ( \40679 , \40673 , \40678 );
not \g134650/U$4 ( \40680 , \40673 );
and \g134650/U$3 ( \40681 , \40680 , \40677 );
nor \g134650/U$1 ( \40682 , \40679 , \40681 );
xor \g456231/U$5 ( \40683 , \40663 , \40682 );
and \g134852/U$2 ( \40684 , \40091 , \40568 );
and \g134852/U$3 ( \40685 , \40525 , \40113 );
nor \g134852/U$1 ( \40686 , \40684 , \40685 );
and \g134180/U$2 ( \40687 , \40686 , \40080 );
not \g134180/U$4 ( \40688 , \40686 );
and \g134180/U$3 ( \40689 , \40688 , \40079 );
nor \g134180/U$1 ( \40690 , \40687 , \40689 );
and \g456231/U$4 ( \40691 , \40683 , \40690 );
and \g456231/U$6 ( \40692 , \40663 , \40682 );
or \g456231/U$3 ( \40693 , \40691 , \40692 );
xor \g456267/U$9 ( \40694 , \40567 , \40570 );
xor \g456267/U$9_r1 ( \40695 , \40694 , \40578 );
and \g456267/U$8 ( \40696 , \40693 , \40695 );
xor \g134041/U$1 ( \40697 , \40536 , \40543 );
xor \g134041/U$1_r1 ( \40698 , \40697 , \40551 );
xor \g456267/U$11 ( \40699 , \40567 , \40570 );
xor \g456267/U$11_r1 ( \40700 , \40699 , \40578 );
and \g456267/U$10 ( \40701 , \40698 , \40700 );
and \g456267/U$12 ( \40702 , \40693 , \40698 );
or \g456267/U$7 ( \40703 , \40696 , \40701 , \40702 );
and \g135017/U$2 ( \40704 , \40301 , \40189 );
and \g135017/U$3 ( \40705 , \40138 , \40391 );
nor \g135017/U$1 ( \40706 , \40704 , \40705 );
and \g134567/U$2 ( \40707 , \40706 , \40220 );
not \g134567/U$4 ( \40708 , \40706 );
and \g134567/U$3 ( \40709 , \40708 , \40219 );
nor \g134567/U$1 ( \40710 , \40707 , \40709 );
xor \g133936/U$4 ( \40711 , \40710 , \40678 );
and \g134791/U$2 ( \40712 , \40513 , \40067 );
not \g135276/U$1 ( \40713 , \40508 );
and \g134791/U$3 ( \40714 , \40064 , \40713 );
nor \g134791/U$1 ( \40715 , \40712 , \40714 );
and \g134375/U$2 ( \40716 , \40715 , \40521 );
not \g134375/U$4 ( \40717 , \40715 );
and \g134375/U$3 ( \40718 , \40717 , \40518 );
nor \g134375/U$1 ( \40719 , \40716 , \40718 );
and \g133936/U$3 ( \40720 , \40711 , \40719 );
and \g133936/U$5 ( \40721 , \40710 , \40678 );
or \g133936/U$2 ( \40722 , \40720 , \40721 );
xor \g133699/U$4 ( \40723 , \40722 , \40523 );
and \g135132/U$2 ( \40724 , \40175 , \40307 );
and \g135132/U$3 ( \40725 , \40278 , \40207 );
nor \g135132/U$1 ( \40726 , \40724 , \40725 );
and \g134550/U$2 ( \40727 , \40726 , \40137 );
not \g134550/U$4 ( \40728 , \40726 );
and \g134550/U$3 ( \40729 , \40728 , \40136 );
nor \g134550/U$1 ( \40730 , \40727 , \40729 );
and \g135449/U$1 ( \40731 , \39912 , \39913 );
not \g135575/U$2 ( \40732 , \40731 );
nor \g135575/U$1 ( \40733 , \40732 , \40062 );
xor \g134047/U$4 ( \40734 , \40730 , \40733 );
and \g135130/U$2 ( \40735 , \40432 , \40158 );
and \g135130/U$3 ( \40736 , \40108 , \40530 );
nor \g135130/U$1 ( \40737 , \40735 , \40736 );
and \g134179/U$2 ( \40738 , \40737 , \40388 );
not \g134179/U$4 ( \40739 , \40737 );
and \g134179/U$3 ( \40740 , \40739 , \40387 );
nor \g134179/U$1 ( \40741 , \40738 , \40740 );
and \g134047/U$3 ( \40742 , \40734 , \40741 );
and \g134047/U$5 ( \40743 , \40730 , \40733 );
or \g134047/U$2 ( \40744 , \40742 , \40743 );
and \g133699/U$3 ( \40745 , \40723 , \40744 );
and \g133699/U$5 ( \40746 , \40722 , \40523 );
or \g133699/U$2 ( \40747 , \40745 , \40746 );
xor \g133565/U$4 ( \40748 , \40703 , \40747 );
xor \g133775/U$1 ( \40749 , \40524 , \40527 );
xor \g133775/U$1_r1 ( \40750 , \40749 , \40554 );
and \g133565/U$3 ( \40751 , \40748 , \40750 );
and \g133565/U$5 ( \40752 , \40703 , \40747 );
or \g133565/U$2 ( \40753 , \40751 , \40752 );
xor \g133793/U$1 ( \40754 , \40633 , \40637 );
xor \g133793/U$1_r1 ( \40755 , \40754 , \40640 );
xor \g133418/U$4 ( \40756 , \40753 , \40755 );
xor \g133588/U$1 ( \40757 , \40557 , \40559 );
xor \g133588/U$1_r1 ( \40758 , \40757 , \40626 );
and \g133418/U$3 ( \40759 , \40756 , \40758 );
and \g133418/U$5 ( \40760 , \40753 , \40755 );
or \g133418/U$2 ( \40761 , \40759 , \40760 );
not \g130180/U$4 ( \40762 , \40761 );
or \g130180/U$2 ( \40763 , \40656 , \40762 );
xor \g133418/U$1 ( \40764 , \40753 , \40755 );
xor \g133418/U$1_r1 ( \40765 , \40764 , \40758 );
xor \g133699/U$1 ( \40766 , \40722 , \40523 );
xor \g133699/U$1_r1 ( \40767 , \40766 , \40744 );
and \g134818/U$2 ( \40768 , \40432 , \40138 );
and \g134818/U$3 ( \40769 , \40158 , \40530 );
nor \g134818/U$1 ( \40770 , \40768 , \40769 );
and \g134268/U$2 ( \40771 , \40770 , \40388 );
not \g134268/U$4 ( \40772 , \40770 );
and \g134268/U$3 ( \40773 , \40772 , \40387 );
nor \g134268/U$1 ( \40774 , \40771 , \40773 );
and \g135087/U$2 ( \40775 , \40175 , \40353 );
and \g135087/U$3 ( \40776 , \40307 , \40207 );
nor \g135087/U$1 ( \40777 , \40775 , \40776 );
and \g134310/U$2 ( \40778 , \40777 , \40137 );
not \g134310/U$4 ( \40779 , \40777 );
and \g134310/U$3 ( \40780 , \40779 , \40136 );
nor \g134310/U$1 ( \40781 , \40778 , \40780 );
xor \g133993/U$4 ( \40782 , \40774 , \40781 );
and \g134704/U$2 ( \40783 , \40147 , \40525 );
and \g134704/U$3 ( \40784 , \40472 , \40149 );
nor \g134704/U$1 ( \40785 , \40783 , \40784 );
and \g134620/U$2 ( \40786 , \40785 , \40107 );
not \g134620/U$4 ( \40787 , \40785 );
and \g134620/U$3 ( \40788 , \40787 , \40106 );
nor \g134620/U$1 ( \40789 , \40786 , \40788 );
and \g133993/U$3 ( \40790 , \40782 , \40789 );
and \g133993/U$5 ( \40791 , \40774 , \40781 );
or \g133993/U$2 ( \40792 , \40790 , \40791 );
and \g135020/U$2 ( \40793 , \40301 , \40278 );
and \g135020/U$3 ( \40794 , \40189 , \40391 );
nor \g135020/U$1 ( \40795 , \40793 , \40794 );
and \g134249/U$2 ( \40796 , \40795 , \40220 );
not \g134249/U$4 ( \40797 , \40795 );
and \g134249/U$3 ( \40798 , \40797 , \40219 );
nor \g134249/U$1 ( \40799 , \40796 , \40798 );
and \g135475/U$1 ( \40800 , \39910 , \39911 );
not \g135588/U$2 ( \40801 , \40800 );
nor \g135588/U$1 ( \40802 , \40801 , \40062 );
xor \g133996/U$4 ( \40803 , \40799 , \40802 );
and \g134860/U$2 ( \40804 , \40513 , \40108 );
and \g134860/U$3 ( \40805 , \40067 , \40713 );
nor \g134860/U$1 ( \40806 , \40804 , \40805 );
and \g134427/U$2 ( \40807 , \40806 , \40521 );
not \g134427/U$4 ( \40808 , \40806 );
and \g134427/U$3 ( \40809 , \40808 , \40518 );
nor \g134427/U$1 ( \40810 , \40807 , \40809 );
and \g133996/U$3 ( \40811 , \40803 , \40810 );
and \g133996/U$5 ( \40812 , \40799 , \40802 );
or \g133996/U$2 ( \40813 , \40811 , \40812 );
xor \g456206/U$5 ( \40814 , \40792 , \40813 );
xor \g133936/U$1 ( \40815 , \40710 , \40678 );
xor \g133936/U$1_r1 ( \40816 , \40815 , \40719 );
and \g456206/U$4 ( \40817 , \40814 , \40816 );
and \g456206/U$6 ( \40818 , \40792 , \40813 );
or \g456206/U$3 ( \40819 , \40817 , \40818 );
xor \g456191/U$5 ( \40820 , \40767 , \40819 );
xor \g456267/U$2 ( \40821 , \40567 , \40570 );
xor \g456267/U$1 ( \40822 , \40821 , \40578 );
xor \g456267/U$1_r1 ( \40823 , \40693 , \40698 );
xor \g456267/U$1_r2 ( \40824 , \40822 , \40823 );
and \g456191/U$4 ( \40825 , \40820 , \40824 );
and \g456191/U$6 ( \40826 , \40767 , \40819 );
or \g456191/U$3 ( \40827 , \40825 , \40826 );
xor \g456255/U$2 ( \40828 , \40588 , \40595 );
xor \g456255/U$1 ( \40829 , \40828 , \40603 );
xor \g456255/U$1_r1 ( \40830 , \40581 , \40621 );
xor \g456255/U$1_r2 ( \40831 , \40829 , \40830 );
xor \g133424/U$4 ( \40832 , \40827 , \40831 );
xor \g133565/U$1 ( \40833 , \40703 , \40747 );
xor \g133565/U$1_r1 ( \40834 , \40833 , \40750 );
and \g133424/U$3 ( \40835 , \40832 , \40834 );
and \g133424/U$5 ( \40836 , \40827 , \40831 );
or \g133424/U$2 ( \40837 , \40835 , \40836 );
and \g130256/U$2 ( \40838 , \40765 , \40837 );
xor \g133379/U$1 ( \40839 , \40837 , \40765 );
xor \g133424/U$1 ( \40840 , \40827 , \40831 );
xor \g133424/U$1_r1 ( \40841 , \40840 , \40834 );
not \g130319/U$3 ( \40842 , \40841 );
xor \g134047/U$1 ( \40843 , \40730 , \40733 );
xor \g134047/U$1_r1 ( \40844 , \40843 , \40741 );
xor \g456231/U$9 ( \40845 , \40663 , \40682 );
xor \g456231/U$9_r1 ( \40846 , \40845 , \40690 );
and \g456231/U$8 ( \40847 , \40844 , \40846 );
and \g134846/U$2 ( \40848 , \40091 , \40731 );
and \g134846/U$3 ( \40849 , \40568 , \40113 );
nor \g134846/U$1 ( \40850 , \40848 , \40849 );
and \g134191/U$2 ( \40851 , \40850 , \40080 );
not \g134191/U$4 ( \40852 , \40850 );
and \g134191/U$3 ( \40853 , \40852 , \40079 );
nor \g134191/U$1 ( \40854 , \40851 , \40853 );
not \g134649/U$1 ( \40855 , \40682 );
xor \g133786/U$4 ( \40856 , \40854 , \40855 );
and \g134808/U$2 ( \40857 , \40672 , \40067 );
not \g135286/U$1 ( \40858 , \40666 );
and \g134808/U$3 ( \40859 , \40064 , \40858 );
nor \g134808/U$1 ( \40860 , \40857 , \40859 );
and \g134357/U$2 ( \40861 , \40860 , \40678 );
not \g134357/U$4 ( \40862 , \40860 );
and \g134357/U$3 ( \40863 , \40862 , \40677 );
nor \g134357/U$1 ( \40864 , \40861 , \40863 );
xnor \g135425/U$1 ( \40865 , \32079 , \31835 );
not \g135243/U$3 ( \40866 , \40865 );
xnor \g135426/U$1 ( \40867 , \32566 , \32321 );
not \g135243/U$4 ( \40868 , \40867 );
and \g135243/U$2 ( \40869 , \40866 , \40868 );
nor \g135243/U$1 ( \40870 , \40869 , \40665 );
not \g135242/U$1 ( \40871 , \40870 );
xor \g133964/U$4 ( \40872 , \40864 , \40871 );
and \g134959/U$2 ( \40873 , \40432 , \40189 );
and \g134959/U$3 ( \40874 , \40138 , \40530 );
nor \g134959/U$1 ( \40875 , \40873 , \40874 );
and \g134585/U$2 ( \40876 , \40875 , \40388 );
not \g134585/U$4 ( \40877 , \40875 );
and \g134585/U$3 ( \40878 , \40877 , \40387 );
nor \g134585/U$1 ( \40879 , \40876 , \40878 );
and \g133964/U$3 ( \40880 , \40872 , \40879 );
and \g133964/U$5 ( \40881 , \40864 , \40871 );
or \g133964/U$2 ( \40882 , \40880 , \40881 );
and \g133786/U$3 ( \40883 , \40856 , \40882 );
and \g133786/U$5 ( \40884 , \40854 , \40855 );
or \g133786/U$2 ( \40885 , \40883 , \40884 );
xor \g456231/U$11 ( \40886 , \40663 , \40682 );
xor \g456231/U$11_r1 ( \40887 , \40886 , \40690 );
and \g456231/U$10 ( \40888 , \40885 , \40887 );
and \g456231/U$12 ( \40889 , \40844 , \40885 );
or \g456231/U$7 ( \40890 , \40847 , \40888 , \40889 );
xor \g456191/U$9 ( \40891 , \40767 , \40819 );
xor \g456191/U$9_r1 ( \40892 , \40891 , \40824 );
and \g456191/U$8 ( \40893 , \40890 , \40892 );
and \g135002/U$2 ( \40894 , \40513 , \40158 );
and \g135002/U$3 ( \40895 , \40108 , \40713 );
nor \g135002/U$1 ( \40896 , \40894 , \40895 );
and \g134421/U$2 ( \40897 , \40896 , \40521 );
not \g134421/U$4 ( \40898 , \40896 );
and \g134421/U$3 ( \40899 , \40898 , \40518 );
nor \g134421/U$1 ( \40900 , \40897 , \40899 );
and \g134886/U$2 ( \40901 , \40175 , \40472 );
and \g134886/U$3 ( \40902 , \40353 , \40207 );
nor \g134886/U$1 ( \40903 , \40901 , \40902 );
and \g134232/U$2 ( \40904 , \40903 , \40137 );
not \g134232/U$4 ( \40905 , \40903 );
and \g134232/U$3 ( \40906 , \40905 , \40136 );
nor \g134232/U$1 ( \40907 , \40904 , \40906 );
xor \g134008/U$4 ( \40908 , \40900 , \40907 );
and \g134827/U$2 ( \40909 , \40147 , \40568 );
and \g134827/U$3 ( \40910 , \40525 , \40149 );
nor \g134827/U$1 ( \40911 , \40909 , \40910 );
and \g134243/U$2 ( \40912 , \40911 , \40107 );
not \g134243/U$4 ( \40913 , \40911 );
and \g134243/U$3 ( \40914 , \40913 , \40106 );
nor \g134243/U$1 ( \40915 , \40912 , \40914 );
and \g134008/U$3 ( \40916 , \40908 , \40915 );
and \g134008/U$5 ( \40917 , \40900 , \40907 );
or \g134008/U$2 ( \40918 , \40916 , \40917 );
and \g134838/U$2 ( \40919 , \40091 , \40800 );
and \g134838/U$3 ( \40920 , \40731 , \40113 );
nor \g134838/U$1 ( \40921 , \40919 , \40920 );
and \g134302/U$2 ( \40922 , \40921 , \40080 );
not \g134302/U$4 ( \40923 , \40921 );
and \g134302/U$3 ( \40924 , \40923 , \40079 );
nor \g134302/U$1 ( \40925 , \40922 , \40924 );
and \g135504/U$1 ( \40926 , \39908 , \39909 );
not \g135601/U$2 ( \40927 , \40926 );
nor \g135601/U$1 ( \40928 , \40927 , \40062 );
xor \g133987/U$4 ( \40929 , \40925 , \40928 );
and \g134792/U$2 ( \40930 , \40301 , \40307 );
and \g134792/U$3 ( \40931 , \40278 , \40391 );
nor \g134792/U$1 ( \40932 , \40930 , \40931 );
and \g134539/U$2 ( \40933 , \40932 , \40220 );
not \g134539/U$4 ( \40934 , \40932 );
and \g134539/U$3 ( \40935 , \40934 , \40219 );
nor \g134539/U$1 ( \40936 , \40933 , \40935 );
and \g133987/U$3 ( \40937 , \40929 , \40936 );
and \g133987/U$5 ( \40938 , \40925 , \40928 );
or \g133987/U$2 ( \40939 , \40937 , \40938 );
xor \g133738/U$4 ( \40940 , \40918 , \40939 );
xor \g133993/U$1 ( \40941 , \40774 , \40781 );
xor \g133993/U$1_r1 ( \40942 , \40941 , \40789 );
and \g133738/U$3 ( \40943 , \40940 , \40942 );
and \g133738/U$5 ( \40944 , \40918 , \40939 );
or \g133738/U$2 ( \40945 , \40943 , \40944 );
xor \g456206/U$9 ( \40946 , \40792 , \40813 );
xor \g456206/U$9_r1 ( \40947 , \40946 , \40816 );
and \g456206/U$8 ( \40948 , \40945 , \40947 );
and \g134789/U$2 ( \40949 , \40091 , \40926 );
and \g134789/U$3 ( \40950 , \40800 , \40113 );
nor \g134789/U$1 ( \40951 , \40949 , \40950 );
and \g134177/U$2 ( \40952 , \40951 , \40080 );
not \g134177/U$4 ( \40953 , \40951 );
and \g134177/U$3 ( \40954 , \40953 , \40079 );
nor \g134177/U$1 ( \40955 , \40952 , \40954 );
and \g135478/U$1 ( \40956 , \39906 , \39907 );
not \g135589/U$2 ( \40957 , \40956 );
nor \g135589/U$1 ( \40958 , \40957 , \40062 );
xor \g133989/U$4 ( \40959 , \40955 , \40958 );
and \g134955/U$2 ( \40960 , \40432 , \40278 );
and \g134955/U$3 ( \40961 , \40189 , \40530 );
nor \g134955/U$1 ( \40962 , \40960 , \40961 );
and \g134293/U$2 ( \40963 , \40962 , \40388 );
not \g134293/U$4 ( \40964 , \40962 );
and \g134293/U$3 ( \40965 , \40964 , \40387 );
nor \g134293/U$1 ( \40966 , \40963 , \40965 );
and \g133989/U$3 ( \40967 , \40959 , \40966 );
and \g133989/U$5 ( \40968 , \40955 , \40958 );
or \g133989/U$2 ( \40969 , \40967 , \40968 );
not \g135424/U$1 ( \40970 , \40865 );
and \g135327/U$2 ( \40971 , \40867 , \40970 );
nor \g135386/U$1 ( \40972 , \40867 , \40970 );
nor \g135327/U$1 ( \40973 , \40971 , \40972 );
not \g135323/U$3 ( \40974 , \40867 );
not \g135323/U$4 ( \40975 , \40665 );
and \g135323/U$2 ( \40976 , \40974 , \40975 );
and \g135323/U$5 ( \40977 , \40665 , \40867 );
nor \g135323/U$1 ( \40978 , \40976 , \40977 );
and \g135236/U$1 ( \40979 , \40973 , \40978 );
nand \g135152/U$1 ( \40980 , \40064 , \40979 );
and \g134671/U$2 ( \40981 , \40980 , \40871 );
not \g134671/U$4 ( \40982 , \40980 );
and \g134671/U$3 ( \40983 , \40982 , \40870 );
nor \g134671/U$1 ( \40984 , \40981 , \40983 );
xor \g133798/U$4 ( \40985 , \40969 , \40984 );
and \g134924/U$2 ( \40986 , \40513 , \40138 );
and \g134924/U$3 ( \40987 , \40158 , \40713 );
nor \g134924/U$1 ( \40988 , \40986 , \40987 );
and \g134507/U$2 ( \40989 , \40988 , \40521 );
not \g134507/U$4 ( \40990 , \40988 );
and \g134507/U$3 ( \40991 , \40990 , \40518 );
nor \g134507/U$1 ( \40992 , \40989 , \40991 );
and \g134984/U$2 ( \40993 , \40672 , \40108 );
and \g134984/U$3 ( \40994 , \40067 , \40858 );
nor \g134984/U$1 ( \40995 , \40993 , \40994 );
and \g134231/U$2 ( \40996 , \40995 , \40678 );
not \g134231/U$4 ( \40997 , \40995 );
and \g134231/U$3 ( \40998 , \40997 , \40677 );
nor \g134231/U$1 ( \40999 , \40996 , \40998 );
xor \g134032/U$4 ( \41000 , \40992 , \40999 );
and \g134733/U$2 ( \41001 , \40301 , \40353 );
and \g134733/U$3 ( \41002 , \40307 , \40391 );
nor \g134733/U$1 ( \41003 , \41001 , \41002 );
and \g134156/U$2 ( \41004 , \41003 , \40220 );
not \g134156/U$4 ( \41005 , \41003 );
and \g134156/U$3 ( \41006 , \41005 , \40219 );
nor \g134156/U$1 ( \41007 , \41004 , \41006 );
and \g134032/U$3 ( \41008 , \41000 , \41007 );
and \g134032/U$5 ( \41009 , \40992 , \40999 );
or \g134032/U$2 ( \41010 , \41008 , \41009 );
and \g133798/U$3 ( \41011 , \40985 , \41010 );
and \g133798/U$5 ( \41012 , \40969 , \40984 );
or \g133798/U$2 ( \41013 , \41011 , \41012 );
xor \g133996/U$1 ( \41014 , \40799 , \40802 );
xor \g133996/U$1_r1 ( \41015 , \41014 , \40810 );
xor \g133609/U$4 ( \41016 , \41013 , \41015 );
xor \g133786/U$1 ( \41017 , \40854 , \40855 );
xor \g133786/U$1_r1 ( \41018 , \41017 , \40882 );
and \g133609/U$3 ( \41019 , \41016 , \41018 );
and \g133609/U$5 ( \41020 , \41013 , \41015 );
or \g133609/U$2 ( \41021 , \41019 , \41020 );
xor \g456206/U$11 ( \41022 , \40792 , \40813 );
xor \g456206/U$11_r1 ( \41023 , \41022 , \40816 );
and \g456206/U$10 ( \41024 , \41021 , \41023 );
and \g456206/U$12 ( \41025 , \40945 , \41021 );
or \g456206/U$7 ( \41026 , \40948 , \41024 , \41025 );
xor \g456191/U$11 ( \41027 , \40767 , \40819 );
xor \g456191/U$11_r1 ( \41028 , \41027 , \40824 );
and \g456191/U$10 ( \41029 , \41026 , \41028 );
and \g456191/U$12 ( \41030 , \40890 , \41026 );
or \g456191/U$7 ( \41031 , \40893 , \41029 , \41030 );
not \g130319/U$4 ( \41032 , \41031 );
or \g130319/U$2 ( \41033 , \40842 , \41032 );
xor \g456191/U$2 ( \41034 , \40767 , \40819 );
xor \g456191/U$1 ( \41035 , \41034 , \40824 );
xor \g456191/U$1_r1 ( \41036 , \40890 , \41026 );
xor \g456191/U$1_r2 ( \41037 , \41035 , \41036 );
xor \g133738/U$1 ( \41038 , \40918 , \40939 );
xor \g133738/U$1_r1 ( \41039 , \41038 , \40942 );
xor \g133964/U$1 ( \41040 , \40864 , \40871 );
xor \g133964/U$1_r1 ( \41041 , \41040 , \40879 );
xor \g134008/U$1 ( \41042 , \40900 , \40907 );
xor \g134008/U$1_r1 ( \41043 , \41042 , \40915 );
xor \g456204/U$5 ( \41044 , \41041 , \41043 );
xor \g133987/U$1 ( \41045 , \40925 , \40928 );
xor \g133987/U$1_r1 ( \41046 , \41045 , \40936 );
and \g456204/U$4 ( \41047 , \41044 , \41046 );
and \g456204/U$6 ( \41048 , \41041 , \41043 );
or \g456204/U$3 ( \41049 , \41047 , \41048 );
xor \g456190/U$5 ( \41050 , \41039 , \41049 );
xor \g133609/U$1 ( \41051 , \41013 , \41015 );
xor \g133609/U$1_r1 ( \41052 , \41051 , \41018 );
and \g456190/U$4 ( \41053 , \41050 , \41052 );
and \g456190/U$6 ( \41054 , \41039 , \41049 );
or \g456190/U$3 ( \41055 , \41053 , \41054 );
xor \g456231/U$2 ( \41056 , \40663 , \40682 );
xor \g456231/U$1 ( \41057 , \41056 , \40690 );
xor \g456231/U$1_r1 ( \41058 , \40844 , \40885 );
xor \g456231/U$1_r2 ( \41059 , \41057 , \41058 );
xor \g133383/U$4 ( \41060 , \41055 , \41059 );
xor \g456206/U$2 ( \41061 , \40792 , \40813 );
xor \g456206/U$1 ( \41062 , \41061 , \40816 );
xor \g456206/U$1_r1 ( \41063 , \40945 , \41021 );
xor \g456206/U$1_r2 ( \41064 , \41062 , \41063 );
and \g133383/U$3 ( \41065 , \41060 , \41064 );
and \g133383/U$5 ( \41066 , \41055 , \41059 );
or \g133383/U$2 ( \41067 , \41065 , \41066 );
and \g130400/U$2 ( \41068 , \41037 , \41067 );
xor \g133329/U$1 ( \41069 , \41067 , \41037 );
and \g134685/U$2 ( \41070 , \40979 , \40138 );
not \g135287/U$1 ( \41071 , \40973 );
and \g134685/U$3 ( \41072 , \40158 , \41071 );
nor \g134685/U$1 ( \41073 , \41070 , \41072 );
and \g134573/U$2 ( \41074 , \41073 , \40871 );
not \g134573/U$4 ( \41075 , \41073 );
and \g134573/U$3 ( \41076 , \41075 , \40870 );
nor \g134573/U$1 ( \41077 , \41074 , \41076 );
xnor \g135417/U$1 ( \41078 , \30625 , \30382 );
xnor \g135400/U$1 ( \41079 , \30137 , \29894 );
xnor \g455963/U$1 ( \41080 , \41078 , \41079 );
xnor \g135437/U$1 ( \41081 , \31108 , \30867 );
and \g135333/U$2 ( \41082 , \41078 , \41081 );
not \g135333/U$4 ( \41083 , \41078 );
not \g135436/U$1 ( \41084 , \41081 );
and \g135333/U$3 ( \41085 , \41083 , \41084 );
nor \g135333/U$1 ( \41086 , \41082 , \41085 );
and \g135230/U$1 ( \41087 , \41080 , \41086 );
nand \g135145/U$1 ( \41088 , \40064 , \41087 );
not \g135249/U$3 ( \41089 , \41079 );
not \g135249/U$4 ( \41090 , \41078 );
and \g135249/U$2 ( \41091 , \41089 , \41090 );
nor \g135249/U$1 ( \41092 , \41091 , \41081 );
not \g135248/U$1 ( \41093 , \41092 );
and \g134668/U$2 ( \41094 , \41088 , \41093 );
not \g134668/U$4 ( \41095 , \41088 );
and \g134668/U$3 ( \41096 , \41095 , \41092 );
nor \g134668/U$1 ( \41097 , \41094 , \41096 );
xor \g133984/U$1 ( \41098 , \41077 , \41097 );
and \g134774/U$2 ( \41099 , \40432 , \40525 );
and \g134774/U$3 ( \41100 , \40472 , \40530 );
nor \g134774/U$1 ( \41101 , \41099 , \41100 );
and \g134388/U$2 ( \41102 , \41101 , \40388 );
not \g134388/U$4 ( \41103 , \41101 );
and \g134388/U$3 ( \41104 , \41103 , \40387 );
nor \g134388/U$1 ( \41105 , \41102 , \41104 );
xor \g133984/U$1_r1 ( \41106 , \41098 , \41105 );
and \g135461/U$1 ( \41107 , \39900 , \39901 );
and \g135135/U$2 ( \41108 , \40091 , \41107 );
and \g135486/U$1 ( \41109 , \39902 , \39903 );
and \g135135/U$3 ( \41110 , \41109 , \40113 );
nor \g135135/U$1 ( \41111 , \41108 , \41110 );
and \g134332/U$2 ( \41112 , \41111 , \40080 );
not \g134332/U$4 ( \41113 , \41111 );
and \g134332/U$3 ( \41114 , \41113 , \40079 );
nor \g134332/U$1 ( \41115 , \41112 , \41114 );
and \g135494/U$1 ( \41116 , \39898 , \39899 );
not \g135596/U$2 ( \41117 , \41116 );
nor \g135596/U$1 ( \41118 , \41117 , \40062 );
xor \g456265/U$9 ( \41119 , \41115 , \41118 );
and \g134795/U$2 ( \41120 , \40513 , \40353 );
and \g134795/U$3 ( \41121 , \40307 , \40713 );
nor \g134795/U$1 ( \41122 , \41120 , \41121 );
and \g134514/U$2 ( \41123 , \41122 , \40521 );
not \g134514/U$4 ( \41124 , \41122 );
and \g134514/U$3 ( \41125 , \41124 , \40518 );
nor \g134514/U$1 ( \41126 , \41123 , \41125 );
xor \g456265/U$9_r1 ( \41127 , \41119 , \41126 );
and \g456265/U$8 ( \41128 , \41106 , \41127 );
and \g134822/U$2 ( \41129 , \40175 , \40926 );
and \g134822/U$3 ( \41130 , \40800 , \40207 );
nor \g134822/U$1 ( \41131 , \41129 , \41130 );
and \g134201/U$2 ( \41132 , \41131 , \40137 );
not \g134201/U$4 ( \41133 , \41131 );
and \g134201/U$3 ( \41134 , \41133 , \40136 );
nor \g134201/U$1 ( \41135 , \41132 , \41134 );
and \g134986/U$2 ( \41136 , \40672 , \40278 );
and \g134986/U$3 ( \41137 , \40189 , \40858 );
nor \g134986/U$1 ( \41138 , \41136 , \41137 );
and \g134254/U$2 ( \41139 , \41138 , \40678 );
not \g134254/U$4 ( \41140 , \41138 );
and \g134254/U$3 ( \41141 , \41140 , \40677 );
nor \g134254/U$1 ( \41142 , \41139 , \41141 );
xor \g134049/U$1 ( \41143 , \41135 , \41142 );
and \g135498/U$1 ( \41144 , \39904 , \39905 );
and \g134909/U$2 ( \41145 , \40147 , \41144 );
and \g134909/U$3 ( \41146 , \40956 , \40149 );
nor \g134909/U$1 ( \41147 , \41145 , \41146 );
and \g134316/U$2 ( \41148 , \41147 , \40107 );
not \g134316/U$4 ( \41149 , \41147 );
and \g134316/U$3 ( \41150 , \41149 , \40106 );
nor \g134316/U$1 ( \41151 , \41148 , \41150 );
xor \g134049/U$1_r1 ( \41152 , \41143 , \41151 );
xor \g456265/U$11 ( \41153 , \41115 , \41118 );
xor \g456265/U$11_r1 ( \41154 , \41153 , \41126 );
and \g456265/U$10 ( \41155 , \41152 , \41154 );
and \g456265/U$12 ( \41156 , \41106 , \41152 );
or \g456265/U$7 ( \41157 , \41128 , \41155 , \41156 );
xor \g134049/U$4 ( \41158 , \41135 , \41142 );
and \g134049/U$3 ( \41159 , \41158 , \41151 );
and \g134049/U$5 ( \41160 , \41135 , \41142 );
or \g134049/U$2 ( \41161 , \41159 , \41160 );
xor \g456265/U$5 ( \41162 , \41115 , \41118 );
and \g456265/U$4 ( \41163 , \41162 , \41126 );
and \g456265/U$6 ( \41164 , \41115 , \41118 );
or \g456265/U$3 ( \41165 , \41163 , \41164 );
xor \g456213/U$9 ( \41166 , \41161 , \41165 );
xor \g133984/U$4 ( \41167 , \41077 , \41097 );
and \g133984/U$3 ( \41168 , \41167 , \41105 );
and \g133984/U$5 ( \41169 , \41077 , \41097 );
or \g133984/U$2 ( \41170 , \41168 , \41169 );
xor \g456213/U$9_r1 ( \41171 , \41166 , \41170 );
and \g456213/U$8 ( \41172 , \41157 , \41171 );
and \g134697/U$2 ( \41173 , \40091 , \41109 );
and \g134697/U$3 ( \41174 , \41144 , \40113 );
nor \g134697/U$1 ( \41175 , \41173 , \41174 );
and \g134269/U$2 ( \41176 , \41175 , \40080 );
not \g134269/U$4 ( \41177 , \41175 );
and \g134269/U$3 ( \41178 , \41177 , \40079 );
nor \g134269/U$1 ( \41179 , \41176 , \41178 );
not \g135581/U$2 ( \41180 , \41107 );
nor \g135581/U$1 ( \41181 , \41180 , \40062 );
xor \g456262/U$2 ( \41182 , \41179 , \41181 );
and \g134865/U$2 ( \41183 , \40979 , \40158 );
and \g134865/U$3 ( \41184 , \40108 , \41071 );
nor \g134865/U$1 ( \41185 , \41183 , \41184 );
and \g134568/U$2 ( \41186 , \41185 , \40871 );
not \g134568/U$4 ( \41187 , \41185 );
and \g134568/U$3 ( \41188 , \41187 , \40870 );
nor \g134568/U$1 ( \41189 , \41186 , \41188 );
xor \g456262/U$1 ( \41190 , \41182 , \41189 );
and \g134710/U$2 ( \41191 , \40672 , \40189 );
and \g134710/U$3 ( \41192 , \40138 , \40858 );
nor \g134710/U$1 ( \41193 , \41191 , \41192 );
or \g134174/U$2 ( \41194 , \41193 , \40677 );
nand \g134632/U$1 ( \41195 , \40677 , \41193 );
nand \g134174/U$1 ( \41196 , \41194 , \41195 );
xor \g133933/U$1 ( \41197 , \41196 , \41093 );
xnor \g135416/U$1 ( \41198 , \31595 , \31351 );
and \g135332/U$2 ( \41199 , \41198 , \41084 );
nor \g135387/U$1 ( \41200 , \41198 , \41084 );
nor \g135332/U$1 ( \41201 , \41199 , \41200 );
and \g135335/U$2 ( \41202 , \41198 , \40865 );
not \g135335/U$4 ( \41203 , \41198 );
and \g135335/U$3 ( \41204 , \41203 , \40970 );
nor \g135335/U$1 ( \41205 , \41202 , \41204 );
and \g135223/U$1 ( \41206 , \41201 , \41205 );
and \g135122/U$2 ( \41207 , \41206 , \40067 );
not \g135274/U$1 ( \41208 , \41201 );
and \g135122/U$3 ( \41209 , \40064 , \41208 );
nor \g135122/U$1 ( \41210 , \41207 , \41209 );
not \g135245/U$3 ( \41211 , \41081 );
not \g135245/U$4 ( \41212 , \41198 );
and \g135245/U$2 ( \41213 , \41211 , \41212 );
nor \g135245/U$1 ( \41214 , \41213 , \40865 );
not \g135244/U$1 ( \41215 , \41214 );
and \g134386/U$2 ( \41216 , \41210 , \41215 );
not \g134386/U$4 ( \41217 , \41210 );
and \g134386/U$3 ( \41218 , \41217 , \41214 );
nor \g134386/U$1 ( \41219 , \41216 , \41218 );
xor \g133933/U$1_r1 ( \41220 , \41197 , \41219 );
and \g134825/U$2 ( \41221 , \40175 , \40800 );
and \g134825/U$3 ( \41222 , \40731 , \40207 );
nor \g134825/U$1 ( \41223 , \41221 , \41222 );
and \g134400/U$2 ( \41224 , \41223 , \40137 );
not \g134400/U$4 ( \41225 , \41223 );
and \g134400/U$3 ( \41226 , \41225 , \40136 );
nor \g134400/U$1 ( \41227 , \41224 , \41226 );
and \g134807/U$2 ( \41228 , \40513 , \40307 );
and \g134807/U$3 ( \41229 , \40278 , \40713 );
nor \g134807/U$1 ( \41230 , \41228 , \41229 );
and \g134158/U$2 ( \41231 , \41230 , \40521 );
not \g134158/U$4 ( \41232 , \41230 );
and \g134158/U$3 ( \41233 , \41232 , \40518 );
nor \g134158/U$1 ( \41234 , \41231 , \41233 );
xor \g134046/U$1 ( \41235 , \41227 , \41234 );
and \g134854/U$2 ( \41236 , \40147 , \40956 );
and \g134854/U$3 ( \41237 , \40926 , \40149 );
nor \g134854/U$1 ( \41238 , \41236 , \41237 );
and \g134591/U$2 ( \41239 , \41238 , \40107 );
not \g134591/U$4 ( \41240 , \41238 );
and \g134591/U$3 ( \41241 , \41240 , \40106 );
nor \g134591/U$1 ( \41242 , \41239 , \41241 );
xor \g134046/U$1_r1 ( \41243 , \41235 , \41242 );
xor \g456262/U$1_r1 ( \41244 , \41220 , \41243 );
xor \g456262/U$1_r2 ( \41245 , \41190 , \41244 );
xor \g456213/U$11 ( \41246 , \41161 , \41165 );
xor \g456213/U$11_r1 ( \41247 , \41246 , \41170 );
and \g456213/U$10 ( \41248 , \41245 , \41247 );
and \g456213/U$12 ( \41249 , \41157 , \41245 );
or \g456213/U$7 ( \41250 , \41172 , \41248 , \41249 );
and \g135001/U$2 ( \41251 , \41206 , \40108 );
and \g135001/U$3 ( \41252 , \40067 , \41208 );
nor \g135001/U$1 ( \41253 , \41251 , \41252 );
and \g134548/U$2 ( \41254 , \41253 , \41214 );
not \g134548/U$4 ( \41255 , \41253 );
and \g134548/U$3 ( \41256 , \41255 , \41215 );
nor \g134548/U$1 ( \41257 , \41254 , \41256 );
and \g134752/U$2 ( \41258 , \40301 , \40731 );
and \g134752/U$3 ( \41259 , \40568 , \40391 );
nor \g134752/U$1 ( \41260 , \41258 , \41259 );
and \g134221/U$2 ( \41261 , \41260 , \40220 );
not \g134221/U$4 ( \41262 , \41260 );
and \g134221/U$3 ( \41263 , \41262 , \40219 );
nor \g134221/U$1 ( \41264 , \41261 , \41263 );
xor \g133801/U$4 ( \41265 , \41257 , \41264 );
and \g134839/U$2 ( \41266 , \41206 , \40158 );
and \g134839/U$3 ( \41267 , \40108 , \41208 );
nor \g134839/U$1 ( \41268 , \41266 , \41267 );
and \g134521/U$2 ( \41269 , \41268 , \41215 );
not \g134521/U$4 ( \41270 , \41268 );
and \g134521/U$3 ( \41271 , \41270 , \41214 );
nor \g134521/U$1 ( \41272 , \41269 , \41271 );
and \g135037/U$2 ( \41273 , \40147 , \41109 );
and \g135037/U$3 ( \41274 , \41144 , \40149 );
nor \g135037/U$1 ( \41275 , \41273 , \41274 );
and \g134237/U$2 ( \41276 , \41275 , \40107 );
not \g134237/U$4 ( \41277 , \41275 );
and \g134237/U$3 ( \41278 , \41277 , \40106 );
nor \g134237/U$1 ( \41279 , \41276 , \41278 );
xor \g133992/U$4 ( \41280 , \41272 , \41279 );
and \g135024/U$2 ( \41281 , \40091 , \41116 );
and \g135024/U$3 ( \41282 , \41107 , \40113 );
nor \g135024/U$1 ( \41283 , \41281 , \41282 );
and \g134235/U$2 ( \41284 , \41283 , \40080 );
not \g134235/U$4 ( \41285 , \41283 );
and \g134235/U$3 ( \41286 , \41285 , \40079 );
nor \g134235/U$1 ( \41287 , \41284 , \41286 );
and \g133992/U$3 ( \41288 , \41280 , \41287 );
and \g133992/U$5 ( \41289 , \41272 , \41279 );
or \g133992/U$2 ( \41290 , \41288 , \41289 );
and \g133801/U$3 ( \41291 , \41265 , \41290 );
and \g133801/U$5 ( \41292 , \41257 , \41264 );
or \g133801/U$2 ( \41293 , \41291 , \41292 );
and \g134856/U$2 ( \41294 , \40301 , \40568 );
and \g134856/U$3 ( \41295 , \40525 , \40391 );
nor \g134856/U$1 ( \41296 , \41294 , \41295 );
and \g134619/U$2 ( \41297 , \41296 , \40220 );
not \g134619/U$4 ( \41298 , \41296 );
and \g134619/U$3 ( \41299 , \41298 , \40219 );
nor \g134619/U$1 ( \41300 , \41297 , \41299 );
and \g135066/U$2 ( \41301 , \40432 , \40472 );
and \g135066/U$3 ( \41302 , \40353 , \40530 );
nor \g135066/U$1 ( \41303 , \41301 , \41302 );
and \g134464/U$2 ( \41304 , \41303 , \40388 );
not \g134464/U$4 ( \41305 , \41303 );
and \g134464/U$3 ( \41306 , \41305 , \40387 );
nor \g134464/U$1 ( \41307 , \41304 , \41306 );
xor \g133982/U$1 ( \41308 , \41300 , \41307 );
not \g134547/U$1 ( \41309 , \41257 );
xor \g133982/U$1_r1 ( \41310 , \41308 , \41309 );
xor \g456194/U$5 ( \41311 , \41293 , \41310 );
and \g135050/U$2 ( \41312 , \40979 , \40189 );
and \g135050/U$3 ( \41313 , \40138 , \41071 );
nor \g135050/U$1 ( \41314 , \41312 , \41313 );
and \g134383/U$2 ( \41315 , \41314 , \40871 );
not \g134383/U$4 ( \41316 , \41314 );
and \g134383/U$3 ( \41317 , \41316 , \40870 );
nor \g134383/U$1 ( \41318 , \41315 , \41317 );
xnor \g135405/U$1 ( \41319 , \29170 , \28925 );
not \g135265/U$3 ( \41320 , \41319 );
xnor \g135438/U$1 ( \41321 , \29653 , \29411 );
not \g135265/U$4 ( \41322 , \41321 );
and \g135265/U$2 ( \41323 , \41320 , \41322 );
nor \g135265/U$1 ( \41324 , \41323 , \41079 );
not \g135264/U$1 ( \41325 , \41324 );
xor \g133921/U$4 ( \41326 , \41318 , \41325 );
and \g134779/U$2 ( \41327 , \41087 , \40067 );
not \g135272/U$1 ( \41328 , \41080 );
and \g134779/U$3 ( \41329 , \40064 , \41328 );
nor \g134779/U$1 ( \41330 , \41327 , \41329 );
and \g134558/U$2 ( \41331 , \41330 , \41093 );
not \g134558/U$4 ( \41332 , \41330 );
and \g134558/U$3 ( \41333 , \41332 , \41092 );
nor \g134558/U$1 ( \41334 , \41331 , \41333 );
and \g133921/U$3 ( \41335 , \41326 , \41334 );
and \g133921/U$5 ( \41336 , \41318 , \41325 );
or \g133921/U$2 ( \41337 , \41335 , \41336 );
and \g134731/U$2 ( \41338 , \40513 , \40472 );
and \g134731/U$3 ( \41339 , \40353 , \40713 );
nor \g134731/U$1 ( \41340 , \41338 , \41339 );
and \g134522/U$2 ( \41341 , \41340 , \40521 );
not \g134522/U$4 ( \41342 , \41340 );
and \g134522/U$3 ( \41343 , \41342 , \40518 );
nor \g134522/U$1 ( \41344 , \41341 , \41343 );
and \g135445/U$1 ( \41345 , \39896 , \39897 );
not \g135573/U$2 ( \41346 , \41345 );
nor \g135573/U$1 ( \41347 , \41346 , \40062 );
xor \g456240/U$5 ( \41348 , \41344 , \41347 );
and \g134768/U$2 ( \41349 , \40432 , \40568 );
and \g134768/U$3 ( \41350 , \40525 , \40530 );
nor \g134768/U$1 ( \41351 , \41349 , \41350 );
and \g134274/U$2 ( \41352 , \41351 , \40388 );
not \g134274/U$4 ( \41353 , \41351 );
and \g134274/U$3 ( \41354 , \41353 , \40387 );
nor \g134274/U$1 ( \41355 , \41352 , \41354 );
and \g456240/U$4 ( \41356 , \41348 , \41355 );
and \g456240/U$6 ( \41357 , \41344 , \41347 );
or \g456240/U$3 ( \41358 , \41356 , \41357 );
xor \g133677/U$4 ( \41359 , \41337 , \41358 );
and \g134711/U$2 ( \41360 , \40175 , \40956 );
and \g134711/U$3 ( \41361 , \40926 , \40207 );
nor \g134711/U$1 ( \41362 , \41360 , \41361 );
and \g134207/U$2 ( \41363 , \41362 , \40137 );
not \g134207/U$4 ( \41364 , \41362 );
and \g134207/U$3 ( \41365 , \41364 , \40136 );
nor \g134207/U$1 ( \41366 , \41363 , \41365 );
and \g135046/U$2 ( \41367 , \40672 , \40307 );
and \g135046/U$3 ( \41368 , \40278 , \40858 );
nor \g135046/U$1 ( \41369 , \41367 , \41368 );
and \g134264/U$2 ( \41370 , \41369 , \40678 );
not \g134264/U$4 ( \41371 , \41369 );
and \g134264/U$3 ( \41372 , \41371 , \40677 );
nor \g134264/U$1 ( \41373 , \41370 , \41372 );
xor \g133888/U$4 ( \41374 , \41366 , \41373 );
and \g135058/U$2 ( \41375 , \40301 , \40800 );
and \g135058/U$3 ( \41376 , \40731 , \40391 );
nor \g135058/U$1 ( \41377 , \41375 , \41376 );
and \g134362/U$2 ( \41378 , \41377 , \40220 );
not \g134362/U$4 ( \41379 , \41377 );
and \g134362/U$3 ( \41380 , \41379 , \40219 );
nor \g134362/U$1 ( \41381 , \41378 , \41380 );
and \g133888/U$3 ( \41382 , \41374 , \41381 );
and \g133888/U$5 ( \41383 , \41366 , \41373 );
or \g133888/U$2 ( \41384 , \41382 , \41383 );
and \g133677/U$3 ( \41385 , \41359 , \41384 );
and \g133677/U$5 ( \41386 , \41337 , \41358 );
or \g133677/U$2 ( \41387 , \41385 , \41386 );
and \g456194/U$4 ( \41388 , \41311 , \41387 );
and \g456194/U$6 ( \41389 , \41293 , \41310 );
or \g456194/U$3 ( \41390 , \41388 , \41389 );
xor \g133414/U$4 ( \41391 , \41250 , \41390 );
and \g134900/U$2 ( \41392 , \40175 , \40731 );
and \g134900/U$3 ( \41393 , \40568 , \40207 );
nor \g134900/U$1 ( \41394 , \41392 , \41393 );
and \g134463/U$2 ( \41395 , \41394 , \40137 );
not \g134463/U$4 ( \41396 , \41394 );
and \g134463/U$3 ( \41397 , \41396 , \40136 );
nor \g134463/U$1 ( \41398 , \41395 , \41397 );
and \g134681/U$2 ( \41399 , \40672 , \40138 );
and \g134681/U$3 ( \41400 , \40158 , \40858 );
nor \g134681/U$1 ( \41401 , \41399 , \41400 );
and \g134618/U$2 ( \41402 , \41401 , \40678 );
not \g134618/U$4 ( \41403 , \41401 );
and \g134618/U$3 ( \41404 , \41403 , \40677 );
nor \g134618/U$1 ( \41405 , \41402 , \41404 );
xor \g456221/U$2 ( \41406 , \41398 , \41405 );
and \g134814/U$2 ( \41407 , \40301 , \40525 );
and \g134814/U$3 ( \41408 , \40472 , \40391 );
nor \g134814/U$1 ( \41409 , \41407 , \41408 );
and \g134417/U$2 ( \41410 , \41409 , \40220 );
not \g134417/U$4 ( \41411 , \41409 );
and \g134417/U$3 ( \41412 , \41411 , \40219 );
nor \g134417/U$1 ( \41413 , \41410 , \41412 );
xor \g456221/U$1 ( \41414 , \41406 , \41413 );
xor \g133982/U$4 ( \41415 , \41300 , \41307 );
and \g133982/U$3 ( \41416 , \41415 , \41309 );
and \g133982/U$5 ( \41417 , \41300 , \41307 );
or \g133982/U$2 ( \41418 , \41416 , \41417 );
xor \g456213/U$5 ( \41419 , \41161 , \41165 );
and \g456213/U$4 ( \41420 , \41419 , \41170 );
and \g456213/U$6 ( \41421 , \41161 , \41165 );
or \g456213/U$3 ( \41422 , \41420 , \41421 );
xor \g456221/U$1_r1 ( \41423 , \41418 , \41422 );
xor \g456221/U$1_r2 ( \41424 , \41414 , \41423 );
and \g133414/U$3 ( \41425 , \41391 , \41424 );
and \g133414/U$5 ( \41426 , \41250 , \41390 );
or \g133414/U$2 ( \41427 , \41425 , \41426 );
xor \g456262/U$5 ( \41428 , \41179 , \41181 );
and \g456262/U$4 ( \41429 , \41428 , \41189 );
and \g456262/U$6 ( \41430 , \41179 , \41181 );
or \g456262/U$3 ( \41431 , \41429 , \41430 );
and \g135042/U$2 ( \41432 , \40432 , \40353 );
and \g135042/U$3 ( \41433 , \40307 , \40530 );
nor \g135042/U$1 ( \41434 , \41432 , \41433 );
or \g134165/U$2 ( \41435 , \41434 , \40387 );
nand \g134631/U$1 ( \41436 , \40387 , \41434 );
nand \g134165/U$1 ( \41437 , \41435 , \41436 );
not \g135593/U$2 ( \41438 , \41109 );
nor \g135593/U$1 ( \41439 , \41438 , \40062 );
xor \g456268/U$9 ( \41440 , \41437 , \41439 );
and \g134892/U$2 ( \41441 , \40979 , \40108 );
and \g134892/U$3 ( \41442 , \40067 , \41071 );
nor \g134892/U$1 ( \41443 , \41441 , \41442 );
and \g134579/U$2 ( \41444 , \41443 , \40871 );
not \g134579/U$4 ( \41445 , \41443 );
and \g134579/U$3 ( \41446 , \41445 , \40870 );
nor \g134579/U$1 ( \41447 , \41444 , \41446 );
xor \g456268/U$9_r1 ( \41448 , \41440 , \41447 );
and \g456268/U$8 ( \41449 , \41431 , \41448 );
and \g135084/U$2 ( \41450 , \40091 , \41144 );
and \g135084/U$3 ( \41451 , \40956 , \40113 );
nor \g135084/U$1 ( \41452 , \41450 , \41451 );
and \g134394/U$2 ( \41453 , \41452 , \40080 );
not \g134394/U$4 ( \41454 , \41452 );
and \g134394/U$3 ( \41455 , \41454 , \40079 );
nor \g134394/U$1 ( \41456 , \41453 , \41455 );
and \g134990/U$2 ( \41457 , \40513 , \40278 );
and \g134990/U$3 ( \41458 , \40189 , \40713 );
nor \g134990/U$1 ( \41459 , \41457 , \41458 );
and \g134553/U$2 ( \41460 , \41459 , \40521 );
not \g134553/U$4 ( \41461 , \41459 );
and \g134553/U$3 ( \41462 , \41461 , \40518 );
nor \g134553/U$1 ( \41463 , \41460 , \41462 );
xor \g133899/U$1 ( \41464 , \41456 , \41463 );
and \g134884/U$2 ( \41465 , \40147 , \40926 );
and \g134884/U$3 ( \41466 , \40800 , \40149 );
nor \g134884/U$1 ( \41467 , \41465 , \41466 );
and \g134377/U$2 ( \41468 , \41467 , \40107 );
not \g134377/U$4 ( \41469 , \41467 );
and \g134377/U$3 ( \41470 , \41469 , \40106 );
nor \g134377/U$1 ( \41471 , \41468 , \41470 );
xor \g133899/U$1_r1 ( \41472 , \41464 , \41471 );
xor \g456268/U$11 ( \41473 , \41437 , \41439 );
xor \g456268/U$11_r1 ( \41474 , \41473 , \41447 );
and \g456268/U$10 ( \41475 , \41472 , \41474 );
and \g456268/U$12 ( \41476 , \41431 , \41472 );
or \g456268/U$7 ( \41477 , \41449 , \41475 , \41476 );
xor \g133933/U$4 ( \41478 , \41196 , \41093 );
and \g133933/U$3 ( \41479 , \41478 , \41219 );
and \g133933/U$5 ( \41480 , \41196 , \41093 );
or \g133933/U$2 ( \41481 , \41479 , \41480 );
nand \g135154/U$1 ( \41482 , \40064 , \41206 );
and \g134657/U$2 ( \41483 , \41482 , \41215 );
not \g134657/U$4 ( \41484 , \41482 );
and \g134657/U$3 ( \41485 , \41484 , \41214 );
nor \g134657/U$1 ( \41486 , \41483 , \41485 );
not \g134656/U$1 ( \41487 , \41486 );
xor \g456217/U$5 ( \41488 , \41481 , \41487 );
xor \g134046/U$4 ( \41489 , \41227 , \41234 );
and \g134046/U$3 ( \41490 , \41489 , \41242 );
and \g134046/U$5 ( \41491 , \41227 , \41234 );
or \g134046/U$2 ( \41492 , \41490 , \41491 );
and \g456217/U$4 ( \41493 , \41488 , \41492 );
and \g456217/U$6 ( \41494 , \41481 , \41487 );
or \g456217/U$3 ( \41495 , \41493 , \41494 );
xor \g133586/U$1 ( \41496 , \41477 , \41495 );
xor \g456221/U$5 ( \41497 , \41398 , \41405 );
and \g456221/U$4 ( \41498 , \41497 , \41413 );
and \g456221/U$6 ( \41499 , \41398 , \41405 );
or \g456221/U$3 ( \41500 , \41498 , \41499 );
xor \g456268/U$5 ( \41501 , \41437 , \41439 );
and \g456268/U$4 ( \41502 , \41501 , \41447 );
and \g456268/U$6 ( \41503 , \41437 , \41439 );
or \g456268/U$3 ( \41504 , \41502 , \41503 );
xor \g133710/U$1 ( \41505 , \41500 , \41504 );
and \g134938/U$2 ( \41506 , \40672 , \40158 );
and \g134938/U$3 ( \41507 , \40108 , \40858 );
nor \g134938/U$1 ( \41508 , \41506 , \41507 );
and \g134530/U$2 ( \41509 , \41508 , \40678 );
not \g134530/U$4 ( \41510 , \41508 );
and \g134530/U$3 ( \41511 , \41510 , \40677 );
nor \g134530/U$1 ( \41512 , \41509 , \41511 );
not \g135598/U$2 ( \41513 , \41144 );
nor \g135598/U$1 ( \41514 , \41513 , \40062 );
xor \g133991/U$1 ( \41515 , \41512 , \41514 );
and \g134730/U$2 ( \41516 , \40301 , \40472 );
and \g134730/U$3 ( \41517 , \40353 , \40391 );
nor \g134730/U$1 ( \41518 , \41516 , \41517 );
and \g134339/U$2 ( \41519 , \41518 , \40220 );
not \g134339/U$4 ( \41520 , \41518 );
and \g134339/U$3 ( \41521 , \41520 , \40219 );
nor \g134339/U$1 ( \41522 , \41519 , \41521 );
xor \g133991/U$1_r1 ( \41523 , \41515 , \41522 );
xor \g133710/U$1_r1 ( \41524 , \41505 , \41523 );
xor \g133586/U$1_r1 ( \41525 , \41496 , \41524 );
xor \g133301/U$1 ( \41526 , \41427 , \41525 );
and \g134917/U$2 ( \41527 , \40432 , \40307 );
and \g134917/U$3 ( \41528 , \40278 , \40530 );
nor \g134917/U$1 ( \41529 , \41527 , \41528 );
and \g134343/U$2 ( \41530 , \41529 , \40388 );
not \g134343/U$4 ( \41531 , \41529 );
and \g134343/U$3 ( \41532 , \41531 , \40387 );
nor \g134343/U$1 ( \41533 , \41530 , \41532 );
and \g134851/U$2 ( \41534 , \40147 , \40800 );
and \g134851/U$3 ( \41535 , \40731 , \40149 );
nor \g134851/U$1 ( \41536 , \41534 , \41535 );
and \g134229/U$2 ( \41537 , \41536 , \40107 );
not \g134229/U$4 ( \41538 , \41536 );
and \g134229/U$3 ( \41539 , \41538 , \40106 );
nor \g134229/U$1 ( \41540 , \41537 , \41539 );
xor \g134004/U$1 ( \41541 , \41533 , \41540 );
and \g135083/U$2 ( \41542 , \40091 , \40956 );
and \g135083/U$3 ( \41543 , \40926 , \40113 );
nor \g135083/U$1 ( \41544 , \41542 , \41543 );
and \g134555/U$2 ( \41545 , \41544 , \40080 );
not \g134555/U$4 ( \41546 , \41544 );
and \g134555/U$3 ( \41547 , \41546 , \40079 );
nor \g134555/U$1 ( \41548 , \41545 , \41547 );
xor \g134004/U$1_r1 ( \41549 , \41541 , \41548 );
and \g134746/U$2 ( \41550 , \40513 , \40189 );
and \g134746/U$3 ( \41551 , \40138 , \40713 );
nor \g134746/U$1 ( \41552 , \41550 , \41551 );
and \g134371/U$2 ( \41553 , \41552 , \40521 );
not \g134371/U$4 ( \41554 , \41552 );
and \g134371/U$3 ( \41555 , \41554 , \40518 );
nor \g134371/U$1 ( \41556 , \41553 , \41555 );
xor \g133937/U$1 ( \41557 , \41556 , \41215 );
and \g135056/U$2 ( \41558 , \40979 , \40067 );
and \g135056/U$3 ( \41559 , \40064 , \41071 );
nor \g135056/U$1 ( \41560 , \41558 , \41559 );
and \g134488/U$2 ( \41561 , \41560 , \40871 );
not \g134488/U$4 ( \41562 , \41560 );
and \g134488/U$3 ( \41563 , \41562 , \40870 );
nor \g134488/U$1 ( \41564 , \41561 , \41563 );
xor \g133937/U$1_r1 ( \41565 , \41557 , \41564 );
xor \g456198/U$2 ( \41566 , \41549 , \41565 );
and \g134742/U$2 ( \41567 , \40175 , \40568 );
and \g134742/U$3 ( \41568 , \40525 , \40207 );
nor \g134742/U$1 ( \41569 , \41567 , \41568 );
and \g134299/U$2 ( \41570 , \41569 , \40137 );
not \g134299/U$4 ( \41571 , \41569 );
and \g134299/U$3 ( \41572 , \41571 , \40136 );
nor \g134299/U$1 ( \41573 , \41570 , \41572 );
xor \g133727/U$1 ( \41574 , \41573 , \41486 );
xor \g133899/U$4 ( \41575 , \41456 , \41463 );
and \g133899/U$3 ( \41576 , \41575 , \41471 );
and \g133899/U$5 ( \41577 , \41456 , \41463 );
or \g133899/U$2 ( \41578 , \41576 , \41577 );
xor \g133727/U$1_r1 ( \41579 , \41574 , \41578 );
xor \g456198/U$1 ( \41580 , \41566 , \41579 );
xor \g456221/U$9 ( \41581 , \41398 , \41405 );
xor \g456221/U$9_r1 ( \41582 , \41581 , \41413 );
and \g456221/U$8 ( \41583 , \41418 , \41582 );
xor \g456221/U$11 ( \41584 , \41398 , \41405 );
xor \g456221/U$11_r1 ( \41585 , \41584 , \41413 );
and \g456221/U$10 ( \41586 , \41422 , \41585 );
and \g456221/U$12 ( \41587 , \41418 , \41422 );
or \g456221/U$7 ( \41588 , \41583 , \41586 , \41587 );
xor \g456262/U$9 ( \41589 , \41179 , \41181 );
xor \g456262/U$9_r1 ( \41590 , \41589 , \41189 );
and \g456262/U$8 ( \41591 , \41220 , \41590 );
xor \g456262/U$11 ( \41592 , \41179 , \41181 );
xor \g456262/U$11_r1 ( \41593 , \41592 , \41189 );
and \g456262/U$10 ( \41594 , \41243 , \41593 );
and \g456262/U$12 ( \41595 , \41220 , \41243 );
or \g456262/U$7 ( \41596 , \41591 , \41594 , \41595 );
xor \g456217/U$9 ( \41597 , \41481 , \41487 );
xor \g456217/U$9_r1 ( \41598 , \41597 , \41492 );
and \g456217/U$8 ( \41599 , \41596 , \41598 );
xor \g456268/U$2 ( \41600 , \41437 , \41439 );
xor \g456268/U$1 ( \41601 , \41600 , \41447 );
xor \g456268/U$1_r1 ( \41602 , \41431 , \41472 );
xor \g456268/U$1_r2 ( \41603 , \41601 , \41602 );
xor \g456217/U$11 ( \41604 , \41481 , \41487 );
xor \g456217/U$11_r1 ( \41605 , \41604 , \41492 );
and \g456217/U$10 ( \41606 , \41603 , \41605 );
and \g456217/U$12 ( \41607 , \41596 , \41603 );
or \g456217/U$7 ( \41608 , \41599 , \41606 , \41607 );
xor \g456198/U$1_r1 ( \41609 , \41588 , \41608 );
xor \g456198/U$1_r2 ( \41610 , \41580 , \41609 );
xor \g133301/U$1_r1 ( \41611 , \41526 , \41610 );
xor \g133801/U$1 ( \41612 , \41257 , \41264 );
xor \g133801/U$1_r1 ( \41613 , \41612 , \41290 );
not \g135404/U$1 ( \41614 , \41319 );
and \g135324/U$2 ( \41615 , \41321 , \41614 );
nor \g135385/U$1 ( \41616 , \41321 , \41614 );
nor \g135324/U$1 ( \41617 , \41615 , \41616 );
not \g135320/U$3 ( \41618 , \41321 );
not \g135320/U$4 ( \41619 , \41079 );
and \g135320/U$2 ( \41620 , \41618 , \41619 );
and \g135320/U$5 ( \41621 , \41079 , \41321 );
nor \g135320/U$1 ( \41622 , \41620 , \41621 );
and \g135237/U$1 ( \41623 , \41617 , \41622 );
nand \g135150/U$1 ( \41624 , \40064 , \41623 );
and \g134661/U$2 ( \41625 , \41624 , \41325 );
not \g134661/U$4 ( \41626 , \41624 );
and \g134661/U$3 ( \41627 , \41626 , \41324 );
nor \g134661/U$1 ( \41628 , \41625 , \41627 );
and \g135469/U$1 ( \41629 , \39894 , \39895 );
not \g135585/U$2 ( \41630 , \41629 );
nor \g135585/U$1 ( \41631 , \41630 , \40062 );
xor \g134021/U$4 ( \41632 , \41628 , \41631 );
and \g135128/U$2 ( \41633 , \41206 , \40138 );
and \g135128/U$3 ( \41634 , \40158 , \41208 );
nor \g135128/U$1 ( \41635 , \41633 , \41634 );
and \g134551/U$2 ( \41636 , \41635 , \41215 );
not \g134551/U$4 ( \41637 , \41635 );
and \g134551/U$3 ( \41638 , \41637 , \41214 );
nor \g134551/U$1 ( \41639 , \41636 , \41638 );
and \g134021/U$3 ( \41640 , \41632 , \41639 );
and \g134021/U$5 ( \41641 , \41628 , \41631 );
or \g134021/U$2 ( \41642 , \41640 , \41641 );
and \g135038/U$2 ( \41643 , \41087 , \40108 );
and \g135038/U$3 ( \41644 , \40067 , \41328 );
nor \g135038/U$1 ( \41645 , \41643 , \41644 );
and \g134510/U$2 ( \41646 , \41645 , \41093 );
not \g134510/U$4 ( \41647 , \41645 );
and \g134510/U$3 ( \41648 , \41647 , \41092 );
nor \g134510/U$1 ( \41649 , \41646 , \41648 );
xor \g133777/U$4 ( \41650 , \41642 , \41649 );
and \g135015/U$2 ( \41651 , \40979 , \40278 );
and \g135015/U$3 ( \41652 , \40189 , \41071 );
nor \g135015/U$1 ( \41653 , \41651 , \41652 );
and \g134272/U$2 ( \41654 , \41653 , \40871 );
not \g134272/U$4 ( \41655 , \41653 );
and \g134272/U$3 ( \41656 , \41655 , \40870 );
nor \g134272/U$1 ( \41657 , \41654 , \41656 );
and \g134686/U$2 ( \41658 , \40301 , \40926 );
and \g134686/U$3 ( \41659 , \40800 , \40391 );
nor \g134686/U$1 ( \41660 , \41658 , \41659 );
and \g134508/U$2 ( \41661 , \41660 , \40220 );
not \g134508/U$4 ( \41662 , \41660 );
and \g134508/U$3 ( \41663 , \41662 , \40219 );
nor \g134508/U$1 ( \41664 , \41661 , \41663 );
xor \g456242/U$5 ( \41665 , \41657 , \41664 );
and \g135044/U$2 ( \41666 , \40175 , \41144 );
and \g135044/U$3 ( \41667 , \40956 , \40207 );
nor \g135044/U$1 ( \41668 , \41666 , \41667 );
and \g134297/U$2 ( \41669 , \41668 , \40137 );
not \g134297/U$4 ( \41670 , \41668 );
and \g134297/U$3 ( \41671 , \41670 , \40136 );
nor \g134297/U$1 ( \41672 , \41669 , \41671 );
and \g456242/U$4 ( \41673 , \41665 , \41672 );
and \g456242/U$6 ( \41674 , \41657 , \41664 );
or \g456242/U$3 ( \41675 , \41673 , \41674 );
and \g133777/U$3 ( \41676 , \41650 , \41675 );
and \g133777/U$5 ( \41677 , \41642 , \41649 );
or \g133777/U$2 ( \41678 , \41676 , \41677 );
xor \g456184/U$5 ( \41679 , \41613 , \41678 );
xor \g133677/U$1 ( \41680 , \41337 , \41358 );
xor \g133677/U$1_r1 ( \41681 , \41680 , \41384 );
and \g456184/U$4 ( \41682 , \41679 , \41681 );
and \g456184/U$6 ( \41683 , \41613 , \41678 );
or \g456184/U$3 ( \41684 , \41682 , \41683 );
xor \g456194/U$9 ( \41685 , \41293 , \41310 );
xor \g456194/U$9_r1 ( \41686 , \41685 , \41387 );
and \g456194/U$8 ( \41687 , \41684 , \41686 );
xor \g456213/U$2 ( \41688 , \41161 , \41165 );
xor \g456213/U$1 ( \41689 , \41688 , \41170 );
xor \g456213/U$1_r1 ( \41690 , \41157 , \41245 );
xor \g456213/U$1_r2 ( \41691 , \41689 , \41690 );
xor \g456194/U$11 ( \41692 , \41293 , \41310 );
xor \g456194/U$11_r1 ( \41693 , \41692 , \41387 );
and \g456194/U$10 ( \41694 , \41691 , \41693 );
and \g456194/U$12 ( \41695 , \41684 , \41691 );
or \g456194/U$7 ( \41696 , \41687 , \41694 , \41695 );
xor \g456217/U$2 ( \41697 , \41481 , \41487 );
xor \g456217/U$1 ( \41698 , \41697 , \41492 );
xor \g456217/U$1_r1 ( \41699 , \41596 , \41603 );
xor \g456217/U$1_r2 ( \41700 , \41698 , \41699 );
xor \g133292/U$4 ( \41701 , \41696 , \41700 );
xor \g133414/U$1 ( \41702 , \41250 , \41390 );
xor \g133414/U$1_r1 ( \41703 , \41702 , \41424 );
and \g133292/U$3 ( \41704 , \41701 , \41703 );
and \g133292/U$5 ( \41705 , \41696 , \41700 );
or \g133292/U$2 ( \41706 , \41704 , \41705 );
and \g130724/U$2 ( \41707 , \41611 , \41706 );
xor \g133272/U$1 ( \41708 , \41706 , \41611 );
and \g134861/U$2 ( \41709 , \40301 , \40956 );
and \g134861/U$3 ( \41710 , \40926 , \40391 );
nor \g134861/U$1 ( \41711 , \41709 , \41710 );
and \g134305/U$2 ( \41712 , \41711 , \40220 );
not \g134305/U$4 ( \41713 , \41711 );
and \g134305/U$3 ( \41714 , \41713 , \40219 );
nor \g134305/U$1 ( \41715 , \41712 , \41714 );
and \g134996/U$2 ( \41716 , \40979 , \40307 );
and \g134996/U$3 ( \41717 , \40278 , \41071 );
nor \g134996/U$1 ( \41718 , \41716 , \41717 );
and \g134217/U$2 ( \41719 , \41718 , \40871 );
not \g134217/U$4 ( \41720 , \41718 );
and \g134217/U$3 ( \41721 , \41720 , \40870 );
nor \g134217/U$1 ( \41722 , \41719 , \41721 );
xor \g133918/U$4 ( \41723 , \41715 , \41722 );
and \g134963/U$2 ( \41724 , \40432 , \40800 );
and \g134963/U$3 ( \41725 , \40731 , \40530 );
nor \g134963/U$1 ( \41726 , \41724 , \41725 );
and \g134456/U$2 ( \41727 , \41726 , \40388 );
not \g134456/U$4 ( \41728 , \41726 );
and \g134456/U$3 ( \41729 , \41728 , \40387 );
nor \g134456/U$1 ( \41730 , \41727 , \41729 );
and \g133918/U$3 ( \41731 , \41723 , \41730 );
and \g133918/U$5 ( \41732 , \41715 , \41722 );
or \g133918/U$2 ( \41733 , \41731 , \41732 );
xor \g456242/U$9 ( \41734 , \41657 , \41664 );
xor \g456242/U$9_r1 ( \41735 , \41734 , \41672 );
and \g456242/U$8 ( \41736 , \41733 , \41735 );
xor \g134021/U$1 ( \41737 , \41628 , \41631 );
xor \g134021/U$1_r1 ( \41738 , \41737 , \41639 );
xor \g456242/U$11 ( \41739 , \41657 , \41664 );
xor \g456242/U$11_r1 ( \41740 , \41739 , \41672 );
and \g456242/U$10 ( \41741 , \41738 , \41740 );
and \g456242/U$12 ( \41742 , \41733 , \41738 );
or \g456242/U$7 ( \41743 , \41736 , \41741 , \41742 );
and \g134761/U$2 ( \41744 , \41623 , \40067 );
not \g135284/U$1 ( \41745 , \41617 );
and \g134761/U$3 ( \41746 , \40064 , \41745 );
nor \g134761/U$1 ( \41747 , \41744 , \41746 );
and \g134226/U$2 ( \41748 , \41747 , \41325 );
not \g134226/U$4 ( \41749 , \41747 );
and \g134226/U$3 ( \41750 , \41749 , \41324 );
nor \g134226/U$1 ( \41751 , \41748 , \41750 );
xor \g135423/U$1 ( \41752 , \28682 , \28439 );
xor \g135431/U$1 ( \41753 , \28197 , \27952 );
and \g135279/U$2 ( \41754 , \41752 , \41753 );
or \g135241/U$1 ( \41755 , \41754 , \41319 );
xor \g456245/U$5 ( \41756 , \41751 , \41755 );
and \g135047/U$2 ( \41757 , \41206 , \40189 );
and \g135047/U$3 ( \41758 , \40138 , \41208 );
nor \g135047/U$1 ( \41759 , \41757 , \41758 );
and \g134589/U$2 ( \41760 , \41759 , \41215 );
not \g134589/U$4 ( \41761 , \41759 );
and \g134589/U$3 ( \41762 , \41761 , \41214 );
nor \g134589/U$1 ( \41763 , \41760 , \41762 );
and \g456245/U$4 ( \41764 , \41756 , \41763 );
and \g456245/U$6 ( \41765 , \41751 , \41755 );
or \g456245/U$3 ( \41766 , \41764 , \41765 );
and \g135126/U$2 ( \41767 , \40672 , \40472 );
and \g135126/U$3 ( \41768 , \40353 , \40858 );
nor \g135126/U$1 ( \41769 , \41767 , \41768 );
and \g134337/U$2 ( \41770 , \41769 , \40678 );
not \g134337/U$4 ( \41771 , \41769 );
and \g134337/U$3 ( \41772 , \41771 , \40677 );
nor \g134337/U$1 ( \41773 , \41770 , \41772 );
and \g135447/U$1 ( \41774 , \39892 , \39893 );
not \g135574/U$2 ( \41775 , \41774 );
nor \g135574/U$1 ( \41776 , \41775 , \40062 );
xor \g134022/U$4 ( \41777 , \41773 , \41776 );
and \g134873/U$2 ( \41778 , \40091 , \41629 );
and \g134873/U$3 ( \41779 , \41345 , \40113 );
nor \g134873/U$1 ( \41780 , \41778 , \41779 );
and \g134485/U$2 ( \41781 , \41780 , \40080 );
not \g134485/U$4 ( \41782 , \41780 );
and \g134485/U$3 ( \41783 , \41782 , \40079 );
nor \g134485/U$1 ( \41784 , \41781 , \41783 );
and \g134022/U$3 ( \41785 , \41777 , \41784 );
and \g134022/U$5 ( \41786 , \41773 , \41776 );
or \g134022/U$2 ( \41787 , \41785 , \41786 );
xor \g133730/U$4 ( \41788 , \41766 , \41787 );
and \g135104/U$2 ( \41789 , \41087 , \40158 );
and \g135104/U$3 ( \41790 , \40108 , \41328 );
nor \g135104/U$1 ( \41791 , \41789 , \41790 );
and \g134422/U$2 ( \41792 , \41791 , \41093 );
not \g134422/U$4 ( \41793 , \41791 );
and \g134422/U$3 ( \41794 , \41793 , \41092 );
nor \g134422/U$1 ( \41795 , \41792 , \41794 );
and \g134906/U$2 ( \41796 , \40175 , \41109 );
and \g134906/U$3 ( \41797 , \41144 , \40207 );
nor \g134906/U$1 ( \41798 , \41796 , \41797 );
and \g134300/U$2 ( \41799 , \41798 , \40137 );
not \g134300/U$4 ( \41800 , \41798 );
and \g134300/U$3 ( \41801 , \41800 , \40136 );
nor \g134300/U$1 ( \41802 , \41799 , \41801 );
xor \g134001/U$4 ( \41803 , \41795 , \41802 );
and \g134869/U$2 ( \41804 , \40147 , \41116 );
and \g134869/U$3 ( \41805 , \41107 , \40149 );
nor \g134869/U$1 ( \41806 , \41804 , \41805 );
and \g134499/U$2 ( \41807 , \41806 , \40107 );
not \g134499/U$4 ( \41808 , \41806 );
and \g134499/U$3 ( \41809 , \41808 , \40106 );
nor \g134499/U$1 ( \41810 , \41807 , \41809 );
and \g134001/U$3 ( \41811 , \41803 , \41810 );
and \g134001/U$5 ( \41812 , \41795 , \41802 );
or \g134001/U$2 ( \41813 , \41811 , \41812 );
and \g133730/U$3 ( \41814 , \41788 , \41813 );
and \g133730/U$5 ( \41815 , \41766 , \41787 );
or \g133730/U$2 ( \41816 , \41814 , \41815 );
xor \g456187/U$5 ( \41817 , \41743 , \41816 );
xor \g133777/U$1 ( \41818 , \41642 , \41649 );
xor \g133777/U$1_r1 ( \41819 , \41818 , \41675 );
and \g456187/U$4 ( \41820 , \41817 , \41819 );
and \g456187/U$6 ( \41821 , \41743 , \41816 );
or \g456187/U$3 ( \41822 , \41820 , \41821 );
xor \g456184/U$9 ( \41823 , \41613 , \41678 );
xor \g456184/U$9_r1 ( \41824 , \41823 , \41681 );
and \g456184/U$8 ( \41825 , \41822 , \41824 );
xor \g456240/U$2 ( \41826 , \41344 , \41347 );
xor \g456240/U$1 ( \41827 , \41826 , \41355 );
and \g135124/U$2 ( \41828 , \40091 , \41345 );
and \g135124/U$3 ( \41829 , \41116 , \40113 );
nor \g135124/U$1 ( \41830 , \41828 , \41829 );
and \g134382/U$2 ( \41831 , \41830 , \40080 );
not \g134382/U$4 ( \41832 , \41830 );
and \g134382/U$3 ( \41833 , \41832 , \40079 );
nor \g134382/U$1 ( \41834 , \41831 , \41833 );
and \g134690/U$2 ( \41835 , \40672 , \40353 );
and \g134690/U$3 ( \41836 , \40307 , \40858 );
nor \g134690/U$1 ( \41837 , \41835 , \41836 );
and \g134600/U$2 ( \41838 , \41837 , \40678 );
not \g134600/U$4 ( \41839 , \41837 );
and \g134600/U$3 ( \41840 , \41839 , \40677 );
nor \g134600/U$1 ( \41841 , \41838 , \41840 );
xor \g133900/U$4 ( \41842 , \41834 , \41841 );
and \g135019/U$2 ( \41843 , \40147 , \41107 );
and \g135019/U$3 ( \41844 , \41109 , \40149 );
nor \g135019/U$1 ( \41845 , \41843 , \41844 );
and \g134404/U$2 ( \41846 , \41845 , \40107 );
not \g134404/U$4 ( \41847 , \41845 );
and \g134404/U$3 ( \41848 , \41847 , \40106 );
nor \g134404/U$1 ( \41849 , \41846 , \41848 );
and \g133900/U$3 ( \41850 , \41842 , \41849 );
and \g133900/U$5 ( \41851 , \41834 , \41841 );
or \g133900/U$2 ( \41852 , \41850 , \41851 );
xor \g133992/U$1 ( \41853 , \41272 , \41279 );
xor \g133992/U$1_r1 ( \41854 , \41853 , \41287 );
xor \g456240/U$1_r1 ( \41855 , \41852 , \41854 );
xor \g456240/U$1_r2 ( \41856 , \41827 , \41855 );
xor \g133888/U$1 ( \41857 , \41366 , \41373 );
xor \g133888/U$1_r1 ( \41858 , \41857 , \41381 );
and \g134971/U$2 ( \41859 , \40513 , \40525 );
and \g134971/U$3 ( \41860 , \40472 , \40713 );
nor \g134971/U$1 ( \41861 , \41859 , \41860 );
and \g134256/U$2 ( \41862 , \41861 , \40521 );
not \g134256/U$4 ( \41863 , \41861 );
and \g134256/U$3 ( \41864 , \41863 , \40518 );
nor \g134256/U$1 ( \41865 , \41862 , \41864 );
and \g134978/U$2 ( \41866 , \40432 , \40731 );
and \g134978/U$3 ( \41867 , \40568 , \40530 );
nor \g134978/U$1 ( \41868 , \41866 , \41867 );
and \g134376/U$2 ( \41869 , \41868 , \40388 );
not \g134376/U$4 ( \41870 , \41868 );
and \g134376/U$3 ( \41871 , \41870 , \40387 );
nor \g134376/U$1 ( \41872 , \41869 , \41871 );
xor \g456220/U$5 ( \41873 , \41865 , \41872 );
not \g134509/U$1 ( \41874 , \41649 );
and \g456220/U$4 ( \41875 , \41873 , \41874 );
and \g456220/U$6 ( \41876 , \41865 , \41872 );
or \g456220/U$3 ( \41877 , \41875 , \41876 );
xor \g456197/U$9 ( \41878 , \41858 , \41877 );
xor \g133921/U$1 ( \41879 , \41318 , \41325 );
xor \g133921/U$1_r1 ( \41880 , \41879 , \41334 );
xor \g456197/U$9_r1 ( \41881 , \41878 , \41880 );
and \g456197/U$8 ( \41882 , \41856 , \41881 );
xor \g133900/U$1 ( \41883 , \41834 , \41841 );
xor \g133900/U$1_r1 ( \41884 , \41883 , \41849 );
xor \g456220/U$9 ( \41885 , \41865 , \41872 );
xor \g456220/U$9_r1 ( \41886 , \41885 , \41874 );
and \g456220/U$8 ( \41887 , \41884 , \41886 );
and \g134855/U$2 ( \41888 , \41206 , \40278 );
and \g134855/U$3 ( \41889 , \40189 , \41208 );
nor \g134855/U$1 ( \41890 , \41888 , \41889 );
and \g134476/U$2 ( \41891 , \41890 , \41215 );
not \g134476/U$4 ( \41892 , \41890 );
and \g134476/U$3 ( \41893 , \41892 , \41214 );
nor \g134476/U$1 ( \41894 , \41891 , \41893 );
and \g134728/U$2 ( \41895 , \40432 , \40926 );
and \g134728/U$3 ( \41896 , \40800 , \40530 );
nor \g134728/U$1 ( \41897 , \41895 , \41896 );
and \g134428/U$2 ( \41898 , \41897 , \40388 );
not \g134428/U$4 ( \41899 , \41897 );
and \g134428/U$3 ( \41900 , \41899 , \40387 );
nor \g134428/U$1 ( \41901 , \41898 , \41900 );
xor \g134010/U$4 ( \41902 , \41894 , \41901 );
and \g135065/U$2 ( \41903 , \40301 , \41144 );
and \g135065/U$3 ( \41904 , \40956 , \40391 );
nor \g135065/U$1 ( \41905 , \41903 , \41904 );
and \g134412/U$2 ( \41906 , \41905 , \40220 );
not \g134412/U$4 ( \41907 , \41905 );
and \g134412/U$3 ( \41908 , \41907 , \40219 );
nor \g134412/U$1 ( \41909 , \41906 , \41908 );
and \g134010/U$3 ( \41910 , \41902 , \41909 );
and \g134010/U$5 ( \41911 , \41894 , \41901 );
or \g134010/U$2 ( \41912 , \41910 , \41911 );
and \g134786/U$2 ( \41913 , \40513 , \40731 );
and \g134786/U$3 ( \41914 , \40568 , \40713 );
nor \g134786/U$1 ( \41915 , \41913 , \41914 );
and \g134323/U$2 ( \41916 , \41915 , \40521 );
not \g134323/U$4 ( \41917 , \41915 );
and \g134323/U$3 ( \41918 , \41917 , \40518 );
nor \g134323/U$1 ( \41919 , \41916 , \41918 );
and \g135484/U$1 ( \41920 , \39890 , \39891 );
not \g135592/U$2 ( \41921 , \41920 );
nor \g135592/U$1 ( \41922 , \41921 , \40062 );
xor \g134044/U$4 ( \41923 , \41919 , \41922 );
and \g134926/U$2 ( \41924 , \41087 , \40138 );
and \g134926/U$3 ( \41925 , \40158 , \41328 );
nor \g134926/U$1 ( \41926 , \41924 , \41925 );
and \g134395/U$2 ( \41927 , \41926 , \41093 );
not \g134395/U$4 ( \41928 , \41926 );
and \g134395/U$3 ( \41929 , \41928 , \41092 );
nor \g134395/U$1 ( \41930 , \41927 , \41929 );
and \g134044/U$3 ( \41931 , \41923 , \41930 );
and \g134044/U$5 ( \41932 , \41919 , \41922 );
or \g134044/U$2 ( \41933 , \41931 , \41932 );
xor \g133724/U$4 ( \41934 , \41912 , \41933 );
and \g135032/U$2 ( \41935 , \40672 , \40525 );
and \g135032/U$3 ( \41936 , \40472 , \40858 );
nor \g135032/U$1 ( \41937 , \41935 , \41936 );
and \g134423/U$2 ( \41938 , \41937 , \40678 );
not \g134423/U$4 ( \41939 , \41937 );
and \g134423/U$3 ( \41940 , \41939 , \40677 );
nor \g134423/U$1 ( \41941 , \41938 , \41940 );
and \g135343/U$2 ( \41942 , \41752 , \41614 );
not \g135343/U$4 ( \41943 , \41752 );
and \g135343/U$3 ( \41944 , \41943 , \41319 );
nor \g135343/U$1 ( \41945 , \41942 , \41944 );
not \g135568/U$2 ( \41946 , \41945 );
xor \g135279/U$1 ( \41947 , \41752 , \41753 );
nor \g135568/U$1 ( \41948 , \41946 , \41947 );
nand \g135144/U$1 ( \41949 , \40064 , \41948 );
and \g134654/U$2 ( \41950 , \41949 , \41755 );
not \g134654/U$4 ( \41951 , \41949 );
not \g135240/U$1 ( \41952 , \41755 );
and \g134654/U$3 ( \41953 , \41951 , \41952 );
nor \g134654/U$1 ( \41954 , \41950 , \41953 );
xor \g134026/U$4 ( \41955 , \41941 , \41954 );
and \g134708/U$2 ( \41956 , \40091 , \41774 );
and \g134708/U$3 ( \41957 , \41629 , \40113 );
nor \g134708/U$1 ( \41958 , \41956 , \41957 );
and \g134173/U$2 ( \41959 , \41958 , \40080 );
not \g134173/U$4 ( \41960 , \41958 );
and \g134173/U$3 ( \41961 , \41960 , \40079 );
nor \g134173/U$1 ( \41962 , \41959 , \41961 );
and \g134026/U$3 ( \41963 , \41955 , \41962 );
and \g134026/U$5 ( \41964 , \41941 , \41954 );
or \g134026/U$2 ( \41965 , \41963 , \41964 );
and \g133724/U$3 ( \41966 , \41934 , \41965 );
and \g133724/U$5 ( \41967 , \41912 , \41933 );
or \g133724/U$2 ( \41968 , \41966 , \41967 );
xor \g456220/U$11 ( \41969 , \41865 , \41872 );
xor \g456220/U$11_r1 ( \41970 , \41969 , \41874 );
and \g456220/U$10 ( \41971 , \41968 , \41970 );
and \g456220/U$12 ( \41972 , \41884 , \41968 );
or \g456220/U$7 ( \41973 , \41887 , \41971 , \41972 );
xor \g456197/U$11 ( \41974 , \41858 , \41877 );
xor \g456197/U$11_r1 ( \41975 , \41974 , \41880 );
and \g456197/U$10 ( \41976 , \41973 , \41975 );
and \g456197/U$12 ( \41977 , \41856 , \41973 );
or \g456197/U$7 ( \41978 , \41882 , \41976 , \41977 );
xor \g456184/U$11 ( \41979 , \41613 , \41678 );
xor \g456184/U$11_r1 ( \41980 , \41979 , \41681 );
and \g456184/U$10 ( \41981 , \41978 , \41980 );
and \g456184/U$12 ( \41982 , \41822 , \41978 );
or \g456184/U$7 ( \41983 , \41825 , \41981 , \41982 );
xor \g456197/U$5 ( \41984 , \41858 , \41877 );
and \g456197/U$4 ( \41985 , \41984 , \41880 );
and \g456197/U$6 ( \41986 , \41858 , \41877 );
or \g456197/U$3 ( \41987 , \41985 , \41986 );
xor \g456240/U$9 ( \41988 , \41344 , \41347 );
xor \g456240/U$9_r1 ( \41989 , \41988 , \41355 );
and \g456240/U$8 ( \41990 , \41852 , \41989 );
xor \g456240/U$11 ( \41991 , \41344 , \41347 );
xor \g456240/U$11_r1 ( \41992 , \41991 , \41355 );
and \g456240/U$10 ( \41993 , \41854 , \41992 );
and \g456240/U$12 ( \41994 , \41852 , \41854 );
or \g456240/U$7 ( \41995 , \41990 , \41993 , \41994 );
xor \g133554/U$4 ( \41996 , \41987 , \41995 );
xor \g456265/U$2 ( \41997 , \41115 , \41118 );
xor \g456265/U$1 ( \41998 , \41997 , \41126 );
xor \g456265/U$1_r1 ( \41999 , \41106 , \41152 );
xor \g456265/U$1_r2 ( \42000 , \41998 , \41999 );
and \g133554/U$3 ( \42001 , \41996 , \42000 );
and \g133554/U$5 ( \42002 , \41987 , \41995 );
or \g133554/U$2 ( \42003 , \42001 , \42002 );
xor \g133246/U$4 ( \42004 , \41983 , \42003 );
xor \g456194/U$2 ( \42005 , \41293 , \41310 );
xor \g456194/U$1 ( \42006 , \42005 , \41387 );
xor \g456194/U$1_r1 ( \42007 , \41684 , \41691 );
xor \g456194/U$1_r2 ( \42008 , \42006 , \42007 );
and \g133246/U$3 ( \42009 , \42004 , \42008 );
and \g133246/U$5 ( \42010 , \41983 , \42003 );
or \g133246/U$2 ( \42011 , \42009 , \42010 );
not \g130777/U$3 ( \42012 , \42011 );
xor \g133292/U$1 ( \42013 , \41696 , \41700 );
xor \g133292/U$1_r1 ( \42014 , \42013 , \41703 );
not \g130777/U$4 ( \42015 , \42014 );
or \g130777/U$2 ( \42016 , \42012 , \42015 );
xor \g133918/U$1 ( \42017 , \41715 , \41722 );
xor \g133918/U$1_r1 ( \42018 , \42017 , \41730 );
xor \g456245/U$9 ( \42019 , \41751 , \41755 );
xor \g456245/U$9_r1 ( \42020 , \42019 , \41763 );
and \g456245/U$8 ( \42021 , \42018 , \42020 );
xor \g134001/U$1 ( \42022 , \41795 , \41802 );
xor \g134001/U$1_r1 ( \42023 , \42022 , \41810 );
xor \g456245/U$11 ( \42024 , \41751 , \41755 );
xor \g456245/U$11_r1 ( \42025 , \42024 , \41763 );
and \g456245/U$10 ( \42026 , \42023 , \42025 );
and \g456245/U$12 ( \42027 , \42018 , \42023 );
or \g456245/U$7 ( \42028 , \42021 , \42026 , \42027 );
and \g134974/U$2 ( \42029 , \41623 , \40108 );
and \g134974/U$3 ( \42030 , \40067 , \41745 );
nor \g134974/U$1 ( \42031 , \42029 , \42030 );
and \g134408/U$2 ( \42032 , \42031 , \41324 );
not \g134408/U$4 ( \42033 , \42031 );
and \g134408/U$3 ( \42034 , \42033 , \41325 );
nor \g134408/U$1 ( \42035 , \42032 , \42034 );
not \g134407/U$1 ( \42036 , \42035 );
and \g134913/U$2 ( \42037 , \40513 , \40568 );
and \g134913/U$3 ( \42038 , \40525 , \40713 );
nor \g134913/U$1 ( \42039 , \42037 , \42038 );
and \g134301/U$2 ( \42040 , \42039 , \40521 );
not \g134301/U$4 ( \42041 , \42039 );
and \g134301/U$3 ( \42042 , \42041 , \40518 );
nor \g134301/U$1 ( \42043 , \42040 , \42042 );
xor \g133769/U$4 ( \42044 , \42036 , \42043 );
and \g134828/U$2 ( \42045 , \40979 , \40353 );
and \g134828/U$3 ( \42046 , \40307 , \41071 );
nor \g134828/U$1 ( \42047 , \42045 , \42046 );
and \g134364/U$2 ( \42048 , \42047 , \40871 );
not \g134364/U$4 ( \42049 , \42047 );
and \g134364/U$3 ( \42050 , \42049 , \40870 );
nor \g134364/U$1 ( \42051 , \42048 , \42050 );
and \g134735/U$2 ( \42052 , \40175 , \41107 );
and \g134735/U$3 ( \42053 , \41109 , \40207 );
nor \g134735/U$1 ( \42054 , \42052 , \42053 );
and \g134170/U$2 ( \42055 , \42054 , \40137 );
not \g134170/U$4 ( \42056 , \42054 );
and \g134170/U$3 ( \42057 , \42056 , \40136 );
nor \g134170/U$1 ( \42058 , \42055 , \42057 );
xor \g456252/U$5 ( \42059 , \42051 , \42058 );
and \g135064/U$2 ( \42060 , \40147 , \41345 );
and \g135064/U$3 ( \42061 , \41116 , \40149 );
nor \g135064/U$1 ( \42062 , \42060 , \42061 );
and \g134503/U$2 ( \42063 , \42062 , \40107 );
not \g134503/U$4 ( \42064 , \42062 );
and \g134503/U$3 ( \42065 , \42064 , \40106 );
nor \g134503/U$1 ( \42066 , \42063 , \42065 );
and \g456252/U$4 ( \42067 , \42059 , \42066 );
and \g456252/U$6 ( \42068 , \42051 , \42058 );
or \g456252/U$3 ( \42069 , \42067 , \42068 );
and \g133769/U$3 ( \42070 , \42044 , \42069 );
and \g133769/U$5 ( \42071 , \42036 , \42043 );
or \g133769/U$2 ( \42072 , \42070 , \42071 );
xor \g456189/U$5 ( \42073 , \42028 , \42072 );
xor \g133730/U$1 ( \42074 , \41766 , \41787 );
xor \g133730/U$1_r1 ( \42075 , \42074 , \41813 );
and \g456189/U$4 ( \42076 , \42073 , \42075 );
and \g456189/U$6 ( \42077 , \42028 , \42072 );
or \g456189/U$3 ( \42078 , \42076 , \42077 );
xor \g456187/U$9 ( \42079 , \41743 , \41816 );
xor \g456187/U$9_r1 ( \42080 , \42079 , \41819 );
and \g456187/U$8 ( \42081 , \42078 , \42080 );
and \g134756/U$2 ( \42082 , \40432 , \40956 );
and \g134756/U$3 ( \42083 , \40926 , \40530 );
nor \g134756/U$1 ( \42084 , \42082 , \42083 );
and \g134571/U$2 ( \42085 , \42084 , \40388 );
not \g134571/U$4 ( \42086 , \42084 );
and \g134571/U$3 ( \42087 , \42086 , \40387 );
nor \g134571/U$1 ( \42088 , \42085 , \42087 );
and \g134796/U$2 ( \42089 , \41206 , \40307 );
and \g134796/U$3 ( \42090 , \40278 , \41208 );
nor \g134796/U$1 ( \42091 , \42089 , \42090 );
and \g134466/U$2 ( \42092 , \42091 , \41215 );
not \g134466/U$4 ( \42093 , \42091 );
and \g134466/U$3 ( \42094 , \42093 , \41214 );
nor \g134466/U$1 ( \42095 , \42092 , \42094 );
xor \g133935/U$4 ( \42096 , \42088 , \42095 );
and \g134903/U$2 ( \42097 , \40513 , \40800 );
and \g134903/U$3 ( \42098 , \40731 , \40713 );
nor \g134903/U$1 ( \42099 , \42097 , \42098 );
and \g134575/U$2 ( \42100 , \42099 , \40521 );
not \g134575/U$4 ( \42101 , \42099 );
and \g134575/U$3 ( \42102 , \42101 , \40518 );
nor \g134575/U$1 ( \42103 , \42100 , \42102 );
and \g133935/U$3 ( \42104 , \42096 , \42103 );
and \g133935/U$5 ( \42105 , \42088 , \42095 );
or \g133935/U$2 ( \42106 , \42104 , \42105 );
xor \g133735/U$4 ( \42107 , \42106 , \42035 );
and \g134896/U$2 ( \42108 , \41623 , \40158 );
and \g134896/U$3 ( \42109 , \40108 , \41745 );
nor \g134896/U$1 ( \42110 , \42108 , \42109 );
and \g134564/U$2 ( \42111 , \42110 , \41325 );
not \g134564/U$4 ( \42112 , \42110 );
and \g134564/U$3 ( \42113 , \42112 , \41324 );
nor \g134564/U$1 ( \42114 , \42111 , \42113 );
and \g135078/U$2 ( \42115 , \40301 , \41109 );
and \g135078/U$3 ( \42116 , \41144 , \40391 );
nor \g135078/U$1 ( \42117 , \42115 , \42116 );
and \g134342/U$2 ( \42118 , \42117 , \40220 );
not \g134342/U$4 ( \42119 , \42117 );
and \g134342/U$3 ( \42120 , \42119 , \40219 );
nor \g134342/U$1 ( \42121 , \42118 , \42120 );
xor \g133941/U$4 ( \42122 , \42114 , \42121 );
and \g134989/U$2 ( \42123 , \40175 , \41116 );
and \g134989/U$3 ( \42124 , \41107 , \40207 );
nor \g134989/U$1 ( \42125 , \42123 , \42124 );
and \g134429/U$2 ( \42126 , \42125 , \40137 );
not \g134429/U$4 ( \42127 , \42125 );
and \g134429/U$3 ( \42128 , \42127 , \40136 );
nor \g134429/U$1 ( \42129 , \42126 , \42128 );
and \g133941/U$3 ( \42130 , \42122 , \42129 );
and \g133941/U$5 ( \42131 , \42114 , \42121 );
or \g133941/U$2 ( \42132 , \42130 , \42131 );
and \g133735/U$3 ( \42133 , \42107 , \42132 );
and \g133735/U$5 ( \42134 , \42106 , \42035 );
or \g133735/U$2 ( \42135 , \42133 , \42134 );
xor \g134022/U$1 ( \42136 , \41773 , \41776 );
xor \g134022/U$1_r1 ( \42137 , \42136 , \41784 );
xor \g133544/U$4 ( \42138 , \42135 , \42137 );
xor \g133769/U$1 ( \42139 , \42036 , \42043 );
xor \g133769/U$1_r1 ( \42140 , \42139 , \42069 );
and \g133544/U$3 ( \42141 , \42138 , \42140 );
and \g133544/U$5 ( \42142 , \42135 , \42137 );
or \g133544/U$2 ( \42143 , \42141 , \42142 );
xor \g456242/U$2 ( \42144 , \41657 , \41664 );
xor \g456242/U$1 ( \42145 , \42144 , \41672 );
xor \g456242/U$1_r1 ( \42146 , \41733 , \41738 );
xor \g456242/U$1_r2 ( \42147 , \42145 , \42146 );
xor \g133420/U$4 ( \42148 , \42143 , \42147 );
xor \g456220/U$2 ( \42149 , \41865 , \41872 );
xor \g456220/U$1 ( \42150 , \42149 , \41874 );
xor \g456220/U$1_r1 ( \42151 , \41884 , \41968 );
xor \g456220/U$1_r2 ( \42152 , \42150 , \42151 );
and \g133420/U$3 ( \42153 , \42148 , \42152 );
and \g133420/U$5 ( \42154 , \42143 , \42147 );
or \g133420/U$2 ( \42155 , \42153 , \42154 );
xor \g456187/U$11 ( \42156 , \41743 , \41816 );
xor \g456187/U$11_r1 ( \42157 , \42156 , \41819 );
and \g456187/U$10 ( \42158 , \42155 , \42157 );
and \g456187/U$12 ( \42159 , \42078 , \42155 );
or \g456187/U$7 ( \42160 , \42081 , \42158 , \42159 );
xor \g133554/U$1 ( \42161 , \41987 , \41995 );
xor \g133554/U$1_r1 ( \42162 , \42161 , \42000 );
xor \g133239/U$4 ( \42163 , \42160 , \42162 );
xor \g456184/U$2 ( \42164 , \41613 , \41678 );
xor \g456184/U$1 ( \42165 , \42164 , \41681 );
xor \g456184/U$1_r1 ( \42166 , \41822 , \41978 );
xor \g456184/U$1_r2 ( \42167 , \42165 , \42166 );
and \g133239/U$3 ( \42168 , \42163 , \42167 );
and \g133239/U$5 ( \42169 , \42160 , \42162 );
or \g133239/U$2 ( \42170 , \42168 , \42169 );
xor \g133246/U$1 ( \42171 , \41983 , \42003 );
xor \g133246/U$1_r1 ( \42172 , \42171 , \42008 );
and \g130836/U$2 ( \42173 , \42170 , \42172 );
xor \g133205/U$1 ( \42174 , \42172 , \42170 );
xor \g134026/U$1 ( \42175 , \41941 , \41954 );
xor \g134026/U$1_r1 ( \42176 , \42175 , \41962 );
xor \g456252/U$9 ( \42177 , \42051 , \42058 );
xor \g456252/U$9_r1 ( \42178 , \42177 , \42066 );
and \g456252/U$8 ( \42179 , \42176 , \42178 );
xor \g134010/U$1 ( \42180 , \41894 , \41901 );
xor \g134010/U$1_r1 ( \42181 , \42180 , \41909 );
xor \g456252/U$11 ( \42182 , \42051 , \42058 );
xor \g456252/U$11_r1 ( \42183 , \42182 , \42066 );
and \g456252/U$10 ( \42184 , \42181 , \42183 );
and \g456252/U$12 ( \42185 , \42176 , \42181 );
or \g456252/U$7 ( \42186 , \42179 , \42184 , \42185 );
and \g135097/U$2 ( \42187 , \40147 , \41629 );
and \g135097/U$3 ( \42188 , \41345 , \40149 );
nor \g135097/U$1 ( \42189 , \42187 , \42188 );
and \g134250/U$2 ( \42190 , \42189 , \40107 );
not \g134250/U$4 ( \42191 , \42189 );
and \g134250/U$3 ( \42192 , \42191 , \40106 );
nor \g134250/U$1 ( \42193 , \42190 , \42192 );
and \g135123/U$2 ( \42194 , \40979 , \40472 );
and \g135123/U$3 ( \42195 , \40353 , \41071 );
nor \g135123/U$1 ( \42196 , \42194 , \42195 );
and \g134356/U$2 ( \42197 , \42196 , \40871 );
not \g134356/U$4 ( \42198 , \42196 );
and \g134356/U$3 ( \42199 , \42198 , \40870 );
nor \g134356/U$1 ( \42200 , \42197 , \42199 );
xor \g133949/U$4 ( \42201 , \42193 , \42200 );
and \g134857/U$2 ( \42202 , \40091 , \41920 );
and \g134857/U$3 ( \42203 , \41774 , \40113 );
nor \g134857/U$1 ( \42204 , \42202 , \42203 );
and \g134181/U$2 ( \42205 , \42204 , \40080 );
not \g134181/U$4 ( \42206 , \42204 );
and \g134181/U$3 ( \42207 , \42206 , \40079 );
nor \g134181/U$1 ( \42208 , \42205 , \42207 );
and \g133949/U$3 ( \42209 , \42201 , \42208 );
and \g133949/U$5 ( \42210 , \42193 , \42200 );
or \g133949/U$2 ( \42211 , \42209 , \42210 );
and \g134806/U$2 ( \42212 , \41948 , \40067 );
and \g134806/U$3 ( \42213 , \40064 , \41947 );
nor \g134806/U$1 ( \42214 , \42212 , \42213 );
and \g134616/U$2 ( \42215 , \42214 , \41755 );
not \g134616/U$4 ( \42216 , \42214 );
and \g134616/U$3 ( \42217 , \42216 , \41952 );
nor \g134616/U$1 ( \42218 , \42215 , \42217 );
xnor \g135435/U$1 ( \42219 , \27220 , \26979 );
not \g135239/U$3 ( \42220 , \42219 );
xnor \g135397/U$1 ( \42221 , \27707 , \27464 );
not \g135239/U$4 ( \42222 , \42221 );
and \g135239/U$2 ( \42223 , \42220 , \42222 );
not \g135430/U$1 ( \42224 , \41753 );
nor \g135239/U$1 ( \42225 , \42223 , \42224 );
not \g135238/U$1 ( \42226 , \42225 );
xor \g456238/U$5 ( \42227 , \42218 , \42226 );
and \g135031/U$2 ( \42228 , \41087 , \40189 );
and \g135031/U$3 ( \42229 , \40138 , \41328 );
nor \g135031/U$1 ( \42230 , \42228 , \42229 );
and \g134594/U$2 ( \42231 , \42230 , \41093 );
not \g134594/U$4 ( \42232 , \42230 );
and \g134594/U$3 ( \42233 , \42232 , \41092 );
nor \g134594/U$1 ( \42234 , \42231 , \42233 );
and \g456238/U$4 ( \42235 , \42227 , \42234 );
and \g456238/U$6 ( \42236 , \42218 , \42226 );
or \g456238/U$3 ( \42237 , \42235 , \42236 );
xor \g133741/U$4 ( \42238 , \42211 , \42237 );
xor \g134044/U$1 ( \42239 , \41919 , \41922 );
xor \g134044/U$1_r1 ( \42240 , \42239 , \41930 );
and \g133741/U$3 ( \42241 , \42238 , \42240 );
and \g133741/U$5 ( \42242 , \42211 , \42237 );
or \g133741/U$2 ( \42243 , \42241 , \42242 );
xor \g456180/U$5 ( \42244 , \42186 , \42243 );
xor \g133724/U$1 ( \42245 , \41912 , \41933 );
xor \g133724/U$1_r1 ( \42246 , \42245 , \41965 );
and \g456180/U$4 ( \42247 , \42244 , \42246 );
and \g456180/U$6 ( \42248 , \42186 , \42243 );
or \g456180/U$3 ( \42249 , \42247 , \42248 );
xor \g456189/U$9 ( \42250 , \42028 , \42072 );
xor \g456189/U$9_r1 ( \42251 , \42250 , \42075 );
and \g456189/U$8 ( \42252 , \42249 , \42251 );
and \g134997/U$2 ( \42253 , \41206 , \40353 );
and \g134997/U$3 ( \42254 , \40307 , \41208 );
nor \g134997/U$1 ( \42255 , \42253 , \42254 );
and \g134303/U$2 ( \42256 , \42255 , \41215 );
not \g134303/U$4 ( \42257 , \42255 );
and \g134303/U$3 ( \42258 , \42257 , \41214 );
nor \g134303/U$1 ( \42259 , \42256 , \42258 );
and \g134720/U$2 ( \42260 , \40301 , \41107 );
and \g134720/U$3 ( \42261 , \41109 , \40391 );
nor \g134720/U$1 ( \42262 , \42260 , \42261 );
and \g134263/U$2 ( \42263 , \42262 , \40220 );
not \g134263/U$4 ( \42264 , \42262 );
and \g134263/U$3 ( \42265 , \42264 , \40219 );
nor \g134263/U$1 ( \42266 , \42263 , \42265 );
xor \g134029/U$4 ( \42267 , \42259 , \42266 );
and \g134724/U$2 ( \42268 , \40175 , \41345 );
and \g134724/U$3 ( \42269 , \41116 , \40207 );
nor \g134724/U$1 ( \42270 , \42268 , \42269 );
and \g134563/U$2 ( \42271 , \42270 , \40137 );
not \g134563/U$4 ( \42272 , \42270 );
and \g134563/U$3 ( \42273 , \42272 , \40136 );
nor \g134563/U$1 ( \42274 , \42271 , \42273 );
and \g134029/U$3 ( \42275 , \42267 , \42274 );
and \g134029/U$5 ( \42276 , \42259 , \42266 );
or \g134029/U$2 ( \42277 , \42275 , \42276 );
and \g134879/U$2 ( \42278 , \40432 , \41144 );
and \g134879/U$3 ( \42279 , \40956 , \40530 );
nor \g134879/U$1 ( \42280 , \42278 , \42279 );
and \g134219/U$2 ( \42281 , \42280 , \40388 );
not \g134219/U$4 ( \42282 , \42280 );
and \g134219/U$3 ( \42283 , \42282 , \40387 );
nor \g134219/U$1 ( \42284 , \42281 , \42283 );
and \g135007/U$2 ( \42285 , \41087 , \40278 );
and \g135007/U$3 ( \42286 , \40189 , \41328 );
nor \g135007/U$1 ( \42287 , \42285 , \42286 );
and \g134267/U$2 ( \42288 , \42287 , \41093 );
not \g134267/U$4 ( \42289 , \42287 );
and \g134267/U$3 ( \42290 , \42289 , \41092 );
nor \g134267/U$1 ( \42291 , \42288 , \42290 );
xor \g133890/U$4 ( \42292 , \42284 , \42291 );
and \g134829/U$2 ( \42293 , \40513 , \40926 );
and \g134829/U$3 ( \42294 , \40800 , \40713 );
nor \g134829/U$1 ( \42295 , \42293 , \42294 );
and \g134448/U$2 ( \42296 , \42295 , \40521 );
not \g134448/U$4 ( \42297 , \42295 );
and \g134448/U$3 ( \42298 , \42297 , \40518 );
nor \g134448/U$1 ( \42299 , \42296 , \42298 );
and \g133890/U$3 ( \42300 , \42292 , \42299 );
and \g133890/U$5 ( \42301 , \42284 , \42291 );
or \g133890/U$2 ( \42302 , \42300 , \42301 );
xor \g133772/U$4 ( \42303 , \42277 , \42302 );
and \g135041/U$2 ( \42304 , \40979 , \40525 );
and \g135041/U$3 ( \42305 , \40472 , \41071 );
nor \g135041/U$1 ( \42306 , \42304 , \42305 );
and \g134433/U$2 ( \42307 , \42306 , \40871 );
not \g134433/U$4 ( \42308 , \42306 );
and \g134433/U$3 ( \42309 , \42308 , \40870 );
nor \g134433/U$1 ( \42310 , \42307 , \42309 );
and \g135346/U$2 ( \42311 , \42221 , \42224 );
not \g135346/U$4 ( \42312 , \42221 );
and \g135346/U$3 ( \42313 , \42312 , \41753 );
nor \g135346/U$1 ( \42314 , \42311 , \42313 );
not \g135567/U$2 ( \42315 , \42314 );
xor \g135348/U$1 ( \42316 , \42221 , \42219 );
nor \g135567/U$1 ( \42317 , \42315 , \42316 );
nand \g135156/U$1 ( \42318 , \40064 , \42317 );
and \g134648/U$2 ( \42319 , \42318 , \42226 );
not \g134648/U$4 ( \42320 , \42318 );
and \g134648/U$3 ( \42321 , \42320 , \42225 );
nor \g134648/U$1 ( \42322 , \42319 , \42321 );
xor \g456234/U$5 ( \42323 , \42310 , \42322 );
and \g134826/U$2 ( \42324 , \40147 , \41774 );
and \g134826/U$3 ( \42325 , \41629 , \40149 );
nor \g134826/U$1 ( \42326 , \42324 , \42325 );
and \g134391/U$2 ( \42327 , \42326 , \40107 );
not \g134391/U$4 ( \42328 , \42326 );
and \g134391/U$3 ( \42329 , \42328 , \40106 );
nor \g134391/U$1 ( \42330 , \42327 , \42329 );
and \g456234/U$4 ( \42331 , \42323 , \42330 );
and \g456234/U$6 ( \42332 , \42310 , \42322 );
or \g456234/U$3 ( \42333 , \42331 , \42332 );
and \g133772/U$3 ( \42334 , \42303 , \42333 );
and \g133772/U$5 ( \42335 , \42277 , \42302 );
or \g133772/U$2 ( \42336 , \42334 , \42335 );
and \g134921/U$2 ( \42337 , \40672 , \40568 );
and \g134921/U$3 ( \42338 , \40525 , \40858 );
nor \g134921/U$1 ( \42339 , \42337 , \42338 );
and \g134531/U$2 ( \42340 , \42339 , \40678 );
not \g134531/U$4 ( \42341 , \42339 );
and \g134531/U$3 ( \42342 , \42341 , \40677 );
nor \g134531/U$1 ( \42343 , \42340 , \42342 );
and \g135471/U$1 ( \42344 , \39888 , \39889 );
not \g135586/U$2 ( \42345 , \42344 );
nor \g135586/U$1 ( \42346 , \42345 , \40062 );
xor \g133983/U$4 ( \42347 , \42343 , \42346 );
and \g134876/U$2 ( \42348 , \41948 , \40108 );
and \g134876/U$3 ( \42349 , \40067 , \41947 );
nor \g134876/U$1 ( \42350 , \42348 , \42349 );
and \g134597/U$2 ( \42351 , \42350 , \41952 );
not \g134597/U$4 ( \42352 , \42350 );
and \g134597/U$3 ( \42353 , \42352 , \41755 );
nor \g134597/U$1 ( \42354 , \42351 , \42353 );
not \g134596/U$1 ( \42355 , \42354 );
and \g133983/U$3 ( \42356 , \42347 , \42355 );
and \g133983/U$5 ( \42357 , \42343 , \42346 );
or \g133983/U$2 ( \42358 , \42356 , \42357 );
xor \g133573/U$4 ( \42359 , \42336 , \42358 );
xor \g133735/U$1 ( \42360 , \42106 , \42035 );
xor \g133735/U$1_r1 ( \42361 , \42360 , \42132 );
and \g133573/U$3 ( \42362 , \42359 , \42361 );
and \g133573/U$5 ( \42363 , \42336 , \42358 );
or \g133573/U$2 ( \42364 , \42362 , \42363 );
xor \g456245/U$2 ( \42365 , \41751 , \41755 );
xor \g456245/U$1 ( \42366 , \42365 , \41763 );
xor \g456245/U$1_r1 ( \42367 , \42018 , \42023 );
xor \g456245/U$1_r2 ( \42368 , \42366 , \42367 );
xor \g133456/U$4 ( \42369 , \42364 , \42368 );
xor \g133544/U$1 ( \42370 , \42135 , \42137 );
xor \g133544/U$1_r1 ( \42371 , \42370 , \42140 );
and \g133456/U$3 ( \42372 , \42369 , \42371 );
and \g133456/U$5 ( \42373 , \42364 , \42368 );
or \g133456/U$2 ( \42374 , \42372 , \42373 );
xor \g456189/U$11 ( \42375 , \42028 , \42072 );
xor \g456189/U$11_r1 ( \42376 , \42375 , \42075 );
and \g456189/U$10 ( \42377 , \42374 , \42376 );
and \g456189/U$12 ( \42378 , \42249 , \42374 );
or \g456189/U$7 ( \42379 , \42252 , \42377 , \42378 );
xor \g456197/U$2 ( \42380 , \41858 , \41877 );
xor \g456197/U$1 ( \42381 , \42380 , \41880 );
xor \g456197/U$1_r1 ( \42382 , \41856 , \41973 );
xor \g456197/U$1_r2 ( \42383 , \42381 , \42382 );
xor \g133248/U$4 ( \42384 , \42379 , \42383 );
xor \g456187/U$2 ( \42385 , \41743 , \41816 );
xor \g456187/U$1 ( \42386 , \42385 , \41819 );
xor \g456187/U$1_r1 ( \42387 , \42078 , \42155 );
xor \g456187/U$1_r2 ( \42388 , \42386 , \42387 );
and \g133248/U$3 ( \42389 , \42384 , \42388 );
and \g133248/U$5 ( \42390 , \42379 , \42383 );
or \g133248/U$2 ( \42391 , \42389 , \42390 );
not \g130890/U$3 ( \42392 , \42391 );
xor \g133239/U$1 ( \42393 , \42160 , \42162 );
xor \g133239/U$1_r1 ( \42394 , \42393 , \42167 );
not \g130890/U$4 ( \42395 , \42394 );
or \g130890/U$2 ( \42396 , \42392 , \42395 );
xor \g133248/U$1 ( \42397 , \42379 , \42383 );
xor \g133248/U$1_r1 ( \42398 , \42397 , \42388 );
xor \g133949/U$1 ( \42399 , \42193 , \42200 );
xor \g133949/U$1_r1 ( \42400 , \42399 , \42208 );
xor \g133941/U$1 ( \42401 , \42114 , \42121 );
xor \g133941/U$1_r1 ( \42402 , \42401 , \42129 );
xor \g456210/U$5 ( \42403 , \42400 , \42402 );
xor \g133983/U$1 ( \42404 , \42343 , \42346 );
xor \g133983/U$1_r1 ( \42405 , \42404 , \42355 );
and \g456210/U$4 ( \42406 , \42403 , \42405 );
and \g456210/U$6 ( \42407 , \42400 , \42402 );
or \g456210/U$3 ( \42408 , \42406 , \42407 );
and \g134837/U$2 ( \42409 , \40091 , \42344 );
and \g134837/U$3 ( \42410 , \41920 , \40113 );
nor \g134837/U$1 ( \42411 , \42409 , \42410 );
and \g134517/U$2 ( \42412 , \42411 , \40080 );
not \g134517/U$4 ( \42413 , \42411 );
and \g134517/U$3 ( \42414 , \42413 , \40079 );
nor \g134517/U$1 ( \42415 , \42412 , \42414 );
and \g135459/U$1 ( \42416 , \39886 , \39887 );
not \g135580/U$2 ( \42417 , \42416 );
nor \g135580/U$1 ( \42418 , \42417 , \40062 );
xor \g133980/U$4 ( \42419 , \42415 , \42418 );
and \g135048/U$2 ( \42420 , \41623 , \40138 );
and \g135048/U$3 ( \42421 , \40158 , \41745 );
nor \g135048/U$1 ( \42422 , \42420 , \42421 );
and \g134455/U$2 ( \42423 , \42422 , \41325 );
not \g134455/U$4 ( \42424 , \42422 );
and \g134455/U$3 ( \42425 , \42424 , \41324 );
nor \g134455/U$1 ( \42426 , \42423 , \42425 );
and \g133980/U$3 ( \42427 , \42419 , \42426 );
and \g133980/U$5 ( \42428 , \42415 , \42418 );
or \g133980/U$2 ( \42429 , \42427 , \42428 );
xor \g456238/U$9 ( \42430 , \42218 , \42226 );
xor \g456238/U$9_r1 ( \42431 , \42430 , \42234 );
and \g456238/U$8 ( \42432 , \42429 , \42431 );
xor \g133935/U$1 ( \42433 , \42088 , \42095 );
xor \g133935/U$1_r1 ( \42434 , \42433 , \42103 );
xor \g456238/U$11 ( \42435 , \42218 , \42226 );
xor \g456238/U$11_r1 ( \42436 , \42435 , \42234 );
and \g456238/U$10 ( \42437 , \42434 , \42436 );
and \g456238/U$12 ( \42438 , \42429 , \42434 );
or \g456238/U$7 ( \42439 , \42432 , \42437 , \42438 );
xor \g456186/U$5 ( \42440 , \42408 , \42439 );
xor \g133741/U$1 ( \42441 , \42211 , \42237 );
xor \g133741/U$1_r1 ( \42442 , \42441 , \42240 );
and \g456186/U$4 ( \42443 , \42440 , \42442 );
and \g456186/U$6 ( \42444 , \42408 , \42439 );
or \g456186/U$3 ( \42445 , \42443 , \42444 );
xor \g456180/U$9 ( \42446 , \42186 , \42243 );
xor \g456180/U$9_r1 ( \42447 , \42446 , \42246 );
and \g456180/U$8 ( \42448 , \42445 , \42447 );
and \g135043/U$2 ( \42449 , \40672 , \40800 );
and \g135043/U$3 ( \42450 , \40731 , \40858 );
nor \g135043/U$1 ( \42451 , \42449 , \42450 );
and \g134496/U$2 ( \42452 , \42451 , \40678 );
not \g134496/U$4 ( \42453 , \42451 );
and \g134496/U$3 ( \42454 , \42453 , \40677 );
nor \g134496/U$1 ( \42455 , \42452 , \42454 );
and \g134688/U$2 ( \42456 , \41087 , \40307 );
and \g134688/U$3 ( \42457 , \40278 , \41328 );
nor \g134688/U$1 ( \42458 , \42456 , \42457 );
and \g134554/U$2 ( \42459 , \42458 , \41093 );
not \g134554/U$4 ( \42460 , \42458 );
and \g134554/U$3 ( \42461 , \42460 , \41092 );
nor \g134554/U$1 ( \42462 , \42459 , \42461 );
xor \g133956/U$4 ( \42463 , \42455 , \42462 );
and \g134927/U$2 ( \42464 , \40513 , \40956 );
and \g134927/U$3 ( \42465 , \40926 , \40713 );
nor \g134927/U$1 ( \42466 , \42464 , \42465 );
and \g134459/U$2 ( \42467 , \42466 , \40521 );
not \g134459/U$4 ( \42468 , \42466 );
and \g134459/U$3 ( \42469 , \42468 , \40518 );
nor \g134459/U$1 ( \42470 , \42467 , \42469 );
and \g133956/U$3 ( \42471 , \42463 , \42470 );
and \g133956/U$5 ( \42472 , \42455 , \42462 );
or \g133956/U$2 ( \42473 , \42471 , \42472 );
and \g134885/U$2 ( \42474 , \41623 , \40189 );
and \g134885/U$3 ( \42475 , \40138 , \41745 );
nor \g134885/U$1 ( \42476 , \42474 , \42475 );
and \g134213/U$2 ( \42477 , \42476 , \41325 );
not \g134213/U$4 ( \42478 , \42476 );
and \g134213/U$3 ( \42479 , \42478 , \41324 );
nor \g134213/U$1 ( \42480 , \42477 , \42479 );
xnor \g135427/U$1 ( \42481 , \26244 , \26002 );
not \g135247/U$3 ( \42482 , \42481 );
xnor \g135403/U$1 ( \42483 , \26736 , \26490 );
not \g135247/U$4 ( \42484 , \42483 );
and \g135247/U$2 ( \42485 , \42482 , \42484 );
nor \g135247/U$1 ( \42486 , \42485 , \42219 );
not \g135246/U$1 ( \42487 , \42486 );
xor \g456254/U$5 ( \42488 , \42480 , \42487 );
and \g134830/U$2 ( \42489 , \42317 , \40067 );
and \g134830/U$3 ( \42490 , \40064 , \42316 );
nor \g134830/U$1 ( \42491 , \42489 , \42490 );
and \g134384/U$2 ( \42492 , \42491 , \42226 );
not \g134384/U$4 ( \42493 , \42491 );
and \g134384/U$3 ( \42494 , \42493 , \42225 );
nor \g134384/U$1 ( \42495 , \42492 , \42494 );
and \g456254/U$4 ( \42496 , \42488 , \42495 );
and \g456254/U$6 ( \42497 , \42480 , \42487 );
or \g456254/U$3 ( \42498 , \42496 , \42497 );
xor \g133685/U$4 ( \42499 , \42473 , \42498 );
and \g134932/U$2 ( \42500 , \40301 , \41116 );
and \g134932/U$3 ( \42501 , \41107 , \40391 );
nor \g134932/U$1 ( \42502 , \42500 , \42501 );
and \g134304/U$2 ( \42503 , \42502 , \40220 );
not \g134304/U$4 ( \42504 , \42502 );
and \g134304/U$3 ( \42505 , \42504 , \40219 );
nor \g134304/U$1 ( \42506 , \42503 , \42505 );
and \g134798/U$2 ( \42507 , \41948 , \40158 );
and \g134798/U$3 ( \42508 , \40108 , \41947 );
nor \g134798/U$1 ( \42509 , \42507 , \42508 );
and \g134613/U$2 ( \42510 , \42509 , \41755 );
not \g134613/U$4 ( \42511 , \42509 );
and \g134613/U$3 ( \42512 , \42511 , \41952 );
nor \g134613/U$1 ( \42513 , \42510 , \42512 );
xor \g456228/U$5 ( \42514 , \42506 , \42513 );
and \g135138/U$2 ( \42515 , \40432 , \41109 );
and \g135138/U$3 ( \42516 , \41144 , \40530 );
nor \g135138/U$1 ( \42517 , \42515 , \42516 );
and \g134242/U$2 ( \42518 , \42517 , \40388 );
not \g134242/U$4 ( \42519 , \42517 );
and \g134242/U$3 ( \42520 , \42519 , \40387 );
nor \g134242/U$1 ( \42521 , \42518 , \42520 );
and \g456228/U$4 ( \42522 , \42514 , \42521 );
and \g456228/U$6 ( \42523 , \42506 , \42513 );
or \g456228/U$3 ( \42524 , \42522 , \42523 );
and \g133685/U$3 ( \42525 , \42499 , \42524 );
and \g133685/U$5 ( \42526 , \42473 , \42498 );
or \g133685/U$2 ( \42527 , \42525 , \42526 );
and \g135068/U$2 ( \42528 , \40672 , \40731 );
and \g135068/U$3 ( \42529 , \40568 , \40858 );
nor \g135068/U$1 ( \42530 , \42528 , \42529 );
and \g134366/U$2 ( \42531 , \42530 , \40678 );
not \g134366/U$4 ( \42532 , \42530 );
and \g134366/U$3 ( \42533 , \42532 , \40677 );
nor \g134366/U$1 ( \42534 , \42531 , \42533 );
xor \g133715/U$4 ( \42535 , \42354 , \42534 );
and \g134820/U$2 ( \42536 , \40147 , \41920 );
and \g134820/U$3 ( \42537 , \41774 , \40149 );
nor \g134820/U$1 ( \42538 , \42536 , \42537 );
and \g134328/U$2 ( \42539 , \42538 , \40107 );
not \g134328/U$4 ( \42540 , \42538 );
and \g134328/U$3 ( \42541 , \42540 , \40106 );
nor \g134328/U$1 ( \42542 , \42539 , \42541 );
and \g134849/U$2 ( \42543 , \41206 , \40472 );
and \g134849/U$3 ( \42544 , \40353 , \41208 );
nor \g134849/U$1 ( \42545 , \42543 , \42544 );
and \g134415/U$2 ( \42546 , \42545 , \41215 );
not \g134415/U$4 ( \42547 , \42545 );
and \g134415/U$3 ( \42548 , \42547 , \41214 );
nor \g134415/U$1 ( \42549 , \42546 , \42548 );
xor \g133895/U$4 ( \42550 , \42542 , \42549 );
and \g135092/U$2 ( \42551 , \40175 , \41629 );
and \g135092/U$3 ( \42552 , \41345 , \40207 );
nor \g135092/U$1 ( \42553 , \42551 , \42552 );
and \g134482/U$2 ( \42554 , \42553 , \40137 );
not \g134482/U$4 ( \42555 , \42553 );
and \g134482/U$3 ( \42556 , \42555 , \40136 );
nor \g134482/U$1 ( \42557 , \42554 , \42556 );
and \g133895/U$3 ( \42558 , \42550 , \42557 );
and \g133895/U$5 ( \42559 , \42542 , \42549 );
or \g133895/U$2 ( \42560 , \42558 , \42559 );
and \g133715/U$3 ( \42561 , \42535 , \42560 );
and \g133715/U$5 ( \42562 , \42354 , \42534 );
or \g133715/U$2 ( \42563 , \42561 , \42562 );
xor \g133514/U$4 ( \42564 , \42527 , \42563 );
xor \g133772/U$1 ( \42565 , \42277 , \42302 );
xor \g133772/U$1_r1 ( \42566 , \42565 , \42333 );
and \g133514/U$3 ( \42567 , \42564 , \42566 );
and \g133514/U$5 ( \42568 , \42527 , \42563 );
or \g133514/U$2 ( \42569 , \42567 , \42568 );
xor \g456252/U$2 ( \42570 , \42051 , \42058 );
xor \g456252/U$1 ( \42571 , \42570 , \42066 );
xor \g456252/U$1_r1 ( \42572 , \42176 , \42181 );
xor \g456252/U$1_r2 ( \42573 , \42571 , \42572 );
xor \g133401/U$4 ( \42574 , \42569 , \42573 );
xor \g133573/U$1 ( \42575 , \42336 , \42358 );
xor \g133573/U$1_r1 ( \42576 , \42575 , \42361 );
and \g133401/U$3 ( \42577 , \42574 , \42576 );
and \g133401/U$5 ( \42578 , \42569 , \42573 );
or \g133401/U$2 ( \42579 , \42577 , \42578 );
xor \g456180/U$11 ( \42580 , \42186 , \42243 );
xor \g456180/U$11_r1 ( \42581 , \42580 , \42246 );
and \g456180/U$10 ( \42582 , \42579 , \42581 );
and \g456180/U$12 ( \42583 , \42445 , \42579 );
or \g456180/U$7 ( \42584 , \42448 , \42582 , \42583 );
xor \g133420/U$1 ( \42585 , \42143 , \42147 );
xor \g133420/U$1_r1 ( \42586 , \42585 , \42152 );
xor \g133217/U$4 ( \42587 , \42584 , \42586 );
xor \g456189/U$2 ( \42588 , \42028 , \42072 );
xor \g456189/U$1 ( \42589 , \42588 , \42075 );
xor \g456189/U$1_r1 ( \42590 , \42249 , \42374 );
xor \g456189/U$1_r2 ( \42591 , \42589 , \42590 );
and \g133217/U$3 ( \42592 , \42587 , \42591 );
and \g133217/U$5 ( \42593 , \42584 , \42586 );
or \g133217/U$2 ( \42594 , \42592 , \42593 );
and \g130945/U$2 ( \42595 , \42398 , \42594 );
xor \g133189/U$1 ( \42596 , \42594 , \42398 );
xor \g133895/U$1 ( \42597 , \42542 , \42549 );
xor \g133895/U$1_r1 ( \42598 , \42597 , \42557 );
xor \g456254/U$9 ( \42599 , \42480 , \42487 );
xor \g456254/U$9_r1 ( \42600 , \42599 , \42495 );
and \g456254/U$8 ( \42601 , \42598 , \42600 );
and \g134911/U$2 ( \42602 , \40979 , \40568 );
and \g134911/U$3 ( \42603 , \40525 , \41071 );
nor \g134911/U$1 ( \42604 , \42602 , \42603 );
and \g134211/U$2 ( \42605 , \42604 , \40871 );
not \g134211/U$4 ( \42606 , \42604 );
and \g134211/U$3 ( \42607 , \42606 , \40870 );
nor \g134211/U$1 ( \42608 , \42605 , \42607 );
and \g135506/U$1 ( \42609 , \39884 , \39885 );
not \g135602/U$2 ( \42610 , \42609 );
nor \g135602/U$1 ( \42611 , \42610 , \40062 );
xor \g133990/U$1 ( \42612 , \42608 , \42611 );
and \g135096/U$2 ( \42613 , \40091 , \42416 );
and \g135096/U$3 ( \42614 , \42344 , \40113 );
nor \g135096/U$1 ( \42615 , \42613 , \42614 );
and \g134282/U$2 ( \42616 , \42615 , \40080 );
not \g134282/U$4 ( \42617 , \42615 );
and \g134282/U$3 ( \42618 , \42617 , \40079 );
nor \g134282/U$1 ( \42619 , \42616 , \42618 );
xor \g133990/U$1_r1 ( \42620 , \42612 , \42619 );
xor \g456254/U$11 ( \42621 , \42480 , \42487 );
xor \g456254/U$11_r1 ( \42622 , \42621 , \42495 );
and \g456254/U$10 ( \42623 , \42620 , \42622 );
and \g456254/U$12 ( \42624 , \42598 , \42620 );
or \g456254/U$7 ( \42625 , \42601 , \42623 , \42624 );
xor \g133980/U$1 ( \42626 , \42415 , \42418 );
xor \g133980/U$1_r1 ( \42627 , \42626 , \42426 );
xor \g133990/U$4 ( \42628 , \42608 , \42611 );
and \g133990/U$3 ( \42629 , \42628 , \42619 );
and \g133990/U$5 ( \42630 , \42608 , \42611 );
or \g133990/U$2 ( \42631 , \42629 , \42630 );
xor \g456200/U$9 ( \42632 , \42627 , \42631 );
xor \g133890/U$1 ( \42633 , \42284 , \42291 );
xor \g133890/U$1_r1 ( \42634 , \42633 , \42299 );
xor \g456200/U$9_r1 ( \42635 , \42632 , \42634 );
and \g456200/U$8 ( \42636 , \42625 , \42635 );
not \g135329/U$3 ( \42637 , \42483 );
not \g135329/U$4 ( \42638 , \42219 );
and \g135329/U$2 ( \42639 , \42637 , \42638 );
and \g135329/U$5 ( \42640 , \42219 , \42483 );
nor \g135329/U$1 ( \42641 , \42639 , \42640 );
not \g135569/U$2 ( \42642 , \42641 );
xor \g135340/U$1 ( \42643 , \42483 , \42481 );
nor \g135569/U$1 ( \42644 , \42642 , \42643 );
nand \g135146/U$1 ( \42645 , \40064 , \42644 );
and \g134652/U$2 ( \42646 , \42645 , \42487 );
not \g134652/U$4 ( \42647 , \42645 );
and \g134652/U$3 ( \42648 , \42647 , \42486 );
nor \g134652/U$1 ( \42649 , \42646 , \42648 );
not \g134651/U$1 ( \42650 , \42649 );
and \g135480/U$1 ( \42651 , \39882 , \39883 );
not \g135590/U$2 ( \42652 , \42651 );
nor \g135590/U$1 ( \42653 , \42652 , \40062 );
xor \g133995/U$4 ( \42654 , \42650 , \42653 );
and \g134679/U$2 ( \42655 , \40091 , \42609 );
and \g134679/U$3 ( \42656 , \42416 , \40113 );
nor \g134679/U$1 ( \42657 , \42655 , \42656 );
and \g134325/U$2 ( \42658 , \42657 , \40080 );
not \g134325/U$4 ( \42659 , \42657 );
and \g134325/U$3 ( \42660 , \42659 , \40079 );
nor \g134325/U$1 ( \42661 , \42658 , \42660 );
and \g133995/U$3 ( \42662 , \42654 , \42661 );
and \g133995/U$5 ( \42663 , \42650 , \42653 );
or \g133995/U$2 ( \42664 , \42662 , \42663 );
xor \g456228/U$9 ( \42665 , \42506 , \42513 );
xor \g456228/U$9_r1 ( \42666 , \42665 , \42521 );
and \g456228/U$8 ( \42667 , \42664 , \42666 );
and \g134883/U$2 ( \42668 , \42644 , \40067 );
and \g134883/U$3 ( \42669 , \40064 , \42643 );
nor \g134883/U$1 ( \42670 , \42668 , \42669 );
and \g134570/U$2 ( \42671 , \42670 , \42487 );
not \g134570/U$4 ( \42672 , \42670 );
and \g134570/U$3 ( \42673 , \42672 , \42486 );
nor \g134570/U$1 ( \42674 , \42671 , \42673 );
xor \g135603/U$1 ( \42675 , \25271 , \25026 );
not \g135409/U$1 ( \42676 , \42675 );
not \g135261/U$3 ( \42677 , \42676 );
xnor \g135418/U$1 ( \42678 , \25759 , \25514 );
not \g135261/U$4 ( \42679 , \42678 );
and \g135261/U$2 ( \42680 , \42677 , \42679 );
nor \g135261/U$1 ( \42681 , \42680 , \42481 );
not \g135260/U$1 ( \42682 , \42681 );
xor \g134024/U$4 ( \42683 , \42674 , \42682 );
and \g134723/U$2 ( \42684 , \41948 , \40189 );
and \g134723/U$3 ( \42685 , \40138 , \41947 );
nor \g134723/U$1 ( \42686 , \42684 , \42685 );
and \g134189/U$2 ( \42687 , \42686 , \41755 );
not \g134189/U$4 ( \42688 , \42686 );
and \g134189/U$3 ( \42689 , \42688 , \41952 );
nor \g134189/U$1 ( \42690 , \42687 , \42689 );
and \g134024/U$3 ( \42691 , \42683 , \42690 );
and \g134024/U$5 ( \42692 , \42674 , \42682 );
or \g134024/U$2 ( \42693 , \42691 , \42692 );
and \g134957/U$2 ( \42694 , \40979 , \40800 );
and \g134957/U$3 ( \42695 , \40731 , \41071 );
nor \g134957/U$1 ( \42696 , \42694 , \42695 );
and \g134236/U$2 ( \42697 , \42696 , \40871 );
not \g134236/U$4 ( \42698 , \42696 );
and \g134236/U$3 ( \42699 , \42698 , \40870 );
nor \g134236/U$1 ( \42700 , \42697 , \42699 );
and \g135488/U$1 ( \42701 , \39880 , \39881 );
not \g135594/U$2 ( \42702 , \42701 );
nor \g135594/U$1 ( \42703 , \42702 , \40062 );
xor \g456256/U$5 ( \42704 , \42700 , \42703 );
and \g135136/U$2 ( \42705 , \40672 , \40956 );
and \g135136/U$3 ( \42706 , \40926 , \40858 );
nor \g135136/U$1 ( \42707 , \42705 , \42706 );
and \g134209/U$2 ( \42708 , \42707 , \40678 );
not \g134209/U$4 ( \42709 , \42707 );
and \g134209/U$3 ( \42710 , \42709 , \40677 );
nor \g134209/U$1 ( \42711 , \42708 , \42710 );
and \g456256/U$4 ( \42712 , \42704 , \42711 );
and \g456256/U$6 ( \42713 , \42700 , \42703 );
or \g456256/U$3 ( \42714 , \42712 , \42713 );
xor \g456223/U$5 ( \42715 , \42693 , \42714 );
and \g134776/U$2 ( \42716 , \40513 , \41109 );
and \g134776/U$3 ( \42717 , \41144 , \40713 );
nor \g134776/U$1 ( \42718 , \42716 , \42717 );
and \g134542/U$2 ( \42719 , \42718 , \40521 );
not \g134542/U$4 ( \42720 , \42718 );
and \g134542/U$3 ( \42721 , \42720 , \40518 );
nor \g134542/U$1 ( \42722 , \42719 , \42721 );
and \g134757/U$2 ( \42723 , \41623 , \40307 );
and \g134757/U$3 ( \42724 , \40278 , \41745 );
nor \g134757/U$1 ( \42725 , \42723 , \42724 );
and \g134194/U$2 ( \42726 , \42725 , \41325 );
not \g134194/U$4 ( \42727 , \42725 );
and \g134194/U$3 ( \42728 , \42727 , \41324 );
nor \g134194/U$1 ( \42729 , \42726 , \42728 );
xor \g133999/U$4 ( \42730 , \42722 , \42729 );
and \g134950/U$2 ( \42731 , \40432 , \41116 );
and \g134950/U$3 ( \42732 , \41107 , \40530 );
nor \g134950/U$1 ( \42733 , \42731 , \42732 );
and \g134216/U$2 ( \42734 , \42733 , \40388 );
not \g134216/U$4 ( \42735 , \42733 );
and \g134216/U$3 ( \42736 , \42735 , \40387 );
nor \g134216/U$1 ( \42737 , \42734 , \42736 );
and \g133999/U$3 ( \42738 , \42730 , \42737 );
and \g133999/U$5 ( \42739 , \42722 , \42729 );
or \g133999/U$2 ( \42740 , \42738 , \42739 );
and \g456223/U$4 ( \42741 , \42715 , \42740 );
and \g456223/U$6 ( \42742 , \42693 , \42714 );
or \g456223/U$3 ( \42743 , \42741 , \42742 );
xor \g456228/U$11 ( \42744 , \42506 , \42513 );
xor \g456228/U$11_r1 ( \42745 , \42744 , \42521 );
and \g456228/U$10 ( \42746 , \42743 , \42745 );
and \g456228/U$12 ( \42747 , \42664 , \42743 );
or \g456228/U$7 ( \42748 , \42667 , \42746 , \42747 );
xor \g456200/U$11 ( \42749 , \42627 , \42631 );
xor \g456200/U$11_r1 ( \42750 , \42749 , \42634 );
and \g456200/U$10 ( \42751 , \42748 , \42750 );
and \g456200/U$12 ( \42752 , \42625 , \42748 );
or \g456200/U$7 ( \42753 , \42636 , \42751 , \42752 );
xor \g456210/U$2 ( \42754 , \42400 , \42402 );
xor \g456210/U$1 ( \42755 , \42754 , \42405 );
xor \g456200/U$5 ( \42756 , \42627 , \42631 );
and \g456200/U$4 ( \42757 , \42756 , \42634 );
and \g456200/U$6 ( \42758 , \42627 , \42631 );
or \g456200/U$3 ( \42759 , \42757 , \42758 );
xor \g456238/U$2 ( \42760 , \42218 , \42226 );
xor \g456238/U$1 ( \42761 , \42760 , \42234 );
xor \g456238/U$1_r1 ( \42762 , \42429 , \42434 );
xor \g456238/U$1_r2 ( \42763 , \42761 , \42762 );
xor \g456210/U$1_r1 ( \42764 , \42759 , \42763 );
xor \g456210/U$1_r2 ( \42765 , \42755 , \42764 );
xor \g133339/U$4 ( \42766 , \42753 , \42765 );
and \g135110/U$2 ( \42767 , \41206 , \40525 );
and \g135110/U$3 ( \42768 , \40472 , \41208 );
nor \g135110/U$1 ( \42769 , \42767 , \42768 );
and \g134406/U$2 ( \42770 , \42769 , \41215 );
not \g134406/U$4 ( \42771 , \42769 );
and \g134406/U$3 ( \42772 , \42771 , \41214 );
nor \g134406/U$1 ( \42773 , \42770 , \42772 );
and \g134804/U$2 ( \42774 , \41948 , \40138 );
and \g134804/U$3 ( \42775 , \40158 , \41947 );
nor \g134804/U$1 ( \42776 , \42774 , \42775 );
and \g134468/U$2 ( \42777 , \42776 , \41755 );
not \g134468/U$4 ( \42778 , \42776 );
and \g134468/U$3 ( \42779 , \42778 , \41952 );
nor \g134468/U$1 ( \42780 , \42777 , \42779 );
xor \g134016/U$4 ( \42781 , \42773 , \42780 );
and \g135034/U$2 ( \42782 , \40301 , \41345 );
and \g135034/U$3 ( \42783 , \41116 , \40391 );
nor \g135034/U$1 ( \42784 , \42782 , \42783 );
and \g134278/U$2 ( \42785 , \42784 , \40220 );
not \g134278/U$4 ( \42786 , \42784 );
and \g134278/U$3 ( \42787 , \42786 , \40219 );
nor \g134278/U$1 ( \42788 , \42785 , \42787 );
and \g134016/U$3 ( \42789 , \42781 , \42788 );
and \g134016/U$5 ( \42790 , \42773 , \42780 );
or \g134016/U$2 ( \42791 , \42789 , \42790 );
and \g134705/U$2 ( \42792 , \40147 , \42344 );
and \g134705/U$3 ( \42793 , \41920 , \40149 );
nor \g134705/U$1 ( \42794 , \42792 , \42793 );
and \g134350/U$2 ( \42795 , \42794 , \40107 );
not \g134350/U$4 ( \42796 , \42794 );
and \g134350/U$3 ( \42797 , \42796 , \40106 );
nor \g134350/U$1 ( \42798 , \42795 , \42797 );
and \g135116/U$2 ( \42799 , \40979 , \40731 );
and \g135116/U$3 ( \42800 , \40568 , \41071 );
nor \g135116/U$1 ( \42801 , \42799 , \42800 );
and \g134556/U$2 ( \42802 , \42801 , \40871 );
not \g134556/U$4 ( \42803 , \42801 );
and \g134556/U$3 ( \42804 , \42803 , \40870 );
nor \g134556/U$1 ( \42805 , \42802 , \42804 );
xor \g133893/U$4 ( \42806 , \42798 , \42805 );
and \g134717/U$2 ( \42807 , \40175 , \41774 );
and \g134717/U$3 ( \42808 , \41629 , \40207 );
nor \g134717/U$1 ( \42809 , \42807 , \42808 );
and \g134168/U$2 ( \42810 , \42809 , \40137 );
not \g134168/U$4 ( \42811 , \42809 );
and \g134168/U$3 ( \42812 , \42811 , \40136 );
nor \g134168/U$1 ( \42813 , \42810 , \42812 );
and \g133893/U$3 ( \42814 , \42806 , \42813 );
and \g133893/U$5 ( \42815 , \42798 , \42805 );
or \g133893/U$2 ( \42816 , \42814 , \42815 );
xor \g133726/U$4 ( \42817 , \42791 , \42816 );
xor \g133956/U$1 ( \42818 , \42455 , \42462 );
xor \g133956/U$1_r1 ( \42819 , \42818 , \42470 );
and \g133726/U$3 ( \42820 , \42817 , \42819 );
and \g133726/U$5 ( \42821 , \42791 , \42816 );
or \g133726/U$2 ( \42822 , \42820 , \42821 );
and \g134930/U$2 ( \42823 , \40432 , \41107 );
and \g134930/U$3 ( \42824 , \41109 , \40530 );
nor \g134930/U$1 ( \42825 , \42823 , \42824 );
and \g134215/U$2 ( \42826 , \42825 , \40388 );
not \g134215/U$4 ( \42827 , \42825 );
and \g134215/U$3 ( \42828 , \42827 , \40387 );
nor \g134215/U$1 ( \42829 , \42826 , \42828 );
and \g134823/U$2 ( \42830 , \41087 , \40353 );
and \g134823/U$3 ( \42831 , \40307 , \41328 );
nor \g134823/U$1 ( \42832 , \42830 , \42831 );
and \g134492/U$2 ( \42833 , \42832 , \41093 );
not \g134492/U$4 ( \42834 , \42832 );
and \g134492/U$3 ( \42835 , \42834 , \41092 );
nor \g134492/U$1 ( \42836 , \42833 , \42835 );
xor \g133926/U$4 ( \42837 , \42829 , \42836 );
and \g134684/U$2 ( \42838 , \40513 , \41144 );
and \g134684/U$3 ( \42839 , \40956 , \40713 );
nor \g134684/U$1 ( \42840 , \42838 , \42839 );
and \g134346/U$2 ( \42841 , \42840 , \40521 );
not \g134346/U$4 ( \42842 , \42840 );
and \g134346/U$3 ( \42843 , \42842 , \40518 );
nor \g134346/U$1 ( \42844 , \42841 , \42843 );
and \g133926/U$3 ( \42845 , \42837 , \42844 );
and \g133926/U$5 ( \42846 , \42829 , \42836 );
or \g133926/U$2 ( \42847 , \42845 , \42846 );
xor \g456229/U$5 ( \42848 , \42847 , \42649 );
and \g135004/U$2 ( \42849 , \40672 , \40926 );
and \g135004/U$3 ( \42850 , \40800 , \40858 );
nor \g135004/U$1 ( \42851 , \42849 , \42850 );
and \g134411/U$2 ( \42852 , \42851 , \40678 );
not \g134411/U$4 ( \42853 , \42851 );
and \g134411/U$3 ( \42854 , \42853 , \40677 );
nor \g134411/U$1 ( \42855 , \42852 , \42854 );
and \g134998/U$2 ( \42856 , \42317 , \40108 );
and \g134998/U$3 ( \42857 , \40067 , \42316 );
nor \g134998/U$1 ( \42858 , \42856 , \42857 );
and \g134171/U$2 ( \42859 , \42858 , \42226 );
not \g134171/U$4 ( \42860 , \42858 );
and \g134171/U$3 ( \42861 , \42860 , \42225 );
nor \g134171/U$1 ( \42862 , \42859 , \42861 );
xor \g133889/U$4 ( \42863 , \42855 , \42862 );
and \g135093/U$2 ( \42864 , \41623 , \40278 );
and \g135093/U$3 ( \42865 , \40189 , \41745 );
nor \g135093/U$1 ( \42866 , \42864 , \42865 );
and \g134515/U$2 ( \42867 , \42866 , \41325 );
not \g134515/U$4 ( \42868 , \42866 );
and \g134515/U$3 ( \42869 , \42868 , \41324 );
nor \g134515/U$1 ( \42870 , \42867 , \42869 );
and \g133889/U$3 ( \42871 , \42863 , \42870 );
and \g133889/U$5 ( \42872 , \42855 , \42862 );
or \g133889/U$2 ( \42873 , \42871 , \42872 );
and \g456229/U$4 ( \42874 , \42848 , \42873 );
and \g456229/U$6 ( \42875 , \42847 , \42649 );
or \g456229/U$3 ( \42876 , \42874 , \42875 );
xor \g133578/U$4 ( \42877 , \42822 , \42876 );
xor \g133685/U$1 ( \42878 , \42473 , \42498 );
xor \g133685/U$1_r1 ( \42879 , \42878 , \42524 );
and \g133578/U$3 ( \42880 , \42877 , \42879 );
and \g133578/U$5 ( \42881 , \42822 , \42876 );
or \g133578/U$2 ( \42882 , \42880 , \42881 );
xor \g134029/U$1 ( \42883 , \42259 , \42266 );
xor \g134029/U$1_r1 ( \42884 , \42883 , \42274 );
xor \g456234/U$9 ( \42885 , \42310 , \42322 );
xor \g456234/U$9_r1 ( \42886 , \42885 , \42330 );
and \g456234/U$8 ( \42887 , \42884 , \42886 );
xor \g133715/U$1 ( \42888 , \42354 , \42534 );
xor \g133715/U$1_r1 ( \42889 , \42888 , \42560 );
xor \g456234/U$11 ( \42890 , \42310 , \42322 );
xor \g456234/U$11_r1 ( \42891 , \42890 , \42330 );
and \g456234/U$10 ( \42892 , \42889 , \42891 );
and \g456234/U$12 ( \42893 , \42884 , \42889 );
or \g456234/U$7 ( \42894 , \42887 , \42892 , \42893 );
xor \g133430/U$1 ( \42895 , \42882 , \42894 );
xor \g133514/U$1 ( \42896 , \42527 , \42563 );
xor \g133514/U$1_r1 ( \42897 , \42896 , \42566 );
xor \g133430/U$1_r1 ( \42898 , \42895 , \42897 );
and \g133339/U$3 ( \42899 , \42766 , \42898 );
and \g133339/U$5 ( \42900 , \42753 , \42765 );
or \g133339/U$2 ( \42901 , \42899 , \42900 );
xor \g133401/U$1 ( \42902 , \42569 , \42573 );
xor \g133401/U$1_r1 ( \42903 , \42902 , \42576 );
xor \g133250/U$4 ( \42904 , \42901 , \42903 );
xor \g456186/U$2 ( \42905 , \42408 , \42439 );
xor \g456186/U$1 ( \42906 , \42905 , \42442 );
xor \g456210/U$9 ( \42907 , \42400 , \42402 );
xor \g456210/U$9_r1 ( \42908 , \42907 , \42405 );
and \g456210/U$8 ( \42909 , \42759 , \42908 );
xor \g456210/U$11 ( \42910 , \42400 , \42402 );
xor \g456210/U$11_r1 ( \42911 , \42910 , \42405 );
and \g456210/U$10 ( \42912 , \42763 , \42911 );
and \g456210/U$12 ( \42913 , \42759 , \42763 );
or \g456210/U$7 ( \42914 , \42909 , \42912 , \42913 );
xor \g133430/U$4 ( \42915 , \42882 , \42894 );
and \g133430/U$3 ( \42916 , \42915 , \42897 );
and \g133430/U$5 ( \42917 , \42882 , \42894 );
or \g133430/U$2 ( \42918 , \42916 , \42917 );
xor \g456186/U$1_r1 ( \42919 , \42914 , \42918 );
xor \g456186/U$1_r2 ( \42920 , \42906 , \42919 );
and \g133250/U$3 ( \42921 , \42904 , \42920 );
and \g133250/U$5 ( \42922 , \42901 , \42903 );
or \g133250/U$2 ( \42923 , \42921 , \42922 );
not \g131082/U$3 ( \42924 , \42923 );
xor \g456186/U$9 ( \42925 , \42408 , \42439 );
xor \g456186/U$9_r1 ( \42926 , \42925 , \42442 );
and \g456186/U$8 ( \42927 , \42914 , \42926 );
xor \g456186/U$11 ( \42928 , \42408 , \42439 );
xor \g456186/U$11_r1 ( \42929 , \42928 , \42442 );
and \g456186/U$10 ( \42930 , \42918 , \42929 );
and \g456186/U$12 ( \42931 , \42914 , \42918 );
or \g456186/U$7 ( \42932 , \42927 , \42930 , \42931 );
xor \g133456/U$1 ( \42933 , \42364 , \42368 );
xor \g133456/U$1_r1 ( \42934 , \42933 , \42371 );
xor \g133244/U$1 ( \42935 , \42932 , \42934 );
xor \g456180/U$2 ( \42936 , \42186 , \42243 );
xor \g456180/U$1 ( \42937 , \42936 , \42246 );
xor \g456180/U$1_r1 ( \42938 , \42445 , \42579 );
xor \g456180/U$1_r2 ( \42939 , \42937 , \42938 );
xor \g133244/U$1_r1 ( \42940 , \42935 , \42939 );
not \g131082/U$4 ( \42941 , \42940 );
or \g131082/U$2 ( \42942 , \42924 , \42941 );
xor \g133250/U$1 ( \42943 , \42901 , \42903 );
xor \g133250/U$1_r1 ( \42944 , \42943 , \42920 );
xor \g456254/U$2 ( \42945 , \42480 , \42487 );
xor \g456254/U$1 ( \42946 , \42945 , \42495 );
xor \g456254/U$1_r1 ( \42947 , \42598 , \42620 );
xor \g456254/U$1_r2 ( \42948 , \42946 , \42947 );
xor \g133926/U$1 ( \42949 , \42829 , \42836 );
xor \g133926/U$1_r1 ( \42950 , \42949 , \42844 );
xor \g134016/U$1 ( \42951 , \42773 , \42780 );
xor \g134016/U$1_r1 ( \42952 , \42951 , \42788 );
xor \g456202/U$5 ( \42953 , \42950 , \42952 );
xor \g133893/U$1 ( \42954 , \42798 , \42805 );
xor \g133893/U$1_r1 ( \42955 , \42954 , \42813 );
and \g456202/U$4 ( \42956 , \42953 , \42955 );
and \g456202/U$6 ( \42957 , \42950 , \42952 );
or \g456202/U$3 ( \42958 , \42956 , \42957 );
xor \g456181/U$5 ( \42959 , \42948 , \42958 );
xor \g456228/U$2 ( \42960 , \42506 , \42513 );
xor \g456228/U$1 ( \42961 , \42960 , \42521 );
xor \g456228/U$1_r1 ( \42962 , \42664 , \42743 );
xor \g456228/U$1_r2 ( \42963 , \42961 , \42962 );
and \g456181/U$4 ( \42964 , \42959 , \42963 );
and \g456181/U$6 ( \42965 , \42948 , \42958 );
or \g456181/U$3 ( \42966 , \42964 , \42965 );
xor \g456200/U$2 ( \42967 , \42627 , \42631 );
xor \g456200/U$1 ( \42968 , \42967 , \42634 );
xor \g456200/U$1_r1 ( \42969 , \42625 , \42748 );
xor \g456200/U$1_r2 ( \42970 , \42968 , \42969 );
xor \g133304/U$4 ( \42971 , \42966 , \42970 );
and \g135057/U$2 ( \42972 , \40175 , \41920 );
and \g135057/U$3 ( \42973 , \41774 , \40207 );
nor \g135057/U$1 ( \42974 , \42972 , \42973 );
or \g134161/U$2 ( \42975 , \42974 , \40136 );
nand \g134644/U$1 ( \42976 , \40136 , \42974 );
nand \g134161/U$1 ( \42977 , \42975 , \42976 );
and \g135003/U$2 ( \42978 , \41206 , \40568 );
and \g135003/U$3 ( \42979 , \40525 , \41208 );
nor \g135003/U$1 ( \42980 , \42978 , \42979 );
and \g134286/U$2 ( \42981 , \42980 , \41215 );
not \g134286/U$4 ( \42982 , \42980 );
and \g134286/U$3 ( \42983 , \42982 , \41214 );
nor \g134286/U$1 ( \42984 , \42981 , \42983 );
xor \g456269/U$5 ( \42985 , \42977 , \42984 );
and \g134895/U$2 ( \42986 , \40147 , \42416 );
and \g134895/U$3 ( \42987 , \42344 , \40149 );
nor \g134895/U$1 ( \42988 , \42986 , \42987 );
and \g134344/U$2 ( \42989 , \42988 , \40107 );
not \g134344/U$4 ( \42990 , \42988 );
and \g134344/U$3 ( \42991 , \42990 , \40106 );
nor \g134344/U$1 ( \42992 , \42989 , \42991 );
and \g456269/U$4 ( \42993 , \42985 , \42992 );
and \g456269/U$6 ( \42994 , \42977 , \42984 );
or \g456269/U$3 ( \42995 , \42993 , \42994 );
and \g134778/U$2 ( \42996 , \42317 , \40158 );
and \g134778/U$3 ( \42997 , \40108 , \42316 );
nor \g134778/U$1 ( \42998 , \42996 , \42997 );
and \g134238/U$2 ( \42999 , \42998 , \42226 );
not \g134238/U$4 ( \43000 , \42998 );
and \g134238/U$3 ( \43001 , \43000 , \42225 );
nor \g134238/U$1 ( \43002 , \42999 , \43001 );
and \g135120/U$2 ( \43003 , \41087 , \40472 );
and \g135120/U$3 ( \43004 , \40353 , \41328 );
nor \g135120/U$1 ( \43005 , \43003 , \43004 );
and \g134560/U$2 ( \43006 , \43005 , \41093 );
not \g134560/U$4 ( \43007 , \43005 );
and \g134560/U$3 ( \43008 , \43007 , \41092 );
nor \g134560/U$1 ( \43009 , \43006 , \43008 );
xor \g134045/U$4 ( \43010 , \43002 , \43009 );
and \g135112/U$2 ( \43011 , \40301 , \41629 );
and \g135112/U$3 ( \43012 , \41345 , \40391 );
nor \g135112/U$1 ( \43013 , \43011 , \43012 );
and \g134505/U$2 ( \43014 , \43013 , \40220 );
not \g134505/U$4 ( \43015 , \43013 );
and \g134505/U$3 ( \43016 , \43015 , \40219 );
nor \g134505/U$1 ( \43017 , \43014 , \43016 );
and \g134045/U$3 ( \43018 , \43010 , \43017 );
and \g134045/U$5 ( \43019 , \43002 , \43009 );
or \g134045/U$2 ( \43020 , \43018 , \43019 );
xor \g133704/U$4 ( \43021 , \42995 , \43020 );
xor \g133889/U$1 ( \43022 , \42855 , \42862 );
xor \g133889/U$1_r1 ( \43023 , \43022 , \42870 );
and \g133704/U$3 ( \43024 , \43021 , \43023 );
and \g133704/U$5 ( \43025 , \42995 , \43020 );
or \g133704/U$2 ( \43026 , \43024 , \43025 );
xor \g456229/U$9 ( \43027 , \42847 , \42649 );
xor \g456229/U$9_r1 ( \43028 , \43027 , \42873 );
and \g456229/U$8 ( \43029 , \43026 , \43028 );
xor \g133726/U$1 ( \43030 , \42791 , \42816 );
xor \g133726/U$1_r1 ( \43031 , \43030 , \42819 );
xor \g456229/U$11 ( \43032 , \42847 , \42649 );
xor \g456229/U$11_r1 ( \43033 , \43032 , \42873 );
and \g456229/U$10 ( \43034 , \43031 , \43033 );
and \g456229/U$12 ( \43035 , \43026 , \43031 );
or \g456229/U$7 ( \43036 , \43029 , \43034 , \43035 );
xor \g456234/U$2 ( \43037 , \42310 , \42322 );
xor \g456234/U$1 ( \43038 , \43037 , \42330 );
xor \g456234/U$1_r1 ( \43039 , \42884 , \42889 );
xor \g456234/U$1_r2 ( \43040 , \43038 , \43039 );
xor \g133423/U$1 ( \43041 , \43036 , \43040 );
xor \g133578/U$1 ( \43042 , \42822 , \42876 );
xor \g133578/U$1_r1 ( \43043 , \43042 , \42879 );
xor \g133423/U$1_r1 ( \43044 , \43041 , \43043 );
and \g133304/U$3 ( \43045 , \42971 , \43044 );
and \g133304/U$5 ( \43046 , \42966 , \42970 );
or \g133304/U$2 ( \43047 , \43045 , \43046 );
xor \g133423/U$4 ( \43048 , \43036 , \43040 );
and \g133423/U$3 ( \43049 , \43048 , \43043 );
and \g133423/U$5 ( \43050 , \43036 , \43040 );
or \g133423/U$2 ( \43051 , \43049 , \43050 );
xor \g133216/U$4 ( \43052 , \43047 , \43051 );
xor \g133339/U$1 ( \43053 , \42753 , \42765 );
xor \g133339/U$1_r1 ( \43054 , \43053 , \42898 );
and \g133216/U$3 ( \43055 , \43052 , \43054 );
and \g133216/U$5 ( \43056 , \43047 , \43051 );
or \g133216/U$2 ( \43057 , \43055 , \43056 );
and \g131166/U$2 ( \43058 , \42944 , \43057 );
xor \g133186/U$1 ( \43059 , \43057 , \42944 );
xor \g134045/U$1 ( \43060 , \43002 , \43009 );
xor \g134045/U$1_r1 ( \43061 , \43060 , \43017 );
xor \g456269/U$9 ( \43062 , \42977 , \42984 );
xor \g456269/U$9_r1 ( \43063 , \43062 , \42992 );
and \g456269/U$8 ( \43064 , \43061 , \43063 );
xor \g133999/U$1 ( \43065 , \42722 , \42729 );
xor \g133999/U$1_r1 ( \43066 , \43065 , \42737 );
xor \g456269/U$11 ( \43067 , \42977 , \42984 );
xor \g456269/U$11_r1 ( \43068 , \43067 , \42992 );
and \g456269/U$10 ( \43069 , \43066 , \43068 );
and \g456269/U$12 ( \43070 , \43061 , \43066 );
or \g456269/U$7 ( \43071 , \43064 , \43069 , \43070 );
xor \g456202/U$9 ( \43072 , \42950 , \42952 );
xor \g456202/U$9_r1 ( \43073 , \43072 , \42955 );
and \g456202/U$8 ( \43074 , \43071 , \43073 );
and \g135105/U$2 ( \43075 , \40979 , \40956 );
and \g135105/U$3 ( \43076 , \40926 , \41071 );
nor \g135105/U$1 ( \43077 , \43075 , \43076 );
and \g134434/U$2 ( \43078 , \43077 , \40871 );
not \g134434/U$4 ( \43079 , \43077 );
and \g134434/U$3 ( \43080 , \43079 , \40870 );
nor \g134434/U$1 ( \43081 , \43078 , \43080 );
and \g134743/U$2 ( \43082 , \42317 , \40189 );
and \g134743/U$3 ( \43083 , \40138 , \42316 );
nor \g134743/U$1 ( \43084 , \43082 , \43083 );
and \g134199/U$2 ( \43085 , \43084 , \42226 );
not \g134199/U$4 ( \43086 , \43084 );
and \g134199/U$3 ( \43087 , \43086 , \42225 );
nor \g134199/U$1 ( \43088 , \43085 , \43087 );
xor \g133962/U$4 ( \43089 , \43081 , \43088 );
and \g135330/U$2 ( \43090 , \42678 , \42675 );
not \g135330/U$4 ( \43091 , \42678 );
and \g135330/U$3 ( \43092 , \43091 , \42676 );
nor \g135330/U$1 ( \43093 , \43090 , \43092 );
not \g135344/U$3 ( \43094 , \42678 );
not \g135344/U$4 ( \43095 , \42481 );
and \g135344/U$2 ( \43096 , \43094 , \43095 );
and \g135344/U$5 ( \43097 , \42481 , \42678 );
nor \g135344/U$1 ( \43098 , \43096 , \43097 );
and \g135229/U$1 ( \43099 , \43093 , \43098 );
and \g134783/U$2 ( \43100 , \43099 , \40067 );
not \g135283/U$1 ( \43101 , \43093 );
and \g134783/U$3 ( \43102 , \40064 , \43101 );
nor \g134783/U$1 ( \43103 , \43100 , \43102 );
and \g134582/U$2 ( \43104 , \43103 , \42682 );
not \g134582/U$4 ( \43105 , \43103 );
and \g134582/U$3 ( \43106 , \43105 , \42681 );
nor \g134582/U$1 ( \43107 , \43104 , \43106 );
and \g133962/U$3 ( \43108 , \43089 , \43107 );
and \g133962/U$5 ( \43109 , \43081 , \43088 );
or \g133962/U$2 ( \43110 , \43108 , \43109 );
and \g134902/U$2 ( \43111 , \40432 , \41629 );
and \g134902/U$3 ( \43112 , \41345 , \40530 );
nor \g134902/U$1 ( \43113 , \43111 , \43112 );
and \g134276/U$2 ( \43114 , \43113 , \40388 );
not \g134276/U$4 ( \43115 , \43113 );
and \g134276/U$3 ( \43116 , \43115 , \40387 );
nor \g134276/U$1 ( \43117 , \43114 , \43116 );
and \g134929/U$2 ( \43118 , \42644 , \40158 );
and \g134929/U$3 ( \43119 , \40108 , \42643 );
nor \g134929/U$1 ( \43120 , \43118 , \43119 );
and \g134208/U$2 ( \43121 , \43120 , \42487 );
not \g134208/U$4 ( \43122 , \43120 );
and \g134208/U$3 ( \43123 , \43122 , \42486 );
nor \g134208/U$1 ( \43124 , \43121 , \43123 );
xor \g133907/U$4 ( \43125 , \43117 , \43124 );
and \g134781/U$2 ( \43126 , \41623 , \40472 );
and \g134781/U$3 ( \43127 , \40353 , \41745 );
nor \g134781/U$1 ( \43128 , \43126 , \43127 );
and \g134190/U$2 ( \43129 , \43128 , \41325 );
not \g134190/U$4 ( \43130 , \43128 );
and \g134190/U$3 ( \43131 , \43130 , \41324 );
nor \g134190/U$1 ( \43132 , \43129 , \43131 );
and \g133907/U$3 ( \43133 , \43125 , \43132 );
and \g133907/U$5 ( \43134 , \43117 , \43124 );
or \g133907/U$2 ( \43135 , \43133 , \43134 );
xor \g133740/U$4 ( \43136 , \43110 , \43135 );
and \g135011/U$2 ( \43137 , \40513 , \41116 );
and \g135011/U$3 ( \43138 , \41107 , \40713 );
nor \g135011/U$1 ( \43139 , \43137 , \43138 );
and \g134234/U$2 ( \43140 , \43139 , \40521 );
not \g134234/U$4 ( \43141 , \43139 );
and \g134234/U$3 ( \43142 , \43141 , \40518 );
nor \g134234/U$1 ( \43143 , \43140 , \43142 );
and \g134759/U$2 ( \43144 , \41948 , \40307 );
and \g134759/U$3 ( \43145 , \40278 , \41947 );
nor \g134759/U$1 ( \43146 , \43144 , \43145 );
and \g134605/U$2 ( \43147 , \43146 , \41755 );
not \g134605/U$4 ( \43148 , \43146 );
and \g134605/U$3 ( \43149 , \43148 , \41952 );
nor \g134605/U$1 ( \43150 , \43147 , \43149 );
xor \g456246/U$5 ( \43151 , \43143 , \43150 );
and \g134918/U$2 ( \43152 , \40672 , \41109 );
and \g134918/U$3 ( \43153 , \41144 , \40858 );
nor \g134918/U$1 ( \43154 , \43152 , \43153 );
and \g134322/U$2 ( \43155 , \43154 , \40678 );
not \g134322/U$4 ( \43156 , \43154 );
and \g134322/U$3 ( \43157 , \43156 , \40677 );
nor \g134322/U$1 ( \43158 , \43155 , \43157 );
and \g456246/U$4 ( \43159 , \43151 , \43158 );
and \g456246/U$6 ( \43160 , \43143 , \43150 );
or \g456246/U$3 ( \43161 , \43159 , \43160 );
and \g133740/U$3 ( \43162 , \43136 , \43161 );
and \g133740/U$5 ( \43163 , \43110 , \43135 );
or \g133740/U$2 ( \43164 , \43162 , \43163 );
nand \g135157/U$1 ( \43165 , \40064 , \43099 );
and \g134660/U$2 ( \43166 , \43165 , \42682 );
not \g134660/U$4 ( \43167 , \43165 );
and \g134660/U$3 ( \43168 , \43167 , \42681 );
nor \g134660/U$1 ( \43169 , \43166 , \43168 );
not \g134659/U$1 ( \43170 , \43169 );
xor \g456226/U$5 ( \43171 , \43170 , \42676 );
and \g135049/U$2 ( \43172 , \41206 , \40800 );
and \g135049/U$3 ( \43173 , \40731 , \41208 );
nor \g135049/U$1 ( \43174 , \43172 , \43173 );
and \g134359/U$2 ( \43175 , \43174 , \41215 );
not \g134359/U$4 ( \43176 , \43174 );
and \g134359/U$3 ( \43177 , \43176 , \41214 );
nor \g134359/U$1 ( \43178 , \43175 , \43177 );
and \g135492/U$1 ( \43179 , \39876 , \39877 );
not \g135595/U$2 ( \43180 , \43179 );
nor \g135595/U$1 ( \43181 , \43180 , \40062 );
xor \g133985/U$4 ( \43182 , \43178 , \43181 );
and \g135502/U$1 ( \43183 , \39878 , \39879 );
and \g135140/U$2 ( \43184 , \40091 , \43183 );
and \g135140/U$3 ( \43185 , \42701 , \40113 );
nor \g135140/U$1 ( \43186 , \43184 , \43185 );
and \g134358/U$2 ( \43187 , \43186 , \40080 );
not \g134358/U$4 ( \43188 , \43186 );
and \g134358/U$3 ( \43189 , \43188 , \40079 );
nor \g134358/U$1 ( \43190 , \43187 , \43189 );
and \g133985/U$3 ( \43191 , \43182 , \43190 );
and \g133985/U$5 ( \43192 , \43178 , \43181 );
or \g133985/U$2 ( \43193 , \43191 , \43192 );
and \g456226/U$4 ( \43194 , \43171 , \43193 );
and \g456226/U$6 ( \43195 , \43170 , \42676 );
or \g456226/U$3 ( \43196 , \43194 , \43195 );
xor \g133545/U$4 ( \43197 , \43164 , \43196 );
and \g134878/U$2 ( \43198 , \40091 , \42651 );
and \g134878/U$3 ( \43199 , \42609 , \40113 );
nor \g134878/U$1 ( \43200 , \43198 , \43199 );
and \g134444/U$2 ( \43201 , \43200 , \40080 );
not \g134444/U$4 ( \43202 , \43200 );
and \g134444/U$3 ( \43203 , \43202 , \40079 );
nor \g134444/U$1 ( \43204 , \43201 , \43203 );
xor \g133792/U$1 ( \43205 , \43169 , \43204 );
and \g134734/U$2 ( \43206 , \41948 , \40278 );
and \g134734/U$3 ( \43207 , \40189 , \41947 );
nor \g134734/U$1 ( \43208 , \43206 , \43207 );
and \g134182/U$2 ( \43209 , \43208 , \41755 );
not \g134182/U$4 ( \43210 , \43208 );
and \g134182/U$3 ( \43211 , \43210 , \41952 );
nor \g134182/U$1 ( \43212 , \43209 , \43211 );
not \g135600/U$2 ( \43213 , \43183 );
nor \g135600/U$1 ( \43214 , \43213 , \40062 );
xor \g133986/U$4 ( \43215 , \43212 , \43214 );
and \g134864/U$2 ( \43216 , \42644 , \40108 );
and \g134864/U$3 ( \43217 , \40067 , \42643 );
nor \g134864/U$1 ( \43218 , \43216 , \43217 );
and \g134580/U$2 ( \43219 , \43218 , \42487 );
not \g134580/U$4 ( \43220 , \43218 );
and \g134580/U$3 ( \43221 , \43220 , \42486 );
nor \g134580/U$1 ( \43222 , \43219 , \43221 );
and \g133986/U$3 ( \43223 , \43215 , \43222 );
and \g133986/U$5 ( \43224 , \43212 , \43214 );
or \g133986/U$2 ( \43225 , \43223 , \43224 );
xor \g133792/U$1_r1 ( \43226 , \43205 , \43225 );
and \g133545/U$3 ( \43227 , \43197 , \43226 );
and \g133545/U$5 ( \43228 , \43164 , \43196 );
or \g133545/U$2 ( \43229 , \43227 , \43228 );
xor \g456202/U$11 ( \43230 , \42950 , \42952 );
xor \g456202/U$11_r1 ( \43231 , \43230 , \42955 );
and \g456202/U$10 ( \43232 , \43229 , \43231 );
and \g456202/U$12 ( \43233 , \43071 , \43229 );
or \g456202/U$7 ( \43234 , \43074 , \43232 , \43233 );
xor \g456181/U$9 ( \43235 , \42948 , \42958 );
xor \g456181/U$9_r1 ( \43236 , \43235 , \42963 );
and \g456181/U$8 ( \43237 , \43234 , \43236 );
xor \g133986/U$1 ( \43238 , \43212 , \43214 );
xor \g133986/U$1_r1 ( \43239 , \43238 , \43222 );
and \g134898/U$2 ( \43240 , \40432 , \41345 );
and \g134898/U$3 ( \43241 , \41116 , \40530 );
nor \g134898/U$1 ( \43242 , \43240 , \43241 );
and \g134367/U$2 ( \43243 , \43242 , \40388 );
not \g134367/U$4 ( \43244 , \43242 );
and \g134367/U$3 ( \43245 , \43244 , \40387 );
nor \g134367/U$1 ( \43246 , \43243 , \43245 );
and \g134766/U$2 ( \43247 , \42317 , \40138 );
and \g134766/U$3 ( \43248 , \40158 , \42316 );
nor \g134766/U$1 ( \43249 , \43247 , \43248 );
and \g134347/U$2 ( \43250 , \43249 , \42226 );
not \g134347/U$4 ( \43251 , \43249 );
and \g134347/U$3 ( \43252 , \43251 , \42225 );
nor \g134347/U$1 ( \43253 , \43250 , \43252 );
xor \g133917/U$1 ( \43254 , \43246 , \43253 );
and \g134725/U$2 ( \43255 , \40513 , \41107 );
and \g134725/U$3 ( \43256 , \41109 , \40713 );
nor \g134725/U$1 ( \43257 , \43255 , \43256 );
and \g134331/U$2 ( \43258 , \43257 , \40521 );
not \g134331/U$4 ( \43259 , \43257 );
and \g134331/U$3 ( \43260 , \43259 , \40518 );
nor \g134331/U$1 ( \43261 , \43258 , \43260 );
xor \g133917/U$1_r1 ( \43262 , \43254 , \43261 );
xor \g456203/U$5 ( \43263 , \43239 , \43262 );
and \g134810/U$2 ( \43264 , \40175 , \42344 );
and \g134810/U$3 ( \43265 , \41920 , \40207 );
nor \g134810/U$1 ( \43266 , \43264 , \43265 );
and \g134471/U$2 ( \43267 , \43266 , \40137 );
not \g134471/U$4 ( \43268 , \43266 );
and \g134471/U$3 ( \43269 , \43268 , \40136 );
nor \g134471/U$1 ( \43270 , \43267 , \43269 );
and \g135073/U$2 ( \43271 , \41087 , \40525 );
and \g135073/U$3 ( \43272 , \40472 , \41328 );
nor \g135073/U$1 ( \43273 , \43271 , \43272 );
and \g134506/U$2 ( \43274 , \43273 , \41093 );
not \g134506/U$4 ( \43275 , \43273 );
and \g134506/U$3 ( \43276 , \43275 , \41092 );
nor \g134506/U$1 ( \43277 , \43274 , \43276 );
xor \g133934/U$1 ( \43278 , \43270 , \43277 );
and \g134925/U$2 ( \43279 , \40301 , \41774 );
and \g134925/U$3 ( \43280 , \41629 , \40391 );
nor \g134925/U$1 ( \43281 , \43279 , \43280 );
and \g134604/U$2 ( \43282 , \43281 , \40220 );
not \g134604/U$4 ( \43283 , \43281 );
and \g134604/U$3 ( \43284 , \43283 , \40219 );
nor \g134604/U$1 ( \43285 , \43282 , \43284 );
xor \g133934/U$1_r1 ( \43286 , \43278 , \43285 );
and \g456203/U$4 ( \43287 , \43263 , \43286 );
and \g456203/U$6 ( \43288 , \43239 , \43262 );
or \g456203/U$3 ( \43289 , \43287 , \43288 );
and \g134863/U$2 ( \43290 , \40175 , \42416 );
and \g134863/U$3 ( \43291 , \42344 , \40207 );
nor \g134863/U$1 ( \43292 , \43290 , \43291 );
and \g134599/U$2 ( \43293 , \43292 , \40137 );
not \g134599/U$4 ( \43294 , \43292 );
and \g134599/U$3 ( \43295 , \43294 , \40136 );
nor \g134599/U$1 ( \43296 , \43293 , \43295 );
and \g135027/U$2 ( \43297 , \41087 , \40568 );
and \g135027/U$3 ( \43298 , \40525 , \41328 );
nor \g135027/U$1 ( \43299 , \43297 , \43298 );
and \g134617/U$2 ( \43300 , \43299 , \41093 );
not \g134617/U$4 ( \43301 , \43299 );
and \g134617/U$3 ( \43302 , \43301 , \41092 );
nor \g134617/U$1 ( \43303 , \43300 , \43302 );
xor \g456251/U$5 ( \43304 , \43296 , \43303 );
and \g134933/U$2 ( \43305 , \40301 , \41920 );
and \g134933/U$3 ( \43306 , \41774 , \40391 );
nor \g134933/U$1 ( \43307 , \43305 , \43306 );
and \g134436/U$2 ( \43308 , \43307 , \40220 );
not \g134436/U$4 ( \43309 , \43307 );
and \g134436/U$3 ( \43310 , \43309 , \40219 );
nor \g134436/U$1 ( \43311 , \43308 , \43310 );
and \g456251/U$4 ( \43312 , \43304 , \43311 );
and \g456251/U$6 ( \43313 , \43296 , \43303 );
or \g456251/U$3 ( \43314 , \43312 , \43313 );
and \g134682/U$2 ( \43315 , \41623 , \40353 );
and \g134682/U$3 ( \43316 , \40307 , \41745 );
nor \g134682/U$1 ( \43317 , \43315 , \43316 );
and \g134473/U$2 ( \43318 , \43317 , \41325 );
not \g134473/U$4 ( \43319 , \43317 );
and \g134473/U$3 ( \43320 , \43319 , \41324 );
nor \g134473/U$1 ( \43321 , \43318 , \43320 );
and \g135075/U$2 ( \43322 , \40979 , \40926 );
and \g135075/U$3 ( \43323 , \40800 , \41071 );
nor \g135075/U$1 ( \43324 , \43322 , \43323 );
and \g134241/U$2 ( \43325 , \43324 , \40871 );
not \g134241/U$4 ( \43326 , \43324 );
and \g134241/U$3 ( \43327 , \43326 , \40870 );
nor \g134241/U$1 ( \43328 , \43325 , \43327 );
xor \g456243/U$9 ( \43329 , \43321 , \43328 );
and \g135030/U$2 ( \43330 , \40672 , \41144 );
and \g135030/U$3 ( \43331 , \40956 , \40858 );
nor \g135030/U$1 ( \43332 , \43330 , \43331 );
and \g134295/U$2 ( \43333 , \43332 , \40678 );
not \g134295/U$4 ( \43334 , \43332 );
and \g134295/U$3 ( \43335 , \43334 , \40677 );
nor \g134295/U$1 ( \43336 , \43333 , \43335 );
xor \g456243/U$9_r1 ( \43337 , \43329 , \43336 );
and \g456243/U$8 ( \43338 , \43314 , \43337 );
and \g134748/U$2 ( \43339 , \41206 , \40731 );
and \g134748/U$3 ( \43340 , \40568 , \41208 );
nor \g134748/U$1 ( \43341 , \43339 , \43340 );
and \g134318/U$2 ( \43342 , \43341 , \41215 );
not \g134318/U$4 ( \43343 , \43341 );
and \g134318/U$3 ( \43344 , \43343 , \41214 );
nor \g134318/U$1 ( \43345 , \43342 , \43344 );
and \g134714/U$2 ( \43346 , \40147 , \42609 );
and \g134714/U$3 ( \43347 , \42416 , \40149 );
nor \g134714/U$1 ( \43348 , \43346 , \43347 );
or \g134183/U$2 ( \43349 , \43348 , \40106 );
nand \g134640/U$1 ( \43350 , \40106 , \43348 );
nand \g134183/U$1 ( \43351 , \43349 , \43350 );
xor \g133974/U$1 ( \43352 , \43345 , \43351 );
and \g135029/U$2 ( \43353 , \40091 , \42701 );
and \g135029/U$3 ( \43354 , \42651 , \40113 );
nor \g135029/U$1 ( \43355 , \43353 , \43354 );
and \g134590/U$2 ( \43356 , \43355 , \40080 );
not \g134590/U$4 ( \43357 , \43355 );
and \g134590/U$3 ( \43358 , \43357 , \40079 );
nor \g134590/U$1 ( \43359 , \43356 , \43358 );
xor \g133974/U$1_r1 ( \43360 , \43352 , \43359 );
xor \g456243/U$11 ( \43361 , \43321 , \43328 );
xor \g456243/U$11_r1 ( \43362 , \43361 , \43336 );
and \g456243/U$10 ( \43363 , \43360 , \43362 );
and \g456243/U$12 ( \43364 , \43314 , \43360 );
or \g456243/U$7 ( \43365 , \43338 , \43363 , \43364 );
xor \g133555/U$4 ( \43366 , \43289 , \43365 );
xor \g133917/U$4 ( \43367 , \43246 , \43253 );
and \g133917/U$3 ( \43368 , \43367 , \43261 );
and \g133917/U$5 ( \43369 , \43246 , \43253 );
or \g133917/U$2 ( \43370 , \43368 , \43369 );
xor \g456243/U$5 ( \43371 , \43321 , \43328 );
and \g456243/U$4 ( \43372 , \43371 , \43336 );
and \g456243/U$6 ( \43373 , \43321 , \43328 );
or \g456243/U$3 ( \43374 , \43372 , \43373 );
xor \g133745/U$1 ( \43375 , \43370 , \43374 );
xor \g133934/U$4 ( \43376 , \43270 , \43277 );
and \g133934/U$3 ( \43377 , \43376 , \43285 );
and \g133934/U$5 ( \43378 , \43270 , \43277 );
or \g133934/U$2 ( \43379 , \43377 , \43378 );
xor \g133745/U$1_r1 ( \43380 , \43375 , \43379 );
and \g133555/U$3 ( \43381 , \43366 , \43380 );
and \g133555/U$5 ( \43382 , \43289 , \43365 );
or \g133555/U$2 ( \43383 , \43381 , \43382 );
xor \g133792/U$4 ( \43384 , \43169 , \43204 );
and \g133792/U$3 ( \43385 , \43384 , \43225 );
and \g133792/U$5 ( \43386 , \43169 , \43204 );
or \g133792/U$2 ( \43387 , \43385 , \43386 );
xor \g133995/U$1 ( \43388 , \42650 , \42653 );
xor \g133995/U$1_r1 ( \43389 , \43388 , \42661 );
xor \g456195/U$9 ( \43390 , \43387 , \43389 );
xor \g133745/U$4 ( \43391 , \43370 , \43374 );
and \g133745/U$3 ( \43392 , \43391 , \43379 );
and \g133745/U$5 ( \43393 , \43370 , \43374 );
or \g133745/U$2 ( \43394 , \43392 , \43393 );
xor \g456195/U$9_r1 ( \43395 , \43390 , \43394 );
and \g456195/U$8 ( \43396 , \43383 , \43395 );
xor \g456223/U$2 ( \43397 , \42693 , \42714 );
xor \g456223/U$1 ( \43398 , \43397 , \42740 );
xor \g133974/U$4 ( \43399 , \43345 , \43351 );
and \g133974/U$3 ( \43400 , \43399 , \43359 );
and \g133974/U$5 ( \43401 , \43345 , \43351 );
or \g133974/U$2 ( \43402 , \43400 , \43401 );
xor \g456256/U$9 ( \43403 , \42700 , \42703 );
xor \g456256/U$9_r1 ( \43404 , \43403 , \42711 );
and \g456256/U$8 ( \43405 , \43402 , \43404 );
xor \g134024/U$1 ( \43406 , \42674 , \42682 );
xor \g134024/U$1_r1 ( \43407 , \43406 , \42690 );
xor \g456256/U$11 ( \43408 , \42700 , \42703 );
xor \g456256/U$11_r1 ( \43409 , \43408 , \42711 );
and \g456256/U$10 ( \43410 , \43407 , \43409 );
and \g456256/U$12 ( \43411 , \43402 , \43407 );
or \g456256/U$7 ( \43412 , \43405 , \43410 , \43411 );
xor \g133704/U$1 ( \43413 , \42995 , \43020 );
xor \g133704/U$1_r1 ( \43414 , \43413 , \43023 );
xor \g456223/U$1_r1 ( \43415 , \43412 , \43414 );
xor \g456223/U$1_r2 ( \43416 , \43398 , \43415 );
xor \g456195/U$11 ( \43417 , \43387 , \43389 );
xor \g456195/U$11_r1 ( \43418 , \43417 , \43394 );
and \g456195/U$10 ( \43419 , \43416 , \43418 );
and \g456195/U$12 ( \43420 , \43383 , \43416 );
or \g456195/U$7 ( \43421 , \43396 , \43419 , \43420 );
xor \g456181/U$11 ( \43422 , \42948 , \42958 );
xor \g456181/U$11_r1 ( \43423 , \43422 , \42963 );
and \g456181/U$10 ( \43424 , \43421 , \43423 );
and \g456181/U$12 ( \43425 , \43234 , \43421 );
or \g456181/U$7 ( \43426 , \43237 , \43424 , \43425 );
xor \g456223/U$9 ( \43427 , \42693 , \42714 );
xor \g456223/U$9_r1 ( \43428 , \43427 , \42740 );
and \g456223/U$8 ( \43429 , \43412 , \43428 );
xor \g456223/U$11 ( \43430 , \42693 , \42714 );
xor \g456223/U$11_r1 ( \43431 , \43430 , \42740 );
and \g456223/U$10 ( \43432 , \43414 , \43431 );
and \g456223/U$12 ( \43433 , \43412 , \43414 );
or \g456223/U$7 ( \43434 , \43429 , \43432 , \43433 );
xor \g456195/U$5 ( \43435 , \43387 , \43389 );
and \g456195/U$4 ( \43436 , \43435 , \43394 );
and \g456195/U$6 ( \43437 , \43387 , \43389 );
or \g456195/U$3 ( \43438 , \43436 , \43437 );
xor \g133421/U$4 ( \43439 , \43434 , \43438 );
xor \g456229/U$2 ( \43440 , \42847 , \42649 );
xor \g456229/U$1 ( \43441 , \43440 , \42873 );
xor \g456229/U$1_r1 ( \43442 , \43026 , \43031 );
xor \g456229/U$1_r2 ( \43443 , \43441 , \43442 );
and \g133421/U$3 ( \43444 , \43439 , \43443 );
and \g133421/U$5 ( \43445 , \43434 , \43438 );
or \g133421/U$2 ( \43446 , \43444 , \43445 );
xor \g133241/U$4 ( \43447 , \43426 , \43446 );
xor \g133304/U$1 ( \43448 , \42966 , \42970 );
xor \g133304/U$1_r1 ( \43449 , \43448 , \43044 );
and \g133241/U$3 ( \43450 , \43447 , \43449 );
and \g133241/U$5 ( \43451 , \43426 , \43446 );
or \g133241/U$2 ( \43452 , \43450 , \43451 );
not \g131224/U$3 ( \43453 , \43452 );
xor \g133216/U$1 ( \43454 , \43047 , \43051 );
xor \g133216/U$1_r1 ( \43455 , \43454 , \43054 );
not \g131224/U$4 ( \43456 , \43455 );
or \g131224/U$2 ( \43457 , \43453 , \43456 );
xor \g133241/U$1 ( \43458 , \43426 , \43446 );
xor \g133241/U$1_r1 ( \43459 , \43458 , \43449 );
and \g134966/U$2 ( \43460 , \41623 , \40525 );
and \g134966/U$3 ( \43461 , \40472 , \41745 );
nor \g134966/U$1 ( \43462 , \43460 , \43461 );
and \g134487/U$2 ( \43463 , \43462 , \41325 );
not \g134487/U$4 ( \43464 , \43462 );
and \g134487/U$3 ( \43465 , \43464 , \41324 );
nor \g134487/U$1 ( \43466 , \43463 , \43465 );
and \g134944/U$2 ( \43467 , \42644 , \40138 );
and \g134944/U$3 ( \43468 , \40158 , \42643 );
nor \g134944/U$1 ( \43469 , \43467 , \43468 );
and \g134405/U$2 ( \43470 , \43469 , \42487 );
not \g134405/U$4 ( \43471 , \43469 );
and \g134405/U$3 ( \43472 , \43471 , \42486 );
nor \g134405/U$1 ( \43473 , \43470 , \43472 );
xor \g134017/U$4 ( \43474 , \43466 , \43473 );
and \g134951/U$2 ( \43475 , \40513 , \41345 );
and \g134951/U$3 ( \43476 , \41116 , \40713 );
nor \g134951/U$1 ( \43477 , \43475 , \43476 );
and \g134186/U$2 ( \43478 , \43477 , \40521 );
not \g134186/U$4 ( \43479 , \43477 );
and \g134186/U$3 ( \43480 , \43479 , \40518 );
nor \g134186/U$1 ( \43481 , \43478 , \43480 );
and \g134017/U$3 ( \43482 , \43474 , \43481 );
and \g134017/U$5 ( \43483 , \43466 , \43473 );
or \g134017/U$2 ( \43484 , \43482 , \43483 );
xor \g456251/U$9 ( \43485 , \43296 , \43303 );
xor \g456251/U$9_r1 ( \43486 , \43485 , \43311 );
and \g456251/U$8 ( \43487 , \43484 , \43486 );
xor \g133985/U$1 ( \43488 , \43178 , \43181 );
xor \g133985/U$1_r1 ( \43489 , \43488 , \43190 );
xor \g456251/U$11 ( \43490 , \43296 , \43303 );
xor \g456251/U$11_r1 ( \43491 , \43490 , \43311 );
and \g456251/U$10 ( \43492 , \43489 , \43491 );
and \g456251/U$12 ( \43493 , \43484 , \43489 );
or \g456251/U$7 ( \43494 , \43487 , \43492 , \43493 );
xor \g456226/U$9 ( \43495 , \43170 , \42676 );
xor \g456226/U$9_r1 ( \43496 , \43495 , \43193 );
and \g456226/U$8 ( \43497 , \43494 , \43496 );
xor \g133907/U$1 ( \43498 , \43117 , \43124 );
xor \g133907/U$1_r1 ( \43499 , \43498 , \43132 );
xor \g456246/U$9 ( \43500 , \43143 , \43150 );
xor \g456246/U$9_r1 ( \43501 , \43500 , \43158 );
and \g456246/U$8 ( \43502 , \43499 , \43501 );
xor \g133962/U$1 ( \43503 , \43081 , \43088 );
xor \g133962/U$1_r1 ( \43504 , \43503 , \43107 );
xor \g456246/U$11 ( \43505 , \43143 , \43150 );
xor \g456246/U$11_r1 ( \43506 , \43505 , \43158 );
and \g456246/U$10 ( \43507 , \43504 , \43506 );
and \g456246/U$12 ( \43508 , \43499 , \43504 );
or \g456246/U$7 ( \43509 , \43502 , \43507 , \43508 );
xor \g456226/U$11 ( \43510 , \43170 , \42676 );
xor \g456226/U$11_r1 ( \43511 , \43510 , \43193 );
and \g456226/U$10 ( \43512 , \43509 , \43511 );
and \g456226/U$12 ( \43513 , \43494 , \43509 );
or \g456226/U$7 ( \43514 , \43497 , \43512 , \43513 );
and \g135118/U$2 ( \43515 , \41206 , \40926 );
and \g135118/U$3 ( \43516 , \40800 , \41208 );
nor \g135118/U$1 ( \43517 , \43515 , \43516 );
and \g134368/U$2 ( \43518 , \43517 , \41215 );
not \g134368/U$4 ( \43519 , \43517 );
and \g134368/U$3 ( \43520 , \43519 , \41214 );
nor \g134368/U$1 ( \43521 , \43518 , \43520 );
and \g134678/U$2 ( \43522 , \42317 , \40278 );
and \g134678/U$3 ( \43523 , \40189 , \42316 );
nor \g134678/U$1 ( \43524 , \43522 , \43523 );
and \g134239/U$2 ( \43525 , \43524 , \42226 );
not \g134239/U$4 ( \43526 , \43524 );
and \g134239/U$3 ( \43527 , \43526 , \42225 );
nor \g134239/U$1 ( \43528 , \43525 , \43527 );
xor \g133957/U$4 ( \43529 , \43521 , \43528 );
and \g135039/U$2 ( \43530 , \40091 , \43179 );
and \g135039/U$3 ( \43531 , \43183 , \40113 );
nor \g135039/U$1 ( \43532 , \43530 , \43531 );
and \g134511/U$2 ( \43533 , \43532 , \40080 );
not \g134511/U$4 ( \43534 , \43532 );
and \g134511/U$3 ( \43535 , \43534 , \40079 );
nor \g134511/U$1 ( \43536 , \43533 , \43535 );
and \g133957/U$3 ( \43537 , \43529 , \43536 );
and \g133957/U$5 ( \43538 , \43521 , \43528 );
or \g133957/U$2 ( \43539 , \43537 , \43538 );
and \g134715/U$2 ( \43540 , \40672 , \41107 );
and \g134715/U$3 ( \43541 , \41109 , \40858 );
nor \g134715/U$1 ( \43542 , \43540 , \43541 );
and \g134210/U$2 ( \43543 , \43542 , \40678 );
not \g134210/U$4 ( \43544 , \43542 );
and \g134210/U$3 ( \43545 , \43544 , \40677 );
nor \g134210/U$1 ( \43546 , \43543 , \43545 );
and \g135045/U$2 ( \43547 , \41948 , \40353 );
and \g135045/U$3 ( \43548 , \40307 , \41947 );
nor \g135045/U$1 ( \43549 , \43547 , \43548 );
and \g134255/U$2 ( \43550 , \43549 , \41755 );
not \g134255/U$4 ( \43551 , \43549 );
and \g134255/U$3 ( \43552 , \43551 , \41952 );
nor \g134255/U$1 ( \43553 , \43550 , \43552 );
xor \g456249/U$5 ( \43554 , \43546 , \43553 );
and \g134897/U$2 ( \43555 , \40979 , \41144 );
and \g134897/U$3 ( \43556 , \40956 , \41071 );
nor \g134897/U$1 ( \43557 , \43555 , \43556 );
and \g134552/U$2 ( \43558 , \43557 , \40871 );
not \g134552/U$4 ( \43559 , \43557 );
and \g134552/U$3 ( \43560 , \43559 , \40870 );
nor \g134552/U$1 ( \43561 , \43558 , \43560 );
and \g456249/U$4 ( \43562 , \43554 , \43561 );
and \g456249/U$6 ( \43563 , \43546 , \43553 );
or \g456249/U$3 ( \43564 , \43562 , \43563 );
xor \g133725/U$4 ( \43565 , \43539 , \43564 );
and \g134919/U$2 ( \43566 , \40301 , \42344 );
and \g134919/U$3 ( \43567 , \41920 , \40391 );
nor \g134919/U$1 ( \43568 , \43566 , \43567 );
and \g134424/U$2 ( \43569 , \43568 , \40220 );
not \g134424/U$4 ( \43570 , \43568 );
and \g134424/U$3 ( \43571 , \43570 , \40219 );
nor \g134424/U$1 ( \43572 , \43569 , \43571 );
and \g134972/U$2 ( \43573 , \41087 , \40731 );
and \g134972/U$3 ( \43574 , \40568 , \41328 );
nor \g134972/U$1 ( \43575 , \43573 , \43574 );
and \g134574/U$2 ( \43576 , \43575 , \41093 );
not \g134574/U$4 ( \43577 , \43575 );
and \g134574/U$3 ( \43578 , \43577 , \41092 );
nor \g134574/U$1 ( \43579 , \43576 , \43578 );
xor \g133913/U$4 ( \43580 , \43572 , \43579 );
and \g134736/U$2 ( \43581 , \40432 , \41774 );
and \g134736/U$3 ( \43582 , \41629 , \40530 );
nor \g134736/U$1 ( \43583 , \43581 , \43582 );
and \g134296/U$2 ( \43584 , \43583 , \40388 );
not \g134296/U$4 ( \43585 , \43583 );
and \g134296/U$3 ( \43586 , \43585 , \40387 );
nor \g134296/U$1 ( \43587 , \43584 , \43586 );
and \g133913/U$3 ( \43588 , \43580 , \43587 );
and \g133913/U$5 ( \43589 , \43572 , \43579 );
or \g133913/U$2 ( \43590 , \43588 , \43589 );
and \g133725/U$3 ( \43591 , \43565 , \43590 );
and \g133725/U$5 ( \43592 , \43539 , \43564 );
or \g133725/U$2 ( \43593 , \43591 , \43592 );
and \g134942/U$2 ( \43594 , \40147 , \42651 );
and \g134942/U$3 ( \43595 , \42609 , \40149 );
nor \g134942/U$1 ( \43596 , \43594 , \43595 );
and \g134462/U$2 ( \43597 , \43596 , \40107 );
not \g134462/U$4 ( \43598 , \43596 );
and \g134462/U$3 ( \43599 , \43598 , \40106 );
nor \g134462/U$1 ( \43600 , \43597 , \43599 );
xor \g456227/U$5 ( \43601 , \43600 , \42675 );
not \g135571/U$2 ( \43602 , \42675 );
xor \g135402/U$1 ( \43603 , \24784 , \24540 );
nor \g135571/U$1 ( \43604 , \43602 , \43603 );
and \g135270/U$2 ( \43605 , \43604 , \40064 );
nor \g135270/U$1 ( \43606 , \43605 , \42676 );
nand \g135490/U$1 ( \43607 , \39875 , \39874 );
nor \g135349/U$1 ( \43608 , \40062 , \43607 );
xor \g134040/U$4 ( \43609 , \43606 , \43608 );
and \g134894/U$2 ( \43610 , \43099 , \40108 );
and \g134894/U$3 ( \43611 , \40067 , \43101 );
nor \g134894/U$1 ( \43612 , \43610 , \43611 );
and \g134193/U$2 ( \43613 , \43612 , \42682 );
not \g134193/U$4 ( \43614 , \43612 );
and \g134193/U$3 ( \43615 , \43614 , \42681 );
nor \g134193/U$1 ( \43616 , \43613 , \43615 );
and \g134040/U$3 ( \43617 , \43609 , \43616 );
and \g134040/U$5 ( \43618 , \43606 , \43608 );
or \g134040/U$2 ( \43619 , \43617 , \43618 );
and \g456227/U$4 ( \43620 , \43601 , \43619 );
and \g456227/U$6 ( \43621 , \43600 , \42675 );
or \g456227/U$3 ( \43622 , \43620 , \43621 );
xor \g456196/U$5 ( \43623 , \43593 , \43622 );
xor \g133740/U$1 ( \43624 , \43110 , \43135 );
xor \g133740/U$1_r1 ( \43625 , \43624 , \43161 );
and \g456196/U$4 ( \43626 , \43623 , \43625 );
and \g456196/U$6 ( \43627 , \43593 , \43622 );
or \g456196/U$3 ( \43628 , \43626 , \43627 );
xor \g133400/U$4 ( \43629 , \43514 , \43628 );
xor \g133555/U$1 ( \43630 , \43289 , \43365 );
xor \g133555/U$1_r1 ( \43631 , \43630 , \43380 );
and \g133400/U$3 ( \43632 , \43629 , \43631 );
and \g133400/U$5 ( \43633 , \43514 , \43628 );
or \g133400/U$2 ( \43634 , \43632 , \43633 );
xor \g456256/U$2 ( \43635 , \42700 , \42703 );
xor \g456256/U$1 ( \43636 , \43635 , \42711 );
xor \g456256/U$1_r1 ( \43637 , \43402 , \43407 );
xor \g456256/U$1_r2 ( \43638 , \43636 , \43637 );
xor \g456269/U$2 ( \43639 , \42977 , \42984 );
xor \g456269/U$1 ( \43640 , \43639 , \42992 );
xor \g456269/U$1_r1 ( \43641 , \43061 , \43066 );
xor \g456269/U$1_r2 ( \43642 , \43640 , \43641 );
xor \g456182/U$5 ( \43643 , \43638 , \43642 );
xor \g133545/U$1 ( \43644 , \43164 , \43196 );
xor \g133545/U$1_r1 ( \43645 , \43644 , \43226 );
and \g456182/U$4 ( \43646 , \43643 , \43645 );
and \g456182/U$6 ( \43647 , \43638 , \43642 );
or \g456182/U$3 ( \43648 , \43646 , \43647 );
xor \g133303/U$4 ( \43649 , \43634 , \43648 );
xor \g456202/U$2 ( \43650 , \42950 , \42952 );
xor \g456202/U$1 ( \43651 , \43650 , \42955 );
xor \g456202/U$1_r1 ( \43652 , \43071 , \43229 );
xor \g456202/U$1_r2 ( \43653 , \43651 , \43652 );
and \g133303/U$3 ( \43654 , \43649 , \43653 );
and \g133303/U$5 ( \43655 , \43634 , \43648 );
or \g133303/U$2 ( \43656 , \43654 , \43655 );
xor \g133421/U$1 ( \43657 , \43434 , \43438 );
xor \g133421/U$1_r1 ( \43658 , \43657 , \43443 );
xor \g133214/U$4 ( \43659 , \43656 , \43658 );
xor \g456181/U$2 ( \43660 , \42948 , \42958 );
xor \g456181/U$1 ( \43661 , \43660 , \42963 );
xor \g456181/U$1_r1 ( \43662 , \43234 , \43421 );
xor \g456181/U$1_r2 ( \43663 , \43661 , \43662 );
and \g133214/U$3 ( \43664 , \43659 , \43663 );
and \g133214/U$5 ( \43665 , \43656 , \43658 );
or \g133214/U$2 ( \43666 , \43664 , \43665 );
and \g131283/U$2 ( \43667 , \43459 , \43666 );
xor \g133184/U$1 ( \43668 , \43666 , \43459 );
xor \g456243/U$2 ( \43669 , \43321 , \43328 );
xor \g456243/U$1 ( \43670 , \43669 , \43336 );
xor \g456243/U$1_r1 ( \43671 , \43314 , \43360 );
xor \g456243/U$1_r2 ( \43672 , \43670 , \43671 );
xor \g456203/U$9 ( \43673 , \43239 , \43262 );
xor \g456203/U$9_r1 ( \43674 , \43673 , \43286 );
and \g456203/U$8 ( \43675 , \43672 , \43674 );
xor \g134017/U$1 ( \43676 , \43466 , \43473 );
xor \g134017/U$1_r1 ( \43677 , \43676 , \43481 );
xor \g456249/U$9 ( \43678 , \43546 , \43553 );
xor \g456249/U$9_r1 ( \43679 , \43678 , \43561 );
and \g456249/U$8 ( \43680 , \43677 , \43679 );
xor \g133913/U$1 ( \43681 , \43572 , \43579 );
xor \g133913/U$1_r1 ( \43682 , \43681 , \43587 );
xor \g456249/U$11 ( \43683 , \43546 , \43553 );
xor \g456249/U$11_r1 ( \43684 , \43683 , \43561 );
and \g456249/U$10 ( \43685 , \43682 , \43684 );
and \g456249/U$12 ( \43686 , \43677 , \43682 );
or \g456249/U$7 ( \43687 , \43680 , \43685 , \43686 );
xor \g456227/U$9 ( \43688 , \43600 , \42675 );
xor \g456227/U$9_r1 ( \43689 , \43688 , \43619 );
and \g456227/U$8 ( \43690 , \43687 , \43689 );
xor \g133725/U$1 ( \43691 , \43539 , \43564 );
xor \g133725/U$1_r1 ( \43692 , \43691 , \43590 );
xor \g456227/U$11 ( \43693 , \43600 , \42675 );
xor \g456227/U$11_r1 ( \43694 , \43693 , \43619 );
and \g456227/U$10 ( \43695 , \43692 , \43694 );
and \g456227/U$12 ( \43696 , \43687 , \43692 );
or \g456227/U$7 ( \43697 , \43690 , \43695 , \43696 );
xor \g456203/U$11 ( \43698 , \43239 , \43262 );
xor \g456203/U$11_r1 ( \43699 , \43698 , \43286 );
and \g456203/U$10 ( \43700 , \43697 , \43699 );
and \g456203/U$12 ( \43701 , \43672 , \43697 );
or \g456203/U$7 ( \43702 , \43675 , \43700 , \43701 );
xor \g456182/U$9 ( \43703 , \43638 , \43642 );
xor \g456182/U$9_r1 ( \43704 , \43703 , \43645 );
and \g456182/U$8 ( \43705 , \43702 , \43704 );
and \g134914/U$2 ( \43706 , \40513 , \41629 );
and \g134914/U$3 ( \43707 , \41345 , \40713 );
nor \g134914/U$1 ( \43708 , \43706 , \43707 );
and \g134490/U$2 ( \43709 , \43708 , \40521 );
not \g134490/U$4 ( \43710 , \43708 );
and \g134490/U$3 ( \43711 , \43710 , \40518 );
nor \g134490/U$1 ( \43712 , \43709 , \43711 );
and \g134790/U$2 ( \43713 , \42644 , \40189 );
and \g134790/U$3 ( \43714 , \40138 , \42643 );
nor \g134790/U$1 ( \43715 , \43713 , \43714 );
and \g134443/U$2 ( \43716 , \43715 , \42487 );
not \g134443/U$4 ( \43717 , \43715 );
and \g134443/U$3 ( \43718 , \43717 , \42486 );
nor \g134443/U$1 ( \43719 , \43716 , \43718 );
xor \g133908/U$4 ( \43720 , \43712 , \43719 );
and \g134890/U$2 ( \43721 , \40672 , \41116 );
and \g134890/U$3 ( \43722 , \41107 , \40858 );
nor \g134890/U$1 ( \43723 , \43721 , \43722 );
and \g134248/U$2 ( \43724 , \43723 , \40678 );
not \g134248/U$4 ( \43725 , \43723 );
and \g134248/U$3 ( \43726 , \43725 , \40677 );
nor \g134248/U$1 ( \43727 , \43724 , \43726 );
and \g133908/U$3 ( \43728 , \43720 , \43727 );
and \g133908/U$5 ( \43729 , \43712 , \43719 );
or \g133908/U$2 ( \43730 , \43728 , \43729 );
and \g134780/U$2 ( \43731 , \41206 , \40956 );
and \g134780/U$3 ( \43732 , \40926 , \41208 );
nor \g134780/U$1 ( \43733 , \43731 , \43732 );
and \g134545/U$2 ( \43734 , \43733 , \41215 );
not \g134545/U$4 ( \43735 , \43733 );
and \g134545/U$3 ( \43736 , \43735 , \41214 );
nor \g134545/U$1 ( \43737 , \43734 , \43736 );
and \g134693/U$2 ( \43738 , \41948 , \40472 );
and \g134693/U$3 ( \43739 , \40353 , \41947 );
nor \g134693/U$1 ( \43740 , \43738 , \43739 );
and \g134537/U$2 ( \43741 , \43740 , \41755 );
not \g134537/U$4 ( \43742 , \43740 );
and \g134537/U$3 ( \43743 , \43742 , \41952 );
nor \g134537/U$1 ( \43744 , \43741 , \43743 );
xor \g456261/U$5 ( \43745 , \43737 , \43744 );
and \g134934/U$2 ( \43746 , \40979 , \41109 );
and \g134934/U$3 ( \43747 , \41144 , \41071 );
nor \g134934/U$1 ( \43748 , \43746 , \43747 );
and \g134220/U$2 ( \43749 , \43748 , \40871 );
not \g134220/U$4 ( \43750 , \43748 );
and \g134220/U$3 ( \43751 , \43750 , \40870 );
nor \g134220/U$1 ( \43752 , \43749 , \43751 );
and \g456261/U$4 ( \43753 , \43745 , \43752 );
and \g456261/U$6 ( \43754 , \43737 , \43744 );
or \g456261/U$3 ( \43755 , \43753 , \43754 );
xor \g133787/U$4 ( \43756 , \43730 , \43755 );
not \g135489/U$1 ( \43757 , \43607 );
and \g134991/U$2 ( \43758 , \40091 , \43757 );
and \g134991/U$3 ( \43759 , \43179 , \40113 );
nor \g134991/U$1 ( \43760 , \43758 , \43759 );
and \g134188/U$2 ( \43761 , \43760 , \40080 );
not \g134188/U$4 ( \43762 , \43760 );
and \g134188/U$3 ( \43763 , \43762 , \40079 );
nor \g134188/U$1 ( \43764 , \43761 , \43763 );
and \g134754/U$2 ( \43765 , \42317 , \40307 );
and \g134754/U$3 ( \43766 , \40278 , \42316 );
nor \g134754/U$1 ( \43767 , \43765 , \43766 );
and \g134240/U$2 ( \43768 , \43767 , \42226 );
not \g134240/U$4 ( \43769 , \43767 );
and \g134240/U$3 ( \43770 , \43769 , \42225 );
nor \g134240/U$1 ( \43771 , \43768 , \43770 );
xor \g133961/U$4 ( \43772 , \43764 , \43771 );
and \g135060/U$2 ( \43773 , \43099 , \40158 );
and \g135060/U$3 ( \43774 , \40108 , \43101 );
nor \g135060/U$1 ( \43775 , \43773 , \43774 );
and \g134534/U$2 ( \43776 , \43775 , \42682 );
not \g134534/U$4 ( \43777 , \43775 );
and \g134534/U$3 ( \43778 , \43777 , \42681 );
nor \g134534/U$1 ( \43779 , \43776 , \43778 );
and \g133961/U$3 ( \43780 , \43772 , \43779 );
and \g133961/U$5 ( \43781 , \43764 , \43771 );
or \g133961/U$2 ( \43782 , \43780 , \43781 );
and \g133787/U$3 ( \43783 , \43756 , \43782 );
and \g133787/U$5 ( \43784 , \43730 , \43755 );
or \g133787/U$2 ( \43785 , \43783 , \43784 );
and \g134980/U$2 ( \43786 , \40175 , \42609 );
and \g134980/U$3 ( \43787 , \42416 , \40207 );
nor \g134980/U$1 ( \43788 , \43786 , \43787 );
and \g134178/U$2 ( \43789 , \43788 , \40137 );
not \g134178/U$4 ( \43790 , \43788 );
and \g134178/U$3 ( \43791 , \43790 , \40136 );
nor \g134178/U$1 ( \43792 , \43789 , \43791 );
nor \g135205/U$1 ( \43793 , \40085 , \43607 );
nor \g135160/U$1 ( \43794 , \43793 , \40080 );
and \g135304/U$2 ( \43795 , \43604 , \40067 );
and \g135304/U$3 ( \43796 , \40064 , \43603 );
nor \g135304/U$1 ( \43797 , \43795 , \43796 );
and \g135186/U$2 ( \43798 , \43797 , \42676 );
not \g135186/U$4 ( \43799 , \43797 );
and \g135186/U$3 ( \43800 , \43799 , \42675 );
nor \g135186/U$1 ( \43801 , \43798 , \43800 );
and \g134626/U$2 ( \43802 , \43794 , \43801 );
xor \g133955/U$4 ( \43803 , \43792 , \43802 );
and \g134689/U$2 ( \43804 , \40147 , \42701 );
and \g134689/U$3 ( \43805 , \42651 , \40149 );
nor \g134689/U$1 ( \43806 , \43804 , \43805 );
and \g134330/U$2 ( \43807 , \43806 , \40107 );
not \g134330/U$4 ( \43808 , \43806 );
and \g134330/U$3 ( \43809 , \43808 , \40106 );
nor \g134330/U$1 ( \43810 , \43807 , \43809 );
and \g133955/U$3 ( \43811 , \43803 , \43810 );
and \g133955/U$5 ( \43812 , \43792 , \43802 );
or \g133955/U$2 ( \43813 , \43811 , \43812 );
xor \g456201/U$5 ( \43814 , \43785 , \43813 );
and \g134719/U$2 ( \43815 , \40301 , \42416 );
and \g134719/U$3 ( \43816 , \42344 , \40391 );
nor \g134719/U$1 ( \43817 , \43815 , \43816 );
or \g134152/U$2 ( \43818 , \43817 , \40219 );
nand \g134630/U$1 ( \43819 , \40219 , \43817 );
nand \g134152/U$1 ( \43820 , \43818 , \43819 );
and \g134782/U$2 ( \43821 , \41623 , \40568 );
and \g134782/U$3 ( \43822 , \40525 , \41745 );
nor \g134782/U$1 ( \43823 , \43821 , \43822 );
and \g134187/U$2 ( \43824 , \43823 , \41325 );
not \g134187/U$4 ( \43825 , \43823 );
and \g134187/U$3 ( \43826 , \43825 , \41324 );
nor \g134187/U$1 ( \43827 , \43824 , \43826 );
xor \g456212/U$5 ( \43828 , \43820 , \43827 );
and \g134848/U$2 ( \43829 , \40432 , \41920 );
and \g134848/U$3 ( \43830 , \41774 , \40530 );
nor \g134848/U$1 ( \43831 , \43829 , \43830 );
and \g134410/U$2 ( \43832 , \43831 , \40388 );
not \g134410/U$4 ( \43833 , \43831 );
and \g134410/U$3 ( \43834 , \43833 , \40387 );
nor \g134410/U$1 ( \43835 , \43832 , \43834 );
and \g456212/U$4 ( \43836 , \43828 , \43835 );
and \g456212/U$6 ( \43837 , \43820 , \43827 );
or \g456212/U$3 ( \43838 , \43836 , \43837 );
and \g135033/U$2 ( \43839 , \40175 , \42651 );
and \g135033/U$3 ( \43840 , \42609 , \40207 );
nor \g135033/U$1 ( \43841 , \43839 , \43840 );
and \g134261/U$2 ( \43842 , \43841 , \40137 );
not \g134261/U$4 ( \43843 , \43841 );
and \g134261/U$3 ( \43844 , \43843 , \40136 );
nor \g134261/U$1 ( \43845 , \43842 , \43844 );
and \g135081/U$2 ( \43846 , \41087 , \40800 );
and \g135081/U$3 ( \43847 , \40731 , \41328 );
nor \g135081/U$1 ( \43848 , \43846 , \43847 );
and \g134327/U$2 ( \43849 , \43848 , \41093 );
not \g134327/U$4 ( \43850 , \43848 );
and \g134327/U$3 ( \43851 , \43850 , \41092 );
nor \g134327/U$1 ( \43852 , \43849 , \43851 );
xor \g133948/U$4 ( \43853 , \43845 , \43852 );
and \g135008/U$2 ( \43854 , \40147 , \43183 );
and \g135008/U$3 ( \43855 , \42701 , \40149 );
nor \g135008/U$1 ( \43856 , \43854 , \43855 );
and \g134365/U$2 ( \43857 , \43856 , \40107 );
not \g134365/U$4 ( \43858 , \43856 );
and \g134365/U$3 ( \43859 , \43858 , \40106 );
nor \g134365/U$1 ( \43860 , \43857 , \43859 );
and \g133948/U$3 ( \43861 , \43853 , \43860 );
and \g133948/U$5 ( \43862 , \43845 , \43852 );
or \g133948/U$2 ( \43863 , \43861 , \43862 );
xor \g456224/U$5 ( \43864 , \43838 , \43863 );
xor \g134040/U$1 ( \43865 , \43606 , \43608 );
xor \g134040/U$1_r1 ( \43866 , \43865 , \43616 );
and \g456224/U$4 ( \43867 , \43864 , \43866 );
and \g456224/U$6 ( \43868 , \43838 , \43863 );
or \g456224/U$3 ( \43869 , \43867 , \43868 );
and \g456201/U$4 ( \43870 , \43814 , \43869 );
and \g456201/U$6 ( \43871 , \43785 , \43813 );
or \g456201/U$3 ( \43872 , \43870 , \43871 );
xor \g456196/U$9 ( \43873 , \43593 , \43622 );
xor \g456196/U$9_r1 ( \43874 , \43873 , \43625 );
and \g456196/U$8 ( \43875 , \43872 , \43874 );
xor \g456226/U$2 ( \43876 , \43170 , \42676 );
xor \g456226/U$1 ( \43877 , \43876 , \43193 );
xor \g456226/U$1_r1 ( \43878 , \43494 , \43509 );
xor \g456226/U$1_r2 ( \43879 , \43877 , \43878 );
xor \g456196/U$11 ( \43880 , \43593 , \43622 );
xor \g456196/U$11_r1 ( \43881 , \43880 , \43625 );
and \g456196/U$10 ( \43882 , \43879 , \43881 );
and \g456196/U$12 ( \43883 , \43872 , \43879 );
or \g456196/U$7 ( \43884 , \43875 , \43882 , \43883 );
xor \g456182/U$11 ( \43885 , \43638 , \43642 );
xor \g456182/U$11_r1 ( \43886 , \43885 , \43645 );
and \g456182/U$10 ( \43887 , \43884 , \43886 );
and \g456182/U$12 ( \43888 , \43702 , \43884 );
or \g456182/U$7 ( \43889 , \43705 , \43887 , \43888 );
xor \g456195/U$2 ( \43890 , \43387 , \43389 );
xor \g456195/U$1 ( \43891 , \43890 , \43394 );
xor \g456195/U$1_r1 ( \43892 , \43383 , \43416 );
xor \g456195/U$1_r2 ( \43893 , \43891 , \43892 );
xor \g133215/U$4 ( \43894 , \43889 , \43893 );
xor \g133303/U$1 ( \43895 , \43634 , \43648 );
xor \g133303/U$1_r1 ( \43896 , \43895 , \43653 );
and \g133215/U$3 ( \43897 , \43894 , \43896 );
and \g133215/U$5 ( \43898 , \43889 , \43893 );
or \g133215/U$2 ( \43899 , \43897 , \43898 );
not \g131337/U$3 ( \43900 , \43899 );
xor \g133214/U$1 ( \43901 , \43656 , \43658 );
xor \g133214/U$1_r1 ( \43902 , \43901 , \43663 );
not \g131337/U$4 ( \43903 , \43902 );
or \g131337/U$2 ( \43904 , \43900 , \43903 );
and \g135299/U$2 ( \43905 , \43604 , \40108 );
and \g135299/U$3 ( \43906 , \40067 , \43603 );
nor \g135299/U$1 ( \43907 , \43905 , \43906 );
and \g135188/U$2 ( \43908 , \43907 , \42676 );
not \g135188/U$4 ( \43909 , \43907 );
and \g135188/U$3 ( \43910 , \43909 , \42675 );
nor \g135188/U$1 ( \43911 , \43908 , \43910 );
xor \g133970/U$4 ( \43912 , \43911 , \43793 );
and \g134799/U$2 ( \43913 , \43099 , \40138 );
and \g134799/U$3 ( \43914 , \40158 , \43101 );
nor \g134799/U$1 ( \43915 , \43913 , \43914 );
and \g134416/U$2 ( \43916 , \43915 , \42682 );
not \g134416/U$4 ( \43917 , \43915 );
and \g134416/U$3 ( \43918 , \43917 , \42681 );
nor \g134416/U$1 ( \43919 , \43916 , \43918 );
and \g133970/U$3 ( \43920 , \43912 , \43919 );
and \g133970/U$5 ( \43921 , \43911 , \43793 );
or \g133970/U$2 ( \43922 , \43920 , \43921 );
xor \g134626/U$1 ( \43923 , \43794 , \43801 );
xor \g133746/U$4 ( \43924 , \43922 , \43923 );
and \g134847/U$2 ( \43925 , \40979 , \41107 );
and \g134847/U$3 ( \43926 , \41109 , \41071 );
nor \g134847/U$1 ( \43927 , \43925 , \43926 );
or \g134163/U$2 ( \43928 , \43927 , \40870 );
nand \g134639/U$1 ( \43929 , \40870 , \43927 );
nand \g134163/U$1 ( \43930 , \43928 , \43929 );
and \g135035/U$2 ( \43931 , \42317 , \40353 );
and \g135035/U$3 ( \43932 , \40307 , \42316 );
nor \g135035/U$1 ( \43933 , \43931 , \43932 );
and \g134478/U$2 ( \43934 , \43933 , \42226 );
not \g134478/U$4 ( \43935 , \43933 );
and \g134478/U$3 ( \43936 , \43935 , \42225 );
nor \g134478/U$1 ( \43937 , \43934 , \43936 );
xor \g456241/U$5 ( \43938 , \43930 , \43937 );
and \g134700/U$2 ( \43939 , \41206 , \41144 );
and \g134700/U$3 ( \43940 , \40956 , \41208 );
nor \g134700/U$1 ( \43941 , \43939 , \43940 );
and \g134479/U$2 ( \43942 , \43941 , \41215 );
not \g134479/U$4 ( \43943 , \43941 );
and \g134479/U$3 ( \43944 , \43943 , \41214 );
nor \g134479/U$1 ( \43945 , \43942 , \43944 );
and \g456241/U$4 ( \43946 , \43938 , \43945 );
and \g456241/U$6 ( \43947 , \43930 , \43937 );
or \g456241/U$3 ( \43948 , \43946 , \43947 );
and \g133746/U$3 ( \43949 , \43924 , \43948 );
and \g133746/U$5 ( \43950 , \43922 , \43923 );
or \g133746/U$2 ( \43951 , \43949 , \43950 );
xor \g456224/U$9 ( \43952 , \43838 , \43863 );
xor \g456224/U$9_r1 ( \43953 , \43952 , \43866 );
and \g456224/U$8 ( \43954 , \43951 , \43953 );
xor \g133948/U$1 ( \43955 , \43845 , \43852 );
xor \g133948/U$1_r1 ( \43956 , \43955 , \43860 );
xor \g456261/U$9 ( \43957 , \43737 , \43744 );
xor \g456261/U$9_r1 ( \43958 , \43957 , \43752 );
and \g456261/U$8 ( \43959 , \43956 , \43958 );
xor \g133961/U$1 ( \43960 , \43764 , \43771 );
xor \g133961/U$1_r1 ( \43961 , \43960 , \43779 );
xor \g456261/U$11 ( \43962 , \43737 , \43744 );
xor \g456261/U$11_r1 ( \43963 , \43962 , \43752 );
and \g456261/U$10 ( \43964 , \43961 , \43963 );
and \g456261/U$12 ( \43965 , \43956 , \43961 );
or \g456261/U$7 ( \43966 , \43959 , \43964 , \43965 );
xor \g456224/U$11 ( \43967 , \43838 , \43863 );
xor \g456224/U$11_r1 ( \43968 , \43967 , \43866 );
and \g456224/U$10 ( \43969 , \43966 , \43968 );
and \g456224/U$12 ( \43970 , \43951 , \43966 );
or \g456224/U$7 ( \43971 , \43954 , \43969 , \43970 );
xor \g456201/U$9 ( \43972 , \43785 , \43813 );
xor \g456201/U$9_r1 ( \43973 , \43972 , \43869 );
and \g456201/U$8 ( \43974 , \43971 , \43973 );
xor \g456227/U$2 ( \43975 , \43600 , \42675 );
xor \g456227/U$1 ( \43976 , \43975 , \43619 );
xor \g456227/U$1_r1 ( \43977 , \43687 , \43692 );
xor \g456227/U$1_r2 ( \43978 , \43976 , \43977 );
xor \g456201/U$11 ( \43979 , \43785 , \43813 );
xor \g456201/U$11_r1 ( \43980 , \43979 , \43869 );
and \g456201/U$10 ( \43981 , \43978 , \43980 );
and \g456201/U$12 ( \43982 , \43971 , \43978 );
or \g456201/U$7 ( \43983 , \43974 , \43981 , \43982 );
xor \g133957/U$1 ( \43984 , \43521 , \43528 );
xor \g133957/U$1_r1 ( \43985 , \43984 , \43536 );
xor \g133955/U$1 ( \43986 , \43792 , \43802 );
xor \g133955/U$1_r1 ( \43987 , \43986 , \43810 );
xor \g456199/U$5 ( \43988 , \43985 , \43987 );
and \g134840/U$2 ( \43989 , \40175 , \42701 );
and \g134840/U$3 ( \43990 , \42651 , \40207 );
nor \g134840/U$1 ( \43991 , \43989 , \43990 );
and \g134524/U$2 ( \43992 , \43991 , \40137 );
not \g134524/U$4 ( \43993 , \43991 );
and \g134524/U$3 ( \43994 , \43993 , \40136 );
nor \g134524/U$1 ( \43995 , \43992 , \43994 );
and \g134874/U$2 ( \43996 , \41087 , \40926 );
and \g134874/U$3 ( \43997 , \40800 , \41328 );
nor \g134874/U$1 ( \43998 , \43996 , \43997 );
and \g134260/U$2 ( \43999 , \43998 , \41093 );
not \g134260/U$4 ( \44000 , \43998 );
and \g134260/U$3 ( \44001 , \44000 , \41092 );
nor \g134260/U$1 ( \44002 , \43999 , \44001 );
xor \g456247/U$5 ( \44003 , \43995 , \44002 );
and \g134977/U$2 ( \44004 , \40301 , \42609 );
and \g134977/U$3 ( \44005 , \42416 , \40391 );
nor \g134977/U$1 ( \44006 , \44004 , \44005 );
and \g134349/U$2 ( \44007 , \44006 , \40220 );
not \g134349/U$4 ( \44008 , \44006 );
and \g134349/U$3 ( \44009 , \44008 , \40219 );
nor \g134349/U$1 ( \44010 , \44007 , \44009 );
and \g456247/U$4 ( \44011 , \44003 , \44010 );
and \g456247/U$6 ( \44012 , \43995 , \44002 );
or \g456247/U$3 ( \44013 , \44011 , \44012 );
and \g134836/U$2 ( \44014 , \40513 , \41774 );
and \g134836/U$3 ( \44015 , \41629 , \40713 );
nor \g134836/U$1 ( \44016 , \44014 , \44015 );
and \g134224/U$2 ( \44017 , \44016 , \40521 );
not \g134224/U$4 ( \44018 , \44016 );
and \g134224/U$3 ( \44019 , \44018 , \40518 );
nor \g134224/U$1 ( \44020 , \44017 , \44019 );
and \g135069/U$2 ( \44021 , \41948 , \40525 );
and \g135069/U$3 ( \44022 , \40472 , \41947 );
nor \g135069/U$1 ( \44023 , \44021 , \44022 );
and \g134396/U$2 ( \44024 , \44023 , \41755 );
not \g134396/U$4 ( \44025 , \44023 );
and \g134396/U$3 ( \44026 , \44025 , \41952 );
nor \g134396/U$1 ( \44027 , \44024 , \44026 );
xor \g133922/U$4 ( \44028 , \44020 , \44027 );
and \g134961/U$2 ( \44029 , \40672 , \41345 );
and \g134961/U$3 ( \44030 , \41116 , \40858 );
nor \g134961/U$1 ( \44031 , \44029 , \44030 );
and \g134262/U$2 ( \44032 , \44031 , \40678 );
not \g134262/U$4 ( \44033 , \44031 );
and \g134262/U$3 ( \44034 , \44033 , \40677 );
nor \g134262/U$1 ( \44035 , \44032 , \44034 );
and \g133922/U$3 ( \44036 , \44028 , \44035 );
and \g133922/U$5 ( \44037 , \44020 , \44027 );
or \g133922/U$2 ( \44038 , \44036 , \44037 );
xor \g133744/U$4 ( \44039 , \44013 , \44038 );
and \g134722/U$2 ( \44040 , \42644 , \40278 );
and \g134722/U$3 ( \44041 , \40189 , \42643 );
nor \g134722/U$1 ( \44042 , \44040 , \44041 );
and \g134317/U$2 ( \44043 , \44042 , \42487 );
not \g134317/U$4 ( \44044 , \44042 );
and \g134317/U$3 ( \44045 , \44044 , \42486 );
nor \g134317/U$1 ( \44046 , \44043 , \44045 );
and \g135103/U$2 ( \44047 , \41623 , \40731 );
and \g135103/U$3 ( \44048 , \40568 , \41745 );
nor \g135103/U$1 ( \44049 , \44047 , \44048 );
and \g134592/U$2 ( \44050 , \44049 , \41325 );
not \g134592/U$4 ( \44051 , \44049 );
and \g134592/U$3 ( \44052 , \44051 , \41324 );
nor \g134592/U$1 ( \44053 , \44050 , \44052 );
xor \g133979/U$4 ( \44054 , \44046 , \44053 );
and \g134773/U$2 ( \44055 , \40432 , \42344 );
and \g134773/U$3 ( \44056 , \41920 , \40530 );
nor \g134773/U$1 ( \44057 , \44055 , \44056 );
and \g134622/U$2 ( \44058 , \44057 , \40388 );
not \g134622/U$4 ( \44059 , \44057 );
and \g134622/U$3 ( \44060 , \44059 , \40387 );
nor \g134622/U$1 ( \44061 , \44058 , \44060 );
and \g133979/U$3 ( \44062 , \44054 , \44061 );
and \g133979/U$5 ( \44063 , \44046 , \44053 );
or \g133979/U$2 ( \44064 , \44062 , \44063 );
and \g133744/U$3 ( \44065 , \44039 , \44064 );
and \g133744/U$5 ( \44066 , \44013 , \44038 );
or \g133744/U$2 ( \44067 , \44065 , \44066 );
and \g456199/U$4 ( \44068 , \43988 , \44067 );
and \g456199/U$6 ( \44069 , \43985 , \43987 );
or \g456199/U$3 ( \44070 , \44068 , \44069 );
xor \g456251/U$2 ( \44071 , \43296 , \43303 );
xor \g456251/U$1 ( \44072 , \44071 , \43311 );
xor \g456251/U$1_r1 ( \44073 , \43484 , \43489 );
xor \g456251/U$1_r2 ( \44074 , \44072 , \44073 );
xor \g456179/U$5 ( \44075 , \44070 , \44074 );
xor \g456246/U$2 ( \44076 , \43143 , \43150 );
xor \g456246/U$1 ( \44077 , \44076 , \43158 );
xor \g456246/U$1_r1 ( \44078 , \43499 , \43504 );
xor \g456246/U$1_r2 ( \44079 , \44077 , \44078 );
and \g456179/U$4 ( \44080 , \44075 , \44079 );
and \g456179/U$6 ( \44081 , \44070 , \44074 );
or \g456179/U$3 ( \44082 , \44080 , \44081 );
xor \g133331/U$4 ( \44083 , \43983 , \44082 );
xor \g456203/U$2 ( \44084 , \43239 , \43262 );
xor \g456203/U$1 ( \44085 , \44084 , \43286 );
xor \g456203/U$1_r1 ( \44086 , \43672 , \43697 );
xor \g456203/U$1_r2 ( \44087 , \44085 , \44086 );
and \g133331/U$3 ( \44088 , \44083 , \44087 );
and \g133331/U$5 ( \44089 , \43983 , \44082 );
or \g133331/U$2 ( \44090 , \44088 , \44089 );
xor \g133400/U$1 ( \44091 , \43514 , \43628 );
xor \g133400/U$1_r1 ( \44092 , \44091 , \43631 );
xor \g133242/U$4 ( \44093 , \44090 , \44092 );
xor \g456182/U$2 ( \44094 , \43638 , \43642 );
xor \g456182/U$1 ( \44095 , \44094 , \43645 );
xor \g456182/U$1_r1 ( \44096 , \43702 , \43884 );
xor \g456182/U$1_r2 ( \44097 , \44095 , \44096 );
and \g133242/U$3 ( \44098 , \44093 , \44097 );
and \g133242/U$5 ( \44099 , \44090 , \44092 );
or \g133242/U$2 ( \44100 , \44098 , \44099 );
xor \g133215/U$1 ( \44101 , \43889 , \43893 );
xor \g133215/U$1_r1 ( \44102 , \44101 , \43896 );
and \g131394/U$2 ( \44103 , \44100 , \44102 );
xor \g133185/U$1 ( \44104 , \44102 , \44100 );
xor \g133242/U$1 ( \44105 , \44090 , \44092 );
xor \g133242/U$1_r1 ( \44106 , \44105 , \44097 );
xor \g456249/U$2 ( \44107 , \43546 , \43553 );
xor \g456249/U$1 ( \44108 , \44107 , \43561 );
xor \g456249/U$1_r1 ( \44109 , \43677 , \43682 );
xor \g456249/U$1_r2 ( \44110 , \44108 , \44109 );
xor \g133787/U$1 ( \44111 , \43730 , \43755 );
xor \g133787/U$1_r1 ( \44112 , \44111 , \43782 );
xor \g456177/U$5 ( \44113 , \44110 , \44112 );
xor \g133908/U$1 ( \44114 , \43712 , \43719 );
xor \g133908/U$1_r1 ( \44115 , \44114 , \43727 );
xor \g456212/U$9 ( \44116 , \43820 , \43827 );
xor \g456212/U$9_r1 ( \44117 , \44116 , \43835 );
and \g456212/U$8 ( \44118 , \44115 , \44117 );
and \g135012/U$2 ( \44119 , \40979 , \41116 );
and \g135012/U$3 ( \44120 , \41107 , \41071 );
nor \g135012/U$1 ( \44121 , \44119 , \44120 );
and \g134185/U$2 ( \44122 , \44121 , \40871 );
not \g134185/U$4 ( \44123 , \44121 );
and \g134185/U$3 ( \44124 , \44123 , \40870 );
nor \g134185/U$1 ( \44125 , \44122 , \44124 );
and \g135074/U$2 ( \44126 , \41948 , \40568 );
and \g135074/U$3 ( \44127 , \40525 , \41947 );
nor \g135074/U$1 ( \44128 , \44126 , \44127 );
and \g134363/U$2 ( \44129 , \44128 , \41755 );
not \g134363/U$4 ( \44130 , \44128 );
and \g134363/U$3 ( \44131 , \44130 , \41952 );
nor \g134363/U$1 ( \44132 , \44129 , \44131 );
xor \g133975/U$4 ( \44133 , \44125 , \44132 );
and \g134843/U$2 ( \44134 , \40672 , \41629 );
and \g134843/U$3 ( \44135 , \41345 , \40858 );
nor \g134843/U$1 ( \44136 , \44134 , \44135 );
and \g134314/U$2 ( \44137 , \44136 , \40678 );
not \g134314/U$4 ( \44138 , \44136 );
and \g134314/U$3 ( \44139 , \44138 , \40677 );
nor \g134314/U$1 ( \44140 , \44137 , \44139 );
and \g133975/U$3 ( \44141 , \44133 , \44140 );
and \g133975/U$5 ( \44142 , \44125 , \44132 );
or \g133975/U$2 ( \44143 , \44141 , \44142 );
and \g134749/U$2 ( \44144 , \40513 , \41920 );
and \g134749/U$3 ( \44145 , \41774 , \40713 );
nor \g134749/U$1 ( \44146 , \44144 , \44145 );
and \g134610/U$2 ( \44147 , \44146 , \40521 );
not \g134610/U$4 ( \44148 , \44146 );
and \g134610/U$3 ( \44149 , \44148 , \40518 );
nor \g134610/U$1 ( \44150 , \44147 , \44149 );
and \g134943/U$2 ( \44151 , \42644 , \40307 );
and \g134943/U$3 ( \44152 , \40278 , \42643 );
nor \g134943/U$1 ( \44153 , \44151 , \44152 );
and \g134621/U$2 ( \44154 , \44153 , \42487 );
not \g134621/U$4 ( \44155 , \44153 );
and \g134621/U$3 ( \44156 , \44155 , \42486 );
nor \g134621/U$1 ( \44157 , \44154 , \44156 );
xor \g456248/U$5 ( \44158 , \44150 , \44157 );
and \g134939/U$2 ( \44159 , \41623 , \40800 );
and \g134939/U$3 ( \44160 , \40731 , \41745 );
nor \g134939/U$1 ( \44161 , \44159 , \44160 );
and \g134474/U$2 ( \44162 , \44161 , \41325 );
not \g134474/U$4 ( \44163 , \44161 );
and \g134474/U$3 ( \44164 , \44163 , \41324 );
nor \g134474/U$1 ( \44165 , \44162 , \44164 );
and \g456248/U$4 ( \44166 , \44158 , \44165 );
and \g456248/U$6 ( \44167 , \44150 , \44157 );
or \g456248/U$3 ( \44168 , \44166 , \44167 );
xor \g133684/U$4 ( \44169 , \44143 , \44168 );
and \g134946/U$2 ( \44170 , \40301 , \42651 );
and \g134946/U$3 ( \44171 , \42609 , \40391 );
nor \g134946/U$1 ( \44172 , \44170 , \44171 );
and \g134157/U$2 ( \44173 , \44172 , \40220 );
not \g134157/U$4 ( \44174 , \44172 );
and \g134157/U$3 ( \44175 , \44174 , \40219 );
nor \g134157/U$1 ( \44176 , \44173 , \44175 );
and \g134967/U$2 ( \44177 , \41087 , \40956 );
and \g134967/U$3 ( \44178 , \40926 , \41328 );
nor \g134967/U$1 ( \44179 , \44177 , \44178 );
or \g134222/U$2 ( \44180 , \44179 , \41092 );
nand \g134638/U$1 ( \44181 , \41092 , \44179 );
nand \g134222/U$1 ( \44182 , \44180 , \44181 );
xor \g133924/U$4 ( \44183 , \44176 , \44182 );
and \g134762/U$2 ( \44184 , \40432 , \42416 );
and \g134762/U$3 ( \44185 , \42344 , \40530 );
nor \g134762/U$1 ( \44186 , \44184 , \44185 );
and \g134452/U$2 ( \44187 , \44186 , \40388 );
not \g134452/U$4 ( \44188 , \44186 );
and \g134452/U$3 ( \44189 , \44188 , \40387 );
nor \g134452/U$1 ( \44190 , \44187 , \44189 );
and \g133924/U$3 ( \44191 , \44183 , \44190 );
and \g133924/U$5 ( \44192 , \44176 , \44182 );
or \g133924/U$2 ( \44193 , \44191 , \44192 );
and \g133684/U$3 ( \44194 , \44169 , \44193 );
and \g133684/U$5 ( \44195 , \44143 , \44168 );
or \g133684/U$2 ( \44196 , \44194 , \44195 );
xor \g456212/U$11 ( \44197 , \43820 , \43827 );
xor \g456212/U$11_r1 ( \44198 , \44197 , \43835 );
and \g456212/U$10 ( \44199 , \44196 , \44198 );
and \g456212/U$12 ( \44200 , \44115 , \44196 );
or \g456212/U$7 ( \44201 , \44118 , \44199 , \44200 );
and \g456177/U$4 ( \44202 , \44113 , \44201 );
and \g456177/U$6 ( \44203 , \44110 , \44112 );
or \g456177/U$3 ( \44204 , \44202 , \44203 );
xor \g456179/U$9 ( \44205 , \44070 , \44074 );
xor \g456179/U$9_r1 ( \44206 , \44205 , \44079 );
and \g456179/U$8 ( \44207 , \44204 , \44206 );
xor \g133746/U$1 ( \44208 , \43922 , \43923 );
xor \g133746/U$1_r1 ( \44209 , \44208 , \43948 );
and \g134831/U$2 ( \44210 , \40147 , \43179 );
and \g134831/U$3 ( \44211 , \43183 , \40149 );
nor \g134831/U$1 ( \44212 , \44210 , \44211 );
and \g134475/U$2 ( \44213 , \44212 , \40107 );
not \g134475/U$4 ( \44214 , \44212 );
and \g134475/U$3 ( \44215 , \44214 , \40106 );
nor \g134475/U$1 ( \44216 , \44213 , \44215 );
nor \g135209/U$1 ( \44217 , \40142 , \43607 );
nor \g135173/U$1 ( \44218 , \44217 , \40107 );
and \g135289/U$2 ( \44219 , \43604 , \40158 );
and \g135289/U$3 ( \44220 , \40108 , \43603 );
nor \g135289/U$1 ( \44221 , \44219 , \44220 );
and \g135174/U$2 ( \44222 , \44221 , \42676 );
not \g135174/U$4 ( \44223 , \44221 );
and \g135174/U$3 ( \44224 , \44223 , \42675 );
nor \g135174/U$1 ( \44225 , \44222 , \44224 );
and \g134624/U$2 ( \44226 , \44218 , \44225 );
xor \g133774/U$4 ( \44227 , \44216 , \44226 );
and \g134696/U$2 ( \44228 , \41206 , \41109 );
and \g134696/U$3 ( \44229 , \41144 , \41208 );
nor \g134696/U$1 ( \44230 , \44228 , \44229 );
and \g134360/U$2 ( \44231 , \44230 , \41215 );
not \g134360/U$4 ( \44232 , \44230 );
and \g134360/U$3 ( \44233 , \44232 , \41214 );
nor \g134360/U$1 ( \44234 , \44231 , \44233 );
and \g135099/U$2 ( \44235 , \42317 , \40472 );
and \g135099/U$3 ( \44236 , \40353 , \42316 );
nor \g135099/U$1 ( \44237 , \44235 , \44236 );
and \g134489/U$2 ( \44238 , \44237 , \42226 );
not \g134489/U$4 ( \44239 , \44237 );
and \g134489/U$3 ( \44240 , \44239 , \42225 );
nor \g134489/U$1 ( \44241 , \44238 , \44240 );
xor \g134014/U$4 ( \44242 , \44234 , \44241 );
and \g134912/U$2 ( \44243 , \43099 , \40189 );
and \g134912/U$3 ( \44244 , \40138 , \43101 );
nor \g134912/U$1 ( \44245 , \44243 , \44244 );
and \g134329/U$2 ( \44246 , \44245 , \42682 );
not \g134329/U$4 ( \44247 , \44245 );
and \g134329/U$3 ( \44248 , \44247 , \42681 );
nor \g134329/U$1 ( \44249 , \44246 , \44248 );
and \g134014/U$3 ( \44250 , \44242 , \44249 );
and \g134014/U$5 ( \44251 , \44234 , \44241 );
or \g134014/U$2 ( \44252 , \44250 , \44251 );
and \g133774/U$3 ( \44253 , \44227 , \44252 );
and \g133774/U$5 ( \44254 , \44216 , \44226 );
or \g133774/U$2 ( \44255 , \44253 , \44254 );
xor \g456185/U$5 ( \44256 , \44209 , \44255 );
xor \g133744/U$1 ( \44257 , \44013 , \44038 );
xor \g133744/U$1_r1 ( \44258 , \44257 , \44064 );
and \g456185/U$4 ( \44259 , \44256 , \44258 );
and \g456185/U$6 ( \44260 , \44209 , \44255 );
or \g456185/U$3 ( \44261 , \44259 , \44260 );
xor \g456199/U$9 ( \44262 , \43985 , \43987 );
xor \g456199/U$9_r1 ( \44263 , \44262 , \44067 );
and \g456199/U$8 ( \44264 , \44261 , \44263 );
xor \g133979/U$1 ( \44265 , \44046 , \44053 );
xor \g133979/U$1_r1 ( \44266 , \44265 , \44061 );
xor \g456247/U$9 ( \44267 , \43995 , \44002 );
xor \g456247/U$9_r1 ( \44268 , \44267 , \44010 );
and \g456247/U$8 ( \44269 , \44266 , \44268 );
xor \g133970/U$1 ( \44270 , \43911 , \43793 );
xor \g133970/U$1_r1 ( \44271 , \44270 , \43919 );
xor \g456247/U$11 ( \44272 , \43995 , \44002 );
xor \g456247/U$11_r1 ( \44273 , \44272 , \44010 );
and \g456247/U$10 ( \44274 , \44271 , \44273 );
and \g456247/U$12 ( \44275 , \44266 , \44271 );
or \g456247/U$7 ( \44276 , \44269 , \44274 , \44275 );
and \g135137/U$2 ( \44277 , \40175 , \43183 );
and \g135137/U$3 ( \44278 , \42701 , \40207 );
nor \g135137/U$1 ( \44279 , \44277 , \44278 );
and \g134583/U$2 ( \44280 , \44279 , \40137 );
not \g134583/U$4 ( \44281 , \44279 );
and \g134583/U$3 ( \44282 , \44281 , \40136 );
nor \g134583/U$1 ( \44283 , \44280 , \44282 );
xor \g134624/U$1 ( \44284 , \44218 , \44225 );
xor \g133897/U$4 ( \44285 , \44283 , \44284 );
and \g134767/U$2 ( \44286 , \40147 , \43757 );
and \g134767/U$3 ( \44287 , \43179 , \40149 );
nor \g134767/U$1 ( \44288 , \44286 , \44287 );
and \g134504/U$2 ( \44289 , \44288 , \40107 );
not \g134504/U$4 ( \44290 , \44288 );
and \g134504/U$3 ( \44291 , \44290 , \40106 );
nor \g134504/U$1 ( \44292 , \44289 , \44291 );
and \g133897/U$3 ( \44293 , \44285 , \44292 );
and \g133897/U$5 ( \44294 , \44283 , \44284 );
or \g133897/U$2 ( \44295 , \44293 , \44294 );
xor \g456241/U$9 ( \44296 , \43930 , \43937 );
xor \g456241/U$9_r1 ( \44297 , \44296 , \43945 );
and \g456241/U$8 ( \44298 , \44295 , \44297 );
xor \g133922/U$1 ( \44299 , \44020 , \44027 );
xor \g133922/U$1_r1 ( \44300 , \44299 , \44035 );
xor \g456241/U$11 ( \44301 , \43930 , \43937 );
xor \g456241/U$11_r1 ( \44302 , \44301 , \43945 );
and \g456241/U$10 ( \44303 , \44300 , \44302 );
and \g456241/U$12 ( \44304 , \44295 , \44300 );
or \g456241/U$7 ( \44305 , \44298 , \44303 , \44304 );
xor \g133538/U$4 ( \44306 , \44276 , \44305 );
xor \g456261/U$2 ( \44307 , \43737 , \43744 );
xor \g456261/U$1 ( \44308 , \44307 , \43752 );
xor \g456261/U$1_r1 ( \44309 , \43956 , \43961 );
xor \g456261/U$1_r2 ( \44310 , \44308 , \44309 );
and \g133538/U$3 ( \44311 , \44306 , \44310 );
and \g133538/U$5 ( \44312 , \44276 , \44305 );
or \g133538/U$2 ( \44313 , \44311 , \44312 );
xor \g456199/U$11 ( \44314 , \43985 , \43987 );
xor \g456199/U$11_r1 ( \44315 , \44314 , \44067 );
and \g456199/U$10 ( \44316 , \44313 , \44315 );
and \g456199/U$12 ( \44317 , \44261 , \44313 );
or \g456199/U$7 ( \44318 , \44264 , \44316 , \44317 );
xor \g456179/U$11 ( \44319 , \44070 , \44074 );
xor \g456179/U$11_r1 ( \44320 , \44319 , \44079 );
and \g456179/U$10 ( \44321 , \44318 , \44320 );
and \g456179/U$12 ( \44322 , \44204 , \44318 );
or \g456179/U$7 ( \44323 , \44207 , \44321 , \44322 );
xor \g456196/U$2 ( \44324 , \43593 , \43622 );
xor \g456196/U$1 ( \44325 , \44324 , \43625 );
xor \g456196/U$1_r1 ( \44326 , \43872 , \43879 );
xor \g456196/U$1_r2 ( \44327 , \44325 , \44326 );
xor \g133218/U$4 ( \44328 , \44323 , \44327 );
xor \g133331/U$1 ( \44329 , \43983 , \44082 );
xor \g133331/U$1_r1 ( \44330 , \44329 , \44087 );
and \g133218/U$3 ( \44331 , \44328 , \44330 );
and \g133218/U$5 ( \44332 , \44323 , \44327 );
or \g133218/U$2 ( \44333 , \44331 , \44332 );
and \g131466/U$2 ( \44334 , \44106 , \44333 );
xor \g133178/U$1 ( \44335 , \44333 , \44106 );
xor \g456224/U$2 ( \44336 , \43838 , \43863 );
xor \g456224/U$1 ( \44337 , \44336 , \43866 );
xor \g456224/U$1_r1 ( \44338 , \43951 , \43966 );
xor \g456224/U$1_r2 ( \44339 , \44337 , \44338 );
xor \g456177/U$9 ( \44340 , \44110 , \44112 );
xor \g456177/U$9_r1 ( \44341 , \44340 , \44201 );
and \g456177/U$8 ( \44342 , \44339 , \44341 );
xor \g456199/U$2 ( \44343 , \43985 , \43987 );
xor \g456199/U$1 ( \44344 , \44343 , \44067 );
xor \g456199/U$1_r1 ( \44345 , \44261 , \44313 );
xor \g456199/U$1_r2 ( \44346 , \44344 , \44345 );
xor \g456177/U$11 ( \44347 , \44110 , \44112 );
xor \g456177/U$11_r1 ( \44348 , \44347 , \44201 );
and \g456177/U$10 ( \44349 , \44346 , \44348 );
and \g456177/U$12 ( \44350 , \44339 , \44346 );
or \g456177/U$7 ( \44351 , \44342 , \44349 , \44350 );
xor \g456201/U$2 ( \44352 , \43785 , \43813 );
xor \g456201/U$1 ( \44353 , \44352 , \43869 );
xor \g456201/U$1_r1 ( \44354 , \43971 , \43978 );
xor \g456201/U$1_r2 ( \44355 , \44353 , \44354 );
xor \g133211/U$4 ( \44356 , \44351 , \44355 );
xor \g456179/U$2 ( \44357 , \44070 , \44074 );
xor \g456179/U$1 ( \44358 , \44357 , \44079 );
xor \g456179/U$1_r1 ( \44359 , \44204 , \44318 );
xor \g456179/U$1_r2 ( \44360 , \44358 , \44359 );
and \g133211/U$3 ( \44361 , \44356 , \44360 );
and \g133211/U$5 ( \44362 , \44351 , \44355 );
or \g133211/U$2 ( \44363 , \44361 , \44362 );
xor \g133218/U$1 ( \44364 , \44323 , \44327 );
xor \g133218/U$1_r1 ( \44365 , \44364 , \44330 );
and \g131534/U$2 ( \44366 , \44363 , \44365 );
xor \g133176/U$1 ( \44367 , \44365 , \44363 );
xor \g133538/U$1 ( \44368 , \44276 , \44305 );
xor \g133538/U$1_r1 ( \44369 , \44368 , \44310 );
xor \g456185/U$9 ( \44370 , \44209 , \44255 );
xor \g456185/U$9_r1 ( \44371 , \44370 , \44258 );
and \g456185/U$8 ( \44372 , \44369 , \44371 );
and \g134958/U$2 ( \44373 , \40979 , \41629 );
and \g134958/U$3 ( \44374 , \41345 , \41071 );
nor \g134958/U$1 ( \44375 , \44373 , \44374 );
and \g134369/U$2 ( \44376 , \44375 , \40871 );
not \g134369/U$4 ( \44377 , \44375 );
and \g134369/U$3 ( \44378 , \44377 , \40870 );
nor \g134369/U$1 ( \44379 , \44376 , \44378 );
and \g134893/U$2 ( \44380 , \42317 , \40568 );
and \g134893/U$3 ( \44381 , \40525 , \42316 );
nor \g134893/U$1 ( \44382 , \44380 , \44381 );
and \g134321/U$2 ( \44383 , \44382 , \42226 );
not \g134321/U$4 ( \44384 , \44382 );
and \g134321/U$3 ( \44385 , \44384 , \42225 );
nor \g134321/U$1 ( \44386 , \44383 , \44385 );
xor \g133923/U$4 ( \44387 , \44379 , \44386 );
and \g134880/U$2 ( \44388 , \41206 , \41116 );
and \g134880/U$3 ( \44389 , \41107 , \41208 );
nor \g134880/U$1 ( \44390 , \44388 , \44389 );
and \g134205/U$2 ( \44391 , \44390 , \41215 );
not \g134205/U$4 ( \44392 , \44390 );
and \g134205/U$3 ( \44393 , \44392 , \41214 );
nor \g134205/U$1 ( \44394 , \44391 , \44393 );
and \g133923/U$3 ( \44395 , \44387 , \44394 );
and \g133923/U$5 ( \44396 , \44379 , \44386 );
or \g133923/U$2 ( \44397 , \44395 , \44396 );
nor \g135207/U$1 ( \44398 , \40169 , \43607 );
nor \g135165/U$1 ( \44399 , \44398 , \40137 );
and \g134937/U$2 ( \44400 , \43099 , \40307 );
and \g134937/U$3 ( \44401 , \40278 , \43101 );
nor \g134937/U$1 ( \44402 , \44400 , \44401 );
and \g134401/U$2 ( \44403 , \44402 , \42682 );
not \g134401/U$4 ( \44404 , \44402 );
and \g134401/U$3 ( \44405 , \44404 , \42681 );
nor \g134401/U$1 ( \44406 , \44403 , \44405 );
and \g134090/U$2 ( \44407 , \44399 , \44406 );
xor \g133689/U$4 ( \44408 , \44397 , \44407 );
and \g135028/U$2 ( \44409 , \40513 , \42416 );
and \g135028/U$3 ( \44410 , \42344 , \40713 );
nor \g135028/U$1 ( \44411 , \44409 , \44410 );
and \g134354/U$2 ( \44412 , \44411 , \40521 );
not \g134354/U$4 ( \44413 , \44411 );
and \g134354/U$3 ( \44414 , \44413 , \40518 );
nor \g134354/U$1 ( \44415 , \44412 , \44414 );
and \g135102/U$2 ( \44416 , \41948 , \40800 );
and \g135102/U$3 ( \44417 , \40731 , \41947 );
nor \g135102/U$1 ( \44418 , \44416 , \44417 );
and \g134484/U$2 ( \44419 , \44418 , \41755 );
not \g134484/U$4 ( \44420 , \44418 );
and \g134484/U$3 ( \44421 , \44420 , \41952 );
nor \g134484/U$1 ( \44422 , \44419 , \44421 );
xor \g133910/U$4 ( \44423 , \44415 , \44422 );
and \g135025/U$2 ( \44424 , \40672 , \41920 );
and \g135025/U$3 ( \44425 , \41774 , \40858 );
nor \g135025/U$1 ( \44426 , \44424 , \44425 );
and \g134446/U$2 ( \44427 , \44426 , \40678 );
not \g134446/U$4 ( \44428 , \44426 );
and \g134446/U$3 ( \44429 , \44428 , \40677 );
nor \g134446/U$1 ( \44430 , \44427 , \44429 );
and \g133910/U$3 ( \44431 , \44423 , \44430 );
and \g133910/U$5 ( \44432 , \44415 , \44422 );
or \g133910/U$2 ( \44433 , \44431 , \44432 );
and \g133689/U$3 ( \44434 , \44408 , \44433 );
and \g133689/U$5 ( \44435 , \44397 , \44407 );
or \g133689/U$2 ( \44436 , \44434 , \44435 );
xor \g133897/U$1 ( \44437 , \44283 , \44284 );
xor \g133897/U$1_r1 ( \44438 , \44437 , \44292 );
xor \g456192/U$5 ( \44439 , \44436 , \44438 );
and \g134908/U$2 ( \44440 , \42644 , \40353 );
and \g134908/U$3 ( \44441 , \40307 , \42643 );
nor \g134908/U$1 ( \44442 , \44440 , \44441 );
and \g134196/U$2 ( \44443 , \44442 , \42487 );
not \g134196/U$4 ( \44444 , \44442 );
and \g134196/U$3 ( \44445 , \44444 , \42486 );
nor \g134196/U$1 ( \44446 , \44443 , \44445 );
and \g135094/U$2 ( \44447 , \41087 , \41144 );
and \g135094/U$3 ( \44448 , \40956 , \41328 );
nor \g135094/U$1 ( \44449 , \44447 , \44448 );
and \g134399/U$2 ( \44450 , \44449 , \41093 );
not \g134399/U$4 ( \44451 , \44449 );
and \g134399/U$3 ( \44452 , \44451 , \41092 );
nor \g134399/U$1 ( \44453 , \44450 , \44452 );
xor \g133981/U$1 ( \44454 , \44446 , \44453 );
and \g134969/U$2 ( \44455 , \40175 , \43179 );
and \g134969/U$3 ( \44456 , \43183 , \40207 );
nor \g134969/U$1 ( \44457 , \44455 , \44456 );
and \g134265/U$2 ( \44458 , \44457 , \40137 );
not \g134265/U$4 ( \44459 , \44457 );
and \g134265/U$3 ( \44460 , \44459 , \40136 );
nor \g134265/U$1 ( \44461 , \44458 , \44460 );
xor \g133981/U$1_r1 ( \44462 , \44454 , \44461 );
and \g134859/U$2 ( \44463 , \40672 , \41774 );
and \g134859/U$3 ( \44464 , \41629 , \40858 );
nor \g134859/U$1 ( \44465 , \44463 , \44464 );
and \g134612/U$2 ( \44466 , \44465 , \40678 );
not \g134612/U$4 ( \44467 , \44465 );
and \g134612/U$3 ( \44468 , \44467 , \40677 );
nor \g134612/U$1 ( \44469 , \44466 , \44468 );
and \g135315/U$2 ( \44470 , \43604 , \40138 );
and \g135315/U$3 ( \44471 , \40158 , \43603 );
nor \g135315/U$1 ( \44472 , \44470 , \44471 );
and \g135177/U$2 ( \44473 , \44472 , \42676 );
not \g135177/U$4 ( \44474 , \44472 );
and \g135177/U$3 ( \44475 , \44474 , \42675 );
nor \g135177/U$1 ( \44476 , \44473 , \44475 );
xor \g456264/U$9 ( \44477 , \44469 , \44476 );
and \g135127/U$2 ( \44478 , \40513 , \42344 );
and \g135127/U$3 ( \44479 , \41920 , \40713 );
nor \g135127/U$1 ( \44480 , \44478 , \44479 );
and \g134494/U$2 ( \44481 , \44480 , \40521 );
not \g134494/U$4 ( \44482 , \44480 );
and \g134494/U$3 ( \44483 , \44482 , \40518 );
nor \g134494/U$1 ( \44484 , \44481 , \44483 );
xor \g456264/U$9_r1 ( \44485 , \44477 , \44484 );
and \g456264/U$8 ( \44486 , \44462 , \44485 );
and \g135054/U$2 ( \44487 , \42317 , \40525 );
and \g135054/U$3 ( \44488 , \40472 , \42316 );
nor \g135054/U$1 ( \44489 , \44487 , \44488 );
and \g134419/U$2 ( \44490 , \44489 , \42226 );
not \g134419/U$4 ( \44491 , \44489 );
and \g134419/U$3 ( \44492 , \44491 , \42225 );
nor \g134419/U$1 ( \44493 , \44490 , \44492 );
xor \g134048/U$1 ( \44494 , \44493 , \44217 );
and \g135095/U$2 ( \44495 , \43099 , \40278 );
and \g135095/U$3 ( \44496 , \40189 , \43101 );
nor \g135095/U$1 ( \44497 , \44495 , \44496 );
and \g134533/U$2 ( \44498 , \44497 , \42682 );
not \g134533/U$4 ( \44499 , \44497 );
and \g134533/U$3 ( \44500 , \44499 , \42681 );
nor \g134533/U$1 ( \44501 , \44498 , \44500 );
xor \g134048/U$1_r1 ( \44502 , \44494 , \44501 );
xor \g456264/U$11 ( \44503 , \44469 , \44476 );
xor \g456264/U$11_r1 ( \44504 , \44503 , \44484 );
and \g456264/U$10 ( \44505 , \44502 , \44504 );
and \g456264/U$12 ( \44506 , \44462 , \44502 );
or \g456264/U$7 ( \44507 , \44486 , \44505 , \44506 );
and \g456192/U$4 ( \44508 , \44439 , \44507 );
and \g456192/U$6 ( \44509 , \44436 , \44438 );
or \g456192/U$3 ( \44510 , \44508 , \44509 );
xor \g456247/U$2 ( \44511 , \43995 , \44002 );
xor \g456247/U$1 ( \44512 , \44511 , \44010 );
xor \g456247/U$1_r1 ( \44513 , \44266 , \44271 );
xor \g456247/U$1_r2 ( \44514 , \44512 , \44513 );
xor \g133416/U$4 ( \44515 , \44510 , \44514 );
and \g134747/U$2 ( \44516 , \40175 , \43757 );
and \g134747/U$3 ( \44517 , \43179 , \40207 );
nor \g134747/U$1 ( \44518 , \44516 , \44517 );
and \g134233/U$2 ( \44519 , \44518 , \40137 );
not \g134233/U$4 ( \44520 , \44518 );
and \g134233/U$3 ( \44521 , \44520 , \40136 );
nor \g134233/U$1 ( \44522 , \44519 , \44521 );
and \g134763/U$2 ( \44523 , \42644 , \40472 );
and \g134763/U$3 ( \44524 , \40353 , \42643 );
nor \g134763/U$1 ( \44525 , \44523 , \44524 );
and \g134352/U$2 ( \44526 , \44525 , \42487 );
not \g134352/U$4 ( \44527 , \44525 );
and \g134352/U$3 ( \44528 , \44527 , \42486 );
nor \g134352/U$1 ( \44529 , \44526 , \44528 );
xor \g456250/U$5 ( \44530 , \44522 , \44529 );
and \g134819/U$2 ( \44531 , \40301 , \43183 );
and \g134819/U$3 ( \44532 , \42701 , \40391 );
nor \g134819/U$1 ( \44533 , \44531 , \44532 );
and \g134414/U$2 ( \44534 , \44533 , \40220 );
not \g134414/U$4 ( \44535 , \44533 );
and \g134414/U$3 ( \44536 , \44535 , \40219 );
nor \g134414/U$1 ( \44537 , \44534 , \44536 );
and \g456250/U$4 ( \44538 , \44530 , \44537 );
and \g456250/U$6 ( \44539 , \44522 , \44529 );
or \g456250/U$3 ( \44540 , \44538 , \44539 );
and \g135108/U$2 ( \44541 , \40432 , \42651 );
and \g135108/U$3 ( \44542 , \42609 , \40530 );
nor \g135108/U$1 ( \44543 , \44541 , \44542 );
and \g134258/U$2 ( \44544 , \44543 , \40388 );
not \g134258/U$4 ( \44545 , \44543 );
and \g134258/U$3 ( \44546 , \44545 , \40387 );
nor \g134258/U$1 ( \44547 , \44544 , \44546 );
and \g135297/U$2 ( \44548 , \43604 , \40189 );
and \g135297/U$3 ( \44549 , \40138 , \43603 );
nor \g135297/U$1 ( \44550 , \44548 , \44549 );
and \g135200/U$2 ( \44551 , \44550 , \42676 );
not \g135200/U$4 ( \44552 , \44550 );
and \g135200/U$3 ( \44553 , \44552 , \42675 );
nor \g135200/U$1 ( \44554 , \44551 , \44553 );
xor \g133928/U$4 ( \44555 , \44547 , \44554 );
and \g134844/U$2 ( \44556 , \41623 , \40956 );
and \g134844/U$3 ( \44557 , \40926 , \41745 );
nor \g134844/U$1 ( \44558 , \44556 , \44557 );
and \g134259/U$2 ( \44559 , \44558 , \41325 );
not \g134259/U$4 ( \44560 , \44558 );
and \g134259/U$3 ( \44561 , \44560 , \41324 );
nor \g134259/U$1 ( \44562 , \44559 , \44561 );
and \g133928/U$3 ( \44563 , \44555 , \44562 );
and \g133928/U$5 ( \44564 , \44547 , \44554 );
or \g133928/U$2 ( \44565 , \44563 , \44564 );
xor \g133711/U$4 ( \44566 , \44540 , \44565 );
and \g134741/U$2 ( \44567 , \41948 , \40731 );
and \g134741/U$3 ( \44568 , \40568 , \41947 );
nor \g134741/U$1 ( \44569 , \44567 , \44568 );
and \g134435/U$2 ( \44570 , \44569 , \41755 );
not \g134435/U$4 ( \44571 , \44569 );
and \g134435/U$3 ( \44572 , \44571 , \41952 );
nor \g134435/U$1 ( \44573 , \44570 , \44572 );
and \g134701/U$2 ( \44574 , \41206 , \41107 );
and \g134701/U$3 ( \44575 , \41109 , \41208 );
nor \g134701/U$1 ( \44576 , \44574 , \44575 );
and \g134501/U$2 ( \44577 , \44576 , \41215 );
not \g134501/U$4 ( \44578 , \44576 );
and \g134501/U$3 ( \44579 , \44578 , \41214 );
nor \g134501/U$1 ( \44580 , \44577 , \44579 );
xor \g133976/U$1 ( \44581 , \44573 , \44580 );
and \g134695/U$2 ( \44582 , \40979 , \41345 );
and \g134695/U$3 ( \44583 , \41116 , \41071 );
nor \g134695/U$1 ( \44584 , \44582 , \44583 );
and \g134306/U$2 ( \44585 , \44584 , \40871 );
not \g134306/U$4 ( \44586 , \44584 );
and \g134306/U$3 ( \44587 , \44586 , \40870 );
nor \g134306/U$1 ( \44588 , \44585 , \44587 );
xor \g133976/U$1_r1 ( \44589 , \44581 , \44588 );
and \g133711/U$3 ( \44590 , \44566 , \44589 );
and \g133711/U$5 ( \44591 , \44540 , \44565 );
or \g133711/U$2 ( \44592 , \44590 , \44591 );
xor \g456264/U$5 ( \44593 , \44469 , \44476 );
and \g456264/U$4 ( \44594 , \44593 , \44484 );
and \g456264/U$6 ( \44595 , \44469 , \44476 );
or \g456264/U$3 ( \44596 , \44594 , \44595 );
xor \g134048/U$4 ( \44597 , \44493 , \44217 );
and \g134048/U$3 ( \44598 , \44597 , \44501 );
and \g134048/U$5 ( \44599 , \44493 , \44217 );
or \g134048/U$2 ( \44600 , \44598 , \44599 );
xor \g456222/U$9 ( \44601 , \44596 , \44600 );
xor \g133976/U$4 ( \44602 , \44573 , \44580 );
and \g133976/U$3 ( \44603 , \44602 , \44588 );
and \g133976/U$5 ( \44604 , \44573 , \44580 );
or \g133976/U$2 ( \44605 , \44603 , \44604 );
xor \g456222/U$9_r1 ( \44606 , \44601 , \44605 );
and \g456222/U$8 ( \44607 , \44592 , \44606 );
and \g135107/U$2 ( \44608 , \41623 , \40926 );
and \g135107/U$3 ( \44609 , \40800 , \41745 );
nor \g135107/U$1 ( \44610 , \44608 , \44609 );
and \g134440/U$2 ( \44611 , \44610 , \41325 );
not \g134440/U$4 ( \44612 , \44610 );
and \g134440/U$3 ( \44613 , \44612 , \41324 );
nor \g134440/U$1 ( \44614 , \44611 , \44613 );
and \g134889/U$2 ( \44615 , \40432 , \42609 );
and \g134889/U$3 ( \44616 , \42416 , \40530 );
nor \g134889/U$1 ( \44617 , \44615 , \44616 );
and \g134389/U$2 ( \44618 , \44617 , \40388 );
not \g134389/U$4 ( \44619 , \44617 );
and \g134389/U$3 ( \44620 , \44619 , \40387 );
nor \g134389/U$1 ( \44621 , \44618 , \44620 );
xor \g133959/U$4 ( \44622 , \44614 , \44621 );
and \g135114/U$2 ( \44623 , \40301 , \42701 );
and \g135114/U$3 ( \44624 , \42651 , \40391 );
nor \g135114/U$1 ( \44625 , \44623 , \44624 );
and \g134247/U$2 ( \44626 , \44625 , \40220 );
not \g134247/U$4 ( \44627 , \44625 );
and \g134247/U$3 ( \44628 , \44627 , \40219 );
nor \g134247/U$1 ( \44629 , \44626 , \44628 );
and \g133959/U$3 ( \44630 , \44622 , \44629 );
and \g133959/U$5 ( \44631 , \44614 , \44621 );
or \g133959/U$2 ( \44632 , \44630 , \44631 );
xor \g133981/U$4 ( \44633 , \44446 , \44453 );
and \g133981/U$3 ( \44634 , \44633 , \44461 );
and \g133981/U$5 ( \44635 , \44446 , \44453 );
or \g133981/U$2 ( \44636 , \44634 , \44635 );
xor \g133789/U$1 ( \44637 , \44632 , \44636 );
xor \g134014/U$1 ( \44638 , \44234 , \44241 );
xor \g134014/U$1_r1 ( \44639 , \44638 , \44249 );
xor \g133789/U$1_r1 ( \44640 , \44637 , \44639 );
xor \g456222/U$11 ( \44641 , \44596 , \44600 );
xor \g456222/U$11_r1 ( \44642 , \44641 , \44605 );
and \g456222/U$10 ( \44643 , \44640 , \44642 );
and \g456222/U$12 ( \44644 , \44592 , \44640 );
or \g456222/U$7 ( \44645 , \44607 , \44643 , \44644 );
and \g133416/U$3 ( \44646 , \44515 , \44645 );
and \g133416/U$5 ( \44647 , \44510 , \44514 );
or \g133416/U$2 ( \44648 , \44646 , \44647 );
xor \g456185/U$11 ( \44649 , \44209 , \44255 );
xor \g456185/U$11_r1 ( \44650 , \44649 , \44258 );
and \g456185/U$10 ( \44651 , \44648 , \44650 );
and \g456185/U$12 ( \44652 , \44369 , \44648 );
or \g456185/U$7 ( \44653 , \44372 , \44651 , \44652 );
xor \g133975/U$1 ( \44654 , \44125 , \44132 );
xor \g133975/U$1_r1 ( \44655 , \44654 , \44140 );
xor \g456248/U$9 ( \44656 , \44150 , \44157 );
xor \g456248/U$9_r1 ( \44657 , \44656 , \44165 );
and \g456248/U$8 ( \44658 , \44655 , \44657 );
xor \g133924/U$1 ( \44659 , \44176 , \44182 );
xor \g133924/U$1_r1 ( \44660 , \44659 , \44190 );
xor \g456248/U$11 ( \44661 , \44150 , \44157 );
xor \g456248/U$11_r1 ( \44662 , \44661 , \44165 );
and \g456248/U$10 ( \44663 , \44660 , \44662 );
and \g456248/U$12 ( \44664 , \44655 , \44660 );
or \g456248/U$7 ( \44665 , \44658 , \44663 , \44664 );
xor \g456222/U$5 ( \44666 , \44596 , \44600 );
and \g456222/U$4 ( \44667 , \44666 , \44605 );
and \g456222/U$6 ( \44668 , \44596 , \44600 );
or \g456222/U$3 ( \44669 , \44667 , \44668 );
xor \g133570/U$4 ( \44670 , \44665 , \44669 );
xor \g133774/U$1 ( \44671 , \44216 , \44226 );
xor \g133774/U$1_r1 ( \44672 , \44671 , \44252 );
and \g133570/U$3 ( \44673 , \44670 , \44672 );
and \g133570/U$5 ( \44674 , \44665 , \44669 );
or \g133570/U$2 ( \44675 , \44673 , \44674 );
xor \g456212/U$2 ( \44676 , \43820 , \43827 );
xor \g456212/U$1 ( \44677 , \44676 , \43835 );
xor \g456212/U$1_r1 ( \44678 , \44115 , \44196 );
xor \g456212/U$1_r2 ( \44679 , \44677 , \44678 );
xor \g456176/U$5 ( \44680 , \44675 , \44679 );
xor \g133789/U$4 ( \44681 , \44632 , \44636 );
and \g133789/U$3 ( \44682 , \44681 , \44639 );
and \g133789/U$5 ( \44683 , \44632 , \44636 );
or \g133789/U$2 ( \44684 , \44682 , \44683 );
xor \g133684/U$1 ( \44685 , \44143 , \44168 );
xor \g133684/U$1_r1 ( \44686 , \44685 , \44193 );
xor \g456183/U$5 ( \44687 , \44684 , \44686 );
xor \g456241/U$2 ( \44688 , \43930 , \43937 );
xor \g456241/U$1 ( \44689 , \44688 , \43945 );
xor \g456241/U$1_r1 ( \44690 , \44295 , \44300 );
xor \g456241/U$1_r2 ( \44691 , \44689 , \44690 );
and \g456183/U$4 ( \44692 , \44687 , \44691 );
and \g456183/U$6 ( \44693 , \44684 , \44686 );
or \g456183/U$3 ( \44694 , \44692 , \44693 );
and \g456176/U$4 ( \44695 , \44680 , \44694 );
and \g456176/U$6 ( \44696 , \44675 , \44679 );
or \g456176/U$3 ( \44697 , \44695 , \44696 );
xor \g133243/U$4 ( \44698 , \44653 , \44697 );
xor \g456177/U$2 ( \44699 , \44110 , \44112 );
xor \g456177/U$1 ( \44700 , \44699 , \44201 );
xor \g456177/U$1_r1 ( \44701 , \44339 , \44346 );
xor \g456177/U$1_r2 ( \44702 , \44700 , \44701 );
and \g133243/U$3 ( \44703 , \44698 , \44702 );
and \g133243/U$5 ( \44704 , \44653 , \44697 );
or \g133243/U$2 ( \44705 , \44703 , \44704 );
not \g131591/U$3 ( \44706 , \44705 );
xor \g133211/U$1 ( \44707 , \44351 , \44355 );
xor \g133211/U$1_r1 ( \44708 , \44707 , \44360 );
not \g131591/U$4 ( \44709 , \44708 );
or \g131591/U$2 ( \44710 , \44706 , \44709 );
xor \g456222/U$2 ( \44711 , \44596 , \44600 );
xor \g456222/U$1 ( \44712 , \44711 , \44605 );
xor \g456222/U$1_r1 ( \44713 , \44592 , \44640 );
xor \g456222/U$1_r2 ( \44714 , \44712 , \44713 );
xor \g456192/U$9 ( \44715 , \44436 , \44438 );
xor \g456192/U$9_r1 ( \44716 , \44715 , \44507 );
and \g456192/U$8 ( \44717 , \44714 , \44716 );
xor \g134090/U$1 ( \44718 , \44399 , \44406 );
and \g134960/U$2 ( \44719 , \41087 , \41109 );
and \g134960/U$3 ( \44720 , \41144 , \41328 );
nor \g134960/U$1 ( \44721 , \44719 , \44720 );
and \g134451/U$2 ( \44722 , \44721 , \41093 );
not \g134451/U$4 ( \44723 , \44721 );
and \g134451/U$3 ( \44724 , \44723 , \41092 );
nor \g134451/U$1 ( \44725 , \44722 , \44724 );
xor \g133770/U$4 ( \44726 , \44718 , \44725 );
and \g134739/U$2 ( \44727 , \42317 , \40731 );
and \g134739/U$3 ( \44728 , \40568 , \42316 );
nor \g134739/U$1 ( \44729 , \44727 , \44728 );
and \g134326/U$2 ( \44730 , \44729 , \42226 );
not \g134326/U$4 ( \44731 , \44729 );
and \g134326/U$3 ( \44732 , \44731 , \42225 );
nor \g134326/U$1 ( \44733 , \44730 , \44732 );
xor \g133994/U$4 ( \44734 , \44733 , \44398 );
and \g134870/U$2 ( \44735 , \43099 , \40353 );
and \g134870/U$3 ( \44736 , \40307 , \43101 );
nor \g134870/U$1 ( \44737 , \44735 , \44736 );
and \g134566/U$2 ( \44738 , \44737 , \42682 );
not \g134566/U$4 ( \44739 , \44737 );
and \g134566/U$3 ( \44740 , \44739 , \42681 );
nor \g134566/U$1 ( \44741 , \44738 , \44740 );
and \g133994/U$3 ( \44742 , \44734 , \44741 );
and \g133994/U$5 ( \44743 , \44733 , \44398 );
or \g133994/U$2 ( \44744 , \44742 , \44743 );
and \g133770/U$3 ( \44745 , \44726 , \44744 );
and \g133770/U$5 ( \44746 , \44718 , \44725 );
or \g133770/U$2 ( \44747 , \44745 , \44746 );
xor \g133959/U$1 ( \44748 , \44614 , \44621 );
xor \g133959/U$1_r1 ( \44749 , \44748 , \44629 );
xor \g133580/U$4 ( \44750 , \44747 , \44749 );
and \g134965/U$2 ( \44751 , \41206 , \41345 );
and \g134965/U$3 ( \44752 , \41116 , \41208 );
nor \g134965/U$1 ( \44753 , \44751 , \44752 );
and \g134288/U$2 ( \44754 , \44753 , \41215 );
not \g134288/U$4 ( \44755 , \44753 );
and \g134288/U$3 ( \44756 , \44755 , \41214 );
nor \g134288/U$1 ( \44757 , \44754 , \44756 );
and \g134687/U$2 ( \44758 , \41948 , \40926 );
and \g134687/U$3 ( \44759 , \40800 , \41947 );
nor \g134687/U$1 ( \44760 , \44758 , \44759 );
and \g134461/U$2 ( \44761 , \44760 , \41755 );
not \g134461/U$4 ( \44762 , \44760 );
and \g134461/U$3 ( \44763 , \44762 , \41952 );
nor \g134461/U$1 ( \44764 , \44761 , \44763 );
xor \g134002/U$4 ( \44765 , \44757 , \44764 );
and \g135062/U$2 ( \44766 , \40979 , \41774 );
and \g135062/U$3 ( \44767 , \41629 , \41071 );
nor \g135062/U$1 ( \44768 , \44766 , \44767 );
and \g134450/U$2 ( \44769 , \44768 , \40871 );
not \g134450/U$4 ( \44770 , \44768 );
and \g134450/U$3 ( \44771 , \44770 , \40870 );
nor \g134450/U$1 ( \44772 , \44769 , \44771 );
and \g134002/U$3 ( \44773 , \44765 , \44772 );
and \g134002/U$5 ( \44774 , \44757 , \44764 );
or \g134002/U$2 ( \44775 , \44773 , \44774 );
and \g134985/U$2 ( \44776 , \40513 , \42609 );
and \g134985/U$3 ( \44777 , \42416 , \40713 );
nor \g134985/U$1 ( \44778 , \44776 , \44777 );
and \g134270/U$2 ( \44779 , \44778 , \40521 );
not \g134270/U$4 ( \44780 , \44778 );
and \g134270/U$3 ( \44781 , \44780 , \40518 );
nor \g134270/U$1 ( \44782 , \44779 , \44781 );
and \g135310/U$2 ( \44783 , \43604 , \40278 );
and \g135310/U$3 ( \44784 , \40189 , \43603 );
nor \g135310/U$1 ( \44785 , \44783 , \44784 );
and \g135191/U$2 ( \44786 , \44785 , \42676 );
not \g135191/U$4 ( \44787 , \44785 );
and \g135191/U$3 ( \44788 , \44787 , \42675 );
nor \g135191/U$1 ( \44789 , \44786 , \44788 );
xor \g456263/U$5 ( \44790 , \44782 , \44789 );
and \g135089/U$2 ( \44791 , \40672 , \42344 );
and \g135089/U$3 ( \44792 , \41920 , \40858 );
nor \g135089/U$1 ( \44793 , \44791 , \44792 );
and \g134409/U$2 ( \44794 , \44793 , \40678 );
not \g134409/U$4 ( \44795 , \44793 );
and \g134409/U$3 ( \44796 , \44795 , \40677 );
nor \g134409/U$1 ( \44797 , \44794 , \44796 );
and \g456263/U$4 ( \44798 , \44790 , \44797 );
and \g456263/U$6 ( \44799 , \44782 , \44789 );
or \g456263/U$3 ( \44800 , \44798 , \44799 );
xor \g456219/U$5 ( \44801 , \44775 , \44800 );
and \g135113/U$2 ( \44802 , \40301 , \43179 );
and \g135113/U$3 ( \44803 , \43183 , \40391 );
nor \g135113/U$1 ( \44804 , \44802 , \44803 );
and \g134284/U$2 ( \44805 , \44804 , \40220 );
not \g134284/U$4 ( \44806 , \44804 );
and \g134284/U$3 ( \44807 , \44806 , \40219 );
nor \g134284/U$1 ( \44808 , \44805 , \44807 );
and \g135009/U$2 ( \44809 , \41623 , \41144 );
and \g135009/U$3 ( \44810 , \40956 , \41745 );
nor \g135009/U$1 ( \44811 , \44809 , \44810 );
and \g134470/U$2 ( \44812 , \44811 , \41325 );
not \g134470/U$4 ( \44813 , \44811 );
and \g134470/U$3 ( \44814 , \44813 , \41324 );
nor \g134470/U$1 ( \44815 , \44812 , \44814 );
xor \g133903/U$4 ( \44816 , \44808 , \44815 );
and \g134899/U$2 ( \44817 , \40432 , \42701 );
and \g134899/U$3 ( \44818 , \42651 , \40530 );
nor \g134899/U$1 ( \44819 , \44817 , \44818 );
and \g134540/U$2 ( \44820 , \44819 , \40388 );
not \g134540/U$4 ( \44821 , \44819 );
and \g134540/U$3 ( \44822 , \44821 , \40387 );
nor \g134540/U$1 ( \44823 , \44820 , \44822 );
and \g133903/U$3 ( \44824 , \44816 , \44823 );
and \g133903/U$5 ( \44825 , \44808 , \44815 );
or \g133903/U$2 ( \44826 , \44824 , \44825 );
and \g456219/U$4 ( \44827 , \44801 , \44826 );
and \g456219/U$6 ( \44828 , \44775 , \44800 );
or \g456219/U$3 ( \44829 , \44827 , \44828 );
and \g133580/U$3 ( \44830 , \44750 , \44829 );
and \g133580/U$5 ( \44831 , \44747 , \44749 );
or \g133580/U$2 ( \44832 , \44830 , \44831 );
xor \g456248/U$2 ( \44833 , \44150 , \44157 );
xor \g456248/U$1 ( \44834 , \44833 , \44165 );
xor \g456248/U$1_r1 ( \44835 , \44655 , \44660 );
xor \g456248/U$1_r2 ( \44836 , \44834 , \44835 );
xor \g133419/U$1 ( \44837 , \44832 , \44836 );
xor \g133689/U$1 ( \44838 , \44397 , \44407 );
xor \g133689/U$1_r1 ( \44839 , \44838 , \44433 );
xor \g133928/U$1 ( \44840 , \44547 , \44554 );
xor \g133928/U$1_r1 ( \44841 , \44840 , \44562 );
xor \g456250/U$9 ( \44842 , \44522 , \44529 );
xor \g456250/U$9_r1 ( \44843 , \44842 , \44537 );
and \g456250/U$8 ( \44844 , \44841 , \44843 );
xor \g133923/U$1 ( \44845 , \44379 , \44386 );
xor \g133923/U$1_r1 ( \44846 , \44845 , \44394 );
xor \g456250/U$11 ( \44847 , \44522 , \44529 );
xor \g456250/U$11_r1 ( \44848 , \44847 , \44537 );
and \g456250/U$10 ( \44849 , \44846 , \44848 );
and \g456250/U$12 ( \44850 , \44841 , \44846 );
or \g456250/U$7 ( \44851 , \44844 , \44849 , \44850 );
xor \g456193/U$5 ( \44852 , \44839 , \44851 );
xor \g133711/U$1 ( \44853 , \44540 , \44565 );
xor \g133711/U$1_r1 ( \44854 , \44853 , \44589 );
and \g456193/U$4 ( \44855 , \44852 , \44854 );
and \g456193/U$6 ( \44856 , \44839 , \44851 );
or \g456193/U$3 ( \44857 , \44855 , \44856 );
xor \g133419/U$1_r1 ( \44858 , \44837 , \44857 );
xor \g456192/U$11 ( \44859 , \44436 , \44438 );
xor \g456192/U$11_r1 ( \44860 , \44859 , \44507 );
and \g456192/U$10 ( \44861 , \44858 , \44860 );
and \g456192/U$12 ( \44862 , \44714 , \44858 );
or \g456192/U$7 ( \44863 , \44717 , \44861 , \44862 );
xor \g133416/U$1 ( \44864 , \44510 , \44514 );
xor \g133416/U$1_r1 ( \44865 , \44864 , \44645 );
xor \g133270/U$4 ( \44866 , \44863 , \44865 );
xor \g456183/U$2 ( \44867 , \44684 , \44686 );
xor \g456183/U$1 ( \44868 , \44867 , \44691 );
xor \g133570/U$1 ( \44869 , \44665 , \44669 );
xor \g133570/U$1_r1 ( \44870 , \44869 , \44672 );
xor \g133419/U$4 ( \44871 , \44832 , \44836 );
and \g133419/U$3 ( \44872 , \44871 , \44857 );
and \g133419/U$5 ( \44873 , \44832 , \44836 );
or \g133419/U$2 ( \44874 , \44872 , \44873 );
xor \g456183/U$1_r1 ( \44875 , \44870 , \44874 );
xor \g456183/U$1_r2 ( \44876 , \44868 , \44875 );
and \g133270/U$3 ( \44877 , \44866 , \44876 );
and \g133270/U$5 ( \44878 , \44863 , \44865 );
or \g133270/U$2 ( \44879 , \44877 , \44878 );
xor \g456176/U$2 ( \44880 , \44675 , \44679 );
xor \g456176/U$1 ( \44881 , \44880 , \44694 );
xor \g456183/U$9 ( \44882 , \44684 , \44686 );
xor \g456183/U$9_r1 ( \44883 , \44882 , \44691 );
and \g456183/U$8 ( \44884 , \44870 , \44883 );
xor \g456183/U$11 ( \44885 , \44684 , \44686 );
xor \g456183/U$11_r1 ( \44886 , \44885 , \44691 );
and \g456183/U$10 ( \44887 , \44874 , \44886 );
and \g456183/U$12 ( \44888 , \44870 , \44874 );
or \g456183/U$7 ( \44889 , \44884 , \44887 , \44888 );
xor \g456185/U$2 ( \44890 , \44209 , \44255 );
xor \g456185/U$1 ( \44891 , \44890 , \44258 );
xor \g456185/U$1_r1 ( \44892 , \44369 , \44648 );
xor \g456185/U$1_r2 ( \44893 , \44891 , \44892 );
xor \g456176/U$1_r1 ( \44894 , \44889 , \44893 );
xor \g456176/U$1_r2 ( \44895 , \44881 , \44894 );
and \g131712/U$2 ( \44896 , \44879 , \44895 );
xor \g133198/U$1 ( \44897 , \44895 , \44879 );
xor \g133580/U$1 ( \44898 , \44747 , \44749 );
xor \g133580/U$1_r1 ( \44899 , \44898 , \44829 );
xor \g456193/U$9 ( \44900 , \44839 , \44851 );
xor \g456193/U$9_r1 ( \44901 , \44900 , \44854 );
and \g456193/U$8 ( \44902 , \44899 , \44901 );
xor \g133903/U$1 ( \44903 , \44808 , \44815 );
xor \g133903/U$1_r1 ( \44904 , \44903 , \44823 );
xor \g134002/U$1 ( \44905 , \44757 , \44764 );
xor \g134002/U$1_r1 ( \44906 , \44905 , \44772 );
xor \g456225/U$5 ( \44907 , \44904 , \44906 );
and \g135106/U$2 ( \44908 , \41087 , \41107 );
and \g135106/U$3 ( \44909 , \41109 , \41328 );
nor \g135106/U$1 ( \44910 , \44908 , \44909 );
and \g134283/U$2 ( \44911 , \44910 , \41093 );
not \g134283/U$4 ( \44912 , \44910 );
and \g134283/U$3 ( \44913 , \44912 , \41092 );
nor \g134283/U$1 ( \44914 , \44911 , \44913 );
and \g134699/U$2 ( \44915 , \42644 , \40525 );
and \g134699/U$3 ( \44916 , \40472 , \42643 );
nor \g134699/U$1 ( \44917 , \44915 , \44916 );
and \g134372/U$2 ( \44918 , \44917 , \42487 );
not \g134372/U$4 ( \44919 , \44917 );
and \g134372/U$3 ( \44920 , \44919 , \42486 );
nor \g134372/U$1 ( \44921 , \44918 , \44920 );
xor \g133848/U$1 ( \44922 , \44914 , \44921 );
nor \g135208/U$1 ( \44923 , \40296 , \43607 );
nor \g135169/U$1 ( \44924 , \44923 , \40220 );
and \g134891/U$2 ( \44925 , \43099 , \40472 );
and \g134891/U$3 ( \44926 , \40353 , \43101 );
nor \g134891/U$1 ( \44927 , \44925 , \44926 );
and \g134538/U$2 ( \44928 , \44927 , \42682 );
not \g134538/U$4 ( \44929 , \44927 );
and \g134538/U$3 ( \44930 , \44929 , \42681 );
nor \g134538/U$1 ( \44931 , \44928 , \44930 );
and \g134089/U$2 ( \44932 , \44924 , \44931 );
xor \g133848/U$1_r1 ( \44933 , \44922 , \44932 );
and \g456225/U$4 ( \44934 , \44907 , \44933 );
and \g456225/U$6 ( \44935 , \44904 , \44906 );
or \g456225/U$3 ( \44936 , \44934 , \44935 );
xor \g456250/U$2 ( \44937 , \44522 , \44529 );
xor \g456250/U$1 ( \44938 , \44937 , \44537 );
xor \g456250/U$1_r1 ( \44939 , \44841 , \44846 );
xor \g456250/U$1_r2 ( \44940 , \44938 , \44939 );
xor \g133510/U$4 ( \44941 , \44936 , \44940 );
xor \g133848/U$4 ( \44942 , \44914 , \44921 );
and \g133848/U$3 ( \44943 , \44942 , \44932 );
and \g133848/U$5 ( \44944 , \44914 , \44921 );
or \g133848/U$2 ( \44945 , \44943 , \44944 );
xor \g133910/U$1 ( \44946 , \44415 , \44422 );
xor \g133910/U$1_r1 ( \44947 , \44946 , \44430 );
xor \g133631/U$1 ( \44948 , \44945 , \44947 );
xor \g133770/U$1 ( \44949 , \44718 , \44725 );
xor \g133770/U$1_r1 ( \44950 , \44949 , \44744 );
xor \g133631/U$1_r1 ( \44951 , \44948 , \44950 );
and \g133510/U$3 ( \44952 , \44941 , \44951 );
and \g133510/U$5 ( \44953 , \44936 , \44940 );
or \g133510/U$2 ( \44954 , \44952 , \44953 );
xor \g456193/U$11 ( \44955 , \44839 , \44851 );
xor \g456193/U$11_r1 ( \44956 , \44955 , \44854 );
and \g456193/U$10 ( \44957 , \44954 , \44956 );
and \g456193/U$12 ( \44958 , \44899 , \44954 );
or \g456193/U$7 ( \44959 , \44902 , \44957 , \44958 );
xor \g133631/U$4 ( \44960 , \44945 , \44947 );
and \g133631/U$3 ( \44961 , \44960 , \44950 );
and \g133631/U$5 ( \44962 , \44945 , \44947 );
or \g133631/U$2 ( \44963 , \44961 , \44962 );
xor \g456264/U$2 ( \44964 , \44469 , \44476 );
xor \g456264/U$1 ( \44965 , \44964 , \44484 );
xor \g456264/U$1_r1 ( \44966 , \44462 , \44502 );
xor \g456264/U$1_r2 ( \44967 , \44965 , \44966 );
xor \g456178/U$5 ( \44968 , \44963 , \44967 );
and \g134824/U$2 ( \44969 , \40979 , \41920 );
and \g134824/U$3 ( \44970 , \41774 , \41071 );
nor \g134824/U$1 ( \44971 , \44969 , \44970 );
and \g134390/U$2 ( \44972 , \44971 , \40871 );
not \g134390/U$4 ( \44973 , \44971 );
and \g134390/U$3 ( \44974 , \44973 , \40870 );
nor \g134390/U$1 ( \44975 , \44972 , \44974 );
and \g134945/U$2 ( \44976 , \42317 , \40800 );
and \g134945/U$3 ( \44977 , \40731 , \42316 );
nor \g134945/U$1 ( \44978 , \44976 , \44977 );
and \g134228/U$2 ( \44979 , \44978 , \42226 );
not \g134228/U$4 ( \44980 , \44978 );
and \g134228/U$3 ( \44981 , \44980 , \42225 );
nor \g134228/U$1 ( \44982 , \44979 , \44981 );
xor \g133914/U$4 ( \44983 , \44975 , \44982 );
and \g134992/U$2 ( \44984 , \41206 , \41629 );
and \g134992/U$3 ( \44985 , \41345 , \41208 );
nor \g134992/U$1 ( \44986 , \44984 , \44985 );
or \g134169/U$2 ( \44987 , \44986 , \41214 );
nand \g134641/U$1 ( \44988 , \41214 , \44986 );
nand \g134169/U$1 ( \44989 , \44987 , \44988 );
and \g133914/U$3 ( \44990 , \44983 , \44989 );
and \g133914/U$5 ( \44991 , \44975 , \44982 );
or \g133914/U$2 ( \44992 , \44990 , \44991 );
and \g135036/U$2 ( \44993 , \40432 , \43183 );
and \g135036/U$3 ( \44994 , \42701 , \40530 );
nor \g135036/U$1 ( \44995 , \44993 , \44994 );
and \g134361/U$2 ( \44996 , \44995 , \40388 );
not \g134361/U$4 ( \44997 , \44995 );
and \g134361/U$3 ( \44998 , \44997 , \40387 );
nor \g134361/U$1 ( \44999 , \44996 , \44998 );
and \g135316/U$2 ( \45000 , \43604 , \40307 );
and \g135316/U$3 ( \45001 , \40278 , \43603 );
nor \g135316/U$1 ( \45002 , \45000 , \45001 );
and \g135184/U$2 ( \45003 , \45002 , \42676 );
not \g135184/U$4 ( \45004 , \45002 );
and \g135184/U$3 ( \45005 , \45004 , \42675 );
nor \g135184/U$1 ( \45006 , \45003 , \45005 );
xor \g456244/U$5 ( \45007 , \44999 , \45006 );
and \g134833/U$2 ( \45008 , \41623 , \41109 );
and \g134833/U$3 ( \45009 , \41144 , \41745 );
nor \g134833/U$1 ( \45010 , \45008 , \45009 );
and \g134252/U$2 ( \45011 , \45010 , \41325 );
not \g134252/U$4 ( \45012 , \45010 );
and \g134252/U$3 ( \45013 , \45012 , \41324 );
nor \g134252/U$1 ( \45014 , \45011 , \45013 );
and \g456244/U$4 ( \45015 , \45007 , \45014 );
and \g456244/U$6 ( \45016 , \44999 , \45006 );
or \g456244/U$3 ( \45017 , \45015 , \45016 );
xor \g133700/U$4 ( \45018 , \44992 , \45017 );
and \g135055/U$2 ( \45019 , \41948 , \40956 );
and \g135055/U$3 ( \45020 , \40926 , \41947 );
nor \g135055/U$1 ( \45021 , \45019 , \45020 );
and \g134266/U$2 ( \45022 , \45021 , \41755 );
not \g134266/U$4 ( \45023 , \45021 );
and \g134266/U$3 ( \45024 , \45023 , \41952 );
nor \g134266/U$1 ( \45025 , \45022 , \45024 );
and \g134718/U$2 ( \45026 , \40672 , \42416 );
and \g134718/U$3 ( \45027 , \42344 , \40858 );
nor \g134718/U$1 ( \45028 , \45026 , \45027 );
and \g134251/U$2 ( \45029 , \45028 , \40678 );
not \g134251/U$4 ( \45030 , \45028 );
and \g134251/U$3 ( \45031 , \45030 , \40677 );
nor \g134251/U$1 ( \45032 , \45029 , \45031 );
xor \g133966/U$4 ( \45033 , \45025 , \45032 );
and \g135026/U$2 ( \45034 , \40513 , \42651 );
and \g135026/U$3 ( \45035 , \42609 , \40713 );
nor \g135026/U$1 ( \45036 , \45034 , \45035 );
and \g134437/U$2 ( \45037 , \45036 , \40521 );
not \g134437/U$4 ( \45038 , \45036 );
and \g134437/U$3 ( \45039 , \45038 , \40518 );
nor \g134437/U$1 ( \45040 , \45037 , \45039 );
and \g133966/U$3 ( \45041 , \45033 , \45040 );
and \g133966/U$5 ( \45042 , \45025 , \45032 );
or \g133966/U$2 ( \45043 , \45041 , \45042 );
and \g133700/U$3 ( \45044 , \45018 , \45043 );
and \g133700/U$5 ( \45045 , \44992 , \45017 );
or \g133700/U$2 ( \45046 , \45044 , \45045 );
xor \g456219/U$9 ( \45047 , \44775 , \44800 );
xor \g456219/U$9_r1 ( \45048 , \45047 , \44826 );
and \g456219/U$8 ( \45049 , \45046 , \45048 );
and \g134750/U$2 ( \45050 , \41087 , \41116 );
and \g134750/U$3 ( \45051 , \41107 , \41328 );
nor \g134750/U$1 ( \45052 , \45050 , \45051 );
and \g134608/U$2 ( \45053 , \45052 , \41093 );
not \g134608/U$4 ( \45054 , \45052 );
and \g134608/U$3 ( \45055 , \45054 , \41092 );
nor \g134608/U$1 ( \45056 , \45053 , \45055 );
and \g134793/U$2 ( \45057 , \42644 , \40568 );
and \g134793/U$3 ( \45058 , \40525 , \42643 );
nor \g134793/U$1 ( \45059 , \45057 , \45058 );
and \g134432/U$2 ( \45060 , \45059 , \42487 );
not \g134432/U$4 ( \45061 , \45059 );
and \g134432/U$3 ( \45062 , \45061 , \42486 );
nor \g134432/U$1 ( \45063 , \45060 , \45062 );
xor \g134019/U$4 ( \45064 , \45056 , \45063 );
and \g135115/U$2 ( \45065 , \40301 , \43757 );
and \g135115/U$3 ( \45066 , \43179 , \40391 );
nor \g135115/U$1 ( \45067 , \45065 , \45066 );
and \g134324/U$2 ( \45068 , \45067 , \40220 );
not \g134324/U$4 ( \45069 , \45067 );
and \g134324/U$3 ( \45070 , \45069 , \40219 );
nor \g134324/U$1 ( \45071 , \45068 , \45070 );
and \g134019/U$3 ( \45072 , \45064 , \45071 );
and \g134019/U$5 ( \45073 , \45056 , \45063 );
or \g134019/U$2 ( \45074 , \45072 , \45073 );
xor \g456263/U$9 ( \45075 , \44782 , \44789 );
xor \g456263/U$9_r1 ( \45076 , \45075 , \44797 );
and \g456263/U$8 ( \45077 , \45074 , \45076 );
xor \g133994/U$1 ( \45078 , \44733 , \44398 );
xor \g133994/U$1_r1 ( \45079 , \45078 , \44741 );
xor \g456263/U$11 ( \45080 , \44782 , \44789 );
xor \g456263/U$11_r1 ( \45081 , \45080 , \44797 );
and \g456263/U$10 ( \45082 , \45079 , \45081 );
and \g456263/U$12 ( \45083 , \45074 , \45079 );
or \g456263/U$7 ( \45084 , \45077 , \45082 , \45083 );
xor \g456219/U$11 ( \45085 , \44775 , \44800 );
xor \g456219/U$11_r1 ( \45086 , \45085 , \44826 );
and \g456219/U$10 ( \45087 , \45084 , \45086 );
and \g456219/U$12 ( \45088 , \45046 , \45084 );
or \g456219/U$7 ( \45089 , \45049 , \45087 , \45088 );
and \g456178/U$4 ( \45090 , \44968 , \45089 );
and \g456178/U$6 ( \45091 , \44963 , \44967 );
or \g456178/U$3 ( \45092 , \45090 , \45091 );
xor \g133293/U$4 ( \45093 , \44959 , \45092 );
xor \g456192/U$2 ( \45094 , \44436 , \44438 );
xor \g456192/U$1 ( \45095 , \45094 , \44507 );
xor \g456192/U$1_r1 ( \45096 , \44714 , \44858 );
xor \g456192/U$1_r2 ( \45097 , \45095 , \45096 );
and \g133293/U$3 ( \45098 , \45093 , \45097 );
and \g133293/U$5 ( \45099 , \44959 , \45092 );
or \g133293/U$2 ( \45100 , \45098 , \45099 );
not \g131774/U$3 ( \45101 , \45100 );
xor \g133270/U$1 ( \45102 , \44863 , \44865 );
xor \g133270/U$1_r1 ( \45103 , \45102 , \44876 );
not \g131774/U$4 ( \45104 , \45103 );
or \g131774/U$2 ( \45105 , \45101 , \45104 );
xor \g133293/U$1 ( \45106 , \44959 , \45092 );
xor \g133293/U$1_r1 ( \45107 , \45106 , \45097 );
xor \g133700/U$1 ( \45108 , \44992 , \45017 );
xor \g133700/U$1_r1 ( \45109 , \45108 , \45043 );
xor \g456225/U$9 ( \45110 , \44904 , \44906 );
xor \g456225/U$9_r1 ( \45111 , \45110 , \44933 );
and \g456225/U$8 ( \45112 , \45109 , \45111 );
xor \g456263/U$2 ( \45113 , \44782 , \44789 );
xor \g456263/U$1 ( \45114 , \45113 , \44797 );
xor \g456263/U$1_r1 ( \45115 , \45074 , \45079 );
xor \g456263/U$1_r2 ( \45116 , \45114 , \45115 );
xor \g456225/U$11 ( \45117 , \44904 , \44906 );
xor \g456225/U$11_r1 ( \45118 , \45117 , \44933 );
and \g456225/U$10 ( \45119 , \45116 , \45118 );
and \g456225/U$12 ( \45120 , \45109 , \45116 );
or \g456225/U$7 ( \45121 , \45112 , \45119 , \45120 );
xor \g133914/U$1 ( \45122 , \44975 , \44982 );
xor \g133914/U$1_r1 ( \45123 , \45122 , \44989 );
xor \g456244/U$9 ( \45124 , \44999 , \45006 );
xor \g456244/U$9_r1 ( \45125 , \45124 , \45014 );
and \g456244/U$8 ( \45126 , \45123 , \45125 );
xor \g133966/U$1 ( \45127 , \45025 , \45032 );
xor \g133966/U$1_r1 ( \45128 , \45127 , \45040 );
xor \g456244/U$11 ( \45129 , \44999 , \45006 );
xor \g456244/U$11_r1 ( \45130 , \45129 , \45014 );
and \g456244/U$10 ( \45131 , \45128 , \45130 );
and \g456244/U$12 ( \45132 , \45123 , \45128 );
or \g456244/U$7 ( \45133 , \45126 , \45131 , \45132 );
and \g134887/U$2 ( \45134 , \40672 , \42609 );
and \g134887/U$3 ( \45135 , \42416 , \40858 );
nor \g134887/U$1 ( \45136 , \45134 , \45135 );
and \g134480/U$2 ( \45137 , \45136 , \40678 );
not \g134480/U$4 ( \45138 , \45136 );
and \g134480/U$3 ( \45139 , \45138 , \40677 );
nor \g134480/U$1 ( \45140 , \45137 , \45139 );
and \g135290/U$2 ( \45141 , \43604 , \40353 );
and \g135290/U$3 ( \45142 , \40307 , \43603 );
nor \g135290/U$1 ( \45143 , \45141 , \45142 );
and \g135203/U$2 ( \45144 , \45143 , \42676 );
not \g135203/U$4 ( \45145 , \45143 );
and \g135203/U$3 ( \45146 , \45145 , \42675 );
nor \g135203/U$1 ( \45147 , \45144 , \45146 );
xor \g134036/U$4 ( \45148 , \45140 , \45147 );
and \g135063/U$2 ( \45149 , \40513 , \42701 );
and \g135063/U$3 ( \45150 , \42651 , \40713 );
nor \g135063/U$1 ( \45151 , \45149 , \45150 );
or \g134150/U$2 ( \45152 , \45151 , \40518 );
nand \g134634/U$1 ( \45153 , \40518 , \45151 );
nand \g134150/U$1 ( \45154 , \45152 , \45153 );
and \g134036/U$3 ( \45155 , \45148 , \45154 );
and \g134036/U$5 ( \45156 , \45140 , \45147 );
or \g134036/U$2 ( \45157 , \45155 , \45156 );
xor \g134089/U$1 ( \45158 , \44924 , \44931 );
xor \g456216/U$5 ( \45159 , \45157 , \45158 );
and \g134916/U$2 ( \45160 , \41948 , \41144 );
and \g134916/U$3 ( \45161 , \40956 , \41947 );
nor \g134916/U$1 ( \45162 , \45160 , \45161 );
and \g134279/U$2 ( \45163 , \45162 , \41755 );
not \g134279/U$4 ( \45164 , \45162 );
and \g134279/U$3 ( \45165 , \45164 , \41952 );
nor \g134279/U$1 ( \45166 , \45163 , \45165 );
and \g134993/U$2 ( \45167 , \41206 , \41774 );
and \g134993/U$3 ( \45168 , \41629 , \41208 );
nor \g134993/U$1 ( \45169 , \45167 , \45168 );
and \g134348/U$2 ( \45170 , \45169 , \41215 );
not \g134348/U$4 ( \45171 , \45169 );
and \g134348/U$3 ( \45172 , \45171 , \41214 );
nor \g134348/U$1 ( \45173 , \45170 , \45172 );
xor \g456266/U$5 ( \45174 , \45166 , \45173 );
and \g134760/U$2 ( \45175 , \40979 , \42344 );
and \g134760/U$3 ( \45176 , \41920 , \41071 );
nor \g134760/U$1 ( \45177 , \45175 , \45176 );
and \g134458/U$2 ( \45178 , \45177 , \40871 );
not \g134458/U$4 ( \45179 , \45177 );
and \g134458/U$3 ( \45180 , \45179 , \40870 );
nor \g134458/U$1 ( \45181 , \45178 , \45180 );
and \g456266/U$4 ( \45182 , \45174 , \45181 );
and \g456266/U$6 ( \45183 , \45166 , \45173 );
or \g456266/U$3 ( \45184 , \45182 , \45183 );
and \g456216/U$4 ( \45185 , \45159 , \45184 );
and \g456216/U$6 ( \45186 , \45157 , \45158 );
or \g456216/U$3 ( \45187 , \45185 , \45186 );
xor \g133513/U$4 ( \45188 , \45133 , \45187 );
and \g135139/U$2 ( \45189 , \42317 , \40926 );
and \g135139/U$3 ( \45190 , \40800 , \42316 );
nor \g135139/U$1 ( \45191 , \45189 , \45190 );
and \g134588/U$2 ( \45192 , \45191 , \42226 );
not \g134588/U$4 ( \45193 , \45191 );
and \g134588/U$3 ( \45194 , \45193 , \42225 );
nor \g134588/U$1 ( \45195 , \45192 , \45194 );
xor \g134009/U$4 ( \45196 , \45195 , \44923 );
and \g135111/U$2 ( \45197 , \43099 , \40525 );
and \g135111/U$3 ( \45198 , \40472 , \43101 );
nor \g135111/U$1 ( \45199 , \45197 , \45198 );
and \g134418/U$2 ( \45200 , \45199 , \42682 );
not \g134418/U$4 ( \45201 , \45199 );
and \g134418/U$3 ( \45202 , \45201 , \42681 );
nor \g134418/U$1 ( \45203 , \45200 , \45202 );
and \g134009/U$3 ( \45204 , \45196 , \45203 );
and \g134009/U$5 ( \45205 , \45195 , \44923 );
or \g134009/U$2 ( \45206 , \45204 , \45205 );
and \g134709/U$2 ( \45207 , \42644 , \40731 );
and \g134709/U$3 ( \45208 , \40568 , \42643 );
nor \g134709/U$1 ( \45209 , \45207 , \45208 );
and \g134469/U$2 ( \45210 , \45209 , \42486 );
not \g134469/U$4 ( \45211 , \45209 );
and \g134469/U$3 ( \45212 , \45211 , \42487 );
nor \g134469/U$1 ( \45213 , \45210 , \45212 );
and \g134964/U$2 ( \45214 , \41623 , \41107 );
and \g134964/U$3 ( \45215 , \41109 , \41745 );
nor \g134964/U$1 ( \45216 , \45214 , \45215 );
and \g134430/U$2 ( \45217 , \45216 , \41324 );
not \g134430/U$4 ( \45218 , \45216 );
and \g134430/U$3 ( \45219 , \45218 , \41325 );
nor \g134430/U$1 ( \45220 , \45217 , \45219 );
xor \g456274/U$4 ( \45221 , \45213 , \45220 );
and \g134928/U$2 ( \45222 , \40432 , \43179 );
and \g134928/U$3 ( \45223 , \43183 , \40530 );
nor \g134928/U$1 ( \45224 , \45222 , \45223 );
and \g134195/U$2 ( \45225 , \45224 , \40387 );
not \g134195/U$4 ( \45226 , \45224 );
and \g134195/U$3 ( \45227 , \45226 , \40388 );
nor \g134195/U$1 ( \45228 , \45225 , \45227 );
and \g456274/U$3 ( \45229 , \45221 , \45228 );
and \g456274/U$5 ( \45230 , \45213 , \45220 );
nor \g456274/U$2 ( \45231 , \45229 , \45230 );
xor \g133675/U$4 ( \45232 , \45206 , \45231 );
xor \g134019/U$1 ( \45233 , \45056 , \45063 );
xor \g134019/U$1_r1 ( \45234 , \45233 , \45071 );
and \g133675/U$3 ( \45235 , \45232 , \45234 );
and \g133675/U$5 ( \45236 , \45206 , \45231 );
or \g133675/U$2 ( \45237 , \45235 , \45236 );
and \g133513/U$3 ( \45238 , \45188 , \45237 );
and \g133513/U$5 ( \45239 , \45133 , \45187 );
or \g133513/U$2 ( \45240 , \45238 , \45239 );
xor \g133406/U$4 ( \45241 , \45121 , \45240 );
xor \g456219/U$2 ( \45242 , \44775 , \44800 );
xor \g456219/U$1 ( \45243 , \45242 , \44826 );
xor \g456219/U$1_r1 ( \45244 , \45046 , \45084 );
xor \g456219/U$1_r2 ( \45245 , \45243 , \45244 );
and \g133406/U$3 ( \45246 , \45241 , \45245 );
and \g133406/U$5 ( \45247 , \45121 , \45240 );
or \g133406/U$2 ( \45248 , \45246 , \45247 );
xor \g456178/U$9 ( \45249 , \44963 , \44967 );
xor \g456178/U$9_r1 ( \45250 , \45249 , \45089 );
and \g456178/U$8 ( \45251 , \45248 , \45250 );
xor \g456193/U$2 ( \45252 , \44839 , \44851 );
xor \g456193/U$1 ( \45253 , \45252 , \44854 );
xor \g456193/U$1_r1 ( \45254 , \44899 , \44954 );
xor \g456193/U$1_r2 ( \45255 , \45253 , \45254 );
xor \g456178/U$11 ( \45256 , \44963 , \44967 );
xor \g456178/U$11_r1 ( \45257 , \45256 , \45089 );
and \g456178/U$10 ( \45258 , \45255 , \45257 );
and \g456178/U$12 ( \45259 , \45248 , \45255 );
or \g456178/U$7 ( \45260 , \45251 , \45258 , \45259 );
and \g131836/U$2 ( \45261 , \45107 , \45260 );
xor \g133260/U$1 ( \45262 , \45260 , \45107 );
xor \g134036/U$1 ( \45263 , \45140 , \45147 );
xor \g134036/U$1_r1 ( \45264 , \45263 , \45154 );
xor \g456266/U$9 ( \45265 , \45166 , \45173 );
xor \g456266/U$9_r1 ( \45266 , \45265 , \45181 );
and \g456266/U$8 ( \45267 , \45264 , \45266 );
xor \g134009/U$1 ( \45268 , \45195 , \44923 );
xor \g134009/U$1_r1 ( \45269 , \45268 , \45203 );
xor \g456266/U$11 ( \45270 , \45166 , \45173 );
xor \g456266/U$11_r1 ( \45271 , \45270 , \45181 );
and \g456266/U$10 ( \45272 , \45269 , \45271 );
and \g456266/U$12 ( \45273 , \45264 , \45269 );
or \g456266/U$7 ( \45274 , \45267 , \45272 , \45273 );
nor \g135216/U$1 ( \45275 , \40426 , \43607 );
nor \g135170/U$1 ( \45276 , \45275 , \40388 );
and \g134962/U$2 ( \45277 , \43099 , \40568 );
and \g134962/U$3 ( \45278 , \40525 , \43101 );
nor \g134962/U$1 ( \45279 , \45277 , \45278 );
and \g134445/U$2 ( \45280 , \45279 , \42682 );
not \g134445/U$4 ( \45281 , \45279 );
and \g134445/U$3 ( \45282 , \45281 , \42681 );
nor \g134445/U$1 ( \45283 , \45280 , \45282 );
and \g134092/U$2 ( \45284 , \45276 , \45283 );
and \g134755/U$2 ( \45285 , \41087 , \41345 );
and \g134755/U$3 ( \45286 , \41116 , \41328 );
nor \g134755/U$1 ( \45287 , \45285 , \45286 );
and \g134502/U$2 ( \45288 , \45287 , \41093 );
not \g134502/U$4 ( \45289 , \45287 );
and \g134502/U$3 ( \45290 , \45289 , \41092 );
nor \g134502/U$1 ( \45291 , \45288 , \45290 );
xor \g133785/U$4 ( \45292 , \45284 , \45291 );
and \g135052/U$2 ( \45293 , \40672 , \42651 );
and \g135052/U$3 ( \45294 , \42609 , \40858 );
nor \g135052/U$1 ( \45295 , \45293 , \45294 );
and \g134309/U$2 ( \45296 , \45295 , \40677 );
not \g134309/U$4 ( \45297 , \45295 );
and \g134309/U$3 ( \45298 , \45297 , \40678 );
nor \g134309/U$1 ( \45299 , \45296 , \45298 );
and \g134976/U$2 ( \45300 , \40513 , \43183 );
and \g134976/U$3 ( \45301 , \42701 , \40713 );
nor \g134976/U$1 ( \45302 , \45300 , \45301 );
and \g134204/U$2 ( \45303 , \45302 , \40518 );
not \g134204/U$4 ( \45304 , \45302 );
and \g134204/U$3 ( \45305 , \45304 , \40521 );
nor \g134204/U$1 ( \45306 , \45303 , \45305 );
or \g134096/U$2 ( \45307 , \45299 , \45306 );
not \g134108/U$3 ( \45308 , \45306 );
not \g134108/U$4 ( \45309 , \45299 );
or \g134108/U$2 ( \45310 , \45308 , \45309 );
and \g134770/U$2 ( \45311 , \41948 , \41109 );
and \g134770/U$3 ( \45312 , \41144 , \41947 );
nor \g134770/U$1 ( \45313 , \45311 , \45312 );
and \g134378/U$2 ( \45314 , \45313 , \41755 );
not \g134378/U$4 ( \45315 , \45313 );
and \g134378/U$3 ( \45316 , \45315 , \41952 );
nor \g134378/U$1 ( \45317 , \45314 , \45316 );
nand \g134108/U$1 ( \45318 , \45310 , \45317 );
nand \g134096/U$1 ( \45319 , \45307 , \45318 );
and \g133785/U$3 ( \45320 , \45292 , \45319 );
and \g133785/U$5 ( \45321 , \45284 , \45291 );
or \g133785/U$2 ( \45322 , \45320 , \45321 );
xor \g133582/U$4 ( \45323 , \45274 , \45322 );
xor \g133675/U$1 ( \45324 , \45206 , \45231 );
xor \g133675/U$1_r1 ( \45325 , \45324 , \45234 );
and \g133582/U$3 ( \45326 , \45323 , \45325 );
and \g133582/U$5 ( \45327 , \45274 , \45322 );
or \g133582/U$2 ( \45328 , \45326 , \45327 );
and \g134726/U$2 ( \45329 , \42644 , \40800 );
and \g134726/U$3 ( \45330 , \40731 , \42643 );
nor \g134726/U$1 ( \45331 , \45329 , \45330 );
and \g134413/U$2 ( \45332 , \45331 , \42486 );
not \g134413/U$4 ( \45333 , \45331 );
and \g134413/U$3 ( \45334 , \45333 , \42487 );
nor \g134413/U$1 ( \45335 , \45332 , \45334 );
and \g135313/U$2 ( \45336 , \43604 , \40472 );
and \g135313/U$3 ( \45337 , \40353 , \43603 );
nor \g135313/U$1 ( \45338 , \45336 , \45337 );
and \g135202/U$2 ( \45339 , \45338 , \42675 );
not \g135202/U$4 ( \45340 , \45338 );
and \g135202/U$3 ( \45341 , \45340 , \42676 );
nor \g135202/U$1 ( \45342 , \45339 , \45341 );
xor \g133947/U$4 ( \45343 , \45335 , \45342 );
and \g134775/U$2 ( \45344 , \40432 , \43757 );
and \g134775/U$3 ( \45345 , \43179 , \40530 );
nor \g134775/U$1 ( \45346 , \45344 , \45345 );
and \g134595/U$2 ( \45347 , \45346 , \40387 );
not \g134595/U$4 ( \45348 , \45346 );
and \g134595/U$3 ( \45349 , \45348 , \40388 );
nor \g134595/U$1 ( \45350 , \45347 , \45349 );
and \g133947/U$3 ( \45351 , \45343 , \45350 );
and \g133947/U$5 ( \45352 , \45335 , \45342 );
or \g133947/U$2 ( \45353 , \45351 , \45352 );
and \g134727/U$2 ( \45354 , \42317 , \40956 );
and \g134727/U$3 ( \45355 , \40926 , \42316 );
nor \g134727/U$1 ( \45356 , \45354 , \45355 );
and \g134527/U$2 ( \45357 , \45356 , \42225 );
not \g134527/U$4 ( \45358 , \45356 );
and \g134527/U$3 ( \45359 , \45358 , \42226 );
nor \g134527/U$1 ( \45360 , \45357 , \45359 );
not \g134100/U$3 ( \45361 , \45360 );
and \g135059/U$2 ( \45362 , \40979 , \42416 );
and \g135059/U$3 ( \45363 , \42344 , \41071 );
nor \g135059/U$1 ( \45364 , \45362 , \45363 );
and \g134439/U$2 ( \45365 , \45364 , \40870 );
not \g134439/U$4 ( \45366 , \45364 );
and \g134439/U$3 ( \45367 , \45366 , \40871 );
nor \g134439/U$1 ( \45368 , \45365 , \45367 );
not \g134100/U$4 ( \45369 , \45368 );
and \g134100/U$2 ( \45370 , \45361 , \45369 );
and \g134111/U$2 ( \45371 , \45368 , \45360 );
and \g135072/U$2 ( \45372 , \41206 , \41920 );
and \g135072/U$3 ( \45373 , \41774 , \41208 );
nor \g135072/U$1 ( \45374 , \45372 , \45373 );
and \g134281/U$2 ( \45375 , \45374 , \41214 );
not \g134281/U$4 ( \45376 , \45374 );
and \g134281/U$3 ( \45377 , \45376 , \41215 );
nor \g134281/U$1 ( \45378 , \45375 , \45377 );
nor \g134111/U$1 ( \45379 , \45371 , \45378 );
nor \g134100/U$1 ( \45380 , \45370 , \45379 );
xor \g456271/U$4 ( \45381 , \45353 , \45380 );
xor \g456274/U$1 ( \45382 , \45213 , \45220 );
xor \g456274/U$1_r1 ( \45383 , \45382 , \45228 );
and \g456271/U$3 ( \45384 , \45381 , \45383 );
and \g456271/U$5 ( \45385 , \45353 , \45380 );
nor \g456271/U$2 ( \45386 , \45384 , \45385 );
xor \g456216/U$9 ( \45387 , \45157 , \45158 );
xor \g456216/U$9_r1 ( \45388 , \45387 , \45184 );
and \g456216/U$8 ( \45389 , \45386 , \45388 );
xor \g456244/U$2 ( \45390 , \44999 , \45006 );
xor \g456244/U$1 ( \45391 , \45390 , \45014 );
xor \g456244/U$1_r1 ( \45392 , \45123 , \45128 );
xor \g456244/U$1_r2 ( \45393 , \45391 , \45392 );
xor \g456216/U$11 ( \45394 , \45157 , \45158 );
xor \g456216/U$11_r1 ( \45395 , \45394 , \45184 );
and \g456216/U$10 ( \45396 , \45393 , \45395 );
and \g456216/U$12 ( \45397 , \45386 , \45393 );
or \g456216/U$7 ( \45398 , \45389 , \45396 , \45397 );
xor \g133426/U$4 ( \45399 , \45328 , \45398 );
xor \g133513/U$1 ( \45400 , \45133 , \45187 );
xor \g133513/U$1_r1 ( \45401 , \45400 , \45237 );
and \g133426/U$3 ( \45402 , \45399 , \45401 );
and \g133426/U$5 ( \45403 , \45328 , \45398 );
or \g133426/U$2 ( \45404 , \45402 , \45403 );
xor \g133510/U$1 ( \45405 , \44936 , \44940 );
xor \g133510/U$1_r1 ( \45406 , \45405 , \44951 );
xor \g133305/U$4 ( \45407 , \45404 , \45406 );
xor \g133406/U$1 ( \45408 , \45121 , \45240 );
xor \g133406/U$1_r1 ( \45409 , \45408 , \45245 );
and \g133305/U$3 ( \45410 , \45407 , \45409 );
and \g133305/U$5 ( \45411 , \45404 , \45406 );
or \g133305/U$2 ( \45412 , \45410 , \45411 );
not \g131911/U$3 ( \45413 , \45412 );
xor \g456178/U$2 ( \45414 , \44963 , \44967 );
xor \g456178/U$1 ( \45415 , \45414 , \45089 );
xor \g456178/U$1_r1 ( \45416 , \45248 , \45255 );
xor \g456178/U$1_r2 ( \45417 , \45415 , \45416 );
not \g131911/U$4 ( \45418 , \45417 );
or \g131911/U$2 ( \45419 , \45413 , \45418 );
xor \g133305/U$1 ( \45420 , \45404 , \45406 );
xor \g133305/U$1_r1 ( \45421 , \45420 , \45409 );
xor \g456271/U$1 ( \45422 , \45353 , \45380 );
xor \g456271/U$1_r1 ( \45423 , \45422 , \45383 );
not \g134117/U$3 ( \45424 , \45299 );
not \g134117/U$4 ( \45425 , \45317 );
or \g134117/U$2 ( \45426 , \45424 , \45425 );
or \g134117/U$5 ( \45427 , \45299 , \45317 );
nand \g134117/U$1 ( \45428 , \45426 , \45427 );
not \g134082/U$3 ( \45429 , \45428 );
not \g134082/U$4 ( \45430 , \45306 );
and \g134082/U$2 ( \45431 , \45429 , \45430 );
and \g134082/U$5 ( \45432 , \45428 , \45306 );
nor \g134082/U$1 ( \45433 , \45431 , \45432 );
not \g133852/U$3 ( \45434 , \45433 );
and \g134817/U$2 ( \45435 , \41948 , \41107 );
and \g134817/U$3 ( \45436 , \41109 , \41947 );
nor \g134817/U$1 ( \45437 , \45435 , \45436 );
and \g134206/U$2 ( \45438 , \45437 , \41952 );
not \g134206/U$4 ( \45439 , \45437 );
and \g134206/U$3 ( \45440 , \45439 , \41755 );
nor \g134206/U$1 ( \45441 , \45438 , \45440 );
not \g134095/U$3 ( \45442 , \45441 );
and \g134907/U$2 ( \45443 , \40979 , \42609 );
and \g134907/U$3 ( \45444 , \42416 , \41071 );
nor \g134907/U$1 ( \45445 , \45443 , \45444 );
and \g134483/U$2 ( \45446 , \45445 , \40870 );
not \g134483/U$4 ( \45447 , \45445 );
and \g134483/U$3 ( \45448 , \45447 , \40871 );
nor \g134483/U$1 ( \45449 , \45446 , \45448 );
not \g134095/U$4 ( \45450 , \45449 );
and \g134095/U$2 ( \45451 , \45442 , \45450 );
and \g134106/U$2 ( \45452 , \45449 , \45441 );
and \g134853/U$2 ( \45453 , \41206 , \42344 );
and \g134853/U$3 ( \45454 , \41920 , \41208 );
nor \g134853/U$1 ( \45455 , \45453 , \45454 );
and \g134290/U$2 ( \45456 , \45455 , \41214 );
not \g134290/U$4 ( \45457 , \45455 );
and \g134290/U$3 ( \45458 , \45457 , \41215 );
nor \g134290/U$1 ( \45459 , \45456 , \45458 );
nor \g134106/U$1 ( \45460 , \45452 , \45459 );
nor \g134095/U$1 ( \45461 , \45451 , \45460 );
not \g133852/U$4 ( \45462 , \45461 );
and \g133852/U$2 ( \45463 , \45434 , \45462 );
and \g133857/U$2 ( \45464 , \45433 , \45461 );
xor \g133947/U$1 ( \45465 , \45335 , \45342 );
xor \g133947/U$1_r1 ( \45466 , \45465 , \45350 );
nor \g133857/U$1 ( \45467 , \45464 , \45466 );
nor \g133852/U$1 ( \45468 , \45463 , \45467 );
or \g133560/U$2 ( \45469 , \45423 , \45468 );
not \g133594/U$3 ( \45470 , \45468 );
not \g133594/U$4 ( \45471 , \45423 );
or \g133594/U$2 ( \45472 , \45470 , \45471 );
xor \g456266/U$2 ( \45473 , \45166 , \45173 );
xor \g456266/U$1 ( \45474 , \45473 , \45181 );
xor \g456266/U$1_r1 ( \45475 , \45264 , \45269 );
xor \g456266/U$1_r2 ( \45476 , \45474 , \45475 );
nand \g133594/U$1 ( \45477 , \45472 , \45476 );
nand \g133560/U$1 ( \45478 , \45469 , \45477 );
and \g134707/U$2 ( \45479 , \42644 , \40926 );
and \g134707/U$3 ( \45480 , \40800 , \42643 );
nor \g134707/U$1 ( \45481 , \45479 , \45480 );
and \g134587/U$2 ( \45482 , \45481 , \42487 );
not \g134587/U$4 ( \45483 , \45481 );
and \g134587/U$3 ( \45484 , \45483 , \42486 );
nor \g134587/U$1 ( \45485 , \45482 , \45484 );
and \g134999/U$2 ( \45486 , \41623 , \41345 );
and \g134999/U$3 ( \45487 , \41116 , \41745 );
nor \g134999/U$1 ( \45488 , \45486 , \45487 );
and \g134246/U$2 ( \45489 , \45488 , \41325 );
not \g134246/U$4 ( \45490 , \45488 );
and \g134246/U$3 ( \45491 , \45490 , \41324 );
nor \g134246/U$1 ( \45492 , \45489 , \45491 );
xor \g134018/U$4 ( \45493 , \45485 , \45492 );
and \g134910/U$2 ( \45494 , \41087 , \41774 );
and \g134910/U$3 ( \45495 , \41629 , \41328 );
nor \g134910/U$1 ( \45496 , \45494 , \45495 );
and \g134380/U$2 ( \45497 , \45496 , \41093 );
not \g134380/U$4 ( \45498 , \45496 );
and \g134380/U$3 ( \45499 , \45498 , \41092 );
nor \g134380/U$1 ( \45500 , \45497 , \45499 );
and \g134018/U$3 ( \45501 , \45493 , \45500 );
and \g134018/U$5 ( \45502 , \45485 , \45492 );
or \g134018/U$2 ( \45503 , \45501 , \45502 );
and \g135006/U$2 ( \45504 , \40513 , \43179 );
and \g135006/U$3 ( \45505 , \43183 , \40713 );
nor \g135006/U$1 ( \45506 , \45504 , \45505 );
and \g134512/U$2 ( \45507 , \45506 , \40521 );
not \g134512/U$4 ( \45508 , \45506 );
and \g134512/U$3 ( \45509 , \45508 , \40518 );
nor \g134512/U$1 ( \45510 , \45507 , \45509 );
and \g135302/U$2 ( \45511 , \43604 , \40525 );
and \g135302/U$3 ( \45512 , \40472 , \43603 );
nor \g135302/U$1 ( \45513 , \45511 , \45512 );
and \g135179/U$2 ( \45514 , \45513 , \42676 );
not \g135179/U$4 ( \45515 , \45513 );
and \g135179/U$3 ( \45516 , \45515 , \42675 );
nor \g135179/U$1 ( \45517 , \45514 , \45516 );
xor \g133930/U$4 ( \45518 , \45510 , \45517 );
and \g134712/U$2 ( \45519 , \40672 , \42701 );
and \g134712/U$3 ( \45520 , \42651 , \40858 );
nor \g134712/U$1 ( \45521 , \45519 , \45520 );
and \g134403/U$2 ( \45522 , \45521 , \40678 );
not \g134403/U$4 ( \45523 , \45521 );
and \g134403/U$3 ( \45524 , \45523 , \40677 );
nor \g134403/U$1 ( \45525 , \45522 , \45524 );
and \g133930/U$3 ( \45526 , \45518 , \45525 );
and \g133930/U$5 ( \45527 , \45510 , \45517 );
or \g133930/U$2 ( \45528 , \45526 , \45527 );
xor \g456214/U$5 ( \45529 , \45503 , \45528 );
and \g134834/U$2 ( \45530 , \42317 , \41144 );
and \g134834/U$3 ( \45531 , \40956 , \42316 );
nor \g134834/U$1 ( \45532 , \45530 , \45531 );
and \g134307/U$2 ( \45533 , \45532 , \42226 );
not \g134307/U$4 ( \45534 , \45532 );
and \g134307/U$3 ( \45535 , \45534 , \42225 );
nor \g134307/U$1 ( \45536 , \45533 , \45535 );
xor \g134003/U$4 ( \45537 , \45536 , \45275 );
and \g134973/U$2 ( \45538 , \43099 , \40731 );
and \g134973/U$3 ( \45539 , \40568 , \43101 );
nor \g134973/U$1 ( \45540 , \45538 , \45539 );
and \g134308/U$2 ( \45541 , \45540 , \42682 );
not \g134308/U$4 ( \45542 , \45540 );
and \g134308/U$3 ( \45543 , \45542 , \42681 );
nor \g134308/U$1 ( \45544 , \45541 , \45543 );
and \g134003/U$3 ( \45545 , \45537 , \45544 );
and \g134003/U$5 ( \45546 , \45536 , \45275 );
or \g134003/U$2 ( \45547 , \45545 , \45546 );
and \g456214/U$4 ( \45548 , \45529 , \45547 );
and \g456214/U$6 ( \45549 , \45503 , \45528 );
or \g456214/U$3 ( \45550 , \45548 , \45549 );
and \g134803/U$2 ( \45551 , \41087 , \41629 );
and \g134803/U$3 ( \45552 , \41345 , \41328 );
nor \g134803/U$1 ( \45553 , \45551 , \45552 );
and \g134298/U$2 ( \45554 , \45553 , \41093 );
not \g134298/U$4 ( \45555 , \45553 );
and \g134298/U$3 ( \45556 , \45555 , \41092 );
nor \g134298/U$1 ( \45557 , \45554 , \45556 );
and \g134740/U$2 ( \45558 , \41623 , \41116 );
and \g134740/U$3 ( \45559 , \41107 , \41745 );
nor \g134740/U$1 ( \45560 , \45558 , \45559 );
and \g134176/U$2 ( \45561 , \45560 , \41325 );
not \g134176/U$4 ( \45562 , \45560 );
and \g134176/U$3 ( \45563 , \45562 , \41324 );
nor \g134176/U$1 ( \45564 , \45561 , \45563 );
xor \g133850/U$4 ( \45565 , \45557 , \45564 );
xor \g134092/U$1 ( \45566 , \45276 , \45283 );
and \g133850/U$3 ( \45567 , \45565 , \45566 );
and \g133850/U$5 ( \45568 , \45557 , \45564 );
or \g133850/U$2 ( \45569 , \45567 , \45568 );
xor \g133516/U$4 ( \45570 , \45550 , \45569 );
xor \g133785/U$1 ( \45571 , \45284 , \45291 );
xor \g133785/U$1_r1 ( \45572 , \45571 , \45319 );
and \g133516/U$3 ( \45573 , \45570 , \45572 );
and \g133516/U$5 ( \45574 , \45550 , \45569 );
or \g133516/U$2 ( \45575 , \45573 , \45574 );
xor \g133402/U$4 ( \45576 , \45478 , \45575 );
xor \g133582/U$1 ( \45577 , \45274 , \45322 );
xor \g133582/U$1_r1 ( \45578 , \45577 , \45325 );
and \g133402/U$3 ( \45579 , \45576 , \45578 );
and \g133402/U$5 ( \45580 , \45478 , \45575 );
or \g133402/U$2 ( \45581 , \45579 , \45580 );
xor \g456225/U$2 ( \45582 , \44904 , \44906 );
xor \g456225/U$1 ( \45583 , \45582 , \44933 );
xor \g456225/U$1_r1 ( \45584 , \45109 , \45116 );
xor \g456225/U$1_r2 ( \45585 , \45583 , \45584 );
xor \g133307/U$4 ( \45586 , \45581 , \45585 );
xor \g133426/U$1 ( \45587 , \45328 , \45398 );
xor \g133426/U$1_r1 ( \45588 , \45587 , \45401 );
and \g133307/U$3 ( \45589 , \45586 , \45588 );
and \g133307/U$5 ( \45590 , \45581 , \45585 );
or \g133307/U$2 ( \45591 , \45589 , \45590 );
and \g131990/U$2 ( \45592 , \45421 , \45591 );
xor \g133278/U$1 ( \45593 , \45591 , \45421 );
not \g134081/U$3 ( \45594 , \45449 );
xor \g134125/U$1 ( \45595 , \45441 , \45459 );
not \g134081/U$4 ( \45596 , \45595 );
or \g134081/U$2 ( \45597 , \45594 , \45596 );
or \g134081/U$5 ( \45598 , \45595 , \45449 );
nand \g134081/U$1 ( \45599 , \45597 , \45598 );
and \g134936/U$2 ( \45600 , \42317 , \41109 );
and \g134936/U$3 ( \45601 , \41144 , \42316 );
nor \g134936/U$1 ( \45602 , \45600 , \45601 );
and \g134277/U$2 ( \45603 , \45602 , \42226 );
not \g134277/U$4 ( \45604 , \45602 );
and \g134277/U$3 ( \45605 , \45604 , \42225 );
nor \g134277/U$1 ( \45606 , \45603 , \45605 );
and \g134811/U$2 ( \45607 , \41206 , \42416 );
and \g134811/U$3 ( \45608 , \42344 , \41208 );
nor \g134811/U$1 ( \45609 , \45607 , \45608 );
and \g134495/U$2 ( \45610 , \45609 , \41215 );
not \g134495/U$4 ( \45611 , \45609 );
and \g134495/U$3 ( \45612 , \45611 , \41214 );
nor \g134495/U$1 ( \45613 , \45610 , \45612 );
xor \g456260/U$5 ( \45614 , \45606 , \45613 );
and \g134888/U$2 ( \45615 , \40979 , \42651 );
and \g134888/U$3 ( \45616 , \42609 , \41071 );
nor \g134888/U$1 ( \45617 , \45615 , \45616 );
and \g134549/U$2 ( \45618 , \45617 , \40871 );
not \g134549/U$4 ( \45619 , \45617 );
and \g134549/U$3 ( \45620 , \45619 , \40870 );
nor \g134549/U$1 ( \45621 , \45618 , \45620 );
and \g456260/U$4 ( \45622 , \45614 , \45621 );
and \g456260/U$6 ( \45623 , \45606 , \45613 );
or \g456260/U$3 ( \45624 , \45622 , \45623 );
xor \g133790/U$4 ( \45625 , \45599 , \45624 );
xor \g134018/U$1 ( \45626 , \45485 , \45492 );
xor \g134018/U$1_r1 ( \45627 , \45626 , \45500 );
and \g133790/U$3 ( \45628 , \45625 , \45627 );
and \g133790/U$5 ( \45629 , \45599 , \45624 );
or \g133790/U$2 ( \45630 , \45628 , \45629 );
xor \g456214/U$9 ( \45631 , \45503 , \45528 );
xor \g456214/U$9_r1 ( \45632 , \45631 , \45547 );
and \g456214/U$8 ( \45633 , \45630 , \45632 );
not \g133829/U$3 ( \45634 , \45433 );
xor \g133871/U$1 ( \45635 , \45461 , \45466 );
not \g133829/U$4 ( \45636 , \45635 );
or \g133829/U$2 ( \45637 , \45634 , \45636 );
or \g133829/U$5 ( \45638 , \45635 , \45433 );
nand \g133829/U$1 ( \45639 , \45637 , \45638 );
xor \g456214/U$11 ( \45640 , \45503 , \45528 );
xor \g456214/U$11_r1 ( \45641 , \45640 , \45547 );
and \g456214/U$10 ( \45642 , \45639 , \45641 );
and \g456214/U$12 ( \45643 , \45630 , \45639 );
or \g456214/U$7 ( \45644 , \45633 , \45642 , \45643 );
and \g134794/U$2 ( \45645 , \42644 , \40956 );
and \g134794/U$3 ( \45646 , \40926 , \42643 );
nor \g134794/U$1 ( \45647 , \45645 , \45646 );
or \g134151/U$2 ( \45648 , \45647 , \42486 );
nand \g134637/U$1 ( \45649 , \42486 , \45647 );
nand \g134151/U$1 ( \45650 , \45648 , \45649 );
and \g135292/U$2 ( \45651 , \43604 , \40568 );
and \g135292/U$3 ( \45652 , \40525 , \43603 );
nor \g135292/U$1 ( \45653 , \45651 , \45652 );
and \g135192/U$2 ( \45654 , \45653 , \42676 );
not \g135192/U$4 ( \45655 , \45653 );
and \g135192/U$3 ( \45656 , \45655 , \42675 );
nor \g135192/U$1 ( \45657 , \45654 , \45656 );
xor \g133965/U$4 ( \45658 , \45650 , \45657 );
and \g135040/U$2 ( \45659 , \41623 , \41629 );
and \g135040/U$3 ( \45660 , \41345 , \41745 );
nor \g135040/U$1 ( \45661 , \45659 , \45660 );
and \g134472/U$2 ( \45662 , \45661 , \41325 );
not \g134472/U$4 ( \45663 , \45661 );
and \g134472/U$3 ( \45664 , \45663 , \41324 );
nor \g134472/U$1 ( \45665 , \45662 , \45664 );
and \g133965/U$3 ( \45666 , \45658 , \45665 );
and \g133965/U$5 ( \45667 , \45650 , \45657 );
or \g133965/U$2 ( \45668 , \45666 , \45667 );
nor \g135219/U$1 ( \45669 , \40508 , \43607 );
nor \g135171/U$1 ( \45670 , \45669 , \40521 );
and \g134772/U$2 ( \45671 , \43099 , \40800 );
and \g134772/U$3 ( \45672 , \40731 , \43101 );
nor \g134772/U$1 ( \45673 , \45671 , \45672 );
and \g134491/U$2 ( \45674 , \45673 , \42682 );
not \g134491/U$4 ( \45675 , \45673 );
and \g134491/U$3 ( \45676 , \45675 , \42681 );
nor \g134491/U$1 ( \45677 , \45674 , \45676 );
and \g134093/U$2 ( \45678 , \45670 , \45677 );
xor \g133773/U$4 ( \45679 , \45668 , \45678 );
and \g135080/U$2 ( \45680 , \41948 , \41116 );
and \g135080/U$3 ( \45681 , \41107 , \41947 );
nor \g135080/U$1 ( \45682 , \45680 , \45681 );
and \g134273/U$2 ( \45683 , \45682 , \41755 );
not \g134273/U$4 ( \45684 , \45682 );
and \g134273/U$3 ( \45685 , \45684 , \41952 );
nor \g134273/U$1 ( \45686 , \45683 , \45685 );
and \g135142/U$2 ( \45687 , \40672 , \43183 );
and \g135142/U$3 ( \45688 , \42701 , \40858 );
nor \g135142/U$1 ( \45689 , \45687 , \45688 );
and \g134584/U$2 ( \45690 , \45689 , \40678 );
not \g134584/U$4 ( \45691 , \45689 );
and \g134584/U$3 ( \45692 , \45691 , \40677 );
nor \g134584/U$1 ( \45693 , \45690 , \45692 );
xor \g133950/U$4 ( \45694 , \45686 , \45693 );
and \g135067/U$2 ( \45695 , \40513 , \43757 );
and \g135067/U$3 ( \45696 , \43179 , \40713 );
nor \g135067/U$1 ( \45697 , \45695 , \45696 );
and \g134536/U$2 ( \45698 , \45697 , \40521 );
not \g134536/U$4 ( \45699 , \45697 );
and \g134536/U$3 ( \45700 , \45699 , \40518 );
nor \g134536/U$1 ( \45701 , \45698 , \45700 );
and \g133950/U$3 ( \45702 , \45694 , \45701 );
and \g133950/U$5 ( \45703 , \45686 , \45693 );
or \g133950/U$2 ( \45704 , \45702 , \45703 );
and \g133773/U$3 ( \45705 , \45679 , \45704 );
and \g133773/U$5 ( \45706 , \45668 , \45678 );
or \g133773/U$2 ( \45707 , \45705 , \45706 );
not \g134080/U$3 ( \45708 , \45368 );
xor \g134128/U$1 ( \45709 , \45360 , \45378 );
not \g134080/U$4 ( \45710 , \45709 );
or \g134080/U$2 ( \45711 , \45708 , \45710 );
or \g134080/U$5 ( \45712 , \45709 , \45368 );
nand \g134080/U$1 ( \45713 , \45711 , \45712 );
xor \g133584/U$4 ( \45714 , \45707 , \45713 );
xor \g133850/U$1 ( \45715 , \45557 , \45564 );
xor \g133850/U$1_r1 ( \45716 , \45715 , \45566 );
and \g133584/U$3 ( \45717 , \45714 , \45716 );
and \g133584/U$5 ( \45718 , \45707 , \45713 );
or \g133584/U$2 ( \45719 , \45717 , \45718 );
xor \g133428/U$4 ( \45720 , \45644 , \45719 );
xor \g133516/U$1 ( \45721 , \45550 , \45569 );
xor \g133516/U$1_r1 ( \45722 , \45721 , \45572 );
and \g133428/U$3 ( \45723 , \45720 , \45722 );
and \g133428/U$5 ( \45724 , \45644 , \45719 );
or \g133428/U$2 ( \45725 , \45723 , \45724 );
xor \g456216/U$2 ( \45726 , \45157 , \45158 );
xor \g456216/U$1 ( \45727 , \45726 , \45184 );
xor \g456216/U$1_r1 ( \45728 , \45386 , \45393 );
xor \g456216/U$1_r2 ( \45729 , \45727 , \45728 );
xor \g133308/U$4 ( \45730 , \45725 , \45729 );
xor \g133402/U$1 ( \45731 , \45478 , \45575 );
xor \g133402/U$1_r1 ( \45732 , \45731 , \45578 );
and \g133308/U$3 ( \45733 , \45730 , \45732 );
and \g133308/U$5 ( \45734 , \45725 , \45729 );
or \g133308/U$2 ( \45735 , \45733 , \45734 );
not \g132057/U$3 ( \45736 , \45735 );
xor \g133307/U$1 ( \45737 , \45581 , \45585 );
xor \g133307/U$1_r1 ( \45738 , \45737 , \45588 );
not \g132057/U$4 ( \45739 , \45738 );
or \g132057/U$2 ( \45740 , \45736 , \45739 );
and \g134800/U$2 ( \45741 , \41087 , \42416 );
and \g134800/U$3 ( \45742 , \42344 , \41328 );
nor \g134800/U$1 ( \45743 , \45741 , \45742 );
and \g134520/U$2 ( \45744 , \45743 , \41093 );
not \g134520/U$4 ( \45745 , \45743 );
and \g134520/U$3 ( \45746 , \45745 , \41092 );
nor \g134520/U$1 ( \45747 , \45744 , \45746 );
and \g134751/U$2 ( \45748 , \42644 , \41109 );
and \g134751/U$3 ( \45749 , \41144 , \42643 );
nor \g134751/U$1 ( \45750 , \45748 , \45749 );
and \g134519/U$2 ( \45751 , \45750 , \42487 );
not \g134519/U$4 ( \45752 , \45750 );
and \g134519/U$3 ( \45753 , \45752 , \42486 );
nor \g134519/U$1 ( \45754 , \45751 , \45753 );
xor \g133911/U$4 ( \45755 , \45747 , \45754 );
and \g134868/U$2 ( \45756 , \41623 , \41920 );
and \g134868/U$3 ( \45757 , \41774 , \41745 );
nor \g134868/U$1 ( \45758 , \45756 , \45757 );
and \g134336/U$2 ( \45759 , \45758 , \41325 );
not \g134336/U$4 ( \45760 , \45758 );
and \g134336/U$3 ( \45761 , \45760 , \41324 );
nor \g134336/U$1 ( \45762 , \45759 , \45761 );
and \g133911/U$3 ( \45763 , \45755 , \45762 );
and \g133911/U$5 ( \45764 , \45747 , \45754 );
or \g133911/U$2 ( \45765 , \45763 , \45764 );
and \g134721/U$2 ( \45766 , \40979 , \43183 );
and \g134721/U$3 ( \45767 , \42701 , \41071 );
nor \g134721/U$1 ( \45768 , \45766 , \45767 );
and \g134257/U$2 ( \45769 , \45768 , \40871 );
not \g134257/U$4 ( \45770 , \45768 );
and \g134257/U$3 ( \45771 , \45770 , \40870 );
nor \g134257/U$1 ( \45772 , \45769 , \45771 );
and \g134680/U$2 ( \45773 , \42317 , \41116 );
and \g134680/U$3 ( \45774 , \41107 , \42316 );
nor \g134680/U$1 ( \45775 , \45773 , \45774 );
and \g134516/U$2 ( \45776 , \45775 , \42226 );
not \g134516/U$4 ( \45777 , \45775 );
and \g134516/U$3 ( \45778 , \45777 , \42225 );
nor \g134516/U$1 ( \45779 , \45776 , \45778 );
xor \g133932/U$4 ( \45780 , \45772 , \45779 );
and \g134785/U$2 ( \45781 , \41206 , \42651 );
and \g134785/U$3 ( \45782 , \42609 , \41208 );
nor \g134785/U$1 ( \45783 , \45781 , \45782 );
and \g134518/U$2 ( \45784 , \45783 , \41215 );
not \g134518/U$4 ( \45785 , \45783 );
and \g134518/U$3 ( \45786 , \45785 , \41214 );
nor \g134518/U$1 ( \45787 , \45784 , \45786 );
and \g133932/U$3 ( \45788 , \45780 , \45787 );
and \g133932/U$5 ( \45789 , \45772 , \45779 );
or \g133932/U$2 ( \45790 , \45788 , \45789 );
xor \g456207/U$2 ( \45791 , \45765 , \45790 );
and \g134787/U$2 ( \45792 , \41948 , \41629 );
and \g134787/U$3 ( \45793 , \41345 , \41947 );
nor \g134787/U$1 ( \45794 , \45792 , \45793 );
and \g134453/U$2 ( \45795 , \45794 , \41952 );
not \g134453/U$4 ( \45796 , \45794 );
and \g134453/U$3 ( \45797 , \45796 , \41755 );
nor \g134453/U$1 ( \45798 , \45795 , \45797 );
and \g134702/U$2 ( \45799 , \43099 , \40956 );
and \g134702/U$3 ( \45800 , \40926 , \43101 );
nor \g134702/U$1 ( \45801 , \45799 , \45800 );
and \g134294/U$2 ( \45802 , \45801 , \42681 );
not \g134294/U$4 ( \45803 , \45801 );
and \g134294/U$3 ( \45804 , \45803 , \42682 );
nor \g134294/U$1 ( \45805 , \45802 , \45804 );
xor \g456275/U$4 ( \45806 , \45798 , \45805 );
and \g134769/U$2 ( \45807 , \40672 , \43757 );
and \g134769/U$3 ( \45808 , \43179 , \40858 );
nor \g134769/U$1 ( \45809 , \45807 , \45808 );
and \g134565/U$2 ( \45810 , \45809 , \40677 );
not \g134565/U$4 ( \45811 , \45809 );
and \g134565/U$3 ( \45812 , \45811 , \40678 );
nor \g134565/U$1 ( \45813 , \45810 , \45812 );
and \g456275/U$3 ( \45814 , \45806 , \45813 );
and \g456275/U$5 ( \45815 , \45798 , \45805 );
nor \g456275/U$2 ( \45816 , \45814 , \45815 );
xor \g456207/U$1 ( \45817 , \45791 , \45816 );
and \g135309/U$2 ( \45818 , \43604 , \40731 );
and \g135309/U$3 ( \45819 , \40568 , \43603 );
nor \g135309/U$1 ( \45820 , \45818 , \45819 );
and \g135182/U$2 ( \45821 , \45820 , \42676 );
not \g135182/U$4 ( \45822 , \45820 );
and \g135182/U$3 ( \45823 , \45822 , \42675 );
nor \g135182/U$1 ( \45824 , \45821 , \45823 );
xor \g456257/U$2 ( \45825 , \45824 , \45669 );
and \g135013/U$2 ( \45826 , \42317 , \41107 );
and \g135013/U$3 ( \45827 , \41109 , \42316 );
nor \g135013/U$1 ( \45828 , \45826 , \45827 );
and \g134230/U$2 ( \45829 , \45828 , \42226 );
not \g134230/U$4 ( \45830 , \45828 );
and \g134230/U$3 ( \45831 , \45830 , \42225 );
nor \g134230/U$1 ( \45832 , \45829 , \45831 );
xor \g456257/U$1 ( \45833 , \45825 , \45832 );
and \g135101/U$2 ( \45834 , \40672 , \43179 );
and \g135101/U$3 ( \45835 , \43183 , \40858 );
nor \g135101/U$1 ( \45836 , \45834 , \45835 );
and \g134523/U$2 ( \45837 , \45836 , \40678 );
not \g134523/U$4 ( \45838 , \45836 );
and \g134523/U$3 ( \45839 , \45838 , \40677 );
nor \g134523/U$1 ( \45840 , \45837 , \45839 );
and \g134940/U$2 ( \45841 , \42644 , \41144 );
and \g134940/U$3 ( \45842 , \40956 , \42643 );
nor \g134940/U$1 ( \45843 , \45841 , \45842 );
and \g134280/U$2 ( \45844 , \45843 , \42487 );
not \g134280/U$4 ( \45845 , \45843 );
and \g134280/U$3 ( \45846 , \45845 , \42486 );
nor \g134280/U$1 ( \45847 , \45844 , \45846 );
xor \g133896/U$1 ( \45848 , \45840 , \45847 );
and \g135131/U$2 ( \45849 , \41948 , \41345 );
and \g135131/U$3 ( \45850 , \41116 , \41947 );
nor \g135131/U$1 ( \45851 , \45849 , \45850 );
and \g134557/U$2 ( \45852 , \45851 , \41755 );
not \g134557/U$4 ( \45853 , \45851 );
and \g134557/U$3 ( \45854 , \45853 , \41952 );
nor \g134557/U$1 ( \45855 , \45852 , \45854 );
xor \g133896/U$1_r1 ( \45856 , \45848 , \45855 );
and \g135077/U$2 ( \45857 , \40979 , \42701 );
and \g135077/U$3 ( \45858 , \42651 , \41071 );
nor \g135077/U$1 ( \45859 , \45857 , \45858 );
and \g134227/U$2 ( \45860 , \45859 , \40871 );
not \g134227/U$4 ( \45861 , \45859 );
and \g134227/U$3 ( \45862 , \45861 , \40870 );
nor \g134227/U$1 ( \45863 , \45860 , \45862 );
and \g134975/U$2 ( \45864 , \41206 , \42609 );
and \g134975/U$3 ( \45865 , \42416 , \41208 );
nor \g134975/U$1 ( \45866 , \45864 , \45865 );
and \g134345/U$2 ( \45867 , \45866 , \41215 );
not \g134345/U$4 ( \45868 , \45866 );
and \g134345/U$3 ( \45869 , \45868 , \41214 );
nor \g134345/U$1 ( \45870 , \45867 , \45869 );
xor \g133998/U$1 ( \45871 , \45863 , \45870 );
and \g135129/U$2 ( \45872 , \43099 , \40926 );
and \g135129/U$3 ( \45873 , \40800 , \43101 );
nor \g135129/U$1 ( \45874 , \45872 , \45873 );
and \g134311/U$2 ( \45875 , \45874 , \42682 );
not \g134311/U$4 ( \45876 , \45874 );
and \g134311/U$3 ( \45877 , \45876 , \42681 );
nor \g134311/U$1 ( \45878 , \45875 , \45877 );
xor \g133998/U$1_r1 ( \45879 , \45871 , \45878 );
xor \g456257/U$1_r1 ( \45880 , \45856 , \45879 );
xor \g456257/U$1_r2 ( \45881 , \45833 , \45880 );
and \g135100/U$2 ( \45882 , \41623 , \41774 );
and \g135100/U$3 ( \45883 , \41629 , \41745 );
nor \g135100/U$1 ( \45884 , \45882 , \45883 );
and \g134576/U$2 ( \45885 , \45884 , \41325 );
not \g134576/U$4 ( \45886 , \45884 );
and \g134576/U$3 ( \45887 , \45886 , \41324 );
nor \g134576/U$1 ( \45888 , \45885 , \45887 );
nor \g135214/U$1 ( \45889 , \40666 , \43607 );
nor \g135172/U$1 ( \45890 , \45889 , \40678 );
and \g135312/U$2 ( \45891 , \43604 , \40800 );
and \g135312/U$3 ( \45892 , \40731 , \43603 );
nor \g135312/U$1 ( \45893 , \45891 , \45892 );
and \g135181/U$2 ( \45894 , \45893 , \42676 );
not \g135181/U$4 ( \45895 , \45893 );
and \g135181/U$3 ( \45896 , \45895 , \42675 );
nor \g135181/U$1 ( \45897 , \45894 , \45896 );
and \g134625/U$2 ( \45898 , \45890 , \45897 );
xor \g133973/U$1 ( \45899 , \45888 , \45898 );
and \g135070/U$2 ( \45900 , \41087 , \42344 );
and \g135070/U$3 ( \45901 , \41920 , \41328 );
nor \g135070/U$1 ( \45902 , \45900 , \45901 );
and \g134341/U$2 ( \45903 , \45902 , \41093 );
not \g134341/U$4 ( \45904 , \45902 );
and \g134341/U$3 ( \45905 , \45904 , \41092 );
nor \g134341/U$1 ( \45906 , \45903 , \45905 );
xor \g133973/U$1_r1 ( \45907 , \45899 , \45906 );
and \g135298/U$2 ( \45908 , \43604 , \40926 );
and \g135298/U$3 ( \45909 , \40800 , \43603 );
nor \g135298/U$1 ( \45910 , \45908 , \45909 );
and \g135189/U$2 ( \45911 , \45910 , \42676 );
not \g135189/U$4 ( \45912 , \45910 );
and \g135189/U$3 ( \45913 , \45912 , \42675 );
nor \g135189/U$1 ( \45914 , \45911 , \45913 );
xor \g456270/U$5 ( \45915 , \45914 , \45889 );
and \g134877/U$2 ( \45916 , \42317 , \41345 );
and \g134877/U$3 ( \45917 , \41116 , \42316 );
nor \g134877/U$1 ( \45918 , \45916 , \45917 );
and \g134544/U$2 ( \45919 , \45918 , \42226 );
not \g134544/U$4 ( \45920 , \45918 );
and \g134544/U$3 ( \45921 , \45920 , \42225 );
nor \g134544/U$1 ( \45922 , \45919 , \45921 );
and \g456270/U$4 ( \45923 , \45915 , \45922 );
and \g456270/U$6 ( \45924 , \45914 , \45889 );
or \g456270/U$3 ( \45925 , \45923 , \45924 );
xor \g134625/U$1 ( \45926 , \45890 , \45897 );
xor \g133778/U$4 ( \45927 , \45925 , \45926 );
and \g134871/U$2 ( \45928 , \41206 , \42701 );
and \g134871/U$3 ( \45929 , \42651 , \41208 );
nor \g134871/U$1 ( \45930 , \45928 , \45929 );
and \g134214/U$2 ( \45931 , \45930 , \41215 );
not \g134214/U$4 ( \45932 , \45930 );
and \g134214/U$3 ( \45933 , \45932 , \41214 );
nor \g134214/U$1 ( \45934 , \45931 , \45933 );
and \g134905/U$2 ( \45935 , \40979 , \43179 );
and \g134905/U$3 ( \45936 , \43183 , \41071 );
nor \g134905/U$1 ( \45937 , \45935 , \45936 );
and \g134543/U$2 ( \45938 , \45937 , \40871 );
not \g134543/U$4 ( \45939 , \45937 );
and \g134543/U$3 ( \45940 , \45939 , \40870 );
nor \g134543/U$1 ( \45941 , \45938 , \45940 );
xor \g456237/U$5 ( \45942 , \45934 , \45941 );
and \g134845/U$2 ( \45943 , \43099 , \41144 );
and \g134845/U$3 ( \45944 , \40956 , \43101 );
nor \g134845/U$1 ( \45945 , \45943 , \45944 );
or \g134153/U$2 ( \45946 , \45945 , \42681 );
nand \g134636/U$1 ( \45947 , \42681 , \45945 );
nand \g134153/U$1 ( \45948 , \45946 , \45947 );
and \g456237/U$4 ( \45949 , \45942 , \45948 );
and \g456237/U$6 ( \45950 , \45934 , \45941 );
or \g456237/U$3 ( \45951 , \45949 , \45950 );
and \g133778/U$3 ( \45952 , \45927 , \45951 );
and \g133778/U$5 ( \45953 , \45925 , \45926 );
or \g133778/U$2 ( \45954 , \45952 , \45953 );
not \g133619/U$3 ( \45955 , \45954 );
xor \g133911/U$1 ( \45956 , \45747 , \45754 );
xor \g133911/U$1_r1 ( \45957 , \45956 , \45762 );
and \g134797/U$2 ( \45958 , \41623 , \42344 );
and \g134797/U$3 ( \45959 , \41920 , \41745 );
nor \g134797/U$1 ( \45960 , \45958 , \45959 );
and \g134546/U$2 ( \45961 , \45960 , \41325 );
not \g134546/U$4 ( \45962 , \45960 );
and \g134546/U$3 ( \45963 , \45962 , \41324 );
nor \g134546/U$1 ( \45964 , \45961 , \45963 );
and \g135076/U$2 ( \45965 , \42644 , \41107 );
and \g135076/U$3 ( \45966 , \41109 , \42643 );
nor \g135076/U$1 ( \45967 , \45965 , \45966 );
and \g134603/U$2 ( \45968 , \45967 , \42487 );
not \g134603/U$4 ( \45969 , \45967 );
and \g134603/U$3 ( \45970 , \45969 , \42486 );
nor \g134603/U$1 ( \45971 , \45968 , \45970 );
xor \g133887/U$4 ( \45972 , \45964 , \45971 );
and \g135141/U$2 ( \45973 , \41948 , \41774 );
and \g135141/U$3 ( \45974 , \41629 , \41947 );
nor \g135141/U$1 ( \45975 , \45973 , \45974 );
and \g134225/U$2 ( \45976 , \45975 , \41755 );
not \g134225/U$4 ( \45977 , \45975 );
and \g134225/U$3 ( \45978 , \45977 , \41952 );
nor \g134225/U$1 ( \45979 , \45976 , \45978 );
and \g133887/U$3 ( \45980 , \45972 , \45979 );
and \g133887/U$5 ( \45981 , \45964 , \45971 );
or \g133887/U$2 ( \45982 , \45980 , \45981 );
xor \g456258/U$4 ( \45983 , \45957 , \45982 );
xor \g133932/U$1 ( \45984 , \45772 , \45779 );
xor \g133932/U$1_r1 ( \45985 , \45984 , \45787 );
and \g456258/U$3 ( \45986 , \45983 , \45985 );
and \g456258/U$5 ( \45987 , \45957 , \45982 );
nor \g456258/U$2 ( \45988 , \45986 , \45987 );
not \g133619/U$4 ( \45989 , \45988 );
or \g133619/U$2 ( \45990 , \45955 , \45989 );
or \g133619/U$5 ( \45991 , \45988 , \45954 );
nand \g133619/U$1 ( \45992 , \45990 , \45991 );
xor \g455959/U$1 ( \45993 , \45907 , \45992 );
xor \g456207/U$1_r1 ( \45994 , \45881 , \45993 );
xor \g456207/U$1_r2 ( \45995 , \45817 , \45994 );
not \g133394/U$3 ( \45996 , \45995 );
and \g134862/U$2 ( \45997 , \41087 , \42609 );
and \g134862/U$3 ( \45998 , \42416 , \41328 );
nor \g134862/U$1 ( \45999 , \45997 , \45998 );
and \g134320/U$2 ( \46000 , \45999 , \41092 );
not \g134320/U$4 ( \46001 , \45999 );
and \g134320/U$3 ( \46002 , \46001 , \41093 );
nor \g134320/U$1 ( \46003 , \46000 , \46002 );
not \g133877/U$3 ( \46004 , \46003 );
and \g135301/U$2 ( \46005 , \43604 , \40956 );
and \g135301/U$3 ( \46006 , \40926 , \43603 );
nor \g135301/U$1 ( \46007 , \46005 , \46006 );
and \g135175/U$2 ( \46008 , \46007 , \42675 );
not \g135175/U$4 ( \46009 , \46007 );
and \g135175/U$3 ( \46010 , \46009 , \42676 );
nor \g135175/U$1 ( \46011 , \46008 , \46010 );
not \g134675/U$2 ( \46012 , \46011 );
nor \g135210/U$1 ( \46013 , \40973 , \43607 );
nor \g135168/U$1 ( \46014 , \46013 , \40871 );
nand \g134675/U$1 ( \46015 , \46012 , \46014 );
not \g133877/U$4 ( \46016 , \46015 );
and \g133877/U$2 ( \46017 , \46004 , \46016 );
and \g133885/U$2 ( \46018 , \46003 , \46015 );
and \g134805/U$2 ( \46019 , \42317 , \41629 );
and \g134805/U$3 ( \46020 , \41345 , \42316 );
nor \g134805/U$1 ( \46021 , \46019 , \46020 );
and \g134447/U$2 ( \46022 , \46021 , \42225 );
not \g134447/U$4 ( \46023 , \46021 );
and \g134447/U$3 ( \46024 , \46023 , \42226 );
nor \g134447/U$1 ( \46025 , \46022 , \46024 );
and \g134703/U$2 ( \46026 , \40979 , \43757 );
and \g134703/U$3 ( \46027 , \43179 , \41071 );
nor \g134703/U$1 ( \46028 , \46026 , \46027 );
and \g134397/U$2 ( \46029 , \46028 , \40870 );
not \g134397/U$4 ( \46030 , \46028 );
and \g134397/U$3 ( \46031 , \46030 , \40871 );
nor \g134397/U$1 ( \46032 , \46029 , \46031 );
or \g134099/U$2 ( \46033 , \46025 , \46032 );
not \g134110/U$3 ( \46034 , \46032 );
not \g134110/U$4 ( \46035 , \46025 );
or \g134110/U$2 ( \46036 , \46034 , \46035 );
and \g134982/U$2 ( \46037 , \41206 , \43183 );
and \g134982/U$3 ( \46038 , \42701 , \41208 );
nor \g134982/U$1 ( \46039 , \46037 , \46038 );
and \g134525/U$2 ( \46040 , \46039 , \41215 );
not \g134525/U$4 ( \46041 , \46039 );
and \g134525/U$3 ( \46042 , \46041 , \41214 );
nor \g134525/U$1 ( \46043 , \46040 , \46042 );
nand \g134110/U$1 ( \46044 , \46036 , \46043 );
nand \g134099/U$1 ( \46045 , \46033 , \46044 );
not \g134020/U$1 ( \46046 , \46045 );
nor \g133885/U$1 ( \46047 , \46018 , \46046 );
nor \g133877/U$1 ( \46048 , \46017 , \46047 );
xor \g456275/U$1 ( \46049 , \45798 , \45805 );
xor \g456275/U$1_r1 ( \46050 , \46049 , \45813 );
or \g133605/U$2 ( \46051 , \46048 , \46050 );
not \g133618/U$3 ( \46052 , \46050 );
not \g133618/U$4 ( \46053 , \46048 );
or \g133618/U$2 ( \46054 , \46052 , \46053 );
xor \g133778/U$1 ( \46055 , \45925 , \45926 );
xor \g133778/U$1_r1 ( \46056 , \46055 , \45951 );
nand \g133618/U$1 ( \46057 , \46054 , \46056 );
nand \g133605/U$1 ( \46058 , \46051 , \46057 );
xor \g456258/U$1 ( \46059 , \45957 , \45982 );
xor \g456258/U$1_r1 ( \46060 , \46059 , \45985 );
and \g134922/U$2 ( \46061 , \41948 , \41920 );
and \g134922/U$3 ( \46062 , \41774 , \41947 );
nor \g134922/U$1 ( \46063 , \46061 , \46062 );
and \g134559/U$2 ( \46064 , \46063 , \41755 );
not \g134559/U$4 ( \46065 , \46063 );
and \g134559/U$3 ( \46066 , \46065 , \41952 );
nor \g134559/U$1 ( \46067 , \46064 , \46066 );
and \g134777/U$2 ( \46068 , \42644 , \41116 );
and \g134777/U$3 ( \46069 , \41107 , \42643 );
nor \g134777/U$1 ( \46070 , \46068 , \46069 );
and \g134541/U$2 ( \46071 , \46070 , \42487 );
not \g134541/U$4 ( \46072 , \46070 );
and \g134541/U$3 ( \46073 , \46072 , \42486 );
nor \g134541/U$1 ( \46074 , \46071 , \46073 );
xor \g134012/U$4 ( \46075 , \46067 , \46074 );
and \g135018/U$2 ( \46076 , \43099 , \41109 );
and \g135018/U$3 ( \46077 , \41144 , \43101 );
nor \g135018/U$1 ( \46078 , \46076 , \46077 );
and \g134561/U$2 ( \46079 , \46078 , \42682 );
not \g134561/U$4 ( \46080 , \46078 );
and \g134561/U$3 ( \46081 , \46080 , \42681 );
nor \g134561/U$1 ( \46082 , \46079 , \46081 );
and \g134012/U$3 ( \46083 , \46075 , \46082 );
and \g134012/U$5 ( \46084 , \46067 , \46074 );
or \g134012/U$2 ( \46085 , \46083 , \46084 );
xor \g456270/U$9 ( \46086 , \45914 , \45889 );
xor \g456270/U$9_r1 ( \46087 , \46086 , \45922 );
and \g456270/U$8 ( \46088 , \46085 , \46087 );
xor \g133887/U$1 ( \46089 , \45964 , \45971 );
xor \g133887/U$1_r1 ( \46090 , \46089 , \45979 );
xor \g456270/U$11 ( \46091 , \45914 , \45889 );
xor \g456270/U$11_r1 ( \46092 , \46091 , \45922 );
and \g456270/U$10 ( \46093 , \46090 , \46092 );
and \g456270/U$12 ( \46094 , \46085 , \46090 );
or \g456270/U$7 ( \46095 , \46088 , \46093 , \46094 );
xor \g133519/U$4 ( \46096 , \46060 , \46095 );
not \g134669/U$3 ( \46097 , \46011 );
not \g134669/U$4 ( \46098 , \46014 );
and \g134669/U$2 ( \46099 , \46097 , \46098 );
and \g134669/U$5 ( \46100 , \46011 , \46014 );
nor \g134669/U$1 ( \46101 , \46099 , \46100 );
and \g134821/U$2 ( \46102 , \41623 , \42416 );
and \g134821/U$3 ( \46103 , \42344 , \41745 );
nor \g134821/U$1 ( \46104 , \46102 , \46103 );
and \g134164/U$2 ( \46105 , \46104 , \41324 );
nor \g134643/U$1 ( \46106 , \46104 , \41324 );
nor \g134164/U$1 ( \46107 , \46105 , \46106 );
xor \g456276/U$4 ( \46108 , \46101 , \46107 );
and \g135098/U$2 ( \46109 , \41087 , \42651 );
and \g135098/U$3 ( \46110 , \42609 , \41328 );
nor \g135098/U$1 ( \46111 , \46109 , \46110 );
and \g134334/U$2 ( \46112 , \46111 , \41092 );
not \g134334/U$4 ( \46113 , \46111 );
and \g134334/U$3 ( \46114 , \46113 , \41093 );
nor \g134334/U$1 ( \46115 , \46112 , \46114 );
and \g456276/U$3 ( \46116 , \46108 , \46115 );
and \g456276/U$5 ( \46117 , \46101 , \46107 );
nor \g456276/U$2 ( \46118 , \46116 , \46117 );
xor \g456237/U$9 ( \46119 , \45934 , \45941 );
xor \g456237/U$9_r1 ( \46120 , \46119 , \45948 );
and \g456237/U$8 ( \46121 , \46118 , \46120 );
not \g133831/U$3 ( \46122 , \46003 );
not \g133870/U$3 ( \46123 , \46015 );
not \g133870/U$4 ( \46124 , \46045 );
or \g133870/U$2 ( \46125 , \46123 , \46124 );
or \g133870/U$5 ( \46126 , \46045 , \46015 );
nand \g133870/U$1 ( \46127 , \46125 , \46126 );
not \g133831/U$4 ( \46128 , \46127 );
or \g133831/U$2 ( \46129 , \46122 , \46128 );
or \g133831/U$5 ( \46130 , \46127 , \46003 );
nand \g133831/U$1 ( \46131 , \46129 , \46130 );
xor \g456237/U$11 ( \46132 , \45934 , \45941 );
xor \g456237/U$11_r1 ( \46133 , \46132 , \45948 );
and \g456237/U$10 ( \46134 , \46131 , \46133 );
and \g456237/U$12 ( \46135 , \46118 , \46131 );
or \g456237/U$7 ( \46136 , \46121 , \46134 , \46135 );
and \g133519/U$3 ( \46137 , \46096 , \46136 );
and \g133519/U$5 ( \46138 , \46060 , \46095 );
or \g133519/U$2 ( \46139 , \46137 , \46138 );
xnor \g133465/U$1 ( \46140 , \46058 , \46139 );
not \g133394/U$4 ( \46141 , \46140 );
or \g133394/U$2 ( \46142 , \45996 , \46141 );
or \g133394/U$5 ( \46143 , \46140 , \45995 );
nand \g133394/U$1 ( \46144 , \46142 , \46143 );
xor \g456270/U$2 ( \46145 , \45914 , \45889 );
xor \g456270/U$1 ( \46146 , \46145 , \45922 );
xor \g456270/U$1_r1 ( \46147 , \46085 , \46090 );
xor \g456270/U$1_r2 ( \46148 , \46146 , \46147 );
and \g135088/U$2 ( \46149 , \41623 , \42609 );
and \g135088/U$3 ( \46150 , \42416 , \41745 );
nor \g135088/U$1 ( \46151 , \46149 , \46150 );
and \g134373/U$2 ( \46152 , \46151 , \41325 );
not \g134373/U$4 ( \46153 , \46151 );
and \g134373/U$3 ( \46154 , \46153 , \41324 );
nor \g134373/U$1 ( \46155 , \46152 , \46154 );
and \g135121/U$2 ( \46156 , \42644 , \41345 );
and \g135121/U$3 ( \46157 , \41116 , \42643 );
nor \g135121/U$1 ( \46158 , \46156 , \46157 );
and \g134529/U$2 ( \46159 , \46158 , \42487 );
not \g134529/U$4 ( \46160 , \46158 );
and \g134529/U$3 ( \46161 , \46160 , \42486 );
nor \g134529/U$1 ( \46162 , \46159 , \46161 );
xor \g134000/U$4 ( \46163 , \46155 , \46162 );
and \g135125/U$2 ( \46164 , \41087 , \42701 );
and \g135125/U$3 ( \46165 , \42651 , \41328 );
nor \g135125/U$1 ( \46166 , \46164 , \46165 );
and \g134460/U$2 ( \46167 , \46166 , \41093 );
not \g134460/U$4 ( \46168 , \46166 );
and \g134460/U$3 ( \46169 , \46168 , \41092 );
nor \g134460/U$1 ( \46170 , \46167 , \46169 );
and \g134000/U$3 ( \46171 , \46163 , \46170 );
and \g134000/U$5 ( \46172 , \46155 , \46162 );
or \g134000/U$2 ( \46173 , \46171 , \46172 );
and \g135293/U$2 ( \46174 , \43604 , \41144 );
and \g135293/U$3 ( \46175 , \40956 , \43603 );
nor \g135293/U$1 ( \46176 , \46174 , \46175 );
and \g135201/U$2 ( \46177 , \46176 , \42676 );
not \g135201/U$4 ( \46178 , \46176 );
and \g135201/U$3 ( \46179 , \46178 , \42675 );
nor \g135201/U$1 ( \46180 , \46177 , \46179 );
xor \g133988/U$4 ( \46181 , \46180 , \46013 );
and \g134931/U$2 ( \46182 , \43099 , \41107 );
and \g134931/U$3 ( \46183 , \41109 , \43101 );
nor \g134931/U$1 ( \46184 , \46182 , \46183 );
and \g134175/U$2 ( \46185 , \46184 , \42682 );
not \g134175/U$4 ( \46186 , \46184 );
and \g134175/U$3 ( \46187 , \46186 , \42681 );
nor \g134175/U$1 ( \46188 , \46185 , \46187 );
and \g133988/U$3 ( \46189 , \46181 , \46188 );
and \g133988/U$5 ( \46190 , \46180 , \46013 );
or \g133988/U$2 ( \46191 , \46189 , \46190 );
xor \g456215/U$5 ( \46192 , \46173 , \46191 );
and \g134875/U$2 ( \46193 , \41206 , \43179 );
and \g134875/U$3 ( \46194 , \43183 , \41208 );
nor \g134875/U$1 ( \46195 , \46193 , \46194 );
and \g134319/U$2 ( \46196 , \46195 , \41215 );
not \g134319/U$4 ( \46197 , \46195 );
and \g134319/U$3 ( \46198 , \46197 , \41214 );
nor \g134319/U$1 ( \46199 , \46196 , \46198 );
and \g134815/U$2 ( \46200 , \42317 , \41774 );
and \g134815/U$3 ( \46201 , \41629 , \42316 );
nor \g134815/U$1 ( \46202 , \46200 , \46201 );
and \g134535/U$2 ( \46203 , \46202 , \42226 );
not \g134535/U$4 ( \46204 , \46202 );
and \g134535/U$3 ( \46205 , \46204 , \42225 );
nor \g134535/U$1 ( \46206 , \46203 , \46205 );
xor \g456239/U$5 ( \46207 , \46199 , \46206 );
and \g135133/U$2 ( \46208 , \41948 , \42344 );
and \g135133/U$3 ( \46209 , \41920 , \41947 );
nor \g135133/U$1 ( \46210 , \46208 , \46209 );
and \g134431/U$2 ( \46211 , \46210 , \41755 );
not \g134431/U$4 ( \46212 , \46210 );
and \g134431/U$3 ( \46213 , \46212 , \41952 );
nor \g134431/U$1 ( \46214 , \46211 , \46213 );
and \g456239/U$4 ( \46215 , \46207 , \46214 );
and \g456239/U$6 ( \46216 , \46199 , \46206 );
or \g456239/U$3 ( \46217 , \46215 , \46216 );
and \g456215/U$4 ( \46218 , \46192 , \46217 );
and \g456215/U$6 ( \46219 , \46173 , \46191 );
or \g456215/U$3 ( \46220 , \46218 , \46219 );
xor \g456232/U$4 ( \46221 , \46148 , \46220 );
not \g134132/U$3 ( \46222 , \46025 );
not \g134132/U$4 ( \46223 , \46043 );
or \g134132/U$2 ( \46224 , \46222 , \46223 );
or \g134132/U$5 ( \46225 , \46025 , \46043 );
nand \g134132/U$1 ( \46226 , \46224 , \46225 );
not \g134083/U$3 ( \46227 , \46226 );
not \g134083/U$4 ( \46228 , \46032 );
and \g134083/U$2 ( \46229 , \46227 , \46228 );
and \g134083/U$5 ( \46230 , \46226 , \46032 );
nor \g134083/U$1 ( \46231 , \46229 , \46230 );
xor \g456276/U$1 ( \46232 , \46101 , \46107 );
xor \g456276/U$1_r1 ( \46233 , \46232 , \46115 );
or \g133828/U$2 ( \46234 , \46231 , \46233 );
not \g133838/U$3 ( \46235 , \46233 );
not \g133838/U$4 ( \46236 , \46231 );
or \g133838/U$2 ( \46237 , \46235 , \46236 );
xor \g134012/U$1 ( \46238 , \46067 , \46074 );
xor \g134012/U$1_r1 ( \46239 , \46238 , \46082 );
nand \g133838/U$1 ( \46240 , \46237 , \46239 );
nand \g133828/U$1 ( \46241 , \46234 , \46240 );
and \g456232/U$3 ( \46242 , \46221 , \46241 );
and \g456232/U$5 ( \46243 , \46148 , \46220 );
nor \g456232/U$2 ( \46244 , \46242 , \46243 );
xnor \g133665/U$1 ( \46245 , \46050 , \46048 );
not \g133607/U$3 ( \46246 , \46245 );
not \g133607/U$4 ( \46247 , \46056 );
and \g133607/U$2 ( \46248 , \46246 , \46247 );
and \g133607/U$5 ( \46249 , \46245 , \46056 );
nor \g133607/U$1 ( \46250 , \46248 , \46249 );
or \g133440/U$2 ( \46251 , \46244 , \46250 );
not \g133463/U$3 ( \46252 , \46250 );
not \g133463/U$4 ( \46253 , \46244 );
or \g133463/U$2 ( \46254 , \46252 , \46253 );
xor \g133519/U$1 ( \46255 , \46060 , \46095 );
xor \g133519/U$1_r1 ( \46256 , \46255 , \46136 );
nand \g133463/U$1 ( \46257 , \46254 , \46256 );
nand \g133440/U$1 ( \46258 , \46251 , \46257 );
and \g132583/U$2 ( \46259 , \46144 , \46258 );
xor \g133345/U$1 ( \46260 , \46258 , \46144 );
and \g134691/U$2 ( \46261 , \41948 , \42416 );
and \g134691/U$3 ( \46262 , \42344 , \41947 );
nor \g134691/U$1 ( \46263 , \46261 , \46262 );
and \g134500/U$2 ( \46264 , \46263 , \41952 );
not \g134500/U$4 ( \46265 , \46263 );
and \g134500/U$3 ( \46266 , \46265 , \41755 );
nor \g134500/U$1 ( \46267 , \46264 , \46266 );
and \g134994/U$2 ( \46268 , \41623 , \42651 );
and \g134994/U$3 ( \46269 , \42609 , \41745 );
nor \g134994/U$1 ( \46270 , \46268 , \46269 );
and \g134253/U$2 ( \46271 , \46270 , \41324 );
not \g134253/U$4 ( \46272 , \46270 );
and \g134253/U$3 ( \46273 , \46272 , \41325 );
nor \g134253/U$1 ( \46274 , \46271 , \46273 );
or \g134101/U$2 ( \46275 , \46267 , \46274 );
not \g134109/U$3 ( \46276 , \46274 );
not \g134109/U$4 ( \46277 , \46267 );
or \g134109/U$2 ( \46278 , \46276 , \46277 );
and \g134866/U$2 ( \46279 , \42644 , \41629 );
and \g134866/U$3 ( \46280 , \41345 , \42643 );
nor \g134866/U$1 ( \46281 , \46279 , \46280 );
and \g134289/U$2 ( \46282 , \46281 , \42487 );
not \g134289/U$4 ( \46283 , \46281 );
and \g134289/U$3 ( \46284 , \46283 , \42486 );
nor \g134289/U$1 ( \46285 , \46282 , \46284 );
nand \g134109/U$1 ( \46286 , \46278 , \46285 );
nand \g134101/U$1 ( \46287 , \46275 , \46286 );
not \g133864/U$3 ( \46288 , \46287 );
and \g135023/U$2 ( \46289 , \41206 , \43757 );
and \g135023/U$3 ( \46290 , \43179 , \41208 );
nor \g135023/U$1 ( \46291 , \46289 , \46290 );
and \g134513/U$2 ( \46292 , \46291 , \41214 );
not \g134513/U$4 ( \46293 , \46291 );
and \g134513/U$3 ( \46294 , \46293 , \41215 );
nor \g134513/U$1 ( \46295 , \46292 , \46294 );
and \g134954/U$2 ( \46296 , \42317 , \41920 );
and \g134954/U$3 ( \46297 , \41774 , \42316 );
nor \g134954/U$1 ( \46298 , \46296 , \46297 );
and \g134275/U$2 ( \46299 , \46298 , \42225 );
not \g134275/U$4 ( \46300 , \46298 );
and \g134275/U$3 ( \46301 , \46300 , \42226 );
nor \g134275/U$1 ( \46302 , \46299 , \46301 );
xor \g134011/U$4 ( \46303 , \46295 , \46302 );
and \g134812/U$2 ( \46304 , \43099 , \41116 );
and \g134812/U$3 ( \46305 , \41107 , \43101 );
nor \g134812/U$1 ( \46306 , \46304 , \46305 );
and \g134313/U$2 ( \46307 , \46306 , \42681 );
not \g134313/U$4 ( \46308 , \46306 );
and \g134313/U$3 ( \46309 , \46308 , \42682 );
nor \g134313/U$1 ( \46310 , \46307 , \46309 );
and \g134011/U$3 ( \46311 , \46303 , \46310 );
and \g134011/U$5 ( \46312 , \46295 , \46302 );
or \g134011/U$2 ( \46313 , \46311 , \46312 );
not \g133864/U$4 ( \46314 , \46313 );
or \g133864/U$2 ( \46315 , \46288 , \46314 );
or \g133864/U$5 ( \46316 , \46313 , \46287 );
nand \g133864/U$1 ( \46317 , \46315 , \46316 );
not \g133832/U$3 ( \46318 , \46317 );
and \g135317/U$2 ( \46319 , \43604 , \41109 );
and \g135317/U$3 ( \46320 , \41144 , \43603 );
nor \g135317/U$1 ( \46321 , \46319 , \46320 );
and \g135185/U$2 ( \46322 , \46321 , \42675 );
not \g135185/U$4 ( \46323 , \46321 );
and \g135185/U$3 ( \46324 , \46323 , \42676 );
nor \g135185/U$1 ( \46325 , \46322 , \46324 );
not \g134676/U$2 ( \46326 , \46325 );
nor \g135213/U$1 ( \46327 , \41201 , \43607 );
nor \g135164/U$1 ( \46328 , \46327 , \41215 );
nand \g134676/U$1 ( \46329 , \46326 , \46328 );
not \g133832/U$4 ( \46330 , \46329 );
and \g133832/U$2 ( \46331 , \46318 , \46330 );
and \g133832/U$5 ( \46332 , \46317 , \46329 );
nor \g133832/U$1 ( \46333 , \46331 , \46332 );
not \g133616/U$3 ( \46334 , \46333 );
and \g134732/U$2 ( \46335 , \41087 , \43183 );
and \g134732/U$3 ( \46336 , \42701 , \41328 );
nor \g134732/U$1 ( \46337 , \46335 , \46336 );
and \g134353/U$2 ( \46338 , \46337 , \41093 );
not \g134353/U$4 ( \46339 , \46337 );
and \g134353/U$3 ( \46340 , \46339 , \41092 );
nor \g134353/U$1 ( \46341 , \46338 , \46340 );
not \g134658/U$3 ( \46342 , \46328 );
not \g134658/U$4 ( \46343 , \46325 );
or \g134658/U$2 ( \46344 , \46342 , \46343 );
or \g134658/U$5 ( \46345 , \46325 , \46328 );
nand \g134658/U$1 ( \46346 , \46344 , \46345 );
xor \g133771/U$4 ( \46347 , \46341 , \46346 );
and \g135303/U$2 ( \46348 , \43604 , \41107 );
and \g135303/U$3 ( \46349 , \41109 , \43603 );
nor \g135303/U$1 ( \46350 , \46348 , \46349 );
and \g135196/U$2 ( \46351 , \46350 , \42676 );
not \g135196/U$4 ( \46352 , \46350 );
and \g135196/U$3 ( \46353 , \46352 , \42675 );
nor \g135196/U$1 ( \46354 , \46351 , \46353 );
xor \g133954/U$4 ( \46355 , \46354 , \46327 );
and \g134953/U$2 ( \46356 , \43099 , \41345 );
and \g134953/U$3 ( \46357 , \41116 , \43101 );
nor \g134953/U$1 ( \46358 , \46356 , \46357 );
and \g134577/U$2 ( \46359 , \46358 , \42682 );
not \g134577/U$4 ( \46360 , \46358 );
and \g134577/U$3 ( \46361 , \46360 , \42681 );
nor \g134577/U$1 ( \46362 , \46359 , \46361 );
and \g133954/U$3 ( \46363 , \46355 , \46362 );
and \g133954/U$5 ( \46364 , \46354 , \46327 );
or \g133954/U$2 ( \46365 , \46363 , \46364 );
and \g133771/U$3 ( \46366 , \46347 , \46365 );
and \g133771/U$5 ( \46367 , \46341 , \46346 );
or \g133771/U$2 ( \46368 , \46366 , \46367 );
not \g133641/U$3 ( \46369 , \46368 );
not \g134121/U$3 ( \46370 , \46267 );
not \g134121/U$4 ( \46371 , \46285 );
or \g134121/U$2 ( \46372 , \46370 , \46371 );
or \g134121/U$5 ( \46373 , \46267 , \46285 );
nand \g134121/U$1 ( \46374 , \46372 , \46373 );
not \g134079/U$3 ( \46375 , \46374 );
not \g134079/U$4 ( \46376 , \46274 );
and \g134079/U$2 ( \46377 , \46375 , \46376 );
and \g134079/U$5 ( \46378 , \46374 , \46274 );
nor \g134079/U$1 ( \46379 , \46377 , \46378 );
and \g134970/U$2 ( \46380 , \41948 , \42609 );
and \g134970/U$3 ( \46381 , \42416 , \41947 );
nor \g134970/U$1 ( \46382 , \46380 , \46381 );
and \g134454/U$2 ( \46383 , \46382 , \41952 );
not \g134454/U$4 ( \46384 , \46382 );
and \g134454/U$3 ( \46385 , \46384 , \41755 );
nor \g134454/U$1 ( \46386 , \46383 , \46385 );
and \g135061/U$2 ( \46387 , \42644 , \41774 );
and \g135061/U$3 ( \46388 , \41629 , \42643 );
nor \g135061/U$1 ( \46389 , \46387 , \46388 );
and \g134287/U$2 ( \46390 , \46389 , \42486 );
not \g134287/U$4 ( \46391 , \46389 );
and \g134287/U$3 ( \46392 , \46391 , \42487 );
nor \g134287/U$1 ( \46393 , \46390 , \46392 );
xor \g133894/U$4 ( \46394 , \46386 , \46393 );
and \g134738/U$2 ( \46395 , \42317 , \42344 );
and \g134738/U$3 ( \46396 , \41920 , \42316 );
nor \g134738/U$1 ( \46397 , \46395 , \46396 );
and \g134335/U$2 ( \46398 , \46397 , \42225 );
not \g134335/U$4 ( \46399 , \46397 );
and \g134335/U$3 ( \46400 , \46399 , \42226 );
nor \g134335/U$1 ( \46401 , \46398 , \46400 );
and \g133894/U$3 ( \46402 , \46394 , \46401 );
and \g133894/U$5 ( \46403 , \46386 , \46393 );
or \g133894/U$2 ( \46404 , \46402 , \46403 );
xor \g133721/U$4 ( \46405 , \46379 , \46404 );
xor \g134011/U$1 ( \46406 , \46295 , \46302 );
xor \g134011/U$1_r1 ( \46407 , \46406 , \46310 );
and \g133721/U$3 ( \46408 , \46405 , \46407 );
and \g133721/U$5 ( \46409 , \46379 , \46404 );
or \g133721/U$2 ( \46410 , \46408 , \46409 );
not \g133641/U$4 ( \46411 , \46410 );
or \g133641/U$2 ( \46412 , \46369 , \46411 );
or \g133641/U$5 ( \46413 , \46410 , \46368 );
nand \g133641/U$1 ( \46414 , \46412 , \46413 );
not \g133616/U$4 ( \46415 , \46414 );
or \g133616/U$2 ( \46416 , \46334 , \46415 );
or \g133616/U$5 ( \46417 , \46414 , \46333 );
nand \g133616/U$1 ( \46418 , \46416 , \46417 );
not \g133462/U$3 ( \46419 , \46418 );
xor \g456239/U$2 ( \46420 , \46199 , \46206 );
xor \g456239/U$1 ( \46421 , \46420 , \46214 );
xor \g134000/U$1 ( \46422 , \46155 , \46162 );
xor \g134000/U$1_r1 ( \46423 , \46422 , \46170 );
xor \g133988/U$1 ( \46424 , \46180 , \46013 );
xor \g133988/U$1_r1 ( \46425 , \46424 , \46188 );
xor \g456239/U$1_r1 ( \46426 , \46423 , \46425 );
xor \g456239/U$1_r2 ( \46427 , \46421 , \46426 );
and \g135091/U$2 ( \46428 , \41948 , \42651 );
and \g135091/U$3 ( \46429 , \42609 , \41947 );
nor \g135091/U$1 ( \46430 , \46428 , \46429 );
and \g134498/U$2 ( \46431 , \46430 , \41755 );
not \g134498/U$4 ( \46432 , \46430 );
and \g134498/U$3 ( \46433 , \46432 , \41952 );
nor \g134498/U$1 ( \46434 , \46431 , \46433 );
and \g134923/U$2 ( \46435 , \42317 , \42416 );
and \g134923/U$3 ( \46436 , \42344 , \42316 );
nor \g134923/U$1 ( \46437 , \46435 , \46436 );
or \g134159/U$2 ( \46438 , \46437 , \42225 );
nand \g134642/U$1 ( \46439 , \42225 , \46437 );
nand \g134159/U$1 ( \46440 , \46438 , \46439 );
xor \g133946/U$4 ( \46441 , \46434 , \46440 );
and \g134692/U$2 ( \46442 , \43099 , \41629 );
and \g134692/U$3 ( \46443 , \41345 , \43101 );
nor \g134692/U$1 ( \46444 , \46442 , \46443 );
and \g134162/U$2 ( \46445 , \46444 , \42682 );
not \g134162/U$4 ( \46446 , \46444 );
and \g134162/U$3 ( \46447 , \46446 , \42681 );
nor \g134162/U$1 ( \46448 , \46445 , \46447 );
and \g133946/U$3 ( \46449 , \46441 , \46448 );
and \g133946/U$5 ( \46450 , \46434 , \46440 );
or \g133946/U$2 ( \46451 , \46449 , \46450 );
and \g135109/U$2 ( \46452 , \41623 , \43183 );
and \g135109/U$3 ( \46453 , \42701 , \41745 );
nor \g135109/U$1 ( \46454 , \46452 , \46453 );
and \g134615/U$2 ( \46455 , \46454 , \41324 );
not \g134615/U$4 ( \46456 , \46454 );
and \g134615/U$3 ( \46457 , \46456 , \41325 );
nor \g134615/U$1 ( \46458 , \46455 , \46457 );
and \g134935/U$2 ( \46459 , \41087 , \43757 );
and \g134935/U$3 ( \46460 , \43179 , \41328 );
nor \g134935/U$1 ( \46461 , \46459 , \46460 );
and \g134602/U$2 ( \46462 , \46461 , \41092 );
not \g134602/U$4 ( \46463 , \46461 );
and \g134602/U$3 ( \46464 , \46463 , \41093 );
nor \g134602/U$1 ( \46465 , \46462 , \46464 );
or \g134102/U$2 ( \46466 , \46458 , \46465 );
not \g134107/U$3 ( \46467 , \46465 );
not \g134107/U$4 ( \46468 , \46458 );
or \g134107/U$2 ( \46469 , \46467 , \46468 );
and \g134981/U$2 ( \46470 , \42644 , \41920 );
and \g134981/U$3 ( \46471 , \41774 , \42643 );
nor \g134981/U$1 ( \46472 , \46470 , \46471 );
and \g134426/U$2 ( \46473 , \46472 , \42487 );
not \g134426/U$4 ( \46474 , \46472 );
and \g134426/U$3 ( \46475 , \46474 , \42486 );
nor \g134426/U$1 ( \46476 , \46473 , \46475 );
nand \g134107/U$1 ( \46477 , \46469 , \46476 );
nand \g134102/U$1 ( \46478 , \46466 , \46477 );
xor \g133733/U$4 ( \46479 , \46451 , \46478 );
xor \g133954/U$1 ( \46480 , \46354 , \46327 );
xor \g133954/U$1_r1 ( \46481 , \46480 , \46362 );
and \g133733/U$3 ( \46482 , \46479 , \46481 );
and \g133733/U$5 ( \46483 , \46451 , \46478 );
or \g133733/U$2 ( \46484 , \46482 , \46483 );
and \g134683/U$2 ( \46485 , \41623 , \42701 );
and \g134683/U$3 ( \46486 , \42651 , \41745 );
nor \g134683/U$1 ( \46487 , \46485 , \46486 );
and \g134387/U$2 ( \46488 , \46487 , \41324 );
not \g134387/U$4 ( \46489 , \46487 );
and \g134387/U$3 ( \46490 , \46489 , \41325 );
nor \g134387/U$1 ( \46491 , \46488 , \46490 );
and \g135016/U$2 ( \46492 , \41087 , \43179 );
and \g135016/U$3 ( \46493 , \43183 , \41328 );
nor \g135016/U$1 ( \46494 , \46492 , \46493 );
and \g134607/U$2 ( \46495 , \46494 , \41092 );
not \g134607/U$4 ( \46496 , \46494 );
and \g134607/U$3 ( \46497 , \46496 , \41093 );
nor \g134607/U$1 ( \46498 , \46495 , \46497 );
or \g134087/U$2 ( \46499 , \46491 , \46498 );
not \g134103/U$3 ( \46500 , \46498 );
not \g134103/U$4 ( \46501 , \46491 );
or \g134103/U$2 ( \46502 , \46500 , \46501 );
nor \g135220/U$1 ( \46503 , \41080 , \43607 );
nor \g135167/U$1 ( \46504 , \46503 , \41093 );
and \g135300/U$2 ( \46505 , \43604 , \41116 );
and \g135300/U$3 ( \46506 , \41107 , \43603 );
nor \g135300/U$1 ( \46507 , \46505 , \46506 );
and \g135190/U$2 ( \46508 , \46507 , \42676 );
not \g135190/U$4 ( \46509 , \46507 );
and \g135190/U$3 ( \46510 , \46509 , \42675 );
nor \g135190/U$1 ( \46511 , \46508 , \46510 );
and \g134623/U$2 ( \46512 , \46504 , \46511 );
nand \g134103/U$1 ( \46513 , \46502 , \46512 );
nand \g134087/U$1 ( \46514 , \46499 , \46513 );
xor \g133572/U$4 ( \46515 , \46484 , \46514 );
xor \g133771/U$1 ( \46516 , \46341 , \46346 );
xor \g133771/U$1_r1 ( \46517 , \46516 , \46365 );
and \g133572/U$3 ( \46518 , \46515 , \46517 );
and \g133572/U$5 ( \46519 , \46484 , \46514 );
or \g133572/U$2 ( \46520 , \46518 , \46519 );
xnor \g133504/U$1 ( \46521 , \46427 , \46520 );
not \g133462/U$4 ( \46522 , \46521 );
or \g133462/U$2 ( \46523 , \46419 , \46522 );
or \g133462/U$5 ( \46524 , \46521 , \46418 );
nand \g133462/U$1 ( \46525 , \46523 , \46524 );
not \g134129/U$3 ( \46526 , \46512 );
not \g134129/U$4 ( \46527 , \46491 );
or \g134129/U$2 ( \46528 , \46526 , \46527 );
or \g134129/U$5 ( \46529 , \46491 , \46512 );
nand \g134129/U$1 ( \46530 , \46528 , \46529 );
not \g134078/U$3 ( \46531 , \46530 );
not \g134078/U$4 ( \46532 , \46498 );
and \g134078/U$2 ( \46533 , \46531 , \46532 );
and \g134078/U$5 ( \46534 , \46530 , \46498 );
nor \g134078/U$1 ( \46535 , \46533 , \46534 );
not \g133671/U$3 ( \46536 , \46535 );
xor \g133894/U$1 ( \46537 , \46386 , \46393 );
xor \g133894/U$1_r1 ( \46538 , \46537 , \46401 );
not \g133671/U$4 ( \46539 , \46538 );
and \g133671/U$2 ( \46540 , \46536 , \46539 );
and \g133695/U$2 ( \46541 , \46535 , \46538 );
xor \g134623/U$1 ( \46542 , \46504 , \46511 );
not \g133843/U$3 ( \46543 , \46542 );
and \g135005/U$2 ( \46544 , \42317 , \42609 );
and \g135005/U$3 ( \46545 , \42416 , \42316 );
nor \g135005/U$1 ( \46546 , \46544 , \46545 );
and \g134614/U$2 ( \46547 , \46546 , \42226 );
not \g134614/U$4 ( \46548 , \46546 );
and \g134614/U$3 ( \46549 , \46548 , \42225 );
nor \g134614/U$1 ( \46550 , \46547 , \46549 );
xor \g133969/U$4 ( \46551 , \46550 , \46503 );
and \g134801/U$2 ( \46552 , \43099 , \41774 );
and \g134801/U$3 ( \46553 , \41629 , \43101 );
nor \g134801/U$1 ( \46554 , \46552 , \46553 );
and \g134578/U$2 ( \46555 , \46554 , \42682 );
not \g134578/U$4 ( \46556 , \46554 );
and \g134578/U$3 ( \46557 , \46556 , \42681 );
nor \g134578/U$1 ( \46558 , \46555 , \46557 );
and \g133969/U$3 ( \46559 , \46551 , \46558 );
and \g133969/U$5 ( \46560 , \46550 , \46503 );
or \g133969/U$2 ( \46561 , \46559 , \46560 );
not \g133843/U$4 ( \46562 , \46561 );
or \g133843/U$2 ( \46563 , \46543 , \46562 );
or \g133855/U$2 ( \46564 , \46561 , \46542 );
and \g134816/U$2 ( \46565 , \41948 , \42701 );
and \g134816/U$3 ( \46566 , \42651 , \41947 );
nor \g134816/U$1 ( \46567 , \46565 , \46566 );
or \g134160/U$2 ( \46568 , \46567 , \41952 );
nand \g134635/U$1 ( \46569 , \41952 , \46567 );
nand \g134160/U$1 ( \46570 , \46568 , \46569 );
and \g135288/U$2 ( \46571 , \43604 , \41345 );
and \g135288/U$3 ( \46572 , \41116 , \43603 );
nor \g135288/U$1 ( \46573 , \46571 , \46572 );
and \g135204/U$2 ( \46574 , \46573 , \42676 );
not \g135204/U$4 ( \46575 , \46573 );
and \g135204/U$3 ( \46576 , \46575 , \42675 );
nor \g135204/U$1 ( \46577 , \46574 , \46576 );
xor \g133978/U$4 ( \46578 , \46570 , \46577 );
and \g134841/U$2 ( \46579 , \41623 , \43179 );
and \g134841/U$3 ( \46580 , \43183 , \41745 );
nor \g134841/U$1 ( \46581 , \46579 , \46580 );
and \g134569/U$2 ( \46582 , \46581 , \41325 );
not \g134569/U$4 ( \46583 , \46581 );
and \g134569/U$3 ( \46584 , \46583 , \41324 );
nor \g134569/U$1 ( \46585 , \46582 , \46584 );
and \g133978/U$3 ( \46586 , \46578 , \46585 );
and \g133978/U$5 ( \46587 , \46570 , \46577 );
or \g133978/U$2 ( \46588 , \46586 , \46587 );
nand \g133855/U$1 ( \46589 , \46564 , \46588 );
nand \g133843/U$1 ( \46590 , \46563 , \46589 );
not \g133795/U$1 ( \46591 , \46590 );
nor \g133695/U$1 ( \46592 , \46541 , \46591 );
nor \g133671/U$1 ( \46593 , \46540 , \46592 );
xor \g133721/U$1 ( \46594 , \46379 , \46404 );
xor \g133721/U$1_r1 ( \46595 , \46594 , \46407 );
or \g133469/U$2 ( \46596 , \46593 , \46595 );
not \g133482/U$3 ( \46597 , \46595 );
not \g133482/U$4 ( \46598 , \46593 );
or \g133482/U$2 ( \46599 , \46597 , \46598 );
xor \g133572/U$1 ( \46600 , \46484 , \46514 );
xor \g133572/U$1_r1 ( \46601 , \46600 , \46517 );
nand \g133482/U$1 ( \46602 , \46599 , \46601 );
nand \g133469/U$1 ( \46603 , \46596 , \46602 );
and \g132868/U$2 ( \46604 , \46525 , \46603 );
xor \g133377/U$1 ( \46605 , \46603 , \46525 );
not \g133470/U$3 ( \46606 , \46601 );
xnor \g133528/U$1 ( \46607 , \46595 , \46593 );
not \g133470/U$4 ( \46608 , \46607 );
and \g133470/U$2 ( \46609 , \46606 , \46608 );
and \g133470/U$5 ( \46610 , \46601 , \46607 );
nor \g133470/U$1 ( \46611 , \46609 , \46610 );
not \g133626/U$3 ( \46612 , \46535 );
not \g133667/U$3 ( \46613 , \46538 );
not \g133667/U$4 ( \46614 , \46590 );
or \g133667/U$2 ( \46615 , \46613 , \46614 );
or \g133667/U$5 ( \46616 , \46590 , \46538 );
nand \g133667/U$1 ( \46617 , \46615 , \46616 );
not \g133626/U$4 ( \46618 , \46617 );
or \g133626/U$2 ( \46619 , \46612 , \46618 );
or \g133626/U$5 ( \46620 , \46617 , \46535 );
nand \g133626/U$1 ( \46621 , \46619 , \46620 );
and \g134941/U$2 ( \46622 , \41948 , \43183 );
and \g134941/U$3 ( \46623 , \42701 , \41947 );
nor \g134941/U$1 ( \46624 , \46622 , \46623 );
and \g134379/U$2 ( \46625 , \46624 , \41952 );
not \g134379/U$4 ( \46626 , \46624 );
and \g134379/U$3 ( \46627 , \46626 , \41755 );
nor \g134379/U$1 ( \46628 , \46625 , \46627 );
and \g135305/U$2 ( \46629 , \43604 , \41629 );
and \g135305/U$3 ( \46630 , \41345 , \43603 );
nor \g135305/U$1 ( \46631 , \46629 , \46630 );
and \g135176/U$2 ( \46632 , \46631 , \42675 );
not \g135176/U$4 ( \46633 , \46631 );
and \g135176/U$3 ( \46634 , \46633 , \42676 );
nor \g135176/U$1 ( \46635 , \46632 , \46634 );
xor \g133905/U$4 ( \46636 , \46628 , \46635 );
and \g134920/U$2 ( \46637 , \42317 , \42651 );
and \g134920/U$3 ( \46638 , \42609 , \42316 );
nor \g134920/U$1 ( \46639 , \46637 , \46638 );
and \g134425/U$2 ( \46640 , \46639 , \42225 );
not \g134425/U$4 ( \46641 , \46639 );
and \g134425/U$3 ( \46642 , \46641 , \42226 );
nor \g134425/U$1 ( \46643 , \46640 , \46642 );
and \g133905/U$3 ( \46644 , \46636 , \46643 );
and \g133905/U$5 ( \46645 , \46628 , \46635 );
or \g133905/U$2 ( \46646 , \46644 , \46645 );
not \g133827/U$3 ( \46647 , \46646 );
and \g134988/U$2 ( \46648 , \42644 , \42344 );
and \g134988/U$3 ( \46649 , \41920 , \42643 );
nor \g134988/U$1 ( \46650 , \46648 , \46649 );
and \g134381/U$2 ( \46651 , \46650 , \42486 );
not \g134381/U$4 ( \46652 , \46650 );
and \g134381/U$3 ( \46653 , \46652 , \42487 );
nor \g134381/U$1 ( \46654 , \46651 , \46653 );
not \g133827/U$4 ( \46655 , \46654 );
and \g133827/U$2 ( \46656 , \46647 , \46655 );
and \g133837/U$2 ( \46657 , \46646 , \46654 );
and \g134813/U$2 ( \46658 , \43099 , \41920 );
and \g134813/U$3 ( \46659 , \41774 , \43101 );
nor \g134813/U$1 ( \46660 , \46658 , \46659 );
and \g134202/U$2 ( \46661 , \46660 , \42681 );
not \g134202/U$4 ( \46662 , \46660 );
and \g134202/U$3 ( \46663 , \46662 , \42682 );
nor \g134202/U$1 ( \46664 , \46661 , \46663 );
not \g134142/U$2 ( \46665 , \46664 );
nor \g135215/U$1 ( \46666 , \41617 , \43607 );
nor \g135163/U$1 ( \46667 , \46666 , \41325 );
nand \g134142/U$1 ( \46668 , \46665 , \46667 );
nor \g133837/U$1 ( \46669 , \46657 , \46668 );
nor \g133827/U$1 ( \46670 , \46656 , \46669 );
not \g134133/U$3 ( \46671 , \46458 );
not \g134133/U$4 ( \46672 , \46476 );
or \g134133/U$2 ( \46673 , \46671 , \46672 );
or \g134133/U$5 ( \46674 , \46458 , \46476 );
nand \g134133/U$1 ( \46675 , \46673 , \46674 );
not \g134076/U$3 ( \46676 , \46675 );
not \g134076/U$4 ( \46677 , \46465 );
and \g134076/U$2 ( \46678 , \46676 , \46677 );
and \g134076/U$5 ( \46679 , \46675 , \46465 );
nor \g134076/U$1 ( \46680 , \46678 , \46679 );
not \g133883/U$2 ( \46681 , \46680 );
xor \g133946/U$1 ( \46682 , \46434 , \46440 );
xor \g133946/U$1_r1 ( \46683 , \46682 , \46448 );
nor \g133883/U$1 ( \46684 , \46681 , \46683 );
or \g133653/U$2 ( \46685 , \46670 , \46684 );
not \g133881/U$2 ( \46686 , \46680 );
nand \g133881/U$1 ( \46687 , \46686 , \46683 );
nand \g133653/U$1 ( \46688 , \46685 , \46687 );
xor \g133733/U$1 ( \46689 , \46451 , \46478 );
xor \g133733/U$1_r1 ( \46690 , \46689 , \46481 );
or \g133523/U$1 ( \46691 , \46688 , \46690 );
and \g133447/U$2 ( \46692 , \46621 , \46691 );
and \g133447/U$3 ( \46693 , \46690 , \46688 );
nor \g133447/U$1 ( \46694 , \46692 , \46693 );
or \g132921/U$2 ( \46695 , \46611 , \46694 );
xnor \g133374/U$1 ( \46696 , \46694 , \46611 );
not \g133452/U$3 ( \46697 , \46621 );
xnor \g133500/U$1 ( \46698 , \46690 , \46688 );
not \g133452/U$4 ( \46699 , \46698 );
or \g133452/U$2 ( \46700 , \46697 , \46699 );
or \g133452/U$5 ( \46701 , \46698 , \46621 );
nand \g133452/U$1 ( \46702 , \46700 , \46701 );
xor \g133969/U$1 ( \46703 , \46550 , \46503 );
xor \g133969/U$1_r1 ( \46704 , \46703 , \46558 );
xor \g133978/U$1 ( \46705 , \46570 , \46577 );
xor \g133978/U$1_r1 ( \46706 , \46705 , \46585 );
and \g133763/U$2 ( \46707 , \46704 , \46706 );
not \g133818/U$3 ( \46708 , \46704 );
not \g133818/U$4 ( \46709 , \46706 );
and \g133818/U$2 ( \46710 , \46708 , \46709 );
and \g135079/U$2 ( \46711 , \41623 , \43757 );
and \g135079/U$3 ( \46712 , \43179 , \41745 );
nor \g135079/U$1 ( \46713 , \46711 , \46712 );
and \g134351/U$2 ( \46714 , \46713 , \41324 );
not \g134351/U$4 ( \46715 , \46713 );
and \g134351/U$3 ( \46716 , \46715 , \41325 );
nor \g134351/U$1 ( \46717 , \46714 , \46716 );
and \g135071/U$2 ( \46718 , \42644 , \42416 );
and \g135071/U$3 ( \46719 , \42344 , \42643 );
nor \g135071/U$1 ( \46720 , \46718 , \46719 );
and \g134562/U$2 ( \46721 , \46720 , \42486 );
not \g134562/U$4 ( \46722 , \46720 );
and \g134562/U$3 ( \46723 , \46722 , \42487 );
nor \g134562/U$1 ( \46724 , \46721 , \46723 );
xor \g133849/U$4 ( \46725 , \46717 , \46724 );
not \g134113/U$3 ( \46726 , \46664 );
not \g134113/U$4 ( \46727 , \46667 );
and \g134113/U$2 ( \46728 , \46726 , \46727 );
and \g134113/U$5 ( \46729 , \46664 , \46667 );
nor \g134113/U$1 ( \46730 , \46728 , \46729 );
and \g133849/U$3 ( \46731 , \46725 , \46730 );
and \g133849/U$5 ( \46732 , \46717 , \46724 );
or \g133849/U$2 ( \46733 , \46731 , \46732 );
nor \g133818/U$1 ( \46734 , \46710 , \46733 );
nor \g133763/U$1 ( \46735 , \46707 , \46734 );
xnor \g133862/U$1 ( \46736 , \46542 , \46588 );
not \g133833/U$3 ( \46737 , \46736 );
not \g133833/U$4 ( \46738 , \46561 );
and \g133833/U$2 ( \46739 , \46737 , \46738 );
and \g133833/U$5 ( \46740 , \46736 , \46561 );
nor \g133833/U$1 ( \46741 , \46739 , \46740 );
or \g133508/U$2 ( \46742 , \46735 , \46741 );
and \g133526/U$2 ( \46743 , \46735 , \46741 );
not \g133637/U$3 ( \46744 , \46683 );
not \g133637/U$4 ( \46745 , \46670 );
or \g133637/U$2 ( \46746 , \46744 , \46745 );
or \g133637/U$5 ( \46747 , \46670 , \46683 );
nand \g133637/U$1 ( \46748 , \46746 , \46747 );
not \g133613/U$3 ( \46749 , \46748 );
not \g133613/U$4 ( \46750 , \46680 );
and \g133613/U$2 ( \46751 , \46749 , \46750 );
and \g133613/U$5 ( \46752 , \46748 , \46680 );
nor \g133613/U$1 ( \46753 , \46751 , \46752 );
nor \g133526/U$1 ( \46754 , \46743 , \46753 );
not \g133525/U$1 ( \46755 , \46754 );
nand \g133508/U$1 ( \46756 , \46742 , \46755 );
and \g132973/U$2 ( \46757 , \46702 , \46756 );
xor \g133375/U$1 ( \46758 , \46756 , \46702 );
and \g135022/U$2 ( \46759 , \42644 , \42609 );
and \g135022/U$3 ( \46760 , \42416 , \42643 );
nor \g135022/U$1 ( \46761 , \46759 , \46760 );
and \g134333/U$2 ( \46762 , \46761 , \42487 );
not \g134333/U$4 ( \46763 , \46761 );
and \g134333/U$3 ( \46764 , \46763 , \42486 );
nor \g134333/U$1 ( \46765 , \46762 , \46764 );
and \g135291/U$2 ( \46766 , \43604 , \41774 );
and \g135291/U$3 ( \46767 , \41629 , \43603 );
nor \g135291/U$1 ( \46768 , \46766 , \46767 );
and \g135198/U$2 ( \46769 , \46768 , \42676 );
not \g135198/U$4 ( \46770 , \46768 );
and \g135198/U$3 ( \46771 , \46770 , \42675 );
nor \g135198/U$1 ( \46772 , \46769 , \46771 );
xor \g456273/U$4 ( \46773 , \46765 , \46772 );
and \g135051/U$2 ( \46774 , \41948 , \43179 );
and \g135051/U$3 ( \46775 , \43183 , \41947 );
nor \g135051/U$1 ( \46776 , \46774 , \46775 );
and \g134449/U$2 ( \46777 , \46776 , \41755 );
not \g134449/U$4 ( \46778 , \46776 );
and \g134449/U$3 ( \46779 , \46778 , \41952 );
nor \g134449/U$1 ( \46780 , \46777 , \46779 );
and \g456273/U$3 ( \46781 , \46773 , \46780 );
and \g456273/U$5 ( \46782 , \46765 , \46772 );
nor \g456273/U$2 ( \46783 , \46781 , \46782 );
and \g134858/U$2 ( \46784 , \42317 , \42701 );
and \g134858/U$3 ( \46785 , \42651 , \42316 );
nor \g134858/U$1 ( \46786 , \46784 , \46785 );
and \g134601/U$2 ( \46787 , \46786 , \42226 );
not \g134601/U$4 ( \46788 , \46786 );
and \g134601/U$3 ( \46789 , \46788 , \42225 );
nor \g134601/U$1 ( \46790 , \46787 , \46789 );
xor \g456277/U$4 ( \46791 , \46666 , \46790 );
and \g135086/U$2 ( \46792 , \43099 , \42344 );
and \g135086/U$3 ( \46793 , \41920 , \43101 );
nor \g135086/U$1 ( \46794 , \46792 , \46793 );
and \g134200/U$2 ( \46795 , \46794 , \42682 );
not \g134200/U$4 ( \46796 , \46794 );
and \g134200/U$3 ( \46797 , \46796 , \42681 );
nor \g134200/U$1 ( \46798 , \46795 , \46797 );
and \g456277/U$3 ( \46799 , \46791 , \46798 );
and \g456277/U$5 ( \46800 , \46666 , \46790 );
nor \g456277/U$2 ( \46801 , \46799 , \46800 );
xor \g456259/U$4 ( \46802 , \46783 , \46801 );
xor \g133905/U$1 ( \46803 , \46628 , \46635 );
xor \g133905/U$1_r1 ( \46804 , \46803 , \46643 );
and \g456259/U$3 ( \46805 , \46802 , \46804 );
and \g456259/U$5 ( \46806 , \46783 , \46801 );
nor \g456259/U$2 ( \46807 , \46805 , \46806 );
not \g133810/U$3 ( \46808 , \46654 );
xor \g133841/U$1 ( \46809 , \46668 , \46646 );
not \g133810/U$4 ( \46810 , \46809 );
or \g133810/U$2 ( \46811 , \46808 , \46810 );
or \g133810/U$5 ( \46812 , \46809 , \46654 );
nand \g133810/U$1 ( \46813 , \46811 , \46812 );
xor \g456211/U$1 ( \46814 , \46807 , \46813 );
not \g133691/U$3 ( \46815 , \46704 );
not \g133760/U$3 ( \46816 , \46733 );
not \g133760/U$4 ( \46817 , \46706 );
and \g133760/U$2 ( \46818 , \46816 , \46817 );
and \g133760/U$5 ( \46819 , \46733 , \46706 );
nor \g133760/U$1 ( \46820 , \46818 , \46819 );
not \g133691/U$4 ( \46821 , \46820 );
or \g133691/U$2 ( \46822 , \46815 , \46821 );
or \g133691/U$5 ( \46823 , \46820 , \46704 );
nand \g133691/U$1 ( \46824 , \46822 , \46823 );
xor \g456211/U$1_r1 ( \46825 , \46814 , \46824 );
xor \g456259/U$1 ( \46826 , \46783 , \46801 );
xor \g456259/U$1_r1 ( \46827 , \46826 , \46804 );
xor \g133849/U$1 ( \46828 , \46717 , \46724 );
xor \g133849/U$1_r1 ( \46829 , \46828 , \46730 );
or \g133604/U$2 ( \46830 , \46827 , \46829 );
not \g133617/U$3 ( \46831 , \46829 );
not \g133617/U$4 ( \46832 , \46827 );
or \g133617/U$2 ( \46833 , \46831 , \46832 );
and \g134881/U$2 ( \46834 , \41948 , \43757 );
and \g134881/U$3 ( \46835 , \43179 , \41947 );
nor \g134881/U$1 ( \46836 , \46834 , \46835 );
and \g134338/U$2 ( \46837 , \46836 , \41952 );
not \g134338/U$4 ( \46838 , \46836 );
and \g134338/U$3 ( \46839 , \46838 , \41755 );
nor \g134338/U$1 ( \46840 , \46837 , \46839 );
and \g135314/U$2 ( \46841 , \43604 , \41920 );
and \g135314/U$3 ( \46842 , \41774 , \43603 );
nor \g135314/U$1 ( \46843 , \46841 , \46842 );
and \g135195/U$2 ( \46844 , \46843 , \42675 );
not \g135195/U$4 ( \46845 , \46843 );
and \g135195/U$3 ( \46846 , \46845 , \42676 );
nor \g135195/U$1 ( \46847 , \46844 , \46846 );
or \g134094/U$2 ( \46848 , \46840 , \46847 );
not \g134105/U$3 ( \46849 , \46847 );
not \g134105/U$4 ( \46850 , \46840 );
or \g134105/U$2 ( \46851 , \46849 , \46850 );
and \g134729/U$2 ( \46852 , \42317 , \43183 );
and \g134729/U$3 ( \46853 , \42701 , \42316 );
nor \g134729/U$1 ( \46854 , \46852 , \46853 );
and \g134218/U$2 ( \46855 , \46854 , \42226 );
not \g134218/U$4 ( \46856 , \46854 );
and \g134218/U$3 ( \46857 , \46856 , \42225 );
nor \g134218/U$1 ( \46858 , \46855 , \46857 );
nand \g134105/U$1 ( \46859 , \46851 , \46858 );
nand \g134094/U$1 ( \46860 , \46848 , \46859 );
nand \g135222/U$1 ( \46861 , \43757 , \41947 );
not \g135221/U$1 ( \46862 , \46861 );
nor \g135166/U$1 ( \46863 , \46862 , \41755 );
and \g134882/U$2 ( \46864 , \43099 , \42416 );
and \g134882/U$3 ( \46865 , \42344 , \43101 );
nor \g134882/U$1 ( \46866 , \46864 , \46865 );
and \g134526/U$2 ( \46867 , \46866 , \42682 );
not \g134526/U$4 ( \46868 , \46866 );
and \g134526/U$3 ( \46869 , \46868 , \42681 );
nor \g134526/U$1 ( \46870 , \46867 , \46869 );
and \g134088/U$2 ( \46871 , \46863 , \46870 );
xor \g133807/U$4 ( \46872 , \46860 , \46871 );
xor \g456277/U$1 ( \46873 , \46666 , \46790 );
xor \g456277/U$1_r1 ( \46874 , \46873 , \46798 );
and \g133807/U$3 ( \46875 , \46872 , \46874 );
and \g133807/U$5 ( \46876 , \46860 , \46871 );
or \g133807/U$2 ( \46877 , \46875 , \46876 );
nand \g133617/U$1 ( \46878 , \46833 , \46877 );
nand \g133604/U$1 ( \46879 , \46830 , \46878 );
and \g133082/U$2 ( \46880 , \46825 , \46879 );
xor \g133466/U$1 ( \46881 , \46879 , \46825 );
and \g135318/U$2 ( \46882 , \43604 , \42344 );
and \g135318/U$3 ( \46883 , \41920 , \43603 );
nor \g135318/U$1 ( \46884 , \46882 , \46883 );
and \g135178/U$2 ( \46885 , \46884 , \42675 );
not \g135178/U$4 ( \46886 , \46884 );
and \g135178/U$3 ( \46887 , \46886 , \42676 );
nor \g135178/U$1 ( \46888 , \46885 , \46887 );
or \g134135/U$2 ( \46889 , \46888 , \46861 );
not \g134146/U$3 ( \46890 , \46861 );
not \g134146/U$4 ( \46891 , \46888 );
or \g134146/U$2 ( \46892 , \46890 , \46891 );
and \g134948/U$2 ( \46893 , \42317 , \43179 );
and \g134948/U$3 ( \46894 , \43183 , \42316 );
nor \g134948/U$1 ( \46895 , \46893 , \46894 );
and \g134497/U$2 ( \46896 , \46895 , \42226 );
not \g134497/U$4 ( \46897 , \46895 );
and \g134497/U$3 ( \46898 , \46897 , \42225 );
nor \g134497/U$1 ( \46899 , \46896 , \46898 );
nand \g134146/U$1 ( \46900 , \46892 , \46899 );
nand \g134135/U$1 ( \46901 , \46889 , \46900 );
and \g134809/U$2 ( \46902 , \42644 , \42651 );
and \g134809/U$3 ( \46903 , \42609 , \42643 );
nor \g134809/U$1 ( \46904 , \46902 , \46903 );
and \g134606/U$2 ( \46905 , \46904 , \42487 );
not \g134606/U$4 ( \46906 , \46904 );
and \g134606/U$3 ( \46907 , \46906 , \42486 );
nor \g134606/U$1 ( \46908 , \46905 , \46907 );
xor \g133805/U$4 ( \46909 , \46901 , \46908 );
xor \g134088/U$1 ( \46910 , \46863 , \46870 );
and \g133805/U$3 ( \46911 , \46909 , \46910 );
and \g133805/U$5 ( \46912 , \46901 , \46908 );
or \g133805/U$2 ( \46913 , \46911 , \46912 );
xor \g456273/U$1 ( \46914 , \46765 , \46772 );
xor \g456273/U$1_r1 ( \46915 , \46914 , \46780 );
xor \g456230/U$1 ( \46916 , \46913 , \46915 );
xor \g133807/U$1 ( \46917 , \46860 , \46871 );
xor \g133807/U$1_r1 ( \46918 , \46917 , \46874 );
xor \g456230/U$1_r1 ( \46919 , \46916 , \46918 );
and \g134784/U$2 ( \46920 , \42644 , \42701 );
and \g134784/U$3 ( \46921 , \42651 , \42643 );
nor \g134784/U$1 ( \46922 , \46920 , \46921 );
and \g134223/U$2 ( \46923 , \46922 , \42486 );
not \g134223/U$4 ( \46924 , \46922 );
and \g134223/U$3 ( \46925 , \46924 , \42487 );
nor \g134223/U$1 ( \46926 , \46923 , \46925 );
and \g135295/U$2 ( \46927 , \43604 , \42416 );
and \g135295/U$3 ( \46928 , \42344 , \43603 );
nor \g135295/U$1 ( \46929 , \46927 , \46928 );
and \g135183/U$2 ( \46930 , \46929 , \42675 );
not \g135183/U$4 ( \46931 , \46929 );
and \g135183/U$3 ( \46932 , \46931 , \42676 );
nor \g135183/U$1 ( \46933 , \46930 , \46932 );
not \g134677/U$2 ( \46934 , \46933 );
nand \g135218/U$1 ( \46935 , \43757 , \42316 );
not \g135217/U$1 ( \46936 , \46935 );
nor \g135162/U$1 ( \46937 , \46936 , \42226 );
nand \g134677/U$1 ( \46938 , \46934 , \46937 );
xor \g134051/U$4 ( \46939 , \46926 , \46938 );
and \g134737/U$2 ( \46940 , \43099 , \42609 );
and \g134737/U$3 ( \46941 , \42416 , \43101 );
nor \g134737/U$1 ( \46942 , \46940 , \46941 );
and \g134245/U$2 ( \46943 , \46942 , \42681 );
not \g134245/U$4 ( \46944 , \46942 );
and \g134245/U$3 ( \46945 , \46944 , \42682 );
nor \g134245/U$1 ( \46946 , \46943 , \46945 );
and \g134051/U$3 ( \46947 , \46939 , \46946 );
and \g134051/U$5 ( \46948 , \46926 , \46938 );
or \g134051/U$2 ( \46949 , \46947 , \46948 );
not \g134130/U$3 ( \46950 , \46847 );
not \g134130/U$4 ( \46951 , \46858 );
or \g134130/U$2 ( \46952 , \46950 , \46951 );
or \g134130/U$5 ( \46953 , \46858 , \46847 );
nand \g134130/U$1 ( \46954 , \46952 , \46953 );
not \g134074/U$3 ( \46955 , \46954 );
not \g134074/U$4 ( \46956 , \46840 );
and \g134074/U$2 ( \46957 , \46955 , \46956 );
and \g134074/U$5 ( \46958 , \46954 , \46840 );
nor \g134074/U$1 ( \46959 , \46957 , \46958 );
or \g133673/U$2 ( \46960 , \46949 , \46959 );
not \g133694/U$3 ( \46961 , \46959 );
not \g133694/U$4 ( \46962 , \46949 );
or \g133694/U$2 ( \46963 , \46961 , \46962 );
xor \g133805/U$1 ( \46964 , \46901 , \46908 );
xor \g133805/U$1_r1 ( \46965 , \46964 , \46910 );
nand \g133694/U$1 ( \46966 , \46963 , \46965 );
nand \g133673/U$1 ( \46967 , \46960 , \46966 );
and \g133179/U$2 ( \46968 , \46919 , \46967 );
xor \g133502/U$1 ( \46969 , \46967 , \46919 );
nor \g135206/U$1 ( \46970 , \43093 , \43607 );
nor \g135158/U$1 ( \46971 , \46970 , \42682 );
not \g134674/U$2 ( \46972 , \46971 );
and \g135308/U$2 ( \46973 , \43604 , \43183 );
and \g135308/U$3 ( \46974 , \42701 , \43603 );
nor \g135308/U$1 ( \46975 , \46973 , \46974 );
and \g135180/U$2 ( \46976 , \46975 , \42675 );
not \g135180/U$4 ( \46977 , \46975 );
and \g135180/U$3 ( \46978 , \46977 , \42676 );
nor \g135180/U$1 ( \46979 , \46976 , \46978 );
nor \g134674/U$1 ( \46980 , \46972 , \46979 );
nand \g135212/U$1 ( \46981 , \43757 , \42643 );
not \g135211/U$1 ( \46982 , \46981 );
not \g134070/U$3 ( \46983 , \46982 );
and \g134802/U$2 ( \46984 , \43099 , \43179 );
and \g134802/U$3 ( \46985 , \43183 , \43101 );
nor \g134802/U$1 ( \46986 , \46984 , \46985 );
and \g134393/U$2 ( \46987 , \46986 , \42681 );
not \g134393/U$4 ( \46988 , \46986 );
and \g134393/U$3 ( \46989 , \46988 , \42682 );
nor \g134393/U$1 ( \46990 , \46987 , \46989 );
and \g135306/U$2 ( \46991 , \43604 , \42701 );
and \g135306/U$3 ( \46992 , \42651 , \43603 );
nor \g135306/U$1 ( \46993 , \46991 , \46992 );
and \g135199/U$2 ( \46994 , \46993 , \42675 );
not \g135199/U$4 ( \46995 , \46993 );
and \g135199/U$3 ( \46996 , \46995 , \42676 );
nor \g135199/U$1 ( \46997 , \46994 , \46996 );
xnor \g455962/U$1 ( \46998 , \46990 , \46997 );
not \g134070/U$4 ( \46999 , \46998 );
or \g134070/U$2 ( \47000 , \46983 , \46999 );
or \g134070/U$5 ( \47001 , \46998 , \46982 );
nand \g134070/U$1 ( \47002 , \47000 , \47001 );
xor \g133866/U$1 ( \47003 , \46980 , \47002 );
not \g134664/U$3 ( \47004 , \46971 );
not \g134664/U$4 ( \47005 , \46979 );
and \g134664/U$2 ( \47006 , \47004 , \47005 );
and \g134664/U$5 ( \47007 , \46971 , \46979 );
nor \g134664/U$1 ( \47008 , \47006 , \47007 );
and \g134698/U$2 ( \47009 , \43099 , \43757 );
and \g134698/U$3 ( \47010 , \43179 , \43101 );
nor \g134698/U$1 ( \47011 , \47009 , \47010 );
and \g134192/U$2 ( \47012 , \47011 , \42681 );
not \g134192/U$4 ( \47013 , \47011 );
and \g134192/U$3 ( \47014 , \47013 , \42682 );
nor \g134192/U$1 ( \47015 , \47012 , \47014 );
xnor \g134124/U$1 ( \47016 , \47008 , \47015 );
and \g135296/U$2 ( \47017 , \43604 , \43179 );
and \g135296/U$3 ( \47018 , \43183 , \43603 );
nor \g135296/U$1 ( \47019 , \47017 , \47018 );
and \g135197/U$2 ( \47020 , \47019 , \42676 );
not \g135197/U$4 ( \47021 , \47019 );
and \g135197/U$3 ( \47022 , \47021 , \42675 );
nor \g135197/U$1 ( \47023 , \47020 , \47022 );
xor \g134672/U$1 ( \47024 , \46970 , \47023 );
nand \g135367/U$1 ( \47025 , \43757 , \43603 );
not \g135366/U$1 ( \47026 , \47025 );
nor \g135319/U$1 ( \47027 , \47026 , \42676 );
and \g135294/U$2 ( \47028 , \43604 , \43757 );
and \g135294/U$3 ( \47029 , \43179 , \43603 );
nor \g135294/U$1 ( \47030 , \47028 , \47029 );
and \g135194/U$2 ( \47031 , \47030 , \42676 );
not \g135194/U$4 ( \47032 , \47030 );
and \g135194/U$3 ( \47033 , \47032 , \42675 );
nor \g135194/U$1 ( \47034 , \47031 , \47033 );
and \g134629/U$2 ( \47035 , \47027 , \47034 );
and \g134069/U$2 ( \47036 , \47024 , \47035 );
and \g134069/U$3 ( \47037 , \46970 , \47023 );
nor \g134069/U$1 ( \47038 , \47036 , \47037 );
or \g133844/U$2 ( \47039 , \47016 , \47038 );
or \g133844/U$3 ( \47040 , \47008 , \47015 );
nand \g133844/U$1 ( \47041 , \47039 , \47040 );
and \g133672/U$2 ( \47042 , \47003 , \47041 );
and \g133672/U$3 ( \47043 , \46980 , \47002 );
nor \g133672/U$1 ( \47044 , \47042 , \47043 );
not \g134136/U$3 ( \47045 , \46997 );
not \g134136/U$4 ( \47046 , \46981 );
and \g134136/U$2 ( \47047 , \47045 , \47046 );
and \g134147/U$2 ( \47048 , \46997 , \46981 );
nor \g134147/U$1 ( \47049 , \47048 , \46990 );
nor \g134136/U$1 ( \47050 , \47047 , \47049 );
nor \g135161/U$1 ( \47051 , \46982 , \42487 );
and \g135311/U$2 ( \47052 , \43604 , \42651 );
and \g135311/U$3 ( \47053 , \42609 , \43603 );
nor \g135311/U$1 ( \47054 , \47052 , \47053 );
and \g135193/U$2 ( \47055 , \47054 , \42676 );
not \g135193/U$4 ( \47056 , \47054 );
and \g135193/U$3 ( \47057 , \47056 , \42675 );
nor \g135193/U$1 ( \47058 , \47055 , \47057 );
xor \g134627/U$1 ( \47059 , \47051 , \47058 );
not \g134116/U$3 ( \47060 , \47059 );
and \g134835/U$2 ( \47061 , \43099 , \43183 );
and \g134835/U$3 ( \47062 , \42701 , \43101 );
nor \g134835/U$1 ( \47063 , \47061 , \47062 );
and \g134203/U$2 ( \47064 , \47063 , \42681 );
not \g134203/U$4 ( \47065 , \47063 );
and \g134203/U$3 ( \47066 , \47065 , \42682 );
nor \g134203/U$1 ( \47067 , \47064 , \47066 );
not \g134116/U$4 ( \47068 , \47067 );
or \g134116/U$2 ( \47069 , \47060 , \47068 );
or \g134116/U$5 ( \47070 , \47067 , \47059 );
nand \g134116/U$1 ( \47071 , \47069 , \47070 );
not \g134077/U$3 ( \47072 , \47071 );
and \g134947/U$2 ( \47073 , \42644 , \43757 );
and \g134947/U$3 ( \47074 , \43179 , \42643 );
nor \g134947/U$1 ( \47075 , \47073 , \47074 );
and \g134197/U$2 ( \47076 , \47075 , \42486 );
not \g134197/U$4 ( \47077 , \47075 );
and \g134197/U$3 ( \47078 , \47077 , \42487 );
nor \g134197/U$1 ( \47079 , \47076 , \47078 );
not \g134077/U$4 ( \47080 , \47079 );
and \g134077/U$2 ( \47081 , \47072 , \47080 );
and \g134077/U$5 ( \47082 , \47071 , \47079 );
nor \g134077/U$1 ( \47083 , \47081 , \47082 );
xnor \g133869/U$1 ( \47084 , \47050 , \47083 );
or \g133559/U$2 ( \47085 , \47044 , \47084 );
or \g133559/U$3 ( \47086 , \47050 , \47083 );
nand \g133559/U$1 ( \47087 , \47085 , \47086 );
or \g134097/U$2 ( \47088 , \47067 , \47079 );
not \g134112/U$3 ( \47089 , \47079 );
not \g134112/U$4 ( \47090 , \47067 );
or \g134112/U$2 ( \47091 , \47089 , \47090 );
nand \g134112/U$1 ( \47092 , \47091 , \47059 );
nand \g134097/U$1 ( \47093 , \47088 , \47092 );
and \g134627/U$2 ( \47094 , \47051 , \47058 );
and \g134901/U$2 ( \47095 , \42644 , \43179 );
and \g134901/U$3 ( \47096 , \43183 , \42643 );
nor \g134901/U$1 ( \47097 , \47095 , \47096 );
and \g134611/U$2 ( \47098 , \47097 , \42487 );
not \g134611/U$4 ( \47099 , \47097 );
and \g134611/U$3 ( \47100 , \47099 , \42486 );
nor \g134611/U$1 ( \47101 , \47098 , \47100 );
xor \g456272/U$1 ( \47102 , \47094 , \47101 );
not \g134071/U$3 ( \47103 , \46936 );
and \g135014/U$2 ( \47104 , \43099 , \42701 );
and \g135014/U$3 ( \47105 , \42651 , \43101 );
nor \g135014/U$1 ( \47106 , \47104 , \47105 );
and \g134442/U$2 ( \47107 , \47106 , \42681 );
not \g134442/U$4 ( \47108 , \47106 );
and \g134442/U$3 ( \47109 , \47108 , \42682 );
nor \g134442/U$1 ( \47110 , \47107 , \47109 );
and \g135307/U$2 ( \47111 , \43604 , \42609 );
and \g135307/U$3 ( \47112 , \42416 , \43603 );
nor \g135307/U$1 ( \47113 , \47111 , \47112 );
and \g135187/U$2 ( \47114 , \47113 , \42675 );
not \g135187/U$4 ( \47115 , \47113 );
and \g135187/U$3 ( \47116 , \47115 , \42676 );
nor \g135187/U$1 ( \47117 , \47114 , \47116 );
xnor \g455961/U$1 ( \47118 , \47110 , \47117 );
not \g134071/U$4 ( \47119 , \47118 );
or \g134071/U$2 ( \47120 , \47103 , \47119 );
or \g134071/U$5 ( \47121 , \47118 , \46936 );
nand \g134071/U$1 ( \47122 , \47120 , \47121 );
xor \g456272/U$1_r1 ( \47123 , \47102 , \47122 );
xor \g133759/U$1 ( \47124 , \47093 , \47123 );
and \g133471/U$2 ( \47125 , \47087 , \47124 );
and \g133471/U$3 ( \47126 , \47093 , \47123 );
nor \g133471/U$1 ( \47127 , \47125 , \47126 );
not \g134653/U$3 ( \47128 , \46933 );
not \g134653/U$4 ( \47129 , \46937 );
and \g134653/U$2 ( \47130 , \47128 , \47129 );
and \g134653/U$5 ( \47131 , \46933 , \46937 );
nor \g134653/U$1 ( \47132 , \47130 , \47131 );
not \g134137/U$3 ( \47133 , \47117 );
not \g134137/U$4 ( \47134 , \46935 );
and \g134137/U$2 ( \47135 , \47133 , \47134 );
and \g134145/U$2 ( \47136 , \47117 , \46935 );
nor \g134145/U$1 ( \47137 , \47136 , \47110 );
nor \g134137/U$1 ( \47138 , \47135 , \47137 );
xnor \g133858/U$1 ( \47139 , \47132 , \47138 );
not \g133811/U$3 ( \47140 , \47139 );
and \g134765/U$2 ( \47141 , \42317 , \43757 );
and \g134765/U$3 ( \47142 , \43179 , \42316 );
nor \g134765/U$1 ( \47143 , \47141 , \47142 );
and \g134285/U$2 ( \47144 , \47143 , \42225 );
not \g134285/U$4 ( \47145 , \47143 );
and \g134285/U$3 ( \47146 , \47145 , \42226 );
nor \g134285/U$1 ( \47147 , \47144 , \47146 );
not \g134075/U$3 ( \47148 , \47147 );
and \g134758/U$2 ( \47149 , \42644 , \43183 );
and \g134758/U$3 ( \47150 , \42701 , \42643 );
nor \g134758/U$1 ( \47151 , \47149 , \47150 );
and \g134486/U$2 ( \47152 , \47151 , \42486 );
not \g134486/U$4 ( \47153 , \47151 );
and \g134486/U$3 ( \47154 , \47153 , \42487 );
nor \g134486/U$1 ( \47155 , \47152 , \47154 );
and \g134832/U$2 ( \47156 , \43099 , \42651 );
and \g134832/U$3 ( \47157 , \42609 , \43101 );
nor \g134832/U$1 ( \47158 , \47156 , \47157 );
and \g134385/U$2 ( \47159 , \47158 , \42681 );
not \g134385/U$4 ( \47160 , \47158 );
and \g134385/U$3 ( \47161 , \47160 , \42682 );
nor \g134385/U$1 ( \47162 , \47159 , \47161 );
xor \g134134/U$1 ( \47163 , \47155 , \47162 );
not \g134075/U$4 ( \47164 , \47163 );
or \g134075/U$2 ( \47165 , \47148 , \47164 );
or \g134075/U$5 ( \47166 , \47163 , \47147 );
nand \g134075/U$1 ( \47167 , \47165 , \47166 );
not \g133811/U$4 ( \47168 , \47167 );
and \g133811/U$2 ( \47169 , \47140 , \47168 );
and \g133811/U$5 ( \47170 , \47139 , \47167 );
nor \g133811/U$1 ( \47171 , \47169 , \47170 );
xor \g456272/U$4 ( \47172 , \47094 , \47101 );
and \g456272/U$3 ( \47173 , \47172 , \47122 );
and \g456272/U$5 ( \47174 , \47094 , \47101 );
nor \g456272/U$2 ( \47175 , \47173 , \47174 );
xnor \g133642/U$1 ( \47176 , \47171 , \47175 );
or \g133380/U$2 ( \47177 , \47127 , \47176 );
or \g133380/U$3 ( \47178 , \47175 , \47171 );
nand \g133380/U$1 ( \47179 , \47177 , \47178 );
or \g133762/U$2 ( \47180 , \47138 , \47132 );
not \g133817/U$3 ( \47181 , \47132 );
not \g133817/U$4 ( \47182 , \47138 );
or \g133817/U$2 ( \47183 , \47181 , \47182 );
nand \g133817/U$1 ( \47184 , \47183 , \47167 );
nand \g133762/U$1 ( \47185 , \47180 , \47184 );
xor \g134051/U$1 ( \47186 , \46926 , \46938 );
xor \g134051/U$1_r1 ( \47187 , \47186 , \46946 );
not \g133823/U$3 ( \47188 , \47187 );
not \g134098/U$3 ( \47189 , \47155 );
not \g134098/U$4 ( \47190 , \47147 );
and \g134098/U$2 ( \47191 , \47189 , \47190 );
and \g134104/U$2 ( \47192 , \47147 , \47155 );
nor \g134104/U$1 ( \47193 , \47192 , \47162 );
nor \g134098/U$1 ( \47194 , \47191 , \47193 );
not \g134120/U$3 ( \47195 , \46899 );
not \g134120/U$4 ( \47196 , \46888 );
and \g134120/U$2 ( \47197 , \47195 , \47196 );
and \g134120/U$5 ( \47198 , \46899 , \46888 );
nor \g134120/U$1 ( \47199 , \47197 , \47198 );
not \g134072/U$3 ( \47200 , \47199 );
not \g134072/U$4 ( \47201 , \46862 );
and \g134072/U$2 ( \47202 , \47200 , \47201 );
and \g134072/U$5 ( \47203 , \47199 , \46862 );
nor \g134072/U$1 ( \47204 , \47202 , \47203 );
xor \g133860/U$1 ( \47205 , \47194 , \47204 );
not \g133823/U$4 ( \47206 , \47205 );
or \g133823/U$2 ( \47207 , \47188 , \47206 );
or \g133823/U$5 ( \47208 , \47205 , \47187 );
nand \g133823/U$1 ( \47209 , \47207 , \47208 );
xor \g133643/U$1 ( \47210 , \47185 , \47209 );
and \g133300/U$2 ( \47211 , \47179 , \47210 );
and \g133300/U$3 ( \47212 , \47185 , \47209 );
nor \g133300/U$1 ( \47213 , \47211 , \47212 );
not \g133842/U$3 ( \47214 , \47187 );
not \g133842/U$4 ( \47215 , \47194 );
and \g133842/U$2 ( \47216 , \47214 , \47215 );
and \g133854/U$2 ( \47217 , \47187 , \47194 );
nor \g133854/U$1 ( \47218 , \47217 , \47204 );
nor \g133842/U$1 ( \47219 , \47216 , \47218 );
not \g133674/U$3 ( \47220 , \46965 );
xnor \g133861/U$1 ( \47221 , \46959 , \46949 );
not \g133674/U$4 ( \47222 , \47221 );
and \g133674/U$2 ( \47223 , \47220 , \47222 );
and \g133674/U$5 ( \47224 , \46965 , \47221 );
nor \g133674/U$1 ( \47225 , \47223 , \47224 );
xnor \g133601/U$1 ( \47226 , \47219 , \47225 );
or \g133245/U$2 ( \47227 , \47213 , \47226 );
or \g133245/U$3 ( \47228 , \47219 , \47225 );
nand \g133245/U$1 ( \47229 , \47227 , \47228 );
and \g133179/U$3 ( \47230 , \46969 , \47229 );
nor \g133179/U$1 ( \47231 , \46968 , \47230 );
xor \g456230/U$4 ( \47232 , \46913 , \46915 );
and \g456230/U$3 ( \47233 , \47232 , \46918 );
and \g456230/U$5 ( \47234 , \46913 , \46915 );
nor \g456230/U$2 ( \47235 , \47233 , \47234 );
not \g133666/U$3 ( \47236 , \46829 );
not \g133666/U$4 ( \47237 , \46877 );
or \g133666/U$2 ( \47238 , \47236 , \47237 );
or \g133666/U$5 ( \47239 , \46877 , \46829 );
nand \g133666/U$1 ( \47240 , \47238 , \47239 );
not \g133627/U$3 ( \47241 , \47240 );
not \g133627/U$4 ( \47242 , \46827 );
and \g133627/U$2 ( \47243 , \47241 , \47242 );
and \g133627/U$5 ( \47244 , \47240 , \46827 );
nor \g133627/U$1 ( \47245 , \47243 , \47244 );
xnor \g133505/U$1 ( \47246 , \47235 , \47245 );
or \g133126/U$2 ( \47247 , \47231 , \47246 );
or \g133126/U$3 ( \47248 , \47235 , \47245 );
nand \g133126/U$1 ( \47249 , \47247 , \47248 );
and \g133082/U$3 ( \47250 , \46881 , \47249 );
nor \g133082/U$1 ( \47251 , \46880 , \47250 );
xor \g456211/U$4 ( \47252 , \46807 , \46813 );
and \g456211/U$3 ( \47253 , \47252 , \46824 );
and \g456211/U$5 ( \47254 , \46807 , \46813 );
nor \g456211/U$2 ( \47255 , \47253 , \47254 );
not \g133520/U$3 ( \47256 , \46753 );
xor \g133602/U$1 ( \47257 , \46741 , \46735 );
not \g133520/U$4 ( \47258 , \47257 );
and \g133520/U$2 ( \47259 , \47256 , \47258 );
and \g133520/U$5 ( \47260 , \46753 , \47257 );
nor \g133520/U$1 ( \47261 , \47259 , \47260 );
xnor \g133439/U$1 ( \47262 , \47255 , \47261 );
or \g133035/U$2 ( \47263 , \47251 , \47262 );
or \g133035/U$3 ( \47264 , \47255 , \47261 );
nand \g133035/U$1 ( \47265 , \47263 , \47264 );
and \g132973/U$3 ( \47266 , \46758 , \47265 );
nor \g132973/U$1 ( \47267 , \46757 , \47266 );
or \g132921/U$3 ( \47268 , \46696 , \47267 );
nand \g132921/U$1 ( \47269 , \46695 , \47268 );
and \g132868/U$3 ( \47270 , \46605 , \47269 );
nor \g132868/U$1 ( \47271 , \46604 , \47270 );
or \g133521/U$1 ( \47272 , \46520 , \46427 );
and \g133442/U$2 ( \47273 , \46418 , \47272 );
and \g133442/U$3 ( \47274 , \46427 , \46520 );
nor \g133442/U$1 ( \47275 , \47273 , \47274 );
not \g133863/U$3 ( \47276 , \46231 );
not \g133863/U$4 ( \47277 , \46239 );
or \g133863/U$2 ( \47278 , \47276 , \47277 );
or \g133863/U$5 ( \47279 , \46239 , \46231 );
nand \g133863/U$1 ( \47280 , \47278 , \47279 );
not \g133830/U$3 ( \47281 , \47280 );
not \g133830/U$4 ( \47282 , \46233 );
and \g133830/U$2 ( \47283 , \47281 , \47282 );
and \g133830/U$5 ( \47284 , \47280 , \46233 );
nor \g133830/U$1 ( \47285 , \47283 , \47284 );
not \g133781/U$1 ( \47286 , \46333 );
and \g133657/U$2 ( \47287 , \47286 , \46368 );
not \g133662/U$3 ( \47288 , \47286 );
not \g133662/U$4 ( \47289 , \46368 );
and \g133662/U$2 ( \47290 , \47288 , \47289 );
nor \g133662/U$1 ( \47291 , \47290 , \46410 );
nor \g133657/U$1 ( \47292 , \47287 , \47291 );
xnor \g133501/U$1 ( \47293 , \47285 , \47292 );
not \g133443/U$3 ( \47294 , \47293 );
xor \g456215/U$2 ( \47295 , \46173 , \46191 );
xor \g456215/U$1 ( \47296 , \47295 , \46217 );
or \g133845/U$2 ( \47297 , \46313 , \46329 );
not \g133856/U$3 ( \47298 , \46329 );
not \g133856/U$4 ( \47299 , \46313 );
or \g133856/U$2 ( \47300 , \47298 , \47299 );
nand \g133856/U$1 ( \47301 , \47300 , \46287 );
nand \g133845/U$1 ( \47302 , \47297 , \47301 );
xor \g456239/U$9 ( \47303 , \46199 , \46206 );
xor \g456239/U$9_r1 ( \47304 , \47303 , \46214 );
and \g456239/U$8 ( \47305 , \46423 , \47304 );
xor \g456239/U$11 ( \47306 , \46199 , \46206 );
xor \g456239/U$11_r1 ( \47307 , \47306 , \46214 );
and \g456239/U$10 ( \47308 , \46425 , \47307 );
and \g456239/U$12 ( \47309 , \46423 , \46425 );
or \g456239/U$7 ( \47310 , \47305 , \47308 , \47309 );
xor \g456215/U$1_r1 ( \47311 , \47302 , \47310 );
xor \g456215/U$1_r2 ( \47312 , \47296 , \47311 );
not \g133443/U$4 ( \47313 , \47312 );
and \g133443/U$2 ( \47314 , \47294 , \47313 );
and \g133443/U$5 ( \47315 , \47293 , \47312 );
nor \g133443/U$1 ( \47316 , \47314 , \47315 );
xnor \g133376/U$1 ( \47317 , \47275 , \47316 );
or \g132794/U$2 ( \47318 , \47271 , \47317 );
or \g132794/U$3 ( \47319 , \47275 , \47316 );
nand \g132794/U$1 ( \47320 , \47318 , \47319 );
or \g133441/U$2 ( \47321 , \47292 , \47285 );
not \g133464/U$3 ( \47322 , \47285 );
not \g133464/U$4 ( \47323 , \47292 );
or \g133464/U$2 ( \47324 , \47322 , \47323 );
nand \g133464/U$1 ( \47325 , \47324 , \47312 );
nand \g133441/U$1 ( \47326 , \47321 , \47325 );
xor \g456232/U$1 ( \47327 , \46148 , \46220 );
xor \g456232/U$1_r1 ( \47328 , \47327 , \46241 );
not \g133413/U$3 ( \47329 , \47328 );
xor \g456237/U$2 ( \47330 , \45934 , \45941 );
xor \g456237/U$1 ( \47331 , \47330 , \45948 );
xor \g456237/U$1_r1 ( \47332 , \46118 , \46131 );
xor \g456237/U$1_r2 ( \47333 , \47331 , \47332 );
xor \g456215/U$9 ( \47334 , \46173 , \46191 );
xor \g456215/U$9_r1 ( \47335 , \47334 , \46217 );
and \g456215/U$8 ( \47336 , \47302 , \47335 );
xor \g456215/U$11 ( \47337 , \46173 , \46191 );
xor \g456215/U$11_r1 ( \47338 , \47337 , \46217 );
and \g456215/U$10 ( \47339 , \47310 , \47338 );
and \g456215/U$12 ( \47340 , \47302 , \47310 );
or \g456215/U$7 ( \47341 , \47336 , \47339 , \47340 );
xnor \g133486/U$1 ( \47342 , \47333 , \47341 );
not \g133413/U$4 ( \47343 , \47342 );
or \g133413/U$2 ( \47344 , \47329 , \47343 );
or \g133413/U$5 ( \47345 , \47342 , \47328 );
nand \g133413/U$1 ( \47346 , \47344 , \47345 );
xor \g133355/U$1 ( \47347 , \47326 , \47346 );
and \g132734/U$2 ( \47348 , \47320 , \47347 );
and \g132734/U$3 ( \47349 , \47326 , \47346 );
nor \g132734/U$1 ( \47350 , \47348 , \47349 );
and \g133412/U$2 ( \47351 , \47341 , \47333 );
or \g133496/U$1 ( \47352 , \47341 , \47333 );
and \g133412/U$3 ( \47353 , \47328 , \47352 );
nor \g133412/U$1 ( \47354 , \47351 , \47353 );
not \g133451/U$3 ( \47355 , \46256 );
xnor \g133503/U$1 ( \47356 , \46250 , \46244 );
not \g133451/U$4 ( \47357 , \47356 );
and \g133451/U$2 ( \47358 , \47355 , \47357 );
and \g133451/U$5 ( \47359 , \46256 , \47356 );
nor \g133451/U$1 ( \47360 , \47358 , \47359 );
xnor \g133356/U$1 ( \47361 , \47354 , \47360 );
or \g132670/U$2 ( \47362 , \47350 , \47361 );
or \g132670/U$3 ( \47363 , \47354 , \47360 );
nand \g132670/U$1 ( \47364 , \47362 , \47363 );
and \g132583/U$3 ( \47365 , \46260 , \47364 );
nor \g132583/U$1 ( \47366 , \46259 , \47365 );
and \g133393/U$2 ( \47367 , \46139 , \46058 );
or \g133481/U$1 ( \47368 , \46139 , \46058 );
and \g133393/U$3 ( \47369 , \47368 , \45995 );
nor \g133393/U$1 ( \47370 , \47367 , \47369 );
xor \g456207/U$9 ( \47371 , \45765 , \45790 );
xor \g456207/U$9_r1 ( \47372 , \47371 , \45816 );
and \g456207/U$8 ( \47373 , \45881 , \47372 );
xor \g456207/U$11 ( \47374 , \45765 , \45790 );
xor \g456207/U$11_r1 ( \47375 , \47374 , \45816 );
and \g456207/U$10 ( \47376 , \45993 , \47375 );
and \g456207/U$12 ( \47377 , \45881 , \45993 );
or \g456207/U$7 ( \47378 , \47373 , \47376 , \47377 );
not \g133410/U$3 ( \47379 , \47378 );
and \g133624/U$2 ( \47380 , \45954 , \45907 );
not \g133636/U$3 ( \47381 , \45954 );
not \g133636/U$4 ( \47382 , \45907 );
and \g133636/U$2 ( \47383 , \47381 , \47382 );
nor \g133636/U$1 ( \47384 , \47383 , \45988 );
nor \g133624/U$1 ( \47385 , \47380 , \47384 );
not \g133410/U$4 ( \47386 , \47385 );
and \g133410/U$2 ( \47387 , \47379 , \47386 );
and \g133410/U$5 ( \47388 , \47378 , \47385 );
nor \g133410/U$1 ( \47389 , \47387 , \47388 );
not \g133381/U$3 ( \47390 , \47389 );
xor \g456257/U$9 ( \47391 , \45824 , \45669 );
xor \g456257/U$9_r1 ( \47392 , \47391 , \45832 );
and \g456257/U$8 ( \47393 , \45856 , \47392 );
xor \g456257/U$11 ( \47394 , \45824 , \45669 );
xor \g456257/U$11_r1 ( \47395 , \47394 , \45832 );
and \g456257/U$10 ( \47396 , \45879 , \47395 );
and \g456257/U$12 ( \47397 , \45856 , \45879 );
or \g456257/U$7 ( \47398 , \47393 , \47396 , \47397 );
xor \g456260/U$2 ( \47399 , \45606 , \45613 );
xor \g456260/U$1 ( \47400 , \47399 , \45621 );
xor \g133973/U$4 ( \47401 , \45888 , \45898 );
and \g133973/U$3 ( \47402 , \47401 , \45906 );
and \g133973/U$5 ( \47403 , \45888 , \45898 );
or \g133973/U$2 ( \47404 , \47402 , \47403 );
xor \g133950/U$1 ( \47405 , \45686 , \45693 );
xor \g133950/U$1_r1 ( \47406 , \47405 , \45701 );
xor \g456260/U$1_r1 ( \47407 , \47404 , \47406 );
xor \g456260/U$1_r2 ( \47408 , \47400 , \47407 );
xor \g133494/U$1 ( \47409 , \47398 , \47408 );
xor \g133896/U$4 ( \47410 , \45840 , \45847 );
and \g133896/U$3 ( \47411 , \47410 , \45855 );
and \g133896/U$5 ( \47412 , \45840 , \45847 );
or \g133896/U$2 ( \47413 , \47411 , \47412 );
xor \g456257/U$5 ( \47414 , \45824 , \45669 );
and \g456257/U$4 ( \47415 , \47414 , \45832 );
and \g456257/U$6 ( \47416 , \45824 , \45669 );
or \g456257/U$3 ( \47417 , \47415 , \47416 );
xor \g456218/U$2 ( \47418 , \47413 , \47417 );
xor \g133965/U$1 ( \47419 , \45650 , \45657 );
xor \g133965/U$1_r1 ( \47420 , \47419 , \45665 );
xor \g456218/U$1 ( \47421 , \47418 , \47420 );
xor \g456207/U$5 ( \47422 , \45765 , \45790 );
and \g456207/U$4 ( \47423 , \47422 , \45816 );
and \g456207/U$6 ( \47424 , \45765 , \45790 );
or \g456207/U$3 ( \47425 , \47423 , \47424 );
xor \g134093/U$1 ( \47426 , \45670 , \45677 );
and \g134716/U$2 ( \47427 , \41087 , \41920 );
and \g134716/U$3 ( \47428 , \41774 , \41328 );
nor \g134716/U$1 ( \47429 , \47427 , \47428 );
and \g134477/U$2 ( \47430 , \47429 , \41093 );
not \g134477/U$4 ( \47431 , \47429 );
and \g134477/U$3 ( \47432 , \47431 , \41092 );
nor \g134477/U$1 ( \47433 , \47430 , \47432 );
xor \g133797/U$1 ( \47434 , \47426 , \47433 );
xor \g133998/U$4 ( \47435 , \45863 , \45870 );
and \g133998/U$3 ( \47436 , \47435 , \45878 );
and \g133998/U$5 ( \47437 , \45863 , \45870 );
or \g133998/U$2 ( \47438 , \47436 , \47437 );
xor \g133797/U$1_r1 ( \47439 , \47434 , \47438 );
xor \g456218/U$1_r1 ( \47440 , \47425 , \47439 );
xor \g456218/U$1_r2 ( \47441 , \47421 , \47440 );
xor \g133494/U$1_r1 ( \47442 , \47409 , \47441 );
not \g133381/U$4 ( \47443 , \47442 );
and \g133381/U$2 ( \47444 , \47390 , \47443 );
and \g133381/U$5 ( \47445 , \47389 , \47442 );
nor \g133381/U$1 ( \47446 , \47444 , \47445 );
xnor \g133325/U$1 ( \47447 , \47370 , \47446 );
or \g132513/U$2 ( \47448 , \47366 , \47447 );
or \g132513/U$3 ( \47449 , \47370 , \47446 );
nand \g132513/U$1 ( \47450 , \47448 , \47449 );
not \g133493/U$1 ( \47451 , \47442 );
or \g133411/U$2 ( \47452 , \47451 , \47385 );
not \g133433/U$3 ( \47453 , \47385 );
not \g133433/U$4 ( \47454 , \47451 );
or \g133433/U$2 ( \47455 , \47453 , \47454 );
nand \g133433/U$1 ( \47456 , \47455 , \47378 );
nand \g133411/U$1 ( \47457 , \47452 , \47456 );
xor \g133494/U$4 ( \47458 , \47398 , \47408 );
and \g133494/U$3 ( \47459 , \47458 , \47441 );
and \g133494/U$5 ( \47460 , \47398 , \47408 );
or \g133494/U$2 ( \47461 , \47459 , \47460 );
xor \g456260/U$9 ( \47462 , \45606 , \45613 );
xor \g456260/U$9_r1 ( \47463 , \47462 , \45621 );
and \g456260/U$8 ( \47464 , \47404 , \47463 );
xor \g456260/U$11 ( \47465 , \45606 , \45613 );
xor \g456260/U$11_r1 ( \47466 , \47465 , \45621 );
and \g456260/U$10 ( \47467 , \47406 , \47466 );
and \g456260/U$12 ( \47468 , \47404 , \47406 );
or \g456260/U$7 ( \47469 , \47464 , \47467 , \47468 );
xor \g456218/U$5 ( \47470 , \47413 , \47417 );
and \g456218/U$4 ( \47471 , \47470 , \47420 );
and \g456218/U$6 ( \47472 , \47413 , \47417 );
or \g456218/U$3 ( \47473 , \47471 , \47472 );
xor \g133536/U$1 ( \47474 , \47469 , \47473 );
xor \g133773/U$1 ( \47475 , \45668 , \45678 );
xor \g133773/U$1_r1 ( \47476 , \47475 , \45704 );
xor \g133536/U$1_r1 ( \47477 , \47474 , \47476 );
xor \g133370/U$1 ( \47478 , \47461 , \47477 );
xor \g134003/U$1 ( \47479 , \45536 , \45275 );
xor \g134003/U$1_r1 ( \47480 , \47479 , \45544 );
xor \g133930/U$1 ( \47481 , \45510 , \45517 );
xor \g133930/U$1_r1 ( \47482 , \47481 , \45525 );
xor \g456205/U$2 ( \47483 , \47480 , \47482 );
xor \g133797/U$4 ( \47484 , \47426 , \47433 );
and \g133797/U$3 ( \47485 , \47484 , \47438 );
and \g133797/U$5 ( \47486 , \47426 , \47433 );
or \g133797/U$2 ( \47487 , \47485 , \47486 );
xor \g456205/U$1 ( \47488 , \47483 , \47487 );
xor \g133790/U$1 ( \47489 , \45599 , \45624 );
xor \g133790/U$1_r1 ( \47490 , \47489 , \45627 );
xor \g456218/U$9 ( \47491 , \47413 , \47417 );
xor \g456218/U$9_r1 ( \47492 , \47491 , \47420 );
and \g456218/U$8 ( \47493 , \47425 , \47492 );
xor \g456218/U$11 ( \47494 , \47413 , \47417 );
xor \g456218/U$11_r1 ( \47495 , \47494 , \47420 );
and \g456218/U$10 ( \47496 , \47439 , \47495 );
and \g456218/U$12 ( \47497 , \47425 , \47439 );
or \g456218/U$7 ( \47498 , \47493 , \47496 , \47497 );
xor \g456205/U$1_r1 ( \47499 , \47490 , \47498 );
xor \g456205/U$1_r2 ( \47500 , \47488 , \47499 );
xor \g133370/U$1_r1 ( \47501 , \47478 , \47500 );
xor \g133326/U$1 ( \47502 , \47457 , \47501 );
and \g132440/U$2 ( \47503 , \47450 , \47502 );
and \g132440/U$3 ( \47504 , \47457 , \47501 );
nor \g132440/U$1 ( \47505 , \47503 , \47504 );
not \g132439/U$1 ( \47506 , \47505 );
xor \g456205/U$9 ( \47507 , \47480 , \47482 );
xor \g456205/U$9_r1 ( \47508 , \47507 , \47487 );
and \g456205/U$8 ( \47509 , \47490 , \47508 );
xor \g456205/U$11 ( \47510 , \47480 , \47482 );
xor \g456205/U$11_r1 ( \47511 , \47510 , \47487 );
and \g456205/U$10 ( \47512 , \47498 , \47511 );
and \g456205/U$12 ( \47513 , \47490 , \47498 );
or \g456205/U$7 ( \47514 , \47509 , \47512 , \47513 );
xor \g133536/U$4 ( \47515 , \47469 , \47473 );
and \g133536/U$3 ( \47516 , \47515 , \47476 );
and \g133536/U$5 ( \47517 , \47469 , \47473 );
or \g133536/U$2 ( \47518 , \47516 , \47517 );
xor \g456188/U$1 ( \47519 , \47514 , \47518 );
xor \g456214/U$2 ( \47520 , \45503 , \45528 );
xor \g456214/U$1 ( \47521 , \47520 , \45547 );
xor \g456214/U$1_r1 ( \47522 , \45630 , \45639 );
xor \g456214/U$1_r2 ( \47523 , \47521 , \47522 );
not \g133450/U$3 ( \47524 , \47523 );
xor \g456205/U$5 ( \47525 , \47480 , \47482 );
and \g456205/U$4 ( \47526 , \47525 , \47487 );
and \g456205/U$6 ( \47527 , \47480 , \47482 );
or \g456205/U$3 ( \47528 , \47526 , \47527 );
xor \g133584/U$1 ( \47529 , \45707 , \45713 );
xor \g133584/U$1_r1 ( \47530 , \47529 , \45716 );
xnor \g133498/U$1 ( \47531 , \47528 , \47530 );
not \g133450/U$4 ( \47532 , \47531 );
or \g133450/U$2 ( \47533 , \47524 , \47532 );
or \g133450/U$5 ( \47534 , \47531 , \47523 );
nand \g133450/U$1 ( \47535 , \47533 , \47534 );
xor \g456188/U$1_r1 ( \47536 , \47519 , \47535 );
xor \g133370/U$4 ( \47537 , \47461 , \47477 );
and \g133370/U$3 ( \47538 , \47537 , \47500 );
and \g133370/U$5 ( \47539 , \47461 , \47477 );
or \g133370/U$2 ( \47540 , \47538 , \47539 );
xor \g133284/U$1 ( \47541 , \47536 , \47540 );
and \g132315/U$2 ( \47542 , \47506 , \47541 );
and \g132315/U$3 ( \47543 , \47536 , \47540 );
nor \g132315/U$1 ( \47544 , \47542 , \47543 );
xor \g456188/U$4 ( \47545 , \47514 , \47518 );
and \g456188/U$3 ( \47546 , \47545 , \47535 );
and \g456188/U$5 ( \47547 , \47514 , \47518 );
nor \g456188/U$2 ( \47548 , \47546 , \47547 );
xnor \g133639/U$1 ( \47549 , \45468 , \45423 );
not \g133561/U$3 ( \47550 , \47549 );
not \g133561/U$4 ( \47551 , \45476 );
and \g133561/U$2 ( \47552 , \47550 , \47551 );
and \g133561/U$5 ( \47553 , \47549 , \45476 );
nor \g133561/U$1 ( \47554 , \47552 , \47553 );
and \g133446/U$2 ( \47555 , \47530 , \47528 );
or \g133522/U$1 ( \47556 , \47530 , \47528 );
and \g133446/U$3 ( \47557 , \47523 , \47556 );
nor \g133446/U$1 ( \47558 , \47555 , \47557 );
xnor \g133373/U$1 ( \47559 , \47554 , \47558 );
not \g133330/U$3 ( \47560 , \47559 );
xor \g133428/U$1 ( \47561 , \45644 , \45719 );
xor \g133428/U$1_r1 ( \47562 , \47561 , \45722 );
not \g133330/U$4 ( \47563 , \47562 );
and \g133330/U$2 ( \47564 , \47560 , \47563 );
and \g133330/U$5 ( \47565 , \47559 , \47562 );
nor \g133330/U$1 ( \47566 , \47564 , \47565 );
xnor \g133275/U$1 ( \47567 , \47548 , \47566 );
or \g132236/U$2 ( \47568 , \47544 , \47567 );
or \g132236/U$3 ( \47569 , \47548 , \47566 );
nand \g132236/U$1 ( \47570 , \47568 , \47569 );
or \g133327/U$2 ( \47571 , \47558 , \47554 );
not \g133343/U$3 ( \47572 , \47554 );
not \g133343/U$4 ( \47573 , \47558 );
or \g133343/U$2 ( \47574 , \47572 , \47573 );
nand \g133343/U$1 ( \47575 , \47574 , \47562 );
nand \g133327/U$1 ( \47576 , \47571 , \47575 );
xor \g133308/U$1 ( \47577 , \45725 , \45729 );
xor \g133308/U$1_r1 ( \47578 , \47577 , \45732 );
xor \g133276/U$1 ( \47579 , \47576 , \47578 );
and \g132142/U$2 ( \47580 , \47570 , \47579 );
and \g132142/U$3 ( \47581 , \47576 , \47578 );
nor \g132142/U$1 ( \47582 , \47580 , \47581 );
xnor \g133277/U$1 ( \47583 , \45735 , \45738 );
or \g132057/U$5 ( \47584 , \47582 , \47583 );
nand \g132057/U$1 ( \47585 , \45740 , \47584 );
and \g131990/U$3 ( \47586 , \45593 , \47585 );
nor \g131990/U$1 ( \47587 , \45592 , \47586 );
xnor \g133259/U$1 ( \47588 , \45412 , \45417 );
or \g131911/U$5 ( \47589 , \47587 , \47588 );
nand \g131911/U$1 ( \47590 , \45419 , \47589 );
and \g131836/U$3 ( \47591 , \45262 , \47590 );
nor \g131836/U$1 ( \47592 , \45261 , \47591 );
xnor \g133231/U$1 ( \47593 , \45100 , \45103 );
or \g131774/U$5 ( \47594 , \47592 , \47593 );
nand \g131774/U$1 ( \47595 , \45105 , \47594 );
and \g131712/U$3 ( \47596 , \44897 , \47595 );
nor \g131712/U$1 ( \47597 , \44896 , \47596 );
not \g131711/U$1 ( \47598 , \47597 );
xor \g456176/U$9 ( \47599 , \44675 , \44679 );
xor \g456176/U$9_r1 ( \47600 , \47599 , \44694 );
and \g456176/U$8 ( \47601 , \44889 , \47600 );
xor \g456176/U$11 ( \47602 , \44675 , \44679 );
xor \g456176/U$11_r1 ( \47603 , \47602 , \44694 );
and \g456176/U$10 ( \47604 , \44893 , \47603 );
and \g456176/U$12 ( \47605 , \44889 , \44893 );
or \g456176/U$7 ( \47606 , \47601 , \47604 , \47605 );
xor \g133243/U$1 ( \47607 , \44653 , \44697 );
xor \g133243/U$1_r1 ( \47608 , \47607 , \44702 );
xor \g133197/U$1 ( \47609 , \47606 , \47608 );
and \g131649/U$2 ( \47610 , \47598 , \47609 );
and \g131649/U$3 ( \47611 , \47606 , \47608 );
nor \g131649/U$1 ( \47612 , \47610 , \47611 );
xnor \g133177/U$1 ( \47613 , \44705 , \44708 );
or \g131591/U$5 ( \47614 , \47612 , \47613 );
nand \g131591/U$1 ( \47615 , \44710 , \47614 );
and \g131534/U$3 ( \47616 , \44367 , \47615 );
nor \g131534/U$1 ( \47617 , \44366 , \47616 );
not \g131533/U$1 ( \47618 , \47617 );
and \g131466/U$3 ( \47619 , \44335 , \47618 );
nor \g131466/U$1 ( \47620 , \44334 , \47619 );
not \g131465/U$1 ( \47621 , \47620 );
and \g131394/U$3 ( \47622 , \44104 , \47621 );
nor \g131394/U$1 ( \47623 , \44103 , \47622 );
xor \g133188/U$1 ( \47624 , \43899 , \43902 );
not \g133174/U$1 ( \47625 , \47624 );
or \g131337/U$5 ( \47626 , \47623 , \47625 );
nand \g131337/U$1 ( \47627 , \43904 , \47626 );
and \g131283/U$3 ( \47628 , \43668 , \47627 );
nor \g131283/U$1 ( \47629 , \43667 , \47628 );
xor \g133183/U$1 ( \47630 , \43455 , \43452 );
not \g133173/U$1 ( \47631 , \47630 );
or \g131224/U$5 ( \47632 , \47629 , \47631 );
nand \g131224/U$1 ( \47633 , \43457 , \47632 );
and \g131166/U$3 ( \47634 , \43059 , \47633 );
nor \g131166/U$1 ( \47635 , \43058 , \47634 );
xor \g133206/U$1 ( \47636 , \42923 , \42940 );
not \g133181/U$1 ( \47637 , \47636 );
or \g131082/U$5 ( \47638 , \47635 , \47637 );
nand \g131082/U$1 ( \47639 , \42942 , \47638 );
xor \g133217/U$1 ( \47640 , \42584 , \42586 );
xor \g133217/U$1_r1 ( \47641 , \47640 , \42591 );
xor \g133244/U$4 ( \47642 , \42932 , \42934 );
and \g133244/U$3 ( \47643 , \47642 , \42939 );
and \g133244/U$5 ( \47644 , \42932 , \42934 );
or \g133244/U$2 ( \47645 , \47643 , \47644 );
xor \g133187/U$1 ( \47646 , \47641 , \47645 );
and \g131002/U$2 ( \47647 , \47639 , \47646 );
and \g131002/U$3 ( \47648 , \47641 , \47645 );
nor \g131002/U$1 ( \47649 , \47647 , \47648 );
not \g131001/U$1 ( \47650 , \47649 );
and \g130945/U$3 ( \47651 , \42596 , \47650 );
nor \g130945/U$1 ( \47652 , \42595 , \47651 );
xor \g133207/U$1 ( \47653 , \42391 , \42394 );
not \g133182/U$1 ( \47654 , \47653 );
or \g130890/U$5 ( \47655 , \47652 , \47654 );
nand \g130890/U$1 ( \47656 , \42396 , \47655 );
and \g130836/U$3 ( \47657 , \42174 , \47656 );
nor \g130836/U$1 ( \47658 , \42173 , \47657 );
xor \g133219/U$1 ( \47659 , \42011 , \42014 );
not \g133204/U$1 ( \47660 , \47659 );
or \g130777/U$5 ( \47661 , \47658 , \47660 );
nand \g130777/U$1 ( \47662 , \42016 , \47661 );
and \g130724/U$3 ( \47663 , \41708 , \47662 );
nor \g130724/U$1 ( \47664 , \41707 , \47663 );
not \g130723/U$1 ( \47665 , \47664 );
xor \g133301/U$4 ( \47666 , \41427 , \41525 );
and \g133301/U$3 ( \47667 , \47666 , \41610 );
and \g133301/U$5 ( \47668 , \41427 , \41525 );
or \g133301/U$2 ( \47669 , \47667 , \47668 );
xor \g456198/U$9 ( \47670 , \41549 , \41565 );
xor \g456198/U$9_r1 ( \47671 , \47670 , \41579 );
and \g456198/U$8 ( \47672 , \41588 , \47671 );
xor \g456198/U$11 ( \47673 , \41549 , \41565 );
xor \g456198/U$11_r1 ( \47674 , \47673 , \41579 );
and \g456198/U$10 ( \47675 , \41608 , \47674 );
and \g456198/U$12 ( \47676 , \41588 , \41608 );
or \g456198/U$7 ( \47677 , \47672 , \47675 , \47676 );
xor \g133710/U$4 ( \47678 , \41500 , \41504 );
and \g133710/U$3 ( \47679 , \47678 , \41523 );
and \g133710/U$5 ( \47680 , \41500 , \41504 );
or \g133710/U$2 ( \47681 , \47679 , \47680 );
xor \g133727/U$4 ( \47682 , \41573 , \41486 );
and \g133727/U$3 ( \47683 , \47682 , \41578 );
and \g133727/U$5 ( \47684 , \41573 , \41486 );
or \g133727/U$2 ( \47685 , \47683 , \47684 );
xor \g133583/U$1 ( \47686 , \47681 , \47685 );
xor \g133937/U$4 ( \47687 , \41556 , \41215 );
and \g133937/U$3 ( \47688 , \47687 , \41564 );
and \g133937/U$5 ( \47689 , \41556 , \41215 );
or \g133937/U$2 ( \47690 , \47688 , \47689 );
xor \g133991/U$4 ( \47691 , \41512 , \41514 );
and \g133991/U$3 ( \47692 , \47691 , \41522 );
and \g133991/U$5 ( \47693 , \41512 , \41514 );
or \g133991/U$2 ( \47694 , \47692 , \47693 );
xor \g133706/U$1 ( \47695 , \47690 , \47694 );
xor \g134004/U$4 ( \47696 , \41533 , \41540 );
and \g134004/U$3 ( \47697 , \47696 , \41548 );
and \g134004/U$5 ( \47698 , \41533 , \41540 );
or \g134004/U$2 ( \47699 , \47697 , \47698 );
xor \g133706/U$1_r1 ( \47700 , \47695 , \47699 );
xor \g133583/U$1_r1 ( \47701 , \47686 , \47700 );
xor \g133332/U$1 ( \47702 , \47677 , \47701 );
xor \g456198/U$5 ( \47703 , \41549 , \41565 );
and \g456198/U$4 ( \47704 , \47703 , \41579 );
and \g456198/U$6 ( \47705 , \41549 , \41565 );
or \g456198/U$3 ( \47706 , \47704 , \47705 );
and \g134744/U$2 ( \47707 , \40175 , \40525 );
and \g134744/U$3 ( \47708 , \40472 , \40207 );
nor \g134744/U$1 ( \47709 , \47707 , \47708 );
and \g134315/U$2 ( \47710 , \47709 , \40137 );
not \g134315/U$4 ( \47711 , \47709 );
and \g134315/U$3 ( \47712 , \47711 , \40136 );
nor \g134315/U$1 ( \47713 , \47710 , \47712 );
not \g134670/U$1 ( \47714 , \40984 );
xor \g456253/U$2 ( \47715 , \47713 , \47714 );
and \g135010/U$2 ( \47716 , \40147 , \40731 );
and \g135010/U$3 ( \47717 , \40568 , \40149 );
nor \g135010/U$1 ( \47718 , \47716 , \47717 );
and \g134420/U$2 ( \47719 , \47718 , \40107 );
not \g134420/U$4 ( \47720 , \47718 );
and \g134420/U$3 ( \47721 , \47720 , \40106 );
nor \g134420/U$1 ( \47722 , \47719 , \47721 );
xor \g456253/U$1 ( \47723 , \47715 , \47722 );
xor \g134032/U$1 ( \47724 , \40992 , \40999 );
xor \g134032/U$1_r1 ( \47725 , \47724 , \41007 );
xor \g133989/U$1 ( \47726 , \40955 , \40958 );
xor \g133989/U$1_r1 ( \47727 , \47726 , \40966 );
xor \g456253/U$1_r1 ( \47728 , \47725 , \47727 );
xor \g456253/U$1_r2 ( \47729 , \47723 , \47728 );
xor \g133461/U$1 ( \47730 , \47706 , \47729 );
xor \g133586/U$4 ( \47731 , \41477 , \41495 );
and \g133586/U$3 ( \47732 , \47731 , \41524 );
and \g133586/U$5 ( \47733 , \41477 , \41495 );
or \g133586/U$2 ( \47734 , \47732 , \47733 );
xor \g133461/U$1_r1 ( \47735 , \47730 , \47734 );
xor \g133332/U$1_r1 ( \47736 , \47702 , \47735 );
xor \g133281/U$1 ( \47737 , \47669 , \47736 );
and \g130666/U$2 ( \47738 , \47665 , \47737 );
and \g130666/U$3 ( \47739 , \47669 , \47736 );
nor \g130666/U$1 ( \47740 , \47738 , \47739 );
not \g130665/U$1 ( \47741 , \47740 );
xor \g133461/U$4 ( \47742 , \47706 , \47729 );
and \g133461/U$3 ( \47743 , \47742 , \47734 );
and \g133461/U$5 ( \47744 , \47706 , \47729 );
or \g133461/U$2 ( \47745 , \47743 , \47744 );
xor \g133706/U$4 ( \47746 , \47690 , \47694 );
and \g133706/U$3 ( \47747 , \47746 , \47699 );
and \g133706/U$5 ( \47748 , \47690 , \47694 );
or \g133706/U$2 ( \47749 , \47747 , \47748 );
xor \g456253/U$5 ( \47750 , \47713 , \47714 );
and \g456253/U$4 ( \47751 , \47750 , \47722 );
and \g456253/U$6 ( \47752 , \47713 , \47714 );
or \g456253/U$3 ( \47753 , \47751 , \47752 );
xor \g133551/U$1 ( \47754 , \47749 , \47753 );
xor \g133798/U$1 ( \47755 , \40969 , \40984 );
xor \g133798/U$1_r1 ( \47756 , \47755 , \41010 );
xor \g133551/U$1_r1 ( \47757 , \47754 , \47756 );
xor \g133341/U$1 ( \47758 , \47745 , \47757 );
xor \g456204/U$2 ( \47759 , \41041 , \41043 );
xor \g456204/U$1 ( \47760 , \47759 , \41046 );
xor \g456253/U$9 ( \47761 , \47713 , \47714 );
xor \g456253/U$9_r1 ( \47762 , \47761 , \47722 );
and \g456253/U$8 ( \47763 , \47725 , \47762 );
xor \g456253/U$11 ( \47764 , \47713 , \47714 );
xor \g456253/U$11_r1 ( \47765 , \47764 , \47722 );
and \g456253/U$10 ( \47766 , \47727 , \47765 );
and \g456253/U$12 ( \47767 , \47725 , \47727 );
or \g456253/U$7 ( \47768 , \47763 , \47766 , \47767 );
xor \g133583/U$4 ( \47769 , \47681 , \47685 );
and \g133583/U$3 ( \47770 , \47769 , \47700 );
and \g133583/U$5 ( \47771 , \47681 , \47685 );
or \g133583/U$2 ( \47772 , \47770 , \47771 );
xor \g456204/U$1_r1 ( \47773 , \47768 , \47772 );
xor \g456204/U$1_r2 ( \47774 , \47760 , \47773 );
xor \g133341/U$1_r1 ( \47775 , \47758 , \47774 );
xor \g133332/U$4 ( \47776 , \47677 , \47701 );
and \g133332/U$3 ( \47777 , \47776 , \47735 );
and \g133332/U$5 ( \47778 , \47677 , \47701 );
or \g133332/U$2 ( \47779 , \47777 , \47778 );
xor \g133298/U$1 ( \47780 , \47775 , \47779 );
and \g130600/U$2 ( \47781 , \47741 , \47780 );
and \g130600/U$3 ( \47782 , \47775 , \47779 );
nor \g130600/U$1 ( \47783 , \47781 , \47782 );
not \g130599/U$1 ( \47784 , \47783 );
xor \g133341/U$4 ( \47785 , \47745 , \47757 );
and \g133341/U$3 ( \47786 , \47785 , \47774 );
and \g133341/U$5 ( \47787 , \47745 , \47757 );
or \g133341/U$2 ( \47788 , \47786 , \47787 );
xor \g456190/U$2 ( \47789 , \41039 , \41049 );
xor \g456190/U$1 ( \47790 , \47789 , \41052 );
xor \g133551/U$4 ( \47791 , \47749 , \47753 );
and \g133551/U$3 ( \47792 , \47791 , \47756 );
and \g133551/U$5 ( \47793 , \47749 , \47753 );
or \g133551/U$2 ( \47794 , \47792 , \47793 );
xor \g456204/U$9 ( \47795 , \41041 , \41043 );
xor \g456204/U$9_r1 ( \47796 , \47795 , \41046 );
and \g456204/U$8 ( \47797 , \47768 , \47796 );
xor \g456204/U$11 ( \47798 , \41041 , \41043 );
xor \g456204/U$11_r1 ( \47799 , \47798 , \41046 );
and \g456204/U$10 ( \47800 , \47772 , \47799 );
and \g456204/U$12 ( \47801 , \47768 , \47772 );
or \g456204/U$7 ( \47802 , \47797 , \47800 , \47801 );
xor \g456190/U$1_r1 ( \47803 , \47794 , \47802 );
xor \g456190/U$1_r2 ( \47804 , \47790 , \47803 );
xor \g133297/U$1 ( \47805 , \47788 , \47804 );
and \g130535/U$2 ( \47806 , \47784 , \47805 );
and \g130535/U$3 ( \47807 , \47788 , \47804 );
nor \g130535/U$1 ( \47808 , \47806 , \47807 );
not \g130534/U$1 ( \47809 , \47808 );
xor \g456190/U$9 ( \47810 , \41039 , \41049 );
xor \g456190/U$9_r1 ( \47811 , \47810 , \41052 );
and \g456190/U$8 ( \47812 , \47794 , \47811 );
xor \g456190/U$11 ( \47813 , \41039 , \41049 );
xor \g456190/U$11_r1 ( \47814 , \47813 , \41052 );
and \g456190/U$10 ( \47815 , \47802 , \47814 );
and \g456190/U$12 ( \47816 , \47794 , \47802 );
or \g456190/U$7 ( \47817 , \47812 , \47815 , \47816 );
xor \g133383/U$1 ( \47818 , \41055 , \41059 );
xor \g133383/U$1_r1 ( \47819 , \47818 , \41064 );
xor \g133311/U$1 ( \47820 , \47817 , \47819 );
and \g130465/U$2 ( \47821 , \47809 , \47820 );
and \g130465/U$3 ( \47822 , \47817 , \47819 );
nor \g130465/U$1 ( \47823 , \47821 , \47822 );
not \g130464/U$1 ( \47824 , \47823 );
and \g130400/U$3 ( \47825 , \41069 , \47824 );
nor \g130400/U$1 ( \47826 , \41068 , \47825 );
xnor \g133328/U$1 ( \47827 , \40841 , \41031 );
or \g130319/U$5 ( \47828 , \47826 , \47827 );
nand \g130319/U$1 ( \47829 , \41033 , \47828 );
and \g130256/U$3 ( \47830 , \40839 , \47829 );
nor \g130256/U$1 ( \47831 , \40838 , \47830 );
xnor \g133378/U$1 ( \47832 , \40655 , \40761 );
or \g130180/U$5 ( \47833 , \47831 , \47832 );
nand \g130180/U$1 ( \47834 , \40763 , \47833 );
and \g130105/U$3 ( \47835 , \40653 , \47834 );
nor \g130105/U$1 ( \47836 , \40652 , \47835 );
xnor \g133468/U$1 ( \47837 , \40494 , \40499 );
or \g130012/U$5 ( \47838 , \47836 , \47837 );
nand \g130012/U$1 ( \47839 , \40501 , \47838 );
and \g129915/U$3 ( \47840 , \40415 , \47839 );
nor \g129915/U$1 ( \47841 , \40414 , \47840 );
or \g129824/U$3 ( \47842 , \40337 , \47841 );
nand \g129824/U$1 ( \47843 , \40336 , \47842 );
and \g129735/U$3 ( \47844 , \40268 , \47843 );
nor \g129735/U$1 ( \47845 , \40267 , \47844 );
xor \g134006/U$4 ( \47846 , \40245 , \40247 );
and \g134006/U$3 ( \47847 , \47846 , \40255 );
and \g134006/U$5 ( \47848 , \40245 , \40247 );
or \g134006/U$2 ( \47849 , \47847 , \47848 );
and \g135566/U$2 ( \47850 , \40245 , \47849 );
not \g135566/U$4 ( \47851 , \40245 );
not \g134005/U$1 ( \47852 , \47849 );
and \g135566/U$3 ( \47853 , \47851 , \47852 );
nor \g135566/U$1 ( \47854 , \47850 , \47853 );
not \g133764/U$3 ( \47855 , \47854 );
xor \g134035/U$1 ( \47856 , \40107 , \40110 );
xor \g134035/U$1_r1 ( \47857 , \47856 , \40119 );
not \g133764/U$4 ( \47858 , \47857 );
and \g133764/U$2 ( \47859 , \47855 , \47858 );
and \g133764/U$5 ( \47860 , \47854 , \47857 );
nor \g133764/U$1 ( \47861 , \47859 , \47860 );
xor \g456235/U$4 ( \47862 , \40256 , \40260 );
and \g456235/U$3 ( \47863 , \47862 , \40265 );
and \g456235/U$5 ( \47864 , \40256 , \40260 );
nor \g456235/U$2 ( \47865 , \47863 , \47864 );
xnor \g133529/U$1 ( \47866 , \47861 , \47865 );
or \g129661/U$2 ( \47867 , \47845 , \47866 );
or \g129661/U$3 ( \47868 , \47861 , \47865 );
nand \g129661/U$1 ( \47869 , \47867 , \47868 );
not \g133825/U$3 ( \47870 , \40069 );
not \g133865/U$3 ( \47871 , \40096 );
not \g133865/U$4 ( \47872 , \40122 );
or \g133865/U$2 ( \47873 , \47871 , \47872 );
or \g133865/U$5 ( \47874 , \40122 , \40096 );
nand \g133865/U$1 ( \47875 , \47873 , \47874 );
not \g133825/U$4 ( \47876 , \47875 );
or \g133825/U$2 ( \47877 , \47870 , \47876 );
or \g133825/U$5 ( \47878 , \47875 , \40069 );
nand \g133825/U$1 ( \47879 , \47877 , \47878 );
or \g133761/U$2 ( \47880 , \47852 , \40245 );
not \g133816/U$3 ( \47881 , \40245 );
not \g133816/U$4 ( \47882 , \47852 );
or \g133816/U$2 ( \47883 , \47881 , \47882 );
nand \g133816/U$1 ( \47884 , \47883 , \47857 );
nand \g133761/U$1 ( \47885 , \47880 , \47884 );
xor \g133638/U$1 ( \47886 , \47879 , \47885 );
and \g129555/U$2 ( \47887 , \47869 , \47886 );
and \g129555/U$3 ( \47888 , \47879 , \47885 );
nor \g129555/U$1 ( \47889 , \47887 , \47888 );
not \g129493/U$4 ( \47890 , \47889 );
or \g129493/U$2 ( \47891 , \40130 , \47890 );
or \g129493/U$5 ( \47892 , \47889 , \40129 );
nand \g129493/U$1 ( \47893 , \47891 , \47892 );
xor \g129455/U$1 ( \47894 , \40073 , \47893 );
nand \g129431/U$1 ( \47895 , \40061 , \47894 );
not \g128583/U$3 ( \47896 , \47895 );
xor \g132578/U$1 ( \47897 , \17412 , \9425 );
xor \g132578/U$1_r1 ( \47898 , \47897 , \40050 );
xor \g132520/U$1 ( \47899 , \17162 , \9169 );
xor \g132520/U$1_r1 ( \47900 , \47899 , \40053 );
and \g132464/U$2 ( \47901 , \47898 , \47900 );
not \g132464/U$4 ( \47902 , \47898 );
not \g132519/U$1 ( \47903 , \47900 );
and \g132464/U$3 ( \47904 , \47902 , \47903 );
nor \g132464/U$1 ( \47905 , \47901 , \47904 );
not \g135533/U$2 ( \47906 , \47905 );
xor \g132633/U$1 ( \47907 , \17661 , \9670 );
xor \g132633/U$1_r1 ( \47908 , \47907 , \40047 );
not \g132632/U$1 ( \47909 , \47908 );
and \g132535/U$2 ( \47910 , \47898 , \47909 );
not \g132535/U$4 ( \47911 , \47898 );
and \g132535/U$3 ( \47912 , \47911 , \47908 );
or \g132535/U$1 ( \47913 , \47910 , \47912 );
nor \g135533/U$1 ( \47914 , \47906 , \47913 );
nand \g129415/U$1 ( \47915 , \47914 , \47894 );
not \g129414/U$1 ( \47916 , \47915 );
xor \g132693/U$1 ( \47917 , \17908 , \9922 );
xor \g132693/U$1_r1 ( \47918 , \47917 , \40044 );
and \g132582/U$2 ( \47919 , \47918 , \47908 );
not \g132582/U$4 ( \47920 , \47918 );
and \g132582/U$3 ( \47921 , \47920 , \47909 );
nor \g132582/U$1 ( \47922 , \47919 , \47921 );
not \g135536/U$2 ( \47923 , \47922 );
xor \g132737/U$1 ( \47924 , \18157 , \10170 );
xor \g132737/U$1_r1 ( \47925 , \47924 , \40041 );
not \g132736/U$1 ( \47926 , \47925 );
and \g132637/U$2 ( \47927 , \47918 , \47926 );
not \g132637/U$4 ( \47928 , \47918 );
and \g132637/U$3 ( \47929 , \47928 , \47925 );
or \g132637/U$1 ( \47930 , \47927 , \47929 );
nor \g135536/U$1 ( \47931 , \47923 , \47930 );
nand \g129417/U$1 ( \47932 , \47931 , \47894 );
not \g129364/U$3 ( \47933 , \47932 );
nand \g132669/U$1 ( \47934 , \47925 , \47918 );
and \g132591/U$1 ( \47935 , \47908 , \47934 );
not \g129364/U$4 ( \47936 , \47935 );
and \g129364/U$2 ( \47937 , \47933 , \47936 );
and \g129364/U$5 ( \47938 , \47932 , \47935 );
nor \g129364/U$1 ( \47939 , \47937 , \47938 );
not \g129363/U$1 ( \47940 , \47939 );
not \g129135/U$3 ( \47941 , \47940 );
xor \g129949/U$1 ( \47942 , \47839 , \40415 );
not \g135512/U$2 ( \47943 , \47942 );
nor \g135512/U$1 ( \47944 , \47943 , \40060 );
xor \g132463/U$1 ( \47945 , \16912 , \8913 );
xor \g132463/U$1_r1 ( \47946 , \47945 , \40056 );
nand \g132438/U$1 ( \47947 , \47900 , \47946 );
and \g132319/U$1 ( \47948 , \40061 , \47947 );
not \g129671/U$3 ( \47949 , \47948 );
xor \g129859/U$1 ( \47950 , \40337 , \47841 );
and \g132348/U$2 ( \47951 , \47946 , \40061 );
not \g132348/U$4 ( \47952 , \47946 );
and \g132348/U$3 ( \47953 , \47952 , \40060 );
nor \g132348/U$1 ( \47954 , \47951 , \47953 );
not \g135531/U$2 ( \47955 , \47954 );
and \g132400/U$2 ( \47956 , \47946 , \47903 );
not \g132400/U$4 ( \47957 , \47946 );
and \g132400/U$3 ( \47958 , \47957 , \47900 );
or \g132400/U$1 ( \47959 , \47956 , \47958 );
nor \g135531/U$1 ( \47960 , \47955 , \47959 );
and \g129706/U$2 ( \47961 , \47950 , \47960 );
xor \g129768/U$1 ( \47962 , \47843 , \40268 );
and \g129706/U$3 ( \47963 , \47959 , \47962 );
nor \g129706/U$1 ( \47964 , \47961 , \47963 );
not \g129671/U$4 ( \47965 , \47964 );
or \g129671/U$2 ( \47966 , \47949 , \47965 );
or \g129671/U$5 ( \47967 , \47964 , \47948 );
nand \g129671/U$1 ( \47968 , \47966 , \47967 );
xor \g456000/U$1 ( \47969 , \47944 , \47968 );
xor \g129692/U$1 ( \47970 , \47866 , \47845 );
and \g129506/U$2 ( \47971 , \47970 , \47914 );
xor \g129592/U$1 ( \47972 , \47869 , \47886 );
and \g129506/U$3 ( \47973 , \47913 , \47972 );
nor \g129506/U$1 ( \47974 , \47971 , \47973 );
nand \g132560/U$1 ( \47975 , \47908 , \47898 );
and \g132470/U$1 ( \47976 , \47900 , \47975 );
not \g132469/U$1 ( \47977 , \47976 );
and \g129463/U$2 ( \47978 , \47974 , \47977 );
not \g129463/U$4 ( \47979 , \47974 );
and \g129463/U$3 ( \47980 , \47979 , \47976 );
nor \g129463/U$1 ( \47981 , \47978 , \47980 );
xor \g456000/U$1_r1 ( \47982 , \47969 , \47981 );
not \g129169/U$3 ( \47983 , \47982 );
and \g129789/U$2 ( \47984 , \47950 , \47959 );
and \g129789/U$3 ( \47985 , \47960 , \47942 );
nor \g129789/U$1 ( \47986 , \47984 , \47985 );
not \g129743/U$3 ( \47987 , \47986 );
not \g129743/U$4 ( \47988 , \47948 );
and \g129743/U$2 ( \47989 , \47987 , \47988 );
and \g129743/U$5 ( \47990 , \47986 , \47948 );
nor \g129743/U$1 ( \47991 , \47989 , \47990 );
xor \g132835/U$1 ( \47992 , \18659 , \10670 );
xor \g132835/U$1_r1 ( \47993 , \47992 , \40035 );
xor \g132792/U$1 ( \47994 , \18405 , \10422 );
xor \g132792/U$1_r1 ( \47995 , \47994 , \40038 );
nand \g132771/U$1 ( \47996 , \47993 , \47995 );
and \g132701/U$1 ( \47997 , \47925 , \47996 );
xor \g129248/U$4 ( \47998 , \47991 , \47997 );
and \g129389/U$2 ( \47999 , \47894 , \47930 );
and \g129389/U$3 ( \48000 , \47931 , \47972 );
nor \g129389/U$1 ( \48001 , \47999 , \48000 );
not \g129331/U$3 ( \48002 , \48001 );
not \g129331/U$4 ( \48003 , \47935 );
and \g129331/U$2 ( \48004 , \48002 , \48003 );
and \g129331/U$5 ( \48005 , \48001 , \47935 );
nor \g129331/U$1 ( \48006 , \48004 , \48005 );
and \g129248/U$3 ( \48007 , \47998 , \48006 );
and \g129248/U$5 ( \48008 , \47991 , \47997 );
or \g129248/U$2 ( \48009 , \48007 , \48008 );
not \g129169/U$4 ( \48010 , \48009 );
or \g129169/U$2 ( \48011 , \47983 , \48010 );
or \g129169/U$5 ( \48012 , \48009 , \47982 );
nand \g129169/U$1 ( \48013 , \48011 , \48012 );
not \g129135/U$4 ( \48014 , \48013 );
or \g129135/U$2 ( \48015 , \47941 , \48014 );
or \g129135/U$5 ( \48016 , \48013 , \47940 );
nand \g129135/U$1 ( \48017 , \48015 , \48016 );
xor \g130041/U$1 ( \48018 , \47837 , \47836 );
and \g129872/U$2 ( \48019 , \48018 , \47960 );
and \g129872/U$3 ( \48020 , \47959 , \47942 );
nor \g129872/U$1 ( \48021 , \48019 , \48020 );
not \g129835/U$3 ( \48022 , \48021 );
not \g129835/U$4 ( \48023 , \47948 );
and \g129835/U$2 ( \48024 , \48022 , \48023 );
and \g129835/U$5 ( \48025 , \48021 , \47948 );
nor \g129835/U$1 ( \48026 , \48024 , \48025 );
nand \g129997/U$1 ( \48027 , \40061 , \48018 );
or \g129530/U$2 ( \48028 , \48026 , \48027 );
and \g129547/U$2 ( \48029 , \48026 , \48027 );
and \g129614/U$2 ( \48030 , \47970 , \47913 );
and \g129614/U$3 ( \48031 , \47914 , \47962 );
nor \g129614/U$1 ( \48032 , \48030 , \48031 );
and \g129569/U$2 ( \48033 , \48032 , \47976 );
not \g129569/U$4 ( \48034 , \48032 );
and \g129569/U$3 ( \48035 , \48034 , \47977 );
nor \g129569/U$1 ( \48036 , \48033 , \48035 );
nor \g129547/U$1 ( \48037 , \48029 , \48036 );
not \g129546/U$1 ( \48038 , \48037 );
nand \g129530/U$1 ( \48039 , \48028 , \48038 );
and \g129046/U$2 ( \48040 , \48017 , \48039 );
not \g129066/U$3 ( \48041 , \48017 );
not \g129066/U$4 ( \48042 , \48039 );
and \g129066/U$2 ( \48043 , \48041 , \48042 );
and \g129705/U$2 ( \48044 , \47950 , \47914 );
and \g129705/U$3 ( \48045 , \47913 , \47962 );
nor \g129705/U$1 ( \48046 , \48044 , \48045 );
and \g129670/U$2 ( \48047 , \48046 , \47976 );
not \g129670/U$4 ( \48048 , \48046 );
and \g129670/U$3 ( \48049 , \48048 , \47977 );
nor \g129670/U$1 ( \48050 , \48047 , \48049 );
xor \g130131/U$1 ( \48051 , \40653 , \47834 );
nand \g130094/U$1 ( \48052 , \40061 , \48051 );
xor \g129282/U$4 ( \48053 , \48050 , \48052 );
and \g132695/U$2 ( \48054 , \47995 , \47925 );
not \g132695/U$4 ( \48055 , \47995 );
and \g132695/U$3 ( \48056 , \48055 , \47926 );
nor \g132695/U$1 ( \48057 , \48054 , \48056 );
not \g135538/U$2 ( \48058 , \48057 );
not \g132834/U$1 ( \48059 , \47993 );
and \g132750/U$2 ( \48060 , \47995 , \48059 );
not \g132750/U$4 ( \48061 , \47995 );
and \g132750/U$3 ( \48062 , \48061 , \47993 );
or \g132750/U$1 ( \48063 , \48060 , \48062 );
nor \g135538/U$1 ( \48064 , \48058 , \48063 );
nand \g129416/U$1 ( \48065 , \48064 , \47894 );
not \g129362/U$3 ( \48066 , \48065 );
not \g129362/U$4 ( \48067 , \47997 );
and \g129362/U$2 ( \48068 , \48066 , \48067 );
and \g129362/U$5 ( \48069 , \48065 , \47997 );
nor \g129362/U$1 ( \48070 , \48068 , \48069 );
and \g129282/U$3 ( \48071 , \48053 , \48070 );
and \g129282/U$5 ( \48072 , \48050 , \48052 );
or \g129282/U$2 ( \48073 , \48071 , \48072 );
not \g129536/U$3 ( \48074 , \48036 );
and \g129785/U$2 ( \48075 , \48027 , \48026 );
not \g129785/U$4 ( \48076 , \48027 );
not \g129834/U$1 ( \48077 , \48026 );
and \g129785/U$3 ( \48078 , \48076 , \48077 );
nor \g129785/U$1 ( \48079 , \48075 , \48078 );
not \g129536/U$4 ( \48080 , \48079 );
and \g129536/U$2 ( \48081 , \48074 , \48080 );
and \g129536/U$5 ( \48082 , \48036 , \48079 );
nor \g129536/U$1 ( \48083 , \48081 , \48082 );
xor \g129115/U$4 ( \48084 , \48073 , \48083 );
xor \g129248/U$1 ( \48085 , \47991 , \47997 );
xor \g129248/U$1_r1 ( \48086 , \48085 , \48006 );
and \g129115/U$3 ( \48087 , \48084 , \48086 );
and \g129115/U$5 ( \48088 , \48073 , \48083 );
or \g129115/U$2 ( \48089 , \48087 , \48088 );
nor \g129066/U$1 ( \48090 , \48043 , \48089 );
nor \g129046/U$1 ( \48091 , \48040 , \48090 );
not \g129037/U$3 ( \48092 , \48039 );
not \g129071/U$3 ( \48093 , \48017 );
not \g129071/U$4 ( \48094 , \48089 );
and \g129071/U$2 ( \48095 , \48093 , \48094 );
and \g129071/U$5 ( \48096 , \48089 , \48017 );
nor \g129071/U$1 ( \48097 , \48095 , \48096 );
not \g129037/U$4 ( \48098 , \48097 );
or \g129037/U$2 ( \48099 , \48092 , \48098 );
or \g129037/U$5 ( \48100 , \48097 , \48039 );
nand \g129037/U$1 ( \48101 , \48099 , \48100 );
and \g129874/U$2 ( \48102 , \48018 , \47914 );
and \g129874/U$3 ( \48103 , \47913 , \47942 );
nor \g129874/U$1 ( \48104 , \48102 , \48103 );
and \g129838/U$2 ( \48105 , \48104 , \47976 );
not \g129838/U$4 ( \48106 , \48104 );
and \g129838/U$3 ( \48107 , \48106 , \47977 );
nor \g129838/U$1 ( \48108 , \48105 , \48107 );
and \g129967/U$2 ( \48109 , \48051 , \47960 );
and \g129967/U$3 ( \48110 , \47959 , \48018 );
nor \g129967/U$1 ( \48111 , \48109 , \48110 );
not \g129924/U$3 ( \48112 , \48111 );
not \g129924/U$4 ( \48113 , \47948 );
and \g129924/U$2 ( \48114 , \48112 , \48113 );
and \g129924/U$5 ( \48115 , \48111 , \47948 );
nor \g129924/U$1 ( \48116 , \48114 , \48115 );
xor \g130213/U$1 ( \48117 , \47832 , \47831 );
nand \g130172/U$1 ( \48118 , \40061 , \48117 );
xor \g455987/U$9 ( \48119 , \48116 , \48118 );
and \g129615/U$2 ( \48120 , \47970 , \47930 );
and \g129615/U$3 ( \48121 , \47931 , \47962 );
nor \g129615/U$1 ( \48122 , \48120 , \48121 );
not \g129570/U$3 ( \48123 , \48122 );
not \g129570/U$4 ( \48124 , \47935 );
and \g129570/U$2 ( \48125 , \48123 , \48124 );
and \g129570/U$5 ( \48126 , \48122 , \47935 );
nor \g129570/U$1 ( \48127 , \48125 , \48126 );
xor \g455987/U$9_r1 ( \48128 , \48119 , \48127 );
and \g455987/U$8 ( \48129 , \48108 , \48128 );
and \g130062/U$2 ( \48130 , \48051 , \47959 );
and \g130062/U$3 ( \48131 , \47960 , \48117 );
nor \g130062/U$1 ( \48132 , \48130 , \48131 );
not \g130020/U$3 ( \48133 , \48132 );
not \g130020/U$4 ( \48134 , \47948 );
and \g130020/U$2 ( \48135 , \48133 , \48134 );
and \g130020/U$5 ( \48136 , \48132 , \47948 );
nor \g130020/U$1 ( \48137 , \48135 , \48136 );
xor \g130285/U$1 ( \48138 , \47829 , \40839 );
nand \g130251/U$1 ( \48139 , \40061 , \48138 );
xor \g129272/U$4 ( \48140 , \48137 , \48139 );
xor \g132885/U$1 ( \48141 , \18910 , \10912 );
xor \g132885/U$1_r1 ( \48142 , \48141 , \40032 );
and \g132793/U$2 ( \48143 , \48142 , \47993 );
not \g132793/U$4 ( \48144 , \48142 );
and \g132793/U$3 ( \48145 , \48144 , \48059 );
nor \g132793/U$1 ( \48146 , \48143 , \48145 );
not \g135540/U$2 ( \48147 , \48146 );
xor \g132923/U$1 ( \48148 , \19156 , \11157 );
xor \g132923/U$1_r1 ( \48149 , \48148 , \40029 );
not \g132922/U$1 ( \48150 , \48149 );
and \g132836/U$2 ( \48151 , \48142 , \48150 );
not \g132836/U$4 ( \48152 , \48142 );
and \g132836/U$3 ( \48153 , \48152 , \48149 );
or \g132836/U$1 ( \48154 , \48151 , \48153 );
nor \g135540/U$1 ( \48155 , \48147 , \48154 );
nand \g129419/U$1 ( \48156 , \48155 , \47894 );
not \g129367/U$3 ( \48157 , \48156 );
nand \g132867/U$1 ( \48158 , \48149 , \48142 );
and \g132800/U$1 ( \48159 , \47993 , \48158 );
not \g129367/U$4 ( \48160 , \48159 );
and \g129367/U$2 ( \48161 , \48157 , \48160 );
and \g129367/U$5 ( \48162 , \48156 , \48159 );
nor \g129367/U$1 ( \48163 , \48161 , \48162 );
and \g129272/U$3 ( \48164 , \48140 , \48163 );
and \g129272/U$5 ( \48165 , \48137 , \48139 );
or \g129272/U$2 ( \48166 , \48164 , \48165 );
xor \g455987/U$11 ( \48167 , \48116 , \48118 );
xor \g455987/U$11_r1 ( \48168 , \48167 , \48127 );
and \g455987/U$10 ( \48169 , \48166 , \48168 );
and \g455987/U$12 ( \48170 , \48108 , \48166 );
or \g455987/U$7 ( \48171 , \48129 , \48169 , \48170 );
not \g128936/U$3 ( \48172 , \48171 );
not \g129465/U$3 ( \48173 , \47997 );
and \g129508/U$2 ( \48174 , \47970 , \48064 );
and \g129508/U$3 ( \48175 , \48063 , \47972 );
nor \g129508/U$1 ( \48176 , \48174 , \48175 );
not \g129465/U$4 ( \48177 , \48176 );
or \g129465/U$2 ( \48178 , \48173 , \48177 );
or \g129465/U$5 ( \48179 , \48176 , \47997 );
nand \g129465/U$1 ( \48180 , \48178 , \48179 );
not \g129673/U$3 ( \48181 , \47935 );
and \g129708/U$2 ( \48182 , \47950 , \47931 );
and \g129708/U$3 ( \48183 , \47930 , \47962 );
nor \g129708/U$1 ( \48184 , \48182 , \48183 );
not \g129673/U$4 ( \48185 , \48184 );
or \g129673/U$2 ( \48186 , \48181 , \48185 );
or \g129673/U$5 ( \48187 , \48184 , \47935 );
nand \g129673/U$1 ( \48188 , \48186 , \48187 );
not \g129650/U$2 ( \48189 , \48188 );
not \g129837/U$1 ( \48190 , \48108 );
nand \g129650/U$1 ( \48191 , \48189 , \48190 );
and \g129438/U$2 ( \48192 , \48180 , \48191 );
and \g129438/U$3 ( \48193 , \48108 , \48188 );
nor \g129438/U$1 ( \48194 , \48192 , \48193 );
and \g129790/U$2 ( \48195 , \47950 , \47913 );
and \g129790/U$3 ( \48196 , \47914 , \47942 );
nor \g129790/U$1 ( \48197 , \48195 , \48196 );
and \g129744/U$2 ( \48198 , \48197 , \47976 );
not \g129744/U$4 ( \48199 , \48197 );
and \g129744/U$3 ( \48200 , \48199 , \47977 );
nor \g129744/U$1 ( \48201 , \48198 , \48200 );
xor \g455985/U$9 ( \48202 , \48201 , \48159 );
and \g129390/U$2 ( \48203 , \47894 , \48063 );
and \g129390/U$3 ( \48204 , \48064 , \47972 );
nor \g129390/U$1 ( \48205 , \48203 , \48204 );
not \g129332/U$3 ( \48206 , \48205 );
not \g129332/U$4 ( \48207 , \47997 );
and \g129332/U$2 ( \48208 , \48206 , \48207 );
and \g129332/U$5 ( \48209 , \48205 , \47997 );
nor \g129332/U$1 ( \48210 , \48208 , \48209 );
xor \g455985/U$9_r1 ( \48211 , \48202 , \48210 );
and \g455985/U$8 ( \48212 , \48194 , \48211 );
xor \g455987/U$2 ( \48213 , \48116 , \48118 );
xor \g455987/U$1 ( \48214 , \48213 , \48127 );
xor \g455987/U$1_r1 ( \48215 , \48108 , \48166 );
xor \g455987/U$1_r2 ( \48216 , \48214 , \48215 );
xor \g455985/U$11 ( \48217 , \48201 , \48159 );
xor \g455985/U$11_r1 ( \48218 , \48217 , \48210 );
and \g455985/U$10 ( \48219 , \48216 , \48218 );
and \g455985/U$12 ( \48220 , \48194 , \48216 );
or \g455985/U$7 ( \48221 , \48212 , \48219 , \48220 );
xor \g129282/U$1 ( \48222 , \48050 , \48052 );
xor \g129282/U$1_r1 ( \48223 , \48222 , \48070 );
not \g129072/U$3 ( \48224 , \48223 );
and \g129507/U$2 ( \48225 , \47970 , \47931 );
and \g129507/U$3 ( \48226 , \47930 , \47972 );
nor \g129507/U$1 ( \48227 , \48225 , \48226 );
not \g129464/U$3 ( \48228 , \48227 );
not \g129464/U$4 ( \48229 , \47935 );
and \g129464/U$2 ( \48230 , \48228 , \48229 );
and \g129464/U$5 ( \48231 , \48227 , \47935 );
nor \g129464/U$1 ( \48232 , \48230 , \48231 );
not \g129136/U$3 ( \48233 , \48232 );
not \g129170/U$3 ( \48234 , \48026 );
xor \g455985/U$5 ( \48235 , \48201 , \48159 );
and \g455985/U$4 ( \48236 , \48235 , \48210 );
and \g455985/U$6 ( \48237 , \48201 , \48159 );
or \g455985/U$3 ( \48238 , \48236 , \48237 );
not \g129170/U$4 ( \48239 , \48238 );
or \g129170/U$2 ( \48240 , \48234 , \48239 );
or \g129170/U$5 ( \48241 , \48238 , \48026 );
nand \g129170/U$1 ( \48242 , \48240 , \48241 );
not \g129136/U$4 ( \48243 , \48242 );
or \g129136/U$2 ( \48244 , \48233 , \48243 );
or \g129136/U$5 ( \48245 , \48242 , \48232 );
nand \g129136/U$1 ( \48246 , \48244 , \48245 );
not \g129072/U$4 ( \48247 , \48246 );
or \g129072/U$2 ( \48248 , \48224 , \48247 );
or \g129072/U$5 ( \48249 , \48246 , \48223 );
nand \g129072/U$1 ( \48250 , \48248 , \48249 );
not \g129030/U$3 ( \48251 , \48250 );
xor \g455987/U$5 ( \48252 , \48116 , \48118 );
and \g455987/U$4 ( \48253 , \48252 , \48127 );
and \g455987/U$6 ( \48254 , \48116 , \48118 );
or \g455987/U$3 ( \48255 , \48253 , \48254 );
not \g129030/U$4 ( \48256 , \48255 );
and \g129030/U$2 ( \48257 , \48251 , \48256 );
and \g129030/U$5 ( \48258 , \48250 , \48255 );
nor \g129030/U$1 ( \48259 , \48257 , \48258 );
xor \g455931/U$1 ( \48260 , \48221 , \48259 );
not \g128936/U$4 ( \48261 , \48260 );
or \g128936/U$2 ( \48262 , \48172 , \48261 );
or \g128936/U$5 ( \48263 , \48260 , \48171 );
nand \g128936/U$1 ( \48264 , \48262 , \48263 );
xor \g455985/U$2 ( \48265 , \48201 , \48159 );
xor \g455985/U$1 ( \48266 , \48265 , \48210 );
xor \g455985/U$1_r1 ( \48267 , \48194 , \48216 );
xor \g455985/U$1_r2 ( \48268 , \48266 , \48267 );
not \g128978/U$3 ( \48269 , \48268 );
and \g129612/U$2 ( \48270 , \48188 , \48190 );
nor \g129649/U$1 ( \48271 , \48188 , \48190 );
nor \g129612/U$1 ( \48272 , \48270 , \48271 );
not \g129444/U$3 ( \48273 , \48272 );
not \g129444/U$4 ( \48274 , \48180 );
or \g129444/U$2 ( \48275 , \48273 , \48274 );
or \g129444/U$5 ( \48276 , \48180 , \48272 );
nand \g129444/U$1 ( \48277 , \48275 , \48276 );
not \g129087/U$3 ( \48278 , \48277 );
and \g129616/U$2 ( \48279 , \47970 , \48063 );
and \g129616/U$3 ( \48280 , \48064 , \47962 );
nor \g129616/U$1 ( \48281 , \48279 , \48280 );
not \g129571/U$3 ( \48282 , \48281 );
not \g129571/U$4 ( \48283 , \47997 );
and \g129571/U$2 ( \48284 , \48282 , \48283 );
and \g129571/U$5 ( \48285 , \48281 , \47997 );
nor \g129571/U$1 ( \48286 , \48284 , \48285 );
and \g130061/U$2 ( \48287 , \48051 , \47913 );
and \g130061/U$3 ( \48288 , \47914 , \48117 );
nor \g130061/U$1 ( \48289 , \48287 , \48288 );
and \g130019/U$2 ( \48290 , \48289 , \47977 );
not \g130019/U$4 ( \48291 , \48289 );
and \g130019/U$3 ( \48292 , \48291 , \47976 );
nor \g130019/U$1 ( \48293 , \48290 , \48292 );
not \g129836/U$3 ( \48294 , \47935 );
and \g129873/U$2 ( \48295 , \48018 , \47931 );
and \g129873/U$3 ( \48296 , \47930 , \47942 );
nor \g129873/U$1 ( \48297 , \48295 , \48296 );
not \g129836/U$4 ( \48298 , \48297 );
or \g129836/U$2 ( \48299 , \48294 , \48298 );
or \g129836/U$5 ( \48300 , \48297 , \47935 );
nand \g129836/U$1 ( \48301 , \48299 , \48300 );
xor \g456018/U$4 ( \48302 , \48293 , \48301 );
not \g129672/U$3 ( \48303 , \47997 );
and \g129707/U$2 ( \48304 , \47950 , \48064 );
and \g129707/U$3 ( \48305 , \48063 , \47962 );
nor \g129707/U$1 ( \48306 , \48304 , \48305 );
not \g129672/U$4 ( \48307 , \48306 );
or \g129672/U$2 ( \48308 , \48303 , \48307 );
or \g129672/U$5 ( \48309 , \48306 , \47997 );
nand \g129672/U$1 ( \48310 , \48308 , \48309 );
and \g456018/U$3 ( \48311 , \48302 , \48310 );
and \g456018/U$5 ( \48312 , \48293 , \48301 );
nor \g456018/U$2 ( \48313 , \48311 , \48312 );
or \g129317/U$2 ( \48314 , \48286 , \48313 );
not \g129324/U$3 ( \48315 , \48313 );
not \g129324/U$4 ( \48316 , \48286 );
or \g129324/U$2 ( \48317 , \48315 , \48316 );
xor \g133005/U$1 ( \48318 , \19652 , \11649 );
xor \g133005/U$1_r1 ( \48319 , \48318 , \40023 );
xor \g132971/U$1 ( \48320 , \19406 , \11400 );
xor \g132971/U$1_r1 ( \48321 , \48320 , \40026 );
nand \g132956/U$1 ( \48322 , \48319 , \48321 );
and \g132893/U$1 ( \48323 , \48149 , \48322 );
not \g129366/U$3 ( \48324 , \48323 );
and \g132886/U$2 ( \48325 , \48321 , \48149 );
not \g132886/U$4 ( \48326 , \48321 );
and \g132886/U$3 ( \48327 , \48326 , \48150 );
nor \g132886/U$1 ( \48328 , \48325 , \48327 );
not \g135541/U$2 ( \48329 , \48328 );
not \g133004/U$1 ( \48330 , \48319 );
and \g132937/U$2 ( \48331 , \48321 , \48330 );
not \g132937/U$4 ( \48332 , \48321 );
and \g132937/U$3 ( \48333 , \48332 , \48319 );
or \g132937/U$1 ( \48334 , \48331 , \48333 );
nor \g135541/U$1 ( \48335 , \48329 , \48334 );
nand \g129418/U$1 ( \48336 , \48335 , \47894 );
not \g129366/U$4 ( \48337 , \48336 );
or \g129366/U$2 ( \48338 , \48324 , \48337 );
or \g129366/U$5 ( \48339 , \48336 , \48323 );
nand \g129366/U$1 ( \48340 , \48338 , \48339 );
nand \g129324/U$1 ( \48341 , \48317 , \48340 );
nand \g129317/U$1 ( \48342 , \48314 , \48341 );
not \g129087/U$4 ( \48343 , \48342 );
or \g129087/U$2 ( \48344 , \48278 , \48343 );
or \g129098/U$2 ( \48345 , \48342 , \48277 );
and \g130426/U$2 ( \48346 , \41069 , \47823 );
not \g130426/U$4 ( \48347 , \41069 );
and \g130426/U$3 ( \48348 , \48347 , \47824 );
or \g130426/U$1 ( \48349 , \48346 , \48348 );
not \g135513/U$2 ( \48350 , \48349 );
nor \g135513/U$1 ( \48351 , \48350 , \40060 );
not \g130189/U$3 ( \48352 , \47948 );
xor \g130355/U$1 ( \48353 , \47827 , \47826 );
and \g130228/U$2 ( \48354 , \48353 , \47960 );
and \g130228/U$3 ( \48355 , \47959 , \48138 );
nor \g130228/U$1 ( \48356 , \48354 , \48355 );
not \g130189/U$4 ( \48357 , \48356 );
or \g130189/U$2 ( \48358 , \48352 , \48357 );
or \g130189/U$5 ( \48359 , \48356 , \47948 );
nand \g130189/U$1 ( \48360 , \48358 , \48359 );
xor \g456001/U$4 ( \48361 , \48351 , \48360 );
not \g129466/U$3 ( \48362 , \48159 );
and \g129509/U$2 ( \48363 , \47970 , \48155 );
and \g129509/U$3 ( \48364 , \48154 , \47972 );
nor \g129509/U$1 ( \48365 , \48363 , \48364 );
not \g129466/U$4 ( \48366 , \48365 );
or \g129466/U$2 ( \48367 , \48362 , \48366 );
or \g129466/U$5 ( \48368 , \48365 , \48159 );
nand \g129466/U$1 ( \48369 , \48367 , \48368 );
and \g456001/U$3 ( \48370 , \48361 , \48369 );
and \g456001/U$5 ( \48371 , \48351 , \48360 );
nor \g456001/U$2 ( \48372 , \48370 , \48371 );
and \g130148/U$2 ( \48373 , \48117 , \47959 );
and \g130148/U$3 ( \48374 , \47960 , \48138 );
nor \g130148/U$1 ( \48375 , \48373 , \48374 );
not \g130110/U$3 ( \48376 , \48375 );
not \g130110/U$4 ( \48377 , \47948 );
and \g130110/U$2 ( \48378 , \48376 , \48377 );
and \g130110/U$5 ( \48379 , \48375 , \47948 );
nor \g130110/U$1 ( \48380 , \48378 , \48379 );
nand \g130316/U$1 ( \48381 , \40061 , \48353 );
xor \g129861/U$1 ( \48382 , \48380 , \48381 );
and \g129968/U$2 ( \48383 , \48051 , \47914 );
and \g129968/U$3 ( \48384 , \47913 , \48018 );
nor \g129968/U$1 ( \48385 , \48383 , \48384 );
and \g129925/U$2 ( \48386 , \48385 , \47976 );
not \g129925/U$4 ( \48387 , \48385 );
and \g129925/U$3 ( \48388 , \48387 , \47977 );
nor \g129925/U$1 ( \48389 , \48386 , \48388 );
xor \g129861/U$1_r1 ( \48390 , \48382 , \48389 );
xor \g129114/U$4 ( \48391 , \48372 , \48390 );
and \g129791/U$2 ( \48392 , \47950 , \47930 );
and \g129791/U$3 ( \48393 , \47931 , \47942 );
nor \g129791/U$1 ( \48394 , \48392 , \48393 );
not \g129745/U$3 ( \48395 , \48394 );
not \g129745/U$4 ( \48396 , \47935 );
and \g129745/U$2 ( \48397 , \48395 , \48396 );
and \g129745/U$5 ( \48398 , \48394 , \47935 );
nor \g129745/U$1 ( \48399 , \48397 , \48398 );
xor \g129249/U$1 ( \48400 , \48399 , \48323 );
and \g129391/U$2 ( \48401 , \47894 , \48154 );
and \g129391/U$3 ( \48402 , \48155 , \47972 );
nor \g129391/U$1 ( \48403 , \48401 , \48402 );
not \g129333/U$3 ( \48404 , \48403 );
not \g129333/U$4 ( \48405 , \48159 );
and \g129333/U$2 ( \48406 , \48404 , \48405 );
and \g129333/U$5 ( \48407 , \48403 , \48159 );
nor \g129333/U$1 ( \48408 , \48406 , \48407 );
xor \g129249/U$1_r1 ( \48409 , \48400 , \48408 );
and \g129114/U$3 ( \48410 , \48391 , \48409 );
and \g129114/U$5 ( \48411 , \48372 , \48390 );
or \g129114/U$2 ( \48412 , \48410 , \48411 );
not \g129113/U$1 ( \48413 , \48412 );
nand \g129098/U$1 ( \48414 , \48345 , \48413 );
nand \g129087/U$1 ( \48415 , \48344 , \48414 );
not \g128978/U$4 ( \48416 , \48415 );
or \g128978/U$2 ( \48417 , \48269 , \48416 );
or \g128978/U$5 ( \48418 , \48415 , \48268 );
nand \g128978/U$1 ( \48419 , \48417 , \48418 );
not \g128947/U$3 ( \48420 , \48419 );
xor \g129249/U$4 ( \48421 , \48399 , \48323 );
and \g129249/U$3 ( \48422 , \48421 , \48408 );
and \g129249/U$5 ( \48423 , \48399 , \48323 );
or \g129249/U$2 ( \48424 , \48422 , \48423 );
xor \g129861/U$4 ( \48425 , \48380 , \48381 );
and \g129861/U$3 ( \48426 , \48425 , \48389 );
and \g129861/U$5 ( \48427 , \48380 , \48381 );
or \g129861/U$2 ( \48428 , \48426 , \48427 );
xor \g129116/U$4 ( \48429 , \48424 , \48428 );
xor \g129272/U$1 ( \48430 , \48137 , \48139 );
xor \g129272/U$1_r1 ( \48431 , \48430 , \48163 );
and \g129116/U$3 ( \48432 , \48429 , \48431 );
and \g129116/U$5 ( \48433 , \48424 , \48428 );
or \g129116/U$2 ( \48434 , \48432 , \48433 );
not \g128947/U$4 ( \48435 , \48434 );
and \g128947/U$2 ( \48436 , \48420 , \48435 );
and \g128947/U$5 ( \48437 , \48419 , \48434 );
nor \g128947/U$1 ( \48438 , \48436 , \48437 );
xor \g456018/U$1 ( \48439 , \48293 , \48301 );
xor \g456018/U$1_r1 ( \48440 , \48439 , \48310 );
xor \g456001/U$1 ( \48441 , \48351 , \48360 );
xor \g456001/U$1_r1 ( \48442 , \48441 , \48369 );
xor \g455996/U$4 ( \48443 , \48440 , \48442 );
and \g129617/U$2 ( \48444 , \47970 , \48154 );
and \g129617/U$3 ( \48445 , \48155 , \47962 );
nor \g129617/U$1 ( \48446 , \48444 , \48445 );
not \g129572/U$3 ( \48447 , \48446 );
not \g129572/U$4 ( \48448 , \48159 );
and \g129572/U$2 ( \48449 , \48447 , \48448 );
and \g129572/U$5 ( \48450 , \48446 , \48159 );
nor \g129572/U$1 ( \48451 , \48449 , \48450 );
not \g130264/U$3 ( \48452 , \47948 );
and \g130298/U$2 ( \48453 , \48349 , \47960 );
and \g130298/U$3 ( \48454 , \47959 , \48353 );
nor \g130298/U$1 ( \48455 , \48453 , \48454 );
not \g130264/U$4 ( \48456 , \48455 );
or \g130264/U$2 ( \48457 , \48452 , \48456 );
or \g130264/U$5 ( \48458 , \48455 , \47948 );
nand \g130264/U$1 ( \48459 , \48457 , \48458 );
not \g130263/U$1 ( \48460 , \48459 );
or \g129318/U$2 ( \48461 , \48451 , \48460 );
not \g129325/U$3 ( \48462 , \48460 );
not \g129325/U$4 ( \48463 , \48451 );
or \g129325/U$2 ( \48464 , \48462 , \48463 );
xor \g133048/U$1 ( \48465 , \19894 , \11898 );
xor \g133048/U$1_r1 ( \48466 , \48465 , \40020 );
and \g132972/U$2 ( \48467 , \48466 , \48319 );
not \g132972/U$4 ( \48468 , \48466 );
and \g132972/U$3 ( \48469 , \48468 , \48330 );
nor \g132972/U$1 ( \48470 , \48467 , \48469 );
not \g135544/U$2 ( \48471 , \48470 );
xor \g133086/U$1 ( \48472 , \20139 , \12140 );
xor \g133086/U$1_r1 ( \48473 , \48472 , \40017 );
not \g133085/U$1 ( \48474 , \48473 );
and \g133007/U$2 ( \48475 , \48466 , \48474 );
not \g133007/U$4 ( \48476 , \48466 );
and \g133007/U$3 ( \48477 , \48476 , \48473 );
or \g133007/U$1 ( \48478 , \48475 , \48477 );
nor \g135544/U$1 ( \48479 , \48471 , \48478 );
nand \g129420/U$1 ( \48480 , \48479 , \47894 );
not \g129369/U$3 ( \48481 , \48480 );
nand \g133034/U$1 ( \48482 , \48473 , \48466 );
and \g132979/U$1 ( \48483 , \48319 , \48482 );
not \g129369/U$4 ( \48484 , \48483 );
and \g129369/U$2 ( \48485 , \48481 , \48484 );
and \g129369/U$5 ( \48486 , \48480 , \48483 );
nor \g129369/U$1 ( \48487 , \48485 , \48486 );
not \g129368/U$1 ( \48488 , \48487 );
nand \g129325/U$1 ( \48489 , \48464 , \48488 );
nand \g129318/U$1 ( \48490 , \48461 , \48489 );
and \g455996/U$3 ( \48491 , \48443 , \48490 );
and \g455996/U$5 ( \48492 , \48440 , \48442 );
nor \g455996/U$2 ( \48493 , \48491 , \48492 );
not \g129365/U$1 ( \48494 , \48340 );
and \g129309/U$2 ( \48495 , \48313 , \48494 );
not \g129309/U$4 ( \48496 , \48313 );
and \g129309/U$3 ( \48497 , \48496 , \48340 );
nor \g129309/U$1 ( \48498 , \48495 , \48497 );
not \g129292/U$3 ( \48499 , \48498 );
not \g129292/U$4 ( \48500 , \48286 );
and \g129292/U$2 ( \48501 , \48499 , \48500 );
and \g129292/U$5 ( \48502 , \48498 , \48286 );
nor \g129292/U$1 ( \48503 , \48501 , \48502 );
xor \g129018/U$1 ( \48504 , \48493 , \48503 );
and \g130149/U$2 ( \48505 , \48117 , \47913 );
and \g130149/U$3 ( \48506 , \47914 , \48138 );
nor \g130149/U$1 ( \48507 , \48505 , \48506 );
and \g130111/U$2 ( \48508 , \48507 , \47976 );
not \g130111/U$4 ( \48509 , \48507 );
and \g130111/U$3 ( \48510 , \48509 , \47977 );
nor \g130111/U$1 ( \48511 , \48508 , \48510 );
and \g130498/U$2 ( \48512 , \47820 , \47808 );
not \g130498/U$4 ( \48513 , \47820 );
and \g130498/U$3 ( \48514 , \48513 , \47809 );
or \g130498/U$1 ( \48515 , \48512 , \48514 );
nand \g130460/U$1 ( \48516 , \40061 , \48515 );
or \g129890/U$2 ( \48517 , \48511 , \48516 );
and \g129910/U$2 ( \48518 , \48511 , \48516 );
and \g129969/U$2 ( \48519 , \48051 , \47931 );
and \g129969/U$3 ( \48520 , \47930 , \48018 );
nor \g129969/U$1 ( \48521 , \48519 , \48520 );
not \g129926/U$3 ( \48522 , \48521 );
not \g129926/U$4 ( \48523 , \47935 );
and \g129926/U$2 ( \48524 , \48522 , \48523 );
and \g129926/U$5 ( \48525 , \48521 , \47935 );
nor \g129926/U$1 ( \48526 , \48524 , \48525 );
nor \g129910/U$1 ( \48527 , \48518 , \48526 );
not \g129909/U$1 ( \48528 , \48527 );
nand \g129890/U$1 ( \48529 , \48517 , \48528 );
and \g129185/U$2 ( \48530 , \48494 , \48529 );
not \g129205/U$3 ( \48531 , \48494 );
not \g129205/U$4 ( \48532 , \48529 );
and \g129205/U$2 ( \48533 , \48531 , \48532 );
and \g129792/U$2 ( \48534 , \47950 , \48063 );
and \g129792/U$3 ( \48535 , \48064 , \47942 );
nor \g129792/U$1 ( \48536 , \48534 , \48535 );
not \g129746/U$3 ( \48537 , \48536 );
not \g129746/U$4 ( \48538 , \47997 );
and \g129746/U$2 ( \48539 , \48537 , \48538 );
and \g129746/U$5 ( \48540 , \48536 , \47997 );
nor \g129746/U$1 ( \48541 , \48539 , \48540 );
xor \g129250/U$4 ( \48542 , \48541 , \48483 );
and \g129392/U$2 ( \48543 , \47894 , \48334 );
and \g129392/U$3 ( \48544 , \48335 , \47972 );
nor \g129392/U$1 ( \48545 , \48543 , \48544 );
not \g129334/U$3 ( \48546 , \48545 );
not \g129334/U$4 ( \48547 , \48323 );
and \g129334/U$2 ( \48548 , \48546 , \48547 );
and \g129334/U$5 ( \48549 , \48545 , \48323 );
nor \g129334/U$1 ( \48550 , \48548 , \48549 );
and \g129250/U$3 ( \48551 , \48542 , \48550 );
and \g129250/U$5 ( \48552 , \48541 , \48483 );
or \g129250/U$2 ( \48553 , \48551 , \48552 );
nor \g129205/U$1 ( \48554 , \48533 , \48553 );
nor \g129185/U$1 ( \48555 , \48530 , \48554 );
xor \g129018/U$1_r1 ( \48556 , \48504 , \48555 );
xor \g129114/U$1 ( \48557 , \48372 , \48390 );
xor \g129114/U$1_r1 ( \48558 , \48557 , \48409 );
or \g128955/U$2 ( \48559 , \48556 , \48558 );
not \g128964/U$3 ( \48560 , \48558 );
not \g128964/U$4 ( \48561 , \48556 );
or \g128964/U$2 ( \48562 , \48560 , \48561 );
xor \g129250/U$1 ( \48563 , \48541 , \48483 );
xor \g129250/U$1_r1 ( \48564 , \48563 , \48550 );
and \g130565/U$2 ( \48565 , \47805 , \47783 );
not \g130565/U$4 ( \48566 , \47805 );
and \g130565/U$3 ( \48567 , \48566 , \47784 );
or \g130565/U$1 ( \48568 , \48565 , \48567 );
not \g135514/U$2 ( \48569 , \48568 );
nor \g135514/U$1 ( \48570 , \48569 , \40060 );
not \g130021/U$3 ( \48571 , \47935 );
and \g130063/U$2 ( \48572 , \48051 , \47930 );
and \g130063/U$3 ( \48573 , \47931 , \48117 );
nor \g130063/U$1 ( \48574 , \48572 , \48573 );
not \g130021/U$4 ( \48575 , \48574 );
or \g130021/U$2 ( \48576 , \48571 , \48575 );
or \g130021/U$5 ( \48577 , \48574 , \47935 );
nand \g130021/U$1 ( \48578 , \48576 , \48577 );
xor \g456032/U$4 ( \48579 , \48570 , \48578 );
not \g129839/U$3 ( \48580 , \47997 );
and \g129875/U$2 ( \48581 , \48018 , \48064 );
and \g129875/U$3 ( \48582 , \48063 , \47942 );
nor \g129875/U$1 ( \48583 , \48581 , \48582 );
not \g129839/U$4 ( \48584 , \48583 );
or \g129839/U$2 ( \48585 , \48580 , \48584 );
or \g129839/U$5 ( \48586 , \48583 , \47997 );
nand \g129839/U$1 ( \48587 , \48585 , \48586 );
and \g456032/U$3 ( \48588 , \48579 , \48587 );
and \g456032/U$5 ( \48589 , \48570 , \48578 );
nor \g456032/U$2 ( \48590 , \48588 , \48589 );
not \g129562/U$2 ( \48591 , \48590 );
and \g130229/U$2 ( \48592 , \48353 , \47914 );
and \g130229/U$3 ( \48593 , \47913 , \48138 );
nor \g130229/U$1 ( \48594 , \48592 , \48593 );
and \g130190/U$2 ( \48595 , \48594 , \47976 );
not \g130190/U$4 ( \48596 , \48594 );
and \g130190/U$3 ( \48597 , \48596 , \47977 );
nor \g130190/U$1 ( \48598 , \48595 , \48597 );
and \g130372/U$2 ( \48599 , \48349 , \47959 );
and \g130372/U$3 ( \48600 , \47960 , \48515 );
nor \g130372/U$1 ( \48601 , \48599 , \48600 );
not \g130331/U$3 ( \48602 , \48601 );
not \g130331/U$4 ( \48603 , \47948 );
and \g130331/U$2 ( \48604 , \48602 , \48603 );
and \g130331/U$5 ( \48605 , \48601 , \47948 );
nor \g130331/U$1 ( \48606 , \48604 , \48605 );
or \g129633/U$2 ( \48607 , \48598 , \48606 );
and \g129653/U$2 ( \48608 , \48598 , \48606 );
and \g129709/U$2 ( \48609 , \47950 , \48155 );
and \g129709/U$3 ( \48610 , \48154 , \47962 );
nor \g129709/U$1 ( \48611 , \48609 , \48610 );
not \g129674/U$3 ( \48612 , \48611 );
not \g129674/U$4 ( \48613 , \48159 );
and \g129674/U$2 ( \48614 , \48612 , \48613 );
and \g129674/U$5 ( \48615 , \48611 , \48159 );
nor \g129674/U$1 ( \48616 , \48614 , \48615 );
nor \g129653/U$1 ( \48617 , \48608 , \48616 );
not \g129652/U$1 ( \48618 , \48617 );
nand \g129633/U$1 ( \48619 , \48607 , \48618 );
nor \g129562/U$1 ( \48620 , \48591 , \48619 );
or \g129186/U$2 ( \48621 , \48564 , \48620 );
not \g129563/U$2 ( \48622 , \48590 );
nand \g129563/U$1 ( \48623 , \48622 , \48619 );
nand \g129186/U$1 ( \48624 , \48621 , \48623 );
xor \g455996/U$1 ( \48625 , \48440 , \48442 );
xor \g455996/U$1_r1 ( \48626 , \48625 , \48490 );
xor \g129005/U$4 ( \48627 , \48624 , \48626 );
not \g129137/U$3 ( \48628 , \48340 );
not \g129171/U$3 ( \48629 , \48529 );
not \g129171/U$4 ( \48630 , \48553 );
or \g129171/U$2 ( \48631 , \48629 , \48630 );
or \g129171/U$5 ( \48632 , \48553 , \48529 );
nand \g129171/U$1 ( \48633 , \48631 , \48632 );
not \g129137/U$4 ( \48634 , \48633 );
or \g129137/U$2 ( \48635 , \48628 , \48634 );
or \g129137/U$5 ( \48636 , \48633 , \48340 );
nand \g129137/U$1 ( \48637 , \48635 , \48636 );
and \g129005/U$3 ( \48638 , \48627 , \48637 );
and \g129005/U$5 ( \48639 , \48624 , \48626 );
or \g129005/U$2 ( \48640 , \48638 , \48639 );
nand \g128964/U$1 ( \48641 , \48562 , \48640 );
nand \g128955/U$1 ( \48642 , \48559 , \48641 );
not \g129310/U$3 ( \48643 , \48459 );
not \g129310/U$4 ( \48644 , \48487 );
or \g129310/U$2 ( \48645 , \48643 , \48644 );
or \g129310/U$5 ( \48646 , \48487 , \48459 );
nand \g129310/U$1 ( \48647 , \48645 , \48646 );
not \g129293/U$3 ( \48648 , \48647 );
not \g129293/U$4 ( \48649 , \48451 );
and \g129293/U$2 ( \48650 , \48648 , \48649 );
and \g129293/U$5 ( \48651 , \48647 , \48451 );
nor \g129293/U$1 ( \48652 , \48650 , \48651 );
not \g129900/U$3 ( \48653 , \48526 );
xor \g130055/U$1 ( \48654 , \48516 , \48511 );
not \g129900/U$4 ( \48655 , \48654 );
and \g129900/U$2 ( \48656 , \48653 , \48655 );
and \g129900/U$5 ( \48657 , \48526 , \48654 );
nor \g129900/U$1 ( \48658 , \48656 , \48657 );
xor \g129007/U$4 ( \48659 , \48652 , \48658 );
not \g129467/U$3 ( \48660 , \48323 );
and \g129510/U$2 ( \48661 , \47970 , \48335 );
and \g129510/U$3 ( \48662 , \48334 , \47972 );
nor \g129510/U$1 ( \48663 , \48661 , \48662 );
not \g129467/U$4 ( \48664 , \48663 );
or \g129467/U$2 ( \48665 , \48660 , \48664 );
or \g129467/U$5 ( \48666 , \48663 , \48323 );
nand \g129467/U$1 ( \48667 , \48665 , \48666 );
and \g129181/U$2 ( \48668 , \48487 , \48667 );
not \g129201/U$3 ( \48669 , \48487 );
not \g129201/U$4 ( \48670 , \48667 );
and \g129201/U$2 ( \48671 , \48669 , \48670 );
and \g129793/U$2 ( \48672 , \47950 , \48154 );
and \g129793/U$3 ( \48673 , \48155 , \47942 );
nor \g129793/U$1 ( \48674 , \48672 , \48673 );
not \g129747/U$3 ( \48675 , \48674 );
not \g129747/U$4 ( \48676 , \48159 );
and \g129747/U$2 ( \48677 , \48675 , \48676 );
and \g129747/U$5 ( \48678 , \48674 , \48159 );
nor \g129747/U$1 ( \48679 , \48677 , \48678 );
xor \g133152/U$1 ( \48680 , \20628 , \12636 );
xor \g133152/U$1_r1 ( \48681 , \48680 , \40011 );
xor \g133124/U$1 ( \48682 , \20384 , \12391 );
xor \g133124/U$1_r1 ( \48683 , \48682 , \40014 );
nand \g133110/U$1 ( \48684 , \48681 , \48683 );
and \g133058/U$1 ( \48685 , \48473 , \48684 );
xor \g129251/U$4 ( \48686 , \48679 , \48685 );
and \g129393/U$2 ( \48687 , \47894 , \48478 );
and \g129393/U$3 ( \48688 , \48479 , \47972 );
nor \g129393/U$1 ( \48689 , \48687 , \48688 );
not \g129336/U$3 ( \48690 , \48689 );
not \g129336/U$4 ( \48691 , \48483 );
and \g129336/U$2 ( \48692 , \48690 , \48691 );
and \g129336/U$5 ( \48693 , \48689 , \48483 );
nor \g129336/U$1 ( \48694 , \48692 , \48693 );
and \g129251/U$3 ( \48695 , \48686 , \48694 );
and \g129251/U$5 ( \48696 , \48679 , \48685 );
or \g129251/U$2 ( \48697 , \48695 , \48696 );
nor \g129201/U$1 ( \48698 , \48671 , \48697 );
nor \g129181/U$1 ( \48699 , \48668 , \48698 );
and \g129007/U$3 ( \48700 , \48659 , \48699 );
and \g129007/U$5 ( \48701 , \48652 , \48658 );
or \g129007/U$2 ( \48702 , \48700 , \48701 );
not \g128872/U$3 ( \48703 , \48702 );
xor \g129005/U$1 ( \48704 , \48624 , \48626 );
xor \g129005/U$1_r1 ( \48705 , \48704 , \48637 );
not \g128897/U$3 ( \48706 , \48705 );
not \g129174/U$3 ( \48707 , \48619 );
not \g129174/U$4 ( \48708 , \48564 );
or \g129174/U$2 ( \48709 , \48707 , \48708 );
or \g129174/U$5 ( \48710 , \48564 , \48619 );
nand \g129174/U$1 ( \48711 , \48709 , \48710 );
not \g129139/U$3 ( \48712 , \48711 );
not \g129139/U$4 ( \48713 , \48590 );
and \g129139/U$2 ( \48714 , \48712 , \48713 );
and \g129139/U$5 ( \48715 , \48711 , \48590 );
nor \g129139/U$1 ( \48716 , \48714 , \48715 );
not \g129641/U$3 ( \48717 , \48616 );
xor \g130145/U$1 ( \48718 , \48606 , \48598 );
not \g129641/U$4 ( \48719 , \48718 );
and \g129641/U$2 ( \48720 , \48717 , \48719 );
and \g129641/U$5 ( \48721 , \48616 , \48718 );
nor \g129641/U$1 ( \48722 , \48720 , \48721 );
and \g130629/U$2 ( \48723 , \47780 , \47740 );
not \g130629/U$4 ( \48724 , \47780 );
and \g130629/U$3 ( \48725 , \48724 , \47741 );
or \g130629/U$1 ( \48726 , \48723 , \48725 );
not \g135515/U$2 ( \48727 , \48726 );
nor \g135515/U$1 ( \48728 , \48727 , \40060 );
not \g130407/U$3 ( \48729 , \47948 );
and \g130436/U$2 ( \48730 , \48568 , \47960 );
and \g130436/U$3 ( \48731 , \47959 , \48515 );
nor \g130436/U$1 ( \48732 , \48730 , \48731 );
not \g130407/U$4 ( \48733 , \48732 );
or \g130407/U$2 ( \48734 , \48729 , \48733 );
or \g130407/U$5 ( \48735 , \48732 , \47948 );
nand \g130407/U$1 ( \48736 , \48734 , \48735 );
xor \g456038/U$4 ( \48737 , \48728 , \48736 );
not \g129927/U$3 ( \48738 , \47997 );
and \g129970/U$2 ( \48739 , \48051 , \48064 );
and \g129970/U$3 ( \48740 , \48063 , \48018 );
nor \g129970/U$1 ( \48741 , \48739 , \48740 );
not \g129927/U$4 ( \48742 , \48741 );
or \g129927/U$2 ( \48743 , \48738 , \48742 );
or \g129927/U$5 ( \48744 , \48741 , \47997 );
nand \g129927/U$1 ( \48745 , \48743 , \48744 );
and \g456038/U$3 ( \48746 , \48737 , \48745 );
and \g456038/U$5 ( \48747 , \48728 , \48736 );
nor \g456038/U$2 ( \48748 , \48746 , \48747 );
xor \g129435/U$4 ( \48749 , \48722 , \48748 );
and \g130299/U$2 ( \48750 , \48349 , \47914 );
and \g130299/U$3 ( \48751 , \47913 , \48353 );
nor \g130299/U$1 ( \48752 , \48750 , \48751 );
and \g130265/U$2 ( \48753 , \48752 , \47977 );
not \g130265/U$4 ( \48754 , \48752 );
and \g130265/U$3 ( \48755 , \48754 , \47976 );
nor \g130265/U$1 ( \48756 , \48753 , \48755 );
not \g130112/U$3 ( \48757 , \47935 );
and \g130150/U$2 ( \48758 , \48117 , \47930 );
and \g130150/U$3 ( \48759 , \47931 , \48138 );
nor \g130150/U$1 ( \48760 , \48758 , \48759 );
not \g130112/U$4 ( \48761 , \48760 );
or \g130112/U$2 ( \48762 , \48757 , \48761 );
or \g130112/U$5 ( \48763 , \48760 , \47935 );
nand \g130112/U$1 ( \48764 , \48762 , \48763 );
xor \g456011/U$4 ( \48765 , \48756 , \48764 );
not \g129573/U$3 ( \48766 , \48323 );
and \g129618/U$2 ( \48767 , \47970 , \48334 );
and \g129618/U$3 ( \48768 , \48335 , \47962 );
nor \g129618/U$1 ( \48769 , \48767 , \48768 );
not \g129573/U$4 ( \48770 , \48769 );
or \g129573/U$2 ( \48771 , \48766 , \48770 );
or \g129573/U$5 ( \48772 , \48769 , \48323 );
nand \g129573/U$1 ( \48773 , \48771 , \48772 );
and \g456011/U$3 ( \48774 , \48765 , \48773 );
and \g456011/U$5 ( \48775 , \48756 , \48764 );
nor \g456011/U$2 ( \48776 , \48774 , \48775 );
and \g129435/U$3 ( \48777 , \48749 , \48776 );
and \g129435/U$5 ( \48778 , \48722 , \48748 );
or \g129435/U$2 ( \48779 , \48777 , \48778 );
xor \g128925/U$4 ( \48780 , \48716 , \48779 );
xor \g456032/U$1 ( \48781 , \48570 , \48578 );
xor \g456032/U$1_r1 ( \48782 , \48781 , \48587 );
not \g129138/U$3 ( \48783 , \48667 );
not \g129172/U$3 ( \48784 , \48697 );
not \g129172/U$4 ( \48785 , \48487 );
and \g129172/U$2 ( \48786 , \48784 , \48785 );
and \g129172/U$5 ( \48787 , \48697 , \48487 );
nor \g129172/U$1 ( \48788 , \48786 , \48787 );
not \g129138/U$4 ( \48789 , \48788 );
or \g129138/U$2 ( \48790 , \48783 , \48789 );
or \g129138/U$5 ( \48791 , \48788 , \48667 );
nand \g129138/U$1 ( \48792 , \48790 , \48791 );
xor \g455981/U$4 ( \48793 , \48782 , \48792 );
not \g130022/U$3 ( \48794 , \47997 );
and \g130064/U$2 ( \48795 , \48051 , \48063 );
and \g130064/U$3 ( \48796 , \48064 , \48117 );
nor \g130064/U$1 ( \48797 , \48795 , \48796 );
not \g130022/U$4 ( \48798 , \48797 );
or \g130022/U$2 ( \48799 , \48794 , \48798 );
or \g130022/U$5 ( \48800 , \48797 , \47997 );
nand \g130022/U$1 ( \48801 , \48799 , \48800 );
not \g130191/U$3 ( \48802 , \47935 );
and \g130230/U$2 ( \48803 , \48353 , \47931 );
and \g130230/U$3 ( \48804 , \47930 , \48138 );
nor \g130230/U$1 ( \48805 , \48803 , \48804 );
not \g130191/U$4 ( \48806 , \48805 );
or \g130191/U$2 ( \48807 , \48802 , \48806 );
or \g130191/U$5 ( \48808 , \48805 , \47935 );
nand \g130191/U$1 ( \48809 , \48807 , \48808 );
xor \g129595/U$4 ( \48810 , \48801 , \48809 );
not \g129675/U$3 ( \48811 , \48323 );
and \g129710/U$2 ( \48812 , \47950 , \48335 );
and \g129710/U$3 ( \48813 , \48334 , \47962 );
nor \g129710/U$1 ( \48814 , \48812 , \48813 );
not \g129675/U$4 ( \48815 , \48814 );
or \g129675/U$2 ( \48816 , \48811 , \48815 );
or \g129675/U$5 ( \48817 , \48814 , \48323 );
nand \g129675/U$1 ( \48818 , \48816 , \48817 );
and \g129595/U$3 ( \48819 , \48810 , \48818 );
and \g129595/U$5 ( \48820 , \48801 , \48809 );
or \g129595/U$2 ( \48821 , \48819 , \48820 );
not \g130478/U$3 ( \48822 , \47948 );
and \g130509/U$2 ( \48823 , \48726 , \47960 );
and \g130509/U$3 ( \48824 , \47959 , \48568 );
nor \g130509/U$1 ( \48825 , \48823 , \48824 );
not \g130478/U$4 ( \48826 , \48825 );
or \g130478/U$2 ( \48827 , \48822 , \48826 );
or \g130478/U$5 ( \48828 , \48825 , \47948 );
nand \g130478/U$1 ( \48829 , \48827 , \48828 );
and \g130693/U$2 ( \48830 , \47737 , \47664 );
not \g130693/U$4 ( \48831 , \47737 );
and \g130693/U$3 ( \48832 , \48831 , \47665 );
or \g130693/U$1 ( \48833 , \48830 , \48832 );
not \g135516/U$2 ( \48834 , \48833 );
nor \g135516/U$1 ( \48835 , \48834 , \40060 );
xor \g129769/U$4 ( \48836 , \48829 , \48835 );
not \g129840/U$3 ( \48837 , \48159 );
and \g129876/U$2 ( \48838 , \48018 , \48155 );
and \g129876/U$3 ( \48839 , \48154 , \47942 );
nor \g129876/U$1 ( \48840 , \48838 , \48839 );
not \g129840/U$4 ( \48841 , \48840 );
or \g129840/U$2 ( \48842 , \48837 , \48841 );
or \g129840/U$5 ( \48843 , \48840 , \48159 );
nand \g129840/U$1 ( \48844 , \48842 , \48843 );
and \g129769/U$3 ( \48845 , \48836 , \48844 );
and \g129769/U$5 ( \48846 , \48829 , \48835 );
or \g129769/U$2 ( \48847 , \48845 , \48846 );
xor \g129304/U$4 ( \48848 , \48821 , \48847 );
not \g129371/U$3 ( \48849 , \48685 );
and \g133053/U$2 ( \48850 , \48683 , \48473 );
not \g133053/U$4 ( \48851 , \48683 );
and \g133053/U$3 ( \48852 , \48851 , \48474 );
nor \g133053/U$1 ( \48853 , \48850 , \48852 );
not \g133151/U$1 ( \48854 , \48681 );
and \g133095/U$2 ( \48855 , \48683 , \48854 );
not \g133095/U$4 ( \48856 , \48683 );
and \g133095/U$3 ( \48857 , \48856 , \48681 );
or \g133095/U$1 ( \48858 , \48855 , \48857 );
not \g133084/U$1 ( \48859 , \48858 );
and \g133037/U$1 ( \48860 , \48853 , \48859 );
nand \g129421/U$1 ( \48861 , \48860 , \47894 );
not \g129371/U$4 ( \48862 , \48861 );
or \g129371/U$2 ( \48863 , \48849 , \48862 );
or \g129371/U$5 ( \48864 , \48861 , \48685 );
nand \g129371/U$1 ( \48865 , \48863 , \48864 );
and \g129304/U$3 ( \48866 , \48848 , \48865 );
and \g129304/U$5 ( \48867 , \48821 , \48847 );
or \g129304/U$2 ( \48868 , \48866 , \48867 );
and \g455981/U$3 ( \48869 , \48793 , \48868 );
and \g455981/U$5 ( \48870 , \48782 , \48792 );
nor \g455981/U$2 ( \48871 , \48869 , \48870 );
and \g128925/U$3 ( \48872 , \48780 , \48871 );
and \g128925/U$5 ( \48873 , \48716 , \48779 );
or \g128925/U$2 ( \48874 , \48872 , \48873 );
not \g128897/U$4 ( \48875 , \48874 );
or \g128897/U$2 ( \48876 , \48706 , \48875 );
or \g128897/U$5 ( \48877 , \48874 , \48705 );
nand \g128897/U$1 ( \48878 , \48876 , \48877 );
not \g128872/U$4 ( \48879 , \48878 );
or \g128872/U$2 ( \48880 , \48703 , \48879 );
or \g128872/U$5 ( \48881 , \48878 , \48702 );
nand \g128872/U$1 ( \48882 , \48880 , \48881 );
xor \g128925/U$1 ( \48883 , \48716 , \48779 );
xor \g128925/U$1_r1 ( \48884 , \48883 , \48871 );
xor \g129007/U$1 ( \48885 , \48652 , \48658 );
xor \g129007/U$1_r1 ( \48886 , \48885 , \48699 );
or \g128888/U$2 ( \48887 , \48884 , \48886 );
not \g128895/U$3 ( \48888 , \48886 );
not \g128895/U$4 ( \48889 , \48884 );
or \g128895/U$2 ( \48890 , \48888 , \48889 );
xor \g456011/U$1 ( \48891 , \48756 , \48764 );
xor \g456011/U$1_r1 ( \48892 , \48891 , \48773 );
xor \g456038/U$1 ( \48893 , \48728 , \48736 );
xor \g456038/U$1_r1 ( \48894 , \48893 , \48745 );
and \g129182/U$2 ( \48895 , \48892 , \48894 );
not \g129202/U$3 ( \48896 , \48892 );
not \g129202/U$4 ( \48897 , \48894 );
and \g129202/U$2 ( \48898 , \48896 , \48897 );
xor \g129251/U$1 ( \48899 , \48679 , \48685 );
xor \g129251/U$1_r1 ( \48900 , \48899 , \48694 );
nor \g129202/U$1 ( \48901 , \48898 , \48900 );
nor \g129182/U$1 ( \48902 , \48895 , \48901 );
xor \g129435/U$1 ( \48903 , \48722 , \48748 );
xor \g129435/U$1_r1 ( \48904 , \48903 , \48776 );
or \g128982/U$2 ( \48905 , \48902 , \48904 );
not \g128992/U$3 ( \48906 , \48904 );
not \g128992/U$4 ( \48907 , \48902 );
or \g128992/U$2 ( \48908 , \48906 , \48907 );
xor \g455981/U$1 ( \48909 , \48782 , \48792 );
xor \g455981/U$1_r1 ( \48910 , \48909 , \48868 );
nand \g128992/U$1 ( \48911 , \48908 , \48910 );
nand \g128982/U$1 ( \48912 , \48905 , \48911 );
nand \g128895/U$1 ( \48913 , \48890 , \48912 );
nand \g128888/U$1 ( \48914 , \48887 , \48913 );
xor \g129453/U$1 ( \48915 , \48894 , \48892 );
not \g129199/U$3 ( \48916 , \48915 );
not \g129199/U$4 ( \48917 , \48900 );
or \g129199/U$2 ( \48918 , \48916 , \48917 );
or \g129199/U$5 ( \48919 , \48900 , \48915 );
nand \g129199/U$1 ( \48920 , \48918 , \48919 );
xor \g129769/U$1 ( \48921 , \48829 , \48835 );
xor \g129769/U$1_r1 ( \48922 , \48921 , \48844 );
not \g129225/U$3 ( \48923 , \48922 );
xor \g129595/U$1 ( \48924 , \48801 , \48809 );
xor \g129595/U$1_r1 ( \48925 , \48924 , \48818 );
not \g129225/U$4 ( \48926 , \48925 );
or \g129225/U$2 ( \48927 , \48923 , \48926 );
or \g129237/U$2 ( \48928 , \48925 , \48922 );
not \g129468/U$3 ( \48929 , \48483 );
and \g129511/U$2 ( \48930 , \47970 , \48479 );
and \g129511/U$3 ( \48931 , \48478 , \47972 );
nor \g129511/U$1 ( \48932 , \48930 , \48931 );
not \g129468/U$4 ( \48933 , \48932 );
or \g129468/U$2 ( \48934 , \48929 , \48933 );
or \g129468/U$5 ( \48935 , \48932 , \48483 );
nand \g129468/U$1 ( \48936 , \48934 , \48935 );
and \g130373/U$2 ( \48937 , \48349 , \47913 );
and \g130373/U$3 ( \48938 , \47914 , \48515 );
nor \g130373/U$1 ( \48939 , \48937 , \48938 );
and \g130332/U$2 ( \48940 , \48939 , \47977 );
not \g130332/U$4 ( \48941 , \48939 );
and \g130332/U$3 ( \48942 , \48941 , \47976 );
nor \g130332/U$1 ( \48943 , \48940 , \48942 );
xor \g129276/U$1 ( \48944 , \48936 , \48943 );
not \g129370/U$1 ( \48945 , \48865 );
xor \g129276/U$1_r1 ( \48946 , \48944 , \48945 );
nand \g129237/U$1 ( \48947 , \48928 , \48946 );
nand \g129225/U$1 ( \48948 , \48927 , \48947 );
xor \g128957/U$4 ( \48949 , \48920 , \48948 );
not \g130546/U$3 ( \48950 , \47948 );
and \g130575/U$2 ( \48951 , \48726 , \47959 );
and \g130575/U$3 ( \48952 , \47960 , \48833 );
nor \g130575/U$1 ( \48953 , \48951 , \48952 );
not \g130546/U$4 ( \48954 , \48953 );
or \g130546/U$2 ( \48955 , \48950 , \48954 );
or \g130546/U$5 ( \48956 , \48953 , \47948 );
nand \g130546/U$1 ( \48957 , \48955 , \48956 );
and \g130437/U$2 ( \48958 , \48568 , \47914 );
and \g130437/U$3 ( \48959 , \47913 , \48515 );
nor \g130437/U$1 ( \48960 , \48958 , \48959 );
and \g130408/U$2 ( \48961 , \48960 , \47977 );
not \g130408/U$4 ( \48962 , \48960 );
and \g130408/U$3 ( \48963 , \48962 , \47976 );
nor \g130408/U$1 ( \48964 , \48961 , \48963 );
xor \g456039/U$4 ( \48965 , \48957 , \48964 );
not \g129928/U$3 ( \48966 , \48159 );
and \g129971/U$2 ( \48967 , \48051 , \48155 );
and \g129971/U$3 ( \48968 , \48154 , \48018 );
nor \g129971/U$1 ( \48969 , \48967 , \48968 );
not \g129928/U$4 ( \48970 , \48969 );
or \g129928/U$2 ( \48971 , \48966 , \48970 );
or \g129928/U$5 ( \48972 , \48969 , \48159 );
nand \g129928/U$1 ( \48973 , \48971 , \48972 );
and \g456039/U$3 ( \48974 , \48965 , \48973 );
and \g456039/U$5 ( \48975 , \48957 , \48964 );
nor \g456039/U$2 ( \48976 , \48974 , \48975 );
xor \g130747/U$1 ( \48977 , \47662 , \41708 );
not \g135517/U$2 ( \48978 , \48977 );
nor \g135517/U$1 ( \48979 , \48978 , \40060 );
not \g130266/U$3 ( \48980 , \47935 );
and \g130300/U$2 ( \48981 , \48349 , \47931 );
and \g130300/U$3 ( \48982 , \47930 , \48353 );
nor \g130300/U$1 ( \48983 , \48981 , \48982 );
not \g130266/U$4 ( \48984 , \48983 );
or \g130266/U$2 ( \48985 , \48980 , \48984 );
or \g130266/U$5 ( \48986 , \48983 , \47935 );
nand \g130266/U$1 ( \48987 , \48985 , \48986 );
xor \g456048/U$4 ( \48988 , \48979 , \48987 );
not \g130113/U$3 ( \48989 , \47997 );
and \g130151/U$2 ( \48990 , \48117 , \48063 );
and \g130151/U$3 ( \48991 , \48064 , \48138 );
nor \g130151/U$1 ( \48992 , \48990 , \48991 );
not \g130113/U$4 ( \48993 , \48992 );
or \g130113/U$2 ( \48994 , \48989 , \48993 );
or \g130113/U$5 ( \48995 , \48992 , \47997 );
nand \g130113/U$1 ( \48996 , \48994 , \48995 );
and \g456048/U$3 ( \48997 , \48988 , \48996 );
and \g456048/U$5 ( \48998 , \48979 , \48987 );
nor \g456048/U$2 ( \48999 , \48997 , \48998 );
xor \g129117/U$1 ( \49000 , \48976 , \48999 );
and \g129794/U$2 ( \49001 , \47950 , \48334 );
and \g129794/U$3 ( \49002 , \48335 , \47942 );
nor \g129794/U$1 ( \49003 , \49001 , \49002 );
not \g129748/U$3 ( \49004 , \49003 );
not \g129748/U$4 ( \49005 , \48323 );
and \g129748/U$2 ( \49006 , \49004 , \49005 );
and \g129748/U$5 ( \49007 , \49003 , \48323 );
nor \g129748/U$1 ( \49008 , \49006 , \49007 );
xor \g133252/U$1 ( \49009 , \21118 , \13123 );
xor \g133252/U$1_r1 ( \49010 , \49009 , \40005 );
xor \g133202/U$1 ( \49011 , \20875 , \12879 );
xor \g133202/U$1_r1 ( \49012 , \49011 , \40008 );
nand \g133175/U$1 ( \49013 , \49010 , \49012 );
and \g133130/U$1 ( \49014 , \48681 , \49013 );
xor \g129252/U$4 ( \49015 , \49008 , \49014 );
and \g129394/U$2 ( \49016 , \47894 , \48858 );
and \g129394/U$3 ( \49017 , \48860 , \47972 );
nor \g129394/U$1 ( \49018 , \49016 , \49017 );
not \g129337/U$3 ( \49019 , \49018 );
not \g129337/U$4 ( \49020 , \48685 );
and \g129337/U$2 ( \49021 , \49019 , \49020 );
and \g129337/U$5 ( \49022 , \49018 , \48685 );
nor \g129337/U$1 ( \49023 , \49021 , \49022 );
and \g129252/U$3 ( \49024 , \49015 , \49023 );
and \g129252/U$5 ( \49025 , \49008 , \49014 );
or \g129252/U$2 ( \49026 , \49024 , \49025 );
xor \g129117/U$1_r1 ( \49027 , \49000 , \49026 );
and \g129619/U$2 ( \49028 , \47970 , \48478 );
and \g129619/U$3 ( \49029 , \48479 , \47962 );
nor \g129619/U$1 ( \49030 , \49028 , \49029 );
not \g129574/U$3 ( \49031 , \49030 );
not \g129574/U$4 ( \49032 , \48483 );
and \g129574/U$2 ( \49033 , \49031 , \49032 );
and \g129574/U$5 ( \49034 , \49030 , \48483 );
nor \g129574/U$1 ( \49035 , \49033 , \49034 );
and \g130510/U$2 ( \49036 , \48726 , \47914 );
and \g130510/U$3 ( \49037 , \47913 , \48568 );
nor \g130510/U$1 ( \49038 , \49036 , \49037 );
and \g130479/U$2 ( \49039 , \49038 , \47976 );
not \g130479/U$4 ( \49040 , \49038 );
and \g130479/U$3 ( \49041 , \49040 , \47977 );
nor \g130479/U$1 ( \49042 , \49039 , \49041 );
and \g130644/U$2 ( \49043 , \48833 , \47959 );
and \g130644/U$3 ( \49044 , \47960 , \48977 );
nor \g130644/U$1 ( \49045 , \49043 , \49044 );
not \g130608/U$3 ( \49046 , \49045 );
not \g130608/U$4 ( \49047 , \47948 );
and \g130608/U$2 ( \49048 , \49046 , \49047 );
and \g130608/U$5 ( \49049 , \49045 , \47948 );
nor \g130608/U$1 ( \49050 , \49048 , \49049 );
xor \g456005/U$5 ( \49051 , \49042 , \49050 );
and \g129877/U$2 ( \49052 , \48018 , \48335 );
and \g129877/U$3 ( \49053 , \48334 , \47942 );
nor \g129877/U$1 ( \49054 , \49052 , \49053 );
not \g129841/U$3 ( \49055 , \49054 );
not \g129841/U$4 ( \49056 , \48323 );
and \g129841/U$2 ( \49057 , \49055 , \49056 );
and \g129841/U$5 ( \49058 , \49054 , \48323 );
nor \g129841/U$1 ( \49059 , \49057 , \49058 );
and \g456005/U$4 ( \49060 , \49051 , \49059 );
and \g456005/U$6 ( \49061 , \49042 , \49050 );
or \g456005/U$3 ( \49062 , \49060 , \49061 );
xor \g129273/U$4 ( \49063 , \49035 , \49062 );
not \g129373/U$3 ( \49064 , \49014 );
and \g133125/U$2 ( \49065 , \49012 , \48681 );
not \g133125/U$4 ( \49066 , \49012 );
and \g133125/U$3 ( \49067 , \49066 , \48854 );
nor \g133125/U$1 ( \49068 , \49065 , \49067 );
not \g135549/U$2 ( \49069 , \49068 );
not \g133251/U$1 ( \49070 , \49010 );
and \g133155/U$2 ( \49071 , \49012 , \49070 );
not \g133155/U$4 ( \49072 , \49012 );
and \g133155/U$3 ( \49073 , \49072 , \49010 );
or \g133155/U$1 ( \49074 , \49071 , \49073 );
nor \g135549/U$1 ( \49075 , \49069 , \49074 );
nand \g129422/U$1 ( \49076 , \49075 , \47894 );
not \g129373/U$4 ( \49077 , \49076 );
or \g129373/U$2 ( \49078 , \49064 , \49077 );
or \g129373/U$5 ( \49079 , \49076 , \49014 );
nand \g129373/U$1 ( \49080 , \49078 , \49079 );
not \g129372/U$1 ( \49081 , \49080 );
and \g129273/U$3 ( \49082 , \49063 , \49081 );
and \g129273/U$5 ( \49083 , \49035 , \49062 );
or \g129273/U$2 ( \49084 , \49082 , \49083 );
or \g129047/U$2 ( \49085 , \49027 , \49084 );
not \g129067/U$3 ( \49086 , \49084 );
not \g129067/U$4 ( \49087 , \49027 );
or \g129067/U$2 ( \49088 , \49086 , \49087 );
xor \g129252/U$1 ( \49089 , \49008 , \49014 );
xor \g129252/U$1_r1 ( \49090 , \49089 , \49023 );
and \g130065/U$2 ( \49091 , \48051 , \48154 );
and \g130065/U$3 ( \49092 , \48155 , \48117 );
nor \g130065/U$1 ( \49093 , \49091 , \49092 );
not \g130023/U$3 ( \49094 , \49093 );
not \g130023/U$4 ( \49095 , \48159 );
and \g130023/U$2 ( \49096 , \49094 , \49095 );
and \g130023/U$5 ( \49097 , \49093 , \48159 );
nor \g130023/U$1 ( \49098 , \49096 , \49097 );
and \g130804/U$2 ( \49099 , \47658 , \47659 );
not \g130804/U$4 ( \49100 , \47658 );
and \g130804/U$3 ( \49101 , \49100 , \47660 );
or \g130804/U$1 ( \49102 , \49099 , \49101 );
nand \g130775/U$1 ( \49103 , \40061 , \49102 );
xor \g129596/U$4 ( \49104 , \49098 , \49103 );
and \g129711/U$2 ( \49105 , \47950 , \48479 );
and \g129711/U$3 ( \49106 , \48478 , \47962 );
nor \g129711/U$1 ( \49107 , \49105 , \49106 );
not \g129676/U$3 ( \49108 , \49107 );
not \g129676/U$4 ( \49109 , \48483 );
and \g129676/U$2 ( \49110 , \49108 , \49109 );
and \g129676/U$5 ( \49111 , \49107 , \48483 );
nor \g129676/U$1 ( \49112 , \49110 , \49111 );
and \g129596/U$3 ( \49113 , \49104 , \49112 );
and \g129596/U$5 ( \49114 , \49098 , \49103 );
or \g129596/U$2 ( \49115 , \49113 , \49114 );
not \g129564/U$2 ( \49116 , \49115 );
xor \g456048/U$1 ( \49117 , \48979 , \48987 );
xor \g456048/U$1_r1 ( \49118 , \49117 , \48996 );
nor \g129564/U$1 ( \49119 , \49116 , \49118 );
or \g129187/U$2 ( \49120 , \49090 , \49119 );
not \g129565/U$2 ( \49121 , \49115 );
nand \g129565/U$1 ( \49122 , \49121 , \49118 );
nand \g129187/U$1 ( \49123 , \49120 , \49122 );
nand \g129067/U$1 ( \49124 , \49088 , \49123 );
nand \g129047/U$1 ( \49125 , \49085 , \49124 );
and \g128957/U$3 ( \49126 , \48949 , \49125 );
and \g128957/U$5 ( \49127 , \48920 , \48948 );
or \g128957/U$2 ( \49128 , \49126 , \49127 );
xor \g129304/U$1 ( \49129 , \48821 , \48847 );
xor \g129304/U$1_r1 ( \49130 , \49129 , \48865 );
xor \g129276/U$4 ( \49131 , \48936 , \48943 );
and \g129276/U$3 ( \49132 , \49131 , \48945 );
and \g129276/U$5 ( \49133 , \48936 , \48943 );
or \g129276/U$2 ( \49134 , \49132 , \49133 );
and \g129088/U$2 ( \49135 , \49130 , \49134 );
not \g129099/U$3 ( \49136 , \49130 );
not \g129099/U$4 ( \49137 , \49134 );
and \g129099/U$2 ( \49138 , \49136 , \49137 );
xor \g129117/U$4 ( \49139 , \48976 , \48999 );
and \g129117/U$3 ( \49140 , \49139 , \49026 );
and \g129117/U$5 ( \49141 , \48976 , \48999 );
or \g129117/U$2 ( \49142 , \49140 , \49141 );
nor \g129099/U$1 ( \49143 , \49138 , \49142 );
nor \g129088/U$1 ( \49144 , \49135 , \49143 );
not \g129008/U$1 ( \49145 , \49144 );
and \g128908/U$2 ( \49146 , \49128 , \49145 );
not \g128915/U$3 ( \49147 , \49128 );
not \g128915/U$4 ( \49148 , \49145 );
and \g128915/U$2 ( \49149 , \49147 , \49148 );
not \g128968/U$3 ( \49150 , \48910 );
not \g128968/U$4 ( \49151 , \48902 );
and \g128968/U$2 ( \49152 , \49150 , \49151 );
and \g128968/U$5 ( \49153 , \48910 , \48902 );
nor \g128968/U$1 ( \49154 , \49152 , \49153 );
xnor \g455930/U$1 ( \49155 , \49154 , \48904 );
nor \g128915/U$1 ( \49156 , \49149 , \49155 );
nor \g128908/U$1 ( \49157 , \49146 , \49156 );
xor \g130860/U$1 ( \49158 , \47656 , \42174 );
not \g135518/U$2 ( \49159 , \49158 );
nor \g135518/U$1 ( \49160 , \49159 , \40060 );
not \g130673/U$3 ( \49161 , \47948 );
and \g130699/U$2 ( \49162 , \49102 , \47960 );
and \g130699/U$3 ( \49163 , \47959 , \48977 );
nor \g130699/U$1 ( \49164 , \49162 , \49163 );
not \g130673/U$4 ( \49165 , \49164 );
or \g130673/U$2 ( \49166 , \49161 , \49165 );
or \g130673/U$5 ( \49167 , \49164 , \47948 );
nand \g130673/U$1 ( \49168 , \49166 , \49167 );
xor \g456049/U$4 ( \49169 , \49160 , \49168 );
not \g130114/U$3 ( \49170 , \48159 );
and \g130152/U$2 ( \49171 , \48117 , \48154 );
and \g130152/U$3 ( \49172 , \48155 , \48138 );
nor \g130152/U$1 ( \49173 , \49171 , \49172 );
not \g130114/U$4 ( \49174 , \49173 );
or \g130114/U$2 ( \49175 , \49170 , \49174 );
or \g130114/U$5 ( \49176 , \49173 , \48159 );
nand \g130114/U$1 ( \49177 , \49175 , \49176 );
and \g456049/U$3 ( \49178 , \49169 , \49177 );
and \g456049/U$5 ( \49179 , \49160 , \49168 );
nor \g456049/U$2 ( \49180 , \49178 , \49179 );
xor \g456005/U$9 ( \49181 , \49042 , \49050 );
xor \g456005/U$9_r1 ( \49182 , \49181 , \49059 );
and \g456005/U$8 ( \49183 , \49180 , \49182 );
xor \g129596/U$1 ( \49184 , \49098 , \49103 );
xor \g129596/U$1_r1 ( \49185 , \49184 , \49112 );
xor \g456005/U$11 ( \49186 , \49042 , \49050 );
xor \g456005/U$11_r1 ( \49187 , \49186 , \49059 );
and \g456005/U$10 ( \49188 , \49185 , \49187 );
and \g456005/U$12 ( \49189 , \49180 , \49185 );
or \g456005/U$7 ( \49190 , \49183 , \49188 , \49189 );
not \g129042/U$3 ( \49191 , \49190 );
and \g130576/U$2 ( \49192 , \48726 , \47913 );
and \g130576/U$3 ( \49193 , \47914 , \48833 );
nor \g130576/U$1 ( \49194 , \49192 , \49193 );
and \g130547/U$2 ( \49195 , \49194 , \47977 );
not \g130547/U$4 ( \49196 , \49194 );
and \g130547/U$3 ( \49197 , \49196 , \47976 );
nor \g130547/U$1 ( \49198 , \49195 , \49197 );
not \g130409/U$3 ( \49199 , \47935 );
and \g130438/U$2 ( \49200 , \48568 , \47931 );
and \g130438/U$3 ( \49201 , \47930 , \48515 );
nor \g130438/U$1 ( \49202 , \49200 , \49201 );
not \g130409/U$4 ( \49203 , \49202 );
or \g130409/U$2 ( \49204 , \49199 , \49203 );
or \g130409/U$5 ( \49205 , \49202 , \47935 );
nand \g130409/U$1 ( \49206 , \49204 , \49205 );
xor \g456040/U$4 ( \49207 , \49198 , \49206 );
not \g129929/U$3 ( \49208 , \48323 );
and \g129972/U$2 ( \49209 , \48051 , \48335 );
and \g129972/U$3 ( \49210 , \48334 , \48018 );
nor \g129972/U$1 ( \49211 , \49209 , \49210 );
not \g129929/U$4 ( \49212 , \49211 );
or \g129929/U$2 ( \49213 , \49208 , \49212 );
or \g129929/U$5 ( \49214 , \49211 , \48323 );
nand \g129929/U$1 ( \49215 , \49213 , \49214 );
and \g456040/U$3 ( \49216 , \49207 , \49215 );
and \g456040/U$5 ( \49217 , \49198 , \49206 );
nor \g456040/U$2 ( \49218 , \49216 , \49217 );
xor \g129118/U$4 ( \49219 , \49080 , \49218 );
and \g129795/U$2 ( \49220 , \47950 , \48478 );
and \g129795/U$3 ( \49221 , \48479 , \47942 );
nor \g129795/U$1 ( \49222 , \49220 , \49221 );
not \g129749/U$3 ( \49223 , \49222 );
not \g129749/U$4 ( \49224 , \48483 );
and \g129749/U$2 ( \49225 , \49223 , \49224 );
and \g129749/U$5 ( \49226 , \49222 , \48483 );
nor \g129749/U$1 ( \49227 , \49225 , \49226 );
xor \g133353/U$1 ( \49228 , \21605 , \13617 );
xor \g133353/U$1_r1 ( \49229 , \49228 , \39999 );
xor \g133295/U$1 ( \49230 , \21361 , \13370 );
xor \g133295/U$1_r1 ( \49231 , \49230 , \40002 );
nand \g133273/U$1 ( \49232 , \49229 , \49231 );
and \g133222/U$1 ( \49233 , \49010 , \49232 );
xor \g129253/U$4 ( \49234 , \49227 , \49233 );
and \g129395/U$2 ( \49235 , \47894 , \49074 );
and \g129395/U$3 ( \49236 , \49075 , \47972 );
nor \g129395/U$1 ( \49237 , \49235 , \49236 );
not \g129338/U$3 ( \49238 , \49237 );
not \g129338/U$4 ( \49239 , \49014 );
and \g129338/U$2 ( \49240 , \49238 , \49239 );
and \g129338/U$5 ( \49241 , \49237 , \49014 );
nor \g129338/U$1 ( \49242 , \49240 , \49241 );
and \g129253/U$3 ( \49243 , \49234 , \49242 );
and \g129253/U$5 ( \49244 , \49227 , \49233 );
or \g129253/U$2 ( \49245 , \49243 , \49244 );
and \g129118/U$3 ( \49246 , \49219 , \49245 );
and \g129118/U$5 ( \49247 , \49080 , \49218 );
or \g129118/U$2 ( \49248 , \49246 , \49247 );
not \g129175/U$3 ( \49249 , \49118 );
not \g129175/U$4 ( \49250 , \49090 );
or \g129175/U$2 ( \49251 , \49249 , \49250 );
or \g129175/U$5 ( \49252 , \49090 , \49118 );
nand \g129175/U$1 ( \49253 , \49251 , \49252 );
not \g129140/U$3 ( \49254 , \49253 );
not \g129140/U$4 ( \49255 , \49115 );
and \g129140/U$2 ( \49256 , \49254 , \49255 );
and \g129140/U$5 ( \49257 , \49253 , \49115 );
nor \g129140/U$1 ( \49258 , \49256 , \49257 );
xor \g129079/U$1 ( \49259 , \49248 , \49258 );
not \g129042/U$4 ( \49260 , \49259 );
or \g129042/U$2 ( \49261 , \49191 , \49260 );
or \g129042/U$5 ( \49262 , \49259 , \49190 );
nand \g129042/U$1 ( \49263 , \49261 , \49262 );
not \g129843/U$3 ( \49264 , \48483 );
and \g129878/U$2 ( \49265 , \48018 , \48479 );
and \g129878/U$3 ( \49266 , \48478 , \47942 );
nor \g129878/U$1 ( \49267 , \49265 , \49266 );
not \g129843/U$4 ( \49268 , \49267 );
or \g129843/U$2 ( \49269 , \49264 , \49268 );
or \g129843/U$5 ( \49270 , \49267 , \48483 );
nand \g129843/U$1 ( \49271 , \49269 , \49270 );
and \g130700/U$2 ( \49272 , \49102 , \47914 );
and \g130700/U$3 ( \49273 , \47913 , \48977 );
nor \g130700/U$1 ( \49274 , \49272 , \49273 );
and \g130674/U$2 ( \49275 , \49274 , \47976 );
not \g130674/U$4 ( \49276 , \49274 );
and \g130674/U$3 ( \49277 , \49276 , \47977 );
nor \g130674/U$1 ( \49278 , \49275 , \49277 );
and \g130914/U$2 ( \49279 , \47652 , \47653 );
not \g130914/U$4 ( \49280 , \47652 );
and \g130914/U$3 ( \49281 , \49280 , \47654 );
or \g130914/U$1 ( \49282 , \49279 , \49281 );
and \g130812/U$2 ( \49283 , \49282 , \47960 );
and \g130812/U$3 ( \49284 , \47959 , \49158 );
nor \g130812/U$1 ( \49285 , \49283 , \49284 );
not \g130784/U$3 ( \49286 , \49285 );
not \g130784/U$4 ( \49287 , \47948 );
and \g130784/U$2 ( \49288 , \49286 , \49287 );
and \g130784/U$5 ( \49289 , \49285 , \47948 );
nor \g130784/U$1 ( \49290 , \49288 , \49289 );
xor \g130043/U$4 ( \49291 , \49278 , \49290 );
and \g130153/U$2 ( \49292 , \48117 , \48334 );
and \g130153/U$3 ( \49293 , \48335 , \48138 );
nor \g130153/U$1 ( \49294 , \49292 , \49293 );
not \g130115/U$3 ( \49295 , \49294 );
not \g130115/U$4 ( \49296 , \48323 );
and \g130115/U$2 ( \49297 , \49295 , \49296 );
and \g130115/U$5 ( \49298 , \49294 , \48323 );
nor \g130115/U$1 ( \49299 , \49297 , \49298 );
and \g130043/U$3 ( \49300 , \49291 , \49299 );
and \g130043/U$5 ( \49301 , \49278 , \49290 );
or \g130043/U$2 ( \49302 , \49300 , \49301 );
xor \g455976/U$5 ( \49303 , \49271 , \49302 );
and \g129514/U$2 ( \49304 , \47970 , \49075 );
and \g129514/U$3 ( \49305 , \49074 , \47972 );
nor \g129514/U$1 ( \49306 , \49304 , \49305 );
not \g129471/U$3 ( \49307 , \49306 );
not \g129471/U$4 ( \49308 , \49014 );
and \g129471/U$2 ( \49309 , \49307 , \49308 );
and \g129471/U$5 ( \49310 , \49306 , \49014 );
nor \g129471/U$1 ( \49311 , \49309 , \49310 );
and \g455976/U$4 ( \49312 , \49303 , \49311 );
and \g455976/U$6 ( \49313 , \49271 , \49302 );
or \g455976/U$3 ( \49314 , \49312 , \49313 );
not \g130267/U$3 ( \49315 , \47997 );
and \g130301/U$2 ( \49316 , \48349 , \48064 );
and \g130301/U$3 ( \49317 , \48063 , \48353 );
nor \g130301/U$1 ( \49318 , \49316 , \49317 );
not \g130267/U$4 ( \49319 , \49318 );
or \g130267/U$2 ( \49320 , \49315 , \49319 );
or \g130267/U$5 ( \49321 , \49318 , \47997 );
nand \g130267/U$1 ( \49322 , \49320 , \49321 );
xor \g129496/U$1 ( \49323 , \49271 , \49322 );
not \g129575/U$3 ( \49324 , \48685 );
and \g129620/U$2 ( \49325 , \47970 , \48858 );
and \g129620/U$3 ( \49326 , \48860 , \47962 );
nor \g129620/U$1 ( \49327 , \49325 , \49326 );
not \g129575/U$4 ( \49328 , \49327 );
or \g129575/U$2 ( \49329 , \49324 , \49328 );
or \g129575/U$5 ( \49330 , \49327 , \48685 );
nand \g129575/U$1 ( \49331 , \49329 , \49330 );
xor \g129496/U$1_r1 ( \49332 , \49323 , \49331 );
not \g129495/U$1 ( \49333 , \49332 );
or \g129134/U$2 ( \49334 , \49314 , \49333 );
and \g129153/U$2 ( \49335 , \49314 , \49333 );
and \g130066/U$2 ( \49336 , \48051 , \48334 );
and \g130066/U$3 ( \49337 , \48335 , \48117 );
nor \g130066/U$1 ( \49338 , \49336 , \49337 );
not \g130024/U$3 ( \49339 , \49338 );
not \g130024/U$4 ( \49340 , \48323 );
and \g130024/U$2 ( \49341 , \49339 , \49340 );
and \g130024/U$5 ( \49342 , \49338 , \48323 );
nor \g130024/U$1 ( \49343 , \49341 , \49342 );
not \g129992/U$3 ( \49344 , \49343 );
and \g130645/U$2 ( \49345 , \48833 , \47913 );
and \g130645/U$3 ( \49346 , \47914 , \48977 );
nor \g130645/U$1 ( \49347 , \49345 , \49346 );
and \g130609/U$2 ( \49348 , \49347 , \47976 );
not \g130609/U$4 ( \49349 , \49347 );
and \g130609/U$3 ( \49350 , \49349 , \47977 );
nor \g130609/U$1 ( \49351 , \49348 , \49350 );
and \g130511/U$2 ( \49352 , \48726 , \47931 );
and \g130511/U$3 ( \49353 , \47930 , \48568 );
nor \g130511/U$1 ( \49354 , \49352 , \49353 );
not \g130480/U$3 ( \49355 , \49354 );
not \g130480/U$4 ( \49356 , \47935 );
and \g130480/U$2 ( \49357 , \49355 , \49356 );
and \g130480/U$5 ( \49358 , \49354 , \47935 );
nor \g130480/U$1 ( \49359 , \49357 , \49358 );
xor \g130431/U$1 ( \49360 , \49351 , \49359 );
not \g129992/U$4 ( \49361 , \49360 );
and \g129992/U$2 ( \49362 , \49344 , \49361 );
and \g129992/U$5 ( \49363 , \49343 , \49360 );
nor \g129992/U$1 ( \49364 , \49362 , \49363 );
and \g130233/U$2 ( \49365 , \48353 , \48155 );
and \g130233/U$3 ( \49366 , \48154 , \48138 );
nor \g130233/U$1 ( \49367 , \49365 , \49366 );
not \g130193/U$3 ( \49368 , \49367 );
not \g130193/U$4 ( \49369 , \48159 );
and \g130193/U$2 ( \49370 , \49368 , \49369 );
and \g130193/U$5 ( \49371 , \49367 , \48159 );
nor \g130193/U$1 ( \49372 , \49370 , \49371 );
and \g130375/U$2 ( \49373 , \48349 , \48063 );
and \g130375/U$3 ( \49374 , \48064 , \48515 );
nor \g130375/U$1 ( \49375 , \49373 , \49374 );
not \g130334/U$3 ( \49376 , \49375 );
not \g130334/U$4 ( \49377 , \47997 );
and \g130334/U$2 ( \49378 , \49376 , \49377 );
and \g130334/U$5 ( \49379 , \49375 , \47997 );
nor \g130334/U$1 ( \49380 , \49378 , \49379 );
xor \g455993/U$9 ( \49381 , \49372 , \49380 );
and \g129712/U$2 ( \49382 , \47950 , \48860 );
and \g129712/U$3 ( \49383 , \48858 , \47962 );
nor \g129712/U$1 ( \49384 , \49382 , \49383 );
not \g129677/U$3 ( \49385 , \49384 );
not \g129677/U$4 ( \49386 , \48685 );
and \g129677/U$2 ( \49387 , \49385 , \49386 );
and \g129677/U$5 ( \49388 , \49384 , \48685 );
nor \g129677/U$1 ( \49389 , \49387 , \49388 );
xor \g455993/U$9_r1 ( \49390 , \49381 , \49389 );
and \g455993/U$8 ( \49391 , \49364 , \49390 );
nand \g130886/U$1 ( \49392 , \40061 , \49282 );
not \g129311/U$3 ( \49393 , \49392 );
not \g129374/U$3 ( \49394 , \49233 );
and \g133210/U$2 ( \49395 , \49231 , \49010 );
not \g133210/U$4 ( \49396 , \49231 );
and \g133210/U$3 ( \49397 , \49396 , \49070 );
nor \g133210/U$1 ( \49398 , \49395 , \49397 );
not \g133352/U$1 ( \49399 , \49229 );
and \g133261/U$2 ( \49400 , \49231 , \49399 );
not \g133261/U$4 ( \49401 , \49231 );
and \g133261/U$3 ( \49402 , \49401 , \49229 );
or \g133261/U$1 ( \49403 , \49400 , \49402 );
not \g133253/U$1 ( \49404 , \49403 );
and \g133190/U$1 ( \49405 , \49398 , \49404 );
nand \g129423/U$1 ( \49406 , \49405 , \47894 );
not \g129374/U$4 ( \49407 , \49406 );
or \g129374/U$2 ( \49408 , \49394 , \49407 );
or \g129374/U$5 ( \49409 , \49406 , \49233 );
nand \g129374/U$1 ( \49410 , \49408 , \49409 );
not \g129311/U$4 ( \49411 , \49410 );
or \g129311/U$2 ( \49412 , \49393 , \49411 );
or \g129311/U$5 ( \49413 , \49410 , \49392 );
nand \g129311/U$1 ( \49414 , \49412 , \49413 );
not \g129294/U$3 ( \49415 , \49414 );
and \g130755/U$2 ( \49416 , \49102 , \47959 );
and \g130755/U$3 ( \49417 , \47960 , \49158 );
nor \g130755/U$1 ( \49418 , \49416 , \49417 );
not \g130729/U$3 ( \49419 , \49418 );
not \g130729/U$4 ( \49420 , \47948 );
and \g130729/U$2 ( \49421 , \49419 , \49420 );
and \g130729/U$5 ( \49422 , \49418 , \47948 );
nor \g130729/U$1 ( \49423 , \49421 , \49422 );
not \g129294/U$4 ( \49424 , \49423 );
and \g129294/U$2 ( \49425 , \49415 , \49424 );
and \g129294/U$5 ( \49426 , \49414 , \49423 );
nor \g129294/U$1 ( \49427 , \49425 , \49426 );
xor \g455993/U$11 ( \49428 , \49372 , \49380 );
xor \g455993/U$11_r1 ( \49429 , \49428 , \49389 );
and \g455993/U$10 ( \49430 , \49427 , \49429 );
and \g455993/U$12 ( \49431 , \49364 , \49427 );
or \g455993/U$7 ( \49432 , \49391 , \49430 , \49431 );
nor \g129153/U$1 ( \49433 , \49335 , \49432 );
not \g129152/U$1 ( \49434 , \49433 );
nand \g129134/U$1 ( \49435 , \49334 , \49434 );
not \g130192/U$3 ( \49436 , \47997 );
and \g130232/U$2 ( \49437 , \48353 , \48064 );
and \g130232/U$3 ( \49438 , \48063 , \48138 );
nor \g130232/U$1 ( \49439 , \49437 , \49438 );
not \g130192/U$4 ( \49440 , \49439 );
or \g130192/U$2 ( \49441 , \49436 , \49440 );
or \g130192/U$5 ( \49442 , \49439 , \47997 );
nand \g130192/U$1 ( \49443 , \49441 , \49442 );
not \g130333/U$3 ( \49444 , \47935 );
and \g130374/U$2 ( \49445 , \48349 , \47930 );
and \g130374/U$3 ( \49446 , \47931 , \48515 );
nor \g130374/U$1 ( \49447 , \49445 , \49446 );
not \g130333/U$4 ( \49448 , \49447 );
or \g130333/U$2 ( \49449 , \49444 , \49448 );
or \g130333/U$5 ( \49450 , \49447 , \47935 );
nand \g130333/U$1 ( \49451 , \49449 , \49450 );
xor \g129405/U$1 ( \49452 , \49443 , \49451 );
not \g129469/U$3 ( \49453 , \48685 );
and \g129512/U$2 ( \49454 , \47970 , \48860 );
and \g129512/U$3 ( \49455 , \48858 , \47972 );
nor \g129512/U$1 ( \49456 , \49454 , \49455 );
not \g129469/U$4 ( \49457 , \49456 );
or \g129469/U$2 ( \49458 , \49453 , \49457 );
or \g129469/U$5 ( \49459 , \49456 , \48685 );
nand \g129469/U$1 ( \49460 , \49458 , \49459 );
xor \g129405/U$1_r1 ( \49461 , \49452 , \49460 );
xor \g129496/U$4 ( \49462 , \49271 , \49322 );
and \g129496/U$3 ( \49463 , \49462 , \49331 );
and \g129496/U$5 ( \49464 , \49271 , \49322 );
or \g129496/U$2 ( \49465 , \49463 , \49464 );
xor \g455975/U$9 ( \49466 , \49461 , \49465 );
xor \g455993/U$5 ( \49467 , \49372 , \49380 );
and \g455993/U$4 ( \49468 , \49467 , \49389 );
and \g455993/U$6 ( \49469 , \49372 , \49380 );
or \g455993/U$3 ( \49470 , \49468 , \49469 );
or \g129985/U$2 ( \49471 , \49359 , \49351 );
and \g130001/U$2 ( \49472 , \49359 , \49351 );
nor \g130001/U$1 ( \49473 , \49472 , \49343 );
not \g130000/U$1 ( \49474 , \49473 );
nand \g129985/U$1 ( \49475 , \49471 , \49474 );
not \g129951/U$1 ( \49476 , \49475 );
or \g129227/U$2 ( \49477 , \49470 , \49476 );
not \g129239/U$3 ( \49478 , \49476 );
not \g129239/U$4 ( \49479 , \49470 );
or \g129239/U$2 ( \49480 , \49478 , \49479 );
or \g129319/U$2 ( \49481 , \49423 , \49392 );
not \g129326/U$3 ( \49482 , \49392 );
not \g129326/U$4 ( \49483 , \49423 );
or \g129326/U$2 ( \49484 , \49482 , \49483 );
nand \g129326/U$1 ( \49485 , \49484 , \49410 );
nand \g129319/U$1 ( \49486 , \49481 , \49485 );
nand \g129239/U$1 ( \49487 , \49480 , \49486 );
nand \g129227/U$1 ( \49488 , \49477 , \49487 );
xor \g455975/U$9_r1 ( \49489 , \49466 , \49488 );
and \g455975/U$8 ( \49490 , \49435 , \49489 );
not \g129213/U$3 ( \49491 , \49486 );
not \g129213/U$4 ( \49492 , \49470 );
and \g129213/U$2 ( \49493 , \49491 , \49492 );
and \g129213/U$5 ( \49494 , \49486 , \49470 );
nor \g129213/U$1 ( \49495 , \49493 , \49494 );
not \g129160/U$3 ( \49496 , \49495 );
not \g129160/U$4 ( \49497 , \49475 );
and \g129160/U$2 ( \49498 , \49496 , \49497 );
and \g129160/U$5 ( \49499 , \49495 , \49475 );
nor \g129160/U$1 ( \49500 , \49498 , \49499 );
and \g130302/U$2 ( \49501 , \48349 , \48155 );
and \g130302/U$3 ( \49502 , \48154 , \48353 );
nor \g130302/U$1 ( \49503 , \49501 , \49502 );
not \g130268/U$3 ( \49504 , \49503 );
not \g130268/U$4 ( \49505 , \48159 );
and \g130268/U$2 ( \49506 , \49504 , \49505 );
and \g130268/U$5 ( \49507 , \49503 , \48159 );
nor \g130268/U$1 ( \49508 , \49506 , \49507 );
and \g130973/U$2 ( \49509 , \42596 , \47649 );
not \g130973/U$4 ( \49510 , \42596 );
and \g130973/U$3 ( \49511 , \49510 , \47650 );
or \g130973/U$1 ( \49512 , \49509 , \49511 );
nand \g130942/U$1 ( \49513 , \40061 , \49512 );
xor \g129497/U$4 ( \49514 , \49508 , \49513 );
and \g129621/U$2 ( \49515 , \47970 , \49074 );
and \g129621/U$3 ( \49516 , \49075 , \47962 );
nor \g129621/U$1 ( \49517 , \49515 , \49516 );
not \g129576/U$3 ( \49518 , \49517 );
not \g129576/U$4 ( \49519 , \49014 );
and \g129576/U$2 ( \49520 , \49518 , \49519 );
and \g129576/U$5 ( \49521 , \49517 , \49014 );
nor \g129576/U$1 ( \49522 , \49520 , \49521 );
and \g129497/U$3 ( \49523 , \49514 , \49522 );
and \g129497/U$5 ( \49524 , \49508 , \49513 );
or \g129497/U$2 ( \49525 , \49523 , \49524 );
and \g130439/U$2 ( \49526 , \48568 , \48064 );
and \g130439/U$3 ( \49527 , \48063 , \48515 );
nor \g130439/U$1 ( \49528 , \49526 , \49527 );
not \g130410/U$3 ( \49529 , \49528 );
not \g130410/U$4 ( \49530 , \47997 );
and \g130410/U$2 ( \49531 , \49529 , \49530 );
and \g130410/U$5 ( \49532 , \49528 , \47997 );
nor \g130410/U$1 ( \49533 , \49531 , \49532 );
and \g130577/U$2 ( \49534 , \48726 , \47930 );
and \g130577/U$3 ( \49535 , \47931 , \48833 );
nor \g130577/U$1 ( \49536 , \49534 , \49535 );
not \g130548/U$3 ( \49537 , \49536 );
not \g130548/U$4 ( \49538 , \47935 );
and \g130548/U$2 ( \49539 , \49537 , \49538 );
and \g130548/U$5 ( \49540 , \49536 , \47935 );
nor \g130548/U$1 ( \49541 , \49539 , \49540 );
xor \g129864/U$4 ( \49542 , \49533 , \49541 );
and \g129973/U$2 ( \49543 , \48051 , \48479 );
and \g129973/U$3 ( \49544 , \48478 , \48018 );
nor \g129973/U$1 ( \49545 , \49543 , \49544 );
not \g129930/U$3 ( \49546 , \49545 );
not \g129930/U$4 ( \49547 , \48483 );
and \g129930/U$2 ( \49548 , \49546 , \49547 );
and \g129930/U$5 ( \49549 , \49545 , \48483 );
nor \g129930/U$1 ( \49550 , \49548 , \49549 );
and \g129864/U$3 ( \49551 , \49542 , \49550 );
and \g129864/U$5 ( \49552 , \49533 , \49541 );
or \g129864/U$2 ( \49553 , \49551 , \49552 );
xor \g129120/U$4 ( \49554 , \49525 , \49553 );
and \g129796/U$2 ( \49555 , \47950 , \48858 );
and \g129796/U$3 ( \49556 , \48860 , \47942 );
nor \g129796/U$1 ( \49557 , \49555 , \49556 );
not \g129750/U$3 ( \49558 , \49557 );
not \g129750/U$4 ( \49559 , \48685 );
and \g129750/U$2 ( \49560 , \49558 , \49559 );
and \g129750/U$5 ( \49561 , \49557 , \48685 );
nor \g129750/U$1 ( \49562 , \49560 , \49561 );
xor \g133476/U$1 ( \49563 , \22092 , \14107 );
xor \g133476/U$1_r1 ( \49564 , \49563 , \39993 );
xor \g133405/U$1 ( \49565 , \21847 , \13864 );
xor \g133405/U$1_r1 ( \49566 , \49565 , \39996 );
nand \g133372/U$1 ( \49567 , \49564 , \49566 );
and \g133313/U$1 ( \49568 , \49229 , \49567 );
xor \g129255/U$4 ( \49569 , \49562 , \49568 );
and \g129396/U$2 ( \49570 , \47894 , \49403 );
and \g129396/U$3 ( \49571 , \49405 , \47972 );
nor \g129396/U$1 ( \49572 , \49570 , \49571 );
not \g129339/U$3 ( \49573 , \49572 );
not \g129339/U$4 ( \49574 , \49233 );
and \g129339/U$2 ( \49575 , \49573 , \49574 );
and \g129339/U$5 ( \49576 , \49572 , \49233 );
nor \g129339/U$1 ( \49577 , \49575 , \49576 );
and \g129255/U$3 ( \49578 , \49569 , \49577 );
and \g129255/U$5 ( \49579 , \49562 , \49568 );
or \g129255/U$2 ( \49580 , \49578 , \49579 );
and \g129120/U$3 ( \49581 , \49554 , \49580 );
and \g129120/U$5 ( \49582 , \49525 , \49553 );
or \g129120/U$2 ( \49583 , \49581 , \49582 );
or \g129050/U$2 ( \49584 , \49500 , \49583 );
not \g129069/U$3 ( \49585 , \49583 );
not \g129069/U$4 ( \49586 , \49500 );
or \g129069/U$2 ( \49587 , \49585 , \49586 );
xor \g456049/U$1 ( \49588 , \49160 , \49168 );
xor \g456049/U$1_r1 ( \49589 , \49588 , \49177 );
not \g129141/U$3 ( \49590 , \49589 );
xor \g129253/U$1 ( \49591 , \49227 , \49233 );
xor \g129253/U$1_r1 ( \49592 , \49591 , \49242 );
not \g129176/U$3 ( \49593 , \49592 );
xor \g456040/U$1 ( \49594 , \49198 , \49206 );
xor \g456040/U$1_r1 ( \49595 , \49594 , \49215 );
not \g129176/U$4 ( \49596 , \49595 );
and \g129176/U$2 ( \49597 , \49593 , \49596 );
and \g129176/U$5 ( \49598 , \49592 , \49595 );
nor \g129176/U$1 ( \49599 , \49597 , \49598 );
not \g129141/U$4 ( \49600 , \49599 );
or \g129141/U$2 ( \49601 , \49590 , \49600 );
or \g129141/U$5 ( \49602 , \49599 , \49589 );
nand \g129141/U$1 ( \49603 , \49601 , \49602 );
nand \g129069/U$1 ( \49604 , \49587 , \49603 );
nand \g129050/U$1 ( \49605 , \49584 , \49604 );
xor \g455975/U$11 ( \49606 , \49461 , \49465 );
xor \g455975/U$11_r1 ( \49607 , \49606 , \49488 );
and \g455975/U$10 ( \49608 , \49605 , \49607 );
and \g455975/U$12 ( \49609 , \49435 , \49605 );
or \g455975/U$7 ( \49610 , \49490 , \49608 , \49609 );
xnor \g128904/U$1 ( \49611 , \49263 , \49610 );
not \g128877/U$3 ( \49612 , \49611 );
xor \g455975/U$5 ( \49613 , \49461 , \49465 );
and \g455975/U$4 ( \49614 , \49613 , \49488 );
and \g455975/U$6 ( \49615 , \49461 , \49465 );
or \g455975/U$3 ( \49616 , \49614 , \49615 );
xor \g129405/U$4 ( \49617 , \49443 , \49451 );
and \g129405/U$3 ( \49618 , \49617 , \49460 );
and \g129405/U$5 ( \49619 , \49443 , \49451 );
or \g129405/U$2 ( \49620 , \49618 , \49619 );
xor \g456039/U$1 ( \49621 , \48957 , \48964 );
xor \g456039/U$1_r1 ( \49622 , \49621 , \48973 );
not \g129212/U$3 ( \49623 , \49622 );
xor \g129273/U$1 ( \49624 , \49035 , \49062 );
xor \g129273/U$1_r1 ( \49625 , \49624 , \49081 );
not \g129212/U$4 ( \49626 , \49625 );
or \g129212/U$2 ( \49627 , \49623 , \49626 );
or \g129212/U$5 ( \49628 , \49625 , \49622 );
nand \g129212/U$1 ( \49629 , \49627 , \49628 );
xor \g455934/U$1 ( \49630 , \49620 , \49629 );
xor \g129000/U$1 ( \49631 , \49616 , \49630 );
not \g128940/U$3 ( \49632 , \49631 );
xor \g129118/U$1 ( \49633 , \49080 , \49218 );
xor \g129118/U$1_r1 ( \49634 , \49633 , \49245 );
not \g129044/U$3 ( \49635 , \49634 );
xor \g456005/U$2 ( \49636 , \49042 , \49050 );
xor \g456005/U$1 ( \49637 , \49636 , \49059 );
xor \g456005/U$1_r1 ( \49638 , \49180 , \49185 );
xor \g456005/U$1_r2 ( \49639 , \49637 , \49638 );
not \g129044/U$4 ( \49640 , \49639 );
and \g129044/U$2 ( \49641 , \49635 , \49640 );
and \g129064/U$2 ( \49642 , \49634 , \49639 );
and \g129183/U$2 ( \49643 , \49595 , \49589 );
not \g129203/U$3 ( \49644 , \49595 );
not \g129203/U$4 ( \49645 , \49589 );
and \g129203/U$2 ( \49646 , \49644 , \49645 );
nor \g129203/U$1 ( \49647 , \49646 , \49592 );
nor \g129183/U$1 ( \49648 , \49643 , \49647 );
nor \g129064/U$1 ( \49649 , \49642 , \49648 );
nor \g129044/U$1 ( \49650 , \49641 , \49649 );
not \g128940/U$4 ( \49651 , \49650 );
or \g128940/U$2 ( \49652 , \49632 , \49651 );
or \g128940/U$5 ( \49653 , \49650 , \49631 );
nand \g128940/U$1 ( \49654 , \49652 , \49653 );
not \g128877/U$4 ( \49655 , \49654 );
and \g128877/U$2 ( \49656 , \49612 , \49655 );
and \g128877/U$5 ( \49657 , \49611 , \49654 );
nor \g128877/U$1 ( \49658 , \49656 , \49657 );
not \g129040/U$3 ( \49659 , \49634 );
xor \g129078/U$1 ( \49660 , \49639 , \49648 );
not \g129040/U$4 ( \49661 , \49660 );
or \g129040/U$2 ( \49662 , \49659 , \49661 );
or \g129040/U$5 ( \49663 , \49660 , \49634 );
nand \g129040/U$1 ( \49664 , \49662 , \49663 );
not \g128870/U$3 ( \49665 , \49664 );
not \g129126/U$3 ( \49666 , \49332 );
not \g129126/U$4 ( \49667 , \49432 );
or \g129126/U$2 ( \49668 , \49666 , \49667 );
or \g129126/U$5 ( \49669 , \49432 , \49332 );
nand \g129126/U$1 ( \49670 , \49668 , \49669 );
not \g129109/U$3 ( \49671 , \49670 );
not \g129109/U$4 ( \49672 , \49314 );
and \g129109/U$2 ( \49673 , \49671 , \49672 );
and \g129109/U$5 ( \49674 , \49670 , \49314 );
nor \g129109/U$1 ( \49675 , \49673 , \49674 );
not \g128956/U$3 ( \49676 , \49675 );
and \g129879/U$2 ( \49677 , \48018 , \48860 );
and \g129879/U$3 ( \49678 , \48858 , \47942 );
nor \g129879/U$1 ( \49679 , \49677 , \49678 );
not \g129846/U$3 ( \49680 , \49679 );
not \g129846/U$4 ( \49681 , \48685 );
and \g129846/U$2 ( \49682 , \49680 , \49681 );
and \g129846/U$5 ( \49683 , \49679 , \48685 );
nor \g129846/U$1 ( \49684 , \49682 , \49683 );
not \g130611/U$3 ( \49685 , \47935 );
and \g130646/U$2 ( \49686 , \48833 , \47930 );
and \g130646/U$3 ( \49687 , \47931 , \48977 );
nor \g130646/U$1 ( \49688 , \49686 , \49687 );
not \g130611/U$4 ( \49689 , \49688 );
or \g130611/U$2 ( \49690 , \49685 , \49689 );
or \g130611/U$5 ( \49691 , \49688 , \47935 );
nand \g130611/U$1 ( \49692 , \49690 , \49691 );
not \g130481/U$3 ( \49693 , \47997 );
and \g130512/U$2 ( \49694 , \48726 , \48064 );
and \g130512/U$3 ( \49695 , \48063 , \48568 );
nor \g130512/U$1 ( \49696 , \49694 , \49695 );
not \g130481/U$4 ( \49697 , \49696 );
or \g130481/U$2 ( \49698 , \49693 , \49697 );
or \g130481/U$5 ( \49699 , \49696 , \47997 );
nand \g130481/U$1 ( \49700 , \49698 , \49699 );
xor \g456046/U$4 ( \49701 , \49692 , \49700 );
not \g130025/U$3 ( \49702 , \48483 );
and \g130067/U$2 ( \49703 , \48051 , \48478 );
and \g130067/U$3 ( \49704 , \48479 , \48117 );
nor \g130067/U$1 ( \49705 , \49703 , \49704 );
not \g130025/U$4 ( \49706 , \49705 );
or \g130025/U$2 ( \49707 , \49702 , \49706 );
or \g130025/U$5 ( \49708 , \49705 , \48483 );
nand \g130025/U$1 ( \49709 , \49707 , \49708 );
and \g456046/U$3 ( \49710 , \49701 , \49709 );
and \g456046/U$5 ( \49711 , \49692 , \49700 );
nor \g456046/U$2 ( \49712 , \49710 , \49711 );
xor \g129482/U$4 ( \49713 , \49684 , \49712 );
xor \g131039/U$1 ( \49714 , \47639 , \47646 );
not \g135519/U$2 ( \49715 , \49714 );
nor \g135519/U$1 ( \49716 , \49715 , \40060 );
not \g130194/U$3 ( \49717 , \48323 );
and \g130234/U$2 ( \49718 , \48353 , \48335 );
and \g130234/U$3 ( \49719 , \48334 , \48138 );
nor \g130234/U$1 ( \49720 , \49718 , \49719 );
not \g130194/U$4 ( \49721 , \49720 );
or \g130194/U$2 ( \49722 , \49717 , \49721 );
or \g130194/U$5 ( \49723 , \49720 , \48323 );
nand \g130194/U$1 ( \49724 , \49722 , \49723 );
xor \g456019/U$4 ( \49725 , \49716 , \49724 );
not \g129678/U$3 ( \49726 , \49014 );
and \g129713/U$2 ( \49727 , \47950 , \49075 );
and \g129713/U$3 ( \49728 , \49074 , \47962 );
nor \g129713/U$1 ( \49729 , \49727 , \49728 );
not \g129678/U$4 ( \49730 , \49729 );
or \g129678/U$2 ( \49731 , \49726 , \49730 );
or \g129678/U$5 ( \49732 , \49729 , \49014 );
nand \g129678/U$1 ( \49733 , \49731 , \49732 );
and \g456019/U$3 ( \49734 , \49725 , \49733 );
and \g456019/U$5 ( \49735 , \49716 , \49724 );
nor \g456019/U$2 ( \49736 , \49734 , \49735 );
and \g129482/U$3 ( \49737 , \49713 , \49736 );
and \g129482/U$5 ( \49738 , \49684 , \49712 );
or \g129482/U$2 ( \49739 , \49737 , \49738 );
xor \g455976/U$9 ( \49740 , \49271 , \49302 );
xor \g455976/U$9_r1 ( \49741 , \49740 , \49311 );
and \g455976/U$8 ( \49742 , \49739 , \49741 );
xor \g129120/U$1 ( \49743 , \49525 , \49553 );
xor \g129120/U$1_r1 ( \49744 , \49743 , \49580 );
xor \g455976/U$11 ( \49745 , \49271 , \49302 );
xor \g455976/U$11_r1 ( \49746 , \49745 , \49311 );
and \g455976/U$10 ( \49747 , \49744 , \49746 );
and \g455976/U$12 ( \49748 , \49739 , \49744 );
or \g455976/U$7 ( \49749 , \49742 , \49747 , \49748 );
not \g128956/U$4 ( \49750 , \49749 );
and \g128956/U$2 ( \49751 , \49676 , \49750 );
and \g128965/U$2 ( \49752 , \49675 , \49749 );
not \g129075/U$3 ( \49753 , \49500 );
not \g129075/U$4 ( \49754 , \49603 );
or \g129075/U$2 ( \49755 , \49753 , \49754 );
or \g129075/U$5 ( \49756 , \49603 , \49500 );
nand \g129075/U$1 ( \49757 , \49755 , \49756 );
not \g129041/U$3 ( \49758 , \49757 );
not \g129041/U$4 ( \49759 , \49583 );
and \g129041/U$2 ( \49760 , \49758 , \49759 );
and \g129041/U$5 ( \49761 , \49757 , \49583 );
nor \g129041/U$1 ( \49762 , \49760 , \49761 );
nor \g128965/U$1 ( \49763 , \49752 , \49762 );
nor \g128956/U$1 ( \49764 , \49751 , \49763 );
not \g128900/U$3 ( \49765 , \49764 );
xor \g455975/U$2 ( \49766 , \49461 , \49465 );
xor \g455975/U$1 ( \49767 , \49766 , \49488 );
xor \g455975/U$1_r1 ( \49768 , \49435 , \49605 );
xor \g455975/U$1_r2 ( \49769 , \49767 , \49768 );
not \g128900/U$4 ( \49770 , \49769 );
and \g128900/U$2 ( \49771 , \49765 , \49770 );
and \g128900/U$5 ( \49772 , \49764 , \49769 );
nor \g128900/U$1 ( \49773 , \49771 , \49772 );
not \g128870/U$4 ( \49774 , \49773 );
or \g128870/U$2 ( \49775 , \49665 , \49774 );
or \g128870/U$5 ( \49776 , \49773 , \49664 );
nand \g128870/U$1 ( \49777 , \49775 , \49776 );
xor \g455993/U$2 ( \49778 , \49372 , \49380 );
xor \g455993/U$1 ( \49779 , \49778 , \49389 );
xor \g455993/U$1_r1 ( \49780 , \49364 , \49427 );
xor \g455993/U$1_r2 ( \49781 , \49779 , \49780 );
xor \g129497/U$1 ( \49782 , \49508 , \49513 );
xor \g129497/U$1_r1 ( \49783 , \49782 , \49522 );
xor \g130043/U$1 ( \49784 , \49278 , \49290 );
xor \g130043/U$1_r1 ( \49785 , \49784 , \49299 );
xor \g455984/U$5 ( \49786 , \49783 , \49785 );
and \g130756/U$2 ( \49787 , \49102 , \47913 );
and \g130756/U$3 ( \49788 , \47914 , \49158 );
nor \g130756/U$1 ( \49789 , \49787 , \49788 );
and \g130730/U$2 ( \49790 , \49789 , \47976 );
not \g130730/U$4 ( \49791 , \49789 );
and \g130730/U$3 ( \49792 , \49791 , \47977 );
nor \g130730/U$1 ( \49793 , \49790 , \49792 );
and \g130867/U$2 ( \49794 , \49512 , \47960 );
and \g130867/U$3 ( \49795 , \47959 , \49282 );
nor \g130867/U$1 ( \49796 , \49794 , \49795 );
not \g130842/U$3 ( \49797 , \49796 );
not \g130842/U$4 ( \49798 , \47948 );
and \g130842/U$2 ( \49799 , \49797 , \49798 );
and \g130842/U$5 ( \49800 , \49796 , \47948 );
nor \g130842/U$1 ( \49801 , \49799 , \49800 );
xor \g129277/U$4 ( \49802 , \49793 , \49801 );
and \g133299/U$2 ( \49803 , \49566 , \49229 );
not \g133299/U$4 ( \49804 , \49566 );
and \g133299/U$3 ( \49805 , \49804 , \49399 );
nor \g133299/U$1 ( \49806 , \49803 , \49805 );
not \g135554/U$2 ( \49807 , \49806 );
not \g133475/U$1 ( \49808 , \49564 );
and \g133357/U$2 ( \49809 , \49566 , \49808 );
not \g133357/U$4 ( \49810 , \49566 );
and \g133357/U$3 ( \49811 , \49810 , \49564 );
or \g133357/U$1 ( \49812 , \49809 , \49811 );
nor \g135554/U$1 ( \49813 , \49807 , \49812 );
nand \g129424/U$1 ( \49814 , \49813 , \47894 );
not \g129375/U$3 ( \49815 , \49814 );
not \g129375/U$4 ( \49816 , \49568 );
and \g129375/U$2 ( \49817 , \49815 , \49816 );
and \g129375/U$5 ( \49818 , \49814 , \49568 );
nor \g129375/U$1 ( \49819 , \49817 , \49818 );
and \g129277/U$3 ( \49820 , \49802 , \49819 );
and \g129277/U$5 ( \49821 , \49793 , \49801 );
or \g129277/U$2 ( \49822 , \49820 , \49821 );
and \g455984/U$4 ( \49823 , \49786 , \49822 );
and \g455984/U$6 ( \49824 , \49783 , \49785 );
or \g455984/U$3 ( \49825 , \49823 , \49824 );
xor \g455974/U$2 ( \49826 , \49781 , \49825 );
not \g129470/U$3 ( \49827 , \49233 );
and \g129513/U$2 ( \49828 , \47970 , \49405 );
and \g129513/U$3 ( \49829 , \49403 , \47972 );
nor \g129513/U$1 ( \49830 , \49828 , \49829 );
not \g129470/U$4 ( \49831 , \49830 );
or \g129470/U$2 ( \49832 , \49827 , \49831 );
or \g129470/U$5 ( \49833 , \49830 , \49233 );
nand \g129470/U$1 ( \49834 , \49832 , \49833 );
not \g130335/U$3 ( \49835 , \48159 );
and \g130376/U$2 ( \49836 , \48349 , \48154 );
and \g130376/U$3 ( \49837 , \48155 , \48515 );
nor \g130376/U$1 ( \49838 , \49836 , \49837 );
not \g130335/U$4 ( \49839 , \49838 );
or \g130335/U$2 ( \49840 , \49835 , \49839 );
or \g130335/U$5 ( \49841 , \49838 , \48159 );
nand \g130335/U$1 ( \49842 , \49840 , \49841 );
not \g129815/U$2 ( \49843 , \49842 );
not \g129845/U$1 ( \49844 , \49684 );
nand \g129815/U$1 ( \49845 , \49843 , \49844 );
and \g129439/U$2 ( \49846 , \49834 , \49845 );
and \g129439/U$3 ( \49847 , \49842 , \49684 );
nor \g129439/U$1 ( \49848 , \49846 , \49847 );
xor \g129864/U$1 ( \49849 , \49533 , \49541 );
xor \g129864/U$1_r1 ( \49850 , \49849 , \49550 );
xor \g129154/U$4 ( \49851 , \49848 , \49850 );
xor \g129255/U$1 ( \49852 , \49562 , \49568 );
xor \g129255/U$1_r1 ( \49853 , \49852 , \49577 );
and \g129154/U$3 ( \49854 , \49851 , \49853 );
and \g129154/U$5 ( \49855 , \49848 , \49850 );
or \g129154/U$2 ( \49856 , \49854 , \49855 );
xor \g455974/U$1 ( \49857 , \49826 , \49856 );
and \g130816/U$2 ( \49858 , \49282 , \47914 );
and \g130816/U$3 ( \49859 , \47913 , \49158 );
nor \g130816/U$1 ( \49860 , \49858 , \49859 );
and \g130785/U$2 ( \49861 , \49860 , \47977 );
not \g130785/U$4 ( \49862 , \49860 );
and \g130785/U$3 ( \49863 , \49862 , \47976 );
nor \g130785/U$1 ( \49864 , \49861 , \49863 );
not \g130675/U$3 ( \49865 , \47935 );
and \g130701/U$2 ( \49866 , \49102 , \47931 );
and \g130701/U$3 ( \49867 , \47930 , \48977 );
nor \g130701/U$1 ( \49868 , \49866 , \49867 );
not \g130675/U$4 ( \49869 , \49868 );
or \g130675/U$2 ( \49870 , \49865 , \49869 );
or \g130675/U$5 ( \49871 , \49868 , \47935 );
nand \g130675/U$1 ( \49872 , \49870 , \49871 );
xor \g456050/U$4 ( \49873 , \49864 , \49872 );
not \g130116/U$3 ( \49874 , \48483 );
and \g130154/U$2 ( \49875 , \48117 , \48478 );
and \g130154/U$3 ( \49876 , \48479 , \48138 );
nor \g130154/U$1 ( \49877 , \49875 , \49876 );
not \g130116/U$4 ( \49878 , \49877 );
or \g130116/U$2 ( \49879 , \49874 , \49878 );
or \g130116/U$5 ( \49880 , \49877 , \48483 );
nand \g130116/U$1 ( \49881 , \49879 , \49880 );
and \g456050/U$3 ( \49882 , \49873 , \49881 );
and \g456050/U$5 ( \49883 , \49864 , \49872 );
nor \g456050/U$2 ( \49884 , \49882 , \49883 );
and \g131117/U$2 ( \49885 , \47635 , \47636 );
not \g131117/U$4 ( \49886 , \47635 );
and \g131117/U$3 ( \49887 , \49886 , \47637 );
or \g131117/U$1 ( \49888 , \49885 , \49887 );
not \g135520/U$2 ( \49889 , \49888 );
nor \g135520/U$1 ( \49890 , \49889 , \40060 );
not \g130897/U$3 ( \49891 , \47948 );
and \g130924/U$2 ( \49892 , \49512 , \47959 );
and \g130924/U$3 ( \49893 , \47960 , \49714 );
nor \g130924/U$1 ( \49894 , \49892 , \49893 );
not \g130897/U$4 ( \49895 , \49894 );
or \g130897/U$2 ( \49896 , \49891 , \49895 );
or \g130897/U$5 ( \49897 , \49894 , \47948 );
nand \g130897/U$1 ( \49898 , \49896 , \49897 );
xor \g456057/U$4 ( \49899 , \49890 , \49898 );
not \g130269/U$3 ( \49900 , \48323 );
and \g130303/U$2 ( \49901 , \48349 , \48335 );
and \g130303/U$3 ( \49902 , \48334 , \48353 );
nor \g130303/U$1 ( \49903 , \49901 , \49902 );
not \g130269/U$4 ( \49904 , \49903 );
or \g130269/U$2 ( \49905 , \49900 , \49904 );
or \g130269/U$5 ( \49906 , \49903 , \48323 );
nand \g130269/U$1 ( \49907 , \49905 , \49906 );
and \g456057/U$3 ( \49908 , \49899 , \49907 );
and \g456057/U$5 ( \49909 , \49890 , \49898 );
nor \g456057/U$2 ( \49910 , \49908 , \49909 );
xor \g129119/U$4 ( \49911 , \49884 , \49910 );
and \g129797/U$2 ( \49912 , \47950 , \49074 );
and \g129797/U$3 ( \49913 , \49075 , \47942 );
nor \g129797/U$1 ( \49914 , \49912 , \49913 );
not \g129751/U$3 ( \49915 , \49914 );
not \g129751/U$4 ( \49916 , \49014 );
and \g129751/U$2 ( \49917 , \49915 , \49916 );
and \g129751/U$5 ( \49918 , \49914 , \49014 );
nor \g129751/U$1 ( \49919 , \49917 , \49918 );
xor \g133630/U$1 ( \49920 , \22585 , \14597 );
xor \g133630/U$1_r1 ( \49921 , \49920 , \39987 );
xor \g133539/U$1 ( \49922 , \22336 , \14354 );
xor \g133539/U$1_r1 ( \49923 , \49922 , \39990 );
nand \g133497/U$1 ( \49924 , \49921 , \49923 );
and \g133432/U$1 ( \49925 , \49564 , \49924 );
xor \g129254/U$4 ( \49926 , \49919 , \49925 );
and \g129397/U$2 ( \49927 , \47894 , \49812 );
and \g129397/U$3 ( \49928 , \49813 , \47972 );
nor \g129397/U$1 ( \49929 , \49927 , \49928 );
not \g129340/U$3 ( \49930 , \49929 );
not \g129340/U$4 ( \49931 , \49568 );
and \g129340/U$2 ( \49932 , \49930 , \49931 );
and \g129340/U$5 ( \49933 , \49929 , \49568 );
nor \g129340/U$1 ( \49934 , \49932 , \49933 );
and \g129254/U$3 ( \49935 , \49926 , \49934 );
and \g129254/U$5 ( \49936 , \49919 , \49925 );
or \g129254/U$2 ( \49937 , \49935 , \49936 );
and \g129119/U$3 ( \49938 , \49911 , \49937 );
and \g129119/U$5 ( \49939 , \49884 , \49910 );
or \g129119/U$2 ( \49940 , \49938 , \49939 );
xor \g129482/U$1 ( \49941 , \49684 , \49712 );
xor \g129482/U$1_r1 ( \49942 , \49941 , \49736 );
xor \g129009/U$4 ( \49943 , \49940 , \49942 );
xor \g456019/U$1 ( \49944 , \49716 , \49724 );
xor \g456019/U$1_r1 ( \49945 , \49944 , \49733 );
not \g130411/U$3 ( \49946 , \48159 );
and \g130440/U$2 ( \49947 , \48568 , \48155 );
and \g130440/U$3 ( \49948 , \48154 , \48515 );
nor \g130440/U$1 ( \49949 , \49947 , \49948 );
not \g130411/U$4 ( \49950 , \49949 );
or \g130411/U$2 ( \49951 , \49946 , \49950 );
or \g130411/U$5 ( \49952 , \49949 , \48159 );
nand \g130411/U$1 ( \49953 , \49951 , \49952 );
not \g130549/U$3 ( \49954 , \47997 );
and \g130578/U$2 ( \49955 , \48726 , \48063 );
and \g130578/U$3 ( \49956 , \48064 , \48833 );
nor \g130578/U$1 ( \49957 , \49955 , \49956 );
not \g130549/U$4 ( \49958 , \49957 );
or \g130549/U$2 ( \49959 , \49954 , \49958 );
or \g130549/U$5 ( \49960 , \49957 , \47997 );
nand \g130549/U$1 ( \49961 , \49959 , \49960 );
xor \g129863/U$4 ( \49962 , \49953 , \49961 );
not \g129931/U$3 ( \49963 , \48685 );
and \g129974/U$2 ( \49964 , \48051 , \48860 );
and \g129974/U$3 ( \49965 , \48858 , \48018 );
nor \g129974/U$1 ( \49966 , \49964 , \49965 );
not \g129931/U$4 ( \49967 , \49966 );
or \g129931/U$2 ( \49968 , \49963 , \49967 );
or \g129931/U$5 ( \49969 , \49966 , \48685 );
nand \g129931/U$1 ( \49970 , \49968 , \49969 );
and \g129863/U$3 ( \49971 , \49962 , \49970 );
and \g129863/U$5 ( \49972 , \49953 , \49961 );
or \g129863/U$2 ( \49973 , \49971 , \49972 );
and \g129228/U$2 ( \49974 , \49945 , \49973 );
not \g129240/U$3 ( \49975 , \49945 );
not \g129240/U$4 ( \49976 , \49973 );
and \g129240/U$2 ( \49977 , \49975 , \49976 );
xor \g129277/U$1 ( \49978 , \49793 , \49801 );
xor \g129277/U$1_r1 ( \49979 , \49978 , \49819 );
nor \g129240/U$1 ( \49980 , \49977 , \49979 );
nor \g129228/U$1 ( \49981 , \49974 , \49980 );
and \g129009/U$3 ( \49982 , \49943 , \49981 );
and \g129009/U$5 ( \49983 , \49940 , \49942 );
or \g129009/U$2 ( \49984 , \49982 , \49983 );
xor \g455976/U$2 ( \49985 , \49271 , \49302 );
xor \g455976/U$1 ( \49986 , \49985 , \49311 );
xor \g455976/U$1_r1 ( \49987 , \49739 , \49744 );
xor \g455976/U$1_r2 ( \49988 , \49986 , \49987 );
xor \g455974/U$1_r1 ( \49989 , \49984 , \49988 );
xor \g455974/U$1_r2 ( \49990 , \49857 , \49989 );
not \g128886/U$3 ( \49991 , \49990 );
not \g130736/U$3 ( \49992 , \47935 );
and \g130761/U$2 ( \49993 , \49102 , \47930 );
and \g130761/U$3 ( \49994 , \47931 , \49158 );
nor \g130761/U$1 ( \49995 , \49993 , \49994 );
not \g130736/U$4 ( \49996 , \49995 );
or \g130736/U$2 ( \49997 , \49992 , \49996 );
or \g130736/U$5 ( \49998 , \49995 , \47935 );
nand \g130736/U$1 ( \49999 , \49997 , \49998 );
and \g130873/U$2 ( \50000 , \49512 , \47914 );
and \g130873/U$3 ( \50001 , \47913 , \49282 );
nor \g130873/U$1 ( \50002 , \50000 , \50001 );
and \g130847/U$2 ( \50003 , \50002 , \47977 );
not \g130847/U$4 ( \50004 , \50002 );
and \g130847/U$3 ( \50005 , \50004 , \47976 );
nor \g130847/U$1 ( \50006 , \50003 , \50005 );
xor \g129956/U$4 ( \50007 , \49999 , \50006 );
not \g130031/U$3 ( \50008 , \48685 );
and \g130073/U$2 ( \50009 , \48051 , \48858 );
and \g130073/U$3 ( \50010 , \48860 , \48117 );
nor \g130073/U$1 ( \50011 , \50009 , \50010 );
not \g130031/U$4 ( \50012 , \50011 );
or \g130031/U$2 ( \50013 , \50008 , \50012 );
or \g130031/U$5 ( \50014 , \50011 , \48685 );
nand \g130031/U$1 ( \50015 , \50013 , \50014 );
and \g129956/U$3 ( \50016 , \50007 , \50015 );
and \g129956/U$5 ( \50017 , \49999 , \50006 );
or \g129956/U$2 ( \50018 , \50016 , \50017 );
xor \g131195/U$1 ( \50019 , \47633 , \43059 );
not \g135521/U$2 ( \50020 , \50019 );
nor \g135521/U$1 ( \50021 , \50020 , \40060 );
xor \g456013/U$4 ( \50022 , \50018 , \50021 );
not \g129584/U$3 ( \50023 , \49233 );
and \g129626/U$2 ( \50024 , \47970 , \49403 );
and \g129626/U$3 ( \50025 , \49405 , \47962 );
nor \g129626/U$1 ( \50026 , \50024 , \50025 );
not \g129584/U$4 ( \50027 , \50026 );
or \g129584/U$2 ( \50028 , \50023 , \50027 );
or \g129584/U$5 ( \50029 , \50026 , \49233 );
nand \g129584/U$1 ( \50030 , \50028 , \50029 );
and \g456013/U$3 ( \50031 , \50022 , \50030 );
and \g456013/U$5 ( \50032 , \50018 , \50021 );
nor \g456013/U$2 ( \50033 , \50031 , \50032 );
not \g129499/U$1 ( \50034 , \50033 );
xor \g456046/U$1 ( \50035 , \49692 , \49700 );
xor \g456046/U$1_r1 ( \50036 , \50035 , \49709 );
and \g129355/U$2 ( \50037 , \50034 , \50036 );
not \g129460/U$2 ( \50038 , \50036 );
nand \g129460/U$1 ( \50039 , \50038 , \50033 );
and \g129787/U$2 ( \50040 , \49844 , \49842 );
nor \g129816/U$1 ( \50041 , \49844 , \49842 );
nor \g129787/U$1 ( \50042 , \50040 , \50041 );
not \g129447/U$3 ( \50043 , \50042 );
not \g129447/U$4 ( \50044 , \49834 );
or \g129447/U$2 ( \50045 , \50043 , \50044 );
or \g129447/U$5 ( \50046 , \49834 , \50042 );
nand \g129447/U$1 ( \50047 , \50045 , \50046 );
and \g129355/U$3 ( \50048 , \50039 , \50047 );
nor \g129355/U$1 ( \50049 , \50037 , \50048 );
xor \g455984/U$9 ( \50050 , \49783 , \49785 );
xor \g455984/U$9_r1 ( \50051 , \50050 , \49822 );
and \g455984/U$8 ( \50052 , \50049 , \50051 );
xor \g129154/U$1 ( \50053 , \49848 , \49850 );
xor \g129154/U$1_r1 ( \50054 , \50053 , \49853 );
xor \g455984/U$11 ( \50055 , \49783 , \49785 );
xor \g455984/U$11_r1 ( \50056 , \50055 , \49822 );
and \g455984/U$10 ( \50057 , \50054 , \50056 );
and \g455984/U$12 ( \50058 , \50049 , \50054 );
or \g455984/U$7 ( \50059 , \50052 , \50057 , \50058 );
not \g128886/U$4 ( \50060 , \50059 );
and \g128886/U$2 ( \50061 , \49991 , \50060 );
and \g128891/U$2 ( \50062 , \49990 , \50059 );
xor \g129009/U$1 ( \50063 , \49940 , \49942 );
xor \g129009/U$1_r1 ( \50064 , \50063 , \49981 );
not \g128953/U$3 ( \50065 , \50064 );
xor \g129863/U$1 ( \50066 , \49953 , \49961 );
xor \g129863/U$1_r1 ( \50067 , \50066 , \49970 );
xor \g456050/U$1 ( \50068 , \49864 , \49872 );
xor \g456050/U$1_r1 ( \50069 , \50068 , \49881 );
and \g129188/U$2 ( \50070 , \50067 , \50069 );
not \g129206/U$3 ( \50071 , \50067 );
not \g129206/U$4 ( \50072 , \50069 );
and \g129206/U$2 ( \50073 , \50071 , \50072 );
xor \g129254/U$1 ( \50074 , \49919 , \49925 );
xor \g129254/U$1_r1 ( \50075 , \50074 , \49934 );
nor \g129206/U$1 ( \50076 , \50073 , \50075 );
nor \g129188/U$1 ( \50077 , \50070 , \50076 );
not \g130202/U$3 ( \50078 , \48483 );
and \g130240/U$2 ( \50079 , \48353 , \48479 );
and \g130240/U$3 ( \50080 , \48478 , \48138 );
nor \g130240/U$1 ( \50081 , \50079 , \50080 );
not \g130202/U$4 ( \50082 , \50081 );
or \g130202/U$2 ( \50083 , \50078 , \50082 );
or \g130202/U$5 ( \50084 , \50081 , \48483 );
nand \g130202/U$1 ( \50085 , \50083 , \50084 );
not \g130959/U$3 ( \50086 , \47948 );
and \g130986/U$2 ( \50087 , \49888 , \47960 );
and \g130986/U$3 ( \50088 , \47959 , \49714 );
nor \g130986/U$1 ( \50089 , \50087 , \50088 );
not \g130959/U$4 ( \50090 , \50089 );
or \g130959/U$2 ( \50091 , \50086 , \50090 );
or \g130959/U$5 ( \50092 , \50089 , \47948 );
nand \g130959/U$1 ( \50093 , \50091 , \50092 );
xor \g455995/U$5 ( \50094 , \50085 , \50093 );
not \g129685/U$3 ( \50095 , \49233 );
and \g129718/U$2 ( \50096 , \47950 , \49405 );
and \g129718/U$3 ( \50097 , \49403 , \47962 );
nor \g129718/U$1 ( \50098 , \50096 , \50097 );
not \g129685/U$4 ( \50099 , \50098 );
or \g129685/U$2 ( \50100 , \50095 , \50099 );
or \g129685/U$5 ( \50101 , \50098 , \49233 );
nand \g129685/U$1 ( \50102 , \50100 , \50101 );
and \g455995/U$4 ( \50103 , \50094 , \50102 );
and \g455995/U$6 ( \50104 , \50085 , \50093 );
or \g455995/U$3 ( \50105 , \50103 , \50104 );
not \g130486/U$3 ( \50106 , \48159 );
and \g130517/U$2 ( \50107 , \48726 , \48155 );
and \g130517/U$3 ( \50108 , \48154 , \48568 );
nor \g130517/U$1 ( \50109 , \50107 , \50108 );
not \g130486/U$4 ( \50110 , \50109 );
or \g130486/U$2 ( \50111 , \50106 , \50110 );
or \g130486/U$5 ( \50112 , \50109 , \48159 );
nand \g130486/U$1 ( \50113 , \50111 , \50112 );
not \g130618/U$3 ( \50114 , \47997 );
and \g130651/U$2 ( \50115 , \48833 , \48063 );
and \g130651/U$3 ( \50116 , \48064 , \48977 );
nor \g130651/U$1 ( \50117 , \50115 , \50116 );
not \g130618/U$4 ( \50118 , \50117 );
or \g130618/U$2 ( \50119 , \50114 , \50118 );
or \g130618/U$5 ( \50120 , \50117 , \47997 );
nand \g130618/U$1 ( \50121 , \50119 , \50120 );
xor \g129777/U$4 ( \50122 , \50113 , \50121 );
not \g129852/U$3 ( \50123 , \49014 );
and \g129885/U$2 ( \50124 , \48018 , \49075 );
and \g129885/U$3 ( \50125 , \49074 , \47942 );
nor \g129885/U$1 ( \50126 , \50124 , \50125 );
not \g129852/U$4 ( \50127 , \50126 );
or \g129852/U$2 ( \50128 , \50123 , \50127 );
or \g129852/U$5 ( \50129 , \50126 , \49014 );
nand \g129852/U$1 ( \50130 , \50128 , \50129 );
and \g129777/U$3 ( \50131 , \50122 , \50130 );
and \g129777/U$5 ( \50132 , \50113 , \50121 );
or \g129777/U$2 ( \50133 , \50131 , \50132 );
and \g129231/U$2 ( \50134 , \50105 , \50133 );
not \g129243/U$3 ( \50135 , \50105 );
not \g129243/U$4 ( \50136 , \50133 );
and \g129243/U$2 ( \50137 , \50135 , \50136 );
and \g130382/U$2 ( \50138 , \48349 , \48334 );
and \g130382/U$3 ( \50139 , \48335 , \48515 );
nor \g130382/U$1 ( \50140 , \50138 , \50139 );
not \g130341/U$3 ( \50141 , \50140 );
not \g130341/U$4 ( \50142 , \48323 );
and \g130341/U$2 ( \50143 , \50141 , \50142 );
and \g130341/U$5 ( \50144 , \50140 , \48323 );
nor \g130341/U$1 ( \50145 , \50143 , \50144 );
not \g129322/U$3 ( \50146 , \50145 );
not \g129322/U$4 ( \50147 , \50021 );
and \g129322/U$2 ( \50148 , \50146 , \50147 );
and \g129329/U$2 ( \50149 , \50145 , \50021 );
and \g133409/U$2 ( \50150 , \49923 , \49564 );
not \g133409/U$4 ( \50151 , \49923 );
and \g133409/U$3 ( \50152 , \50151 , \49808 );
nor \g133409/U$1 ( \50153 , \50150 , \50152 );
not \g135555/U$2 ( \50154 , \50153 );
not \g133629/U$1 ( \50155 , \49921 );
and \g133487/U$2 ( \50156 , \49923 , \50155 );
not \g133487/U$4 ( \50157 , \49923 );
and \g133487/U$3 ( \50158 , \50157 , \49921 );
or \g133487/U$1 ( \50159 , \50156 , \50158 );
nor \g135555/U$1 ( \50160 , \50154 , \50159 );
nand \g129427/U$1 ( \50161 , \50160 , \47894 );
not \g129382/U$3 ( \50162 , \50161 );
not \g129382/U$4 ( \50163 , \49925 );
and \g129382/U$2 ( \50164 , \50162 , \50163 );
and \g129382/U$5 ( \50165 , \50161 , \49925 );
nor \g129382/U$1 ( \50166 , \50164 , \50165 );
nor \g129329/U$1 ( \50167 , \50149 , \50166 );
nor \g129322/U$1 ( \50168 , \50148 , \50167 );
nor \g129243/U$1 ( \50169 , \50137 , \50168 );
nor \g129231/U$1 ( \50170 , \50134 , \50169 );
xor \g129017/U$4 ( \50171 , \50077 , \50170 );
xor \g129119/U$1 ( \50172 , \49884 , \49910 );
xor \g129119/U$1_r1 ( \50173 , \50172 , \49937 );
and \g129017/U$3 ( \50174 , \50171 , \50173 );
and \g129017/U$5 ( \50175 , \50077 , \50170 );
or \g129017/U$2 ( \50176 , \50174 , \50175 );
not \g128953/U$4 ( \50177 , \50176 );
and \g128953/U$2 ( \50178 , \50065 , \50177 );
and \g128962/U$2 ( \50179 , \50064 , \50176 );
xor \g455984/U$2 ( \50180 , \49783 , \49785 );
xor \g455984/U$1 ( \50181 , \50180 , \49822 );
xor \g455984/U$1_r1 ( \50182 , \50049 , \50054 );
xor \g455984/U$1_r2 ( \50183 , \50181 , \50182 );
nor \g128962/U$1 ( \50184 , \50179 , \50183 );
nor \g128953/U$1 ( \50185 , \50178 , \50184 );
nor \g128891/U$1 ( \50186 , \50062 , \50185 );
nor \g128886/U$1 ( \50187 , \50061 , \50186 );
xor \g456013/U$1 ( \50188 , \50018 , \50021 );
xor \g456013/U$1_r1 ( \50189 , \50188 , \50030 );
xor \g456057/U$1 ( \50190 , \49890 , \49898 );
xor \g456057/U$1_r1 ( \50191 , \50190 , \49907 );
xor \g455983/U$5 ( \50192 , \50189 , \50191 );
and \g130446/U$2 ( \50193 , \48568 , \48335 );
and \g130446/U$3 ( \50194 , \48334 , \48515 );
nor \g130446/U$1 ( \50195 , \50193 , \50194 );
not \g130417/U$3 ( \50196 , \50195 );
not \g130417/U$4 ( \50197 , \48323 );
and \g130417/U$2 ( \50198 , \50196 , \50197 );
and \g130417/U$5 ( \50199 , \50195 , \48323 );
nor \g130417/U$1 ( \50200 , \50198 , \50199 );
and \g130583/U$2 ( \50201 , \48726 , \48154 );
and \g130583/U$3 ( \50202 , \48155 , \48833 );
nor \g130583/U$1 ( \50203 , \50201 , \50202 );
not \g130554/U$3 ( \50204 , \50203 );
not \g130554/U$4 ( \50205 , \48159 );
and \g130554/U$2 ( \50206 , \50204 , \50205 );
and \g130554/U$5 ( \50207 , \50203 , \48159 );
nor \g130554/U$1 ( \50208 , \50206 , \50207 );
or \g129722/U$2 ( \50209 , \50200 , \50208 );
and \g129731/U$2 ( \50210 , \50200 , \50208 );
and \g129802/U$2 ( \50211 , \47950 , \49403 );
and \g129802/U$3 ( \50212 , \49405 , \47942 );
nor \g129802/U$1 ( \50213 , \50211 , \50212 );
not \g129757/U$3 ( \50214 , \50213 );
not \g129757/U$4 ( \50215 , \49233 );
and \g129757/U$2 ( \50216 , \50214 , \50215 );
and \g129757/U$5 ( \50217 , \50213 , \49233 );
nor \g129757/U$1 ( \50218 , \50216 , \50217 );
nor \g129731/U$1 ( \50219 , \50210 , \50218 );
not \g129730/U$1 ( \50220 , \50219 );
nand \g129722/U$1 ( \50221 , \50209 , \50220 );
and \g130706/U$2 ( \50222 , \49102 , \48064 );
and \g130706/U$3 ( \50223 , \48063 , \48977 );
nor \g130706/U$1 ( \50224 , \50222 , \50223 );
not \g130681/U$3 ( \50225 , \50224 );
not \g130681/U$4 ( \50226 , \47997 );
and \g130681/U$2 ( \50227 , \50225 , \50226 );
and \g130681/U$5 ( \50228 , \50224 , \47997 );
nor \g130681/U$1 ( \50229 , \50227 , \50228 );
and \g130817/U$2 ( \50230 , \49282 , \47931 );
and \g130817/U$3 ( \50231 , \47930 , \49158 );
nor \g130817/U$1 ( \50232 , \50230 , \50231 );
not \g130791/U$3 ( \50233 , \50232 );
not \g130791/U$4 ( \50234 , \47935 );
and \g130791/U$2 ( \50235 , \50233 , \50234 );
and \g130791/U$5 ( \50236 , \50232 , \47935 );
nor \g130791/U$1 ( \50237 , \50235 , \50236 );
or \g129896/U$2 ( \50238 , \50229 , \50237 );
and \g129912/U$2 ( \50239 , \50229 , \50237 );
and \g129975/U$2 ( \50240 , \48051 , \49075 );
and \g129975/U$3 ( \50241 , \49074 , \48018 );
nor \g129975/U$1 ( \50242 , \50240 , \50241 );
not \g129936/U$3 ( \50243 , \50242 );
not \g129936/U$4 ( \50244 , \49014 );
and \g129936/U$2 ( \50245 , \50243 , \50244 );
and \g129936/U$5 ( \50246 , \50242 , \49014 );
nor \g129936/U$1 ( \50247 , \50245 , \50246 );
nor \g129912/U$1 ( \50248 , \50239 , \50247 );
not \g129911/U$1 ( \50249 , \50248 );
nand \g129896/U$1 ( \50250 , \50238 , \50249 );
xor \g129411/U$4 ( \50251 , \50221 , \50250 );
not \g129477/U$3 ( \50252 , \49568 );
and \g129518/U$2 ( \50253 , \47970 , \49813 );
and \g129518/U$3 ( \50254 , \49812 , \47972 );
nor \g129518/U$1 ( \50255 , \50253 , \50254 );
not \g129477/U$4 ( \50256 , \50255 );
or \g129477/U$2 ( \50257 , \50252 , \50256 );
or \g129477/U$5 ( \50258 , \50255 , \49568 );
nand \g129477/U$1 ( \50259 , \50257 , \50258 );
and \g129411/U$3 ( \50260 , \50251 , \50259 );
and \g129411/U$5 ( \50261 , \50221 , \50250 );
or \g129411/U$2 ( \50262 , \50260 , \50261 );
and \g455983/U$4 ( \50263 , \50192 , \50262 );
and \g455983/U$6 ( \50264 , \50189 , \50191 );
or \g455983/U$3 ( \50265 , \50263 , \50264 );
not \g129307/U$3 ( \50266 , \50036 );
not \g129346/U$3 ( \50267 , \50047 );
not \g129346/U$4 ( \50268 , \50033 );
and \g129346/U$2 ( \50269 , \50267 , \50268 );
and \g129346/U$5 ( \50270 , \50047 , \50033 );
nor \g129346/U$1 ( \50271 , \50269 , \50270 );
not \g129307/U$4 ( \50272 , \50271 );
or \g129307/U$2 ( \50273 , \50266 , \50272 );
or \g129307/U$5 ( \50274 , \50271 , \50036 );
nand \g129307/U$1 ( \50275 , \50273 , \50274 );
xor \g455986/U$1 ( \50276 , \50265 , \50275 );
not \g129219/U$3 ( \50277 , \49945 );
not \g129219/U$4 ( \50278 , \49979 );
or \g129219/U$2 ( \50279 , \50277 , \50278 );
or \g129219/U$5 ( \50280 , \49979 , \49945 );
nand \g129219/U$1 ( \50281 , \50279 , \50280 );
xor \g455936/U$1 ( \50282 , \49973 , \50281 );
xor \g455986/U$1_r1 ( \50283 , \50276 , \50282 );
not \g129163/U$3 ( \50284 , \50133 );
not \g129216/U$3 ( \50285 , \50168 );
not \g129216/U$4 ( \50286 , \50105 );
and \g129216/U$2 ( \50287 , \50285 , \50286 );
and \g129216/U$5 ( \50288 , \50168 , \50105 );
nor \g129216/U$1 ( \50289 , \50287 , \50288 );
not \g129163/U$4 ( \50290 , \50289 );
or \g129163/U$2 ( \50291 , \50284 , \50290 );
or \g129163/U$5 ( \50292 , \50289 , \50133 );
nand \g129163/U$1 ( \50293 , \50291 , \50292 );
and \g130308/U$2 ( \50294 , \48349 , \48479 );
and \g130308/U$3 ( \50295 , \48478 , \48353 );
nor \g130308/U$1 ( \50296 , \50294 , \50295 );
not \g130274/U$3 ( \50297 , \50296 );
not \g130274/U$4 ( \50298 , \48483 );
and \g130274/U$2 ( \50299 , \50297 , \50298 );
and \g130274/U$5 ( \50300 , \50296 , \48483 );
nor \g130274/U$1 ( \50301 , \50299 , \50300 );
and \g131249/U$2 ( \50302 , \47629 , \47630 );
not \g131249/U$4 ( \50303 , \47629 );
and \g131249/U$3 ( \50304 , \50303 , \47631 );
or \g131249/U$1 ( \50305 , \50302 , \50304 );
and \g131138/U$2 ( \50306 , \50305 , \47960 );
and \g131138/U$3 ( \50307 , \47959 , \50019 );
nor \g131138/U$1 ( \50308 , \50306 , \50307 );
not \g131104/U$3 ( \50309 , \50308 );
not \g131104/U$4 ( \50310 , \47948 );
and \g131104/U$2 ( \50311 , \50309 , \50310 );
and \g131104/U$5 ( \50312 , \50308 , \47948 );
nor \g131104/U$1 ( \50313 , \50311 , \50312 );
or \g129533/U$2 ( \50314 , \50301 , \50313 );
and \g129549/U$2 ( \50315 , \50301 , \50313 );
and \g129625/U$2 ( \50316 , \47970 , \49812 );
and \g129625/U$3 ( \50317 , \49813 , \47962 );
nor \g129625/U$1 ( \50318 , \50316 , \50317 );
not \g129583/U$3 ( \50319 , \50318 );
not \g129583/U$4 ( \50320 , \49568 );
and \g129583/U$2 ( \50321 , \50319 , \50320 );
and \g129583/U$5 ( \50322 , \50318 , \49568 );
nor \g129583/U$1 ( \50323 , \50321 , \50322 );
nor \g129549/U$1 ( \50324 , \50315 , \50323 );
not \g129548/U$1 ( \50325 , \50324 );
nand \g129533/U$1 ( \50326 , \50314 , \50325 );
and \g130929/U$2 ( \50327 , \49512 , \47913 );
and \g130929/U$3 ( \50328 , \47914 , \49714 );
nor \g130929/U$1 ( \50329 , \50327 , \50328 );
and \g130901/U$2 ( \50330 , \50329 , \47976 );
not \g130901/U$4 ( \50331 , \50329 );
and \g130901/U$3 ( \50332 , \50331 , \47977 );
nor \g130901/U$1 ( \50333 , \50330 , \50332 );
and \g131065/U$2 ( \50334 , \49888 , \47959 );
and \g131065/U$3 ( \50335 , \47960 , \50019 );
nor \g131065/U$1 ( \50336 , \50334 , \50335 );
not \g131024/U$3 ( \50337 , \50336 );
not \g131024/U$4 ( \50338 , \47948 );
and \g131024/U$2 ( \50339 , \50337 , \50338 );
and \g131024/U$5 ( \50340 , \50336 , \47948 );
nor \g131024/U$1 ( \50341 , \50339 , \50340 );
or \g130082/U$2 ( \50342 , \50333 , \50341 );
and \g130100/U$2 ( \50343 , \50333 , \50341 );
and \g130159/U$2 ( \50344 , \48117 , \48858 );
and \g130159/U$3 ( \50345 , \48860 , \48138 );
nor \g130159/U$1 ( \50346 , \50344 , \50345 );
not \g130121/U$3 ( \50347 , \50346 );
not \g130121/U$4 ( \50348 , \48685 );
and \g130121/U$2 ( \50349 , \50347 , \50348 );
and \g130121/U$5 ( \50350 , \50346 , \48685 );
nor \g130121/U$1 ( \50351 , \50349 , \50350 );
nor \g130100/U$1 ( \50352 , \50343 , \50351 );
not \g130099/U$1 ( \50353 , \50352 );
nand \g130082/U$1 ( \50354 , \50342 , \50353 );
xor \g129125/U$4 ( \50355 , \50326 , \50354 );
nand \g131223/U$1 ( \50356 , \40061 , \50305 );
xor \g133847/U$1 ( \50357 , \23076 , \15087 );
xor \g133847/U$1_r1 ( \50358 , \50357 , \39981 );
xor \g133728/U$1 ( \50359 , \22831 , \14840 );
xor \g133728/U$1_r1 ( \50360 , \50359 , \39984 );
nand \g133660/U$1 ( \50361 , \50358 , \50360 );
and \g133593/U$1 ( \50362 , \49921 , \50361 );
or \g129302/U$2 ( \50363 , \50356 , \50362 );
not \g129308/U$3 ( \50364 , \50362 );
not \g129308/U$4 ( \50365 , \50356 );
or \g129308/U$2 ( \50366 , \50364 , \50365 );
not \g129344/U$3 ( \50367 , \49925 );
and \g129401/U$2 ( \50368 , \47894 , \50159 );
and \g129401/U$3 ( \50369 , \50160 , \47972 );
nor \g129401/U$1 ( \50370 , \50368 , \50369 );
not \g129344/U$4 ( \50371 , \50370 );
or \g129344/U$2 ( \50372 , \50367 , \50371 );
or \g129344/U$5 ( \50373 , \50370 , \49925 );
nand \g129344/U$1 ( \50374 , \50372 , \50373 );
nand \g129308/U$1 ( \50375 , \50366 , \50374 );
nand \g129302/U$1 ( \50376 , \50363 , \50375 );
and \g129125/U$3 ( \50377 , \50355 , \50376 );
and \g129125/U$5 ( \50378 , \50326 , \50354 );
or \g129125/U$2 ( \50379 , \50377 , \50378 );
xor \g455982/U$4 ( \50380 , \50293 , \50379 );
xor \g129956/U$1 ( \50381 , \49999 , \50006 );
xor \g129956/U$1_r1 ( \50382 , \50381 , \50015 );
xor \g455995/U$9 ( \50383 , \50085 , \50093 );
xor \g455995/U$9_r1 ( \50384 , \50383 , \50102 );
and \g455995/U$8 ( \50385 , \50382 , \50384 );
not \g129298/U$3 ( \50386 , \50145 );
xor \g455942/U$1 ( \50387 , \50021 , \50166 );
not \g129298/U$4 ( \50388 , \50387 );
or \g129298/U$2 ( \50389 , \50386 , \50388 );
or \g129298/U$5 ( \50390 , \50387 , \50145 );
nand \g129298/U$1 ( \50391 , \50389 , \50390 );
xor \g455995/U$11 ( \50392 , \50085 , \50093 );
xor \g455995/U$11_r1 ( \50393 , \50392 , \50102 );
and \g455995/U$10 ( \50394 , \50391 , \50393 );
and \g455995/U$12 ( \50395 , \50382 , \50391 );
or \g455995/U$7 ( \50396 , \50385 , \50394 , \50395 );
and \g455982/U$3 ( \50397 , \50380 , \50396 );
and \g455982/U$5 ( \50398 , \50293 , \50379 );
nor \g455982/U$2 ( \50399 , \50397 , \50398 );
not \g129028/U$1 ( \50400 , \50399 );
and \g128984/U$2 ( \50401 , \50283 , \50400 );
not \g128995/U$3 ( \50402 , \50283 );
not \g128995/U$4 ( \50403 , \50400 );
and \g128995/U$2 ( \50404 , \50402 , \50403 );
xor \g129017/U$1 ( \50405 , \50077 , \50170 );
xor \g129017/U$1_r1 ( \50406 , \50405 , \50173 );
nor \g128995/U$1 ( \50407 , \50404 , \50406 );
nor \g128984/U$1 ( \50408 , \50401 , \50407 );
xor \g455986/U$4 ( \50409 , \50265 , \50275 );
and \g455986/U$3 ( \50410 , \50409 , \50282 );
and \g455986/U$5 ( \50411 , \50265 , \50275 );
nor \g455986/U$2 ( \50412 , \50410 , \50411 );
or \g128885/U$2 ( \50413 , \50408 , \50412 );
not \g128890/U$3 ( \50414 , \50412 );
not \g128890/U$4 ( \50415 , \50408 );
or \g128890/U$2 ( \50416 , \50414 , \50415 );
not \g128945/U$3 ( \50417 , \50176 );
xor \g128975/U$1 ( \50418 , \50064 , \50183 );
not \g128945/U$4 ( \50419 , \50418 );
or \g128945/U$2 ( \50420 , \50417 , \50419 );
or \g128945/U$5 ( \50421 , \50418 , \50176 );
nand \g128945/U$1 ( \50422 , \50420 , \50421 );
nand \g128890/U$1 ( \50423 , \50416 , \50422 );
nand \g128885/U$1 ( \50424 , \50413 , \50423 );
not \g128939/U$3 ( \50425 , \50399 );
not \g128974/U$3 ( \50426 , \50283 );
not \g128974/U$4 ( \50427 , \50406 );
or \g128974/U$2 ( \50428 , \50426 , \50427 );
or \g128974/U$5 ( \50429 , \50406 , \50283 );
nand \g128974/U$1 ( \50430 , \50428 , \50429 );
not \g128939/U$4 ( \50431 , \50430 );
or \g128939/U$2 ( \50432 , \50425 , \50431 );
or \g128939/U$5 ( \50433 , \50430 , \50399 );
nand \g128939/U$1 ( \50434 , \50432 , \50433 );
and \g130515/U$2 ( \50435 , \48726 , \48335 );
and \g130515/U$3 ( \50436 , \48334 , \48568 );
nor \g130515/U$1 ( \50437 , \50435 , \50436 );
not \g130484/U$3 ( \50438 , \50437 );
not \g130484/U$4 ( \50439 , \48323 );
and \g130484/U$2 ( \50440 , \50438 , \50439 );
and \g130484/U$5 ( \50441 , \50437 , \48323 );
nor \g130484/U$1 ( \50442 , \50440 , \50441 );
xor \g131307/U$1 ( \50443 , \47627 , \43668 );
nand \g131280/U$1 ( \50444 , \40061 , \50443 );
xor \g455988/U$5 ( \50445 , \50442 , \50444 );
and \g129882/U$2 ( \50446 , \48018 , \49405 );
and \g129882/U$3 ( \50447 , \49403 , \47942 );
nor \g129882/U$1 ( \50448 , \50446 , \50447 );
not \g129849/U$3 ( \50449 , \50448 );
not \g129849/U$4 ( \50450 , \49233 );
and \g129849/U$2 ( \50451 , \50449 , \50450 );
and \g129849/U$5 ( \50452 , \50448 , \49233 );
nor \g129849/U$1 ( \50453 , \50451 , \50452 );
and \g455988/U$4 ( \50454 , \50445 , \50453 );
and \g455988/U$6 ( \50455 , \50442 , \50444 );
or \g455988/U$3 ( \50456 , \50454 , \50455 );
and \g130649/U$2 ( \50457 , \48833 , \48154 );
and \g130649/U$3 ( \50458 , \48155 , \48977 );
nor \g130649/U$1 ( \50459 , \50457 , \50458 );
not \g130614/U$3 ( \50460 , \50459 );
not \g130614/U$4 ( \50461 , \48159 );
and \g130614/U$2 ( \50462 , \50460 , \50461 );
and \g130614/U$5 ( \50463 , \50459 , \48159 );
nor \g130614/U$1 ( \50464 , \50462 , \50463 );
and \g130760/U$2 ( \50465 , \49102 , \48063 );
and \g130760/U$3 ( \50466 , \48064 , \49158 );
nor \g130760/U$1 ( \50467 , \50465 , \50466 );
not \g130733/U$3 ( \50468 , \50467 );
not \g130733/U$4 ( \50469 , \47997 );
and \g130733/U$2 ( \50470 , \50468 , \50469 );
and \g130733/U$5 ( \50471 , \50467 , \47997 );
nor \g130733/U$1 ( \50472 , \50470 , \50471 );
xor \g129955/U$4 ( \50473 , \50464 , \50472 );
and \g130070/U$2 ( \50474 , \48051 , \49074 );
and \g130070/U$3 ( \50475 , \49075 , \48117 );
nor \g130070/U$1 ( \50476 , \50474 , \50475 );
not \g130028/U$3 ( \50477 , \50476 );
not \g130028/U$4 ( \50478 , \49014 );
and \g130028/U$2 ( \50479 , \50477 , \50478 );
and \g130028/U$5 ( \50480 , \50476 , \49014 );
nor \g130028/U$1 ( \50481 , \50479 , \50480 );
and \g129955/U$3 ( \50482 , \50473 , \50481 );
and \g129955/U$5 ( \50483 , \50464 , \50472 );
or \g129955/U$2 ( \50484 , \50482 , \50483 );
xor \g129527/U$4 ( \50485 , \50456 , \50484 );
and \g130870/U$2 ( \50486 , \49512 , \47931 );
and \g130870/U$3 ( \50487 , \47930 , \49282 );
nor \g130870/U$1 ( \50488 , \50486 , \50487 );
not \g130844/U$3 ( \50489 , \50488 );
not \g130844/U$4 ( \50490 , \47935 );
and \g130844/U$2 ( \50491 , \50489 , \50490 );
and \g130844/U$5 ( \50492 , \50488 , \47935 );
nor \g130844/U$1 ( \50493 , \50491 , \50492 );
and \g130983/U$2 ( \50494 , \49888 , \47914 );
and \g130983/U$3 ( \50495 , \47913 , \49714 );
nor \g130983/U$1 ( \50496 , \50494 , \50495 );
and \g130955/U$2 ( \50497 , \50496 , \47976 );
not \g130955/U$4 ( \50498 , \50496 );
and \g130955/U$3 ( \50499 , \50498 , \47977 );
nor \g130955/U$1 ( \50500 , \50497 , \50499 );
xor \g455998/U$5 ( \50501 , \50493 , \50500 );
and \g129715/U$2 ( \50502 , \47950 , \49813 );
and \g129715/U$3 ( \50503 , \49812 , \47962 );
nor \g129715/U$1 ( \50504 , \50502 , \50503 );
not \g129680/U$3 ( \50505 , \50504 );
not \g129680/U$4 ( \50506 , \49568 );
and \g129680/U$2 ( \50507 , \50505 , \50506 );
and \g129680/U$5 ( \50508 , \50504 , \49568 );
nor \g129680/U$1 ( \50509 , \50507 , \50508 );
and \g455998/U$4 ( \50510 , \50501 , \50509 );
and \g455998/U$6 ( \50511 , \50493 , \50500 );
or \g455998/U$3 ( \50512 , \50510 , \50511 );
and \g129527/U$3 ( \50513 , \50485 , \50512 );
and \g129527/U$5 ( \50514 , \50456 , \50484 );
or \g129527/U$2 ( \50515 , \50513 , \50514 );
xor \g129777/U$1 ( \50516 , \50113 , \50121 );
xor \g129777/U$1_r1 ( \50517 , \50516 , \50130 );
not \g129776/U$1 ( \50518 , \50517 );
or \g129354/U$2 ( \50519 , \50515 , \50518 );
not \g129359/U$3 ( \50520 , \50518 );
not \g129359/U$4 ( \50521 , \50515 );
or \g129359/U$2 ( \50522 , \50520 , \50521 );
xor \g129411/U$1 ( \50523 , \50221 , \50250 );
xor \g129411/U$1_r1 ( \50524 , \50523 , \50259 );
nand \g129359/U$1 ( \50525 , \50522 , \50524 );
nand \g129354/U$1 ( \50526 , \50519 , \50525 );
xor \g455983/U$9 ( \50527 , \50189 , \50191 );
xor \g455983/U$9_r1 ( \50528 , \50527 , \50262 );
and \g455983/U$8 ( \50529 , \50526 , \50528 );
not \g129146/U$3 ( \50530 , \50069 );
not \g129179/U$3 ( \50531 , \50075 );
not \g129179/U$4 ( \50532 , \50067 );
and \g129179/U$2 ( \50533 , \50531 , \50532 );
and \g129179/U$5 ( \50534 , \50075 , \50067 );
nor \g129179/U$1 ( \50535 , \50533 , \50534 );
not \g129146/U$4 ( \50536 , \50535 );
or \g129146/U$2 ( \50537 , \50530 , \50536 );
or \g129146/U$5 ( \50538 , \50535 , \50069 );
nand \g129146/U$1 ( \50539 , \50537 , \50538 );
xor \g455983/U$11 ( \50540 , \50189 , \50191 );
xor \g455983/U$11_r1 ( \50541 , \50540 , \50262 );
and \g455983/U$10 ( \50542 , \50539 , \50541 );
and \g455983/U$12 ( \50543 , \50526 , \50539 );
or \g455983/U$7 ( \50544 , \50529 , \50542 , \50543 );
and \g128856/U$2 ( \50545 , \50434 , \50544 );
not \g128864/U$3 ( \50546 , \50434 );
not \g128864/U$4 ( \50547 , \50544 );
and \g128864/U$2 ( \50548 , \50546 , \50547 );
xor \g455982/U$1 ( \50549 , \50293 , \50379 );
xor \g455982/U$1_r1 ( \50550 , \50549 , \50396 );
xor \g455995/U$2 ( \50551 , \50085 , \50093 );
xor \g455995/U$1 ( \50552 , \50551 , \50102 );
xor \g455995/U$1_r1 ( \50553 , \50382 , \50391 );
xor \g455995/U$1_r2 ( \50554 , \50552 , \50553 );
not \g129048/U$3 ( \50555 , \50554 );
xor \g129125/U$1 ( \50556 , \50326 , \50354 );
xor \g129125/U$1_r1 ( \50557 , \50556 , \50376 );
not \g129048/U$4 ( \50558 , \50557 );
or \g129048/U$2 ( \50559 , \50555 , \50558 );
or \g129068/U$2 ( \50560 , \50557 , \50554 );
and \g130236/U$2 ( \50561 , \48353 , \48860 );
and \g130236/U$3 ( \50562 , \48858 , \48138 );
nor \g130236/U$1 ( \50563 , \50561 , \50562 );
not \g130196/U$3 ( \50564 , \50563 );
not \g130196/U$4 ( \50565 , \48685 );
and \g130196/U$2 ( \50566 , \50564 , \50565 );
and \g130196/U$5 ( \50567 , \50563 , \48685 );
nor \g130196/U$1 ( \50568 , \50566 , \50567 );
and \g130378/U$2 ( \50569 , \48349 , \48478 );
and \g130378/U$3 ( \50570 , \48479 , \48515 );
nor \g130378/U$1 ( \50571 , \50569 , \50570 );
not \g130337/U$3 ( \50572 , \50571 );
not \g130337/U$4 ( \50573 , \48483 );
and \g130337/U$2 ( \50574 , \50572 , \50573 );
and \g130337/U$5 ( \50575 , \50571 , \48483 );
nor \g130337/U$1 ( \50576 , \50574 , \50575 );
xor \g129280/U$4 ( \50577 , \50568 , \50576 );
and \g133558/U$2 ( \50578 , \50360 , \49921 );
not \g133558/U$4 ( \50579 , \50360 );
and \g133558/U$3 ( \50580 , \50579 , \50155 );
nor \g133558/U$1 ( \50581 , \50578 , \50580 );
not \g135558/U$2 ( \50582 , \50581 );
not \g133846/U$1 ( \50583 , \50358 );
and \g133645/U$2 ( \50584 , \50360 , \50583 );
not \g133645/U$4 ( \50585 , \50360 );
and \g133645/U$3 ( \50586 , \50585 , \50358 );
or \g133645/U$1 ( \50587 , \50584 , \50586 );
nor \g135558/U$1 ( \50588 , \50582 , \50587 );
nand \g129426/U$1 ( \50589 , \50588 , \47894 );
not \g129377/U$3 ( \50590 , \50589 );
not \g129377/U$4 ( \50591 , \50362 );
and \g129377/U$2 ( \50592 , \50590 , \50591 );
and \g129377/U$5 ( \50593 , \50589 , \50362 );
nor \g129377/U$1 ( \50594 , \50592 , \50593 );
and \g129280/U$3 ( \50595 , \50577 , \50594 );
and \g129280/U$5 ( \50596 , \50568 , \50576 );
or \g129280/U$2 ( \50597 , \50595 , \50596 );
not \g129725/U$3 ( \50598 , \50218 );
xor \g130370/U$1 ( \50599 , \50208 , \50200 );
not \g129725/U$4 ( \50600 , \50599 );
and \g129725/U$2 ( \50601 , \50598 , \50600 );
and \g129725/U$5 ( \50602 , \50218 , \50599 );
nor \g129725/U$1 ( \50603 , \50601 , \50602 );
or \g129128/U$2 ( \50604 , \50597 , \50603 );
and \g129149/U$2 ( \50605 , \50597 , \50603 );
not \g129300/U$3 ( \50606 , \50362 );
not \g129300/U$4 ( \50607 , \50374 );
or \g129300/U$2 ( \50608 , \50606 , \50607 );
or \g129300/U$5 ( \50609 , \50374 , \50362 );
nand \g129300/U$1 ( \50610 , \50608 , \50609 );
not \g129271/U$3 ( \50611 , \50610 );
not \g129271/U$4 ( \50612 , \50356 );
and \g129271/U$2 ( \50613 , \50611 , \50612 );
and \g129271/U$5 ( \50614 , \50610 , \50356 );
nor \g129271/U$1 ( \50615 , \50613 , \50614 );
nor \g129149/U$1 ( \50616 , \50605 , \50615 );
not \g129148/U$1 ( \50617 , \50616 );
nand \g129128/U$1 ( \50618 , \50604 , \50617 );
nand \g129068/U$1 ( \50619 , \50560 , \50618 );
nand \g129048/U$1 ( \50620 , \50559 , \50619 );
and \g128907/U$2 ( \50621 , \50550 , \50620 );
not \g128916/U$3 ( \50622 , \50550 );
not \g128916/U$4 ( \50623 , \50620 );
and \g128916/U$2 ( \50624 , \50622 , \50623 );
not \g129347/U$3 ( \50625 , \50524 );
not \g129347/U$4 ( \50626 , \50515 );
and \g129347/U$2 ( \50627 , \50625 , \50626 );
and \g129347/U$5 ( \50628 , \50524 , \50515 );
nor \g129347/U$1 ( \50629 , \50627 , \50628 );
not \g129306/U$3 ( \50630 , \50629 );
not \g129306/U$4 ( \50631 , \50517 );
and \g129306/U$2 ( \50632 , \50630 , \50631 );
and \g129306/U$5 ( \50633 , \50629 , \50517 );
nor \g129306/U$1 ( \50634 , \50632 , \50633 );
not \g129899/U$3 ( \50635 , \50247 );
xor \g130638/U$1 ( \50636 , \50237 , \50229 );
not \g129899/U$4 ( \50637 , \50636 );
and \g129899/U$2 ( \50638 , \50635 , \50637 );
and \g129899/U$5 ( \50639 , \50247 , \50636 );
nor \g129899/U$1 ( \50640 , \50638 , \50639 );
not \g130091/U$3 ( \50641 , \50351 );
xor \g130864/U$1 ( \50642 , \50341 , \50333 );
not \g130091/U$4 ( \50643 , \50642 );
and \g130091/U$2 ( \50644 , \50641 , \50643 );
and \g130091/U$5 ( \50645 , \50351 , \50642 );
nor \g130091/U$1 ( \50646 , \50644 , \50645 );
xor \g129385/U$4 ( \50647 , \50640 , \50646 );
not \g129539/U$3 ( \50648 , \50323 );
and \g130225/U$2 ( \50649 , \50301 , \50313 );
not \g130225/U$4 ( \50650 , \50301 );
not \g131103/U$1 ( \50651 , \50313 );
and \g130225/U$3 ( \50652 , \50650 , \50651 );
nor \g130225/U$1 ( \50653 , \50649 , \50652 );
not \g129539/U$4 ( \50654 , \50653 );
and \g129539/U$2 ( \50655 , \50648 , \50654 );
and \g129539/U$5 ( \50656 , \50323 , \50653 );
nor \g129539/U$1 ( \50657 , \50655 , \50656 );
and \g129385/U$3 ( \50658 , \50647 , \50657 );
and \g129385/U$5 ( \50659 , \50640 , \50646 );
or \g129385/U$2 ( \50660 , \50658 , \50659 );
xor \g128930/U$4 ( \50661 , \50634 , \50660 );
and \g130580/U$2 ( \50662 , \48726 , \48334 );
and \g130580/U$3 ( \50663 , \48335 , \48833 );
nor \g130580/U$1 ( \50664 , \50662 , \50663 );
not \g130551/U$3 ( \50665 , \50664 );
not \g130551/U$4 ( \50666 , \48323 );
and \g130551/U$2 ( \50667 , \50665 , \50666 );
and \g130551/U$5 ( \50668 , \50664 , \48323 );
nor \g130551/U$1 ( \50669 , \50667 , \50668 );
and \g130703/U$2 ( \50670 , \49102 , \48155 );
and \g130703/U$3 ( \50671 , \48154 , \48977 );
nor \g130703/U$1 ( \50672 , \50670 , \50671 );
not \g130677/U$3 ( \50673 , \50672 );
not \g130677/U$4 ( \50674 , \48159 );
and \g130677/U$2 ( \50675 , \50673 , \50674 );
and \g130677/U$5 ( \50676 , \50672 , \48159 );
nor \g130677/U$1 ( \50677 , \50675 , \50676 );
xor \g129866/U$4 ( \50678 , \50669 , \50677 );
and \g129977/U$2 ( \50679 , \48051 , \49405 );
and \g129977/U$3 ( \50680 , \49403 , \48018 );
nor \g129977/U$1 ( \50681 , \50679 , \50680 );
not \g129933/U$3 ( \50682 , \50681 );
not \g129933/U$4 ( \50683 , \49233 );
and \g129933/U$2 ( \50684 , \50682 , \50683 );
and \g129933/U$5 ( \50685 , \50681 , \49233 );
nor \g129933/U$1 ( \50686 , \50684 , \50685 );
and \g129866/U$3 ( \50687 , \50678 , \50686 );
and \g129866/U$5 ( \50688 , \50669 , \50677 );
or \g129866/U$2 ( \50689 , \50687 , \50688 );
and \g130925/U$2 ( \50690 , \49512 , \47930 );
and \g130925/U$3 ( \50691 , \47931 , \49714 );
nor \g130925/U$1 ( \50692 , \50690 , \50691 );
not \g130898/U$3 ( \50693 , \50692 );
not \g130898/U$4 ( \50694 , \47935 );
and \g130898/U$2 ( \50695 , \50693 , \50694 );
and \g130898/U$5 ( \50696 , \50692 , \47935 );
nor \g130898/U$1 ( \50697 , \50695 , \50696 );
and \g131060/U$2 ( \50698 , \49888 , \47913 );
and \g131060/U$3 ( \50699 , \47914 , \50019 );
nor \g131060/U$1 ( \50700 , \50698 , \50699 );
and \g131019/U$2 ( \50701 , \50700 , \47976 );
not \g131019/U$4 ( \50702 , \50700 );
and \g131019/U$3 ( \50703 , \50702 , \47977 );
nor \g131019/U$1 ( \50704 , \50701 , \50703 );
xor \g130748/U$4 ( \50705 , \50697 , \50704 );
and \g130814/U$2 ( \50706 , \49282 , \48064 );
and \g130814/U$3 ( \50707 , \48063 , \49158 );
nor \g130814/U$1 ( \50708 , \50706 , \50707 );
not \g130786/U$3 ( \50709 , \50708 );
not \g130786/U$4 ( \50710 , \47997 );
and \g130786/U$2 ( \50711 , \50709 , \50710 );
and \g130786/U$5 ( \50712 , \50708 , \47997 );
nor \g130786/U$1 ( \50713 , \50711 , \50712 );
and \g130748/U$3 ( \50714 , \50705 , \50713 );
and \g130748/U$5 ( \50715 , \50697 , \50704 );
or \g130748/U$2 ( \50716 , \50714 , \50715 );
xor \g129124/U$4 ( \50717 , \50689 , \50716 );
and \g129799/U$2 ( \50718 , \47950 , \49812 );
and \g129799/U$3 ( \50719 , \49813 , \47942 );
nor \g129799/U$1 ( \50720 , \50718 , \50719 );
not \g129753/U$3 ( \50721 , \50720 );
not \g129753/U$4 ( \50722 , \49568 );
and \g129753/U$2 ( \50723 , \50721 , \50722 );
and \g129753/U$5 ( \50724 , \50720 , \49568 );
nor \g129753/U$1 ( \50725 , \50723 , \50724 );
and \g130442/U$2 ( \50726 , \48568 , \48479 );
and \g130442/U$3 ( \50727 , \48478 , \48515 );
nor \g130442/U$1 ( \50728 , \50726 , \50727 );
not \g130413/U$3 ( \50729 , \50728 );
not \g130413/U$4 ( \50730 , \48483 );
and \g130413/U$2 ( \50731 , \50729 , \50730 );
and \g130413/U$5 ( \50732 , \50728 , \48483 );
nor \g130413/U$1 ( \50733 , \50731 , \50732 );
xor \g455977/U$5 ( \50734 , \50725 , \50733 );
and \g129399/U$2 ( \50735 , \47894 , \50587 );
and \g129399/U$3 ( \50736 , \50588 , \47972 );
nor \g129399/U$1 ( \50737 , \50735 , \50736 );
not \g129342/U$3 ( \50738 , \50737 );
not \g129342/U$4 ( \50739 , \50362 );
and \g129342/U$2 ( \50740 , \50738 , \50739 );
and \g129342/U$5 ( \50741 , \50737 , \50362 );
nor \g129342/U$1 ( \50742 , \50740 , \50741 );
and \g455977/U$4 ( \50743 , \50734 , \50742 );
and \g455977/U$6 ( \50744 , \50725 , \50733 );
or \g455977/U$3 ( \50745 , \50743 , \50744 );
and \g129124/U$3 ( \50746 , \50717 , \50745 );
and \g129124/U$5 ( \50747 , \50689 , \50716 );
or \g129124/U$2 ( \50748 , \50746 , \50747 );
and \g131365/U$2 ( \50749 , \47623 , \47624 );
not \g131365/U$4 ( \50750 , \47623 );
and \g131365/U$3 ( \50751 , \50750 , \47625 );
or \g131365/U$1 ( \50752 , \50749 , \50751 );
nand \g131336/U$1 ( \50753 , \40061 , \50752 );
xor \g134140/U$1 ( \50754 , \23562 , \15573 );
xor \g134140/U$1_r1 ( \50755 , \50754 , \39975 );
xor \g134037/U$1 ( \50756 , \23318 , \15330 );
xor \g134037/U$1_r1 ( \50757 , \50756 , \39978 );
nand \g133882/U$1 ( \50758 , \50755 , \50757 );
and \g133815/U$1 ( \50759 , \50358 , \50758 );
xor \g131122/U$4 ( \50760 , \50753 , \50759 );
and \g131209/U$2 ( \50761 , \50305 , \47959 );
and \g131209/U$3 ( \50762 , \47960 , \50443 );
nor \g131209/U$1 ( \50763 , \50761 , \50762 );
not \g131180/U$3 ( \50764 , \50763 );
not \g131180/U$4 ( \50765 , \47948 );
and \g131180/U$2 ( \50766 , \50764 , \50765 );
and \g131180/U$5 ( \50767 , \50763 , \47948 );
nor \g131180/U$1 ( \50768 , \50766 , \50767 );
and \g131122/U$3 ( \50769 , \50760 , \50768 );
and \g131122/U$5 ( \50770 , \50753 , \50759 );
or \g131122/U$2 ( \50771 , \50769 , \50770 );
xor \g129410/U$4 ( \50772 , \50651 , \50771 );
and \g129516/U$2 ( \50773 , \47970 , \50160 );
and \g129516/U$3 ( \50774 , \50159 , \47972 );
nor \g129516/U$1 ( \50775 , \50773 , \50774 );
not \g129473/U$3 ( \50776 , \50775 );
not \g129473/U$4 ( \50777 , \49925 );
and \g129473/U$2 ( \50778 , \50776 , \50777 );
and \g129473/U$5 ( \50779 , \50775 , \49925 );
nor \g129473/U$1 ( \50780 , \50778 , \50779 );
and \g129410/U$3 ( \50781 , \50772 , \50780 );
and \g129410/U$5 ( \50782 , \50651 , \50771 );
or \g129410/U$2 ( \50783 , \50781 , \50782 );
xor \g129016/U$4 ( \50784 , \50748 , \50783 );
not \g129144/U$3 ( \50785 , \50615 );
xor \g129218/U$1 ( \50786 , \50603 , \50597 );
not \g129144/U$4 ( \50787 , \50786 );
and \g129144/U$2 ( \50788 , \50785 , \50787 );
and \g129144/U$5 ( \50789 , \50615 , \50786 );
nor \g129144/U$1 ( \50790 , \50788 , \50789 );
and \g129016/U$3 ( \50791 , \50784 , \50790 );
and \g129016/U$5 ( \50792 , \50748 , \50783 );
or \g129016/U$2 ( \50793 , \50791 , \50792 );
and \g128930/U$3 ( \50794 , \50661 , \50793 );
and \g128930/U$5 ( \50795 , \50634 , \50660 );
or \g128930/U$2 ( \50796 , \50794 , \50795 );
nor \g128916/U$1 ( \50797 , \50624 , \50796 );
nor \g128907/U$1 ( \50798 , \50621 , \50797 );
nor \g128864/U$1 ( \50799 , \50548 , \50798 );
nor \g128856/U$1 ( \50800 , \50545 , \50799 );
not \g128855/U$3 ( \50801 , \50798 );
not \g128855/U$4 ( \50802 , \50434 );
or \g128855/U$2 ( \50803 , \50801 , \50802 );
or \g128855/U$5 ( \50804 , \50434 , \50798 );
nand \g128855/U$1 ( \50805 , \50803 , \50804 );
xor \g455929/U$1 ( \50806 , \50544 , \50805 );
xor \g455983/U$2 ( \50807 , \50189 , \50191 );
xor \g455983/U$1 ( \50808 , \50807 , \50262 );
xor \g455983/U$1_r1 ( \50809 , \50526 , \50539 );
xor \g455983/U$1_r2 ( \50810 , \50808 , \50809 );
not \g128845/U$3 ( \50811 , \50810 );
not \g128912/U$3 ( \50812 , \50796 );
xor \g128977/U$1 ( \50813 , \50620 , \50550 );
not \g128912/U$4 ( \50814 , \50813 );
or \g128912/U$2 ( \50815 , \50812 , \50814 );
or \g128912/U$5 ( \50816 , \50813 , \50796 );
nand \g128912/U$1 ( \50817 , \50815 , \50816 );
not \g128845/U$4 ( \50818 , \50817 );
or \g128845/U$2 ( \50819 , \50811 , \50818 );
or \g128849/U$2 ( \50820 , \50817 , \50810 );
xnor \g129077/U$1 ( \50821 , \50554 , \50618 );
not \g129039/U$3 ( \50822 , \50821 );
not \g129039/U$4 ( \50823 , \50557 );
and \g129039/U$2 ( \50824 , \50822 , \50823 );
and \g129039/U$5 ( \50825 , \50821 , \50557 );
nor \g129039/U$1 ( \50826 , \50824 , \50825 );
xor \g129955/U$1 ( \50827 , \50464 , \50472 );
xor \g129955/U$1_r1 ( \50828 , \50827 , \50481 );
xor \g455998/U$9 ( \50829 , \50493 , \50500 );
xor \g455998/U$9_r1 ( \50830 , \50829 , \50509 );
and \g455998/U$8 ( \50831 , \50828 , \50830 );
xor \g129410/U$1 ( \50832 , \50651 , \50771 );
xor \g129410/U$1_r1 ( \50833 , \50832 , \50780 );
xor \g455998/U$11 ( \50834 , \50493 , \50500 );
xor \g455998/U$11_r1 ( \50835 , \50834 , \50509 );
and \g455998/U$10 ( \50836 , \50833 , \50835 );
and \g455998/U$12 ( \50837 , \50828 , \50833 );
or \g455998/U$7 ( \50838 , \50831 , \50836 , \50837 );
xor \g129527/U$1 ( \50839 , \50456 , \50484 );
xor \g129527/U$1_r1 ( \50840 , \50839 , \50512 );
xor \g455970/U$5 ( \50841 , \50838 , \50840 );
and \g130304/U$2 ( \50842 , \48349 , \48860 );
and \g130304/U$3 ( \50843 , \48858 , \48353 );
nor \g130304/U$1 ( \50844 , \50842 , \50843 );
not \g130270/U$3 ( \50845 , \50844 );
not \g130270/U$4 ( \50846 , \48685 );
and \g130270/U$2 ( \50847 , \50845 , \50846 );
and \g130270/U$5 ( \50848 , \50844 , \48685 );
nor \g130270/U$1 ( \50849 , \50847 , \50848 );
and \g131137/U$2 ( \50850 , \50305 , \47914 );
and \g131137/U$3 ( \50851 , \47913 , \50019 );
nor \g131137/U$1 ( \50852 , \50850 , \50851 );
and \g131102/U$2 ( \50853 , \50852 , \47977 );
not \g131102/U$4 ( \50854 , \50852 );
and \g131102/U$3 ( \50855 , \50854 , \47976 );
nor \g131102/U$1 ( \50856 , \50853 , \50855 );
not \g131101/U$1 ( \50857 , \50856 );
xor \g455994/U$5 ( \50858 , \50849 , \50857 );
and \g130156/U$2 ( \50859 , \48117 , \49074 );
and \g130156/U$3 ( \50860 , \49075 , \48138 );
nor \g130156/U$1 ( \50861 , \50859 , \50860 );
not \g130118/U$3 ( \50862 , \50861 );
not \g130118/U$4 ( \50863 , \49014 );
and \g130118/U$2 ( \50864 , \50862 , \50863 );
and \g130118/U$5 ( \50865 , \50861 , \49014 );
nor \g130118/U$1 ( \50866 , \50864 , \50865 );
and \g455994/U$4 ( \50867 , \50858 , \50866 );
and \g455994/U$6 ( \50868 , \50849 , \50857 );
or \g455994/U$3 ( \50869 , \50867 , \50868 );
xor \g455988/U$9 ( \50870 , \50442 , \50444 );
xor \g455988/U$9_r1 ( \50871 , \50870 , \50453 );
and \g455988/U$8 ( \50872 , \50869 , \50871 );
xor \g129280/U$1 ( \50873 , \50568 , \50576 );
xor \g129280/U$1_r1 ( \50874 , \50873 , \50594 );
xor \g455988/U$11 ( \50875 , \50442 , \50444 );
xor \g455988/U$11_r1 ( \50876 , \50875 , \50453 );
and \g455988/U$10 ( \50877 , \50874 , \50876 );
and \g455988/U$12 ( \50878 , \50869 , \50874 );
or \g455988/U$7 ( \50879 , \50872 , \50877 , \50878 );
and \g455970/U$4 ( \50880 , \50841 , \50879 );
and \g455970/U$6 ( \50881 , \50838 , \50840 );
or \g455970/U$3 ( \50882 , \50880 , \50881 );
xor \g128861/U$4 ( \50883 , \50826 , \50882 );
and \g130377/U$2 ( \50884 , \48349 , \48858 );
and \g130377/U$3 ( \50885 , \48860 , \48515 );
nor \g130377/U$1 ( \50886 , \50884 , \50885 );
not \g130336/U$3 ( \50887 , \50886 );
not \g130336/U$4 ( \50888 , \48685 );
and \g130336/U$2 ( \50889 , \50887 , \50888 );
and \g130336/U$5 ( \50890 , \50886 , \48685 );
nor \g130336/U$1 ( \50891 , \50889 , \50890 );
and \g130982/U$2 ( \50892 , \49888 , \47931 );
and \g130982/U$3 ( \50893 , \47930 , \49714 );
nor \g130982/U$1 ( \50894 , \50892 , \50893 );
not \g130954/U$3 ( \50895 , \50894 );
not \g130954/U$4 ( \50896 , \47935 );
and \g130954/U$2 ( \50897 , \50895 , \50896 );
and \g130954/U$5 ( \50898 , \50894 , \47935 );
nor \g130954/U$1 ( \50899 , \50897 , \50898 );
xor \g130134/U$4 ( \50900 , \50891 , \50899 );
and \g130235/U$2 ( \50901 , \48353 , \49075 );
and \g130235/U$3 ( \50902 , \49074 , \48138 );
nor \g130235/U$1 ( \50903 , \50901 , \50902 );
not \g130195/U$3 ( \50904 , \50903 );
not \g130195/U$4 ( \50905 , \49014 );
and \g130195/U$2 ( \50906 , \50904 , \50905 );
and \g130195/U$5 ( \50907 , \50903 , \49014 );
nor \g130195/U$1 ( \50908 , \50906 , \50907 );
and \g130134/U$3 ( \50909 , \50900 , \50908 );
and \g130134/U$5 ( \50910 , \50891 , \50899 );
or \g130134/U$2 ( \50911 , \50909 , \50910 );
xor \g131122/U$1 ( \50912 , \50753 , \50759 );
xor \g131122/U$1_r1 ( \50913 , \50912 , \50768 );
xor \g129484/U$4 ( \50914 , \50911 , \50913 );
and \g130759/U$2 ( \50915 , \49102 , \48154 );
and \g130759/U$3 ( \50916 , \48155 , \49158 );
nor \g130759/U$1 ( \50917 , \50915 , \50916 );
not \g130732/U$3 ( \50918 , \50917 );
not \g130732/U$4 ( \50919 , \48159 );
and \g130732/U$2 ( \50920 , \50918 , \50919 );
and \g130732/U$5 ( \50921 , \50917 , \48159 );
nor \g130732/U$1 ( \50922 , \50920 , \50921 );
and \g130869/U$2 ( \50923 , \49512 , \48064 );
and \g130869/U$3 ( \50924 , \48063 , \49282 );
nor \g130869/U$1 ( \50925 , \50923 , \50924 );
not \g130843/U$3 ( \50926 , \50925 );
not \g130843/U$4 ( \50927 , \47997 );
and \g130843/U$2 ( \50928 , \50926 , \50927 );
and \g130843/U$5 ( \50929 , \50925 , \47997 );
nor \g130843/U$1 ( \50930 , \50928 , \50929 );
xor \g129598/U$4 ( \50931 , \50922 , \50930 );
and \g129714/U$2 ( \50932 , \47950 , \50160 );
and \g129714/U$3 ( \50933 , \50159 , \47962 );
nor \g129714/U$1 ( \50934 , \50932 , \50933 );
not \g129679/U$3 ( \50935 , \50934 );
not \g129679/U$4 ( \50936 , \49925 );
and \g129679/U$2 ( \50937 , \50935 , \50936 );
and \g129679/U$5 ( \50938 , \50934 , \49925 );
nor \g129679/U$1 ( \50939 , \50937 , \50938 );
and \g129598/U$3 ( \50940 , \50931 , \50939 );
and \g129598/U$5 ( \50941 , \50922 , \50930 );
or \g129598/U$2 ( \50942 , \50940 , \50941 );
and \g129484/U$3 ( \50943 , \50914 , \50942 );
and \g129484/U$5 ( \50944 , \50911 , \50913 );
or \g129484/U$2 ( \50945 , \50943 , \50944 );
and \g131265/U$2 ( \50946 , \50752 , \47960 );
and \g131265/U$3 ( \50947 , \47959 , \50443 );
nor \g131265/U$1 ( \50948 , \50946 , \50947 );
not \g131233/U$3 ( \50949 , \50948 );
not \g131233/U$4 ( \50950 , \47948 );
and \g131233/U$2 ( \50951 , \50949 , \50950 );
and \g131233/U$5 ( \50952 , \50948 , \47948 );
nor \g131233/U$1 ( \50953 , \50951 , \50952 );
and \g131423/U$2 ( \50954 , \44104 , \47620 );
not \g131423/U$4 ( \50955 , \44104 );
and \g131423/U$3 ( \50956 , \50955 , \47621 );
or \g131423/U$1 ( \50957 , \50954 , \50956 );
nand \g131392/U$1 ( \50958 , \40061 , \50957 );
xor \g129773/U$4 ( \50959 , \50953 , \50958 );
and \g129881/U$2 ( \50960 , \48018 , \49813 );
and \g129881/U$3 ( \50961 , \49812 , \47942 );
nor \g129881/U$1 ( \50962 , \50960 , \50961 );
not \g129848/U$3 ( \50963 , \50962 );
not \g129848/U$4 ( \50964 , \49568 );
and \g129848/U$2 ( \50965 , \50963 , \50964 );
and \g129848/U$5 ( \50966 , \50962 , \49568 );
nor \g129848/U$1 ( \50967 , \50965 , \50966 );
and \g129773/U$3 ( \50968 , \50959 , \50967 );
and \g129773/U$5 ( \50969 , \50953 , \50958 );
or \g129773/U$2 ( \50970 , \50968 , \50969 );
and \g130514/U$2 ( \50971 , \48726 , \48479 );
and \g130514/U$3 ( \50972 , \48478 , \48568 );
nor \g130514/U$1 ( \50973 , \50971 , \50972 );
not \g130483/U$3 ( \50974 , \50973 );
not \g130483/U$4 ( \50975 , \48483 );
and \g130483/U$2 ( \50976 , \50974 , \50975 );
and \g130483/U$5 ( \50977 , \50973 , \48483 );
nor \g130483/U$1 ( \50978 , \50976 , \50977 );
and \g130648/U$2 ( \50979 , \48833 , \48334 );
and \g130648/U$3 ( \50980 , \48335 , \48977 );
nor \g130648/U$1 ( \50981 , \50979 , \50980 );
not \g130613/U$3 ( \50982 , \50981 );
not \g130613/U$4 ( \50983 , \48323 );
and \g130613/U$2 ( \50984 , \50982 , \50983 );
and \g130613/U$5 ( \50985 , \50981 , \48323 );
nor \g130613/U$1 ( \50986 , \50984 , \50985 );
xor \g456008/U$5 ( \50987 , \50978 , \50986 );
and \g130069/U$2 ( \50988 , \48051 , \49403 );
and \g130069/U$3 ( \50989 , \49405 , \48117 );
nor \g130069/U$1 ( \50990 , \50988 , \50989 );
not \g130027/U$3 ( \50991 , \50990 );
not \g130027/U$4 ( \50992 , \49233 );
and \g130027/U$2 ( \50993 , \50991 , \50992 );
and \g130027/U$5 ( \50994 , \50990 , \49233 );
nor \g130027/U$1 ( \50995 , \50993 , \50994 );
and \g456008/U$4 ( \50996 , \50987 , \50995 );
and \g456008/U$6 ( \50997 , \50978 , \50986 );
or \g456008/U$3 ( \50998 , \50996 , \50997 );
xor \g129498/U$4 ( \50999 , \50970 , \50998 );
and \g129623/U$2 ( \51000 , \47970 , \50159 );
and \g129623/U$3 ( \51001 , \50160 , \47962 );
nor \g129623/U$1 ( \51002 , \51000 , \51001 );
not \g129578/U$3 ( \51003 , \51002 );
not \g129578/U$4 ( \51004 , \49925 );
and \g129578/U$2 ( \51005 , \51003 , \51004 );
and \g129578/U$5 ( \51006 , \51002 , \49925 );
nor \g129578/U$1 ( \51007 , \51005 , \51006 );
and \g129498/U$3 ( \51008 , \50999 , \51007 );
and \g129498/U$5 ( \51009 , \50970 , \50998 );
or \g129498/U$2 ( \51010 , \51008 , \51009 );
xor \g129056/U$4 ( \51011 , \50945 , \51010 );
xor \g129124/U$1 ( \51012 , \50689 , \50716 );
xor \g129124/U$1_r1 ( \51013 , \51012 , \50745 );
and \g129056/U$3 ( \51014 , \51011 , \51013 );
and \g129056/U$5 ( \51015 , \50945 , \51010 );
or \g129056/U$2 ( \51016 , \51014 , \51015 );
xor \g129385/U$1 ( \51017 , \50640 , \50646 );
xor \g129385/U$1_r1 ( \51018 , \51017 , \50657 );
xor \g128929/U$4 ( \51019 , \51016 , \51018 );
xor \g129016/U$1 ( \51020 , \50748 , \50783 );
xor \g129016/U$1_r1 ( \51021 , \51020 , \50790 );
and \g128929/U$3 ( \51022 , \51019 , \51021 );
and \g128929/U$5 ( \51023 , \51016 , \51018 );
or \g128929/U$2 ( \51024 , \51022 , \51023 );
and \g128861/U$3 ( \51025 , \50883 , \51024 );
and \g128861/U$5 ( \51026 , \50826 , \50882 );
or \g128861/U$2 ( \51027 , \51025 , \51026 );
not \g128860/U$1 ( \51028 , \51027 );
nand \g128849/U$1 ( \51029 , \50820 , \51028 );
nand \g128845/U$1 ( \51030 , \50819 , \51029 );
xor \g130748/U$1 ( \51031 , \50697 , \50704 );
xor \g130748/U$1_r1 ( \51032 , \51031 , \50713 );
xor \g455994/U$9 ( \51033 , \50849 , \50857 );
xor \g455994/U$9_r1 ( \51034 , \51033 , \50866 );
and \g455994/U$8 ( \51035 , \51032 , \51034 );
and \g129515/U$2 ( \51036 , \47970 , \50588 );
and \g129515/U$3 ( \51037 , \50587 , \47972 );
nor \g129515/U$1 ( \51038 , \51036 , \51037 );
not \g129472/U$3 ( \51039 , \51038 );
not \g129472/U$4 ( \51040 , \50362 );
and \g129472/U$2 ( \51041 , \51039 , \51040 );
and \g129472/U$5 ( \51042 , \51038 , \50362 );
nor \g129472/U$1 ( \51043 , \51041 , \51042 );
xor \g129278/U$4 ( \51044 , \51043 , \50856 );
and \g133758/U$2 ( \51045 , \50757 , \50358 );
not \g133758/U$4 ( \51046 , \50757 );
and \g133758/U$3 ( \51047 , \51046 , \50583 );
nor \g133758/U$1 ( \51048 , \51045 , \51047 );
not \g134139/U$1 ( \51049 , \50755 );
and \g133872/U$2 ( \51050 , \50757 , \51049 );
not \g133872/U$4 ( \51051 , \50757 );
and \g133872/U$3 ( \51052 , \51051 , \50755 );
or \g133872/U$1 ( \51053 , \51050 , \51052 );
not \g133851/U$1 ( \51054 , \51053 );
and \g133693/U$1 ( \51055 , \51048 , \51054 );
nand \g129425/U$1 ( \51056 , \51055 , \47894 );
not \g129376/U$3 ( \51057 , \51056 );
not \g129376/U$4 ( \51058 , \50759 );
and \g129376/U$2 ( \51059 , \51057 , \51058 );
and \g129376/U$5 ( \51060 , \51056 , \50759 );
nor \g129376/U$1 ( \51061 , \51059 , \51060 );
and \g129278/U$3 ( \51062 , \51044 , \51061 );
and \g129278/U$5 ( \51063 , \51043 , \50856 );
or \g129278/U$2 ( \51064 , \51062 , \51063 );
xor \g455994/U$11 ( \51065 , \50849 , \50857 );
xor \g455994/U$11_r1 ( \51066 , \51065 , \50866 );
and \g455994/U$10 ( \51067 , \51064 , \51066 );
and \g455994/U$12 ( \51068 , \51032 , \51064 );
or \g455994/U$7 ( \51069 , \51035 , \51067 , \51068 );
xor \g455998/U$2 ( \51070 , \50493 , \50500 );
xor \g455998/U$1 ( \51071 , \51070 , \50509 );
xor \g455998/U$1_r1 ( \51072 , \50828 , \50833 );
xor \g455998/U$1_r2 ( \51073 , \51071 , \51072 );
xor \g129026/U$4 ( \51074 , \51069 , \51073 );
xor \g455988/U$2 ( \51075 , \50442 , \50444 );
xor \g455988/U$1 ( \51076 , \51075 , \50453 );
xor \g455988/U$1_r1 ( \51077 , \50869 , \50874 );
xor \g455988/U$1_r2 ( \51078 , \51076 , \51077 );
and \g129026/U$3 ( \51079 , \51074 , \51078 );
and \g129026/U$5 ( \51080 , \51069 , \51073 );
or \g129026/U$2 ( \51081 , \51079 , \51080 );
xor \g455970/U$9 ( \51082 , \50838 , \50840 );
xor \g455970/U$9_r1 ( \51083 , \51082 , \50879 );
and \g455970/U$8 ( \51084 , \51081 , \51083 );
xor \g129866/U$1 ( \51085 , \50669 , \50677 );
xor \g129866/U$1_r1 ( \51086 , \51085 , \50686 );
xor \g455977/U$9 ( \51087 , \50725 , \50733 );
xor \g455977/U$9_r1 ( \51088 , \51087 , \50742 );
and \g455977/U$8 ( \51089 , \51086 , \51088 );
not \g130550/U$3 ( \51090 , \48483 );
and \g130579/U$2 ( \51091 , \48726 , \48478 );
and \g130579/U$3 ( \51092 , \48479 , \48833 );
nor \g130579/U$1 ( \51093 , \51091 , \51092 );
not \g130550/U$4 ( \51094 , \51093 );
or \g130550/U$2 ( \51095 , \51090 , \51094 );
or \g130550/U$5 ( \51096 , \51093 , \48483 );
nand \g130550/U$1 ( \51097 , \51095 , \51096 );
xor \g131559/U$1 ( \51098 , \44367 , \47615 );
nand \g131528/U$1 ( \51099 , \40061 , \51098 );
not \g131527/U$1 ( \51100 , \51099 );
and \g130388/U$2 ( \51101 , \51097 , \51100 );
not \g130532/U$2 ( \51102 , \51097 );
nand \g130532/U$1 ( \51103 , \51102 , \51099 );
not \g130412/U$3 ( \51104 , \48685 );
and \g130441/U$2 ( \51105 , \48568 , \48860 );
and \g130441/U$3 ( \51106 , \48858 , \48515 );
nor \g130441/U$1 ( \51107 , \51105 , \51106 );
not \g130412/U$4 ( \51108 , \51107 );
or \g130412/U$2 ( \51109 , \51104 , \51108 );
or \g130412/U$5 ( \51110 , \51107 , \48685 );
nand \g130412/U$1 ( \51111 , \51109 , \51110 );
and \g130388/U$3 ( \51112 , \51103 , \51111 );
nor \g130388/U$1 ( \51113 , \51101 , \51112 );
and \g131492/U$2 ( \51114 , \44335 , \47617 );
not \g131492/U$4 ( \51115 , \44335 );
and \g131492/U$3 ( \51116 , \51115 , \47618 );
or \g131492/U$1 ( \51117 , \51114 , \51116 );
nand \g131459/U$1 ( \51118 , \40061 , \51117 );
xor \g135269/U$1 ( \51119 , \24050 , \16062 );
xor \g135269/U$1_r1 ( \51120 , \51119 , \39969 );
xor \g134673/U$1 ( \51121 , \15818 , \23804 );
xor \g134673/U$1_r1 ( \51122 , \51121 , \39972 );
nand \g134149/U$1 ( \51123 , \51120 , \51122 );
and \g134085/U$1 ( \51124 , \50755 , \51123 );
xor \g131121/U$4 ( \51125 , \51118 , \51124 );
and \g131208/U$2 ( \51126 , \50305 , \47913 );
and \g131208/U$3 ( \51127 , \47914 , \50443 );
nor \g131208/U$1 ( \51128 , \51126 , \51127 );
and \g131179/U$2 ( \51129 , \51128 , \47976 );
not \g131179/U$4 ( \51130 , \51128 );
and \g131179/U$3 ( \51131 , \51130 , \47977 );
nor \g131179/U$1 ( \51132 , \51129 , \51131 );
and \g131121/U$3 ( \51133 , \51125 , \51132 );
and \g131121/U$5 ( \51134 , \51118 , \51124 );
or \g131121/U$2 ( \51135 , \51133 , \51134 );
xor \g129121/U$4 ( \51136 , \51113 , \51135 );
and \g129798/U$2 ( \51137 , \47950 , \50159 );
and \g129798/U$3 ( \51138 , \50160 , \47942 );
nor \g129798/U$1 ( \51139 , \51137 , \51138 );
not \g129752/U$3 ( \51140 , \51139 );
not \g129752/U$4 ( \51141 , \49925 );
and \g129752/U$2 ( \51142 , \51140 , \51141 );
and \g129752/U$5 ( \51143 , \51139 , \49925 );
nor \g129752/U$1 ( \51144 , \51142 , \51143 );
and \g131317/U$2 ( \51145 , \50957 , \47960 );
and \g131317/U$3 ( \51146 , \47959 , \50752 );
nor \g131317/U$1 ( \51147 , \51145 , \51146 );
not \g131295/U$3 ( \51148 , \51147 );
not \g131295/U$4 ( \51149 , \47948 );
and \g131295/U$2 ( \51150 , \51148 , \51149 );
and \g131295/U$5 ( \51151 , \51147 , \47948 );
nor \g131295/U$1 ( \51152 , \51150 , \51151 );
xor \g129256/U$4 ( \51153 , \51144 , \51152 );
and \g129398/U$2 ( \51154 , \47894 , \51053 );
and \g129398/U$3 ( \51155 , \51055 , \47972 );
nor \g129398/U$1 ( \51156 , \51154 , \51155 );
not \g129341/U$3 ( \51157 , \51156 );
not \g129341/U$4 ( \51158 , \50759 );
and \g129341/U$2 ( \51159 , \51157 , \51158 );
and \g129341/U$5 ( \51160 , \51156 , \50759 );
nor \g129341/U$1 ( \51161 , \51159 , \51160 );
and \g129256/U$3 ( \51162 , \51153 , \51161 );
and \g129256/U$5 ( \51163 , \51144 , \51152 );
or \g129256/U$2 ( \51164 , \51162 , \51163 );
and \g129121/U$3 ( \51165 , \51136 , \51164 );
and \g129121/U$5 ( \51166 , \51113 , \51135 );
or \g129121/U$2 ( \51167 , \51165 , \51166 );
xor \g455977/U$11 ( \51168 , \50725 , \50733 );
xor \g455977/U$11_r1 ( \51169 , \51168 , \50742 );
and \g455977/U$10 ( \51170 , \51167 , \51169 );
and \g455977/U$12 ( \51171 , \51086 , \51167 );
or \g455977/U$7 ( \51172 , \51089 , \51170 , \51171 );
xor \g130134/U$1 ( \51173 , \50891 , \50899 );
xor \g130134/U$1_r1 ( \51174 , \51173 , \50908 );
xor \g456008/U$9 ( \51175 , \50978 , \50986 );
xor \g456008/U$9_r1 ( \51176 , \51175 , \50995 );
and \g456008/U$8 ( \51177 , \51174 , \51176 );
xor \g129598/U$1 ( \51178 , \50922 , \50930 );
xor \g129598/U$1_r1 ( \51179 , \51178 , \50939 );
xor \g456008/U$11 ( \51180 , \50978 , \50986 );
xor \g456008/U$11_r1 ( \51181 , \51180 , \50995 );
and \g456008/U$10 ( \51182 , \51179 , \51181 );
and \g456008/U$12 ( \51183 , \51174 , \51179 );
or \g456008/U$7 ( \51184 , \51177 , \51182 , \51183 );
not \g130787/U$3 ( \51185 , \48159 );
and \g130815/U$2 ( \51186 , \49282 , \48155 );
and \g130815/U$3 ( \51187 , \48154 , \49158 );
nor \g130815/U$1 ( \51188 , \51186 , \51187 );
not \g130787/U$4 ( \51189 , \51188 );
or \g130787/U$2 ( \51190 , \51185 , \51189 );
or \g130787/U$5 ( \51191 , \51188 , \48159 );
nand \g130787/U$1 ( \51192 , \51190 , \51191 );
not \g130676/U$3 ( \51193 , \48323 );
and \g130702/U$2 ( \51194 , \49102 , \48335 );
and \g130702/U$3 ( \51195 , \48334 , \48977 );
nor \g130702/U$1 ( \51196 , \51194 , \51195 );
not \g130676/U$4 ( \51197 , \51196 );
or \g130676/U$2 ( \51198 , \51193 , \51197 );
or \g130676/U$5 ( \51199 , \51196 , \48323 );
nand \g130676/U$1 ( \51200 , \51198 , \51199 );
xor \g456041/U$4 ( \51201 , \51192 , \51200 );
not \g129932/U$3 ( \51202 , \49568 );
and \g129976/U$2 ( \51203 , \48051 , \49813 );
and \g129976/U$3 ( \51204 , \49812 , \48018 );
nor \g129976/U$1 ( \51205 , \51203 , \51204 );
not \g129932/U$4 ( \51206 , \51205 );
or \g129932/U$2 ( \51207 , \51202 , \51206 );
or \g129932/U$5 ( \51208 , \51205 , \49568 );
nand \g129932/U$1 ( \51209 , \51207 , \51208 );
and \g456041/U$3 ( \51210 , \51201 , \51209 );
and \g456041/U$5 ( \51211 , \51192 , \51200 );
nor \g456041/U$2 ( \51212 , \51210 , \51211 );
not \g131020/U$3 ( \51213 , \47935 );
and \g131061/U$2 ( \51214 , \49888 , \47930 );
and \g131061/U$3 ( \51215 , \47931 , \50019 );
nor \g131061/U$1 ( \51216 , \51214 , \51215 );
not \g131020/U$4 ( \51217 , \51216 );
or \g131020/U$2 ( \51218 , \51213 , \51217 );
or \g131020/U$5 ( \51219 , \51216 , \47935 );
nand \g131020/U$1 ( \51220 , \51218 , \51219 );
not \g130899/U$3 ( \51221 , \47997 );
and \g130926/U$2 ( \51222 , \49512 , \48063 );
and \g130926/U$3 ( \51223 , \48064 , \49714 );
nor \g130926/U$1 ( \51224 , \51222 , \51223 );
not \g130899/U$4 ( \51225 , \51224 );
or \g130899/U$2 ( \51226 , \51221 , \51225 );
or \g130899/U$5 ( \51227 , \51224 , \47997 );
nand \g130899/U$1 ( \51228 , \51226 , \51227 );
xor \g456056/U$4 ( \51229 , \51220 , \51228 );
not \g130271/U$3 ( \51230 , \49014 );
and \g130305/U$2 ( \51231 , \48349 , \49075 );
and \g130305/U$3 ( \51232 , \49074 , \48353 );
nor \g130305/U$1 ( \51233 , \51231 , \51232 );
not \g130271/U$4 ( \51234 , \51233 );
or \g130271/U$2 ( \51235 , \51230 , \51234 );
or \g130271/U$5 ( \51236 , \51233 , \49014 );
nand \g130271/U$1 ( \51237 , \51235 , \51236 );
and \g456056/U$3 ( \51238 , \51229 , \51237 );
and \g456056/U$5 ( \51239 , \51220 , \51228 );
nor \g456056/U$2 ( \51240 , \51238 , \51239 );
xor \g129687/U$4 ( \51241 , \51212 , \51240 );
xor \g129773/U$1 ( \51242 , \50953 , \50958 );
xor \g129773/U$1_r1 ( \51243 , \51242 , \50967 );
and \g129687/U$3 ( \51244 , \51241 , \51243 );
and \g129687/U$5 ( \51245 , \51212 , \51240 );
or \g129687/U$2 ( \51246 , \51244 , \51245 );
xor \g129349/U$4 ( \51247 , \51184 , \51246 );
xor \g129484/U$1 ( \51248 , \50911 , \50913 );
xor \g129484/U$1_r1 ( \51249 , \51248 , \50942 );
and \g129349/U$3 ( \51250 , \51247 , \51249 );
and \g129349/U$5 ( \51251 , \51184 , \51246 );
or \g129349/U$2 ( \51252 , \51250 , \51251 );
xor \g128920/U$4 ( \51253 , \51172 , \51252 );
xor \g129056/U$1 ( \51254 , \50945 , \51010 );
xor \g129056/U$1_r1 ( \51255 , \51254 , \51013 );
and \g128920/U$3 ( \51256 , \51253 , \51255 );
and \g128920/U$5 ( \51257 , \51172 , \51252 );
or \g128920/U$2 ( \51258 , \51256 , \51257 );
xor \g455970/U$11 ( \51259 , \50838 , \50840 );
xor \g455970/U$11_r1 ( \51260 , \51259 , \50879 );
and \g455970/U$10 ( \51261 , \51258 , \51260 );
and \g455970/U$12 ( \51262 , \51081 , \51258 );
or \g455970/U$7 ( \51263 , \51084 , \51261 , \51262 );
not \g128828/U$3 ( \51264 , \51263 );
xor \g128930/U$1 ( \51265 , \50634 , \50660 );
xor \g128930/U$1_r1 ( \51266 , \51265 , \50793 );
not \g128828/U$4 ( \51267 , \51266 );
and \g128828/U$2 ( \51268 , \51264 , \51267 );
and \g128834/U$2 ( \51269 , \51263 , \51266 );
xor \g128861/U$1 ( \51270 , \50826 , \50882 );
xor \g128861/U$1_r1 ( \51271 , \51270 , \51024 );
nor \g128834/U$1 ( \51272 , \51269 , \51271 );
nor \g128828/U$1 ( \51273 , \51268 , \51272 );
xor \g455970/U$2 ( \51274 , \50838 , \50840 );
xor \g455970/U$1 ( \51275 , \51274 , \50879 );
xor \g455970/U$1_r1 ( \51276 , \51081 , \51258 );
xor \g455970/U$1_r2 ( \51277 , \51275 , \51276 );
xor \g128929/U$1 ( \51278 , \51016 , \51018 );
xor \g128929/U$1_r1 ( \51279 , \51278 , \51021 );
or \g128827/U$2 ( \51280 , \51277 , \51279 );
not \g128833/U$3 ( \51281 , \51279 );
not \g128833/U$4 ( \51282 , \51277 );
or \g128833/U$2 ( \51283 , \51281 , \51282 );
xor \g455994/U$2 ( \51284 , \50849 , \50857 );
xor \g455994/U$1 ( \51285 , \51284 , \50866 );
xor \g455994/U$1_r1 ( \51286 , \51032 , \51064 );
xor \g455994/U$1_r2 ( \51287 , \51285 , \51286 );
xor \g129498/U$1 ( \51288 , \50970 , \50998 );
xor \g129498/U$1_r1 ( \51289 , \51288 , \51007 );
xor \g455973/U$5 ( \51290 , \51287 , \51289 );
and \g131264/U$2 ( \51291 , \50752 , \47914 );
and \g131264/U$3 ( \51292 , \47913 , \50443 );
nor \g131264/U$1 ( \51293 , \51291 , \51292 );
and \g131232/U$2 ( \51294 , \51293 , \47977 );
not \g131232/U$4 ( \51295 , \51293 );
and \g131232/U$3 ( \51296 , \51295 , \47976 );
nor \g131232/U$1 ( \51297 , \51294 , \51296 );
not \g131353/U$3 ( \51298 , \47948 );
and \g131373/U$2 ( \51299 , \51117 , \47960 );
and \g131373/U$3 ( \51300 , \47959 , \50957 );
nor \g131373/U$1 ( \51301 , \51299 , \51300 );
not \g131353/U$4 ( \51302 , \51301 );
or \g131353/U$2 ( \51303 , \51298 , \51302 );
or \g131353/U$5 ( \51304 , \51301 , \47948 );
nand \g131353/U$1 ( \51305 , \51303 , \51304 );
xor \g131040/U$4 ( \51306 , \51297 , \51305 );
not \g131100/U$3 ( \51307 , \47935 );
and \g131136/U$2 ( \51308 , \50305 , \47931 );
and \g131136/U$3 ( \51309 , \47930 , \50019 );
nor \g131136/U$1 ( \51310 , \51308 , \51309 );
not \g131100/U$4 ( \51311 , \51310 );
or \g131100/U$2 ( \51312 , \51307 , \51311 );
or \g131100/U$5 ( \51313 , \51310 , \47935 );
nand \g131100/U$1 ( \51314 , \51312 , \51313 );
and \g131040/U$3 ( \51315 , \51306 , \51314 );
and \g131040/U$5 ( \51316 , \51297 , \51305 );
or \g131040/U$2 ( \51317 , \51315 , \51316 );
not \g130117/U$3 ( \51318 , \49233 );
and \g130155/U$2 ( \51319 , \48117 , \49403 );
and \g130155/U$3 ( \51320 , \49405 , \48138 );
nor \g130155/U$1 ( \51321 , \51319 , \51320 );
not \g130117/U$4 ( \51322 , \51321 );
or \g130117/U$2 ( \51323 , \51318 , \51322 );
or \g130117/U$5 ( \51324 , \51321 , \49233 );
nand \g130117/U$1 ( \51325 , \51323 , \51324 );
xor \g456012/U$4 ( \51326 , \51317 , \51325 );
not \g129577/U$3 ( \51327 , \50362 );
and \g129622/U$2 ( \51328 , \47970 , \50587 );
and \g129622/U$3 ( \51329 , \50588 , \47962 );
nor \g129622/U$1 ( \51330 , \51328 , \51329 );
not \g129577/U$4 ( \51331 , \51330 );
or \g129577/U$2 ( \51332 , \51327 , \51331 );
or \g129577/U$5 ( \51333 , \51330 , \50362 );
nand \g129577/U$1 ( \51334 , \51332 , \51333 );
and \g456012/U$3 ( \51335 , \51326 , \51334 );
and \g456012/U$5 ( \51336 , \51317 , \51325 );
nor \g456012/U$2 ( \51337 , \51335 , \51336 );
not \g130731/U$3 ( \51338 , \48323 );
and \g130758/U$2 ( \51339 , \49102 , \48334 );
and \g130758/U$3 ( \51340 , \48335 , \49158 );
nor \g130758/U$1 ( \51341 , \51339 , \51340 );
not \g130731/U$4 ( \51342 , \51341 );
or \g130731/U$2 ( \51343 , \51338 , \51342 );
or \g130731/U$5 ( \51344 , \51341 , \48323 );
nand \g130731/U$1 ( \51345 , \51343 , \51344 );
not \g130612/U$3 ( \51346 , \48483 );
and \g130647/U$2 ( \51347 , \48833 , \48478 );
and \g130647/U$3 ( \51348 , \48479 , \48977 );
nor \g130647/U$1 ( \51349 , \51347 , \51348 );
not \g130612/U$4 ( \51350 , \51349 );
or \g130612/U$2 ( \51351 , \51346 , \51350 );
or \g130612/U$5 ( \51352 , \51349 , \48483 );
nand \g130612/U$1 ( \51353 , \51351 , \51352 );
xor \g456045/U$4 ( \51354 , \51345 , \51353 );
not \g130026/U$3 ( \51355 , \49568 );
and \g130068/U$2 ( \51356 , \48051 , \49812 );
and \g130068/U$3 ( \51357 , \49813 , \48117 );
nor \g130068/U$1 ( \51358 , \51356 , \51357 );
not \g130026/U$4 ( \51359 , \51358 );
or \g130026/U$2 ( \51360 , \51355 , \51359 );
or \g130026/U$5 ( \51361 , \51358 , \49568 );
nand \g130026/U$1 ( \51362 , \51360 , \51361 );
and \g456045/U$3 ( \51363 , \51354 , \51362 );
and \g456045/U$5 ( \51364 , \51345 , \51353 );
nor \g456045/U$2 ( \51365 , \51363 , \51364 );
not \g129736/U$3 ( \51366 , \51365 );
xor \g131121/U$1 ( \51367 , \51118 , \51124 );
xor \g131121/U$1_r1 ( \51368 , \51367 , \51132 );
not \g129736/U$4 ( \51369 , \51368 );
and \g129736/U$2 ( \51370 , \51366 , \51369 );
and \g129740/U$2 ( \51371 , \51365 , \51368 );
not \g130482/U$3 ( \51372 , \48685 );
and \g130513/U$2 ( \51373 , \48726 , \48860 );
and \g130513/U$3 ( \51374 , \48858 , \48568 );
nor \g130513/U$1 ( \51375 , \51373 , \51374 );
not \g130482/U$4 ( \51376 , \51375 );
or \g130482/U$2 ( \51377 , \51372 , \51376 );
or \g130482/U$5 ( \51378 , \51375 , \48685 );
nand \g130482/U$1 ( \51379 , \51377 , \51378 );
xor \g129772/U$4 ( \51380 , \51379 , \51099 );
not \g129847/U$3 ( \51381 , \49925 );
and \g129880/U$2 ( \51382 , \48018 , \50160 );
and \g129880/U$3 ( \51383 , \50159 , \47942 );
nor \g129880/U$1 ( \51384 , \51382 , \51383 );
not \g129847/U$4 ( \51385 , \51384 );
or \g129847/U$2 ( \51386 , \51381 , \51385 );
or \g129847/U$5 ( \51387 , \51384 , \49925 );
nand \g129847/U$1 ( \51388 , \51386 , \51387 );
and \g129772/U$3 ( \51389 , \51380 , \51388 );
and \g129772/U$5 ( \51390 , \51379 , \51099 );
or \g129772/U$2 ( \51391 , \51389 , \51390 );
not \g129771/U$1 ( \51392 , \51391 );
nor \g129740/U$1 ( \51393 , \51371 , \51392 );
nor \g129736/U$1 ( \51394 , \51370 , \51393 );
xor \g129130/U$4 ( \51395 , \51337 , \51394 );
xor \g129278/U$1 ( \51396 , \51043 , \50856 );
xor \g129278/U$1_r1 ( \51397 , \51396 , \51061 );
and \g129130/U$3 ( \51398 , \51395 , \51397 );
and \g129130/U$5 ( \51399 , \51337 , \51394 );
or \g129130/U$2 ( \51400 , \51398 , \51399 );
and \g455973/U$4 ( \51401 , \51290 , \51400 );
and \g455973/U$6 ( \51402 , \51287 , \51289 );
or \g455973/U$3 ( \51403 , \51401 , \51402 );
xor \g455977/U$2 ( \51404 , \50725 , \50733 );
xor \g455977/U$1 ( \51405 , \51404 , \50742 );
xor \g455977/U$1_r1 ( \51406 , \51086 , \51167 );
xor \g455977/U$1_r2 ( \51407 , \51405 , \51406 );
not \g128954/U$3 ( \51408 , \51407 );
xor \g129349/U$1 ( \51409 , \51184 , \51246 );
xor \g129349/U$1_r1 ( \51410 , \51409 , \51249 );
not \g128954/U$4 ( \51411 , \51410 );
and \g128954/U$2 ( \51412 , \51408 , \51411 );
and \g128963/U$2 ( \51413 , \51407 , \51410 );
xor \g456041/U$1 ( \51414 , \51192 , \51200 );
xor \g456041/U$1_r1 ( \51415 , \51414 , \51209 );
and \g130506/U$2 ( \51416 , \51097 , \51099 );
not \g130506/U$4 ( \51417 , \51097 );
and \g130506/U$3 ( \51418 , \51417 , \51100 );
nor \g130506/U$1 ( \51419 , \51416 , \51418 );
not \g130391/U$3 ( \51420 , \51419 );
not \g130391/U$4 ( \51421 , \51111 );
or \g130391/U$2 ( \51422 , \51420 , \51421 );
or \g130391/U$5 ( \51423 , \51111 , \51419 );
nand \g130391/U$1 ( \51424 , \51422 , \51423 );
and \g129196/U$2 ( \51425 , \51415 , \51424 );
not \g129209/U$3 ( \51426 , \51415 );
not \g129209/U$4 ( \51427 , \51424 );
and \g129209/U$2 ( \51428 , \51426 , \51427 );
xor \g129256/U$1 ( \51429 , \51144 , \51152 );
xor \g129256/U$1_r1 ( \51430 , \51429 , \51161 );
nor \g129209/U$1 ( \51431 , \51428 , \51430 );
nor \g129196/U$1 ( \51432 , \51425 , \51431 );
xor \g129687/U$1 ( \51433 , \51212 , \51240 );
xor \g129687/U$1_r1 ( \51434 , \51433 , \51243 );
xor \g129011/U$4 ( \51435 , \51432 , \51434 );
xor \g129121/U$1 ( \51436 , \51113 , \51135 );
xor \g129121/U$1_r1 ( \51437 , \51436 , \51164 );
and \g129011/U$3 ( \51438 , \51435 , \51437 );
and \g129011/U$5 ( \51439 , \51432 , \51434 );
or \g129011/U$2 ( \51440 , \51438 , \51439 );
nor \g128963/U$1 ( \51441 , \51413 , \51440 );
nor \g128954/U$1 ( \51442 , \51412 , \51441 );
xor \g455972/U$4 ( \51443 , \51403 , \51442 );
xor \g129026/U$1 ( \51444 , \51069 , \51073 );
xor \g129026/U$1_r1 ( \51445 , \51444 , \51078 );
and \g455972/U$3 ( \51446 , \51443 , \51445 );
and \g455972/U$5 ( \51447 , \51403 , \51442 );
nor \g455972/U$2 ( \51448 , \51446 , \51447 );
nand \g128833/U$1 ( \51449 , \51283 , \51448 );
nand \g128827/U$1 ( \51450 , \51280 , \51449 );
xor \g128920/U$1 ( \51451 , \51172 , \51252 );
xor \g128920/U$1_r1 ( \51452 , \51451 , \51255 );
not \g128823/U$3 ( \51453 , \51452 );
not \g130845/U$3 ( \51454 , \48159 );
and \g130871/U$2 ( \51455 , \49512 , \48155 );
and \g130871/U$3 ( \51456 , \48154 , \49282 );
nor \g130871/U$1 ( \51457 , \51455 , \51456 );
not \g130845/U$4 ( \51458 , \51457 );
or \g130845/U$2 ( \51459 , \51454 , \51458 );
or \g130845/U$5 ( \51460 , \51457 , \48159 );
nand \g130845/U$1 ( \51461 , \51459 , \51460 );
not \g130956/U$3 ( \51462 , \47997 );
and \g130984/U$2 ( \51463 , \49888 , \48064 );
and \g130984/U$3 ( \51464 , \48063 , \49714 );
nor \g130984/U$1 ( \51465 , \51463 , \51464 );
not \g130956/U$4 ( \51466 , \51465 );
or \g130956/U$2 ( \51467 , \51462 , \51466 );
or \g130956/U$5 ( \51468 , \51465 , \47997 );
nand \g130956/U$1 ( \51469 , \51467 , \51468 );
xor \g129600/U$4 ( \51470 , \51461 , \51469 );
not \g129681/U$3 ( \51471 , \50362 );
and \g129716/U$2 ( \51472 , \47950 , \50588 );
and \g129716/U$3 ( \51473 , \50587 , \47962 );
nor \g129716/U$1 ( \51474 , \51472 , \51473 );
not \g129681/U$4 ( \51475 , \51474 );
or \g129681/U$2 ( \51476 , \51471 , \51475 );
or \g129681/U$5 ( \51477 , \51474 , \50362 );
nand \g129681/U$1 ( \51478 , \51476 , \51477 );
and \g129600/U$3 ( \51479 , \51470 , \51478 );
and \g129600/U$5 ( \51480 , \51461 , \51469 );
or \g129600/U$2 ( \51481 , \51479 , \51480 );
xor \g456056/U$1 ( \51482 , \51220 , \51228 );
xor \g456056/U$1_r1 ( \51483 , \51482 , \51237 );
and \g129229/U$2 ( \51484 , \51481 , \51483 );
not \g129241/U$3 ( \51485 , \51481 );
not \g129241/U$4 ( \51486 , \51483 );
and \g129241/U$2 ( \51487 , \51485 , \51486 );
not \g130198/U$3 ( \51488 , \49233 );
and \g130237/U$2 ( \51489 , \48353 , \49405 );
and \g130237/U$3 ( \51490 , \49403 , \48138 );
nor \g130237/U$1 ( \51491 , \51489 , \51490 );
not \g130198/U$4 ( \51492 , \51491 );
or \g130198/U$2 ( \51493 , \51488 , \51492 );
or \g130198/U$5 ( \51494 , \51491 , \49233 );
nand \g130198/U$1 ( \51495 , \51493 , \51494 );
not \g130338/U$3 ( \51496 , \49014 );
and \g130379/U$2 ( \51497 , \48349 , \49074 );
and \g130379/U$3 ( \51498 , \49075 , \48515 );
nor \g130379/U$1 ( \51499 , \51497 , \51498 );
not \g130338/U$4 ( \51500 , \51499 );
or \g130338/U$2 ( \51501 , \51496 , \51500 );
or \g130338/U$5 ( \51502 , \51499 , \49014 );
nand \g130338/U$1 ( \51503 , \51501 , \51502 );
and \g129320/U$2 ( \51504 , \51495 , \51503 );
not \g129327/U$3 ( \51505 , \51495 );
not \g129327/U$4 ( \51506 , \51503 );
and \g129327/U$2 ( \51507 , \51505 , \51506 );
and \g134068/U$2 ( \51508 , \51122 , \50755 );
not \g134068/U$4 ( \51509 , \51122 );
and \g134068/U$3 ( \51510 , \51509 , \51049 );
nor \g134068/U$1 ( \51511 , \51508 , \51510 );
not \g135564/U$2 ( \51512 , \51511 );
not \g135268/U$1 ( \51513 , \51120 );
and \g134148/U$2 ( \51514 , \51122 , \51513 );
not \g134148/U$4 ( \51515 , \51122 );
and \g134148/U$3 ( \51516 , \51515 , \51120 );
or \g134148/U$1 ( \51517 , \51514 , \51516 );
nor \g135564/U$1 ( \51518 , \51512 , \51517 );
nand \g129429/U$1 ( \51519 , \51518 , \47894 );
not \g129378/U$3 ( \51520 , \51519 );
not \g129378/U$4 ( \51521 , \51124 );
and \g129378/U$2 ( \51522 , \51520 , \51521 );
and \g129378/U$5 ( \51523 , \51519 , \51124 );
nor \g129378/U$1 ( \51524 , \51522 , \51523 );
nor \g129327/U$1 ( \51525 , \51507 , \51524 );
nor \g129320/U$1 ( \51526 , \51504 , \51525 );
nor \g129241/U$1 ( \51527 , \51487 , \51526 );
nor \g129229/U$1 ( \51528 , \51484 , \51527 );
not \g129003/U$3 ( \51529 , \51528 );
xor \g456008/U$2 ( \51530 , \50978 , \50986 );
xor \g456008/U$1 ( \51531 , \51530 , \50995 );
xor \g456008/U$1_r1 ( \51532 , \51174 , \51179 );
xor \g456008/U$1_r2 ( \51533 , \51531 , \51532 );
not \g129003/U$4 ( \51534 , \51533 );
and \g129003/U$2 ( \51535 , \51529 , \51534 );
and \g129020/U$2 ( \51536 , \51528 , \51533 );
and \g131318/U$2 ( \51537 , \50957 , \47914 );
and \g131318/U$3 ( \51538 , \47913 , \50752 );
nor \g131318/U$1 ( \51539 , \51537 , \51538 );
and \g131293/U$2 ( \51540 , \51539 , \47977 );
not \g131293/U$4 ( \51541 , \51539 );
and \g131293/U$3 ( \51542 , \51541 , \47976 );
nor \g131293/U$1 ( \51543 , \51540 , \51542 );
not \g131409/U$3 ( \51544 , \47948 );
and \g131442/U$2 ( \51545 , \51117 , \47959 );
and \g131442/U$3 ( \51546 , \47960 , \51098 );
nor \g131442/U$1 ( \51547 , \51545 , \51546 );
not \g131409/U$4 ( \51548 , \51547 );
or \g131409/U$2 ( \51549 , \51544 , \51548 );
or \g131409/U$5 ( \51550 , \51547 , \47948 );
nand \g131409/U$1 ( \51551 , \51549 , \51550 );
xor \g131123/U$4 ( \51552 , \51543 , \51551 );
not \g131181/U$3 ( \51553 , \47935 );
and \g131210/U$2 ( \51554 , \50305 , \47930 );
and \g131210/U$3 ( \51555 , \47931 , \50443 );
nor \g131210/U$1 ( \51556 , \51554 , \51555 );
not \g131181/U$4 ( \51557 , \51556 );
or \g131181/U$2 ( \51558 , \51553 , \51557 );
or \g131181/U$5 ( \51559 , \51556 , \47935 );
nand \g131181/U$1 ( \51560 , \51558 , \51559 );
and \g131123/U$3 ( \51561 , \51552 , \51560 );
and \g131123/U$5 ( \51562 , \51543 , \51551 );
or \g131123/U$2 ( \51563 , \51561 , \51562 );
xor \g131613/U$1 ( \51564 , \47613 , \47612 );
not \g135522/U$2 ( \51565 , \51564 );
nor \g135522/U$1 ( \51566 , \51565 , \40060 );
nor \g131566/U$1 ( \51567 , \51566 , \51513 );
not \g131565/U$1 ( \51568 , \51567 );
xor \g129407/U$4 ( \51569 , \51563 , \51568 );
not \g129474/U$3 ( \51570 , \50759 );
and \g129517/U$2 ( \51571 , \47970 , \51055 );
and \g129517/U$3 ( \51572 , \51053 , \47972 );
nor \g129517/U$1 ( \51573 , \51571 , \51572 );
not \g129474/U$4 ( \51574 , \51573 );
or \g129474/U$2 ( \51575 , \51570 , \51574 );
or \g129474/U$5 ( \51576 , \51573 , \50759 );
nand \g129474/U$1 ( \51577 , \51575 , \51576 );
and \g129407/U$3 ( \51578 , \51569 , \51577 );
and \g129407/U$5 ( \51579 , \51563 , \51568 );
or \g129407/U$2 ( \51580 , \51578 , \51579 );
xor \g456012/U$1 ( \51581 , \51317 , \51325 );
xor \g456012/U$1_r1 ( \51582 , \51581 , \51334 );
xor \g129054/U$4 ( \51583 , \51580 , \51582 );
not \g130552/U$3 ( \51584 , \48685 );
and \g130581/U$2 ( \51585 , \48726 , \48858 );
and \g130581/U$3 ( \51586 , \48860 , \48833 );
nor \g130581/U$1 ( \51587 , \51585 , \51586 );
not \g130552/U$4 ( \51588 , \51587 );
or \g130552/U$2 ( \51589 , \51584 , \51588 );
or \g130552/U$5 ( \51590 , \51587 , \48685 );
nand \g130552/U$1 ( \51591 , \51589 , \51590 );
not \g131480/U$3 ( \51592 , \47948 );
and \g131508/U$2 ( \51593 , \51564 , \47960 );
and \g131508/U$3 ( \51594 , \47959 , \51098 );
nor \g131508/U$1 ( \51595 , \51593 , \51594 );
not \g131480/U$4 ( \51596 , \51595 );
or \g131480/U$2 ( \51597 , \51592 , \51596 );
or \g131480/U$5 ( \51598 , \51595 , \47948 );
nand \g131480/U$1 ( \51599 , \51597 , \51598 );
not \g131460/U$2 ( \51600 , \51599 );
and \g131671/U$2 ( \51601 , \47609 , \47597 );
not \g131671/U$4 ( \51602 , \47609 );
and \g131671/U$3 ( \51603 , \51602 , \47598 );
or \g131671/U$1 ( \51604 , \51601 , \51603 );
nand \g131646/U$1 ( \51605 , \40061 , \51604 );
nor \g131460/U$1 ( \51606 , \51600 , \51605 );
xor \g129865/U$4 ( \51607 , \51591 , \51606 );
not \g129934/U$3 ( \51608 , \49925 );
and \g129978/U$2 ( \51609 , \48051 , \50160 );
and \g129978/U$3 ( \51610 , \50159 , \48018 );
nor \g129978/U$1 ( \51611 , \51609 , \51610 );
not \g129934/U$4 ( \51612 , \51611 );
or \g129934/U$2 ( \51613 , \51608 , \51612 );
or \g129934/U$5 ( \51614 , \51611 , \49925 );
nand \g129934/U$1 ( \51615 , \51613 , \51614 );
and \g129865/U$3 ( \51616 , \51607 , \51615 );
and \g129865/U$5 ( \51617 , \51591 , \51606 );
or \g129865/U$2 ( \51618 , \51616 , \51617 );
xor \g131040/U$1 ( \51619 , \51297 , \51305 );
xor \g131040/U$1_r1 ( \51620 , \51619 , \51314 );
xor \g129155/U$4 ( \51621 , \51618 , \51620 );
not \g129754/U$3 ( \51622 , \50362 );
and \g129800/U$2 ( \51623 , \47950 , \50587 );
and \g129800/U$3 ( \51624 , \50588 , \47942 );
nor \g129800/U$1 ( \51625 , \51623 , \51624 );
not \g129754/U$4 ( \51626 , \51625 );
or \g129754/U$2 ( \51627 , \51622 , \51626 );
or \g129754/U$5 ( \51628 , \51625 , \50362 );
nand \g129754/U$1 ( \51629 , \51627 , \51628 );
not \g130414/U$3 ( \51630 , \49014 );
and \g130443/U$2 ( \51631 , \48568 , \49075 );
and \g130443/U$3 ( \51632 , \49074 , \48515 );
nor \g130443/U$1 ( \51633 , \51631 , \51632 );
not \g130414/U$4 ( \51634 , \51633 );
or \g130414/U$2 ( \51635 , \51630 , \51634 );
or \g130414/U$5 ( \51636 , \51633 , \49014 );
nand \g130414/U$1 ( \51637 , \51635 , \51636 );
xor \g129258/U$4 ( \51638 , \51629 , \51637 );
not \g129343/U$3 ( \51639 , \51124 );
and \g129402/U$2 ( \51640 , \47894 , \51517 );
and \g129402/U$3 ( \51641 , \51518 , \47972 );
nor \g129402/U$1 ( \51642 , \51640 , \51641 );
not \g129343/U$4 ( \51643 , \51642 );
or \g129343/U$2 ( \51644 , \51639 , \51643 );
or \g129343/U$5 ( \51645 , \51642 , \51124 );
nand \g129343/U$1 ( \51646 , \51644 , \51645 );
and \g129258/U$3 ( \51647 , \51638 , \51646 );
and \g129258/U$5 ( \51648 , \51629 , \51637 );
or \g129258/U$2 ( \51649 , \51647 , \51648 );
and \g129155/U$3 ( \51650 , \51621 , \51649 );
and \g129155/U$5 ( \51651 , \51618 , \51620 );
or \g129155/U$2 ( \51652 , \51650 , \51651 );
and \g129054/U$3 ( \51653 , \51583 , \51652 );
and \g129054/U$5 ( \51654 , \51580 , \51582 );
or \g129054/U$2 ( \51655 , \51653 , \51654 );
not \g129053/U$1 ( \51656 , \51655 );
nor \g129020/U$1 ( \51657 , \51536 , \51656 );
nor \g129003/U$1 ( \51658 , \51535 , \51657 );
xor \g455973/U$9 ( \51659 , \51287 , \51289 );
xor \g455973/U$9_r1 ( \51660 , \51659 , \51400 );
and \g455973/U$8 ( \51661 , \51658 , \51660 );
not \g129214/U$3 ( \51662 , \51483 );
not \g129214/U$4 ( \51663 , \51526 );
or \g129214/U$2 ( \51664 , \51662 , \51663 );
or \g129214/U$5 ( \51665 , \51526 , \51483 );
nand \g129214/U$1 ( \51666 , \51664 , \51665 );
xor \g455935/U$1 ( \51667 , \51481 , \51666 );
xor \g129772/U$1 ( \51668 , \51379 , \51099 );
xor \g129772/U$1_r1 ( \51669 , \51668 , \51388 );
xor \g456045/U$1 ( \51670 , \51345 , \51353 );
xor \g456045/U$1_r1 ( \51671 , \51670 , \51362 );
xor \g455990/U$5 ( \51672 , \51669 , \51671 );
xor \g129600/U$1 ( \51673 , \51461 , \51469 );
xor \g129600/U$1_r1 ( \51674 , \51673 , \51478 );
and \g455990/U$4 ( \51675 , \51672 , \51674 );
and \g455990/U$6 ( \51676 , \51669 , \51671 );
or \g455990/U$3 ( \51677 , \51675 , \51676 );
xor \g455980/U$4 ( \51678 , \51667 , \51677 );
not \g130272/U$3 ( \51679 , \49233 );
and \g130306/U$2 ( \51680 , \48349 , \49405 );
and \g130306/U$3 ( \51681 , \49403 , \48353 );
nor \g130306/U$1 ( \51682 , \51680 , \51681 );
not \g130272/U$4 ( \51683 , \51682 );
or \g130272/U$2 ( \51684 , \51679 , \51683 );
or \g130272/U$5 ( \51685 , \51682 , \49233 );
nand \g130272/U$1 ( \51686 , \51684 , \51685 );
not \g131021/U$3 ( \51687 , \47997 );
and \g131062/U$2 ( \51688 , \49888 , \48063 );
and \g131062/U$3 ( \51689 , \48064 , \50019 );
nor \g131062/U$1 ( \51690 , \51688 , \51689 );
not \g131021/U$4 ( \51691 , \51690 );
or \g131021/U$2 ( \51692 , \51687 , \51691 );
or \g131021/U$5 ( \51693 , \51690 , \47997 );
nand \g131021/U$1 ( \51694 , \51692 , \51693 );
xor \g456009/U$5 ( \51695 , \51686 , \51694 );
not \g130119/U$3 ( \51696 , \49568 );
and \g130157/U$2 ( \51697 , \48117 , \49812 );
and \g130157/U$3 ( \51698 , \49813 , \48138 );
nor \g130157/U$1 ( \51699 , \51697 , \51698 );
not \g130119/U$4 ( \51700 , \51699 );
or \g130119/U$2 ( \51701 , \51696 , \51700 );
or \g130119/U$5 ( \51702 , \51699 , \49568 );
nand \g130119/U$1 ( \51703 , \51701 , \51702 );
and \g456009/U$4 ( \51704 , \51695 , \51703 );
and \g456009/U$6 ( \51705 , \51686 , \51694 );
or \g456009/U$3 ( \51706 , \51704 , \51705 );
not \g130793/U$3 ( \51707 , \48323 );
and \g130813/U$2 ( \51708 , \49282 , \48335 );
and \g130813/U$3 ( \51709 , \48334 , \49158 );
nor \g130813/U$1 ( \51710 , \51708 , \51709 );
not \g130793/U$4 ( \51711 , \51710 );
or \g130793/U$2 ( \51712 , \51707 , \51711 );
or \g130793/U$5 ( \51713 , \51710 , \48323 );
nand \g130793/U$1 ( \51714 , \51712 , \51713 );
not \g130900/U$3 ( \51715 , \48159 );
and \g130927/U$2 ( \51716 , \49512 , \48154 );
and \g130927/U$3 ( \51717 , \48155 , \49714 );
nor \g130927/U$1 ( \51718 , \51716 , \51717 );
not \g130900/U$4 ( \51719 , \51718 );
or \g130900/U$2 ( \51720 , \51715 , \51719 );
or \g130900/U$5 ( \51721 , \51718 , \48159 );
nand \g130900/U$1 ( \51722 , \51720 , \51721 );
xor \g130630/U$4 ( \51723 , \51714 , \51722 );
not \g130678/U$3 ( \51724 , \48483 );
and \g130704/U$2 ( \51725 , \49102 , \48479 );
and \g130704/U$3 ( \51726 , \48478 , \48977 );
nor \g130704/U$1 ( \51727 , \51725 , \51726 );
not \g130678/U$4 ( \51728 , \51727 );
or \g130678/U$2 ( \51729 , \51724 , \51728 );
or \g130678/U$5 ( \51730 , \51727 , \48483 );
nand \g130678/U$1 ( \51731 , \51729 , \51730 );
and \g130630/U$3 ( \51732 , \51723 , \51731 );
and \g130630/U$5 ( \51733 , \51714 , \51722 );
or \g130630/U$2 ( \51734 , \51732 , \51733 );
xor \g129131/U$4 ( \51735 , \51706 , \51734 );
not \g129312/U$3 ( \51736 , \51503 );
not \g129312/U$4 ( \51737 , \51524 );
or \g129312/U$2 ( \51738 , \51736 , \51737 );
or \g129312/U$5 ( \51739 , \51524 , \51503 );
nand \g129312/U$1 ( \51740 , \51738 , \51739 );
xor \g455940/U$1 ( \51741 , \51495 , \51740 );
and \g129131/U$3 ( \51742 , \51735 , \51741 );
and \g129131/U$5 ( \51743 , \51706 , \51734 );
or \g129131/U$2 ( \51744 , \51742 , \51743 );
and \g455980/U$3 ( \51745 , \51678 , \51744 );
and \g455980/U$5 ( \51746 , \51667 , \51677 );
nor \g455980/U$2 ( \51747 , \51745 , \51746 );
not \g128951/U$3 ( \51748 , \51747 );
xor \g129130/U$1 ( \51749 , \51337 , \51394 );
xor \g129130/U$1_r1 ( \51750 , \51749 , \51397 );
not \g128951/U$4 ( \51751 , \51750 );
and \g128951/U$2 ( \51752 , \51748 , \51751 );
and \g128960/U$2 ( \51753 , \51747 , \51750 );
xor \g129011/U$1 ( \51754 , \51432 , \51434 );
xor \g129011/U$1_r1 ( \51755 , \51754 , \51437 );
nor \g128960/U$1 ( \51756 , \51753 , \51755 );
nor \g128951/U$1 ( \51757 , \51752 , \51756 );
xor \g455973/U$11 ( \51758 , \51287 , \51289 );
xor \g455973/U$11_r1 ( \51759 , \51758 , \51400 );
and \g455973/U$10 ( \51760 , \51757 , \51759 );
and \g455973/U$12 ( \51761 , \51658 , \51757 );
or \g455973/U$7 ( \51762 , \51661 , \51760 , \51761 );
xor \g455972/U$1 ( \51763 , \51403 , \51442 );
xor \g455972/U$1_r1 ( \51764 , \51763 , \51445 );
xor \g128836/U$1 ( \51765 , \51762 , \51764 );
not \g128823/U$4 ( \51766 , \51765 );
or \g128823/U$2 ( \51767 , \51453 , \51766 );
or \g128823/U$5 ( \51768 , \51765 , \51452 );
nand \g128823/U$1 ( \51769 , \51767 , \51768 );
xor \g455973/U$2 ( \51770 , \51287 , \51289 );
xor \g455973/U$1 ( \51771 , \51770 , \51400 );
xor \g455973/U$1_r1 ( \51772 , \51658 , \51757 );
xor \g455973/U$1_r2 ( \51773 , \51771 , \51772 );
not \g128943/U$3 ( \51774 , \51407 );
xor \g128971/U$1 ( \51775 , \51410 , \51440 );
not \g128943/U$4 ( \51776 , \51775 );
or \g128943/U$2 ( \51777 , \51774 , \51776 );
or \g128943/U$5 ( \51778 , \51775 , \51407 );
nand \g128943/U$1 ( \51779 , \51777 , \51778 );
not \g128927/U$1 ( \51780 , \51779 );
or \g128844/U$2 ( \51781 , \51773 , \51780 );
not \g128848/U$3 ( \51782 , \51780 );
not \g128848/U$4 ( \51783 , \51773 );
or \g128848/U$2 ( \51784 , \51782 , \51783 );
not \g128980/U$3 ( \51785 , \51528 );
not \g129001/U$3 ( \51786 , \51533 );
not \g129001/U$4 ( \51787 , \51655 );
or \g129001/U$2 ( \51788 , \51786 , \51787 );
or \g129001/U$5 ( \51789 , \51655 , \51533 );
nand \g129001/U$1 ( \51790 , \51788 , \51789 );
not \g128980/U$4 ( \51791 , \51790 );
or \g128980/U$2 ( \51792 , \51785 , \51791 );
or \g128980/U$5 ( \51793 , \51790 , \51528 );
nand \g128980/U$1 ( \51794 , \51792 , \51793 );
and \g131266/U$2 ( \51795 , \50752 , \47931 );
and \g131266/U$3 ( \51796 , \47930 , \50443 );
nor \g131266/U$1 ( \51797 , \51795 , \51796 );
not \g131234/U$3 ( \51798 , \51797 );
not \g131234/U$4 ( \51799 , \47935 );
and \g131234/U$2 ( \51800 , \51798 , \51799 );
and \g131234/U$5 ( \51801 , \51797 , \47935 );
nor \g131234/U$1 ( \51802 , \51800 , \51801 );
and \g131375/U$2 ( \51803 , \51117 , \47914 );
and \g131375/U$3 ( \51804 , \47913 , \50957 );
nor \g131375/U$1 ( \51805 , \51803 , \51804 );
and \g131354/U$2 ( \51806 , \51805 , \47976 );
not \g131354/U$4 ( \51807 , \51805 );
and \g131354/U$3 ( \51808 , \51807 , \47977 );
nor \g131354/U$1 ( \51809 , \51806 , \51808 );
xor \g131042/U$4 ( \51810 , \51802 , \51809 );
and \g131139/U$2 ( \51811 , \50305 , \48064 );
and \g131139/U$3 ( \51812 , \48063 , \50019 );
nor \g131139/U$1 ( \51813 , \51811 , \51812 );
not \g131105/U$3 ( \51814 , \51813 );
not \g131105/U$4 ( \51815 , \47997 );
and \g131105/U$2 ( \51816 , \51814 , \51815 );
and \g131105/U$5 ( \51817 , \51813 , \47997 );
nor \g131105/U$1 ( \51818 , \51816 , \51817 );
and \g131042/U$3 ( \51819 , \51810 , \51818 );
and \g131042/U$5 ( \51820 , \51802 , \51809 );
or \g131042/U$2 ( \51821 , \51819 , \51820 );
and \g131558/U$2 ( \51822 , \51566 , \51513 );
nor \g131558/U$1 ( \51823 , \51822 , \51567 );
or \g129520/U$2 ( \51824 , \51821 , \51823 );
and \g129545/U$2 ( \51825 , \51821 , \51823 );
and \g129624/U$2 ( \51826 , \47970 , \51053 );
and \g129624/U$3 ( \51827 , \51055 , \47962 );
nor \g129624/U$1 ( \51828 , \51826 , \51827 );
not \g129579/U$3 ( \51829 , \51828 );
not \g129579/U$4 ( \51830 , \50759 );
and \g129579/U$2 ( \51831 , \51829 , \51830 );
and \g129579/U$5 ( \51832 , \51828 , \50759 );
nor \g129579/U$1 ( \51833 , \51831 , \51832 );
nor \g129545/U$1 ( \51834 , \51825 , \51833 );
not \g129544/U$1 ( \51835 , \51834 );
nand \g129520/U$1 ( \51836 , \51824 , \51835 );
and \g130650/U$2 ( \51837 , \48833 , \48858 );
and \g130650/U$3 ( \51838 , \48860 , \48977 );
nor \g130650/U$1 ( \51839 , \51837 , \51838 );
not \g130615/U$3 ( \51840 , \51839 );
not \g130615/U$4 ( \51841 , \48685 );
and \g130615/U$2 ( \51842 , \51840 , \51841 );
and \g130615/U$5 ( \51843 , \51839 , \48685 );
nor \g130615/U$1 ( \51844 , \51842 , \51843 );
and \g131577/U$2 ( \51845 , \51604 , \47960 );
and \g131577/U$3 ( \51846 , \47959 , \51564 );
nor \g131577/U$1 ( \51847 , \51845 , \51846 );
not \g131546/U$3 ( \51848 , \51847 );
not \g131546/U$4 ( \51849 , \47948 );
and \g131546/U$2 ( \51850 , \51848 , \51849 );
and \g131546/U$5 ( \51851 , \51847 , \47948 );
nor \g131546/U$1 ( \51852 , \51850 , \51851 );
not \g131526/U$2 ( \51853 , \51852 );
xor \g131744/U$1 ( \51854 , \47595 , \44897 );
not \g135523/U$2 ( \51855 , \51854 );
nor \g135523/U$1 ( \51856 , \51855 , \40060 );
nand \g131526/U$1 ( \51857 , \51853 , \51856 );
or \g129988/U$2 ( \51858 , \51844 , \51857 );
and \g130003/U$2 ( \51859 , \51844 , \51857 );
and \g130071/U$2 ( \51860 , \48051 , \50159 );
and \g130071/U$3 ( \51861 , \50160 , \48117 );
nor \g130071/U$1 ( \51862 , \51860 , \51861 );
not \g130029/U$3 ( \51863 , \51862 );
not \g130029/U$4 ( \51864 , \49925 );
and \g130029/U$2 ( \51865 , \51863 , \51864 );
and \g130029/U$5 ( \51866 , \51862 , \49925 );
nor \g130029/U$1 ( \51867 , \51865 , \51866 );
nor \g130003/U$1 ( \51868 , \51859 , \51867 );
not \g130002/U$1 ( \51869 , \51868 );
nand \g129988/U$1 ( \51870 , \51858 , \51869 );
xor \g131123/U$1 ( \51871 , \51543 , \51551 );
xor \g131123/U$1_r1 ( \51872 , \51871 , \51560 );
xor \g129688/U$4 ( \51873 , \51870 , \51872 );
and \g130516/U$2 ( \51874 , \48726 , \49075 );
and \g130516/U$3 ( \51875 , \49074 , \48568 );
nor \g130516/U$1 ( \51876 , \51874 , \51875 );
not \g130485/U$3 ( \51877 , \51876 );
not \g130485/U$4 ( \51878 , \49014 );
and \g130485/U$2 ( \51879 , \51877 , \51878 );
and \g130485/U$5 ( \51880 , \51876 , \49014 );
nor \g130485/U$1 ( \51881 , \51879 , \51880 );
not \g131435/U$3 ( \51882 , \51599 );
not \g131435/U$4 ( \51883 , \51605 );
and \g131435/U$2 ( \51884 , \51882 , \51883 );
and \g131435/U$5 ( \51885 , \51599 , \51605 );
nor \g131435/U$1 ( \51886 , \51884 , \51885 );
or \g129809/U$2 ( \51887 , \51881 , \51886 );
and \g129820/U$2 ( \51888 , \51881 , \51886 );
and \g129883/U$2 ( \51889 , \48018 , \50588 );
and \g129883/U$3 ( \51890 , \50587 , \47942 );
nor \g129883/U$1 ( \51891 , \51889 , \51890 );
not \g129850/U$3 ( \51892 , \51891 );
not \g129850/U$4 ( \51893 , \50362 );
and \g129850/U$2 ( \51894 , \51892 , \51893 );
and \g129850/U$5 ( \51895 , \51891 , \50362 );
nor \g129850/U$1 ( \51896 , \51894 , \51895 );
nor \g129820/U$1 ( \51897 , \51888 , \51896 );
not \g129819/U$1 ( \51898 , \51897 );
nand \g129809/U$1 ( \51899 , \51887 , \51898 );
and \g129688/U$3 ( \51900 , \51873 , \51899 );
and \g129688/U$5 ( \51901 , \51870 , \51872 );
or \g129688/U$2 ( \51902 , \51900 , \51901 );
xor \g129287/U$4 ( \51903 , \51836 , \51902 );
xor \g129407/U$1 ( \51904 , \51563 , \51568 );
xor \g129407/U$1_r1 ( \51905 , \51904 , \51577 );
and \g129287/U$3 ( \51906 , \51903 , \51905 );
and \g129287/U$5 ( \51907 , \51836 , \51902 );
or \g129287/U$2 ( \51908 , \51906 , \51907 );
not \g129698/U$3 ( \51909 , \51368 );
not \g129732/U$3 ( \51910 , \51365 );
not \g129732/U$4 ( \51911 , \51391 );
or \g129732/U$2 ( \51912 , \51910 , \51911 );
or \g129732/U$5 ( \51913 , \51391 , \51365 );
nand \g129732/U$1 ( \51914 , \51912 , \51913 );
not \g129698/U$4 ( \51915 , \51914 );
or \g129698/U$2 ( \51916 , \51909 , \51915 );
or \g129698/U$5 ( \51917 , \51914 , \51368 );
nand \g129698/U$1 ( \51918 , \51916 , \51917 );
xor \g455971/U$5 ( \51919 , \51908 , \51918 );
not \g129142/U$3 ( \51920 , \51415 );
not \g129177/U$3 ( \51921 , \51430 );
not \g129177/U$4 ( \51922 , \51424 );
and \g129177/U$2 ( \51923 , \51921 , \51922 );
and \g129177/U$5 ( \51924 , \51430 , \51424 );
nor \g129177/U$1 ( \51925 , \51923 , \51924 );
not \g129142/U$4 ( \51926 , \51925 );
or \g129142/U$2 ( \51927 , \51920 , \51926 );
or \g129142/U$5 ( \51928 , \51925 , \51415 );
nand \g129142/U$1 ( \51929 , \51927 , \51928 );
and \g455971/U$4 ( \51930 , \51919 , \51929 );
and \g455971/U$6 ( \51931 , \51908 , \51918 );
or \g455971/U$3 ( \51932 , \51930 , \51931 );
xor \g128858/U$4 ( \51933 , \51794 , \51932 );
not \g128941/U$3 ( \51934 , \51750 );
xor \g128970/U$1 ( \51935 , \51747 , \51755 );
not \g128941/U$4 ( \51936 , \51935 );
or \g128941/U$2 ( \51937 , \51934 , \51936 );
or \g128941/U$5 ( \51938 , \51935 , \51750 );
nand \g128941/U$1 ( \51939 , \51937 , \51938 );
and \g128858/U$3 ( \51940 , \51933 , \51939 );
and \g128858/U$5 ( \51941 , \51794 , \51932 );
or \g128858/U$2 ( \51942 , \51940 , \51941 );
nand \g128848/U$1 ( \51943 , \51784 , \51942 );
nand \g128844/U$1 ( \51944 , \51781 , \51943 );
xor \g455990/U$2 ( \51945 , \51669 , \51671 );
xor \g455990/U$1 ( \51946 , \51945 , \51674 );
and \g130385/U$2 ( \51947 , \48349 , \49403 );
and \g130385/U$3 ( \51948 , \49405 , \48515 );
nor \g130385/U$1 ( \51949 , \51947 , \51948 );
not \g130339/U$3 ( \51950 , \51949 );
not \g130339/U$4 ( \51951 , \49233 );
and \g130339/U$2 ( \51952 , \51950 , \51951 );
and \g130339/U$5 ( \51953 , \51949 , \49233 );
nor \g130339/U$1 ( \51954 , \51952 , \51953 );
and \g130981/U$2 ( \51955 , \49888 , \48155 );
and \g130981/U$3 ( \51956 , \48154 , \49714 );
nor \g130981/U$1 ( \51957 , \51955 , \51956 );
not \g130957/U$3 ( \51958 , \51957 );
not \g130957/U$4 ( \51959 , \48159 );
and \g130957/U$2 ( \51960 , \51958 , \51959 );
and \g130957/U$5 ( \51961 , \51957 , \48159 );
nor \g130957/U$1 ( \51962 , \51960 , \51961 );
or \g130164/U$2 ( \51963 , \51954 , \51962 );
and \g130178/U$2 ( \51964 , \51954 , \51962 );
and \g130238/U$2 ( \51965 , \48353 , \49813 );
and \g130238/U$3 ( \51966 , \49812 , \48138 );
nor \g130238/U$1 ( \51967 , \51965 , \51966 );
not \g130201/U$3 ( \51968 , \51967 );
not \g130201/U$4 ( \51969 , \49568 );
and \g130201/U$2 ( \51970 , \51968 , \51969 );
and \g130201/U$5 ( \51971 , \51967 , \49568 );
nor \g130201/U$1 ( \51972 , \51970 , \51971 );
nor \g130178/U$1 ( \51973 , \51964 , \51972 );
not \g130177/U$1 ( \51974 , \51973 );
nand \g130164/U$1 ( \51975 , \51963 , \51974 );
xor \g456009/U$9 ( \51976 , \51686 , \51694 );
xor \g456009/U$9_r1 ( \51977 , \51976 , \51703 );
and \g456009/U$8 ( \51978 , \51975 , \51977 );
and \g130754/U$2 ( \51979 , \49102 , \48478 );
and \g130754/U$3 ( \51980 , \48479 , \49158 );
nor \g130754/U$1 ( \51981 , \51979 , \51980 );
not \g130735/U$3 ( \51982 , \51981 );
not \g130735/U$4 ( \51983 , \48483 );
and \g130735/U$2 ( \51984 , \51982 , \51983 );
and \g130735/U$5 ( \51985 , \51981 , \48483 );
nor \g130735/U$1 ( \51986 , \51984 , \51985 );
and \g130872/U$2 ( \51987 , \49512 , \48335 );
and \g130872/U$3 ( \51988 , \48334 , \49282 );
nor \g130872/U$1 ( \51989 , \51987 , \51988 );
not \g130846/U$3 ( \51990 , \51989 );
not \g130846/U$4 ( \51991 , \48323 );
and \g130846/U$2 ( \51992 , \51990 , \51991 );
and \g130846/U$5 ( \51993 , \51989 , \48323 );
nor \g130846/U$1 ( \51994 , \51992 , \51993 );
or \g129635/U$2 ( \51995 , \51986 , \51994 );
and \g129655/U$2 ( \51996 , \51986 , \51994 );
and \g129717/U$2 ( \51997 , \47950 , \51055 );
and \g129717/U$3 ( \51998 , \51053 , \47962 );
nor \g129717/U$1 ( \51999 , \51997 , \51998 );
not \g129683/U$3 ( \52000 , \51999 );
not \g129683/U$4 ( \52001 , \50759 );
and \g129683/U$2 ( \52002 , \52000 , \52001 );
and \g129683/U$5 ( \52003 , \51999 , \50759 );
nor \g129683/U$1 ( \52004 , \52002 , \52003 );
nor \g129655/U$1 ( \52005 , \51996 , \52004 );
not \g129654/U$1 ( \52006 , \52005 );
nand \g129635/U$1 ( \52007 , \51995 , \52006 );
xor \g456009/U$11 ( \52008 , \51686 , \51694 );
xor \g456009/U$11_r1 ( \52009 , \52008 , \51703 );
and \g456009/U$10 ( \52010 , \52007 , \52009 );
and \g456009/U$12 ( \52011 , \51975 , \52007 );
or \g456009/U$7 ( \52012 , \51978 , \52010 , \52011 );
xor \g129287/U$1 ( \52013 , \51836 , \51902 );
xor \g129287/U$1_r1 ( \52014 , \52013 , \51905 );
xor \g455990/U$1_r1 ( \52015 , \52012 , \52014 );
xor \g455990/U$1_r2 ( \52016 , \51946 , \52015 );
not \g128979/U$3 ( \52017 , \52016 );
not \g130169/U$3 ( \52018 , \51972 );
xor \g130296/U$1 ( \52019 , \51962 , \51954 );
not \g130169/U$4 ( \52020 , \52019 );
and \g130169/U$2 ( \52021 , \52018 , \52020 );
and \g130169/U$5 ( \52022 , \51972 , \52019 );
nor \g130169/U$1 ( \52023 , \52021 , \52022 );
not \g131023/U$3 ( \52024 , \48159 );
and \g131063/U$2 ( \52025 , \49888 , \48154 );
and \g131063/U$3 ( \52026 , \48155 , \50019 );
nor \g131063/U$1 ( \52027 , \52025 , \52026 );
not \g131023/U$4 ( \52028 , \52027 );
or \g131023/U$2 ( \52029 , \52024 , \52028 );
or \g131023/U$5 ( \52030 , \52027 , \48159 );
nand \g131023/U$1 ( \52031 , \52029 , \52030 );
not \g130416/U$3 ( \52032 , \49233 );
and \g130444/U$2 ( \52033 , \48568 , \49405 );
and \g130444/U$3 ( \52034 , \49403 , \48515 );
nor \g130444/U$1 ( \52035 , \52033 , \52034 );
not \g130416/U$4 ( \52036 , \52035 );
or \g130416/U$2 ( \52037 , \52032 , \52036 );
or \g130416/U$5 ( \52038 , \52035 , \49233 );
nand \g130416/U$1 ( \52039 , \52037 , \52038 );
xor \g456058/U$4 ( \52040 , \52031 , \52039 );
not \g130273/U$3 ( \52041 , \49568 );
and \g130307/U$2 ( \52042 , \48349 , \49813 );
and \g130307/U$3 ( \52043 , \49812 , \48353 );
nor \g130307/U$1 ( \52044 , \52042 , \52043 );
not \g130273/U$4 ( \52045 , \52044 );
or \g130273/U$2 ( \52046 , \52041 , \52045 );
or \g130273/U$5 ( \52047 , \52044 , \49568 );
nand \g130273/U$1 ( \52048 , \52046 , \52047 );
and \g456058/U$3 ( \52049 , \52040 , \52048 );
and \g456058/U$5 ( \52050 , \52031 , \52039 );
nor \g456058/U$2 ( \52051 , \52049 , \52050 );
or \g129663/U$2 ( \52052 , \52023 , \52051 );
and \g129669/U$2 ( \52053 , \52023 , \52051 );
and \g130820/U$2 ( \52054 , \49282 , \48479 );
and \g130820/U$3 ( \52055 , \48478 , \49158 );
nor \g130820/U$1 ( \52056 , \52054 , \52055 );
not \g130789/U$3 ( \52057 , \52056 );
not \g130789/U$4 ( \52058 , \48483 );
and \g130789/U$2 ( \52059 , \52057 , \52058 );
and \g130789/U$5 ( \52060 , \52056 , \48483 );
nor \g130789/U$1 ( \52061 , \52059 , \52060 );
and \g130928/U$2 ( \52062 , \49512 , \48334 );
and \g130928/U$3 ( \52063 , \48335 , \49714 );
nor \g130928/U$1 ( \52064 , \52062 , \52063 );
not \g130902/U$3 ( \52065 , \52064 );
not \g130902/U$4 ( \52066 , \48323 );
and \g130902/U$2 ( \52067 , \52065 , \52066 );
and \g130902/U$5 ( \52068 , \52064 , \48323 );
nor \g130902/U$1 ( \52069 , \52067 , \52068 );
xor \g129693/U$4 ( \52070 , \52061 , \52069 );
and \g129801/U$2 ( \52071 , \47950 , \51053 );
and \g129801/U$3 ( \52072 , \51055 , \47942 );
nor \g129801/U$1 ( \52073 , \52071 , \52072 );
not \g129756/U$3 ( \52074 , \52073 );
not \g129756/U$4 ( \52075 , \50759 );
and \g129756/U$2 ( \52076 , \52074 , \52075 );
and \g129756/U$5 ( \52077 , \52073 , \50759 );
nor \g129756/U$1 ( \52078 , \52076 , \52077 );
and \g129693/U$3 ( \52079 , \52070 , \52078 );
and \g129693/U$5 ( \52080 , \52061 , \52069 );
or \g129693/U$2 ( \52081 , \52079 , \52080 );
nor \g129669/U$1 ( \52082 , \52053 , \52081 );
not \g129668/U$1 ( \52083 , \52082 );
nand \g129663/U$1 ( \52084 , \52052 , \52083 );
xor \g129688/U$1 ( \52085 , \51870 , \51872 );
xor \g129688/U$1_r1 ( \52086 , \52085 , \51899 );
xor \g129409/U$1 ( \52087 , \52084 , \52086 );
xor \g456009/U$2 ( \52088 , \51686 , \51694 );
xor \g456009/U$1 ( \52089 , \52088 , \51703 );
xor \g456009/U$1_r1 ( \52090 , \51975 , \52007 );
xor \g456009/U$1_r2 ( \52091 , \52089 , \52090 );
xor \g129409/U$1_r1 ( \52092 , \52087 , \52091 );
not \g129408/U$1 ( \52093 , \52092 );
not \g129666/U$3 ( \52094 , \52081 );
xor \g130107/U$1 ( \52095 , \52051 , \52023 );
not \g129666/U$4 ( \52096 , \52095 );
and \g129666/U$2 ( \52097 , \52094 , \52096 );
and \g129666/U$5 ( \52098 , \52081 , \52095 );
nor \g129666/U$1 ( \52099 , \52097 , \52098 );
and \g130705/U$2 ( \52100 , \49102 , \48860 );
and \g130705/U$3 ( \52101 , \48858 , \48977 );
nor \g130705/U$1 ( \52102 , \52100 , \52101 );
not \g130680/U$3 ( \52103 , \52102 );
not \g130680/U$4 ( \52104 , \48685 );
and \g130680/U$2 ( \52105 , \52103 , \52104 );
and \g130680/U$5 ( \52106 , \52102 , \48685 );
nor \g130680/U$1 ( \52107 , \52105 , \52106 );
xor \g131805/U$1 ( \52108 , \47593 , \47592 );
nand \g131771/U$1 ( \52109 , \40061 , \52108 );
not \g131461/U$2 ( \52110 , \52109 );
and \g131509/U$2 ( \52111 , \51564 , \47914 );
and \g131509/U$3 ( \52112 , \47913 , \51098 );
nor \g131509/U$1 ( \52113 , \52111 , \52112 );
and \g131482/U$2 ( \52114 , \52113 , \47977 );
not \g131482/U$4 ( \52115 , \52113 );
and \g131482/U$3 ( \52116 , \52115 , \47976 );
nor \g131482/U$1 ( \52117 , \52114 , \52116 );
nand \g131461/U$1 ( \52118 , \52110 , \52117 );
xor \g130046/U$4 ( \52119 , \52107 , \52118 );
and \g130158/U$2 ( \52120 , \48117 , \50159 );
and \g130158/U$3 ( \52121 , \50160 , \48138 );
nor \g130158/U$1 ( \52122 , \52120 , \52121 );
not \g130120/U$3 ( \52123 , \52122 );
not \g130120/U$4 ( \52124 , \49925 );
and \g130120/U$2 ( \52125 , \52123 , \52124 );
and \g130120/U$5 ( \52126 , \52122 , \49925 );
nor \g130120/U$1 ( \52127 , \52125 , \52126 );
and \g130046/U$3 ( \52128 , \52119 , \52127 );
and \g130046/U$5 ( \52129 , \52107 , \52118 );
or \g130046/U$2 ( \52130 , \52128 , \52129 );
xor \g131042/U$1 ( \52131 , \51802 , \51809 );
xor \g131042/U$1_r1 ( \52132 , \52131 , \51818 );
xor \g129805/U$1 ( \52133 , \52130 , \52132 );
and \g130582/U$2 ( \52134 , \48726 , \49074 );
and \g130582/U$3 ( \52135 , \49075 , \48833 );
nor \g130582/U$1 ( \52136 , \52134 , \52135 );
not \g130553/U$3 ( \52137 , \52136 );
not \g130553/U$4 ( \52138 , \49014 );
and \g130553/U$2 ( \52139 , \52137 , \52138 );
and \g130553/U$5 ( \52140 , \52136 , \49014 );
nor \g130553/U$1 ( \52141 , \52139 , \52140 );
not \g131501/U$3 ( \52142 , \51852 );
not \g131501/U$4 ( \52143 , \51856 );
and \g131501/U$2 ( \52144 , \52142 , \52143 );
and \g131501/U$5 ( \52145 , \51852 , \51856 );
nor \g131501/U$1 ( \52146 , \52144 , \52145 );
xor \g456015/U$5 ( \52147 , \52141 , \52146 );
and \g129979/U$2 ( \52148 , \48051 , \50588 );
and \g129979/U$3 ( \52149 , \50587 , \48018 );
nor \g129979/U$1 ( \52150 , \52148 , \52149 );
not \g129935/U$3 ( \52151 , \52150 );
not \g129935/U$4 ( \52152 , \50362 );
and \g129935/U$2 ( \52153 , \52151 , \52152 );
and \g129935/U$5 ( \52154 , \52150 , \50362 );
nor \g129935/U$1 ( \52155 , \52153 , \52154 );
and \g456015/U$4 ( \52156 , \52147 , \52155 );
and \g456015/U$6 ( \52157 , \52141 , \52146 );
or \g456015/U$3 ( \52158 , \52156 , \52157 );
xor \g129805/U$1_r1 ( \52159 , \52133 , \52158 );
xor \g455978/U$5 ( \52160 , \52099 , \52159 );
and \g130868/U$2 ( \52161 , \49512 , \48479 );
and \g130868/U$3 ( \52162 , \48478 , \49282 );
nor \g130868/U$1 ( \52163 , \52161 , \52162 );
not \g130850/U$3 ( \52164 , \52163 );
not \g130850/U$4 ( \52165 , \48483 );
and \g130850/U$2 ( \52166 , \52164 , \52165 );
and \g130850/U$5 ( \52167 , \52163 , \48483 );
nor \g130850/U$1 ( \52168 , \52166 , \52167 );
and \g130987/U$2 ( \52169 , \49888 , \48335 );
and \g130987/U$3 ( \52170 , \48334 , \49714 );
nor \g130987/U$1 ( \52171 , \52169 , \52170 );
not \g130958/U$3 ( \52172 , \52171 );
not \g130958/U$4 ( \52173 , \48323 );
and \g130958/U$2 ( \52174 , \52172 , \52173 );
and \g130958/U$5 ( \52175 , \52171 , \48323 );
nor \g130958/U$1 ( \52176 , \52174 , \52175 );
or \g130165/U$2 ( \52177 , \52168 , \52176 );
and \g130176/U$2 ( \52178 , \52168 , \52176 );
and \g130239/U$2 ( \52179 , \48353 , \50160 );
and \g130239/U$3 ( \52180 , \50159 , \48138 );
nor \g130239/U$1 ( \52181 , \52179 , \52180 );
not \g130200/U$3 ( \52182 , \52181 );
not \g130200/U$4 ( \52183 , \49925 );
and \g130200/U$2 ( \52184 , \52182 , \52183 );
and \g130200/U$5 ( \52185 , \52181 , \49925 );
nor \g130200/U$1 ( \52186 , \52184 , \52185 );
nor \g130176/U$1 ( \52187 , \52178 , \52186 );
not \g130175/U$1 ( \52188 , \52187 );
nand \g130165/U$1 ( \52189 , \52177 , \52188 );
xor \g456058/U$1 ( \52190 , \52031 , \52039 );
xor \g456058/U$1_r1 ( \52191 , \52190 , \52048 );
and \g129558/U$2 ( \52192 , \52189 , \52191 );
not \g129567/U$3 ( \52193 , \52189 );
not \g129567/U$4 ( \52194 , \52191 );
and \g129567/U$2 ( \52195 , \52193 , \52194 );
not \g130340/U$3 ( \52196 , \49568 );
and \g130380/U$2 ( \52197 , \48349 , \49812 );
and \g130380/U$3 ( \52198 , \49813 , \48515 );
nor \g130380/U$1 ( \52199 , \52197 , \52198 );
not \g130340/U$4 ( \52200 , \52199 );
or \g130340/U$2 ( \52201 , \52196 , \52200 );
or \g130340/U$5 ( \52202 , \52199 , \49568 );
nand \g130340/U$1 ( \52203 , \52201 , \52202 );
not \g129851/U$3 ( \52204 , \50759 );
and \g129884/U$2 ( \52205 , \48018 , \51055 );
and \g129884/U$3 ( \52206 , \51053 , \47942 );
nor \g129884/U$1 ( \52207 , \52205 , \52206 );
not \g129851/U$4 ( \52208 , \52207 );
or \g129851/U$2 ( \52209 , \52204 , \52208 );
or \g129851/U$5 ( \52210 , \52207 , \50759 );
nand \g129851/U$1 ( \52211 , \52209 , \52210 );
xor \g456020/U$4 ( \52212 , \52203 , \52211 );
not \g129684/U$3 ( \52213 , \51124 );
and \g129719/U$2 ( \52214 , \47950 , \51518 );
and \g129719/U$3 ( \52215 , \51517 , \47962 );
nor \g129719/U$1 ( \52216 , \52214 , \52215 );
not \g129684/U$4 ( \52217 , \52216 );
or \g129684/U$2 ( \52218 , \52213 , \52217 );
or \g129684/U$5 ( \52219 , \52216 , \51124 );
nand \g129684/U$1 ( \52220 , \52218 , \52219 );
and \g456020/U$3 ( \52221 , \52212 , \52220 );
and \g456020/U$5 ( \52222 , \52203 , \52211 );
nor \g456020/U$2 ( \52223 , \52221 , \52222 );
nor \g129567/U$1 ( \52224 , \52195 , \52223 );
nor \g129558/U$1 ( \52225 , \52192 , \52224 );
and \g455978/U$4 ( \52226 , \52160 , \52225 );
and \g455978/U$6 ( \52227 , \52099 , \52159 );
or \g455978/U$3 ( \52228 , \52226 , \52227 );
or \g129107/U$2 ( \52229 , \52093 , \52228 );
not \g129112/U$3 ( \52230 , \52228 );
not \g129112/U$4 ( \52231 , \52093 );
or \g129112/U$2 ( \52232 , \52230 , \52231 );
and \g129628/U$2 ( \52233 , \47970 , \51517 );
and \g129628/U$3 ( \52234 , \51518 , \47962 );
nor \g129628/U$1 ( \52235 , \52233 , \52234 );
not \g129582/U$3 ( \52236 , \52235 );
not \g129582/U$4 ( \52237 , \51124 );
and \g129582/U$2 ( \52238 , \52236 , \52237 );
and \g129582/U$5 ( \52239 , \52235 , \51124 );
nor \g129582/U$1 ( \52240 , \52238 , \52239 );
and \g131267/U$2 ( \52241 , \50752 , \48064 );
and \g131267/U$3 ( \52242 , \48063 , \50443 );
nor \g131267/U$1 ( \52243 , \52241 , \52242 );
not \g131235/U$3 ( \52244 , \52243 );
not \g131235/U$4 ( \52245 , \47997 );
and \g131235/U$2 ( \52246 , \52244 , \52245 );
and \g131235/U$5 ( \52247 , \52243 , \47997 );
nor \g131235/U$1 ( \52248 , \52246 , \52247 );
and \g131627/U$2 ( \52249 , \51604 , \47959 );
and \g131627/U$3 ( \52250 , \47960 , \51854 );
nor \g131627/U$1 ( \52251 , \52249 , \52250 );
not \g131598/U$3 ( \52252 , \52251 );
not \g131598/U$4 ( \52253 , \47948 );
and \g131598/U$2 ( \52254 , \52252 , \52253 );
and \g131598/U$5 ( \52255 , \52251 , \47948 );
nor \g131598/U$1 ( \52256 , \52254 , \52255 );
xor \g131043/U$4 ( \52257 , \52248 , \52256 );
and \g131140/U$2 ( \52258 , \50305 , \48155 );
and \g131140/U$3 ( \52259 , \48154 , \50019 );
nor \g131140/U$1 ( \52260 , \52258 , \52259 );
not \g131106/U$3 ( \52261 , \52260 );
not \g131106/U$4 ( \52262 , \48159 );
and \g131106/U$2 ( \52263 , \52261 , \52262 );
and \g131106/U$5 ( \52264 , \52260 , \48159 );
nor \g131106/U$1 ( \52265 , \52263 , \52264 );
and \g131043/U$3 ( \52266 , \52257 , \52265 );
and \g131043/U$5 ( \52267 , \52248 , \52256 );
or \g131043/U$2 ( \52268 , \52266 , \52267 );
xor \g129260/U$4 ( \52269 , \52240 , \52268 );
xor \g135396/U$1 ( \52270 , \24296 , \16306 );
and \g129403/U$2 ( \52271 , \47894 , \52270 );
not \g135570/U$2 ( \52272 , \51120 );
nor \g135570/U$1 ( \52273 , \52272 , \52270 );
and \g129403/U$3 ( \52274 , \52273 , \47972 );
nor \g129403/U$1 ( \52275 , \52271 , \52274 );
not \g129345/U$3 ( \52276 , \52275 );
not \g129345/U$4 ( \52277 , \51120 );
and \g129345/U$2 ( \52278 , \52276 , \52277 );
and \g129345/U$5 ( \52279 , \52275 , \51120 );
nor \g129345/U$1 ( \52280 , \52278 , \52279 );
and \g129260/U$3 ( \52281 , \52269 , \52280 );
and \g129260/U$5 ( \52282 , \52240 , \52268 );
or \g129260/U$2 ( \52283 , \52281 , \52282 );
and \g131443/U$2 ( \52284 , \51117 , \47913 );
and \g131443/U$3 ( \52285 , \47914 , \51098 );
nor \g131443/U$1 ( \52286 , \52284 , \52285 );
and \g131410/U$2 ( \52287 , \52286 , \47977 );
not \g131410/U$4 ( \52288 , \52286 );
and \g131410/U$3 ( \52289 , \52288 , \47976 );
nor \g131410/U$1 ( \52290 , \52287 , \52289 );
not \g131296/U$3 ( \52291 , \47935 );
and \g131320/U$2 ( \52292 , \50957 , \47931 );
and \g131320/U$3 ( \52293 , \47930 , \50752 );
nor \g131320/U$1 ( \52294 , \52292 , \52293 );
not \g131296/U$4 ( \52295 , \52294 );
or \g131296/U$2 ( \52296 , \52291 , \52295 );
or \g131296/U$5 ( \52297 , \52294 , \47935 );
nand \g131296/U$1 ( \52298 , \52296 , \52297 );
xor \g456103/U$1 ( \52299 , \52290 , \52298 );
not \g131182/U$3 ( \52300 , \47997 );
and \g131211/U$2 ( \52301 , \50305 , \48063 );
and \g131211/U$3 ( \52302 , \48064 , \50443 );
nor \g131211/U$1 ( \52303 , \52301 , \52302 );
not \g131182/U$4 ( \52304 , \52303 );
or \g131182/U$2 ( \52305 , \52300 , \52304 );
or \g131182/U$5 ( \52306 , \52303 , \47997 );
nand \g131182/U$1 ( \52307 , \52305 , \52306 );
xor \g456103/U$1_r1 ( \52308 , \52299 , \52307 );
and \g130643/U$2 ( \52309 , \48833 , \49074 );
and \g130643/U$3 ( \52310 , \49075 , \48977 );
nor \g130643/U$1 ( \52311 , \52309 , \52310 );
not \g130617/U$3 ( \52312 , \52311 );
not \g130617/U$4 ( \52313 , \49014 );
and \g130617/U$2 ( \52314 , \52312 , \52313 );
and \g130617/U$5 ( \52315 , \52311 , \49014 );
nor \g130617/U$1 ( \52316 , \52314 , \52315 );
and \g131374/U$2 ( \52317 , \51117 , \47931 );
and \g131374/U$3 ( \52318 , \47930 , \50957 );
nor \g131374/U$1 ( \52319 , \52317 , \52318 );
not \g131355/U$3 ( \52320 , \52319 );
not \g131355/U$4 ( \52321 , \47935 );
and \g131355/U$2 ( \52322 , \52320 , \52321 );
and \g131355/U$5 ( \52323 , \52319 , \47935 );
nor \g131355/U$1 ( \52324 , \52322 , \52323 );
or \g129989/U$2 ( \52325 , \52316 , \52324 );
and \g130005/U$2 ( \52326 , \52316 , \52324 );
and \g130072/U$2 ( \52327 , \48051 , \50587 );
and \g130072/U$3 ( \52328 , \50588 , \48117 );
nor \g130072/U$1 ( \52329 , \52327 , \52328 );
not \g130030/U$3 ( \52330 , \52329 );
not \g130030/U$4 ( \52331 , \50362 );
and \g130030/U$2 ( \52332 , \52330 , \52331 );
and \g130030/U$5 ( \52333 , \52329 , \50362 );
nor \g130030/U$1 ( \52334 , \52332 , \52333 );
nor \g130005/U$1 ( \52335 , \52326 , \52334 );
not \g130004/U$1 ( \52336 , \52335 );
nand \g129989/U$1 ( \52337 , \52325 , \52336 );
xor \g456036/U$4 ( \52338 , \52308 , \52337 );
not \g131436/U$3 ( \52339 , \52117 );
not \g131436/U$4 ( \52340 , \52109 );
and \g131436/U$2 ( \52341 , \52339 , \52340 );
and \g131436/U$5 ( \52342 , \52117 , \52109 );
nor \g131436/U$1 ( \52343 , \52341 , \52342 );
and \g131576/U$2 ( \52344 , \51604 , \47914 );
and \g131576/U$3 ( \52345 , \47913 , \51564 );
nor \g131576/U$1 ( \52346 , \52344 , \52345 );
and \g131547/U$2 ( \52347 , \52346 , \47976 );
not \g131547/U$4 ( \52348 , \52346 );
and \g131547/U$3 ( \52349 , \52348 , \47977 );
nor \g131547/U$1 ( \52350 , \52347 , \52349 );
not \g131529/U$2 ( \52351 , \52350 );
xor \g131866/U$1 ( \52352 , \47590 , \45262 );
not \g135524/U$2 ( \52353 , \52352 );
nor \g135524/U$1 ( \52354 , \52353 , \40060 );
nand \g131529/U$1 ( \52355 , \52351 , \52354 );
or \g130716/U$2 ( \52356 , \52343 , \52355 );
and \g130726/U$2 ( \52357 , \52343 , \52355 );
and \g130757/U$2 ( \52358 , \49102 , \48858 );
and \g130757/U$3 ( \52359 , \48860 , \49158 );
nor \g130757/U$1 ( \52360 , \52358 , \52359 );
not \g130734/U$3 ( \52361 , \52360 );
not \g130734/U$4 ( \52362 , \48685 );
and \g130734/U$2 ( \52363 , \52361 , \52362 );
and \g130734/U$5 ( \52364 , \52360 , \48685 );
nor \g130734/U$1 ( \52365 , \52363 , \52364 );
nor \g130726/U$1 ( \52366 , \52357 , \52365 );
not \g130725/U$1 ( \52367 , \52366 );
nand \g130716/U$1 ( \52368 , \52356 , \52367 );
and \g456036/U$3 ( \52369 , \52338 , \52368 );
and \g456036/U$5 ( \52370 , \52308 , \52337 );
nor \g456036/U$2 ( \52371 , \52369 , \52370 );
or \g129157/U$2 ( \52372 , \52283 , \52371 );
not \g129168/U$3 ( \52373 , \52371 );
not \g129168/U$4 ( \52374 , \52283 );
or \g129168/U$2 ( \52375 , \52373 , \52374 );
and \g129521/U$2 ( \52376 , \47970 , \51518 );
and \g129521/U$3 ( \52377 , \51517 , \47972 );
nor \g129521/U$1 ( \52378 , \52376 , \52377 );
not \g129475/U$3 ( \52379 , \52378 );
not \g129475/U$4 ( \52380 , \51124 );
and \g129475/U$2 ( \52381 , \52379 , \52380 );
and \g129475/U$5 ( \52382 , \52378 , \51124 );
nor \g129475/U$1 ( \52383 , \52381 , \52382 );
not \g129297/U$3 ( \52384 , \52383 );
xor \g456103/U$4 ( \52385 , \52290 , \52298 );
and \g456103/U$3 ( \52386 , \52385 , \52307 );
and \g456103/U$5 ( \52387 , \52290 , \52298 );
nor \g456103/U$2 ( \52388 , \52386 , \52387 );
nand \g129430/U$1 ( \52389 , \52273 , \47894 );
and \g129380/U$5 ( \52390 , \52389 , \51120 );
nor \g129380/U$1 ( \52391 , 1'b0 , \52390 );
xor \g455941/U$1 ( \52392 , \52388 , \52391 );
not \g129297/U$4 ( \52393 , \52392 );
or \g129297/U$2 ( \52394 , \52384 , \52393 );
or \g129297/U$5 ( \52395 , \52392 , \52383 );
nand \g129297/U$1 ( \52396 , \52394 , \52395 );
nand \g129168/U$1 ( \52397 , \52375 , \52396 );
nand \g129157/U$1 ( \52398 , \52372 , \52397 );
nand \g129112/U$1 ( \52399 , \52232 , \52398 );
nand \g129107/U$1 ( \52400 , \52229 , \52399 );
not \g128979/U$4 ( \52401 , \52400 );
or \g128979/U$2 ( \52402 , \52017 , \52401 );
or \g128990/U$2 ( \52403 , \52400 , \52016 );
not \g129321/U$3 ( \52404 , \52383 );
not \g129321/U$4 ( \52405 , \52388 );
and \g129321/U$2 ( \52406 , \52404 , \52405 );
and \g129328/U$2 ( \52407 , \52383 , \52388 );
nor \g129328/U$1 ( \52408 , \52407 , \52391 );
nor \g129321/U$1 ( \52409 , \52406 , \52408 );
not \g129233/U$3 ( \52410 , \52409 );
xor \g129805/U$4 ( \52411 , \52130 , \52132 );
and \g129805/U$3 ( \52412 , \52411 , \52158 );
and \g129805/U$5 ( \52413 , \52130 , \52132 );
or \g129805/U$2 ( \52414 , \52412 , \52413 );
not \g129542/U$3 ( \52415 , \51833 );
xor \g131004/U$1 ( \52416 , \51823 , \51821 );
not \g129542/U$4 ( \52417 , \52416 );
and \g129542/U$2 ( \52418 , \52415 , \52417 );
and \g129542/U$5 ( \52419 , \51833 , \52416 );
nor \g129542/U$1 ( \52420 , \52418 , \52419 );
xor \g129454/U$1 ( \52421 , \52414 , \52420 );
not \g129233/U$4 ( \52422 , \52421 );
and \g129233/U$2 ( \52423 , \52410 , \52422 );
and \g129233/U$5 ( \52424 , \52409 , \52421 );
nor \g129233/U$1 ( \52425 , \52423 , \52424 );
not \g129812/U$3 ( \52426 , \51896 );
xor \g130432/U$1 ( \52427 , \51886 , \51881 );
not \g129812/U$4 ( \52428 , \52427 );
and \g129812/U$2 ( \52429 , \52426 , \52428 );
and \g129812/U$5 ( \52430 , \51896 , \52427 );
nor \g129812/U$1 ( \52431 , \52429 , \52430 );
not \g129995/U$3 ( \52432 , \51867 );
xor \g130573/U$1 ( \52433 , \51857 , \51844 );
not \g129995/U$4 ( \52434 , \52433 );
and \g129995/U$2 ( \52435 , \52432 , \52434 );
and \g129995/U$5 ( \52436 , \51867 , \52433 );
nor \g129995/U$1 ( \52437 , \52435 , \52436 );
xor \g455979/U$5 ( \52438 , \52431 , \52437 );
not \g129643/U$3 ( \52439 , \52004 );
xor \g130697/U$1 ( \52440 , \51994 , \51986 );
not \g129643/U$4 ( \52441 , \52440 );
and \g129643/U$2 ( \52442 , \52439 , \52441 );
and \g129643/U$5 ( \52443 , \52004 , \52440 );
nor \g129643/U$1 ( \52444 , \52442 , \52443 );
and \g455979/U$4 ( \52445 , \52438 , \52444 );
and \g455979/U$6 ( \52446 , \52431 , \52437 );
or \g455979/U$3 ( \52447 , \52445 , \52446 );
or \g129085/U$2 ( \52448 , \52425 , \52447 );
and \g129096/U$2 ( \52449 , \52425 , \52447 );
xor \g129258/U$1 ( \52450 , \51629 , \51637 );
xor \g129258/U$1_r1 ( \52451 , \52450 , \51646 );
xor \g129865/U$1 ( \52452 , \51591 , \51606 );
xor \g129865/U$1_r1 ( \52453 , \52452 , \51615 );
xnor \g455938/U$1 ( \52454 , \52451 , \52453 );
not \g129145/U$3 ( \52455 , \52454 );
xor \g130630/U$1 ( \52456 , \51714 , \51722 );
xor \g130630/U$1_r1 ( \52457 , \52456 , \51731 );
not \g129145/U$4 ( \52458 , \52457 );
and \g129145/U$2 ( \52459 , \52455 , \52458 );
and \g129145/U$5 ( \52460 , \52454 , \52457 );
nor \g129145/U$1 ( \52461 , \52459 , \52460 );
nor \g129096/U$1 ( \52462 , \52449 , \52461 );
not \g129095/U$1 ( \52463 , \52462 );
nand \g129085/U$1 ( \52464 , \52448 , \52463 );
nand \g128990/U$1 ( \52465 , \52403 , \52464 );
nand \g128979/U$1 ( \52466 , \52402 , \52465 );
not \g129197/U$3 ( \52467 , \52457 );
not \g129197/U$4 ( \52468 , \52453 );
or \g129197/U$2 ( \52469 , \52467 , \52468 );
or \g129210/U$2 ( \52470 , \52453 , \52457 );
nand \g129210/U$1 ( \52471 , \52470 , \52451 );
nand \g129197/U$1 ( \52472 , \52469 , \52471 );
xor \g129155/U$1 ( \52473 , \51618 , \51620 );
xor \g129155/U$1_r1 ( \52474 , \52473 , \51649 );
xor \g129014/U$4 ( \52475 , \52472 , \52474 );
xor \g129131/U$1 ( \52476 , \51706 , \51734 );
xor \g129131/U$1_r1 ( \52477 , \52476 , \51741 );
and \g129014/U$3 ( \52478 , \52475 , \52477 );
and \g129014/U$5 ( \52479 , \52472 , \52474 );
or \g129014/U$2 ( \52480 , \52478 , \52479 );
xor \g129054/U$1 ( \52481 , \51580 , \51582 );
xor \g129054/U$1_r1 ( \52482 , \52481 , \51652 );
xor \g455969/U$9 ( \52483 , \52480 , \52482 );
xor \g455980/U$1 ( \52484 , \51667 , \51677 );
xor \g455980/U$1_r1 ( \52485 , \52484 , \51744 );
xor \g455969/U$9_r1 ( \52486 , \52483 , \52485 );
and \g455969/U$8 ( \52487 , \52466 , \52486 );
xor \g455971/U$2 ( \52488 , \51908 , \51918 );
xor \g455971/U$1 ( \52489 , \52488 , \51929 );
xor \g455990/U$9 ( \52490 , \51669 , \51671 );
xor \g455990/U$9_r1 ( \52491 , \52490 , \51674 );
and \g455990/U$8 ( \52492 , \52012 , \52491 );
xor \g455990/U$11 ( \52493 , \51669 , \51671 );
xor \g455990/U$11_r1 ( \52494 , \52493 , \51674 );
and \g455990/U$10 ( \52495 , \52014 , \52494 );
and \g455990/U$12 ( \52496 , \52012 , \52014 );
or \g455990/U$7 ( \52497 , \52492 , \52495 , \52496 );
or \g129222/U$2 ( \52498 , \52420 , \52414 );
and \g129236/U$2 ( \52499 , \52420 , \52414 );
nor \g129236/U$1 ( \52500 , \52499 , \52409 );
not \g129235/U$1 ( \52501 , \52500 );
nand \g129222/U$1 ( \52502 , \52498 , \52501 );
xor \g129409/U$4 ( \52503 , \52084 , \52086 );
and \g129409/U$3 ( \52504 , \52503 , \52091 );
and \g129409/U$5 ( \52505 , \52084 , \52086 );
or \g129409/U$2 ( \52506 , \52504 , \52505 );
xor \g128928/U$4 ( \52507 , \52502 , \52506 );
xor \g129014/U$1 ( \52508 , \52472 , \52474 );
xor \g129014/U$1_r1 ( \52509 , \52508 , \52477 );
and \g128928/U$3 ( \52510 , \52507 , \52509 );
and \g128928/U$5 ( \52511 , \52502 , \52506 );
or \g128928/U$2 ( \52512 , \52510 , \52511 );
xor \g455971/U$1_r1 ( \52513 , \52497 , \52512 );
xor \g455971/U$1_r2 ( \52514 , \52489 , \52513 );
xor \g455969/U$11 ( \52515 , \52480 , \52482 );
xor \g455969/U$11_r1 ( \52516 , \52515 , \52485 );
and \g455969/U$10 ( \52517 , \52514 , \52516 );
and \g455969/U$12 ( \52518 , \52466 , \52514 );
or \g455969/U$7 ( \52519 , \52487 , \52517 , \52518 );
xor \g130046/U$1 ( \52520 , \52107 , \52118 );
xor \g130046/U$1_r1 ( \52521 , \52520 , \52127 );
xor \g456015/U$9 ( \52522 , \52141 , \52146 );
xor \g456015/U$9_r1 ( \52523 , \52522 , \52155 );
and \g456015/U$8 ( \52524 , \52521 , \52523 );
xor \g129693/U$1 ( \52525 , \52061 , \52069 );
xor \g129693/U$1_r1 ( \52526 , \52525 , \52078 );
xor \g456015/U$11 ( \52527 , \52141 , \52146 );
xor \g456015/U$11_r1 ( \52528 , \52527 , \52155 );
and \g456015/U$10 ( \52529 , \52526 , \52528 );
and \g456015/U$12 ( \52530 , \52521 , \52526 );
or \g456015/U$7 ( \52531 , \52524 , \52529 , \52530 );
xor \g455979/U$9 ( \52532 , \52431 , \52437 );
xor \g455979/U$9_r1 ( \52533 , \52532 , \52444 );
and \g455979/U$8 ( \52534 , \52531 , \52533 );
not \g129217/U$3 ( \52535 , \52371 );
not \g129217/U$4 ( \52536 , \52396 );
or \g129217/U$2 ( \52537 , \52535 , \52536 );
or \g129217/U$5 ( \52538 , \52396 , \52371 );
nand \g129217/U$1 ( \52539 , \52537 , \52538 );
not \g129162/U$3 ( \52540 , \52539 );
not \g129162/U$4 ( \52541 , \52283 );
and \g129162/U$2 ( \52542 , \52540 , \52541 );
and \g129162/U$5 ( \52543 , \52539 , \52283 );
nor \g129162/U$1 ( \52544 , \52542 , \52543 );
xor \g455979/U$11 ( \52545 , \52431 , \52437 );
xor \g455979/U$11_r1 ( \52546 , \52545 , \52444 );
and \g455979/U$10 ( \52547 , \52544 , \52546 );
and \g455979/U$12 ( \52548 , \52531 , \52544 );
or \g455979/U$7 ( \52549 , \52534 , \52547 , \52548 );
not \g129552/U$3 ( \52550 , \52191 );
not \g129552/U$4 ( \52551 , \52223 );
or \g129552/U$2 ( \52552 , \52550 , \52551 );
or \g129552/U$5 ( \52553 , \52223 , \52191 );
nand \g129552/U$1 ( \52554 , \52552 , \52553 );
xor \g455944/U$1 ( \52555 , \52189 , \52554 );
and \g129980/U$2 ( \52556 , \48051 , \51055 );
and \g129980/U$3 ( \52557 , \51053 , \48018 );
nor \g129980/U$1 ( \52558 , \52556 , \52557 );
not \g129939/U$3 ( \52559 , \52558 );
not \g129939/U$4 ( \52560 , \50759 );
and \g129939/U$2 ( \52561 , \52559 , \52560 );
and \g129939/U$5 ( \52562 , \52558 , \50759 );
nor \g129939/U$1 ( \52563 , \52561 , \52562 );
and \g130448/U$2 ( \52564 , \48568 , \49813 );
and \g130448/U$3 ( \52565 , \49812 , \48515 );
nor \g130448/U$1 ( \52566 , \52564 , \52565 );
not \g130419/U$3 ( \52567 , \52566 );
not \g130419/U$4 ( \52568 , \49568 );
and \g130419/U$2 ( \52569 , \52567 , \52568 );
and \g130419/U$5 ( \52570 , \52566 , \49568 );
nor \g130419/U$1 ( \52571 , \52569 , \52570 );
xor \g129694/U$4 ( \52572 , \52563 , \52571 );
and \g129803/U$2 ( \52573 , \47950 , \51517 );
and \g129803/U$3 ( \52574 , \51518 , \47942 );
nor \g129803/U$1 ( \52575 , \52573 , \52574 );
not \g129759/U$3 ( \52576 , \52575 );
not \g129759/U$4 ( \52577 , \51124 );
and \g129759/U$2 ( \52578 , \52576 , \52577 );
and \g129759/U$5 ( \52579 , \52575 , \51124 );
nor \g129759/U$1 ( \52580 , \52578 , \52579 );
and \g129694/U$3 ( \52581 , \52572 , \52580 );
and \g129694/U$5 ( \52582 , \52563 , \52571 );
or \g129694/U$2 ( \52583 , \52581 , \52582 );
xor \g131043/U$1 ( \52584 , \52248 , \52256 );
xor \g131043/U$1_r1 ( \52585 , \52584 , \52265 );
or \g129557/U$2 ( \52586 , \52583 , \52585 );
not \g129566/U$3 ( \52587 , \52585 );
not \g129566/U$4 ( \52588 , \52583 );
or \g129566/U$2 ( \52589 , \52587 , \52588 );
xor \g456020/U$1 ( \52590 , \52203 , \52211 );
xor \g456020/U$1_r1 ( \52591 , \52590 , \52220 );
nand \g129566/U$1 ( \52592 , \52589 , \52591 );
nand \g129557/U$1 ( \52593 , \52586 , \52592 );
xor \g456036/U$1 ( \52594 , \52308 , \52337 );
xor \g456036/U$1_r1 ( \52595 , \52594 , \52368 );
or \g129450/U$1 ( \52596 , \52593 , \52595 );
and \g129353/U$2 ( \52597 , \52555 , \52596 );
and \g129353/U$3 ( \52598 , \52595 , \52593 );
nor \g129353/U$1 ( \52599 , \52597 , \52598 );
xor \g455978/U$9 ( \52600 , \52099 , \52159 );
xor \g455978/U$9_r1 ( \52601 , \52600 , \52225 );
and \g455978/U$8 ( \52602 , \52599 , \52601 );
and \g131692/U$2 ( \52603 , \52108 , \47960 );
and \g131692/U$3 ( \52604 , \47959 , \51854 );
nor \g131692/U$1 ( \52605 , \52603 , \52604 );
not \g131660/U$3 ( \52606 , \52605 );
not \g131660/U$4 ( \52607 , \47948 );
and \g131660/U$2 ( \52608 , \52606 , \52607 );
and \g131660/U$5 ( \52609 , \52605 , \47948 );
nor \g131660/U$1 ( \52610 , \52608 , \52609 );
and \g131759/U$2 ( \52611 , \52108 , \47959 );
and \g131759/U$3 ( \52612 , \47960 , \52352 );
nor \g131759/U$1 ( \52613 , \52611 , \52612 );
not \g131728/U$3 ( \52614 , \52613 );
not \g131728/U$4 ( \52615 , \47948 );
and \g131728/U$2 ( \52616 , \52614 , \52615 );
and \g131728/U$5 ( \52617 , \52613 , \47948 );
nor \g131728/U$1 ( \52618 , \52616 , \52617 );
not \g131707/U$2 ( \52619 , \52618 );
xor \g131946/U$1 ( \52620 , \47588 , \47587 );
not \g135525/U$2 ( \52621 , \52620 );
nor \g135525/U$1 ( \52622 , \52621 , \40060 );
nand \g131707/U$1 ( \52623 , \52619 , \52622 );
or \g131155/U$2 ( \52624 , \52610 , \52623 );
and \g131169/U$2 ( \52625 , \52610 , \52623 );
and \g131214/U$2 ( \52626 , \50305 , \48154 );
and \g131214/U$3 ( \52627 , \48155 , \50443 );
nor \g131214/U$1 ( \52628 , \52626 , \52627 );
not \g131184/U$3 ( \52629 , \52628 );
not \g131184/U$4 ( \52630 , \48159 );
and \g131184/U$2 ( \52631 , \52629 , \52630 );
and \g131184/U$5 ( \52632 , \52628 , \48159 );
nor \g131184/U$1 ( \52633 , \52631 , \52632 );
nor \g131169/U$1 ( \52634 , \52625 , \52633 );
not \g131168/U$1 ( \52635 , \52634 );
nand \g131155/U$1 ( \52636 , \52624 , \52635 );
not \g130489/U$3 ( \52637 , \49233 );
and \g130520/U$2 ( \52638 , \48726 , \49405 );
and \g130520/U$3 ( \52639 , \49403 , \48568 );
nor \g130520/U$1 ( \52640 , \52638 , \52639 );
not \g130489/U$4 ( \52641 , \52640 );
or \g130489/U$2 ( \52642 , \52637 , \52641 );
or \g130489/U$5 ( \52643 , \52640 , \49233 );
nand \g130489/U$1 ( \52644 , \52642 , \52643 );
xor \g456002/U$4 ( \52645 , \52636 , \52644 );
not \g129479/U$3 ( \52646 , \51120 );
and \g129522/U$2 ( \52647 , \47970 , \52273 );
and \g129522/U$3 ( \52648 , \52270 , \47972 );
nor \g129522/U$1 ( \52649 , \52647 , \52648 );
not \g129479/U$4 ( \52650 , \52649 );
or \g129479/U$2 ( \52651 , \52646 , \52650 );
or \g129479/U$5 ( \52652 , \52649 , \51120 );
nand \g129479/U$1 ( \52653 , \52651 , \52652 );
and \g456002/U$3 ( \52654 , \52645 , \52653 );
and \g456002/U$5 ( \52655 , \52636 , \52644 );
nor \g456002/U$2 ( \52656 , \52654 , \52655 );
and \g130932/U$2 ( \52657 , \49512 , \48478 );
and \g130932/U$3 ( \52658 , \48479 , \49714 );
nor \g130932/U$1 ( \52659 , \52657 , \52658 );
not \g130904/U$3 ( \52660 , \52659 );
not \g130904/U$4 ( \52661 , \48483 );
and \g130904/U$2 ( \52662 , \52660 , \52661 );
and \g130904/U$5 ( \52663 , \52659 , \48483 );
nor \g130904/U$1 ( \52664 , \52662 , \52663 );
and \g131067/U$2 ( \52665 , \49888 , \48334 );
and \g131067/U$3 ( \52666 , \48335 , \50019 );
nor \g131067/U$1 ( \52667 , \52665 , \52666 );
not \g131026/U$3 ( \52668 , \52667 );
not \g131026/U$4 ( \52669 , \48323 );
and \g131026/U$2 ( \52670 , \52668 , \52669 );
and \g131026/U$5 ( \52671 , \52667 , \48323 );
nor \g131026/U$1 ( \52672 , \52670 , \52671 );
xor \g456017/U$5 ( \52673 , \52664 , \52672 );
and \g130310/U$2 ( \52674 , \48349 , \50160 );
and \g130310/U$3 ( \52675 , \50159 , \48353 );
nor \g130310/U$1 ( \52676 , \52674 , \52675 );
not \g130276/U$3 ( \52677 , \52676 );
not \g130276/U$4 ( \52678 , \49925 );
and \g130276/U$2 ( \52679 , \52677 , \52678 );
and \g130276/U$5 ( \52680 , \52676 , \49925 );
nor \g130276/U$1 ( \52681 , \52679 , \52680 );
and \g456017/U$4 ( \52682 , \52673 , \52681 );
and \g456017/U$6 ( \52683 , \52664 , \52672 );
or \g456017/U$3 ( \52684 , \52682 , \52683 );
and \g130819/U$2 ( \52685 , \49282 , \48860 );
and \g130819/U$3 ( \52686 , \48858 , \49158 );
nor \g130819/U$1 ( \52687 , \52685 , \52686 );
not \g130792/U$3 ( \52688 , \52687 );
not \g130792/U$4 ( \52689 , \48685 );
and \g130792/U$2 ( \52690 , \52688 , \52689 );
and \g130792/U$5 ( \52691 , \52687 , \48685 );
nor \g130792/U$1 ( \52692 , \52690 , \52691 );
not \g131502/U$3 ( \52693 , \52350 );
not \g131502/U$4 ( \52694 , \52354 );
and \g131502/U$2 ( \52695 , \52693 , \52694 );
and \g131502/U$5 ( \52696 , \52350 , \52354 );
nor \g131502/U$1 ( \52697 , \52695 , \52696 );
xor \g130631/U$4 ( \52698 , \52692 , \52697 );
and \g130709/U$2 ( \52699 , \49102 , \49075 );
and \g130709/U$3 ( \52700 , \49074 , \48977 );
nor \g130709/U$1 ( \52701 , \52699 , \52700 );
not \g130683/U$3 ( \52702 , \52701 );
not \g130683/U$4 ( \52703 , \49014 );
and \g130683/U$2 ( \52704 , \52702 , \52703 );
and \g130683/U$5 ( \52705 , \52701 , \49014 );
nor \g130683/U$1 ( \52706 , \52704 , \52705 );
and \g130631/U$3 ( \52707 , \52698 , \52706 );
and \g130631/U$5 ( \52708 , \52692 , \52697 );
or \g130631/U$2 ( \52709 , \52707 , \52708 );
xor \g129983/U$4 ( \52710 , \52684 , \52709 );
and \g131322/U$2 ( \52711 , \50957 , \48064 );
and \g131322/U$3 ( \52712 , \48063 , \50752 );
nor \g131322/U$1 ( \52713 , \52711 , \52712 );
not \g131298/U$3 ( \52714 , \52713 );
not \g131298/U$4 ( \52715 , \47997 );
and \g131298/U$2 ( \52716 , \52714 , \52715 );
and \g131298/U$5 ( \52717 , \52713 , \47997 );
nor \g131298/U$1 ( \52718 , \52716 , \52717 );
and \g131445/U$2 ( \52719 , \51117 , \47930 );
and \g131445/U$3 ( \52720 , \47931 , \51098 );
nor \g131445/U$1 ( \52721 , \52719 , \52720 );
not \g131413/U$3 ( \52722 , \52721 );
not \g131413/U$4 ( \52723 , \47935 );
and \g131413/U$2 ( \52724 , \52722 , \52723 );
and \g131413/U$5 ( \52725 , \52721 , \47935 );
nor \g131413/U$1 ( \52726 , \52724 , \52725 );
xor \g130049/U$4 ( \52727 , \52718 , \52726 );
and \g130161/U$2 ( \52728 , \48117 , \50587 );
and \g130161/U$3 ( \52729 , \50588 , \48138 );
nor \g130161/U$1 ( \52730 , \52728 , \52729 );
not \g130124/U$3 ( \52731 , \52730 );
not \g130124/U$4 ( \52732 , \50362 );
and \g130124/U$2 ( \52733 , \52731 , \52732 );
and \g130124/U$5 ( \52734 , \52730 , \50362 );
nor \g130124/U$1 ( \52735 , \52733 , \52734 );
and \g130049/U$3 ( \52736 , \52727 , \52735 );
and \g130049/U$5 ( \52737 , \52718 , \52726 );
or \g130049/U$2 ( \52738 , \52736 , \52737 );
and \g129983/U$3 ( \52739 , \52710 , \52738 );
and \g129983/U$5 ( \52740 , \52684 , \52709 );
or \g129983/U$2 ( \52741 , \52739 , \52740 );
xor \g129123/U$4 ( \52742 , \52656 , \52741 );
xor \g129260/U$1 ( \52743 , \52240 , \52268 );
xor \g129260/U$1_r1 ( \52744 , \52743 , \52280 );
and \g129123/U$3 ( \52745 , \52742 , \52744 );
and \g129123/U$5 ( \52746 , \52656 , \52741 );
or \g129123/U$2 ( \52747 , \52745 , \52746 );
xor \g455978/U$11 ( \52748 , \52099 , \52159 );
xor \g455978/U$11_r1 ( \52749 , \52748 , \52225 );
and \g455978/U$10 ( \52750 , \52747 , \52749 );
and \g455978/U$12 ( \52751 , \52599 , \52747 );
or \g455978/U$7 ( \52752 , \52602 , \52750 , \52751 );
xor \g128918/U$1 ( \52753 , \52549 , \52752 );
not \g129093/U$3 ( \52754 , \52461 );
xor \g129127/U$1 ( \52755 , \52447 , \52425 );
not \g129093/U$4 ( \52756 , \52755 );
and \g129093/U$2 ( \52757 , \52754 , \52756 );
and \g129093/U$5 ( \52758 , \52461 , \52755 );
nor \g129093/U$1 ( \52759 , \52757 , \52758 );
xor \g128918/U$1_r1 ( \52760 , \52753 , \52759 );
not \g128867/U$3 ( \52761 , \52760 );
not \g129104/U$3 ( \52762 , \52398 );
not \g129104/U$4 ( \52763 , \52228 );
and \g129104/U$2 ( \52764 , \52762 , \52763 );
and \g129104/U$5 ( \52765 , \52398 , \52228 );
nor \g129104/U$1 ( \52766 , \52764 , \52765 );
not \g129060/U$3 ( \52767 , \52766 );
not \g129060/U$4 ( \52768 , \52092 );
and \g129060/U$2 ( \52769 , \52767 , \52768 );
and \g129060/U$5 ( \52770 , \52766 , \52092 );
nor \g129060/U$1 ( \52771 , \52769 , \52770 );
not \g128867/U$4 ( \52772 , \52771 );
and \g128867/U$2 ( \52773 , \52761 , \52772 );
and \g128879/U$2 ( \52774 , \52760 , \52771 );
xor \g456015/U$2 ( \52775 , \52141 , \52146 );
xor \g456015/U$1 ( \52776 , \52775 , \52155 );
xor \g456015/U$1_r1 ( \52777 , \52521 , \52526 );
xor \g456015/U$1_r2 ( \52778 , \52776 , \52777 );
not \g129092/U$3 ( \52779 , \52778 );
not \g130170/U$3 ( \52780 , \52186 );
xor \g130808/U$1 ( \52781 , \52176 , \52168 );
not \g130170/U$4 ( \52782 , \52781 );
and \g130170/U$2 ( \52783 , \52780 , \52782 );
and \g130170/U$5 ( \52784 , \52186 , \52781 );
nor \g130170/U$1 ( \52785 , \52783 , \52784 );
not \g130719/U$3 ( \52786 , \52365 );
xor \g131396/U$1 ( \52787 , \52355 , \52343 );
not \g130719/U$4 ( \52788 , \52787 );
and \g130719/U$2 ( \52789 , \52786 , \52788 );
and \g130719/U$5 ( \52790 , \52365 , \52787 );
nor \g130719/U$1 ( \52791 , \52789 , \52790 );
xor \g129854/U$4 ( \52792 , \52785 , \52791 );
not \g129996/U$3 ( \52793 , \52334 );
xor \g130574/U$1 ( \52794 , \52324 , \52316 );
not \g129996/U$4 ( \52795 , \52794 );
and \g129996/U$2 ( \52796 , \52793 , \52795 );
and \g129996/U$5 ( \52797 , \52334 , \52794 );
nor \g129996/U$1 ( \52798 , \52796 , \52797 );
and \g129854/U$3 ( \52799 , \52792 , \52798 );
and \g129854/U$5 ( \52800 , \52785 , \52791 );
or \g129854/U$2 ( \52801 , \52799 , \52800 );
not \g129092/U$4 ( \52802 , \52801 );
and \g129092/U$2 ( \52803 , \52779 , \52802 );
and \g129101/U$2 ( \52804 , \52778 , \52801 );
xor \g129123/U$1 ( \52805 , \52656 , \52741 );
xor \g129123/U$1_r1 ( \52806 , \52805 , \52744 );
nor \g129101/U$1 ( \52807 , \52804 , \52806 );
nor \g129092/U$1 ( \52808 , \52803 , \52807 );
not \g128959/U$3 ( \52809 , \52808 );
xor \g455978/U$2 ( \52810 , \52099 , \52159 );
xor \g455978/U$1 ( \52811 , \52810 , \52225 );
xor \g455978/U$1_r1 ( \52812 , \52599 , \52747 );
xor \g455978/U$1_r2 ( \52813 , \52811 , \52812 );
not \g128959/U$4 ( \52814 , \52813 );
and \g128959/U$2 ( \52815 , \52809 , \52814 );
and \g128966/U$2 ( \52816 , \52808 , \52813 );
xor \g455979/U$2 ( \52817 , \52431 , \52437 );
xor \g455979/U$1 ( \52818 , \52817 , \52444 );
xor \g455979/U$1_r1 ( \52819 , \52531 , \52544 );
xor \g455979/U$1_r2 ( \52820 , \52818 , \52819 );
nor \g128966/U$1 ( \52821 , \52816 , \52820 );
nor \g128959/U$1 ( \52822 , \52815 , \52821 );
nor \g128879/U$1 ( \52823 , \52774 , \52822 );
nor \g128867/U$1 ( \52824 , \52773 , \52823 );
not \g129554/U$3 ( \52825 , \52585 );
not \g129554/U$4 ( \52826 , \52591 );
or \g129554/U$2 ( \52827 , \52825 , \52826 );
or \g129554/U$5 ( \52828 , \52591 , \52585 );
nand \g129554/U$1 ( \52829 , \52827 , \52828 );
not \g129505/U$3 ( \52830 , \52829 );
not \g129505/U$4 ( \52831 , \52583 );
and \g129505/U$2 ( \52832 , \52830 , \52831 );
and \g129505/U$5 ( \52833 , \52829 , \52583 );
nor \g129505/U$1 ( \52834 , \52832 , \52833 );
not \g129448/U$3 ( \52835 , \52834 );
xor \g129983/U$1 ( \52836 , \52684 , \52709 );
xor \g129983/U$1_r1 ( \52837 , \52836 , \52738 );
and \g130519/U$2 ( \52838 , \48726 , \49813 );
and \g130519/U$3 ( \52839 , \49812 , \48568 );
nor \g130519/U$1 ( \52840 , \52838 , \52839 );
not \g130488/U$3 ( \52841 , \52840 );
not \g130488/U$4 ( \52842 , \49568 );
and \g130488/U$2 ( \52843 , \52841 , \52842 );
and \g130488/U$5 ( \52844 , \52840 , \49568 );
nor \g130488/U$1 ( \52845 , \52843 , \52844 );
and \g130988/U$2 ( \52846 , \49888 , \48479 );
and \g130988/U$3 ( \52847 , \48478 , \49714 );
nor \g130988/U$1 ( \52848 , \52846 , \52847 );
not \g130961/U$3 ( \52849 , \52848 );
not \g130961/U$4 ( \52850 , \48483 );
and \g130961/U$2 ( \52851 , \52849 , \52850 );
and \g130961/U$5 ( \52852 , \52848 , \48483 );
nor \g130961/U$1 ( \52853 , \52851 , \52852 );
xor \g130287/U$4 ( \52854 , \52845 , \52853 );
and \g130383/U$2 ( \52855 , \48349 , \50159 );
and \g130383/U$3 ( \52856 , \50160 , \48515 );
nor \g130383/U$1 ( \52857 , \52855 , \52856 );
not \g130343/U$3 ( \52858 , \52857 );
not \g130343/U$4 ( \52859 , \49925 );
and \g130343/U$2 ( \52860 , \52858 , \52859 );
and \g130343/U$5 ( \52861 , \52857 , \49925 );
nor \g130343/U$1 ( \52862 , \52860 , \52861 );
and \g130287/U$3 ( \52863 , \52854 , \52862 );
and \g130287/U$5 ( \52864 , \52845 , \52853 );
or \g130287/U$2 ( \52865 , \52863 , \52864 );
not \g131161/U$3 ( \52866 , \52633 );
xor \g131621/U$1 ( \52867 , \52623 , \52610 );
not \g131161/U$4 ( \52868 , \52867 );
and \g131161/U$2 ( \52869 , \52866 , \52868 );
and \g131161/U$5 ( \52870 , \52633 , \52867 );
nor \g131161/U$1 ( \52871 , \52869 , \52870 );
xor \g129940/U$4 ( \52872 , \52865 , \52871 );
xor \g130049/U$1 ( \52873 , \52718 , \52726 );
xor \g130049/U$1_r1 ( \52874 , \52873 , \52735 );
and \g129940/U$3 ( \52875 , \52872 , \52874 );
and \g129940/U$5 ( \52876 , \52865 , \52871 );
or \g129940/U$2 ( \52877 , \52875 , \52876 );
xor \g129871/U$1 ( \52878 , \52837 , \52877 );
not \g129448/U$4 ( \52879 , \52878 );
and \g129448/U$2 ( \52880 , \52835 , \52879 );
and \g129448/U$5 ( \52881 , \52834 , \52878 );
nor \g129448/U$1 ( \52882 , \52880 , \52881 );
xor \g132024/U$1 ( \52883 , \47585 , \45593 );
not \g135526/U$2 ( \52884 , \52883 );
nor \g135526/U$1 ( \52885 , \52884 , \40060 );
not \g131751/U$3 ( \52886 , \52885 );
and \g131817/U$2 ( \52887 , \47960 , \52620 );
and \g131817/U$3 ( \52888 , \47959 , \52352 );
nor \g131817/U$1 ( \52889 , \52887 , \52888 );
not \g131790/U$3 ( \52890 , \52889 );
not \g131790/U$4 ( \52891 , \47948 );
and \g131790/U$2 ( \52892 , \52890 , \52891 );
and \g131790/U$5 ( \52893 , \52889 , \47948 );
nor \g131790/U$1 ( \52894 , \52892 , \52893 );
not \g131751/U$4 ( \52895 , \52894 );
or \g131751/U$2 ( \52896 , \52886 , \52895 );
or \g131751/U$5 ( \52897 , \52894 , \52885 );
nand \g131751/U$1 ( \52898 , \52896 , \52897 );
not \g131411/U$3 ( \52899 , \47997 );
and \g131444/U$2 ( \52900 , \51117 , \48063 );
and \g131444/U$3 ( \52901 , \48064 , \51098 );
nor \g131444/U$1 ( \52902 , \52900 , \52901 );
not \g131411/U$4 ( \52903 , \52902 );
or \g131411/U$2 ( \52904 , \52899 , \52903 );
or \g131411/U$5 ( \52905 , \52902 , \47997 );
nand \g131411/U$1 ( \52906 , \52904 , \52905 );
xor \g456104/U$4 ( \52907 , \52898 , \52906 );
not \g131183/U$3 ( \52908 , \48323 );
and \g131212/U$2 ( \52909 , \50305 , \48334 );
and \g131212/U$3 ( \52910 , \48335 , \50443 );
nor \g131212/U$1 ( \52911 , \52909 , \52910 );
not \g131183/U$4 ( \52912 , \52911 );
or \g131183/U$2 ( \52913 , \52908 , \52912 );
or \g131183/U$5 ( \52914 , \52911 , \48323 );
nand \g131183/U$1 ( \52915 , \52913 , \52914 );
and \g456104/U$3 ( \52916 , \52907 , \52915 );
and \g456104/U$5 ( \52917 , \52898 , \52906 );
nor \g456104/U$2 ( \52918 , \52916 , \52917 );
and \g131629/U$2 ( \52919 , \51604 , \47913 );
and \g131629/U$3 ( \52920 , \47914 , \51854 );
nor \g131629/U$1 ( \52921 , \52919 , \52920 );
and \g131600/U$2 ( \52922 , \52921 , \47976 );
not \g131600/U$4 ( \52923 , \52921 );
and \g131600/U$3 ( \52924 , \52923 , \47977 );
nor \g131600/U$1 ( \52925 , \52922 , \52924 );
not \g131772/U$2 ( \52926 , \52894 );
nand \g131772/U$1 ( \52927 , \52926 , \52885 );
xor \g131426/U$1 ( \52928 , \52925 , \52927 );
and \g131511/U$2 ( \52929 , \51564 , \47931 );
and \g131511/U$3 ( \52930 , \47930 , \51098 );
nor \g131511/U$1 ( \52931 , \52929 , \52930 );
not \g131483/U$3 ( \52932 , \52931 );
not \g131483/U$4 ( \52933 , \47935 );
and \g131483/U$2 ( \52934 , \52932 , \52933 );
and \g131483/U$5 ( \52935 , \52931 , \47935 );
nor \g131483/U$1 ( \52936 , \52934 , \52935 );
xor \g131426/U$1_r1 ( \52937 , \52928 , \52936 );
xor \g129630/U$4 ( \52938 , \52918 , \52937 );
not \g131297/U$3 ( \52939 , \48159 );
and \g131321/U$2 ( \52940 , \50957 , \48155 );
and \g131321/U$3 ( \52941 , \48154 , \50752 );
nor \g131321/U$1 ( \52942 , \52940 , \52941 );
not \g131297/U$4 ( \52943 , \52942 );
or \g131297/U$2 ( \52944 , \52939 , \52943 );
or \g131297/U$5 ( \52945 , \52942 , \48159 );
nand \g131297/U$1 ( \52946 , \52944 , \52945 );
not \g130790/U$3 ( \52947 , \49014 );
and \g130818/U$2 ( \52948 , \49282 , \49075 );
and \g130818/U$3 ( \52949 , \49074 , \49158 );
nor \g130818/U$1 ( \52950 , \52948 , \52949 );
not \g130790/U$4 ( \52951 , \52950 );
or \g130790/U$2 ( \52952 , \52947 , \52951 );
or \g130790/U$5 ( \52953 , \52950 , \49014 );
nand \g130790/U$1 ( \52954 , \52952 , \52953 );
xor \g456027/U$4 ( \52955 , \52946 , \52954 );
not \g129758/U$3 ( \52956 , \51120 );
and \g129804/U$2 ( \52957 , \47950 , \52270 );
and \g129804/U$3 ( \52958 , \52273 , \47942 );
nor \g129804/U$1 ( \52959 , \52957 , \52958 );
not \g129758/U$4 ( \52960 , \52959 );
or \g129758/U$2 ( \52961 , \52956 , \52960 );
or \g129758/U$5 ( \52962 , \52959 , \51120 );
nand \g129758/U$1 ( \52963 , \52961 , \52962 );
and \g456027/U$3 ( \52964 , \52955 , \52963 );
and \g456027/U$5 ( \52965 , \52946 , \52954 );
nor \g456027/U$2 ( \52966 , \52964 , \52965 );
and \g129630/U$3 ( \52967 , \52938 , \52966 );
and \g129630/U$5 ( \52968 , \52918 , \52937 );
or \g129630/U$2 ( \52969 , \52967 , \52968 );
and \g130653/U$2 ( \52970 , \48833 , \49403 );
and \g130653/U$3 ( \52971 , \49405 , \48977 );
nor \g130653/U$1 ( \52972 , \52970 , \52971 );
not \g130619/U$3 ( \52973 , \52972 );
not \g130619/U$4 ( \52974 , \49233 );
and \g130619/U$2 ( \52975 , \52973 , \52974 );
and \g130619/U$5 ( \52976 , \52972 , \49233 );
nor \g130619/U$1 ( \52977 , \52975 , \52976 );
xor \g132103/U$1 ( \52978 , \47583 , \47582 );
not \g135527/U$2 ( \52979 , \52978 );
nor \g135527/U$1 ( \52980 , \52979 , \40060 );
and \g131757/U$2 ( \52981 , \52108 , \47913 );
and \g131757/U$3 ( \52982 , \47914 , \52352 );
nor \g131757/U$1 ( \52983 , \52981 , \52982 );
and \g131727/U$2 ( \52984 , \52983 , \47977 );
not \g131727/U$4 ( \52985 , \52983 );
and \g131727/U$3 ( \52986 , \52985 , \47976 );
nor \g131727/U$1 ( \52987 , \52984 , \52986 );
and \g131677/U$2 ( \52988 , \52980 , \52987 );
and \g131691/U$2 ( \52989 , \52108 , \47914 );
and \g131691/U$3 ( \52990 , \47913 , \51854 );
nor \g131691/U$1 ( \52991 , \52989 , \52990 );
and \g131658/U$2 ( \52992 , \52991 , \47977 );
not \g131658/U$4 ( \52993 , \52991 );
and \g131658/U$3 ( \52994 , \52993 , \47976 );
nor \g131658/U$1 ( \52995 , \52992 , \52994 );
xor \g456130/U$4 ( \52996 , \52988 , \52995 );
not \g131548/U$3 ( \52997 , \47935 );
and \g131578/U$2 ( \52998 , \51604 , \47931 );
and \g131578/U$3 ( \52999 , \47930 , \51564 );
nor \g131578/U$1 ( \53000 , \52998 , \52999 );
not \g131548/U$4 ( \53001 , \53000 );
or \g131548/U$2 ( \53002 , \52997 , \53001 );
or \g131548/U$5 ( \53003 , \53000 , \47935 );
nand \g131548/U$1 ( \53004 , \53002 , \53003 );
and \g456130/U$3 ( \53005 , \52996 , \53004 );
and \g456130/U$5 ( \53006 , \52988 , \52995 );
nor \g456130/U$2 ( \53007 , \53005 , \53006 );
xor \g456006/U$5 ( \53008 , \52977 , \53007 );
and \g130074/U$2 ( \53009 , \48051 , \51053 );
and \g130074/U$3 ( \53010 , \51055 , \48117 );
nor \g130074/U$1 ( \53011 , \53009 , \53010 );
not \g130033/U$3 ( \53012 , \53011 );
not \g130033/U$4 ( \53013 , \50759 );
and \g130033/U$2 ( \53014 , \53012 , \53013 );
and \g130033/U$5 ( \53015 , \53011 , \50759 );
nor \g130033/U$1 ( \53016 , \53014 , \53015 );
and \g456006/U$4 ( \53017 , \53008 , \53016 );
and \g456006/U$6 ( \53018 , \52977 , \53007 );
or \g456006/U$3 ( \53019 , \53017 , \53018 );
xor \g455997/U$5 ( \53020 , \52969 , \53019 );
and \g129629/U$2 ( \53021 , \47970 , \52270 );
and \g129629/U$3 ( \53022 , \52273 , \47962 );
nor \g129629/U$1 ( \53023 , \53021 , \53022 );
not \g129585/U$3 ( \53024 , \53023 );
not \g129585/U$4 ( \53025 , \51120 );
and \g129585/U$2 ( \53026 , \53024 , \53025 );
and \g129585/U$5 ( \53027 , \53023 , \51120 );
nor \g129585/U$1 ( \53028 , \53026 , \53027 );
not \g129541/U$3 ( \53029 , \53028 );
xor \g131426/U$4 ( \53030 , \52925 , \52927 );
and \g131426/U$3 ( \53031 , \53030 , \52936 );
and \g131426/U$5 ( \53032 , \52925 , \52927 );
or \g131426/U$2 ( \53033 , \53031 , \53032 );
and \g130586/U$2 ( \53034 , \48726 , \49403 );
and \g130586/U$3 ( \53035 , \49405 , \48833 );
nor \g130586/U$1 ( \53036 , \53034 , \53035 );
not \g130557/U$3 ( \53037 , \53036 );
not \g130557/U$4 ( \53038 , \49233 );
and \g130557/U$2 ( \53039 , \53037 , \53038 );
and \g130557/U$5 ( \53040 , \53036 , \49233 );
nor \g130557/U$1 ( \53041 , \53039 , \53040 );
xor \g130508/U$1 ( \53042 , \53033 , \53041 );
not \g129541/U$4 ( \53043 , \53042 );
and \g129541/U$2 ( \53044 , \53029 , \53043 );
and \g129541/U$5 ( \53045 , \53028 , \53042 );
nor \g129541/U$1 ( \53046 , \53044 , \53045 );
and \g455997/U$4 ( \53047 , \53020 , \53046 );
and \g455997/U$6 ( \53048 , \52969 , \53019 );
or \g455997/U$3 ( \53049 , \53047 , \53048 );
xor \g129262/U$1 ( \53050 , \52882 , \53049 );
not \g131022/U$3 ( \53051 , \48483 );
and \g131064/U$2 ( \53052 , \49888 , \48478 );
and \g131064/U$3 ( \53053 , \48479 , \50019 );
nor \g131064/U$1 ( \53054 , \53052 , \53053 );
not \g131022/U$4 ( \53055 , \53054 );
or \g131022/U$2 ( \53056 , \53051 , \53055 );
or \g131022/U$5 ( \53057 , \53054 , \48483 );
nand \g131022/U$1 ( \53058 , \53056 , \53057 );
not \g130556/U$3 ( \53059 , \49568 );
and \g130585/U$2 ( \53060 , \48726 , \49812 );
and \g130585/U$3 ( \53061 , \49813 , \48833 );
nor \g130585/U$1 ( \53062 , \53060 , \53061 );
not \g130556/U$4 ( \53063 , \53062 );
or \g130556/U$2 ( \53064 , \53059 , \53063 );
or \g130556/U$5 ( \53065 , \53062 , \49568 );
nand \g130556/U$1 ( \53066 , \53064 , \53065 );
xor \g456064/U$4 ( \53067 , \53058 , \53066 );
not \g130418/U$3 ( \53068 , \49925 );
and \g130445/U$2 ( \53069 , \48568 , \50160 );
and \g130445/U$3 ( \53070 , \50159 , \48515 );
nor \g130445/U$1 ( \53071 , \53069 , \53070 );
not \g130418/U$4 ( \53072 , \53071 );
or \g130418/U$2 ( \53073 , \53068 , \53072 );
or \g130418/U$5 ( \53074 , \53071 , \49925 );
nand \g130418/U$1 ( \53075 , \53073 , \53074 );
and \g456064/U$3 ( \53076 , \53067 , \53075 );
and \g456064/U$5 ( \53077 , \53058 , \53066 );
nor \g456064/U$2 ( \53078 , \53076 , \53077 );
and \g131377/U$2 ( \53079 , \51117 , \48064 );
and \g131377/U$3 ( \53080 , \48063 , \50957 );
nor \g131377/U$1 ( \53081 , \53079 , \53080 );
not \g131356/U$3 ( \53082 , \53081 );
not \g131356/U$4 ( \53083 , \47997 );
and \g131356/U$2 ( \53084 , \53082 , \53083 );
and \g131356/U$5 ( \53085 , \53081 , \47997 );
nor \g131356/U$1 ( \53086 , \53084 , \53085 );
not \g131682/U$3 ( \53087 , \52618 );
not \g131682/U$4 ( \53088 , \52622 );
and \g131682/U$2 ( \53089 , \53087 , \53088 );
and \g131682/U$5 ( \53090 , \52618 , \52622 );
nor \g131682/U$1 ( \53091 , \53089 , \53090 );
xor \g131044/U$1 ( \53092 , \53086 , \53091 );
and \g131142/U$2 ( \53093 , \50305 , \48335 );
and \g131142/U$3 ( \53094 , \48334 , \50019 );
nor \g131142/U$1 ( \53095 , \53093 , \53094 );
not \g131108/U$3 ( \53096 , \53095 );
not \g131108/U$4 ( \53097 , \48323 );
and \g131108/U$2 ( \53098 , \53096 , \53097 );
and \g131108/U$5 ( \53099 , \53095 , \48323 );
nor \g131108/U$1 ( \53100 , \53098 , \53099 );
xor \g131044/U$1_r1 ( \53101 , \53092 , \53100 );
xor \g456014/U$5 ( \53102 , \53078 , \53101 );
not \g130903/U$3 ( \53103 , \48685 );
and \g130930/U$2 ( \53104 , \49512 , \48858 );
and \g130930/U$3 ( \53105 , \48860 , \49714 );
nor \g130930/U$1 ( \53106 , \53104 , \53105 );
not \g130903/U$4 ( \53107 , \53106 );
or \g130903/U$2 ( \53108 , \53103 , \53107 );
or \g130903/U$5 ( \53109 , \53106 , \48685 );
nand \g130903/U$1 ( \53110 , \53108 , \53109 );
not \g130275/U$3 ( \53111 , \50362 );
and \g130309/U$2 ( \53112 , \48349 , \50588 );
and \g130309/U$3 ( \53113 , \50587 , \48353 );
nor \g130309/U$1 ( \53114 , \53112 , \53113 );
not \g130275/U$4 ( \53115 , \53114 );
or \g130275/U$2 ( \53116 , \53111 , \53115 );
or \g130275/U$5 ( \53117 , \53114 , \50362 );
nand \g130275/U$1 ( \53118 , \53116 , \53117 );
xor \g456042/U$4 ( \53119 , \53110 , \53118 );
not \g129938/U$3 ( \53120 , \51124 );
and \g129981/U$2 ( \53121 , \48051 , \51518 );
and \g129981/U$3 ( \53122 , \51517 , \48018 );
nor \g129981/U$1 ( \53123 , \53121 , \53122 );
not \g129938/U$4 ( \53124 , \53123 );
or \g129938/U$2 ( \53125 , \53120 , \53124 );
or \g129938/U$5 ( \53126 , \53123 , \51124 );
nand \g129938/U$1 ( \53127 , \53125 , \53126 );
and \g456042/U$3 ( \53128 , \53119 , \53127 );
and \g456042/U$5 ( \53129 , \53110 , \53118 );
nor \g456042/U$2 ( \53130 , \53128 , \53129 );
and \g456014/U$4 ( \53131 , \53102 , \53130 );
and \g456014/U$6 ( \53132 , \53078 , \53101 );
or \g456014/U$3 ( \53133 , \53131 , \53132 );
xor \g129940/U$1 ( \53134 , \52865 , \52871 );
xor \g129940/U$1_r1 ( \53135 , \53134 , \52874 );
xor \g129351/U$4 ( \53136 , \53133 , \53135 );
and \g130231/U$2 ( \53137 , \48353 , \50588 );
and \g130231/U$3 ( \53138 , \50587 , \48138 );
nor \g130231/U$1 ( \53139 , \53137 , \53138 );
not \g130203/U$3 ( \53140 , \53139 );
not \g130203/U$4 ( \53141 , \50362 );
and \g130203/U$2 ( \53142 , \53140 , \53141 );
and \g130203/U$5 ( \53143 , \53139 , \50362 );
nor \g130203/U$1 ( \53144 , \53142 , \53143 );
and \g130874/U$2 ( \53145 , \49512 , \48860 );
and \g130874/U$3 ( \53146 , \48858 , \49282 );
nor \g130874/U$1 ( \53147 , \53145 , \53146 );
not \g130849/U$3 ( \53148 , \53147 );
not \g130849/U$4 ( \53149 , \48685 );
and \g130849/U$2 ( \53150 , \53148 , \53149 );
and \g130849/U$5 ( \53151 , \53147 , \48685 );
nor \g130849/U$1 ( \53152 , \53150 , \53151 );
xor \g456010/U$5 ( \53153 , \53144 , \53152 );
and \g129886/U$2 ( \53154 , \48018 , \51518 );
and \g129886/U$3 ( \53155 , \51517 , \47942 );
nor \g129886/U$1 ( \53156 , \53154 , \53155 );
not \g129842/U$3 ( \53157 , \53156 );
not \g129842/U$4 ( \53158 , \51124 );
and \g129842/U$2 ( \53159 , \53157 , \53158 );
and \g129842/U$5 ( \53160 , \53156 , \51124 );
nor \g129842/U$1 ( \53161 , \53159 , \53160 );
and \g456010/U$4 ( \53162 , \53153 , \53161 );
and \g456010/U$6 ( \53163 , \53144 , \53152 );
or \g456010/U$3 ( \53164 , \53162 , \53163 );
not \g129553/U$3 ( \53165 , \53164 );
and \g130762/U$2 ( \53166 , \49102 , \49074 );
and \g130762/U$3 ( \53167 , \49075 , \49158 );
nor \g130762/U$1 ( \53168 , \53166 , \53167 );
not \g130737/U$3 ( \53169 , \53168 );
not \g130737/U$4 ( \53170 , \49014 );
and \g130737/U$2 ( \53171 , \53169 , \53170 );
and \g130737/U$5 ( \53172 , \53168 , \49014 );
nor \g130737/U$1 ( \53173 , \53171 , \53172 );
and \g131268/U$2 ( \53174 , \50752 , \48155 );
and \g131268/U$3 ( \53175 , \48154 , \50443 );
nor \g131268/U$1 ( \53176 , \53174 , \53175 );
not \g131237/U$3 ( \53177 , \53176 );
not \g131237/U$4 ( \53178 , \48159 );
and \g131237/U$2 ( \53179 , \53177 , \53178 );
and \g131237/U$5 ( \53180 , \53176 , \48159 );
nor \g131237/U$1 ( \53181 , \53179 , \53180 );
or \g129638/U$2 ( \53182 , \53173 , \53181 );
and \g129658/U$2 ( \53183 , \53173 , \53181 );
and \g129720/U$2 ( \53184 , \47950 , \52273 );
and \g129720/U$3 ( \53185 , \52270 , \47962 );
nor \g129720/U$1 ( \53186 , \53184 , \53185 );
not \g129686/U$3 ( \53187 , \53186 );
not \g129686/U$4 ( \53188 , \51120 );
and \g129686/U$2 ( \53189 , \53187 , \53188 );
and \g129686/U$5 ( \53190 , \53186 , \51120 );
nor \g129686/U$1 ( \53191 , \53189 , \53190 );
nor \g129658/U$1 ( \53192 , \53183 , \53191 );
not \g129657/U$1 ( \53193 , \53192 );
nand \g129638/U$1 ( \53194 , \53182 , \53193 );
not \g129553/U$4 ( \53195 , \53194 );
or \g129553/U$2 ( \53196 , \53165 , \53195 );
or \g129553/U$5 ( \53197 , \53194 , \53164 );
nand \g129553/U$1 ( \53198 , \53196 , \53197 );
not \g129504/U$3 ( \53199 , \53198 );
xor \g131044/U$4 ( \53200 , \53086 , \53091 );
and \g131044/U$3 ( \53201 , \53200 , \53100 );
and \g131044/U$5 ( \53202 , \53086 , \53091 );
or \g131044/U$2 ( \53203 , \53201 , \53202 );
not \g129504/U$4 ( \53204 , \53203 );
and \g129504/U$2 ( \53205 , \53199 , \53204 );
and \g129504/U$5 ( \53206 , \53198 , \53203 );
nor \g129504/U$1 ( \53207 , \53205 , \53206 );
and \g129351/U$3 ( \53208 , \53136 , \53207 );
and \g129351/U$5 ( \53209 , \53133 , \53135 );
or \g129351/U$2 ( \53210 , \53208 , \53209 );
xor \g129262/U$1_r1 ( \53211 , \53050 , \53210 );
not \g129261/U$1 ( \53212 , \53211 );
xor \g130287/U$1 ( \53213 , \52845 , \52853 );
xor \g130287/U$1_r1 ( \53214 , \53213 , \52862 );
xor \g456006/U$9 ( \53215 , \52977 , \53007 );
xor \g456006/U$9_r1 ( \53216 , \53215 , \53016 );
and \g456006/U$8 ( \53217 , \53214 , \53216 );
xor \g129630/U$1 ( \53218 , \52918 , \52937 );
xor \g129630/U$1_r1 ( \53219 , \53218 , \52966 );
xor \g456006/U$11 ( \53220 , \52977 , \53007 );
xor \g456006/U$11_r1 ( \53221 , \53220 , \53016 );
and \g456006/U$10 ( \53222 , \53219 , \53221 );
and \g456006/U$12 ( \53223 , \53214 , \53219 );
or \g456006/U$7 ( \53224 , \53217 , \53222 , \53223 );
xor \g456017/U$2 ( \53225 , \52664 , \52672 );
xor \g456017/U$1 ( \53226 , \53225 , \52681 );
xor \g130631/U$1 ( \53227 , \52692 , \52697 );
xor \g130631/U$1_r1 ( \53228 , \53227 , \52706 );
xor \g129694/U$1 ( \53229 , \52563 , \52571 );
xor \g129694/U$1_r1 ( \53230 , \53229 , \52580 );
xor \g456017/U$1_r1 ( \53231 , \53228 , \53230 );
xor \g456017/U$1_r2 ( \53232 , \53226 , \53231 );
xor \g129352/U$1 ( \53233 , \53224 , \53232 );
not \g131599/U$3 ( \53234 , \47935 );
and \g131628/U$2 ( \53235 , \51604 , \47930 );
and \g131628/U$3 ( \53236 , \47931 , \51854 );
nor \g131628/U$1 ( \53237 , \53235 , \53236 );
not \g131599/U$4 ( \53238 , \53237 );
or \g131599/U$2 ( \53239 , \53234 , \53238 );
or \g131599/U$5 ( \53240 , \53237 , \47935 );
nand \g131599/U$1 ( \53241 , \53239 , \53240 );
not \g131854/U$3 ( \53242 , \47948 );
and \g131890/U$2 ( \53243 , \52620 , \47959 );
and \g131890/U$3 ( \53244 , \52883 , \47960 );
nor \g131890/U$1 ( \53245 , \53243 , \53244 );
not \g131854/U$4 ( \53246 , \53245 );
or \g131854/U$2 ( \53247 , \53242 , \53246 );
or \g131854/U$5 ( \53248 , \53245 , \47948 );
nand \g131854/U$1 ( \53249 , \53247 , \53248 );
xor \g131425/U$4 ( \53250 , \53241 , \53249 );
not \g131478/U$3 ( \53251 , \47997 );
and \g131510/U$2 ( \53252 , \51564 , \48064 );
and \g131510/U$3 ( \53253 , \48063 , \51098 );
nor \g131510/U$1 ( \53254 , \53252 , \53253 );
not \g131478/U$4 ( \53255 , \53254 );
or \g131478/U$2 ( \53256 , \53251 , \53255 );
or \g131478/U$5 ( \53257 , \53254 , \47997 );
nand \g131478/U$1 ( \53258 , \53256 , \53257 );
and \g131425/U$3 ( \53259 , \53250 , \53258 );
and \g131425/U$5 ( \53260 , \53241 , \53249 );
or \g131425/U$2 ( \53261 , \53259 , \53260 );
not \g130682/U$3 ( \53262 , \49233 );
and \g130708/U$2 ( \53263 , \49102 , \49405 );
and \g130708/U$3 ( \53264 , \49403 , \48977 );
nor \g130708/U$1 ( \53265 , \53263 , \53264 );
not \g130682/U$4 ( \53266 , \53265 );
or \g130682/U$2 ( \53267 , \53262 , \53266 );
or \g130682/U$5 ( \53268 , \53265 , \49233 );
nand \g130682/U$1 ( \53269 , \53267 , \53268 );
xor \g456051/U$4 ( \53270 , \53261 , \53269 );
not \g130123/U$3 ( \53271 , \50759 );
and \g130160/U$2 ( \53272 , \48117 , \51053 );
and \g130160/U$3 ( \53273 , \51055 , \48138 );
nor \g130160/U$1 ( \53274 , \53272 , \53273 );
not \g130123/U$4 ( \53275 , \53274 );
or \g130123/U$2 ( \53276 , \53271 , \53275 );
or \g130123/U$5 ( \53277 , \53274 , \50759 );
nand \g130123/U$1 ( \53278 , \53276 , \53277 );
and \g456051/U$3 ( \53279 , \53270 , \53278 );
and \g456051/U$5 ( \53280 , \53261 , \53269 );
nor \g456051/U$2 ( \53281 , \53279 , \53280 );
xor \g456010/U$9 ( \53282 , \53144 , \53152 );
xor \g456010/U$9_r1 ( \53283 , \53282 , \53161 );
and \g456010/U$8 ( \53284 , \53281 , \53283 );
not \g129644/U$3 ( \53285 , \53191 );
xor \g130698/U$1 ( \53286 , \53181 , \53173 );
not \g129644/U$4 ( \53287 , \53286 );
and \g129644/U$2 ( \53288 , \53285 , \53287 );
and \g129644/U$5 ( \53289 , \53191 , \53286 );
nor \g129644/U$1 ( \53290 , \53288 , \53289 );
xor \g456010/U$11 ( \53291 , \53144 , \53152 );
xor \g456010/U$11_r1 ( \53292 , \53291 , \53161 );
and \g456010/U$10 ( \53293 , \53290 , \53292 );
and \g456010/U$12 ( \53294 , \53281 , \53290 );
or \g456010/U$7 ( \53295 , \53284 , \53293 , \53294 );
xor \g129352/U$1_r1 ( \53296 , \53233 , \53295 );
xor \g456014/U$2 ( \53297 , \53078 , \53101 );
xor \g456014/U$1 ( \53298 , \53297 , \53130 );
xor \g131677/U$1 ( \53299 , \52980 , \52987 );
xor \g132181/U$1 ( \53300 , \47570 , \47579 );
not \g135528/U$2 ( \53301 , \53300 );
nor \g135528/U$1 ( \53302 , \53301 , \40060 );
and \g131818/U$2 ( \53303 , \52620 , \47914 );
and \g131818/U$3 ( \53304 , \47913 , \52352 );
nor \g131818/U$1 ( \53305 , \53303 , \53304 );
and \g131787/U$2 ( \53306 , \53305 , \47977 );
not \g131787/U$4 ( \53307 , \53305 );
and \g131787/U$3 ( \53308 , \53307 , \47976 );
nor \g131787/U$1 ( \53309 , \53306 , \53308 );
and \g131745/U$2 ( \53310 , \53302 , \53309 );
xor \g131200/U$4 ( \53311 , \53299 , \53310 );
not \g131236/U$3 ( \53312 , \48323 );
and \g131271/U$2 ( \53313 , \50752 , \48335 );
and \g131271/U$3 ( \53314 , \48334 , \50443 );
nor \g131271/U$1 ( \53315 , \53313 , \53314 );
not \g131236/U$4 ( \53316 , \53315 );
or \g131236/U$2 ( \53317 , \53312 , \53316 );
or \g131236/U$5 ( \53318 , \53315 , \48323 );
nand \g131236/U$1 ( \53319 , \53317 , \53318 );
and \g131200/U$3 ( \53320 , \53311 , \53319 );
and \g131200/U$5 ( \53321 , \53299 , \53310 );
or \g131200/U$2 ( \53322 , \53320 , \53321 );
xor \g456130/U$1 ( \53323 , \52988 , \52995 );
xor \g456130/U$1_r1 ( \53324 , \53323 , \53004 );
and \g130780/U$2 ( \53325 , \53322 , \53324 );
not \g130781/U$3 ( \53326 , \53322 );
not \g130781/U$4 ( \53327 , \53324 );
and \g130781/U$2 ( \53328 , \53326 , \53327 );
not \g131352/U$3 ( \53329 , \48159 );
and \g131376/U$2 ( \53330 , \51117 , \48155 );
and \g131376/U$3 ( \53331 , \48154 , \50957 );
nor \g131376/U$1 ( \53332 , \53330 , \53331 );
not \g131352/U$4 ( \53333 , \53332 );
or \g131352/U$2 ( \53334 , \53329 , \53333 );
or \g131352/U$5 ( \53335 , \53332 , \48159 );
nand \g131352/U$1 ( \53336 , \53334 , \53335 );
not \g131107/U$3 ( \53337 , \48483 );
and \g131141/U$2 ( \53338 , \50305 , \48479 );
and \g131141/U$3 ( \53339 , \48478 , \50019 );
nor \g131141/U$1 ( \53340 , \53338 , \53339 );
not \g131107/U$4 ( \53341 , \53340 );
or \g131107/U$2 ( \53342 , \53337 , \53341 );
or \g131107/U$5 ( \53343 , \53340 , \48483 );
nand \g131107/U$1 ( \53344 , \53342 , \53343 );
xor \g456087/U$4 ( \53345 , \53336 , \53344 );
not \g130848/U$3 ( \53346 , \49014 );
and \g130866/U$2 ( \53347 , \49512 , \49075 );
and \g130866/U$3 ( \53348 , \49074 , \49282 );
nor \g130866/U$1 ( \53349 , \53347 , \53348 );
not \g130848/U$4 ( \53350 , \53349 );
or \g130848/U$2 ( \53351 , \53346 , \53350 );
or \g130848/U$5 ( \53352 , \53349 , \49014 );
nand \g130848/U$1 ( \53353 , \53351 , \53352 );
and \g456087/U$3 ( \53354 , \53345 , \53353 );
and \g456087/U$5 ( \53355 , \53336 , \53344 );
nor \g456087/U$2 ( \53356 , \53354 , \53355 );
nor \g130781/U$1 ( \53357 , \53328 , \53356 );
nor \g130780/U$1 ( \53358 , \53325 , \53357 );
not \g130487/U$3 ( \53359 , \49925 );
and \g130518/U$2 ( \53360 , \48726 , \50160 );
and \g130518/U$3 ( \53361 , \50159 , \48568 );
nor \g130518/U$1 ( \53362 , \53360 , \53361 );
not \g130487/U$4 ( \53363 , \53362 );
or \g130487/U$2 ( \53364 , \53359 , \53363 );
or \g130487/U$5 ( \53365 , \53362 , \49925 );
nand \g130487/U$1 ( \53366 , \53364 , \53365 );
not \g130610/U$3 ( \53367 , \49568 );
and \g130652/U$2 ( \53368 , \48833 , \49812 );
and \g130652/U$3 ( \53369 , \49813 , \48977 );
nor \g130652/U$1 ( \53370 , \53368 , \53369 );
not \g130610/U$4 ( \53371 , \53370 );
or \g130610/U$2 ( \53372 , \53367 , \53371 );
or \g130610/U$5 ( \53373 , \53370 , \49568 );
nand \g130610/U$1 ( \53374 , \53372 , \53373 );
xor \g129954/U$4 ( \53375 , \53366 , \53374 );
not \g130032/U$3 ( \53376 , \51124 );
and \g130076/U$2 ( \53377 , \48051 , \51517 );
and \g130076/U$3 ( \53378 , \51518 , \48117 );
nor \g130076/U$1 ( \53379 , \53377 , \53378 );
not \g130032/U$4 ( \53380 , \53379 );
or \g130032/U$2 ( \53381 , \53376 , \53380 );
or \g130032/U$5 ( \53382 , \53379 , \51124 );
nand \g130032/U$1 ( \53383 , \53381 , \53382 );
and \g129954/U$3 ( \53384 , \53375 , \53383 );
and \g129954/U$5 ( \53385 , \53366 , \53374 );
or \g129954/U$2 ( \53386 , \53384 , \53385 );
xor \g456104/U$1 ( \53387 , \52898 , \52906 );
xor \g456104/U$1_r1 ( \53388 , \53387 , \52915 );
and \g129737/U$2 ( \53389 , \53386 , \53388 );
not \g129741/U$3 ( \53390 , \53386 );
not \g129741/U$4 ( \53391 , \53388 );
and \g129741/U$2 ( \53392 , \53390 , \53391 );
not \g130960/U$3 ( \53393 , \48685 );
and \g130985/U$2 ( \53394 , \49888 , \48860 );
and \g130985/U$3 ( \53395 , \48858 , \49714 );
nor \g130985/U$1 ( \53396 , \53394 , \53395 );
not \g130960/U$4 ( \53397 , \53396 );
or \g130960/U$2 ( \53398 , \53393 , \53397 );
or \g130960/U$5 ( \53399 , \53396 , \48685 );
nand \g130960/U$1 ( \53400 , \53398 , \53399 );
not \g130342/U$3 ( \53401 , \50362 );
and \g130381/U$2 ( \53402 , \48349 , \50587 );
and \g130381/U$3 ( \53403 , \50588 , \48515 );
nor \g130381/U$1 ( \53404 , \53402 , \53403 );
not \g130342/U$4 ( \53405 , \53404 );
or \g130342/U$2 ( \53406 , \53401 , \53405 );
or \g130342/U$5 ( \53407 , \53404 , \50362 );
nand \g130342/U$1 ( \53408 , \53406 , \53407 );
xor \g456033/U$4 ( \53409 , \53400 , \53408 );
not \g129853/U$3 ( \53410 , \51120 );
and \g129887/U$2 ( \53411 , \48018 , \52273 );
and \g129887/U$3 ( \53412 , \52270 , \47942 );
nor \g129887/U$1 ( \53413 , \53411 , \53412 );
not \g129853/U$4 ( \53414 , \53413 );
or \g129853/U$2 ( \53415 , \53410 , \53414 );
or \g129853/U$5 ( \53416 , \53413 , \51120 );
nand \g129853/U$1 ( \53417 , \53415 , \53416 );
and \g456033/U$3 ( \53418 , \53409 , \53417 );
and \g456033/U$5 ( \53419 , \53400 , \53408 );
nor \g456033/U$2 ( \53420 , \53418 , \53419 );
nor \g129741/U$1 ( \53421 , \53392 , \53420 );
nor \g129737/U$1 ( \53422 , \53389 , \53421 );
xor \g456014/U$1_r1 ( \53423 , \53358 , \53422 );
xor \g456014/U$1_r2 ( \53424 , \53298 , \53423 );
not \g129487/U$3 ( \53425 , \53424 );
not \g130752/U$3 ( \53426 , \53324 );
not \g130778/U$3 ( \53427 , \53356 );
not \g130778/U$4 ( \53428 , \53322 );
and \g130778/U$2 ( \53429 , \53427 , \53428 );
and \g130778/U$5 ( \53430 , \53356 , \53322 );
nor \g130778/U$1 ( \53431 , \53429 , \53430 );
not \g130752/U$4 ( \53432 , \53431 );
or \g130752/U$2 ( \53433 , \53426 , \53432 );
or \g130752/U$5 ( \53434 , \53431 , \53324 );
nand \g130752/U$1 ( \53435 , \53433 , \53434 );
xor \g456064/U$1 ( \53436 , \53058 , \53066 );
xor \g456064/U$1_r1 ( \53437 , \53436 , \53075 );
xor \g456022/U$4 ( \53438 , \53435 , \53437 );
xor \g456027/U$1 ( \53439 , \52946 , \52954 );
xor \g456027/U$1_r1 ( \53440 , \53439 , \52963 );
and \g456022/U$3 ( \53441 , \53438 , \53440 );
and \g456022/U$5 ( \53442 , \53435 , \53437 );
nor \g456022/U$2 ( \53443 , \53441 , \53442 );
not \g129487/U$4 ( \53444 , \53443 );
and \g129487/U$2 ( \53445 , \53425 , \53444 );
and \g129490/U$2 ( \53446 , \53424 , \53443 );
xor \g456087/U$1 ( \53447 , \53336 , \53344 );
xor \g456087/U$1_r1 ( \53448 , \53447 , \53353 );
not \g130415/U$3 ( \53449 , \50362 );
and \g130447/U$2 ( \53450 , \48568 , \50588 );
and \g130447/U$3 ( \53451 , \50587 , \48515 );
nor \g130447/U$1 ( \53452 , \53450 , \53451 );
not \g130415/U$4 ( \53453 , \53452 );
or \g130415/U$2 ( \53454 , \53449 , \53453 );
or \g130415/U$5 ( \53455 , \53452 , \50362 );
nand \g130415/U$1 ( \53456 , \53454 , \53455 );
not \g131025/U$3 ( \53457 , \48685 );
and \g131066/U$2 ( \53458 , \49888 , \48858 );
and \g131066/U$3 ( \53459 , \48860 , \50019 );
nor \g131066/U$1 ( \53460 , \53458 , \53459 );
not \g131025/U$4 ( \53461 , \53460 );
or \g131025/U$2 ( \53462 , \53457 , \53461 );
or \g131025/U$5 ( \53463 , \53460 , \48685 );
nand \g131025/U$1 ( \53464 , \53462 , \53463 );
xor \g129869/U$4 ( \53465 , \53456 , \53464 );
not \g129937/U$3 ( \53466 , \51120 );
and \g129982/U$2 ( \53467 , \48051 , \52273 );
and \g129982/U$3 ( \53468 , \52270 , \48018 );
nor \g129982/U$1 ( \53469 , \53467 , \53468 );
not \g129937/U$4 ( \53470 , \53469 );
or \g129937/U$2 ( \53471 , \53466 , \53470 );
or \g129937/U$5 ( \53472 , \53469 , \51120 );
nand \g129937/U$1 ( \53473 , \53471 , \53472 );
and \g129869/U$3 ( \53474 , \53465 , \53473 );
and \g129869/U$5 ( \53475 , \53456 , \53464 );
or \g129869/U$2 ( \53476 , \53474 , \53475 );
xor \g456031/U$4 ( \53477 , \53448 , \53476 );
not \g130555/U$3 ( \53478 , \49925 );
and \g130584/U$2 ( \53479 , \48726 , \50159 );
and \g130584/U$3 ( \53480 , \50160 , \48833 );
nor \g130584/U$1 ( \53481 , \53479 , \53480 );
not \g130555/U$4 ( \53482 , \53481 );
or \g130555/U$2 ( \53483 , \53478 , \53482 );
or \g130555/U$5 ( \53484 , \53481 , \49925 );
nand \g130555/U$1 ( \53485 , \53483 , \53484 );
not \g130679/U$3 ( \53486 , \49568 );
and \g130707/U$2 ( \53487 , \49102 , \49813 );
and \g130707/U$3 ( \53488 , \49812 , \48977 );
nor \g130707/U$1 ( \53489 , \53487 , \53488 );
not \g130679/U$4 ( \53490 , \53489 );
or \g130679/U$2 ( \53491 , \53486 , \53490 );
or \g130679/U$5 ( \53492 , \53489 , \49568 );
nand \g130679/U$1 ( \53493 , \53491 , \53492 );
xor \g130048/U$4 ( \53494 , \53485 , \53493 );
not \g130122/U$3 ( \53495 , \51124 );
and \g130162/U$2 ( \53496 , \48117 , \51517 );
and \g130162/U$3 ( \53497 , \51518 , \48138 );
nor \g130162/U$1 ( \53498 , \53496 , \53497 );
not \g130122/U$4 ( \53499 , \53498 );
or \g130122/U$2 ( \53500 , \53495 , \53499 );
or \g130122/U$5 ( \53501 , \53498 , \51124 );
nand \g130122/U$1 ( \53502 , \53500 , \53501 );
and \g130048/U$3 ( \53503 , \53494 , \53502 );
and \g130048/U$5 ( \53504 , \53485 , \53493 );
or \g130048/U$2 ( \53505 , \53503 , \53504 );
and \g456031/U$3 ( \53506 , \53477 , \53505 );
and \g456031/U$5 ( \53507 , \53448 , \53476 );
nor \g456031/U$2 ( \53508 , \53506 , \53507 );
not \g129637/U$3 ( \53509 , \53508 );
xor \g131425/U$1 ( \53510 , \53241 , \53249 );
xor \g131425/U$1_r1 ( \53511 , \53510 , \53258 );
and \g131213/U$2 ( \53512 , \50305 , \48478 );
and \g131213/U$3 ( \53513 , \48479 , \50443 );
nor \g131213/U$1 ( \53514 , \53512 , \53513 );
not \g131176/U$3 ( \53515 , \53514 );
not \g131176/U$4 ( \53516 , \48483 );
and \g131176/U$2 ( \53517 , \53515 , \53516 );
and \g131176/U$5 ( \53518 , \53514 , \48483 );
nor \g131176/U$1 ( \53519 , \53517 , \53518 );
and \g131439/U$2 ( \53520 , \51117 , \48154 );
and \g131439/U$3 ( \53521 , \48155 , \51098 );
nor \g131439/U$1 ( \53522 , \53520 , \53521 );
not \g131412/U$3 ( \53523 , \53522 );
not \g131412/U$4 ( \53524 , \48159 );
and \g131412/U$2 ( \53525 , \53523 , \53524 );
and \g131412/U$5 ( \53526 , \53522 , \48159 );
nor \g131412/U$1 ( \53527 , \53525 , \53526 );
or \g130882/U$2 ( \53528 , \53519 , \53527 );
and \g130892/U$2 ( \53529 , \53519 , \53527 );
and \g130931/U$2 ( \53530 , \49512 , \49074 );
and \g130931/U$3 ( \53531 , \49075 , \49714 );
nor \g130931/U$1 ( \53532 , \53530 , \53531 );
not \g130896/U$3 ( \53533 , \53532 );
not \g130896/U$4 ( \53534 , \49014 );
and \g130896/U$2 ( \53535 , \53533 , \53534 );
and \g130896/U$5 ( \53536 , \53532 , \49014 );
nor \g130896/U$1 ( \53537 , \53535 , \53536 );
nor \g130892/U$1 ( \53538 , \53529 , \53537 );
not \g130891/U$1 ( \53539 , \53538 );
nand \g130882/U$1 ( \53540 , \53528 , \53539 );
xor \g456086/U$4 ( \53541 , \53511 , \53540 );
not \g131659/U$3 ( \53542 , \47935 );
and \g131690/U$2 ( \53543 , \52108 , \47931 );
and \g131690/U$3 ( \53544 , \47930 , \51854 );
nor \g131690/U$1 ( \53545 , \53543 , \53544 );
not \g131659/U$4 ( \53546 , \53545 );
or \g131659/U$2 ( \53547 , \53542 , \53546 );
or \g131659/U$5 ( \53548 , \53545 , \47935 );
nand \g131659/U$1 ( \53549 , \53547 , \53548 );
xor \g131745/U$1 ( \53550 , \53302 , \53309 );
xor \g131252/U$4 ( \53551 , \53549 , \53550 );
not \g131294/U$3 ( \53552 , \48323 );
and \g131319/U$2 ( \53553 , \50957 , \48335 );
and \g131319/U$3 ( \53554 , \48334 , \50752 );
nor \g131319/U$1 ( \53555 , \53553 , \53554 );
not \g131294/U$4 ( \53556 , \53555 );
or \g131294/U$2 ( \53557 , \53552 , \53556 );
or \g131294/U$5 ( \53558 , \53555 , \48323 );
nand \g131294/U$1 ( \53559 , \53557 , \53558 );
and \g131252/U$3 ( \53560 , \53551 , \53559 );
and \g131252/U$5 ( \53561 , \53549 , \53550 );
or \g131252/U$2 ( \53562 , \53560 , \53561 );
and \g456086/U$3 ( \53563 , \53541 , \53562 );
and \g456086/U$5 ( \53564 , \53511 , \53540 );
nor \g456086/U$2 ( \53565 , \53563 , \53564 );
not \g129637/U$4 ( \53566 , \53565 );
and \g129637/U$2 ( \53567 , \53509 , \53566 );
and \g129656/U$2 ( \53568 , \53508 , \53565 );
not \g129733/U$3 ( \53569 , \53388 );
not \g129733/U$4 ( \53570 , \53420 );
or \g129733/U$2 ( \53571 , \53569 , \53570 );
or \g129733/U$5 ( \53572 , \53420 , \53388 );
nand \g129733/U$1 ( \53573 , \53571 , \53572 );
xor \g455946/U$1 ( \53574 , \53386 , \53573 );
not \g129689/U$1 ( \53575 , \53574 );
nor \g129656/U$1 ( \53576 , \53568 , \53575 );
nor \g129637/U$1 ( \53577 , \53567 , \53576 );
nor \g129490/U$1 ( \53578 , \53446 , \53577 );
nor \g129487/U$1 ( \53579 , \53445 , \53578 );
or \g129291/U$2 ( \53580 , \53296 , \53579 );
not \g129299/U$3 ( \53581 , \53579 );
not \g129299/U$4 ( \53582 , \53296 );
or \g129299/U$2 ( \53583 , \53581 , \53582 );
xor \g456010/U$2 ( \53584 , \53144 , \53152 );
xor \g456010/U$1 ( \53585 , \53584 , \53161 );
xor \g456010/U$1_r1 ( \53586 , \53281 , \53290 );
xor \g456010/U$1_r2 ( \53587 , \53585 , \53586 );
xor \g456006/U$2 ( \53588 , \52977 , \53007 );
xor \g456006/U$1 ( \53589 , \53588 , \53016 );
xor \g456006/U$1_r1 ( \53590 , \53214 , \53219 );
xor \g456006/U$1_r2 ( \53591 , \53589 , \53590 );
xor \g455999/U$4 ( \53592 , \53587 , \53591 );
not \g130738/U$3 ( \53593 , \49233 );
and \g130763/U$2 ( \53594 , \49102 , \49403 );
and \g130763/U$3 ( \53595 , \49405 , \49158 );
nor \g130763/U$1 ( \53596 , \53594 , \53595 );
not \g130738/U$4 ( \53597 , \53596 );
or \g130738/U$2 ( \53598 , \53593 , \53597 );
or \g130738/U$5 ( \53599 , \53596 , \49233 );
nand \g130738/U$1 ( \53600 , \53598 , \53599 );
and \g132047/U$2 ( \53601 , \47959 , \52978 );
and \g132047/U$3 ( \53602 , \53300 , \47960 );
nor \g132047/U$1 ( \53603 , \53601 , \53602 );
not \g132008/U$3 ( \53604 , \53603 );
not \g132008/U$4 ( \53605 , \47948 );
and \g132008/U$2 ( \53606 , \53604 , \53605 );
and \g132008/U$5 ( \53607 , \53603 , \47948 );
nor \g132008/U$1 ( \53608 , \53606 , \53607 );
not \g131989/U$2 ( \53609 , \53608 );
xor \g132265/U$1 ( \53610 , \47567 , \47544 );
not \g135529/U$2 ( \53611 , \53610 );
nor \g135529/U$1 ( \53612 , \53611 , \40060 );
nand \g131989/U$1 ( \53613 , \53609 , \53612 );
and \g131962/U$2 ( \53614 , \47960 , \52978 );
and \g131962/U$3 ( \53615 , \47959 , \52883 );
nor \g131962/U$1 ( \53616 , \53614 , \53615 );
not \g131927/U$3 ( \53617 , \53616 );
not \g131927/U$4 ( \53618 , \47948 );
and \g131927/U$2 ( \53619 , \53617 , \53618 );
and \g131927/U$5 ( \53620 , \53616 , \47948 );
nor \g131927/U$1 ( \53621 , \53619 , \53620 );
or \g131522/U$2 ( \53622 , \53613 , \53621 );
and \g131532/U$2 ( \53623 , \53613 , \53621 );
and \g131579/U$2 ( \53624 , \51604 , \48064 );
and \g131579/U$3 ( \53625 , \48063 , \51564 );
nor \g131579/U$1 ( \53626 , \53624 , \53625 );
not \g131549/U$3 ( \53627 , \53626 );
not \g131549/U$4 ( \53628 , \47997 );
and \g131549/U$2 ( \53629 , \53627 , \53628 );
and \g131549/U$5 ( \53630 , \53626 , \47997 );
nor \g131549/U$1 ( \53631 , \53629 , \53630 );
nor \g131532/U$1 ( \53632 , \53623 , \53631 );
not \g131531/U$1 ( \53633 , \53632 );
nand \g131522/U$1 ( \53634 , \53622 , \53633 );
xor \g130138/U$4 ( \53635 , \53600 , \53634 );
not \g130204/U$3 ( \53636 , \50759 );
and \g130241/U$2 ( \53637 , \48353 , \51055 );
and \g130241/U$3 ( \53638 , \51053 , \48138 );
nor \g130241/U$1 ( \53639 , \53637 , \53638 );
not \g130204/U$4 ( \53640 , \53639 );
or \g130204/U$2 ( \53641 , \53636 , \53640 );
or \g130204/U$5 ( \53642 , \53639 , \50759 );
nand \g130204/U$1 ( \53643 , \53641 , \53642 );
and \g130138/U$3 ( \53644 , \53635 , \53643 );
and \g130138/U$5 ( \53645 , \53600 , \53634 );
or \g130138/U$2 ( \53646 , \53644 , \53645 );
xor \g456051/U$1 ( \53647 , \53261 , \53269 );
xor \g456051/U$1_r1 ( \53648 , \53647 , \53278 );
xor \g456035/U$4 ( \53649 , \53646 , \53648 );
xor \g456042/U$1 ( \53650 , \53110 , \53118 );
xor \g456042/U$1_r1 ( \53651 , \53650 , \53127 );
and \g456035/U$3 ( \53652 , \53649 , \53651 );
and \g456035/U$5 ( \53653 , \53646 , \53648 );
nor \g456035/U$2 ( \53654 , \53652 , \53653 );
and \g455999/U$3 ( \53655 , \53592 , \53654 );
and \g455999/U$5 ( \53656 , \53587 , \53591 );
nor \g455999/U$2 ( \53657 , \53655 , \53656 );
nand \g129299/U$1 ( \53658 , \53583 , \53657 );
nand \g129291/U$1 ( \53659 , \53580 , \53658 );
and \g129019/U$2 ( \53660 , \53212 , \53659 );
not \g129021/U$3 ( \53661 , \53212 );
not \g129021/U$4 ( \53662 , \53659 );
and \g129021/U$2 ( \53663 , \53661 , \53662 );
xor \g456014/U$9 ( \53664 , \53078 , \53101 );
xor \g456014/U$9_r1 ( \53665 , \53664 , \53130 );
and \g456014/U$8 ( \53666 , \53358 , \53665 );
xor \g456014/U$11 ( \53667 , \53078 , \53101 );
xor \g456014/U$11_r1 ( \53668 , \53667 , \53130 );
and \g456014/U$10 ( \53669 , \53422 , \53668 );
and \g456014/U$12 ( \53670 , \53358 , \53422 );
or \g456014/U$7 ( \53671 , \53666 , \53669 , \53670 );
xor \g455997/U$9 ( \53672 , \52969 , \53019 );
xor \g455997/U$9_r1 ( \53673 , \53672 , \53046 );
and \g455997/U$8 ( \53674 , \53671 , \53673 );
xor \g129351/U$1 ( \53675 , \53133 , \53135 );
xor \g129351/U$1_r1 ( \53676 , \53675 , \53207 );
xor \g455997/U$11 ( \53677 , \52969 , \53019 );
xor \g455997/U$11_r1 ( \53678 , \53677 , \53046 );
and \g455997/U$10 ( \53679 , \53676 , \53678 );
and \g455997/U$12 ( \53680 , \53671 , \53676 );
or \g455997/U$7 ( \53681 , \53674 , \53679 , \53680 );
xor \g129352/U$4 ( \53682 , \53224 , \53232 );
and \g129352/U$3 ( \53683 , \53682 , \53295 );
and \g129352/U$5 ( \53684 , \53224 , \53232 );
or \g129352/U$2 ( \53685 , \53683 , \53684 );
xor \g129055/U$1 ( \53686 , \53681 , \53685 );
xor \g129854/U$1 ( \53687 , \52785 , \52791 );
xor \g129854/U$1_r1 ( \53688 , \53687 , \52798 );
not \g129246/U$3 ( \53689 , \53688 );
or \g129535/U$2 ( \53690 , \53041 , \53033 );
and \g129551/U$2 ( \53691 , \53041 , \53033 );
nor \g129551/U$1 ( \53692 , \53691 , \53028 );
not \g129550/U$1 ( \53693 , \53692 );
nand \g129535/U$1 ( \53694 , \53690 , \53693 );
or \g129559/U$2 ( \53695 , \53164 , \53203 );
not \g129568/U$3 ( \53696 , \53203 );
not \g129568/U$4 ( \53697 , \53164 );
or \g129568/U$2 ( \53698 , \53696 , \53697 );
nand \g129568/U$1 ( \53699 , \53698 , \53194 );
nand \g129559/U$1 ( \53700 , \53695 , \53699 );
xor \g129288/U$1 ( \53701 , \53694 , \53700 );
xor \g456002/U$1 ( \53702 , \52636 , \52644 );
xor \g456002/U$1_r1 ( \53703 , \53702 , \52653 );
xor \g129288/U$1_r1 ( \53704 , \53701 , \53703 );
not \g129246/U$4 ( \53705 , \53704 );
or \g129246/U$2 ( \53706 , \53689 , \53705 );
or \g129246/U$5 ( \53707 , \53704 , \53688 );
nand \g129246/U$1 ( \53708 , \53706 , \53707 );
not \g129200/U$3 ( \53709 , \53708 );
xor \g456017/U$9 ( \53710 , \52664 , \52672 );
xor \g456017/U$9_r1 ( \53711 , \53710 , \52681 );
and \g456017/U$8 ( \53712 , \53228 , \53711 );
xor \g456017/U$11 ( \53713 , \52664 , \52672 );
xor \g456017/U$11_r1 ( \53714 , \53713 , \52681 );
and \g456017/U$10 ( \53715 , \53230 , \53714 );
and \g456017/U$12 ( \53716 , \53228 , \53230 );
or \g456017/U$7 ( \53717 , \53712 , \53715 , \53716 );
not \g129200/U$4 ( \53718 , \53717 );
and \g129200/U$2 ( \53719 , \53709 , \53718 );
and \g129200/U$5 ( \53720 , \53708 , \53717 );
nor \g129200/U$1 ( \53721 , \53719 , \53720 );
xor \g129055/U$1_r1 ( \53722 , \53686 , \53721 );
nor \g129021/U$1 ( \53723 , \53663 , \53722 );
nor \g129019/U$1 ( \53724 , \53660 , \53723 );
not \g128988/U$3 ( \53725 , \53211 );
not \g129002/U$3 ( \53726 , \53659 );
not \g129002/U$4 ( \53727 , \53722 );
or \g129002/U$2 ( \53728 , \53726 , \53727 );
or \g129002/U$5 ( \53729 , \53722 , \53659 );
nand \g129002/U$1 ( \53730 , \53728 , \53729 );
not \g128988/U$4 ( \53731 , \53730 );
or \g128988/U$2 ( \53732 , \53725 , \53731 );
or \g128988/U$5 ( \53733 , \53730 , \53211 );
nand \g128988/U$1 ( \53734 , \53732 , \53733 );
not \g129313/U$3 ( \53735 , \53579 );
not \g129313/U$4 ( \53736 , \53657 );
or \g129313/U$2 ( \53737 , \53735 , \53736 );
or \g129313/U$5 ( \53738 , \53657 , \53579 );
nand \g129313/U$1 ( \53739 , \53737 , \53738 );
not \g129296/U$3 ( \53740 , \53739 );
not \g129296/U$4 ( \53741 , \53296 );
and \g129296/U$2 ( \53742 , \53740 , \53741 );
and \g129296/U$5 ( \53743 , \53739 , \53296 );
nor \g129296/U$1 ( \53744 , \53742 , \53743 );
not \g130962/U$3 ( \53745 , \49014 );
and \g130989/U$2 ( \53746 , \49888 , \49075 );
and \g130989/U$3 ( \53747 , \49074 , \49714 );
nor \g130989/U$1 ( \53748 , \53746 , \53747 );
not \g130962/U$4 ( \53749 , \53748 );
or \g130962/U$2 ( \53750 , \53745 , \53749 );
or \g130962/U$5 ( \53751 , \53748 , \49014 );
nand \g130962/U$1 ( \53752 , \53750 , \53751 );
not \g130490/U$3 ( \53753 , \50362 );
and \g130521/U$2 ( \53754 , \48726 , \50588 );
and \g130521/U$3 ( \53755 , \50587 , \48568 );
nor \g130521/U$1 ( \53756 , \53754 , \53755 );
not \g130490/U$4 ( \53757 , \53756 );
or \g130490/U$2 ( \53758 , \53753 , \53757 );
or \g130490/U$5 ( \53759 , \53756 , \50362 );
nand \g130490/U$1 ( \53760 , \53758 , \53759 );
xor \g456053/U$4 ( \53761 , \53752 , \53760 );
not \g130205/U$3 ( \53762 , \51124 );
and \g130242/U$2 ( \53763 , \48353 , \51518 );
and \g130242/U$3 ( \53764 , \51517 , \48138 );
nor \g130242/U$1 ( \53765 , \53763 , \53764 );
not \g130205/U$4 ( \53766 , \53765 );
or \g130205/U$2 ( \53767 , \53762 , \53766 );
or \g130205/U$5 ( \53768 , \53765 , \51124 );
nand \g130205/U$1 ( \53769 , \53767 , \53768 );
and \g456053/U$3 ( \53770 , \53761 , \53769 );
and \g456053/U$5 ( \53771 , \53752 , \53760 );
nor \g456053/U$2 ( \53772 , \53770 , \53771 );
not \g130885/U$3 ( \53773 , \53537 );
xor \g131133/U$1 ( \53774 , \53527 , \53519 );
not \g130885/U$4 ( \53775 , \53774 );
and \g130885/U$2 ( \53776 , \53773 , \53775 );
and \g130885/U$5 ( \53777 , \53537 , \53774 );
nor \g130885/U$1 ( \53778 , \53776 , \53777 );
or \g129918/U$2 ( \53779 , \53772 , \53778 );
not \g129923/U$3 ( \53780 , \53778 );
not \g129923/U$4 ( \53781 , \53772 );
or \g129923/U$2 ( \53782 , \53780 , \53781 );
not \g130620/U$3 ( \53783 , \49925 );
and \g130654/U$2 ( \53784 , \48833 , \50159 );
and \g130654/U$3 ( \53785 , \50160 , \48977 );
nor \g130654/U$1 ( \53786 , \53784 , \53785 );
not \g130620/U$4 ( \53787 , \53786 );
or \g130620/U$2 ( \53788 , \53783 , \53787 );
or \g130620/U$5 ( \53789 , \53786 , \49925 );
nand \g130620/U$1 ( \53790 , \53788 , \53789 );
not \g130739/U$3 ( \53791 , \49568 );
and \g130764/U$2 ( \53792 , \49102 , \49812 );
and \g130764/U$3 ( \53793 , \49813 , \49158 );
nor \g130764/U$1 ( \53794 , \53792 , \53793 );
not \g130739/U$4 ( \53795 , \53794 );
or \g130739/U$2 ( \53796 , \53791 , \53795 );
or \g130739/U$5 ( \53797 , \53794 , \49568 );
nand \g130739/U$1 ( \53798 , \53796 , \53797 );
xor \g129958/U$4 ( \53799 , \53790 , \53798 );
not \g130034/U$3 ( \53800 , \51120 );
and \g130077/U$2 ( \53801 , \48051 , \52270 );
and \g130077/U$3 ( \53802 , \52273 , \48117 );
nor \g130077/U$1 ( \53803 , \53801 , \53802 );
not \g130034/U$4 ( \53804 , \53803 );
or \g130034/U$2 ( \53805 , \53800 , \53804 );
or \g130034/U$5 ( \53806 , \53803 , \51120 );
nand \g130034/U$1 ( \53807 , \53805 , \53806 );
and \g129958/U$3 ( \53808 , \53799 , \53807 );
and \g129958/U$5 ( \53809 , \53790 , \53798 );
or \g129958/U$2 ( \53810 , \53808 , \53809 );
nand \g129923/U$1 ( \53811 , \53782 , \53810 );
nand \g129918/U$1 ( \53812 , \53779 , \53811 );
xor \g456086/U$1 ( \53813 , \53511 , \53540 );
xor \g456086/U$1_r1 ( \53814 , \53813 , \53562 );
xor \g129695/U$4 ( \53815 , \53812 , \53814 );
xor \g456031/U$1 ( \53816 , \53448 , \53476 );
xor \g456031/U$1_r1 ( \53817 , \53816 , \53505 );
and \g129695/U$3 ( \53818 , \53815 , \53817 );
and \g129695/U$5 ( \53819 , \53812 , \53814 );
or \g129695/U$2 ( \53820 , \53818 , \53819 );
xor \g456022/U$1 ( \53821 , \53435 , \53437 );
xor \g456022/U$1_r1 ( \53822 , \53821 , \53440 );
xor \g456007/U$4 ( \53823 , \53820 , \53822 );
not \g129589/U$3 ( \53824 , \53565 );
not \g129613/U$3 ( \53825 , \53508 );
not \g129613/U$4 ( \53826 , \53574 );
or \g129613/U$2 ( \53827 , \53825 , \53826 );
or \g129613/U$5 ( \53828 , \53574 , \53508 );
nand \g129613/U$1 ( \53829 , \53827 , \53828 );
not \g129589/U$4 ( \53830 , \53829 );
or \g129589/U$2 ( \53831 , \53824 , \53830 );
or \g129589/U$5 ( \53832 , \53829 , \53565 );
nand \g129589/U$1 ( \53833 , \53831 , \53832 );
and \g456007/U$3 ( \53834 , \53823 , \53833 );
and \g456007/U$5 ( \53835 , \53820 , \53822 );
nor \g456007/U$2 ( \53836 , \53834 , \53835 );
not \g130794/U$3 ( \53837 , \49233 );
and \g130821/U$2 ( \53838 , \49282 , \49405 );
and \g130821/U$3 ( \53839 , \49403 , \49158 );
nor \g130821/U$1 ( \53840 , \53838 , \53839 );
not \g130794/U$4 ( \53841 , \53840 );
or \g130794/U$2 ( \53842 , \53837 , \53841 );
or \g130794/U$5 ( \53843 , \53840 , \49233 );
nand \g130794/U$1 ( \53844 , \53842 , \53843 );
and \g132387/U$2 ( \53845 , \47541 , \47505 );
not \g132387/U$4 ( \53846 , \47541 );
and \g132387/U$3 ( \53847 , \53846 , \47506 );
or \g132387/U$1 ( \53848 , \53845 , \53847 );
not \g135530/U$2 ( \53849 , \53848 );
nor \g135530/U$1 ( \53850 , \53849 , \40060 );
not \g132088/U$3 ( \53851 , \47948 );
and \g132128/U$2 ( \53852 , \47960 , \53610 );
and \g132128/U$3 ( \53853 , \53300 , \47959 );
nor \g132128/U$1 ( \53854 , \53852 , \53853 );
not \g132088/U$4 ( \53855 , \53854 );
or \g132088/U$2 ( \53856 , \53851 , \53855 );
or \g132088/U$5 ( \53857 , \53854 , \47948 );
nand \g132088/U$1 ( \53858 , \53856 , \53857 );
and \g132029/U$2 ( \53859 , \53850 , \53858 );
and \g131893/U$2 ( \53860 , \52620 , \47913 );
and \g131893/U$3 ( \53861 , \47914 , \52883 );
nor \g131893/U$1 ( \53862 , \53860 , \53861 );
and \g131855/U$2 ( \53863 , \53862 , \47977 );
not \g131855/U$4 ( \53864 , \53862 );
and \g131855/U$3 ( \53865 , \53864 , \47976 );
nor \g131855/U$1 ( \53866 , \53863 , \53865 );
xor \g131675/U$4 ( \53867 , \53859 , \53866 );
not \g131729/U$3 ( \53868 , \47935 );
and \g131760/U$2 ( \53869 , \52108 , \47930 );
and \g131760/U$3 ( \53870 , \47931 , \52352 );
nor \g131760/U$1 ( \53871 , \53869 , \53870 );
not \g131729/U$4 ( \53872 , \53871 );
or \g131729/U$2 ( \53873 , \53868 , \53872 );
or \g131729/U$5 ( \53874 , \53871 , \47935 );
nand \g131729/U$1 ( \53875 , \53873 , \53874 );
and \g131675/U$3 ( \53876 , \53867 , \53875 );
and \g131675/U$5 ( \53877 , \53859 , \53866 );
or \g131675/U$2 ( \53878 , \53876 , \53877 );
xor \g130216/U$4 ( \53879 , \53844 , \53878 );
not \g130277/U$3 ( \53880 , \50759 );
and \g130311/U$2 ( \53881 , \48349 , \51055 );
and \g130311/U$3 ( \53882 , \51053 , \48353 );
nor \g130311/U$1 ( \53883 , \53881 , \53882 );
not \g130277/U$4 ( \53884 , \53883 );
or \g130277/U$2 ( \53885 , \53880 , \53884 );
or \g130277/U$5 ( \53886 , \53883 , \50759 );
nand \g130277/U$1 ( \53887 , \53885 , \53886 );
and \g130216/U$3 ( \53888 , \53879 , \53887 );
and \g130216/U$5 ( \53889 , \53844 , \53878 );
or \g130216/U$2 ( \53890 , \53888 , \53889 );
not \g131951/U$3 ( \53891 , \53612 );
not \g131951/U$4 ( \53892 , \53608 );
or \g131951/U$2 ( \53893 , \53891 , \53892 );
or \g131951/U$5 ( \53894 , \53608 , \53612 );
nand \g131951/U$1 ( \53895 , \53893 , \53894 );
not \g131601/U$3 ( \53896 , \47997 );
and \g131631/U$2 ( \53897 , \51604 , \48063 );
and \g131631/U$3 ( \53898 , \48064 , \51854 );
nor \g131631/U$1 ( \53899 , \53897 , \53898 );
not \g131601/U$4 ( \53900 , \53899 );
or \g131601/U$2 ( \53901 , \53896 , \53900 );
or \g131601/U$5 ( \53902 , \53899 , \47997 );
nand \g131601/U$1 ( \53903 , \53901 , \53902 );
xor \g456124/U$4 ( \53904 , \53895 , \53903 );
not \g131484/U$3 ( \53905 , \48159 );
and \g131512/U$2 ( \53906 , \51564 , \48155 );
and \g131512/U$3 ( \53907 , \48154 , \51098 );
nor \g131512/U$1 ( \53908 , \53906 , \53907 );
not \g131484/U$4 ( \53909 , \53908 );
or \g131484/U$2 ( \53910 , \53905 , \53909 );
or \g131484/U$5 ( \53911 , \53908 , \48159 );
nand \g131484/U$1 ( \53912 , \53910 , \53911 );
and \g456124/U$3 ( \53913 , \53904 , \53912 );
and \g456124/U$5 ( \53914 , \53895 , \53903 );
nor \g456124/U$2 ( \53915 , \53913 , \53914 );
not \g131525/U$3 ( \53916 , \53631 );
xor \g131884/U$1 ( \53917 , \53621 , \53613 );
not \g131525/U$4 ( \53918 , \53917 );
and \g131525/U$2 ( \53919 , \53916 , \53918 );
and \g131525/U$5 ( \53920 , \53631 , \53917 );
nor \g131525/U$1 ( \53921 , \53919 , \53920 );
or \g131009/U$2 ( \53922 , \53915 , \53921 );
not \g131014/U$3 ( \53923 , \53921 );
not \g131014/U$4 ( \53924 , \53915 );
or \g131014/U$2 ( \53925 , \53923 , \53924 );
not \g131238/U$3 ( \53926 , \48483 );
and \g131269/U$2 ( \53927 , \50752 , \48479 );
and \g131269/U$3 ( \53928 , \48478 , \50443 );
nor \g131269/U$1 ( \53929 , \53927 , \53928 );
not \g131238/U$4 ( \53930 , \53929 );
or \g131238/U$2 ( \53931 , \53926 , \53930 );
or \g131238/U$5 ( \53932 , \53929 , \48483 );
nand \g131238/U$1 ( \53933 , \53931 , \53932 );
not \g131357/U$3 ( \53934 , \48323 );
and \g131378/U$2 ( \53935 , \51117 , \48335 );
and \g131378/U$3 ( \53936 , \48334 , \50957 );
nor \g131378/U$1 ( \53937 , \53935 , \53936 );
not \g131357/U$4 ( \53938 , \53937 );
or \g131357/U$2 ( \53939 , \53934 , \53938 );
or \g131357/U$5 ( \53940 , \53937 , \48323 );
nand \g131357/U$1 ( \53941 , \53939 , \53940 );
xor \g131045/U$4 ( \53942 , \53933 , \53941 );
not \g131109/U$3 ( \53943 , \48685 );
and \g131143/U$2 ( \53944 , \50305 , \48860 );
and \g131143/U$3 ( \53945 , \48858 , \50019 );
nor \g131143/U$1 ( \53946 , \53944 , \53945 );
not \g131109/U$4 ( \53947 , \53946 );
or \g131109/U$2 ( \53948 , \53943 , \53947 );
or \g131109/U$5 ( \53949 , \53946 , \48685 );
nand \g131109/U$1 ( \53950 , \53948 , \53949 );
and \g131045/U$3 ( \53951 , \53942 , \53950 );
and \g131045/U$5 ( \53952 , \53933 , \53941 );
or \g131045/U$2 ( \53953 , \53951 , \53952 );
nand \g131014/U$1 ( \53954 , \53925 , \53953 );
nand \g131009/U$1 ( \53955 , \53922 , \53954 );
xor \g456024/U$5 ( \53956 , \53890 , \53955 );
xor \g129954/U$1 ( \53957 , \53366 , \53374 );
xor \g129954/U$1_r1 ( \53958 , \53957 , \53383 );
and \g456024/U$4 ( \53959 , \53956 , \53958 );
and \g456024/U$6 ( \53960 , \53890 , \53955 );
or \g456024/U$3 ( \53961 , \53959 , \53960 );
xor \g456035/U$1 ( \53962 , \53646 , \53648 );
xor \g456035/U$1_r1 ( \53963 , \53962 , \53651 );
xor \g456003/U$5 ( \53964 , \53961 , \53963 );
xor \g131200/U$1 ( \53965 , \53299 , \53310 );
xor \g131200/U$1_r1 ( \53966 , \53965 , \53319 );
not \g129738/U$3 ( \53967 , \53966 );
xor \g130138/U$1 ( \53968 , \53600 , \53634 );
xor \g130138/U$1_r1 ( \53969 , \53968 , \53643 );
not \g129738/U$4 ( \53970 , \53969 );
or \g129738/U$2 ( \53971 , \53967 , \53970 );
or \g129742/U$2 ( \53972 , \53969 , \53966 );
xor \g456033/U$1 ( \53973 , \53400 , \53408 );
xor \g456033/U$1_r1 ( \53974 , \53973 , \53417 );
nand \g129742/U$1 ( \53975 , \53972 , \53974 );
nand \g129738/U$1 ( \53976 , \53971 , \53975 );
and \g456003/U$4 ( \53977 , \53964 , \53976 );
and \g456003/U$6 ( \53978 , \53961 , \53963 );
or \g456003/U$3 ( \53979 , \53977 , \53978 );
not \g456004/U$1 ( \53980 , \53979 );
xor \g129279/U$4 ( \53981 , \53836 , \53980 );
xor \g455999/U$1 ( \53982 , \53587 , \53591 );
xor \g455999/U$1_r1 ( \53983 , \53982 , \53654 );
and \g129279/U$3 ( \53984 , \53981 , \53983 );
and \g129279/U$5 ( \53985 , \53836 , \53980 );
or \g129279/U$2 ( \53986 , \53984 , \53985 );
xor \g455989/U$4 ( \53987 , \53744 , \53986 );
xor \g455997/U$2 ( \53988 , \52969 , \53019 );
xor \g455997/U$1 ( \53989 , \53988 , \53046 );
xor \g455997/U$1_r1 ( \53990 , \53671 , \53676 );
xor \g455997/U$1_r2 ( \53991 , \53989 , \53990 );
and \g455989/U$3 ( \53992 , \53987 , \53991 );
and \g455989/U$5 ( \53993 , \53744 , \53986 );
nor \g455989/U$2 ( \53994 , \53992 , \53993 );
xor \g456007/U$1 ( \53995 , \53820 , \53822 );
xor \g456007/U$1_r1 ( \53996 , \53995 , \53833 );
not \g129486/U$1 ( \53997 , \53996 );
xor \g456024/U$2 ( \53998 , \53890 , \53955 );
xor \g456024/U$1 ( \53999 , \53998 , \53958 );
not \g130851/U$3 ( \54000 , \49233 );
and \g130875/U$2 ( \54001 , \49512 , \49405 );
and \g130875/U$3 ( \54002 , \49403 , \49282 );
nor \g130875/U$1 ( \54003 , \54001 , \54002 );
not \g130851/U$4 ( \54004 , \54003 );
or \g130851/U$2 ( \54005 , \54000 , \54004 );
or \g130851/U$5 ( \54006 , \54003 , \49233 );
nand \g130851/U$1 ( \54007 , \54005 , \54006 );
and \g131963/U$2 ( \54008 , \47914 , \52978 );
and \g131963/U$3 ( \54009 , \47913 , \52883 );
nor \g131963/U$1 ( \54010 , \54008 , \54009 );
and \g131928/U$2 ( \54011 , \54010 , \47977 );
not \g131928/U$4 ( \54012 , \54010 );
and \g131928/U$3 ( \54013 , \54012 , \47976 );
nor \g131928/U$1 ( \54014 , \54011 , \54013 );
xor \g132465/U$1 ( \54015 , \47450 , \47502 );
not \g135532/U$2 ( \54016 , \54015 );
nor \g135532/U$1 ( \54017 , \54016 , \40060 );
and \g132048/U$2 ( \54018 , \52978 , \47913 );
and \g132048/U$3 ( \54019 , \53300 , \47914 );
nor \g132048/U$1 ( \54020 , \54018 , \54019 );
and \g132009/U$2 ( \54021 , \54020 , \47977 );
not \g132009/U$4 ( \54022 , \54020 );
and \g132009/U$3 ( \54023 , \54022 , \47976 );
nor \g132009/U$1 ( \54024 , \54021 , \54023 );
and \g131947/U$2 ( \54025 , \54017 , \54024 );
xor \g131747/U$4 ( \54026 , \54014 , \54025 );
not \g131788/U$3 ( \54027 , \47935 );
and \g131820/U$2 ( \54028 , \52620 , \47931 );
and \g131820/U$3 ( \54029 , \47930 , \52352 );
nor \g131820/U$1 ( \54030 , \54028 , \54029 );
not \g131788/U$4 ( \54031 , \54030 );
or \g131788/U$2 ( \54032 , \54027 , \54031 );
or \g131788/U$5 ( \54033 , \54030 , \47935 );
nand \g131788/U$1 ( \54034 , \54032 , \54033 );
and \g131747/U$3 ( \54035 , \54026 , \54034 );
and \g131747/U$5 ( \54036 , \54014 , \54025 );
or \g131747/U$2 ( \54037 , \54035 , \54036 );
xor \g130288/U$4 ( \54038 , \54007 , \54037 );
not \g130344/U$3 ( \54039 , \50759 );
and \g130384/U$2 ( \54040 , \48349 , \51053 );
and \g130384/U$3 ( \54041 , \51055 , \48515 );
nor \g130384/U$1 ( \54042 , \54040 , \54041 );
not \g130344/U$4 ( \54043 , \54042 );
or \g130344/U$2 ( \54044 , \54039 , \54043 );
or \g130344/U$5 ( \54045 , \54042 , \50759 );
nand \g130344/U$1 ( \54046 , \54044 , \54045 );
and \g130288/U$3 ( \54047 , \54038 , \54046 );
and \g130288/U$5 ( \54048 , \54007 , \54037 );
or \g130288/U$2 ( \54049 , \54047 , \54048 );
not \g131661/U$3 ( \54050 , \47997 );
and \g131693/U$2 ( \54051 , \52108 , \48064 );
and \g131693/U$3 ( \54052 , \48063 , \51854 );
nor \g131693/U$1 ( \54053 , \54051 , \54052 );
not \g131661/U$4 ( \54054 , \54053 );
or \g131661/U$2 ( \54055 , \54050 , \54054 );
or \g131661/U$5 ( \54056 , \54053 , \47997 );
nand \g131661/U$1 ( \54057 , \54055 , \54056 );
xor \g132029/U$1 ( \54058 , \53850 , \53858 );
xor \g131496/U$4 ( \54059 , \54057 , \54058 );
not \g131550/U$3 ( \54060 , \48159 );
and \g131580/U$2 ( \54061 , \51604 , \48155 );
and \g131580/U$3 ( \54062 , \48154 , \51564 );
nor \g131580/U$1 ( \54063 , \54061 , \54062 );
not \g131550/U$4 ( \54064 , \54063 );
or \g131550/U$2 ( \54065 , \54060 , \54064 );
or \g131550/U$5 ( \54066 , \54063 , \48159 );
nand \g131550/U$1 ( \54067 , \54065 , \54066 );
and \g131496/U$3 ( \54068 , \54059 , \54067 );
and \g131496/U$5 ( \54069 , \54057 , \54058 );
or \g131496/U$2 ( \54070 , \54068 , \54069 );
xor \g131675/U$1 ( \54071 , \53859 , \53866 );
xor \g131675/U$1_r1 ( \54072 , \54071 , \53875 );
xor \g131033/U$4 ( \54073 , \54070 , \54072 );
and \g131323/U$2 ( \54074 , \50957 , \48479 );
and \g131323/U$3 ( \54075 , \48478 , \50752 );
nor \g131323/U$1 ( \54076 , \54074 , \54075 );
not \g131299/U$3 ( \54077 , \54076 );
not \g131299/U$4 ( \54078 , \48483 );
and \g131299/U$2 ( \54079 , \54077 , \54078 );
and \g131299/U$5 ( \54080 , \54076 , \48483 );
nor \g131299/U$1 ( \54081 , \54079 , \54080 );
and \g131446/U$2 ( \54082 , \51117 , \48334 );
and \g131446/U$3 ( \54083 , \48335 , \51098 );
nor \g131446/U$1 ( \54084 , \54082 , \54083 );
not \g131414/U$3 ( \54085 , \54084 );
not \g131414/U$4 ( \54086 , \48323 );
and \g131414/U$2 ( \54087 , \54085 , \54086 );
and \g131414/U$5 ( \54088 , \54084 , \48323 );
nor \g131414/U$1 ( \54089 , \54087 , \54088 );
or \g131156/U$2 ( \54090 , \54081 , \54089 );
and \g131171/U$2 ( \54091 , \54081 , \54089 );
and \g131215/U$2 ( \54092 , \50305 , \48858 );
and \g131215/U$3 ( \54093 , \48860 , \50443 );
nor \g131215/U$1 ( \54094 , \54092 , \54093 );
not \g131185/U$3 ( \54095 , \54094 );
not \g131185/U$4 ( \54096 , \48685 );
and \g131185/U$2 ( \54097 , \54095 , \54096 );
and \g131185/U$5 ( \54098 , \54094 , \48685 );
nor \g131185/U$1 ( \54099 , \54097 , \54098 );
nor \g131171/U$1 ( \54100 , \54091 , \54099 );
not \g131170/U$1 ( \54101 , \54100 );
nand \g131156/U$1 ( \54102 , \54090 , \54101 );
and \g131033/U$3 ( \54103 , \54073 , \54102 );
and \g131033/U$5 ( \54104 , \54070 , \54072 );
or \g131033/U$2 ( \54105 , \54103 , \54104 );
xor \g456029/U$5 ( \54106 , \54049 , \54105 );
xor \g130048/U$1 ( \54107 , \53485 , \53493 );
xor \g130048/U$1_r1 ( \54108 , \54107 , \53502 );
and \g456029/U$4 ( \54109 , \54106 , \54108 );
and \g456029/U$6 ( \54110 , \54049 , \54105 );
or \g456029/U$3 ( \54111 , \54109 , \54110 );
xor \g131252/U$1 ( \54112 , \53549 , \53550 );
xor \g131252/U$1_r1 ( \54113 , \54112 , \53559 );
not \g129829/U$3 ( \54114 , \54113 );
xor \g130216/U$1 ( \54115 , \53844 , \53878 );
xor \g130216/U$1_r1 ( \54116 , \54115 , \53887 );
not \g129829/U$4 ( \54117 , \54116 );
or \g129829/U$2 ( \54118 , \54114 , \54117 );
or \g129833/U$2 ( \54119 , \54116 , \54113 );
xor \g129869/U$1 ( \54120 , \53456 , \53464 );
xor \g129869/U$1_r1 ( \54121 , \54120 , \53473 );
nand \g129833/U$1 ( \54122 , \54119 , \54121 );
nand \g129829/U$1 ( \54123 , \54118 , \54122 );
xor \g456024/U$1_r1 ( \54124 , \54111 , \54123 );
xor \g456024/U$1_r2 ( \54125 , \53999 , \54124 );
not \g130795/U$3 ( \54126 , \49568 );
and \g130822/U$2 ( \54127 , \49282 , \49813 );
and \g130822/U$3 ( \54128 , \49812 , \49158 );
nor \g130822/U$1 ( \54129 , \54127 , \54128 );
not \g130795/U$4 ( \54130 , \54129 );
or \g130795/U$2 ( \54131 , \54126 , \54130 );
or \g130795/U$5 ( \54132 , \54129 , \49568 );
nand \g130795/U$1 ( \54133 , \54131 , \54132 );
not \g130905/U$3 ( \54134 , \49233 );
and \g130933/U$2 ( \54135 , \49512 , \49403 );
and \g130933/U$3 ( \54136 , \49405 , \49714 );
nor \g130933/U$1 ( \54137 , \54135 , \54136 );
not \g130905/U$4 ( \54138 , \54137 );
or \g130905/U$2 ( \54139 , \54134 , \54138 );
or \g130905/U$5 ( \54140 , \54137 , \49233 );
nand \g130905/U$1 ( \54141 , \54139 , \54140 );
xor \g130357/U$4 ( \54142 , \54133 , \54141 );
not \g130420/U$3 ( \54143 , \50759 );
and \g130449/U$2 ( \54144 , \48568 , \51055 );
and \g130449/U$3 ( \54145 , \51053 , \48515 );
nor \g130449/U$1 ( \54146 , \54144 , \54145 );
not \g130420/U$4 ( \54147 , \54146 );
or \g130420/U$2 ( \54148 , \54143 , \54147 );
or \g130420/U$5 ( \54149 , \54146 , \50759 );
nand \g130420/U$1 ( \54150 , \54148 , \54149 );
and \g130357/U$3 ( \54151 , \54142 , \54150 );
and \g130357/U$5 ( \54152 , \54133 , \54141 );
or \g130357/U$2 ( \54153 , \54151 , \54152 );
xor \g131045/U$1 ( \54154 , \53933 , \53941 );
xor \g131045/U$1_r1 ( \54155 , \54154 , \53950 );
xor \g456034/U$5 ( \54156 , \54153 , \54155 );
xor \g456053/U$1 ( \54157 , \53752 , \53760 );
xor \g456053/U$1_r1 ( \54158 , \54157 , \53769 );
and \g456034/U$4 ( \54159 , \54156 , \54158 );
and \g456034/U$6 ( \54160 , \54153 , \54155 );
or \g456034/U$3 ( \54161 , \54159 , \54160 );
xor \g456029/U$9 ( \54162 , \54049 , \54105 );
xor \g456029/U$9_r1 ( \54163 , \54162 , \54108 );
and \g456029/U$8 ( \54164 , \54161 , \54163 );
xor \g130288/U$1 ( \54165 , \54007 , \54037 );
xor \g130288/U$1_r1 ( \54166 , \54165 , \54046 );
xor \g131033/U$1 ( \54167 , \54070 , \54072 );
xor \g131033/U$1_r1 ( \54168 , \54167 , \54102 );
xor \g456028/U$5 ( \54169 , \54166 , \54168 );
xor \g129958/U$1 ( \54170 , \53790 , \53798 );
xor \g129958/U$1_r1 ( \54171 , \54170 , \53807 );
and \g456028/U$4 ( \54172 , \54169 , \54171 );
and \g456028/U$6 ( \54173 , \54166 , \54168 );
or \g456028/U$3 ( \54174 , \54172 , \54173 );
xor \g456029/U$11 ( \54175 , \54049 , \54105 );
xor \g456029/U$11_r1 ( \54176 , \54175 , \54108 );
and \g456029/U$10 ( \54177 , \54174 , \54176 );
and \g456029/U$12 ( \54178 , \54161 , \54174 );
or \g456029/U$7 ( \54179 , \54164 , \54177 , \54178 );
and \g129603/U$2 ( \54180 , \54125 , \54179 );
not \g129609/U$3 ( \54181 , \54125 );
not \g129609/U$4 ( \54182 , \54179 );
and \g129609/U$2 ( \54183 , \54181 , \54182 );
xor \g131947/U$1 ( \54184 , \54017 , \54024 );
xor \g132561/U$1 ( \54185 , \47447 , \47366 );
not \g135534/U$2 ( \54186 , \54185 );
nor \g135534/U$1 ( \54187 , \54186 , \40060 );
and \g132129/U$2 ( \54188 , \47914 , \53610 );
and \g132129/U$3 ( \54189 , \47913 , \53300 );
nor \g132129/U$1 ( \54190 , \54188 , \54189 );
and \g132089/U$2 ( \54191 , \54190 , \47977 );
not \g132089/U$4 ( \54192 , \54190 );
and \g132089/U$3 ( \54193 , \54192 , \47976 );
nor \g132089/U$1 ( \54194 , \54191 , \54193 );
and \g132031/U$2 ( \54195 , \54187 , \54194 );
xor \g131563/U$4 ( \54196 , \54184 , \54195 );
not \g131602/U$3 ( \54197 , \48159 );
and \g131632/U$2 ( \54198 , \51604 , \48154 );
and \g131632/U$3 ( \54199 , \48155 , \51854 );
nor \g131632/U$1 ( \54200 , \54198 , \54199 );
not \g131602/U$4 ( \54201 , \54200 );
or \g131602/U$2 ( \54202 , \54197 , \54201 );
or \g131602/U$5 ( \54203 , \54200 , \48159 );
nand \g131602/U$1 ( \54204 , \54202 , \54203 );
and \g131563/U$3 ( \54205 , \54196 , \54204 );
and \g131563/U$5 ( \54206 , \54184 , \54195 );
or \g131563/U$2 ( \54207 , \54205 , \54206 );
xor \g131747/U$1 ( \54208 , \54014 , \54025 );
xor \g131747/U$1_r1 ( \54209 , \54208 , \54034 );
xor \g130970/U$4 ( \54210 , \54207 , \54209 );
and \g131270/U$2 ( \54211 , \50752 , \48860 );
and \g131270/U$3 ( \54212 , \48858 , \50443 );
nor \g131270/U$1 ( \54213 , \54211 , \54212 );
not \g131239/U$3 ( \54214 , \54213 );
not \g131239/U$4 ( \54215 , \48685 );
and \g131239/U$2 ( \54216 , \54214 , \54215 );
and \g131239/U$5 ( \54217 , \54213 , \48685 );
nor \g131239/U$1 ( \54218 , \54216 , \54217 );
and \g131513/U$2 ( \54219 , \51564 , \48335 );
and \g131513/U$3 ( \54220 , \48334 , \51098 );
nor \g131513/U$1 ( \54221 , \54219 , \54220 );
not \g131485/U$3 ( \54222 , \54221 );
not \g131485/U$4 ( \54223 , \48323 );
and \g131485/U$2 ( \54224 , \54222 , \54223 );
and \g131485/U$5 ( \54225 , \54221 , \48323 );
nor \g131485/U$1 ( \54226 , \54224 , \54225 );
or \g131078/U$2 ( \54227 , \54218 , \54226 );
and \g131084/U$2 ( \54228 , \54218 , \54226 );
and \g131144/U$2 ( \54229 , \50305 , \49075 );
and \g131144/U$3 ( \54230 , \49074 , \50019 );
nor \g131144/U$1 ( \54231 , \54229 , \54230 );
not \g131110/U$3 ( \54232 , \54231 );
not \g131110/U$4 ( \54233 , \49014 );
and \g131110/U$2 ( \54234 , \54232 , \54233 );
and \g131110/U$5 ( \54235 , \54231 , \49014 );
nor \g131110/U$1 ( \54236 , \54234 , \54235 );
nor \g131084/U$1 ( \54237 , \54228 , \54236 );
not \g131083/U$1 ( \54238 , \54237 );
nand \g131078/U$1 ( \54239 , \54227 , \54238 );
and \g130970/U$3 ( \54240 , \54210 , \54239 );
and \g130970/U$5 ( \54241 , \54207 , \54209 );
or \g130970/U$2 ( \54242 , \54240 , \54241 );
not \g130740/U$3 ( \54243 , \49925 );
and \g130765/U$2 ( \54244 , \49102 , \50159 );
and \g130765/U$3 ( \54245 , \50160 , \49158 );
nor \g130765/U$1 ( \54246 , \54244 , \54245 );
not \g130740/U$4 ( \54247 , \54246 );
or \g130740/U$2 ( \54248 , \54243 , \54247 );
or \g130740/U$5 ( \54249 , \54246 , \49925 );
nand \g130740/U$1 ( \54250 , \54248 , \54249 );
xor \g132629/U$1 ( \54251 , \46260 , \47364 );
not \g135535/U$2 ( \54252 , \54251 );
nor \g135535/U$1 ( \54253 , \54252 , \40060 );
not \g132226/U$3 ( \54254 , \47948 );
and \g132279/U$2 ( \54255 , \47960 , \54185 );
and \g132279/U$3 ( \54256 , \54015 , \47959 );
nor \g132279/U$1 ( \54257 , \54255 , \54256 );
not \g132226/U$4 ( \54258 , \54257 );
or \g132226/U$2 ( \54259 , \54254 , \54258 );
or \g132226/U$5 ( \54260 , \54257 , \47948 );
nand \g132226/U$1 ( \54261 , \54259 , \54260 );
and \g132179/U$2 ( \54262 , \54253 , \54261 );
not \g132227/U$3 ( \54263 , \47948 );
and \g132280/U$2 ( \54264 , \47959 , \53848 );
and \g132280/U$3 ( \54265 , \54015 , \47960 );
nor \g132280/U$1 ( \54266 , \54264 , \54265 );
not \g132227/U$4 ( \54267 , \54266 );
or \g132227/U$2 ( \54268 , \54263 , \54267 );
or \g132227/U$5 ( \54269 , \54266 , \47948 );
nand \g132227/U$1 ( \54270 , \54268 , \54269 );
xor \g131738/U$4 ( \54271 , \54262 , \54270 );
not \g131789/U$3 ( \54272 , \47997 );
and \g131821/U$2 ( \54273 , \52620 , \48064 );
and \g131821/U$3 ( \54274 , \48063 , \52352 );
nor \g131821/U$1 ( \54275 , \54273 , \54274 );
not \g131789/U$4 ( \54276 , \54275 );
or \g131789/U$2 ( \54277 , \54272 , \54276 );
or \g131789/U$5 ( \54278 , \54275 , \47997 );
nand \g131789/U$1 ( \54279 , \54277 , \54278 );
and \g131738/U$3 ( \54280 , \54271 , \54279 );
and \g131738/U$5 ( \54281 , \54262 , \54270 );
or \g131738/U$2 ( \54282 , \54280 , \54281 );
xor \g456047/U$5 ( \54283 , \54250 , \54282 );
not \g130345/U$3 ( \54284 , \51124 );
and \g130386/U$2 ( \54285 , \48349 , \51517 );
and \g130386/U$3 ( \54286 , \51518 , \48515 );
nor \g130386/U$1 ( \54287 , \54285 , \54286 );
not \g130345/U$4 ( \54288 , \54287 );
or \g130345/U$2 ( \54289 , \54284 , \54288 );
or \g130345/U$5 ( \54290 , \54287 , \51124 );
nand \g130345/U$1 ( \54291 , \54289 , \54290 );
and \g456047/U$4 ( \54292 , \54283 , \54291 );
and \g456047/U$6 ( \54293 , \54250 , \54282 );
or \g456047/U$3 ( \54294 , \54292 , \54293 );
xor \g131496/U$1 ( \54295 , \54057 , \54058 );
xor \g131496/U$1_r1 ( \54296 , \54295 , \54067 );
xor \g130036/U$4 ( \54297 , \54294 , \54296 );
not \g130621/U$3 ( \54298 , \50362 );
and \g130655/U$2 ( \54299 , \48833 , \50587 );
and \g130655/U$3 ( \54300 , \50588 , \48977 );
nor \g130655/U$1 ( \54301 , \54299 , \54300 );
not \g130621/U$4 ( \54302 , \54301 );
or \g130621/U$2 ( \54303 , \54298 , \54302 );
or \g130621/U$5 ( \54304 , \54301 , \50362 );
nand \g130621/U$1 ( \54305 , \54303 , \54304 );
not \g131358/U$3 ( \54306 , \48483 );
and \g131379/U$2 ( \54307 , \51117 , \48479 );
and \g131379/U$3 ( \54308 , \48478 , \50957 );
nor \g131379/U$1 ( \54309 , \54307 , \54308 );
not \g131358/U$4 ( \54310 , \54309 );
or \g131358/U$2 ( \54311 , \54306 , \54310 );
or \g131358/U$5 ( \54312 , \54309 , \48483 );
nand \g131358/U$1 ( \54313 , \54311 , \54312 );
xor \g130139/U$4 ( \54314 , \54305 , \54313 );
not \g130206/U$3 ( \54315 , \51120 );
and \g130243/U$2 ( \54316 , \48353 , \52273 );
and \g130243/U$3 ( \54317 , \52270 , \48138 );
nor \g130243/U$1 ( \54318 , \54316 , \54317 );
not \g130206/U$4 ( \54319 , \54318 );
or \g130206/U$2 ( \54320 , \54315 , \54319 );
or \g130206/U$5 ( \54321 , \54318 , \51120 );
nand \g130206/U$1 ( \54322 , \54320 , \54321 );
and \g130139/U$3 ( \54323 , \54314 , \54322 );
and \g130139/U$5 ( \54324 , \54305 , \54313 );
or \g130139/U$2 ( \54325 , \54323 , \54324 );
and \g130036/U$3 ( \54326 , \54297 , \54325 );
and \g130036/U$5 ( \54327 , \54294 , \54296 );
or \g130036/U$2 ( \54328 , \54326 , \54327 );
xor \g456043/U$4 ( \54329 , \54242 , \54328 );
xor \g456124/U$1 ( \54330 , \53895 , \53903 );
xor \g456124/U$1_r1 ( \54331 , \54330 , \53912 );
not \g130684/U$3 ( \54332 , \49925 );
and \g130710/U$2 ( \54333 , \49102 , \50160 );
and \g130710/U$3 ( \54334 , \50159 , \48977 );
nor \g130710/U$1 ( \54335 , \54333 , \54334 );
not \g130684/U$4 ( \54336 , \54335 );
or \g130684/U$2 ( \54337 , \54332 , \54336 );
or \g130684/U$5 ( \54338 , \54335 , \49925 );
nand \g130684/U$1 ( \54339 , \54337 , \54338 );
and \g132201/U$2 ( \54340 , \47959 , \53610 );
and \g132201/U$3 ( \54341 , \53848 , \47960 );
nor \g132201/U$1 ( \54342 , \54340 , \54341 );
not \g132155/U$3 ( \54343 , \54342 );
not \g132155/U$4 ( \54344 , \47948 );
and \g132155/U$2 ( \54345 , \54343 , \54344 );
and \g132155/U$5 ( \54346 , \54342 , \47948 );
nor \g132155/U$1 ( \54347 , \54345 , \54346 );
and \g131894/U$2 ( \54348 , \52620 , \47930 );
and \g131894/U$3 ( \54349 , \47931 , \52883 );
nor \g131894/U$1 ( \54350 , \54348 , \54349 );
not \g131856/U$3 ( \54351 , \54350 );
not \g131856/U$4 ( \54352 , \47935 );
and \g131856/U$2 ( \54353 , \54351 , \54352 );
and \g131856/U$5 ( \54354 , \54350 , \47935 );
nor \g131856/U$1 ( \54355 , \54353 , \54354 );
or \g131703/U$2 ( \54356 , \54347 , \54355 );
and \g131710/U$2 ( \54357 , \54347 , \54355 );
and \g131761/U$2 ( \54358 , \52108 , \48063 );
and \g131761/U$3 ( \54359 , \48064 , \52352 );
nor \g131761/U$1 ( \54360 , \54358 , \54359 );
not \g131730/U$3 ( \54361 , \54360 );
not \g131730/U$4 ( \54362 , \47997 );
and \g131730/U$2 ( \54363 , \54361 , \54362 );
and \g131730/U$5 ( \54364 , \54360 , \47997 );
nor \g131730/U$1 ( \54365 , \54363 , \54364 );
nor \g131710/U$1 ( \54366 , \54357 , \54365 );
not \g131709/U$1 ( \54367 , \54366 );
nand \g131703/U$1 ( \54368 , \54356 , \54367 );
xor \g130050/U$4 ( \54369 , \54339 , \54368 );
not \g130125/U$3 ( \54370 , \51120 );
and \g130163/U$2 ( \54371 , \48117 , \52270 );
and \g130163/U$3 ( \54372 , \52273 , \48138 );
nor \g130163/U$1 ( \54373 , \54371 , \54372 );
not \g130125/U$4 ( \54374 , \54373 );
or \g130125/U$2 ( \54375 , \54370 , \54374 );
or \g130125/U$5 ( \54376 , \54373 , \51120 );
nand \g130125/U$1 ( \54377 , \54375 , \54376 );
and \g130050/U$3 ( \54378 , \54369 , \54377 );
and \g130050/U$5 ( \54379 , \54339 , \54368 );
or \g130050/U$2 ( \54380 , \54378 , \54379 );
xor \g456044/U$1 ( \54381 , \54331 , \54380 );
not \g130558/U$3 ( \54382 , \50362 );
and \g130587/U$2 ( \54383 , \48726 , \50587 );
and \g130587/U$3 ( \54384 , \50588 , \48833 );
nor \g130587/U$1 ( \54385 , \54383 , \54384 );
not \g130558/U$4 ( \54386 , \54385 );
or \g130558/U$2 ( \54387 , \54382 , \54386 );
or \g130558/U$5 ( \54388 , \54385 , \50362 );
nand \g130558/U$1 ( \54389 , \54387 , \54388 );
not \g131027/U$3 ( \54390 , \49014 );
and \g131068/U$2 ( \54391 , \49888 , \49074 );
and \g131068/U$3 ( \54392 , \49075 , \50019 );
nor \g131068/U$1 ( \54393 , \54391 , \54392 );
not \g131027/U$4 ( \54394 , \54393 );
or \g131027/U$2 ( \54395 , \54390 , \54394 );
or \g131027/U$5 ( \54396 , \54393 , \49014 );
nand \g131027/U$1 ( \54397 , \54395 , \54396 );
xor \g130219/U$4 ( \54398 , \54389 , \54397 );
not \g130278/U$3 ( \54399 , \51124 );
and \g130312/U$2 ( \54400 , \48349 , \51518 );
and \g130312/U$3 ( \54401 , \51517 , \48353 );
nor \g130312/U$1 ( \54402 , \54400 , \54401 );
not \g130278/U$4 ( \54403 , \54402 );
or \g130278/U$2 ( \54404 , \54399 , \54403 );
or \g130278/U$5 ( \54405 , \54402 , \51124 );
nand \g130278/U$1 ( \54406 , \54404 , \54405 );
and \g130219/U$3 ( \54407 , \54398 , \54406 );
and \g130219/U$5 ( \54408 , \54389 , \54397 );
or \g130219/U$2 ( \54409 , \54407 , \54408 );
xor \g456044/U$1_r1 ( \54410 , \54381 , \54409 );
and \g456043/U$3 ( \54411 , \54329 , \54410 );
and \g456043/U$5 ( \54412 , \54242 , \54328 );
nor \g456043/U$2 ( \54413 , \54411 , \54412 );
xor \g456044/U$4 ( \54414 , \54331 , \54380 );
and \g456044/U$3 ( \54415 , \54414 , \54409 );
and \g456044/U$5 ( \54416 , \54331 , \54380 );
nor \g456044/U$2 ( \54417 , \54415 , \54416 );
not \g131011/U$3 ( \54418 , \53953 );
xnor \g131397/U$1 ( \54419 , \53921 , \53915 );
not \g131011/U$4 ( \54420 , \54419 );
and \g131011/U$2 ( \54421 , \54418 , \54420 );
and \g131011/U$5 ( \54422 , \53953 , \54419 );
nor \g131011/U$1 ( \54423 , \54421 , \54422 );
xor \g456021/U$9 ( \54424 , \54417 , \54423 );
not \g129919/U$3 ( \54425 , \53810 );
xnor \g130108/U$1 ( \54426 , \53778 , \53772 );
not \g129919/U$4 ( \54427 , \54426 );
and \g129919/U$2 ( \54428 , \54425 , \54427 );
and \g129919/U$5 ( \54429 , \53810 , \54426 );
nor \g129919/U$1 ( \54430 , \54428 , \54429 );
xor \g456021/U$9_r1 ( \54431 , \54424 , \54430 );
and \g456021/U$8 ( \54432 , \54413 , \54431 );
xnor \g455949/U$1 ( \54433 , \54121 , \54116 );
not \g129784/U$3 ( \54434 , \54433 );
not \g129784/U$4 ( \54435 , \54113 );
and \g129784/U$2 ( \54436 , \54434 , \54435 );
and \g129784/U$5 ( \54437 , \54433 , \54113 );
nor \g129784/U$1 ( \54438 , \54436 , \54437 );
xor \g456021/U$11 ( \54439 , \54417 , \54423 );
xor \g456021/U$11_r1 ( \54440 , \54439 , \54430 );
and \g456021/U$10 ( \54441 , \54438 , \54440 );
and \g456021/U$12 ( \54442 , \54413 , \54438 );
or \g456021/U$7 ( \54443 , \54432 , \54441 , \54442 );
nor \g129609/U$1 ( \54444 , \54183 , \54443 );
nor \g129603/U$1 ( \54445 , \54180 , \54444 );
or \g129412/U$2 ( \54446 , \53997 , \54445 );
not \g129432/U$3 ( \54447 , \54445 );
not \g129432/U$4 ( \54448 , \53997 );
or \g129432/U$2 ( \54449 , \54447 , \54448 );
xor \g456003/U$2 ( \54450 , \53961 , \53963 );
xor \g456003/U$1 ( \54451 , \54450 , \53976 );
xor \g456024/U$9 ( \54452 , \53890 , \53955 );
xor \g456024/U$9_r1 ( \54453 , \54452 , \53958 );
and \g456024/U$8 ( \54454 , \54111 , \54453 );
xor \g456024/U$11 ( \54455 , \53890 , \53955 );
xor \g456024/U$11_r1 ( \54456 , \54455 , \53958 );
and \g456024/U$10 ( \54457 , \54123 , \54456 );
and \g456024/U$12 ( \54458 , \54111 , \54123 );
or \g456024/U$7 ( \54459 , \54454 , \54457 , \54458 );
xnor \g455948/U$1 ( \54460 , \53974 , \53969 );
not \g129701/U$3 ( \54461 , \54460 );
not \g129701/U$4 ( \54462 , \53966 );
and \g129701/U$2 ( \54463 , \54461 , \54462 );
and \g129701/U$5 ( \54464 , \54460 , \53966 );
nor \g129701/U$1 ( \54465 , \54463 , \54464 );
xor \g456021/U$5 ( \54466 , \54417 , \54423 );
and \g456021/U$4 ( \54467 , \54466 , \54430 );
and \g456021/U$6 ( \54468 , \54417 , \54423 );
or \g456021/U$3 ( \54469 , \54467 , \54468 );
or \g129604/U$2 ( \54470 , \54465 , \54469 );
not \g129610/U$3 ( \54471 , \54469 );
not \g129610/U$4 ( \54472 , \54465 );
or \g129610/U$2 ( \54473 , \54471 , \54472 );
xor \g129695/U$1 ( \54474 , \53812 , \53814 );
xor \g129695/U$1_r1 ( \54475 , \54474 , \53817 );
nand \g129610/U$1 ( \54476 , \54473 , \54475 );
nand \g129604/U$1 ( \54477 , \54470 , \54476 );
xor \g456003/U$1_r1 ( \54478 , \54459 , \54477 );
xor \g456003/U$1_r2 ( \54479 , \54451 , \54478 );
nand \g129432/U$1 ( \54480 , \54449 , \54479 );
nand \g129412/U$1 ( \54481 , \54446 , \54480 );
and \g131634/U$2 ( \54482 , \51604 , \48478 );
and \g131634/U$3 ( \54483 , \48479 , \51854 );
nor \g131634/U$1 ( \54484 , \54482 , \54483 );
not \g131605/U$3 ( \54485 , \54484 );
not \g131605/U$4 ( \54486 , \48483 );
and \g131605/U$2 ( \54487 , \54485 , \54486 );
and \g131605/U$5 ( \54488 , \54484 , \48483 );
nor \g131605/U$1 ( \54489 , \54487 , \54488 );
and \g131763/U$2 ( \54490 , \52108 , \48334 );
and \g131763/U$3 ( \54491 , \48335 , \52352 );
nor \g131763/U$1 ( \54492 , \54490 , \54491 );
not \g131732/U$3 ( \54493 , \54492 );
not \g131732/U$4 ( \54494 , \48323 );
and \g131732/U$2 ( \54495 , \54493 , \54494 );
and \g131732/U$5 ( \54496 , \54492 , \48323 );
nor \g131732/U$1 ( \54497 , \54495 , \54496 );
or \g131455/U$2 ( \54498 , \54489 , \54497 );
and \g131463/U$2 ( \54499 , \54489 , \54497 );
and \g131515/U$2 ( \54500 , \51564 , \48860 );
and \g131515/U$3 ( \54501 , \48858 , \51098 );
nor \g131515/U$1 ( \54502 , \54500 , \54501 );
not \g131487/U$3 ( \54503 , \54502 );
not \g131487/U$4 ( \54504 , \48685 );
and \g131487/U$2 ( \54505 , \54503 , \54504 );
and \g131487/U$5 ( \54506 , \54502 , \48685 );
nor \g131487/U$1 ( \54507 , \54505 , \54506 );
nor \g131463/U$1 ( \54508 , \54499 , \54507 );
not \g131462/U$1 ( \54509 , \54508 );
nand \g131455/U$1 ( \54510 , \54498 , \54509 );
and \g132304/U$2 ( \54511 , \47913 , \53848 );
and \g132304/U$3 ( \54512 , \54015 , \47914 );
nor \g132304/U$1 ( \54513 , \54511 , \54512 );
and \g132255/U$2 ( \54514 , \54513 , \47977 );
not \g132255/U$4 ( \54515 , \54513 );
and \g132255/U$3 ( \54516 , \54515 , \47976 );
nor \g132255/U$1 ( \54517 , \54514 , \54516 );
not \g132090/U$3 ( \54518 , \47935 );
and \g132130/U$2 ( \54519 , \47931 , \53610 );
and \g132130/U$3 ( \54520 , \47930 , \53300 );
nor \g132130/U$1 ( \54521 , \54519 , \54520 );
not \g132090/U$4 ( \54522 , \54521 );
or \g132090/U$2 ( \54523 , \54518 , \54522 );
or \g132090/U$5 ( \54524 , \54521 , \47935 );
nand \g132090/U$1 ( \54525 , \54523 , \54524 );
xor \g132019/U$1 ( \54526 , \54517 , \54525 );
not \g132229/U$3 ( \54527 , \47948 );
and \g132282/U$2 ( \54528 , \47959 , \54251 );
xor \g132696/U$1 ( \54529 , \47350 , \47361 );
and \g132282/U$3 ( \54530 , \54529 , \47960 );
nor \g132282/U$1 ( \54531 , \54528 , \54530 );
not \g132229/U$4 ( \54532 , \54531 );
or \g132229/U$2 ( \54533 , \54527 , \54532 );
or \g132229/U$5 ( \54534 , \54531 , \47948 );
nand \g132229/U$1 ( \54535 , \54533 , \54534 );
not \g132189/U$2 ( \54536 , \54535 );
xor \g132772/U$1 ( \54537 , \47347 , \47320 );
nand \g132380/U$1 ( \54538 , \54537 , \40061 );
nor \g132189/U$1 ( \54539 , \54536 , \54538 );
xor \g132019/U$1_r1 ( \54540 , \54526 , \54539 );
xor \g130632/U$4 ( \54541 , \54510 , \54540 );
not \g130686/U$3 ( \54542 , \50759 );
and \g130712/U$2 ( \54543 , \49102 , \51055 );
and \g130712/U$3 ( \54544 , \51053 , \48977 );
nor \g130712/U$1 ( \54545 , \54543 , \54544 );
not \g130686/U$4 ( \54546 , \54545 );
or \g130686/U$2 ( \54547 , \54542 , \54546 );
or \g130686/U$5 ( \54548 , \54545 , \50759 );
nand \g130686/U$1 ( \54549 , \54547 , \54548 );
and \g130632/U$3 ( \54550 , \54541 , \54549 );
and \g130632/U$5 ( \54551 , \54510 , \54540 );
or \g130632/U$2 ( \54552 , \54550 , \54551 );
not \g130741/U$3 ( \54553 , \50362 );
and \g130766/U$2 ( \54554 , \49102 , \50587 );
and \g130766/U$3 ( \54555 , \50588 , \49158 );
nor \g130766/U$1 ( \54556 , \54554 , \54555 );
not \g130741/U$4 ( \54557 , \54556 );
or \g130741/U$2 ( \54558 , \54553 , \54557 );
or \g130741/U$5 ( \54559 , \54556 , \50362 );
nand \g130741/U$1 ( \54560 , \54558 , \54559 );
xor \g132179/U$1 ( \54561 , \54253 , \54261 );
not \g131857/U$3 ( \54562 , \47997 );
and \g131895/U$2 ( \54563 , \52620 , \48063 );
and \g131895/U$3 ( \54564 , \48064 , \52883 );
nor \g131895/U$1 ( \54565 , \54563 , \54564 );
not \g131857/U$4 ( \54566 , \54565 );
or \g131857/U$2 ( \54567 , \54562 , \54566 );
or \g131857/U$5 ( \54568 , \54565 , \47997 );
nand \g131857/U$1 ( \54569 , \54567 , \54568 );
xor \g131676/U$1 ( \54570 , \54561 , \54569 );
not \g131731/U$3 ( \54571 , \48159 );
and \g131762/U$2 ( \54572 , \52108 , \48154 );
and \g131762/U$3 ( \54573 , \48155 , \52352 );
nor \g131762/U$1 ( \54574 , \54572 , \54573 );
not \g131731/U$4 ( \54575 , \54574 );
or \g131731/U$2 ( \54576 , \54571 , \54575 );
or \g131731/U$5 ( \54577 , \54574 , \48159 );
nand \g131731/U$1 ( \54578 , \54576 , \54577 );
xor \g131676/U$1_r1 ( \54579 , \54570 , \54578 );
xor \g130567/U$1 ( \54580 , \54560 , \54579 );
not \g130622/U$3 ( \54581 , \50759 );
and \g130656/U$2 ( \54582 , \48833 , \51053 );
and \g130656/U$3 ( \54583 , \51055 , \48977 );
nor \g130656/U$1 ( \54584 , \54582 , \54583 );
not \g130622/U$4 ( \54585 , \54584 );
or \g130622/U$2 ( \54586 , \54581 , \54585 );
or \g130622/U$5 ( \54587 , \54584 , \50759 );
nand \g130622/U$1 ( \54588 , \54586 , \54587 );
xor \g130567/U$1_r1 ( \54589 , \54580 , \54588 );
xor \g456059/U$4 ( \54590 , \54552 , \54589 );
not \g130964/U$3 ( \54591 , \49568 );
and \g130991/U$2 ( \54592 , \49888 , \49813 );
and \g130991/U$3 ( \54593 , \49812 , \49714 );
nor \g130991/U$1 ( \54594 , \54592 , \54593 );
not \g130964/U$4 ( \54595 , \54594 );
or \g130964/U$2 ( \54596 , \54591 , \54595 );
or \g130964/U$5 ( \54597 , \54594 , \49568 );
nand \g130964/U$1 ( \54598 , \54596 , \54597 );
and \g132202/U$2 ( \54599 , \47913 , \53610 );
and \g132202/U$3 ( \54600 , \53848 , \47914 );
nor \g132202/U$1 ( \54601 , \54599 , \54600 );
and \g132157/U$2 ( \54602 , \54601 , \47977 );
not \g132157/U$4 ( \54603 , \54601 );
and \g132157/U$3 ( \54604 , \54603 , \47976 );
nor \g132157/U$1 ( \54605 , \54602 , \54604 );
not \g132011/U$3 ( \54606 , \47935 );
and \g132049/U$2 ( \54607 , \52978 , \47930 );
and \g132049/U$3 ( \54608 , \47931 , \53300 );
nor \g132049/U$1 ( \54609 , \54607 , \54608 );
not \g132011/U$4 ( \54610 , \54609 );
or \g132011/U$2 ( \54611 , \54606 , \54610 );
or \g132011/U$5 ( \54612 , \54609 , \47935 );
nand \g132011/U$1 ( \54613 , \54611 , \54612 );
xor \g131936/U$1 ( \54614 , \54605 , \54613 );
not \g135537/U$2 ( \54615 , \54529 );
nor \g135537/U$1 ( \54616 , \54615 , \40060 );
not \g132228/U$3 ( \54617 , \47948 );
and \g132281/U$2 ( \54618 , \47959 , \54185 );
and \g132281/U$3 ( \54619 , \54251 , \47960 );
nor \g132281/U$1 ( \54620 , \54618 , \54619 );
not \g132228/U$4 ( \54621 , \54620 );
or \g132228/U$2 ( \54622 , \54617 , \54621 );
or \g132228/U$5 ( \54623 , \54620 , \47948 );
nand \g132228/U$1 ( \54624 , \54622 , \54623 );
and \g132170/U$2 ( \54625 , \54616 , \54624 );
xor \g131936/U$1_r1 ( \54626 , \54614 , \54625 );
xor \g130290/U$1 ( \54627 , \54598 , \54626 );
not \g130346/U$3 ( \54628 , \51120 );
and \g130387/U$2 ( \54629 , \48349 , \52270 );
and \g130387/U$3 ( \54630 , \52273 , \48515 );
nor \g130387/U$1 ( \54631 , \54629 , \54630 );
not \g130346/U$4 ( \54632 , \54631 );
or \g130346/U$2 ( \54633 , \54628 , \54632 );
or \g130346/U$5 ( \54634 , \54631 , \51120 );
nand \g130346/U$1 ( \54635 , \54633 , \54634 );
xor \g130290/U$1_r1 ( \54636 , \54627 , \54635 );
and \g456059/U$3 ( \54637 , \54590 , \54636 );
and \g456059/U$5 ( \54638 , \54552 , \54589 );
nor \g456059/U$2 ( \54639 , \54637 , \54638 );
xor \g132031/U$1 ( \54640 , \54187 , \54194 );
not \g131929/U$3 ( \54641 , \47935 );
and \g131964/U$2 ( \54642 , \52978 , \47931 );
and \g131964/U$3 ( \54643 , \47930 , \52883 );
nor \g131964/U$1 ( \54644 , \54642 , \54643 );
not \g131929/U$4 ( \54645 , \54644 );
or \g131929/U$2 ( \54646 , \54641 , \54645 );
or \g131929/U$5 ( \54647 , \54644 , \47935 );
nand \g131929/U$1 ( \54648 , \54646 , \54647 );
xor \g456137/U$1 ( \54649 , \54640 , \54648 );
not \g131662/U$3 ( \54650 , \48159 );
and \g131694/U$2 ( \54651 , \52108 , \48155 );
and \g131694/U$3 ( \54652 , \48154 , \51854 );
nor \g131694/U$1 ( \54653 , \54651 , \54652 );
not \g131662/U$4 ( \54654 , \54653 );
or \g131662/U$2 ( \54655 , \54650 , \54654 );
or \g131662/U$5 ( \54656 , \54653 , \48159 );
nand \g131662/U$1 ( \54657 , \54655 , \54656 );
xor \g456137/U$1_r1 ( \54658 , \54649 , \54657 );
and \g130877/U$2 ( \54659 , \49512 , \50160 );
and \g130877/U$3 ( \54660 , \50159 , \49282 );
nor \g130877/U$1 ( \54661 , \54659 , \54660 );
not \g130853/U$3 ( \54662 , \54661 );
not \g130853/U$4 ( \54663 , \49925 );
and \g130853/U$2 ( \54664 , \54662 , \54663 );
and \g130853/U$5 ( \54665 , \54661 , \49925 );
nor \g130853/U$1 ( \54666 , \54664 , \54665 );
not \g131791/U$3 ( \54667 , \48159 );
and \g131822/U$2 ( \54668 , \52620 , \48155 );
and \g131822/U$3 ( \54669 , \48154 , \52352 );
nor \g131822/U$1 ( \54670 , \54668 , \54669 );
not \g131791/U$4 ( \54671 , \54670 );
or \g131791/U$2 ( \54672 , \54667 , \54671 );
or \g131791/U$5 ( \54673 , \54670 , \48159 );
nand \g131791/U$1 ( \54674 , \54672 , \54673 );
not \g131930/U$3 ( \54675 , \47997 );
and \g131965/U$2 ( \54676 , \52978 , \48064 );
and \g131965/U$3 ( \54677 , \48063 , \52883 );
nor \g131965/U$1 ( \54678 , \54676 , \54677 );
not \g131930/U$4 ( \54679 , \54678 );
or \g131930/U$2 ( \54680 , \54675 , \54679 );
or \g131930/U$5 ( \54681 , \54678 , \47997 );
nand \g131930/U$1 ( \54682 , \54680 , \54681 );
xor \g456143/U$4 ( \54683 , \54674 , \54682 );
xor \g132170/U$1 ( \54684 , \54616 , \54624 );
and \g456143/U$3 ( \54685 , \54683 , \54684 );
and \g456143/U$5 ( \54686 , \54674 , \54682 );
nor \g456143/U$2 ( \54687 , \54685 , \54686 );
or \g130456/U$2 ( \54688 , \54666 , \54687 );
and \g130468/U$2 ( \54689 , \54666 , \54687 );
and \g130523/U$2 ( \54690 , \48726 , \51518 );
and \g130523/U$3 ( \54691 , \51517 , \48568 );
nor \g130523/U$1 ( \54692 , \54690 , \54691 );
not \g130492/U$3 ( \54693 , \54692 );
not \g130492/U$4 ( \54694 , \51124 );
and \g130492/U$2 ( \54695 , \54693 , \54694 );
and \g130492/U$5 ( \54696 , \54692 , \51124 );
nor \g130492/U$1 ( \54697 , \54695 , \54696 );
nor \g130468/U$1 ( \54698 , \54689 , \54697 );
not \g130467/U$1 ( \54699 , \54698 );
nand \g130456/U$1 ( \54700 , \54688 , \54699 );
xor \g456063/U$1 ( \54701 , \54658 , \54700 );
not \g131240/U$3 ( \54702 , \49014 );
and \g131272/U$2 ( \54703 , \50752 , \49075 );
and \g131272/U$3 ( \54704 , \49074 , \50443 );
nor \g131272/U$1 ( \54705 , \54703 , \54704 );
not \g131240/U$4 ( \54706 , \54705 );
or \g131240/U$2 ( \54707 , \54702 , \54706 );
or \g131240/U$5 ( \54708 , \54705 , \49014 );
nand \g131240/U$1 ( \54709 , \54707 , \54708 );
xor \g132019/U$4 ( \54710 , \54517 , \54525 );
and \g132019/U$3 ( \54711 , \54710 , \54539 );
and \g132019/U$5 ( \54712 , \54517 , \54525 );
or \g132019/U$2 ( \54713 , \54711 , \54712 );
xor \g131048/U$4 ( \54714 , \54709 , \54713 );
not \g131111/U$3 ( \54715 , \49233 );
and \g131145/U$2 ( \54716 , \50305 , \49405 );
and \g131145/U$3 ( \54717 , \49403 , \50019 );
nor \g131145/U$1 ( \54718 , \54716 , \54717 );
not \g131111/U$4 ( \54719 , \54718 );
or \g131111/U$2 ( \54720 , \54715 , \54719 );
or \g131111/U$5 ( \54721 , \54718 , \49233 );
nand \g131111/U$1 ( \54722 , \54720 , \54721 );
and \g131048/U$3 ( \54723 , \54714 , \54722 );
and \g131048/U$5 ( \54724 , \54709 , \54713 );
or \g131048/U$2 ( \54725 , \54723 , \54724 );
xor \g456063/U$1_r1 ( \54726 , \54701 , \54725 );
not \g130348/U$1 ( \54727 , \54726 );
or \g130167/U$2 ( \54728 , \54639 , \54727 );
not \g130179/U$3 ( \54729 , \54727 );
not \g130179/U$4 ( \54730 , \54639 );
or \g130179/U$2 ( \54731 , \54729 , \54730 );
not \g131551/U$3 ( \54732 , \48323 );
and \g131581/U$2 ( \54733 , \51604 , \48335 );
and \g131581/U$3 ( \54734 , \48334 , \51564 );
nor \g131581/U$1 ( \54735 , \54733 , \54734 );
not \g131551/U$4 ( \54736 , \54735 );
or \g131551/U$2 ( \54737 , \54732 , \54736 );
or \g131551/U$5 ( \54738 , \54735 , \48323 );
nand \g131551/U$1 ( \54739 , \54737 , \54738 );
not \g131300/U$3 ( \54740 , \48685 );
and \g131324/U$2 ( \54741 , \50957 , \48860 );
and \g131324/U$3 ( \54742 , \48858 , \50752 );
nor \g131324/U$1 ( \54743 , \54741 , \54742 );
not \g131300/U$4 ( \54744 , \54743 );
or \g131300/U$2 ( \54745 , \54740 , \54744 );
or \g131300/U$5 ( \54746 , \54743 , \48685 );
nand \g131300/U$1 ( \54747 , \54745 , \54746 );
xor \g456105/U$1 ( \54748 , \54739 , \54747 );
not \g131186/U$3 ( \54749 , \49014 );
and \g131216/U$2 ( \54750 , \50305 , \49074 );
and \g131216/U$3 ( \54751 , \49075 , \50443 );
nor \g131216/U$1 ( \54752 , \54750 , \54751 );
not \g131186/U$4 ( \54753 , \54752 );
or \g131186/U$2 ( \54754 , \54749 , \54753 );
or \g131186/U$5 ( \54755 , \54752 , \49014 );
nand \g131186/U$1 ( \54756 , \54754 , \54755 );
xor \g456105/U$1_r1 ( \54757 , \54748 , \54756 );
xor \g130290/U$4 ( \54758 , \54598 , \54626 );
and \g130290/U$3 ( \54759 , \54758 , \54635 );
and \g130290/U$5 ( \54760 , \54598 , \54626 );
or \g130290/U$2 ( \54761 , \54759 , \54760 );
xor \g456055/U$1 ( \54762 , \54757 , \54761 );
xor \g130567/U$4 ( \54763 , \54560 , \54579 );
and \g130567/U$3 ( \54764 , \54763 , \54588 );
and \g130567/U$5 ( \54765 , \54560 , \54579 );
or \g130567/U$2 ( \54766 , \54764 , \54765 );
xor \g456055/U$1_r1 ( \54767 , \54762 , \54766 );
nand \g130179/U$1 ( \54768 , \54731 , \54767 );
nand \g130167/U$1 ( \54769 , \54728 , \54768 );
not \g131486/U$3 ( \54770 , \48483 );
and \g131514/U$2 ( \54771 , \51564 , \48479 );
and \g131514/U$3 ( \54772 , \48478 , \51098 );
nor \g131514/U$1 ( \54773 , \54771 , \54772 );
not \g131486/U$4 ( \54774 , \54773 );
or \g131486/U$2 ( \54775 , \54770 , \54774 );
or \g131486/U$5 ( \54776 , \54773 , \48483 );
nand \g131486/U$1 ( \54777 , \54775 , \54776 );
not \g131603/U$3 ( \54778 , \48323 );
and \g131633/U$2 ( \54779 , \51604 , \48334 );
and \g131633/U$3 ( \54780 , \48335 , \51854 );
nor \g131633/U$1 ( \54781 , \54779 , \54780 );
not \g131603/U$4 ( \54782 , \54781 );
or \g131603/U$2 ( \54783 , \54778 , \54782 );
or \g131603/U$5 ( \54784 , \54781 , \48323 );
nand \g131603/U$1 ( \54785 , \54783 , \54784 );
xor \g131312/U$1 ( \54786 , \54777 , \54785 );
not \g131359/U$3 ( \54787 , \48685 );
and \g131380/U$2 ( \54788 , \51117 , \48860 );
and \g131380/U$3 ( \54789 , \48858 , \50957 );
nor \g131380/U$1 ( \54790 , \54788 , \54789 );
not \g131359/U$4 ( \54791 , \54790 );
or \g131359/U$2 ( \54792 , \54787 , \54791 );
or \g131359/U$5 ( \54793 , \54790 , \48685 );
nand \g131359/U$1 ( \54794 , \54792 , \54793 );
xor \g131312/U$1_r1 ( \54795 , \54786 , \54794 );
not \g131311/U$1 ( \54796 , \54795 );
not \g131663/U$3 ( \54797 , \48323 );
and \g131695/U$2 ( \54798 , \52108 , \48335 );
and \g131695/U$3 ( \54799 , \48334 , \51854 );
nor \g131695/U$1 ( \54800 , \54798 , \54799 );
not \g131663/U$4 ( \54801 , \54800 );
or \g131663/U$2 ( \54802 , \54797 , \54801 );
or \g131663/U$5 ( \54803 , \54800 , \48323 );
nand \g131663/U$1 ( \54804 , \54802 , \54803 );
not \g131552/U$3 ( \54805 , \48483 );
and \g131582/U$2 ( \54806 , \51604 , \48479 );
and \g131582/U$3 ( \54807 , \48478 , \51564 );
nor \g131582/U$1 ( \54808 , \54806 , \54807 );
not \g131552/U$4 ( \54809 , \54808 );
or \g131552/U$2 ( \54810 , \54805 , \54809 );
or \g131552/U$5 ( \54811 , \54808 , \48483 );
nand \g131552/U$1 ( \54812 , \54810 , \54811 );
xor \g456120/U$4 ( \54813 , \54804 , \54812 );
not \g131416/U$3 ( \54814 , \48685 );
and \g131448/U$2 ( \54815 , \51117 , \48858 );
and \g131448/U$3 ( \54816 , \48860 , \51098 );
nor \g131448/U$1 ( \54817 , \54815 , \54816 );
not \g131416/U$4 ( \54818 , \54817 );
or \g131416/U$2 ( \54819 , \54814 , \54818 );
or \g131416/U$5 ( \54820 , \54817 , \48685 );
nand \g131416/U$1 ( \54821 , \54819 , \54820 );
and \g456120/U$3 ( \54822 , \54813 , \54821 );
and \g456120/U$5 ( \54823 , \54804 , \54812 );
nor \g456120/U$2 ( \54824 , \54822 , \54823 );
or \g131090/U$2 ( \54825 , \54796 , \54824 );
not \g131094/U$3 ( \54826 , \54824 );
not \g131094/U$4 ( \54827 , \54796 );
or \g131094/U$2 ( \54828 , \54826 , \54827 );
not \g131301/U$3 ( \54829 , \49014 );
and \g131325/U$2 ( \54830 , \50957 , \49075 );
and \g131325/U$3 ( \54831 , \49074 , \50752 );
nor \g131325/U$1 ( \54832 , \54830 , \54831 );
not \g131301/U$4 ( \54833 , \54832 );
or \g131301/U$2 ( \54834 , \54829 , \54833 );
or \g131301/U$5 ( \54835 , \54832 , \49014 );
nand \g131301/U$1 ( \54836 , \54834 , \54835 );
not \g132182/U$3 ( \54837 , \54535 );
not \g132182/U$4 ( \54838 , \54538 );
and \g132182/U$2 ( \54839 , \54837 , \54838 );
and \g132182/U$5 ( \54840 , \54535 , \54538 );
nor \g132182/U$1 ( \54841 , \54839 , \54840 );
and \g132429/U$2 ( \54842 , \47914 , \54185 );
and \g132429/U$3 ( \54843 , \54015 , \47913 );
nor \g132429/U$1 ( \54844 , \54842 , \54843 );
and \g132350/U$2 ( \54845 , \54844 , \47976 );
not \g132350/U$4 ( \54846 , \54844 );
and \g132350/U$3 ( \54847 , \54846 , \47977 );
nor \g132350/U$1 ( \54848 , \54845 , \54847 );
or \g132111/U$2 ( \54849 , \54841 , \54848 );
not \g132114/U$3 ( \54850 , \54848 );
not \g132114/U$4 ( \54851 , \54841 );
or \g132114/U$2 ( \54852 , \54850 , \54851 );
xor \g132831/U$1 ( \54853 , \47317 , \47271 );
not \g135539/U$2 ( \54854 , \54853 );
nor \g135539/U$1 ( \54855 , \54854 , \40060 );
not \g132190/U$2 ( \54856 , \54855 );
and \g132283/U$2 ( \54857 , \47960 , \54537 );
and \g132283/U$3 ( \54858 , \54529 , \47959 );
nor \g132283/U$1 ( \54859 , \54857 , \54858 );
not \g132230/U$3 ( \54860 , \54859 );
not \g132230/U$4 ( \54861 , \47948 );
and \g132230/U$2 ( \54862 , \54860 , \54861 );
and \g132230/U$5 ( \54863 , \54859 , \47948 );
nor \g132230/U$1 ( \54864 , \54862 , \54863 );
nor \g132190/U$1 ( \54865 , \54856 , \54864 );
nand \g132114/U$1 ( \54866 , \54852 , \54865 );
nand \g132111/U$1 ( \54867 , \54849 , \54866 );
xor \g131124/U$4 ( \54868 , \54836 , \54867 );
not \g131187/U$3 ( \54869 , \49233 );
and \g131217/U$2 ( \54870 , \50305 , \49403 );
and \g131217/U$3 ( \54871 , \49405 , \50443 );
nor \g131217/U$1 ( \54872 , \54870 , \54871 );
not \g131187/U$4 ( \54873 , \54872 );
or \g131187/U$2 ( \54874 , \54869 , \54873 );
or \g131187/U$5 ( \54875 , \54872 , \49233 );
nand \g131187/U$1 ( \54876 , \54874 , \54875 );
and \g131124/U$3 ( \54877 , \54868 , \54876 );
and \g131124/U$5 ( \54878 , \54836 , \54867 );
or \g131124/U$2 ( \54879 , \54877 , \54878 );
nand \g131094/U$1 ( \54880 , \54828 , \54879 );
nand \g131090/U$1 ( \54881 , \54825 , \54880 );
not \g130247/U$3 ( \54882 , \54881 );
xor \g131312/U$4 ( \54883 , \54777 , \54785 );
and \g131312/U$3 ( \54884 , \54883 , \54794 );
and \g131312/U$5 ( \54885 , \54777 , \54785 );
or \g131312/U$2 ( \54886 , \54884 , \54885 );
xor \g131738/U$1 ( \54887 , \54262 , \54270 );
xor \g131738/U$1_r1 ( \54888 , \54887 , \54279 );
xor \g130975/U$1 ( \54889 , \54886 , \54888 );
not \g131028/U$3 ( \54890 , \49233 );
and \g131069/U$2 ( \54891 , \49888 , \49403 );
and \g131069/U$3 ( \54892 , \49405 , \50019 );
nor \g131069/U$1 ( \54893 , \54891 , \54892 );
not \g131028/U$4 ( \54894 , \54893 );
or \g131028/U$2 ( \54895 , \54890 , \54894 );
or \g131028/U$5 ( \54896 , \54893 , \49233 );
nand \g131028/U$1 ( \54897 , \54895 , \54896 );
xor \g130975/U$1_r1 ( \54898 , \54889 , \54897 );
not \g130247/U$4 ( \54899 , \54898 );
or \g130247/U$2 ( \54900 , \54882 , \54899 );
or \g130254/U$2 ( \54901 , \54898 , \54881 );
and \g130824/U$2 ( \54902 , \49282 , \50588 );
and \g130824/U$3 ( \54903 , \50587 , \49158 );
nor \g130824/U$1 ( \54904 , \54902 , \54903 );
not \g130797/U$3 ( \54905 , \54904 );
not \g130797/U$4 ( \54906 , \50362 );
and \g130797/U$2 ( \54907 , \54905 , \54906 );
and \g130797/U$5 ( \54908 , \54904 , \50362 );
nor \g130797/U$1 ( \54909 , \54907 , \54908 );
and \g130935/U$2 ( \54910 , \49512 , \50159 );
and \g130935/U$3 ( \54911 , \50160 , \49714 );
nor \g130935/U$1 ( \54912 , \54910 , \54911 );
not \g130907/U$3 ( \54913 , \54912 );
not \g130907/U$4 ( \54914 , \49925 );
and \g130907/U$2 ( \54915 , \54913 , \54914 );
and \g130907/U$5 ( \54916 , \54912 , \49925 );
nor \g130907/U$1 ( \54917 , \54915 , \54916 );
xor \g130501/U$4 ( \54918 , \54909 , \54917 );
and \g130589/U$2 ( \54919 , \48726 , \51517 );
and \g130589/U$3 ( \54920 , \51518 , \48833 );
nor \g130589/U$1 ( \54921 , \54919 , \54920 );
not \g130560/U$3 ( \54922 , \54921 );
not \g130560/U$4 ( \54923 , \51124 );
and \g130560/U$2 ( \54924 , \54922 , \54923 );
and \g130560/U$5 ( \54925 , \54921 , \51124 );
nor \g130560/U$1 ( \54926 , \54924 , \54925 );
and \g130501/U$3 ( \54927 , \54918 , \54926 );
and \g130501/U$5 ( \54928 , \54909 , \54917 );
or \g130501/U$2 ( \54929 , \54927 , \54928 );
xor \g131048/U$1 ( \54930 , \54709 , \54713 );
xor \g131048/U$1_r1 ( \54931 , \54930 , \54722 );
not \g131046/U$1 ( \54932 , \54931 );
or \g130324/U$2 ( \54933 , \54929 , \54932 );
not \g130330/U$3 ( \54934 , \54932 );
not \g130330/U$4 ( \54935 , \54929 );
or \g130330/U$2 ( \54936 , \54934 , \54935 );
not \g131029/U$3 ( \54937 , \49568 );
and \g131070/U$2 ( \54938 , \49888 , \49812 );
and \g131070/U$3 ( \54939 , \49813 , \50019 );
nor \g131070/U$1 ( \54940 , \54938 , \54939 );
not \g131029/U$4 ( \54941 , \54940 );
or \g131029/U$2 ( \54942 , \54937 , \54941 );
or \g131029/U$5 ( \54943 , \54940 , \49568 );
nand \g131029/U$1 ( \54944 , \54942 , \54943 );
and \g132050/U$2 ( \54945 , \52978 , \48063 );
and \g132050/U$3 ( \54946 , \48064 , \53300 );
nor \g132050/U$1 ( \54947 , \54945 , \54946 );
not \g132012/U$3 ( \54948 , \54947 );
not \g132012/U$4 ( \54949 , \47997 );
and \g132012/U$2 ( \54950 , \54948 , \54949 );
and \g132012/U$5 ( \54951 , \54947 , \47997 );
nor \g132012/U$1 ( \54952 , \54950 , \54951 );
and \g132203/U$2 ( \54953 , \53610 , \47930 );
and \g132203/U$3 ( \54954 , \53848 , \47931 );
nor \g132203/U$1 ( \54955 , \54953 , \54954 );
not \g132158/U$3 ( \54956 , \54955 );
not \g132158/U$4 ( \54957 , \47935 );
and \g132158/U$2 ( \54958 , \54956 , \54957 );
and \g132158/U$5 ( \54959 , \54955 , \47935 );
nor \g132158/U$1 ( \54960 , \54958 , \54959 );
or \g131829/U$2 ( \54961 , \54952 , \54960 );
and \g131833/U$2 ( \54962 , \54952 , \54960 );
and \g131897/U$2 ( \54963 , \52620 , \48154 );
and \g131897/U$3 ( \54964 , \48155 , \52883 );
nor \g131897/U$1 ( \54965 , \54963 , \54964 );
not \g131858/U$3 ( \54966 , \54965 );
not \g131858/U$4 ( \54967 , \48159 );
and \g131858/U$2 ( \54968 , \54966 , \54967 );
and \g131858/U$5 ( \54969 , \54965 , \48159 );
nor \g131858/U$1 ( \54970 , \54968 , \54969 );
nor \g131833/U$1 ( \54971 , \54962 , \54970 );
not \g131832/U$1 ( \54972 , \54971 );
nand \g131829/U$1 ( \54973 , \54961 , \54972 );
xor \g130360/U$4 ( \54974 , \54944 , \54973 );
not \g130422/U$3 ( \54975 , \51120 );
and \g130451/U$2 ( \54976 , \48568 , \52273 );
and \g130451/U$3 ( \54977 , \52270 , \48515 );
nor \g130451/U$1 ( \54978 , \54976 , \54977 );
not \g130422/U$4 ( \54979 , \54978 );
or \g130422/U$2 ( \54980 , \54975 , \54979 );
or \g130422/U$5 ( \54981 , \54978 , \51120 );
nand \g130422/U$1 ( \54982 , \54980 , \54981 );
and \g130360/U$3 ( \54983 , \54974 , \54982 );
and \g130360/U$5 ( \54984 , \54944 , \54973 );
or \g130360/U$2 ( \54985 , \54983 , \54984 );
nand \g130330/U$1 ( \54986 , \54936 , \54985 );
nand \g130324/U$1 ( \54987 , \54933 , \54986 );
nand \g130254/U$1 ( \54988 , \54901 , \54987 );
nand \g130247/U$1 ( \54989 , \54900 , \54988 );
xor \g129959/U$1 ( \54990 , \54769 , \54989 );
xor \g456047/U$2 ( \54991 , \54250 , \54282 );
xor \g456047/U$1 ( \54992 , \54991 , \54291 );
xor \g130975/U$4 ( \54993 , \54886 , \54888 );
and \g130975/U$3 ( \54994 , \54993 , \54897 );
and \g130975/U$5 ( \54995 , \54886 , \54888 );
or \g130975/U$2 ( \54996 , \54994 , \54995 );
xor \g130139/U$1 ( \54997 , \54305 , \54313 );
xor \g130139/U$1_r1 ( \54998 , \54997 , \54322 );
xor \g456047/U$1_r1 ( \54999 , \54996 , \54998 );
xor \g456047/U$1_r2 ( \55000 , \54992 , \54999 );
xor \g129959/U$1_r1 ( \55001 , \54990 , \55000 );
xor \g456137/U$4 ( \55002 , \54640 , \54648 );
and \g456137/U$3 ( \55003 , \55002 , \54657 );
and \g456137/U$5 ( \55004 , \54640 , \54648 );
nor \g456137/U$2 ( \55005 , \55003 , \55004 );
not \g131704/U$3 ( \55006 , \54365 );
xor \g131810/U$1 ( \55007 , \54355 , \54347 );
not \g131704/U$4 ( \55008 , \55007 );
and \g131704/U$2 ( \55009 , \55006 , \55008 );
and \g131704/U$5 ( \55010 , \54365 , \55007 );
nor \g131704/U$1 ( \55011 , \55009 , \55010 );
xor \g131034/U$1 ( \55012 , \55005 , \55011 );
xor \g456105/U$4 ( \55013 , \54739 , \54747 );
and \g456105/U$3 ( \55014 , \55013 , \54756 );
and \g456105/U$5 ( \55015 , \54739 , \54747 );
nor \g456105/U$2 ( \55016 , \55014 , \55015 );
xor \g131034/U$1_r1 ( \55017 , \55012 , \55016 );
not \g130038/U$3 ( \55018 , \55017 );
xor \g456063/U$4 ( \55019 , \54658 , \54700 );
and \g456063/U$3 ( \55020 , \55019 , \54725 );
and \g456063/U$5 ( \55021 , \54658 , \54700 );
nor \g456063/U$2 ( \55022 , \55020 , \55021 );
not \g130059/U$3 ( \55023 , \55022 );
xor \g131563/U$1 ( \55024 , \54184 , \54195 );
xor \g131563/U$1_r1 ( \55025 , \55024 , \54204 );
not \g130685/U$3 ( \55026 , \50362 );
and \g130711/U$2 ( \55027 , \49102 , \50588 );
and \g130711/U$3 ( \55028 , \50587 , \48977 );
nor \g130711/U$1 ( \55029 , \55027 , \55028 );
not \g130685/U$4 ( \55030 , \55029 );
or \g130685/U$2 ( \55031 , \55026 , \55030 );
or \g130685/U$5 ( \55032 , \55029 , \50362 );
nand \g130685/U$1 ( \55033 , \55031 , \55032 );
not \g131415/U$3 ( \55034 , \48483 );
and \g131447/U$2 ( \55035 , \51117 , \48478 );
and \g131447/U$3 ( \55036 , \48479 , \51098 );
nor \g131447/U$1 ( \55037 , \55035 , \55036 );
not \g131415/U$4 ( \55038 , \55037 );
or \g131415/U$2 ( \55039 , \55034 , \55038 );
or \g131415/U$5 ( \55040 , \55037 , \48483 );
nand \g131415/U$1 ( \55041 , \55039 , \55040 );
xor \g130221/U$4 ( \55042 , \55033 , \55041 );
not \g130279/U$3 ( \55043 , \51120 );
and \g130313/U$2 ( \55044 , \48349 , \52273 );
and \g130313/U$3 ( \55045 , \52270 , \48353 );
nor \g130313/U$1 ( \55046 , \55044 , \55045 );
not \g130279/U$4 ( \55047 , \55046 );
or \g130279/U$2 ( \55048 , \55043 , \55047 );
or \g130279/U$5 ( \55049 , \55046 , \51120 );
nand \g130279/U$1 ( \55050 , \55048 , \55049 );
and \g130221/U$3 ( \55051 , \55042 , \55050 );
and \g130221/U$5 ( \55052 , \55033 , \55041 );
or \g130221/U$2 ( \55053 , \55051 , \55052 );
xor \g456052/U$1 ( \55054 , \55025 , \55053 );
not \g130796/U$3 ( \55055 , \49925 );
and \g130823/U$2 ( \55056 , \49282 , \50160 );
and \g130823/U$3 ( \55057 , \50159 , \49158 );
nor \g130823/U$1 ( \55058 , \55056 , \55057 );
not \g130796/U$4 ( \55059 , \55058 );
or \g130796/U$2 ( \55060 , \55055 , \55059 );
or \g130796/U$5 ( \55061 , \55058 , \49925 );
nand \g130796/U$1 ( \55062 , \55060 , \55061 );
xor \g131936/U$4 ( \55063 , \54605 , \54613 );
and \g131936/U$3 ( \55064 , \55063 , \54625 );
and \g131936/U$5 ( \55065 , \54605 , \54613 );
or \g131936/U$2 ( \55066 , \55064 , \55065 );
xor \g130359/U$4 ( \55067 , \55062 , \55066 );
not \g130421/U$3 ( \55068 , \51124 );
and \g130450/U$2 ( \55069 , \48568 , \51518 );
and \g130450/U$3 ( \55070 , \51517 , \48515 );
nor \g130450/U$1 ( \55071 , \55069 , \55070 );
not \g130421/U$4 ( \55072 , \55071 );
or \g130421/U$2 ( \55073 , \55068 , \55072 );
or \g130421/U$5 ( \55074 , \55071 , \51124 );
nand \g130421/U$1 ( \55075 , \55073 , \55074 );
and \g130359/U$3 ( \55076 , \55067 , \55075 );
and \g130359/U$5 ( \55077 , \55062 , \55066 );
or \g130359/U$2 ( \55078 , \55076 , \55077 );
xor \g456052/U$1_r1 ( \55079 , \55054 , \55078 );
not \g130059/U$4 ( \55080 , \55079 );
or \g130059/U$2 ( \55081 , \55023 , \55080 );
or \g130059/U$5 ( \55082 , \55079 , \55022 );
nand \g130059/U$1 ( \55083 , \55081 , \55082 );
not \g130038/U$4 ( \55084 , \55083 );
or \g130038/U$2 ( \55085 , \55018 , \55084 );
or \g130038/U$5 ( \55086 , \55083 , \55017 );
nand \g130038/U$1 ( \55087 , \55085 , \55086 );
not \g129907/U$3 ( \55088 , \55087 );
xnor \g455951/U$1 ( \55089 , \54987 , \54898 );
not \g130209/U$3 ( \55090 , \55089 );
not \g130209/U$4 ( \55091 , \54881 );
and \g130209/U$2 ( \55092 , \55090 , \55091 );
and \g130209/U$5 ( \55093 , \55089 , \54881 );
nor \g130209/U$1 ( \55094 , \55092 , \55093 );
xor \g456120/U$1 ( \55095 , \54804 , \54812 );
xor \g456120/U$1_r1 ( \55096 , \55095 , \54821 );
xor \g456143/U$1 ( \55097 , \54674 , \54682 );
xor \g456143/U$1_r1 ( \55098 , \55097 , \54684 );
and \g131010/U$2 ( \55099 , \55096 , \55098 );
not \g131015/U$3 ( \55100 , \55096 );
not \g131015/U$4 ( \55101 , \55098 );
and \g131015/U$2 ( \55102 , \55100 , \55101 );
and \g131381/U$2 ( \55103 , \51117 , \49075 );
and \g131381/U$3 ( \55104 , \49074 , \50957 );
nor \g131381/U$1 ( \55105 , \55103 , \55104 );
not \g131360/U$3 ( \55106 , \55105 );
not \g131360/U$4 ( \55107 , \49014 );
and \g131360/U$2 ( \55108 , \55106 , \55107 );
and \g131360/U$5 ( \55109 , \55105 , \49014 );
nor \g131360/U$1 ( \55110 , \55108 , \55109 );
not \g132184/U$3 ( \55111 , \54864 );
not \g132184/U$4 ( \55112 , \54855 );
and \g132184/U$2 ( \55113 , \55111 , \55112 );
and \g132184/U$5 ( \55114 , \54864 , \54855 );
nor \g132184/U$1 ( \55115 , \55113 , \55114 );
not \g132112/U$3 ( \55116 , \55115 );
and \g132432/U$2 ( \55117 , \47913 , \54185 );
and \g132432/U$3 ( \55118 , \54251 , \47914 );
nor \g132432/U$1 ( \55119 , \55117 , \55118 );
and \g132352/U$2 ( \55120 , \55119 , \47976 );
not \g132352/U$4 ( \55121 , \55119 );
and \g132352/U$3 ( \55122 , \55121 , \47977 );
nor \g132352/U$1 ( \55123 , \55120 , \55122 );
not \g132112/U$4 ( \55124 , \55123 );
and \g132112/U$2 ( \55125 , \55116 , \55124 );
and \g132115/U$2 ( \55126 , \55115 , \55123 );
xor \g132887/U$1 ( \55127 , \46605 , \47269 );
nand \g132382/U$1 ( \55128 , \55127 , \40061 );
not \g132191/U$2 ( \55129 , \55128 );
not \g132231/U$3 ( \55130 , \47948 );
and \g132284/U$2 ( \55131 , \47960 , \54853 );
and \g132284/U$3 ( \55132 , \54537 , \47959 );
nor \g132284/U$1 ( \55133 , \55131 , \55132 );
not \g132231/U$4 ( \55134 , \55133 );
or \g132231/U$2 ( \55135 , \55130 , \55134 );
or \g132231/U$5 ( \55136 , \55133 , \47948 );
nand \g132231/U$1 ( \55137 , \55135 , \55136 );
nand \g132191/U$1 ( \55138 , \55129 , \55137 );
nor \g132115/U$1 ( \55139 , \55126 , \55138 );
nor \g132112/U$1 ( \55140 , \55125 , \55139 );
xor \g456081/U$5 ( \55141 , \55110 , \55140 );
and \g131146/U$2 ( \55142 , \50305 , \49813 );
and \g131146/U$3 ( \55143 , \49812 , \50019 );
nor \g131146/U$1 ( \55144 , \55142 , \55143 );
not \g131112/U$3 ( \55145 , \55144 );
not \g131112/U$4 ( \55146 , \49568 );
and \g131112/U$2 ( \55147 , \55145 , \55146 );
and \g131112/U$5 ( \55148 , \55144 , \49568 );
nor \g131112/U$1 ( \55149 , \55147 , \55148 );
and \g456081/U$4 ( \55150 , \55141 , \55149 );
and \g456081/U$6 ( \55151 , \55110 , \55140 );
or \g456081/U$3 ( \55152 , \55150 , \55151 );
nor \g131015/U$1 ( \55153 , \55102 , \55152 );
nor \g131010/U$1 ( \55154 , \55099 , \55153 );
not \g131087/U$3 ( \55155 , \54879 );
not \g131087/U$4 ( \55156 , \54824 );
and \g131087/U$2 ( \55157 , \55155 , \55156 );
and \g131087/U$5 ( \55158 , \54879 , \54824 );
nor \g131087/U$1 ( \55159 , \55157 , \55158 );
not \g131056/U$3 ( \55160 , \55159 );
not \g131056/U$4 ( \55161 , \54795 );
and \g131056/U$2 ( \55162 , \55160 , \55161 );
and \g131056/U$5 ( \55163 , \55159 , \54795 );
nor \g131056/U$1 ( \55164 , \55162 , \55163 );
xor \g130350/U$4 ( \55165 , \55154 , \55164 );
not \g130458/U$3 ( \55166 , \54697 );
xor \g130810/U$1 ( \55167 , \54687 , \54666 );
not \g130458/U$4 ( \55168 , \55167 );
and \g130458/U$2 ( \55169 , \55166 , \55168 );
and \g130458/U$5 ( \55170 , \54697 , \55167 );
nor \g130458/U$1 ( \55171 , \55169 , \55170 );
and \g130350/U$3 ( \55172 , \55165 , \55171 );
and \g130350/U$5 ( \55173 , \55154 , \55164 );
or \g130350/U$2 ( \55174 , \55172 , \55173 );
or \g130086/U$2 ( \55175 , \55094 , \55174 );
and \g130104/U$2 ( \55176 , \55094 , \55174 );
xor \g130221/U$1 ( \55177 , \55033 , \55041 );
xor \g130221/U$1_r1 ( \55178 , \55177 , \55050 );
xor \g131676/U$4 ( \55179 , \54561 , \54569 );
and \g131676/U$3 ( \55180 , \55179 , \54578 );
and \g131676/U$5 ( \55181 , \54561 , \54569 );
or \g131676/U$2 ( \55182 , \55180 , \55181 );
not \g130906/U$3 ( \55183 , \49568 );
and \g130934/U$2 ( \55184 , \49512 , \49812 );
and \g130934/U$3 ( \55185 , \49813 , \49714 );
nor \g130934/U$1 ( \55186 , \55184 , \55185 );
not \g130906/U$4 ( \55187 , \55186 );
or \g130906/U$2 ( \55188 , \55183 , \55187 );
or \g130906/U$5 ( \55189 , \55186 , \49568 );
nand \g130906/U$1 ( \55190 , \55188 , \55189 );
xor \g456071/U$1 ( \55191 , \55182 , \55190 );
not \g130559/U$3 ( \55192 , \50759 );
and \g130588/U$2 ( \55193 , \48726 , \51053 );
and \g130588/U$3 ( \55194 , \51055 , \48833 );
nor \g130588/U$1 ( \55195 , \55193 , \55194 );
not \g130559/U$4 ( \55196 , \55195 );
or \g130559/U$2 ( \55197 , \55192 , \55196 );
or \g130559/U$5 ( \55198 , \55195 , \50759 );
nand \g130559/U$1 ( \55199 , \55197 , \55198 );
xor \g456071/U$1_r1 ( \55200 , \55191 , \55199 );
xnor \g455950/U$1 ( \55201 , \55178 , \55200 );
not \g130142/U$3 ( \55202 , \55201 );
xor \g130359/U$1 ( \55203 , \55062 , \55066 );
xor \g130359/U$1_r1 ( \55204 , \55203 , \55075 );
not \g130142/U$4 ( \55205 , \55204 );
and \g130142/U$2 ( \55206 , \55202 , \55205 );
and \g130142/U$5 ( \55207 , \55201 , \55204 );
nor \g130142/U$1 ( \55208 , \55206 , \55207 );
nor \g130104/U$1 ( \55209 , \55176 , \55208 );
not \g130103/U$1 ( \55210 , \55209 );
nand \g130086/U$1 ( \55211 , \55175 , \55210 );
xor \g456055/U$4 ( \55212 , \54757 , \54761 );
and \g456055/U$3 ( \55213 , \55212 , \54766 );
and \g456055/U$5 ( \55214 , \54757 , \54761 );
nor \g456055/U$2 ( \55215 , \55213 , \55214 );
not \g130039/U$3 ( \55216 , \55215 );
not \g131079/U$3 ( \55217 , \54236 );
xor \g131204/U$1 ( \55218 , \54226 , \54218 );
not \g131079/U$4 ( \55219 , \55218 );
and \g131079/U$2 ( \55220 , \55217 , \55219 );
and \g131079/U$5 ( \55221 , \54236 , \55218 );
nor \g131079/U$1 ( \55222 , \55220 , \55221 );
not \g130401/U$3 ( \55223 , \55222 );
not \g130963/U$3 ( \55224 , \49233 );
and \g130990/U$2 ( \55225 , \49888 , \49405 );
and \g130990/U$3 ( \55226 , \49403 , \49714 );
nor \g130990/U$1 ( \55227 , \55225 , \55226 );
not \g130963/U$4 ( \55228 , \55227 );
or \g130963/U$2 ( \55229 , \55224 , \55228 );
or \g130963/U$5 ( \55230 , \55227 , \49233 );
nand \g130963/U$1 ( \55231 , \55229 , \55230 );
not \g130852/U$3 ( \55232 , \49568 );
and \g130876/U$2 ( \55233 , \49512 , \49813 );
and \g130876/U$3 ( \55234 , \49812 , \49282 );
nor \g130876/U$1 ( \55235 , \55233 , \55234 );
not \g130852/U$4 ( \55236 , \55235 );
or \g130852/U$2 ( \55237 , \55232 , \55236 );
or \g130852/U$5 ( \55238 , \55235 , \49568 );
nand \g130852/U$1 ( \55239 , \55237 , \55238 );
xor \g456067/U$1 ( \55240 , \55231 , \55239 );
not \g130491/U$3 ( \55241 , \50759 );
and \g130522/U$2 ( \55242 , \48726 , \51055 );
and \g130522/U$3 ( \55243 , \51053 , \48568 );
nor \g130522/U$1 ( \55244 , \55242 , \55243 );
not \g130491/U$4 ( \55245 , \55244 );
or \g130491/U$2 ( \55246 , \55241 , \55245 );
or \g130491/U$5 ( \55247 , \55244 , \50759 );
nand \g130491/U$1 ( \55248 , \55246 , \55247 );
xor \g456067/U$1_r1 ( \55249 , \55240 , \55248 );
not \g130401/U$4 ( \55250 , \55249 );
or \g130401/U$2 ( \55251 , \55223 , \55250 );
or \g130401/U$5 ( \55252 , \55249 , \55222 );
nand \g130401/U$1 ( \55253 , \55251 , \55252 );
not \g130361/U$3 ( \55254 , \55253 );
xor \g456071/U$4 ( \55255 , \55182 , \55190 );
and \g456071/U$3 ( \55256 , \55255 , \55199 );
and \g456071/U$5 ( \55257 , \55182 , \55190 );
nor \g456071/U$2 ( \55258 , \55256 , \55257 );
not \g130361/U$4 ( \55259 , \55258 );
and \g130361/U$2 ( \55260 , \55254 , \55259 );
and \g130361/U$5 ( \55261 , \55253 , \55258 );
nor \g130361/U$1 ( \55262 , \55260 , \55261 );
not \g130060/U$3 ( \55263 , \55262 );
not \g130185/U$3 ( \55264 , \55200 );
not \g130185/U$4 ( \55265 , \55204 );
or \g130185/U$2 ( \55266 , \55264 , \55265 );
or \g130188/U$2 ( \55267 , \55204 , \55200 );
nand \g130188/U$1 ( \55268 , \55267 , \55178 );
nand \g130185/U$1 ( \55269 , \55266 , \55268 );
not \g130060/U$4 ( \55270 , \55269 );
or \g130060/U$2 ( \55271 , \55263 , \55270 );
or \g130060/U$5 ( \55272 , \55269 , \55262 );
nand \g130060/U$1 ( \55273 , \55271 , \55272 );
not \g130039/U$4 ( \55274 , \55273 );
or \g130039/U$2 ( \55275 , \55216 , \55274 );
or \g130039/U$5 ( \55276 , \55273 , \55215 );
nand \g130039/U$1 ( \55277 , \55275 , \55276 );
xnor \g129950/U$1 ( \55278 , \55211 , \55277 );
not \g129907/U$4 ( \55279 , \55278 );
or \g129907/U$2 ( \55280 , \55088 , \55279 );
or \g129907/U$5 ( \55281 , \55278 , \55087 );
nand \g129907/U$1 ( \55282 , \55280 , \55281 );
xor \g456030/U$4 ( \55283 , \55001 , \55282 );
not \g131792/U$3 ( \55284 , \48323 );
and \g131823/U$2 ( \55285 , \52620 , \48335 );
and \g131823/U$3 ( \55286 , \48334 , \52352 );
nor \g131823/U$1 ( \55287 , \55285 , \55286 );
not \g131792/U$4 ( \55288 , \55287 );
or \g131792/U$2 ( \55289 , \55284 , \55288 );
or \g131792/U$5 ( \55290 , \55287 , \48323 );
nand \g131792/U$1 ( \55291 , \55289 , \55290 );
not \g131931/U$3 ( \55292 , \48159 );
and \g131961/U$2 ( \55293 , \52978 , \48155 );
and \g131961/U$3 ( \55294 , \48154 , \52883 );
nor \g131961/U$1 ( \55295 , \55293 , \55294 );
not \g131931/U$4 ( \55296 , \55295 );
or \g131931/U$2 ( \55297 , \55292 , \55296 );
or \g131931/U$5 ( \55298 , \55295 , \48159 );
nand \g131931/U$1 ( \55299 , \55297 , \55298 );
xor \g131497/U$4 ( \55300 , \55291 , \55299 );
not \g131553/U$3 ( \55301 , \48685 );
and \g131583/U$2 ( \55302 , \51604 , \48860 );
and \g131583/U$3 ( \55303 , \48858 , \51564 );
nor \g131583/U$1 ( \55304 , \55302 , \55303 );
not \g131553/U$4 ( \55305 , \55304 );
or \g131553/U$2 ( \55306 , \55301 , \55305 );
or \g131553/U$5 ( \55307 , \55304 , \48685 );
nand \g131553/U$1 ( \55308 , \55306 , \55307 );
and \g131497/U$3 ( \55309 , \55300 , \55308 );
and \g131497/U$5 ( \55310 , \55291 , \55299 );
or \g131497/U$2 ( \55311 , \55309 , \55310 );
not \g131091/U$3 ( \55312 , \55311 );
not \g131664/U$3 ( \55313 , \48483 );
and \g131696/U$2 ( \55314 , \52108 , \48479 );
and \g131696/U$3 ( \55315 , \48478 , \51854 );
nor \g131696/U$1 ( \55316 , \55314 , \55315 );
not \g131664/U$4 ( \55317 , \55316 );
or \g131664/U$2 ( \55318 , \55313 , \55317 );
or \g131664/U$5 ( \55319 , \55316 , \48483 );
nand \g131664/U$1 ( \55320 , \55318 , \55319 );
not \g132353/U$3 ( \55321 , \47935 );
and \g132433/U$2 ( \55322 , \47931 , \54185 );
and \g132433/U$3 ( \55323 , \54015 , \47930 );
nor \g132433/U$1 ( \55324 , \55322 , \55323 );
not \g132353/U$4 ( \55325 , \55324 );
or \g132353/U$2 ( \55326 , \55321 , \55325 );
or \g132353/U$5 ( \55327 , \55324 , \47935 );
nand \g132353/U$1 ( \55328 , \55326 , \55327 );
not \g132160/U$3 ( \55329 , \47997 );
and \g132204/U$2 ( \55330 , \53610 , \48063 );
and \g132204/U$3 ( \55331 , \48064 , \53848 );
nor \g132204/U$1 ( \55332 , \55330 , \55331 );
not \g132160/U$4 ( \55333 , \55332 );
or \g132160/U$2 ( \55334 , \55329 , \55333 );
or \g132160/U$5 ( \55335 , \55332 , \47997 );
nand \g132160/U$1 ( \55336 , \55334 , \55335 );
xor \g131948/U$4 ( \55337 , \55328 , \55336 );
not \g132013/U$3 ( \55338 , \48159 );
and \g132051/U$2 ( \55339 , \52978 , \48154 );
and \g132051/U$3 ( \55340 , \48155 , \53300 );
nor \g132051/U$1 ( \55341 , \55339 , \55340 );
not \g132013/U$4 ( \55342 , \55341 );
or \g132013/U$2 ( \55343 , \55338 , \55342 );
or \g132013/U$5 ( \55344 , \55341 , \48159 );
nand \g132013/U$1 ( \55345 , \55343 , \55344 );
and \g131948/U$3 ( \55346 , \55337 , \55345 );
and \g131948/U$5 ( \55347 , \55328 , \55336 );
or \g131948/U$2 ( \55348 , \55346 , \55347 );
xor \g131367/U$4 ( \55349 , \55320 , \55348 );
not \g131417/U$3 ( \55350 , \49014 );
and \g131449/U$2 ( \55351 , \51117 , \49074 );
and \g131449/U$3 ( \55352 , \49075 , \51098 );
nor \g131449/U$1 ( \55353 , \55351 , \55352 );
not \g131417/U$4 ( \55354 , \55353 );
or \g131417/U$2 ( \55355 , \55350 , \55354 );
or \g131417/U$5 ( \55356 , \55353 , \49014 );
nand \g131417/U$1 ( \55357 , \55355 , \55356 );
and \g131367/U$3 ( \55358 , \55349 , \55357 );
and \g131367/U$5 ( \55359 , \55320 , \55348 );
or \g131367/U$2 ( \55360 , \55358 , \55359 );
not \g131091/U$4 ( \55361 , \55360 );
or \g131091/U$2 ( \55362 , \55312 , \55361 );
or \g131095/U$2 ( \55363 , \55360 , \55311 );
not \g131302/U$3 ( \55364 , \49233 );
and \g131326/U$2 ( \55365 , \50957 , \49405 );
and \g131326/U$3 ( \55366 , \49403 , \50752 );
nor \g131326/U$1 ( \55367 , \55365 , \55366 );
not \g131302/U$4 ( \55368 , \55367 );
or \g131302/U$2 ( \55369 , \55364 , \55368 );
or \g131302/U$5 ( \55370 , \55367 , \49233 );
nand \g131302/U$1 ( \55371 , \55369 , \55370 );
not \g132102/U$3 ( \55372 , \55123 );
xor \g132118/U$1 ( \55373 , \55138 , \55115 );
not \g132102/U$4 ( \55374 , \55373 );
or \g132102/U$2 ( \55375 , \55372 , \55374 );
or \g132102/U$5 ( \55376 , \55373 , \55123 );
nand \g132102/U$1 ( \55377 , \55375 , \55376 );
xor \g131126/U$4 ( \55378 , \55371 , \55377 );
not \g131188/U$3 ( \55379 , \49568 );
and \g131218/U$2 ( \55380 , \50305 , \49812 );
and \g131218/U$3 ( \55381 , \49813 , \50443 );
nor \g131218/U$1 ( \55382 , \55380 , \55381 );
not \g131188/U$4 ( \55383 , \55382 );
or \g131188/U$2 ( \55384 , \55379 , \55383 );
or \g131188/U$5 ( \55385 , \55382 , \49568 );
nand \g131188/U$1 ( \55386 , \55384 , \55385 );
and \g131126/U$3 ( \55387 , \55378 , \55386 );
and \g131126/U$5 ( \55388 , \55371 , \55377 );
or \g131126/U$2 ( \55389 , \55387 , \55388 );
nand \g131095/U$1 ( \55390 , \55363 , \55389 );
nand \g131091/U$1 ( \55391 , \55362 , \55390 );
not \g131005/U$3 ( \55392 , \55096 );
not \g131005/U$4 ( \55393 , \55152 );
or \g131005/U$2 ( \55394 , \55392 , \55393 );
or \g131005/U$5 ( \55395 , \55152 , \55096 );
nand \g131005/U$1 ( \55396 , \55394 , \55395 );
xor \g455954/U$1 ( \55397 , \55098 , \55396 );
xor \g456061/U$4 ( \55398 , \55391 , \55397 );
xor \g130360/U$1 ( \55399 , \54944 , \54973 );
xor \g130360/U$1_r1 ( \55400 , \55399 , \54982 );
and \g456061/U$3 ( \55401 , \55398 , \55400 );
and \g456061/U$5 ( \55402 , \55391 , \55397 );
nor \g456061/U$2 ( \55403 , \55401 , \55402 );
xor \g130350/U$1 ( \55404 , \55154 , \55164 );
xor \g130350/U$1_r1 ( \55405 , \55404 , \55171 );
or \g130208/U$2 ( \55406 , \55403 , \55405 );
not \g130211/U$3 ( \55407 , \55405 );
not \g130211/U$4 ( \55408 , \55403 );
or \g130211/U$2 ( \55409 , \55407 , \55408 );
xor \g456059/U$1 ( \55410 , \54552 , \54589 );
xor \g456059/U$1_r1 ( \55411 , \55410 , \54636 );
nand \g130211/U$1 ( \55412 , \55409 , \55411 );
nand \g130208/U$1 ( \55413 , \55406 , \55412 );
not \g130140/U$1 ( \55414 , \55413 );
not \g131241/U$3 ( \55415 , \49233 );
and \g131273/U$2 ( \55416 , \50752 , \49405 );
and \g131273/U$3 ( \55417 , \49403 , \50443 );
nor \g131273/U$1 ( \55418 , \55416 , \55417 );
not \g131241/U$4 ( \55419 , \55418 );
or \g131241/U$2 ( \55420 , \55415 , \55419 );
or \g131241/U$5 ( \55421 , \55418 , \49233 );
nand \g131241/U$1 ( \55422 , \55420 , \55421 );
not \g130854/U$3 ( \55423 , \50362 );
and \g130878/U$2 ( \55424 , \49512 , \50588 );
and \g130878/U$3 ( \55425 , \50587 , \49282 );
nor \g130878/U$1 ( \55426 , \55424 , \55425 );
not \g130854/U$4 ( \55427 , \55426 );
or \g130854/U$2 ( \55428 , \55423 , \55427 );
or \g130854/U$5 ( \55429 , \55426 , \50362 );
nand \g130854/U$1 ( \55430 , \55428 , \55429 );
xor \g456078/U$4 ( \55431 , \55422 , \55430 );
not \g130623/U$3 ( \55432 , \51124 );
and \g130657/U$2 ( \55433 , \48833 , \51517 );
and \g130657/U$3 ( \55434 , \51518 , \48977 );
nor \g130657/U$1 ( \55435 , \55433 , \55434 );
not \g130623/U$4 ( \55436 , \55435 );
or \g130623/U$2 ( \55437 , \55432 , \55436 );
or \g130623/U$5 ( \55438 , \55435 , \51124 );
nand \g130623/U$1 ( \55439 , \55437 , \55438 );
and \g456078/U$3 ( \55440 , \55431 , \55439 );
and \g456078/U$5 ( \55441 , \55422 , \55430 );
nor \g456078/U$2 ( \55442 , \55440 , \55441 );
not \g132091/U$3 ( \55443 , \47997 );
and \g132131/U$2 ( \55444 , \53610 , \48064 );
and \g132131/U$3 ( \55445 , \48063 , \53300 );
nor \g132131/U$1 ( \55446 , \55444 , \55445 );
not \g132091/U$4 ( \55447 , \55446 );
or \g132091/U$2 ( \55448 , \55443 , \55447 );
or \g132091/U$5 ( \55449 , \55446 , \47997 );
nand \g132091/U$1 ( \55450 , \55448 , \55449 );
not \g132256/U$3 ( \55451 , \47935 );
and \g132305/U$2 ( \55452 , \53848 , \47930 );
and \g132305/U$3 ( \55453 , \54015 , \47931 );
nor \g132305/U$1 ( \55454 , \55452 , \55453 );
not \g132256/U$4 ( \55455 , \55454 );
or \g132256/U$2 ( \55456 , \55451 , \55455 );
or \g132256/U$5 ( \55457 , \55454 , \47935 );
nand \g132256/U$1 ( \55458 , \55456 , \55457 );
xor \g131981/U$4 ( \55459 , \55450 , \55458 );
xor \g132957/U$1 ( \55460 , \46696 , \47267 );
not \g135542/U$2 ( \55461 , \55460 );
nor \g135542/U$1 ( \55462 , \55461 , \40060 );
not \g132232/U$3 ( \55463 , \47948 );
and \g132285/U$2 ( \55464 , \47959 , \54853 );
and \g132285/U$3 ( \55465 , \55127 , \47960 );
nor \g132285/U$1 ( \55466 , \55464 , \55465 );
not \g132232/U$4 ( \55467 , \55466 );
or \g132232/U$2 ( \55468 , \55463 , \55467 );
or \g132232/U$5 ( \55469 , \55466 , \47948 );
nand \g132232/U$1 ( \55470 , \55468 , \55469 );
and \g132171/U$2 ( \55471 , \55462 , \55470 );
and \g132431/U$2 ( \55472 , \47913 , \54251 );
and \g132431/U$3 ( \55473 , \54529 , \47914 );
nor \g132431/U$1 ( \55474 , \55472 , \55473 );
and \g132351/U$2 ( \55475 , \55474 , \47977 );
not \g132351/U$4 ( \55476 , \55474 );
and \g132351/U$3 ( \55477 , \55476 , \47976 );
nor \g132351/U$1 ( \55478 , \55475 , \55477 );
xor \g132070/U$4 ( \55479 , \55471 , \55478 );
not \g132183/U$3 ( \55480 , \55128 );
not \g132183/U$4 ( \55481 , \55137 );
or \g132183/U$2 ( \55482 , \55480 , \55481 );
or \g132183/U$5 ( \55483 , \55137 , \55128 );
nand \g132183/U$1 ( \55484 , \55482 , \55483 );
and \g132070/U$3 ( \55485 , \55479 , \55484 );
and \g132070/U$5 ( \55486 , \55471 , \55478 );
or \g132070/U$2 ( \55487 , \55485 , \55486 );
and \g131981/U$3 ( \55488 , \55459 , \55487 );
and \g131981/U$5 ( \55489 , \55450 , \55458 );
or \g131981/U$2 ( \55490 , \55488 , \55489 );
not \g130965/U$3 ( \55491 , \49925 );
and \g130992/U$2 ( \55492 , \49888 , \50160 );
and \g130992/U$3 ( \55493 , \50159 , \49714 );
nor \g130992/U$1 ( \55494 , \55492 , \55493 );
not \g130965/U$4 ( \55495 , \55494 );
or \g130965/U$2 ( \55496 , \55491 , \55495 );
or \g130965/U$5 ( \55497 , \55494 , \49925 );
nand \g130965/U$1 ( \55498 , \55496 , \55497 );
xor \g456084/U$4 ( \55499 , \55490 , \55498 );
not \g130742/U$3 ( \55500 , \50759 );
and \g130767/U$2 ( \55501 , \49102 , \51053 );
and \g130767/U$3 ( \55502 , \51055 , \49158 );
nor \g130767/U$1 ( \55503 , \55501 , \55502 );
not \g130742/U$4 ( \55504 , \55503 );
or \g130742/U$2 ( \55505 , \55500 , \55504 );
or \g130742/U$5 ( \55506 , \55503 , \50759 );
nand \g130742/U$1 ( \55507 , \55505 , \55506 );
and \g456084/U$3 ( \55508 , \55499 , \55507 );
and \g456084/U$5 ( \55509 , \55490 , \55498 );
nor \g456084/U$2 ( \55510 , \55508 , \55509 );
xor \g130349/U$4 ( \55511 , \55442 , \55510 );
not \g132116/U$3 ( \55512 , \54865 );
not \g132116/U$4 ( \55513 , \54841 );
or \g132116/U$2 ( \55514 , \55512 , \55513 );
or \g132116/U$5 ( \55515 , \54841 , \54865 );
nand \g132116/U$1 ( \55516 , \55514 , \55515 );
not \g132101/U$3 ( \55517 , \55516 );
not \g132101/U$4 ( \55518 , \54848 );
and \g132101/U$2 ( \55519 , \55517 , \55518 );
and \g132101/U$5 ( \55520 , \55516 , \54848 );
nor \g132101/U$1 ( \55521 , \55519 , \55520 );
not \g131830/U$3 ( \55522 , \54970 );
xor \g131952/U$1 ( \55523 , \54960 , \54952 );
not \g131830/U$4 ( \55524 , \55523 );
and \g131830/U$2 ( \55525 , \55522 , \55524 );
and \g131830/U$5 ( \55526 , \54970 , \55523 );
nor \g131830/U$1 ( \55527 , \55525 , \55526 );
xor \g130427/U$4 ( \55528 , \55521 , \55527 );
and \g130524/U$2 ( \55529 , \48726 , \52273 );
and \g130524/U$3 ( \55530 , \52270 , \48568 );
nor \g130524/U$1 ( \55531 , \55529 , \55530 );
not \g130493/U$3 ( \55532 , \55531 );
not \g130493/U$4 ( \55533 , \51120 );
and \g130493/U$2 ( \55534 , \55532 , \55533 );
and \g130493/U$5 ( \55535 , \55531 , \51120 );
nor \g130493/U$1 ( \55536 , \55534 , \55535 );
and \g130427/U$3 ( \55537 , \55528 , \55536 );
and \g130427/U$5 ( \55538 , \55521 , \55527 );
or \g130427/U$2 ( \55539 , \55537 , \55538 );
and \g130349/U$3 ( \55540 , \55511 , \55539 );
and \g130349/U$5 ( \55541 , \55442 , \55510 );
or \g130349/U$2 ( \55542 , \55540 , \55541 );
xor \g130632/U$1 ( \55543 , \54510 , \54540 );
xor \g130632/U$1_r1 ( \55544 , \55543 , \54549 );
xor \g131124/U$1 ( \55545 , \54836 , \54867 );
xor \g131124/U$1_r1 ( \55546 , \55545 , \54876 );
and \g130475/U$2 ( \55547 , \55544 , \55546 );
not \g130477/U$3 ( \55548 , \55544 );
not \g130477/U$4 ( \55549 , \55546 );
and \g130477/U$2 ( \55550 , \55548 , \55549 );
xor \g130501/U$1 ( \55551 , \54909 , \54917 );
xor \g130501/U$1_r1 ( \55552 , \55551 , \54926 );
nor \g130477/U$1 ( \55553 , \55550 , \55552 );
nor \g130475/U$1 ( \55554 , \55547 , \55553 );
xor \g130222/U$4 ( \55555 , \55542 , \55554 );
not \g130322/U$3 ( \55556 , \54985 );
not \g130322/U$4 ( \55557 , \54929 );
and \g130322/U$2 ( \55558 , \55556 , \55557 );
and \g130322/U$5 ( \55559 , \54985 , \54929 );
nor \g130322/U$1 ( \55560 , \55558 , \55559 );
not \g130293/U$3 ( \55561 , \55560 );
not \g130293/U$4 ( \55562 , \54931 );
and \g130293/U$2 ( \55563 , \55561 , \55562 );
and \g130293/U$5 ( \55564 , \55560 , \54931 );
nor \g130293/U$1 ( \55565 , \55563 , \55564 );
and \g130222/U$3 ( \55566 , \55555 , \55565 );
and \g130222/U$5 ( \55567 , \55542 , \55554 );
or \g130222/U$2 ( \55568 , \55566 , \55567 );
or \g130051/U$2 ( \55569 , \55414 , \55568 );
and \g130054/U$2 ( \55570 , \55414 , \55568 );
not \g130147/U$3 ( \55571 , \54767 );
not \g130147/U$4 ( \55572 , \54639 );
and \g130147/U$2 ( \55573 , \55571 , \55572 );
and \g130147/U$5 ( \55574 , \54767 , \54639 );
nor \g130147/U$1 ( \55575 , \55573 , \55574 );
not \g130129/U$3 ( \55576 , \55575 );
not \g130129/U$4 ( \55577 , \54726 );
and \g130129/U$2 ( \55578 , \55576 , \55577 );
and \g130129/U$5 ( \55579 , \55575 , \54726 );
nor \g130129/U$1 ( \55580 , \55578 , \55579 );
nor \g130054/U$1 ( \55581 , \55570 , \55580 );
not \g130053/U$1 ( \55582 , \55581 );
nand \g130051/U$1 ( \55583 , \55569 , \55582 );
and \g456030/U$3 ( \55584 , \55283 , \55583 );
and \g456030/U$5 ( \55585 , \55001 , \55282 );
nor \g456030/U$2 ( \55586 , \55584 , \55585 );
xor \g456030/U$1 ( \55587 , \55001 , \55282 );
xor \g456030/U$1_r1 ( \55588 , \55587 , \55583 );
not \g130090/U$3 ( \55589 , \55208 );
xor \g130132/U$1 ( \55590 , \55174 , \55094 );
not \g130090/U$4 ( \55591 , \55590 );
and \g130090/U$2 ( \55592 , \55589 , \55591 );
and \g130090/U$5 ( \55593 , \55208 , \55590 );
nor \g130090/U$1 ( \55594 , \55592 , \55593 );
xor \g456084/U$1 ( \55595 , \55490 , \55498 );
xor \g456084/U$1_r1 ( \55596 , \55595 , \55507 );
not \g130695/U$1 ( \55597 , \55596 );
xnor \g455955/U$1 ( \55598 , \55389 , \55360 );
not \g131057/U$3 ( \55599 , \55598 );
not \g131057/U$4 ( \55600 , \55311 );
and \g131057/U$2 ( \55601 , \55599 , \55600 );
and \g131057/U$5 ( \55602 , \55598 , \55311 );
nor \g131057/U$1 ( \55603 , \55601 , \55602 );
or \g130541/U$2 ( \55604 , \55597 , \55603 );
not \g130545/U$3 ( \55605 , \55603 );
not \g130545/U$4 ( \55606 , \55597 );
or \g130545/U$2 ( \55607 , \55605 , \55606 );
xor \g456078/U$1 ( \55608 , \55422 , \55430 );
xor \g456078/U$1_r1 ( \55609 , \55608 , \55439 );
nand \g130545/U$1 ( \55610 , \55607 , \55609 );
nand \g130541/U$1 ( \55611 , \55604 , \55610 );
not \g130430/U$3 ( \55612 , \55546 );
not \g130471/U$3 ( \55613 , \55552 );
not \g130471/U$4 ( \55614 , \55544 );
and \g130471/U$2 ( \55615 , \55613 , \55614 );
and \g130471/U$5 ( \55616 , \55552 , \55544 );
nor \g130471/U$1 ( \55617 , \55615 , \55616 );
not \g130430/U$4 ( \55618 , \55617 );
or \g130430/U$2 ( \55619 , \55612 , \55618 );
or \g130430/U$5 ( \55620 , \55617 , \55546 );
nand \g130430/U$1 ( \55621 , \55619 , \55620 );
xor \g456060/U$4 ( \55622 , \55611 , \55621 );
xor \g456061/U$1 ( \55623 , \55391 , \55397 );
xor \g456061/U$1_r1 ( \55624 , \55623 , \55400 );
and \g456060/U$3 ( \55625 , \55622 , \55624 );
and \g456060/U$5 ( \55626 , \55611 , \55621 );
nor \g456060/U$2 ( \55627 , \55625 , \55626 );
xor \g131497/U$1 ( \55628 , \55291 , \55299 );
xor \g131497/U$1_r1 ( \55629 , \55628 , \55308 );
not \g131606/U$3 ( \55630 , \48685 );
and \g131635/U$2 ( \55631 , \51604 , \48858 );
and \g131635/U$3 ( \55632 , \48860 , \51854 );
nor \g131635/U$1 ( \55633 , \55631 , \55632 );
not \g131606/U$4 ( \55634 , \55633 );
or \g131606/U$2 ( \55635 , \55630 , \55634 );
or \g131606/U$5 ( \55636 , \55633 , \48685 );
nand \g131606/U$1 ( \55637 , \55635 , \55636 );
xor \g132070/U$1 ( \55638 , \55471 , \55478 );
xor \g132070/U$1_r1 ( \55639 , \55638 , \55484 );
xor \g131429/U$4 ( \55640 , \55637 , \55639 );
not \g131488/U$3 ( \55641 , \49014 );
and \g131516/U$2 ( \55642 , \51564 , \49075 );
and \g131516/U$3 ( \55643 , \49074 , \51098 );
nor \g131516/U$1 ( \55644 , \55642 , \55643 );
not \g131488/U$4 ( \55645 , \55644 );
or \g131488/U$2 ( \55646 , \55641 , \55645 );
or \g131488/U$5 ( \55647 , \55644 , \49014 );
nand \g131488/U$1 ( \55648 , \55646 , \55647 );
and \g131429/U$3 ( \55649 , \55640 , \55648 );
and \g131429/U$5 ( \55650 , \55637 , \55639 );
or \g131429/U$2 ( \55651 , \55649 , \55650 );
xor \g456072/U$4 ( \55652 , \55629 , \55651 );
not \g130561/U$3 ( \55653 , \51120 );
and \g130590/U$2 ( \55654 , \48726 , \52270 );
and \g130590/U$3 ( \55655 , \52273 , \48833 );
nor \g130590/U$1 ( \55656 , \55654 , \55655 );
not \g130561/U$4 ( \55657 , \55656 );
or \g130561/U$2 ( \55658 , \55653 , \55657 );
or \g130561/U$5 ( \55659 , \55656 , \51120 );
nand \g130561/U$1 ( \55660 , \55658 , \55659 );
and \g456072/U$3 ( \55661 , \55652 , \55660 );
and \g456072/U$5 ( \55662 , \55629 , \55651 );
nor \g456072/U$2 ( \55663 , \55661 , \55662 );
and \g130937/U$2 ( \55664 , \49512 , \50587 );
and \g130937/U$3 ( \55665 , \50588 , \49714 );
nor \g130937/U$1 ( \55666 , \55664 , \55665 );
not \g130909/U$3 ( \55667 , \55666 );
not \g130909/U$4 ( \55668 , \50362 );
and \g130909/U$2 ( \55669 , \55667 , \55668 );
and \g130909/U$5 ( \55670 , \55666 , \50362 );
nor \g130909/U$1 ( \55671 , \55669 , \55670 );
and \g131072/U$2 ( \55672 , \49888 , \50159 );
and \g131072/U$3 ( \55673 , \50160 , \50019 );
nor \g131072/U$1 ( \55674 , \55672 , \55673 );
not \g131031/U$3 ( \55675 , \55674 );
not \g131031/U$4 ( \55676 , \49925 );
and \g131031/U$2 ( \55677 , \55675 , \55676 );
and \g131031/U$5 ( \55678 , \55674 , \49925 );
nor \g131031/U$1 ( \55679 , \55677 , \55678 );
xor \g130635/U$4 ( \55680 , \55671 , \55679 );
and \g130713/U$2 ( \55681 , \49102 , \51518 );
and \g130713/U$3 ( \55682 , \51517 , \48977 );
nor \g130713/U$1 ( \55683 , \55681 , \55682 );
not \g130688/U$3 ( \55684 , \55683 );
not \g130688/U$4 ( \55685 , \51124 );
and \g130688/U$2 ( \55686 , \55684 , \55685 );
and \g130688/U$5 ( \55687 , \55683 , \51124 );
nor \g130688/U$1 ( \55688 , \55686 , \55687 );
and \g130635/U$3 ( \55689 , \55680 , \55688 );
and \g130635/U$5 ( \55690 , \55671 , \55679 );
or \g130635/U$2 ( \55691 , \55689 , \55690 );
xor \g130351/U$4 ( \55692 , \55663 , \55691 );
xor \g130427/U$1 ( \55693 , \55521 , \55527 );
xor \g130427/U$1_r1 ( \55694 , \55693 , \55536 );
and \g130351/U$3 ( \55695 , \55692 , \55694 );
and \g130351/U$5 ( \55696 , \55663 , \55691 );
or \g130351/U$2 ( \55697 , \55695 , \55696 );
not \g131458/U$3 ( \55698 , \54507 );
xor \g131570/U$1 ( \55699 , \54497 , \54489 );
not \g131458/U$4 ( \55700 , \55699 );
and \g131458/U$2 ( \55701 , \55698 , \55700 );
and \g131458/U$5 ( \55702 , \54507 , \55699 );
nor \g131458/U$1 ( \55703 , \55701 , \55702 );
xor \g456081/U$9 ( \55704 , \55110 , \55140 );
xor \g456081/U$9_r1 ( \55705 , \55704 , \55149 );
and \g456081/U$8 ( \55706 , \55703 , \55705 );
xor \g133003/U$1 ( \55707 , \47265 , \46758 );
not \g135543/U$2 ( \55708 , \55707 );
nor \g135543/U$1 ( \55709 , \55708 , \40060 );
and \g132434/U$2 ( \55710 , \47914 , \54853 );
and \g132434/U$3 ( \55711 , \54537 , \47913 );
nor \g132434/U$1 ( \55712 , \55710 , \55711 );
and \g132354/U$2 ( \55713 , \55712 , \47977 );
not \g132354/U$4 ( \55714 , \55712 );
and \g132354/U$3 ( \55715 , \55714 , \47976 );
nor \g132354/U$1 ( \55716 , \55713 , \55715 );
and \g132290/U$2 ( \55717 , \55709 , \55716 );
and \g132427/U$2 ( \55718 , \47914 , \54537 );
and \g132427/U$3 ( \55719 , \54529 , \47913 );
nor \g132427/U$1 ( \55720 , \55718 , \55719 );
and \g132356/U$2 ( \55721 , \55720 , \47977 );
not \g132356/U$4 ( \55722 , \55720 );
and \g132356/U$3 ( \55723 , \55722 , \47976 );
nor \g132356/U$1 ( \55724 , \55721 , \55723 );
xor \g132071/U$4 ( \55725 , \55717 , \55724 );
xor \g132171/U$1 ( \55726 , \55462 , \55470 );
and \g132071/U$3 ( \55727 , \55725 , \55726 );
and \g132071/U$5 ( \55728 , \55717 , \55724 );
or \g132071/U$2 ( \55729 , \55727 , \55728 );
not \g131852/U$3 ( \55730 , \48323 );
and \g131898/U$2 ( \55731 , \52620 , \48334 );
and \g131898/U$3 ( \55732 , \48335 , \52883 );
nor \g131898/U$1 ( \55733 , \55731 , \55732 );
not \g131852/U$4 ( \55734 , \55733 );
or \g131852/U$2 ( \55735 , \55730 , \55734 );
or \g131852/U$5 ( \55736 , \55733 , \48323 );
nand \g131852/U$1 ( \55737 , \55735 , \55736 );
xor \g131667/U$4 ( \55738 , \55729 , \55737 );
not \g131733/U$3 ( \55739 , \48483 );
and \g131764/U$2 ( \55740 , \52108 , \48478 );
and \g131764/U$3 ( \55741 , \48479 , \52352 );
nor \g131764/U$1 ( \55742 , \55740 , \55741 );
not \g131733/U$4 ( \55743 , \55742 );
or \g131733/U$2 ( \55744 , \55739 , \55743 );
or \g131733/U$5 ( \55745 , \55742 , \48483 );
nand \g131733/U$1 ( \55746 , \55744 , \55745 );
and \g131667/U$3 ( \55747 , \55738 , \55746 );
and \g131667/U$5 ( \55748 , \55729 , \55737 );
or \g131667/U$2 ( \55749 , \55747 , \55748 );
xor \g131981/U$1 ( \55750 , \55450 , \55458 );
xor \g131981/U$1_r1 ( \55751 , \55750 , \55487 );
xor \g456085/U$4 ( \55752 , \55749 , \55751 );
not \g130798/U$3 ( \55753 , \50759 );
and \g130825/U$2 ( \55754 , \49282 , \51055 );
and \g130825/U$3 ( \55755 , \51053 , \49158 );
nor \g130825/U$1 ( \55756 , \55754 , \55755 );
not \g130798/U$4 ( \55757 , \55756 );
or \g130798/U$2 ( \55758 , \55753 , \55757 );
or \g130798/U$5 ( \55759 , \55756 , \50759 );
nand \g130798/U$1 ( \55760 , \55758 , \55759 );
and \g456085/U$3 ( \55761 , \55752 , \55760 );
and \g456085/U$5 ( \55762 , \55749 , \55751 );
nor \g456085/U$2 ( \55763 , \55761 , \55762 );
xor \g456081/U$11 ( \55764 , \55110 , \55140 );
xor \g456081/U$11_r1 ( \55765 , \55764 , \55149 );
and \g456081/U$10 ( \55766 , \55763 , \55765 );
and \g456081/U$12 ( \55767 , \55703 , \55763 );
or \g456081/U$7 ( \55768 , \55706 , \55766 , \55767 );
xor \g130258/U$4 ( \55769 , \55697 , \55768 );
xor \g130349/U$1 ( \55770 , \55442 , \55510 );
xor \g130349/U$1_r1 ( \55771 , \55770 , \55539 );
and \g130258/U$3 ( \55772 , \55769 , \55771 );
and \g130258/U$5 ( \55773 , \55697 , \55768 );
or \g130258/U$2 ( \55774 , \55772 , \55773 );
xor \g130137/U$4 ( \55775 , \55627 , \55774 );
xor \g130222/U$1 ( \55776 , \55542 , \55554 );
xor \g130222/U$1_r1 ( \55777 , \55776 , \55565 );
and \g130137/U$3 ( \55778 , \55775 , \55777 );
and \g130137/U$5 ( \55779 , \55627 , \55774 );
or \g130137/U$2 ( \55780 , \55778 , \55779 );
or \g129943/U$2 ( \55781 , \55594 , \55780 );
and \g129948/U$2 ( \55782 , \55594 , \55780 );
not \g130042/U$3 ( \55783 , \55413 );
not \g130042/U$4 ( \55784 , \55580 );
or \g130042/U$2 ( \55785 , \55783 , \55784 );
or \g130042/U$5 ( \55786 , \55580 , \55413 );
nand \g130042/U$1 ( \55787 , \55785 , \55786 );
not \g130015/U$3 ( \55788 , \55787 );
not \g130015/U$4 ( \55789 , \55568 );
and \g130015/U$2 ( \55790 , \55788 , \55789 );
and \g130015/U$5 ( \55791 , \55787 , \55568 );
nor \g130015/U$1 ( \55792 , \55790 , \55791 );
nor \g129948/U$1 ( \55793 , \55782 , \55792 );
not \g129947/U$1 ( \55794 , \55793 );
nand \g129943/U$1 ( \55795 , \55781 , \55794 );
not \g130199/U$3 ( \55796 , \55403 );
not \g130199/U$4 ( \55797 , \55411 );
or \g130199/U$2 ( \55798 , \55796 , \55797 );
or \g130199/U$5 ( \55799 , \55411 , \55403 );
nand \g130199/U$1 ( \55800 , \55798 , \55799 );
not \g130168/U$3 ( \55801 , \55800 );
not \g130168/U$4 ( \55802 , \55405 );
and \g130168/U$2 ( \55803 , \55801 , \55802 );
and \g130168/U$5 ( \55804 , \55800 , \55405 );
nor \g130168/U$1 ( \55805 , \55803 , \55804 );
not \g130052/U$3 ( \55806 , \55805 );
xor \g130635/U$1 ( \55807 , \55671 , \55679 );
xor \g130635/U$1_r1 ( \55808 , \55807 , \55688 );
xor \g131667/U$1 ( \55809 , \55729 , \55737 );
xor \g131667/U$1_r1 ( \55810 , \55809 , \55746 );
not \g131665/U$3 ( \55811 , \48685 );
and \g131697/U$2 ( \55812 , \52108 , \48860 );
and \g131697/U$3 ( \55813 , \48858 , \51854 );
nor \g131697/U$1 ( \55814 , \55812 , \55813 );
not \g131665/U$4 ( \55815 , \55814 );
or \g131665/U$2 ( \55816 , \55811 , \55815 );
or \g131665/U$5 ( \55817 , \55814 , \48685 );
nand \g131665/U$1 ( \55818 , \55816 , \55817 );
xor \g132071/U$1 ( \55819 , \55717 , \55724 );
xor \g132071/U$1_r1 ( \55820 , \55819 , \55726 );
xor \g131498/U$4 ( \55821 , \55818 , \55820 );
not \g131554/U$3 ( \55822 , \49014 );
and \g131584/U$2 ( \55823 , \51604 , \49075 );
and \g131584/U$3 ( \55824 , \49074 , \51564 );
nor \g131584/U$1 ( \55825 , \55823 , \55824 );
not \g131554/U$4 ( \55826 , \55825 );
or \g131554/U$2 ( \55827 , \55822 , \55826 );
or \g131554/U$5 ( \55828 , \55825 , \49014 );
nand \g131554/U$1 ( \55829 , \55827 , \55828 );
and \g131498/U$3 ( \55830 , \55821 , \55829 );
and \g131498/U$5 ( \55831 , \55818 , \55820 );
or \g131498/U$2 ( \55832 , \55830 , \55831 );
xor \g456088/U$4 ( \55833 , \55810 , \55832 );
not \g130855/U$3 ( \55834 , \50759 );
and \g130879/U$2 ( \55835 , \49512 , \51055 );
and \g130879/U$3 ( \55836 , \51053 , \49282 );
nor \g130879/U$1 ( \55837 , \55835 , \55836 );
not \g130855/U$4 ( \55838 , \55837 );
or \g130855/U$2 ( \55839 , \55834 , \55838 );
or \g130855/U$5 ( \55840 , \55837 , \50759 );
nand \g130855/U$1 ( \55841 , \55839 , \55840 );
and \g456088/U$3 ( \55842 , \55833 , \55841 );
and \g456088/U$5 ( \55843 , \55810 , \55832 );
nor \g456088/U$2 ( \55844 , \55842 , \55843 );
or \g130474/U$2 ( \55845 , \55808 , \55844 );
not \g130476/U$3 ( \55846 , \55844 );
not \g130476/U$4 ( \55847 , \55808 );
or \g130476/U$2 ( \55848 , \55846 , \55847 );
xor \g456072/U$1 ( \55849 , \55629 , \55651 );
xor \g456072/U$1_r1 ( \55850 , \55849 , \55660 );
nand \g130476/U$1 ( \55851 , \55848 , \55850 );
nand \g130474/U$1 ( \55852 , \55845 , \55851 );
not \g130536/U$3 ( \55853 , \55609 );
not \g130536/U$4 ( \55854 , \55603 );
and \g130536/U$2 ( \55855 , \55853 , \55854 );
and \g130536/U$5 ( \55856 , \55609 , \55603 );
nor \g130536/U$1 ( \55857 , \55855 , \55856 );
not \g130504/U$3 ( \55858 , \55857 );
not \g130504/U$4 ( \55859 , \55596 );
and \g130504/U$2 ( \55860 , \55858 , \55859 );
and \g130504/U$5 ( \55861 , \55857 , \55596 );
nor \g130504/U$1 ( \55862 , \55860 , \55861 );
not \g130495/U$1 ( \55863 , \55862 );
and \g130315/U$2 ( \55864 , \55852 , \55863 );
not \g130318/U$3 ( \55865 , \55852 );
not \g130318/U$4 ( \55866 , \55863 );
and \g130318/U$2 ( \55867 , \55865 , \55866 );
xor \g130351/U$1 ( \55868 , \55663 , \55691 );
xor \g130351/U$1_r1 ( \55869 , \55868 , \55694 );
nor \g130318/U$1 ( \55870 , \55867 , \55869 );
nor \g130315/U$1 ( \55871 , \55864 , \55870 );
not \g130207/U$3 ( \55872 , \55871 );
xor \g456085/U$1 ( \55873 , \55749 , \55751 );
xor \g456085/U$1_r1 ( \55874 , \55873 , \55760 );
xor \g131367/U$1 ( \55875 , \55320 , \55348 );
xor \g131367/U$1_r1 ( \55876 , \55875 , \55357 );
and \g130670/U$2 ( \55877 , \55874 , \55876 );
not \g130672/U$3 ( \55878 , \55874 );
not \g130672/U$4 ( \55879 , \55876 );
and \g130672/U$2 ( \55880 , \55878 , \55879 );
xor \g131948/U$1 ( \55881 , \55328 , \55336 );
xor \g131948/U$1_r1 ( \55882 , \55881 , \55345 );
xor \g132290/U$1 ( \55883 , \55709 , \55716 );
xor \g133054/U$1 ( \55884 , \47262 , \47251 );
not \g135545/U$2 ( \55885 , \55884 );
nor \g135545/U$1 ( \55886 , \55885 , \40060 );
and \g132426/U$2 ( \55887 , \47913 , \54853 );
and \g132426/U$3 ( \55888 , \55127 , \47914 );
nor \g132426/U$1 ( \55889 , \55887 , \55888 );
and \g132355/U$2 ( \55890 , \55889 , \47977 );
not \g132355/U$4 ( \55891 , \55889 );
and \g132355/U$3 ( \55892 , \55891 , \47976 );
nor \g132355/U$1 ( \55893 , \55890 , \55892 );
and \g132292/U$2 ( \55894 , \55886 , \55893 );
xor \g132145/U$4 ( \55895 , \55883 , \55894 );
not \g132233/U$3 ( \55896 , \47948 );
and \g132286/U$2 ( \55897 , \47959 , \55127 );
and \g132286/U$3 ( \55898 , \55460 , \47960 );
nor \g132286/U$1 ( \55899 , \55897 , \55898 );
not \g132233/U$4 ( \55900 , \55899 );
or \g132233/U$2 ( \55901 , \55896 , \55900 );
or \g132233/U$5 ( \55902 , \55899 , \47948 );
nand \g132233/U$1 ( \55903 , \55901 , \55902 );
and \g132145/U$3 ( \55904 , \55895 , \55903 );
and \g132145/U$5 ( \55905 , \55883 , \55894 );
or \g132145/U$2 ( \55906 , \55904 , \55905 );
not \g131932/U$3 ( \55907 , \48323 );
and \g131966/U$2 ( \55908 , \52978 , \48335 );
and \g131966/U$3 ( \55909 , \48334 , \52883 );
nor \g131966/U$1 ( \55910 , \55908 , \55909 );
not \g131932/U$4 ( \55911 , \55910 );
or \g131932/U$2 ( \55912 , \55907 , \55911 );
or \g131932/U$5 ( \55913 , \55910 , \48323 );
nand \g131932/U$1 ( \55914 , \55912 , \55913 );
xor \g131741/U$4 ( \55915 , \55906 , \55914 );
not \g131793/U$3 ( \55916 , \48483 );
and \g131824/U$2 ( \55917 , \52620 , \48479 );
and \g131824/U$3 ( \55918 , \48478 , \52352 );
nor \g131824/U$1 ( \55919 , \55917 , \55918 );
not \g131793/U$4 ( \55920 , \55919 );
or \g131793/U$2 ( \55921 , \55916 , \55920 );
or \g131793/U$5 ( \55922 , \55919 , \48483 );
nand \g131793/U$1 ( \55923 , \55921 , \55922 );
and \g131741/U$3 ( \55924 , \55915 , \55923 );
and \g131741/U$5 ( \55925 , \55906 , \55914 );
or \g131741/U$2 ( \55926 , \55924 , \55925 );
xor \g456083/U$4 ( \55927 , \55882 , \55926 );
not \g130743/U$3 ( \55928 , \51124 );
and \g130768/U$2 ( \55929 , \49102 , \51517 );
and \g130768/U$3 ( \55930 , \51518 , \49158 );
nor \g130768/U$1 ( \55931 , \55929 , \55930 );
not \g130743/U$4 ( \55932 , \55931 );
or \g130743/U$2 ( \55933 , \55928 , \55932 );
or \g130743/U$5 ( \55934 , \55931 , \51124 );
nand \g130743/U$1 ( \55935 , \55933 , \55934 );
and \g456083/U$3 ( \55936 , \55927 , \55935 );
and \g456083/U$5 ( \55937 , \55882 , \55926 );
nor \g456083/U$2 ( \55938 , \55936 , \55937 );
nor \g130672/U$1 ( \55939 , \55880 , \55938 );
nor \g130670/U$1 ( \55940 , \55877 , \55939 );
not \g130496/U$3 ( \55941 , \55940 );
xor \g456081/U$2 ( \55942 , \55110 , \55140 );
xor \g456081/U$1 ( \55943 , \55942 , \55149 );
xor \g456081/U$1_r1 ( \55944 , \55703 , \55763 );
xor \g456081/U$1_r2 ( \55945 , \55943 , \55944 );
not \g130496/U$4 ( \55946 , \55945 );
and \g130496/U$2 ( \55947 , \55941 , \55946 );
and \g130497/U$2 ( \55948 , \55940 , \55945 );
not \g131242/U$3 ( \55949 , \49568 );
and \g131274/U$2 ( \55950 , \50752 , \49813 );
and \g131274/U$3 ( \55951 , \49812 , \50443 );
nor \g131274/U$1 ( \55952 , \55950 , \55951 );
not \g131242/U$4 ( \55953 , \55952 );
or \g131242/U$2 ( \55954 , \55949 , \55953 );
or \g131242/U$5 ( \55955 , \55952 , \49568 );
nand \g131242/U$1 ( \55956 , \55954 , \55955 );
not \g132458/U$3 ( \55957 , \47935 );
and \g132502/U$2 ( \55958 , \47930 , \54185 );
and \g132502/U$3 ( \55959 , \54251 , \47931 );
nor \g132502/U$1 ( \55960 , \55958 , \55959 );
not \g132458/U$4 ( \55961 , \55960 );
or \g132458/U$2 ( \55962 , \55957 , \55961 );
or \g132458/U$5 ( \55963 , \55960 , \47935 );
nand \g132458/U$1 ( \55964 , \55962 , \55963 );
not \g132257/U$3 ( \55965 , \47997 );
and \g132306/U$2 ( \55966 , \53848 , \48063 );
and \g132306/U$3 ( \55967 , \54015 , \48064 );
nor \g132306/U$1 ( \55968 , \55966 , \55967 );
not \g132257/U$4 ( \55969 , \55968 );
or \g132257/U$2 ( \55970 , \55965 , \55969 );
or \g132257/U$5 ( \55971 , \55968 , \47997 );
nand \g132257/U$1 ( \55972 , \55970 , \55971 );
xor \g132030/U$4 ( \55973 , \55964 , \55972 );
not \g132092/U$3 ( \55974 , \48159 );
and \g132132/U$2 ( \55975 , \53610 , \48155 );
and \g132132/U$3 ( \55976 , \48154 , \53300 );
nor \g132132/U$1 ( \55977 , \55975 , \55976 );
not \g132092/U$4 ( \55978 , \55977 );
or \g132092/U$2 ( \55979 , \55974 , \55978 );
or \g132092/U$5 ( \55980 , \55977 , \48159 );
nand \g132092/U$1 ( \55981 , \55979 , \55980 );
and \g132030/U$3 ( \55982 , \55973 , \55981 );
and \g132030/U$5 ( \55983 , \55964 , \55972 );
or \g132030/U$2 ( \55984 , \55982 , \55983 );
xor \g131051/U$4 ( \55985 , \55956 , \55984 );
not \g131113/U$3 ( \55986 , \49925 );
and \g131147/U$2 ( \55987 , \50305 , \50160 );
and \g131147/U$3 ( \55988 , \50159 , \50019 );
nor \g131147/U$1 ( \55989 , \55987 , \55988 );
not \g131113/U$4 ( \55990 , \55989 );
or \g131113/U$2 ( \55991 , \55986 , \55990 );
or \g131113/U$5 ( \55992 , \55989 , \49925 );
nand \g131113/U$1 ( \55993 , \55991 , \55992 );
and \g131051/U$3 ( \55994 , \55985 , \55993 );
and \g131051/U$5 ( \55995 , \55956 , \55984 );
or \g131051/U$2 ( \55996 , \55994 , \55995 );
xor \g131126/U$1 ( \55997 , \55371 , \55377 );
xor \g131126/U$1_r1 ( \55998 , \55997 , \55386 );
xor \g130526/U$4 ( \55999 , \55996 , \55998 );
and \g130993/U$2 ( \56000 , \49888 , \50588 );
and \g130993/U$3 ( \56001 , \50587 , \49714 );
nor \g130993/U$1 ( \56002 , \56000 , \56001 );
not \g130966/U$3 ( \56003 , \56002 );
not \g130966/U$4 ( \56004 , \50362 );
and \g130966/U$2 ( \56005 , \56003 , \56004 );
and \g130966/U$5 ( \56006 , \56002 , \50362 );
nor \g130966/U$1 ( \56007 , \56005 , \56006 );
and \g131382/U$2 ( \56008 , \51117 , \49405 );
and \g131382/U$3 ( \56009 , \49403 , \50957 );
nor \g131382/U$1 ( \56010 , \56008 , \56009 );
not \g131361/U$3 ( \56011 , \56010 );
not \g131361/U$4 ( \56012 , \49233 );
and \g131361/U$2 ( \56013 , \56011 , \56012 );
and \g131361/U$5 ( \56014 , \56010 , \49233 );
nor \g131361/U$1 ( \56015 , \56013 , \56014 );
or \g130594/U$2 ( \56016 , \56007 , \56015 );
and \g130602/U$2 ( \56017 , \56007 , \56015 );
and \g130658/U$2 ( \56018 , \48833 , \52270 );
and \g130658/U$3 ( \56019 , \52273 , \48977 );
nor \g130658/U$1 ( \56020 , \56018 , \56019 );
not \g130624/U$3 ( \56021 , \56020 );
not \g130624/U$4 ( \56022 , \51120 );
and \g130624/U$2 ( \56023 , \56021 , \56022 );
and \g130624/U$5 ( \56024 , \56020 , \51120 );
nor \g130624/U$1 ( \56025 , \56023 , \56024 );
nor \g130602/U$1 ( \56026 , \56017 , \56025 );
not \g130601/U$1 ( \56027 , \56026 );
nand \g130594/U$1 ( \56028 , \56016 , \56027 );
and \g130526/U$3 ( \56029 , \55999 , \56028 );
and \g130526/U$5 ( \56030 , \55996 , \55998 );
or \g130526/U$2 ( \56031 , \56029 , \56030 );
not \g130525/U$1 ( \56032 , \56031 );
nor \g130497/U$1 ( \56033 , \55948 , \56032 );
nor \g130496/U$1 ( \56034 , \55947 , \56033 );
not \g130207/U$4 ( \56035 , \56034 );
and \g130207/U$2 ( \56036 , \55872 , \56035 );
and \g130210/U$2 ( \56037 , \55871 , \56034 );
xor \g130258/U$1 ( \56038 , \55697 , \55768 );
xor \g130258/U$1_r1 ( \56039 , \56038 , \55771 );
nor \g130210/U$1 ( \56040 , \56037 , \56039 );
nor \g130207/U$1 ( \56041 , \56036 , \56040 );
xor \g130137/U$1 ( \56042 , \55627 , \55774 );
xor \g130137/U$1_r1 ( \56043 , \56042 , \55777 );
xor \g130106/U$1 ( \56044 , \56041 , \56043 );
not \g130052/U$4 ( \56045 , \56044 );
or \g130052/U$2 ( \56046 , \55806 , \56045 );
or \g130052/U$5 ( \56047 , \56044 , \55805 );
nand \g130052/U$1 ( \56048 , \56046 , \56047 );
xor \g456060/U$1 ( \56049 , \55611 , \55621 );
xor \g456060/U$1_r1 ( \56050 , \56049 , \55624 );
not \g130257/U$1 ( \56051 , \56050 );
not \g130459/U$3 ( \56052 , \55945 );
not \g130494/U$3 ( \56053 , \55940 );
not \g130494/U$4 ( \56054 , \56031 );
or \g130494/U$2 ( \56055 , \56053 , \56054 );
or \g130494/U$5 ( \56056 , \56031 , \55940 );
nand \g130494/U$1 ( \56057 , \56055 , \56056 );
not \g130459/U$4 ( \56058 , \56057 );
or \g130459/U$2 ( \56059 , \56052 , \56058 );
or \g130459/U$5 ( \56060 , \56057 , \55945 );
nand \g130459/U$1 ( \56061 , \56059 , \56060 );
not \g130637/U$3 ( \56062 , \55876 );
not \g130667/U$3 ( \56063 , \55938 );
not \g130667/U$4 ( \56064 , \55874 );
and \g130667/U$2 ( \56065 , \56063 , \56064 );
and \g130667/U$5 ( \56066 , \55938 , \55874 );
nor \g130667/U$1 ( \56067 , \56065 , \56066 );
not \g130637/U$4 ( \56068 , \56067 );
or \g130637/U$2 ( \56069 , \56062 , \56068 );
or \g130637/U$5 ( \56070 , \56067 , \55876 );
nand \g130637/U$1 ( \56071 , \56069 , \56070 );
not \g131303/U$3 ( \56072 , \49568 );
and \g131327/U$2 ( \56073 , \50957 , \49813 );
and \g131327/U$3 ( \56074 , \49812 , \50752 );
nor \g131327/U$1 ( \56075 , \56073 , \56074 );
not \g131303/U$4 ( \56076 , \56075 );
or \g131303/U$2 ( \56077 , \56072 , \56076 );
or \g131303/U$5 ( \56078 , \56075 , \49568 );
nand \g131303/U$1 ( \56079 , \56077 , \56078 );
not \g132490/U$3 ( \56080 , \47935 );
and \g132555/U$2 ( \56081 , \47930 , \54251 );
and \g132555/U$3 ( \56082 , \54529 , \47931 );
nor \g132555/U$1 ( \56083 , \56081 , \56082 );
not \g132490/U$4 ( \56084 , \56083 );
or \g132490/U$2 ( \56085 , \56080 , \56084 );
or \g132490/U$5 ( \56086 , \56083 , \47935 );
nand \g132490/U$1 ( \56087 , \56085 , \56086 );
not \g132357/U$3 ( \56088 , \47997 );
and \g132417/U$2 ( \56089 , \48064 , \54185 );
and \g132417/U$3 ( \56090 , \48063 , \54015 );
nor \g132417/U$1 ( \56091 , \56089 , \56090 );
not \g132357/U$4 ( \56092 , \56091 );
or \g132357/U$2 ( \56093 , \56088 , \56092 );
or \g132357/U$5 ( \56094 , \56091 , \47997 );
nand \g132357/U$1 ( \56095 , \56093 , \56094 );
xor \g132099/U$4 ( \56096 , \56087 , \56095 );
not \g132161/U$3 ( \56097 , \48159 );
and \g132205/U$2 ( \56098 , \53610 , \48154 );
and \g132205/U$3 ( \56099 , \48155 , \53848 );
nor \g132205/U$1 ( \56100 , \56098 , \56099 );
not \g132161/U$4 ( \56101 , \56100 );
or \g132161/U$2 ( \56102 , \56097 , \56101 );
or \g132161/U$5 ( \56103 , \56100 , \48159 );
nand \g132161/U$1 ( \56104 , \56102 , \56103 );
and \g132099/U$3 ( \56105 , \56096 , \56104 );
and \g132099/U$5 ( \56106 , \56087 , \56095 );
or \g132099/U$2 ( \56107 , \56105 , \56106 );
xor \g131127/U$4 ( \56108 , \56079 , \56107 );
not \g131189/U$3 ( \56109 , \49925 );
and \g131219/U$2 ( \56110 , \50305 , \50159 );
and \g131219/U$3 ( \56111 , \50160 , \50443 );
nor \g131219/U$1 ( \56112 , \56110 , \56111 );
not \g131189/U$4 ( \56113 , \56112 );
or \g131189/U$2 ( \56114 , \56109 , \56113 );
or \g131189/U$5 ( \56115 , \56112 , \49925 );
nand \g131189/U$1 ( \56116 , \56114 , \56115 );
and \g131127/U$3 ( \56117 , \56108 , \56116 );
and \g131127/U$5 ( \56118 , \56079 , \56107 );
or \g131127/U$2 ( \56119 , \56117 , \56118 );
xor \g131429/U$1 ( \56120 , \55637 , \55639 );
xor \g131429/U$1_r1 ( \56121 , \56120 , \55648 );
xor \g130971/U$4 ( \56122 , \56119 , \56121 );
xor \g131051/U$1 ( \56123 , \55956 , \55984 );
xor \g131051/U$1_r1 ( \56124 , \56123 , \55993 );
and \g130971/U$3 ( \56125 , \56122 , \56124 );
and \g130971/U$5 ( \56126 , \56119 , \56121 );
or \g130971/U$2 ( \56127 , \56125 , \56126 );
xor \g130473/U$4 ( \56128 , \56071 , \56127 );
xor \g130526/U$1 ( \56129 , \55996 , \55998 );
xor \g130526/U$1_r1 ( \56130 , \56129 , \56028 );
and \g130473/U$3 ( \56131 , \56128 , \56130 );
and \g130473/U$5 ( \56132 , \56071 , \56127 );
or \g130473/U$2 ( \56133 , \56131 , \56132 );
and \g130291/U$2 ( \56134 , \56061 , \56133 );
not \g130294/U$3 ( \56135 , \56061 );
not \g130294/U$4 ( \56136 , \56133 );
and \g130294/U$2 ( \56137 , \56135 , \56136 );
xor \g456083/U$1 ( \56138 , \55882 , \55926 );
xor \g456083/U$1_r1 ( \56139 , \56138 , \55935 );
xor \g456088/U$1 ( \56140 , \55810 , \55832 );
xor \g456088/U$1_r1 ( \56141 , \56140 , \55841 );
and \g130540/U$2 ( \56142 , \56139 , \56141 );
not \g130544/U$3 ( \56143 , \56139 );
not \g130544/U$4 ( \56144 , \56141 );
and \g130544/U$2 ( \56145 , \56143 , \56144 );
not \g130595/U$3 ( \56146 , \56025 );
xor \g130921/U$1 ( \56147 , \56015 , \56007 );
not \g130595/U$4 ( \56148 , \56147 );
and \g130595/U$2 ( \56149 , \56146 , \56148 );
and \g130595/U$5 ( \56150 , \56025 , \56147 );
nor \g130595/U$1 ( \56151 , \56149 , \56150 );
nor \g130544/U$1 ( \56152 , \56145 , \56151 );
nor \g130540/U$1 ( \56153 , \56142 , \56152 );
not \g130390/U$3 ( \56154 , \56153 );
xor \g132030/U$1 ( \56155 , \55964 , \55972 );
xor \g132030/U$1_r1 ( \56156 , \56155 , \55981 );
not \g132234/U$3 ( \56157 , \47948 );
and \g132287/U$2 ( \56158 , \47959 , \55460 );
and \g132287/U$3 ( \56159 , \55707 , \47960 );
nor \g132287/U$1 ( \56160 , \56158 , \56159 );
not \g132234/U$4 ( \56161 , \56160 );
or \g132234/U$2 ( \56162 , \56157 , \56161 );
or \g132234/U$5 ( \56163 , \56160 , \47948 );
nand \g132234/U$1 ( \56164 , \56162 , \56163 );
xor \g132292/U$1 ( \56165 , \55886 , \55893 );
xor \g456134/U$5 ( \56166 , \56164 , \56165 );
xor \g133111/U$1 ( \56167 , \46881 , \47249 );
not \g135547/U$2 ( \56168 , \56167 );
nor \g135547/U$1 ( \56169 , \56168 , \40060 );
not \g132235/U$3 ( \56170 , \47948 );
and \g132288/U$2 ( \56171 , \47960 , \55884 );
and \g132288/U$3 ( \56172 , \55707 , \47959 );
nor \g132288/U$1 ( \56173 , \56171 , \56172 );
not \g132235/U$4 ( \56174 , \56173 );
or \g132235/U$2 ( \56175 , \56170 , \56174 );
or \g132235/U$5 ( \56176 , \56173 , \47948 );
nand \g132235/U$1 ( \56177 , \56175 , \56176 );
and \g132172/U$2 ( \56178 , \56169 , \56177 );
and \g456134/U$4 ( \56179 , \56166 , \56178 );
and \g456134/U$6 ( \56180 , \56164 , \56165 );
or \g456134/U$3 ( \56181 , \56179 , \56180 );
not \g132014/U$3 ( \56182 , \48323 );
and \g132052/U$2 ( \56183 , \52978 , \48334 );
and \g132052/U$3 ( \56184 , \48335 , \53300 );
nor \g132052/U$1 ( \56185 , \56183 , \56184 );
not \g132014/U$4 ( \56186 , \56185 );
or \g132014/U$2 ( \56187 , \56182 , \56186 );
or \g132014/U$5 ( \56188 , \56185 , \48323 );
nand \g132014/U$1 ( \56189 , \56187 , \56188 );
xor \g131668/U$4 ( \56190 , \56181 , \56189 );
not \g131734/U$3 ( \56191 , \48685 );
and \g131765/U$2 ( \56192 , \52108 , \48858 );
and \g131765/U$3 ( \56193 , \48860 , \52352 );
nor \g131765/U$1 ( \56194 , \56192 , \56193 );
not \g131734/U$4 ( \56195 , \56194 );
or \g131734/U$2 ( \56196 , \56191 , \56195 );
or \g131734/U$5 ( \56197 , \56194 , \48685 );
nand \g131734/U$1 ( \56198 , \56196 , \56197 );
and \g131668/U$3 ( \56199 , \56190 , \56198 );
and \g131668/U$5 ( \56200 , \56181 , \56189 );
or \g131668/U$2 ( \56201 , \56199 , \56200 );
xor \g456073/U$5 ( \56202 , \56156 , \56201 );
not \g130799/U$3 ( \56203 , \51124 );
and \g130826/U$2 ( \56204 , \49282 , \51518 );
and \g130826/U$3 ( \56205 , \51517 , \49158 );
nor \g130826/U$1 ( \56206 , \56204 , \56205 );
not \g130799/U$4 ( \56207 , \56206 );
or \g130799/U$2 ( \56208 , \56203 , \56207 );
or \g130799/U$5 ( \56209 , \56206 , \51124 );
nand \g130799/U$1 ( \56210 , \56208 , \56209 );
and \g456073/U$4 ( \56211 , \56202 , \56210 );
and \g456073/U$6 ( \56212 , \56156 , \56201 );
or \g456073/U$3 ( \56213 , \56211 , \56212 );
not \g456074/U$1 ( \56214 , \56213 );
not \g130606/U$3 ( \56215 , \56214 );
xor \g131741/U$1 ( \56216 , \55906 , \55914 );
xor \g131741/U$1_r1 ( \56217 , \56216 , \55923 );
not \g131607/U$3 ( \56218 , \49014 );
and \g131636/U$2 ( \56219 , \51604 , \49074 );
and \g131636/U$3 ( \56220 , \49075 , \51854 );
nor \g131636/U$1 ( \56221 , \56219 , \56220 );
not \g131607/U$4 ( \56222 , \56221 );
or \g131607/U$2 ( \56223 , \56218 , \56222 );
or \g131607/U$5 ( \56224 , \56221 , \49014 );
nand \g131607/U$1 ( \56225 , \56223 , \56224 );
not \g131859/U$3 ( \56226 , \48483 );
and \g131900/U$2 ( \56227 , \52620 , \48478 );
and \g131900/U$3 ( \56228 , \48479 , \52883 );
nor \g131900/U$1 ( \56229 , \56227 , \56228 );
not \g131859/U$4 ( \56230 , \56229 );
or \g131859/U$2 ( \56231 , \56226 , \56230 );
or \g131859/U$5 ( \56232 , \56229 , \48483 );
nand \g131859/U$1 ( \56233 , \56231 , \56232 );
xor \g131428/U$4 ( \56234 , \56225 , \56233 );
not \g131489/U$3 ( \56235 , \49233 );
and \g131517/U$2 ( \56236 , \51564 , \49405 );
and \g131517/U$3 ( \56237 , \49403 , \51098 );
nor \g131517/U$1 ( \56238 , \56236 , \56237 );
not \g131489/U$4 ( \56239 , \56238 );
or \g131489/U$2 ( \56240 , \56235 , \56239 );
or \g131489/U$5 ( \56241 , \56238 , \49233 );
nand \g131489/U$1 ( \56242 , \56240 , \56241 );
and \g131428/U$3 ( \56243 , \56234 , \56242 );
and \g131428/U$5 ( \56244 , \56225 , \56233 );
or \g131428/U$2 ( \56245 , \56243 , \56244 );
xor \g456092/U$4 ( \56246 , \56217 , \56245 );
not \g130908/U$3 ( \56247 , \50759 );
and \g130936/U$2 ( \56248 , \49512 , \51053 );
and \g130936/U$3 ( \56249 , \51055 , \49714 );
nor \g130936/U$1 ( \56250 , \56248 , \56249 );
not \g130908/U$4 ( \56251 , \56250 );
or \g130908/U$2 ( \56252 , \56247 , \56251 );
or \g130908/U$5 ( \56253 , \56250 , \50759 );
nand \g130908/U$1 ( \56254 , \56252 , \56253 );
and \g456092/U$3 ( \56255 , \56246 , \56254 );
and \g456092/U$5 ( \56256 , \56217 , \56245 );
nor \g456092/U$2 ( \56257 , \56255 , \56256 );
not \g130606/U$4 ( \56258 , \56257 );
and \g130606/U$2 ( \56259 , \56215 , \56258 );
and \g130607/U$2 ( \56260 , \56214 , \56257 );
not \g131030/U$3 ( \56261 , \50362 );
and \g131071/U$2 ( \56262 , \49888 , \50587 );
and \g131071/U$3 ( \56263 , \50588 , \50019 );
nor \g131071/U$1 ( \56264 , \56262 , \56263 );
not \g131030/U$4 ( \56265 , \56264 );
or \g131030/U$2 ( \56266 , \56261 , \56265 );
or \g131030/U$5 ( \56267 , \56264 , \50362 );
nand \g131030/U$1 ( \56268 , \56266 , \56267 );
not \g131418/U$3 ( \56269 , \49233 );
and \g131450/U$2 ( \56270 , \51117 , \49403 );
and \g131450/U$3 ( \56271 , \49405 , \51098 );
nor \g131450/U$1 ( \56272 , \56270 , \56271 );
not \g131418/U$4 ( \56273 , \56272 );
or \g131418/U$2 ( \56274 , \56269 , \56273 );
or \g131418/U$5 ( \56275 , \56272 , \49233 );
nand \g131418/U$1 ( \56276 , \56274 , \56275 );
xor \g130634/U$4 ( \56277 , \56268 , \56276 );
not \g130687/U$3 ( \56278 , \51120 );
and \g130714/U$2 ( \56279 , \49102 , \52273 );
and \g130714/U$3 ( \56280 , \52270 , \48977 );
nor \g130714/U$1 ( \56281 , \56279 , \56280 );
not \g130687/U$4 ( \56282 , \56281 );
or \g130687/U$2 ( \56283 , \56278 , \56282 );
or \g130687/U$5 ( \56284 , \56281 , \51120 );
nand \g130687/U$1 ( \56285 , \56283 , \56284 );
and \g130634/U$3 ( \56286 , \56277 , \56285 );
and \g130634/U$5 ( \56287 , \56268 , \56276 );
or \g130634/U$2 ( \56288 , \56286 , \56287 );
not \g130633/U$1 ( \56289 , \56288 );
nor \g130607/U$1 ( \56290 , \56260 , \56289 );
nor \g130606/U$1 ( \56291 , \56259 , \56290 );
not \g130390/U$4 ( \56292 , \56291 );
and \g130390/U$2 ( \56293 , \56154 , \56292 );
and \g130399/U$2 ( \56294 , \56153 , \56291 );
not \g130470/U$3 ( \56295 , \55808 );
not \g130470/U$4 ( \56296 , \55850 );
or \g130470/U$2 ( \56297 , \56295 , \56296 );
or \g130470/U$5 ( \56298 , \55850 , \55808 );
nand \g130470/U$1 ( \56299 , \56297 , \56298 );
not \g130429/U$3 ( \56300 , \56299 );
not \g130429/U$4 ( \56301 , \55844 );
and \g130429/U$2 ( \56302 , \56300 , \56301 );
and \g130429/U$5 ( \56303 , \56299 , \55844 );
nor \g130429/U$1 ( \56304 , \56302 , \56303 );
nor \g130399/U$1 ( \56305 , \56294 , \56304 );
nor \g130390/U$1 ( \56306 , \56293 , \56305 );
nor \g130294/U$1 ( \56307 , \56137 , \56306 );
nor \g130291/U$1 ( \56308 , \56134 , \56307 );
or \g130128/U$2 ( \56309 , \56051 , \56308 );
not \g130130/U$3 ( \56310 , \56308 );
not \g130130/U$4 ( \56311 , \56051 );
or \g130130/U$2 ( \56312 , \56310 , \56311 );
not \g130186/U$3 ( \56313 , \56034 );
xor \g130212/U$1 ( \56314 , \55871 , \56039 );
not \g130186/U$4 ( \56315 , \56314 );
or \g130186/U$2 ( \56316 , \56313 , \56315 );
or \g130186/U$5 ( \56317 , \56314 , \56034 );
nand \g130186/U$1 ( \56318 , \56316 , \56317 );
nand \g130130/U$1 ( \56319 , \56312 , \56318 );
nand \g130128/U$1 ( \56320 , \56309 , \56319 );
not \g132149/U$3 ( \56321 , \49925 );
and \g132197/U$2 ( \56322 , \53610 , \50159 );
and \g132197/U$3 ( \56323 , \50160 , \53848 );
nor \g132197/U$1 ( \56324 , \56322 , \56323 );
not \g132149/U$4 ( \56325 , \56324 );
or \g132149/U$2 ( \56326 , \56321 , \56325 );
or \g132149/U$5 ( \56327 , \56324 , \49925 );
nand \g132149/U$1 ( \56328 , \56326 , \56327 );
not \g132680/U$3 ( \56329 , \49014 );
and \g132723/U$2 ( \56330 , \54853 , \49075 );
and \g132723/U$3 ( \56331 , \49074 , \54537 );
nor \g132723/U$1 ( \56332 , \56330 , \56331 );
not \g132680/U$4 ( \56333 , \56332 );
or \g132680/U$2 ( \56334 , \56329 , \56333 );
or \g132680/U$5 ( \56335 , \56332 , \49014 );
nand \g132680/U$1 ( \56336 , \56334 , \56335 );
not \g132807/U$3 ( \56337 , \48685 );
and \g132843/U$2 ( \56338 , \55127 , \48858 );
and \g132843/U$3 ( \56339 , \48860 , \55460 );
nor \g132843/U$1 ( \56340 , \56338 , \56339 );
not \g132807/U$4 ( \56341 , \56340 );
or \g132807/U$2 ( \56342 , \56337 , \56341 );
or \g132807/U$5 ( \56343 , \56340 , \48685 );
nand \g132807/U$1 ( \56344 , \56342 , \56343 );
xor \g456145/U$9 ( \56345 , \56336 , \56344 );
not \g132607/U$3 ( \56346 , \47997 );
xor \g133408/U$1 ( \56347 , \47176 , \47127 );
and \g132654/U$2 ( \56348 , \48063 , \56347 );
xor \g133499/U$1 ( \56349 , \47124 , \47087 );
and \g132654/U$3 ( \56350 , \56349 , \48064 );
nor \g132654/U$1 ( \56351 , \56348 , \56350 );
not \g132607/U$4 ( \56352 , \56351 );
or \g132607/U$2 ( \56353 , \56346 , \56352 );
or \g132607/U$5 ( \56354 , \56351 , \47997 );
nand \g132607/U$1 ( \56355 , \56353 , \56354 );
not \g132709/U$3 ( \56356 , \48159 );
xor \g133274/U$1 ( \56357 , \47226 , \47213 );
and \g132759/U$2 ( \56358 , \48154 , \56357 );
xor \g133344/U$1 ( \56359 , \47179 , \47210 );
and \g132759/U$3 ( \56360 , \56359 , \48155 );
nor \g132759/U$1 ( \56361 , \56358 , \56360 );
not \g132709/U$4 ( \56362 , \56361 );
or \g132709/U$2 ( \56363 , \56356 , \56362 );
or \g132709/U$5 ( \56364 , \56361 , \48159 );
nand \g132709/U$1 ( \56365 , \56363 , \56364 );
xor \g132175/U$4 ( \56366 , \56355 , \56365 );
not \g132485/U$3 ( \56367 , \47935 );
xor \g133757/U$1 ( \56368 , \47041 , \47003 );
and \g132554/U$2 ( \56369 , \47930 , \56368 );
xor \g133886/U$1 ( \56370 , \47038 , \47016 );
and \g132554/U$3 ( \56371 , \56370 , \47931 );
nor \g132554/U$1 ( \56372 , \56369 , \56371 );
not \g132485/U$4 ( \56373 , \56372 );
or \g132485/U$2 ( \56374 , \56367 , \56373 );
or \g132485/U$5 ( \56375 , \56372 , \47935 );
nand \g132485/U$1 ( \56376 , \56374 , \56375 );
xor \g134629/U$1 ( \56377 , \47027 , \47034 );
and \g132422/U$2 ( \56378 , \47914 , \56377 );
xor \g134119/U$1 ( \56379 , \47035 , \47024 );
and \g132422/U$3 ( \56380 , \56379 , \47913 );
nor \g132422/U$1 ( \56381 , \56378 , \56380 );
and \g132339/U$2 ( \56382 , \56381 , \47977 );
not \g132339/U$4 ( \56383 , \56381 );
and \g132339/U$3 ( \56384 , \56383 , \47976 );
nor \g132339/U$1 ( \56385 , \56382 , \56384 );
and \g132289/U$2 ( \56386 , \56376 , \56385 );
and \g132175/U$3 ( \56387 , \56366 , \56386 );
and \g132175/U$5 ( \56388 , \56355 , \56365 );
or \g132175/U$2 ( \56389 , \56387 , \56388 );
xor \g456145/U$9_r1 ( \56390 , \56345 , \56389 );
and \g456145/U$8 ( \56391 , \56328 , \56390 );
not \g132748/U$3 ( \56392 , \49014 );
and \g132782/U$2 ( \56393 , \54853 , \49074 );
and \g132782/U$3 ( \56394 , \49075 , \55127 );
nor \g132782/U$1 ( \56395 , \56393 , \56394 );
not \g132748/U$4 ( \56396 , \56395 );
or \g132748/U$2 ( \56397 , \56392 , \56396 );
or \g132748/U$5 ( \56398 , \56395 , \49014 );
nand \g132748/U$1 ( \56399 , \56397 , \56398 );
not \g132873/U$3 ( \56400 , \48685 );
and \g132914/U$2 ( \56401 , \55460 , \48858 );
and \g132914/U$3 ( \56402 , \55707 , \48860 );
nor \g132914/U$1 ( \56403 , \56401 , \56402 );
not \g132873/U$4 ( \56404 , \56403 );
or \g132873/U$2 ( \56405 , \56400 , \56404 );
or \g132873/U$5 ( \56406 , \56403 , \48685 );
nand \g132873/U$1 ( \56407 , \56405 , \56406 );
xor \g131869/U$4 ( \56408 , \56399 , \56407 );
not \g132608/U$3 ( \56409 , \47997 );
and \g132650/U$2 ( \56410 , \48063 , \56349 );
xor \g133621/U$1 ( \56411 , \47084 , \47044 );
and \g132650/U$3 ( \56412 , \56411 , \48064 );
nor \g132650/U$1 ( \56413 , \56410 , \56412 );
not \g132608/U$4 ( \56414 , \56413 );
or \g132608/U$2 ( \56415 , \56409 , \56414 );
or \g132608/U$5 ( \56416 , \56413 , \47997 );
nand \g132608/U$1 ( \56417 , \56415 , \56416 );
not \g132710/U$3 ( \56418 , \48159 );
and \g132760/U$2 ( \56419 , \48155 , \56347 );
and \g132760/U$3 ( \56420 , \56359 , \48154 );
nor \g132760/U$1 ( \56421 , \56419 , \56420 );
not \g132710/U$4 ( \56422 , \56421 );
or \g132710/U$2 ( \56423 , \56418 , \56422 );
or \g132710/U$5 ( \56424 , \56421 , \48159 );
nand \g132710/U$1 ( \56425 , \56423 , \56424 );
xor \g132186/U$4 ( \56426 , \56417 , \56425 );
not \g132486/U$3 ( \56427 , \47935 );
and \g132553/U$2 ( \56428 , \47930 , \56370 );
and \g132553/U$3 ( \56429 , \56379 , \47931 );
nor \g132553/U$1 ( \56430 , \56428 , \56429 );
not \g132486/U$4 ( \56431 , \56430 );
or \g132486/U$2 ( \56432 , \56427 , \56431 );
or \g132486/U$5 ( \56433 , \56430 , \47935 );
nand \g132486/U$1 ( \56434 , \56432 , \56433 );
nand \g132468/U$1 ( \56435 , \47026 , \47913 );
and \g132451/U$2 ( \56436 , \56435 , \47977 );
not \g132451/U$4 ( \56437 , \56435 );
and \g132451/U$3 ( \56438 , \56437 , \47976 );
nor \g132451/U$1 ( \56439 , \56436 , \56438 );
and \g132390/U$2 ( \56440 , \47976 , \56439 );
and \g132309/U$2 ( \56441 , \56434 , \56440 );
and \g132186/U$3 ( \56442 , \56426 , \56441 );
and \g132186/U$5 ( \56443 , \56417 , \56425 );
or \g132186/U$2 ( \56444 , \56442 , \56443 );
not \g132808/U$3 ( \56445 , \48323 );
xor \g133148/U$1 ( \56446 , \47246 , \47231 );
and \g132844/U$2 ( \56447 , \48334 , \56446 );
xor \g133209/U$1 ( \56448 , \47229 , \46969 );
and \g132844/U$3 ( \56449 , \56448 , \48335 );
nor \g132844/U$1 ( \56450 , \56447 , \56449 );
not \g132808/U$4 ( \56451 , \56450 );
or \g132808/U$2 ( \56452 , \56445 , \56451 );
or \g132808/U$5 ( \56453 , \56450 , \48323 );
nand \g132808/U$1 ( \56454 , \56452 , \56453 );
xor \g131972/U$1 ( \56455 , \56444 , \56454 );
not \g132225/U$3 ( \56456 , \47948 );
and \g132266/U$2 ( \56457 , \47960 , \47026 );
and \g132266/U$3 ( \56458 , \56377 , \47959 );
nor \g132266/U$1 ( \56459 , \56457 , \56458 );
not \g132225/U$4 ( \56460 , \56459 );
or \g132225/U$2 ( \56461 , \56456 , \56460 );
or \g132225/U$5 ( \56462 , \56459 , \47948 );
nand \g132225/U$1 ( \56463 , \56461 , \56462 );
not \g132484/U$3 ( \56464 , \47935 );
and \g132548/U$2 ( \56465 , \47930 , \56411 );
and \g132548/U$3 ( \56466 , \56368 , \47931 );
nor \g132548/U$1 ( \56467 , \56465 , \56466 );
not \g132484/U$4 ( \56468 , \56467 );
or \g132484/U$2 ( \56469 , \56464 , \56468 );
or \g132484/U$5 ( \56470 , \56467 , \47935 );
nand \g132484/U$1 ( \56471 , \56469 , \56470 );
xor \g132061/U$1 ( \56472 , \56463 , \56471 );
and \g132420/U$2 ( \56473 , \47913 , \56370 );
and \g132420/U$3 ( \56474 , \56379 , \47914 );
nor \g132420/U$1 ( \56475 , \56473 , \56474 );
and \g132337/U$2 ( \56476 , \56475 , \47977 );
not \g132337/U$4 ( \56477 , \56475 );
and \g132337/U$3 ( \56478 , \56477 , \47976 );
nor \g132337/U$1 ( \56479 , \56476 , \56478 );
nand \g132318/U$1 ( \56480 , \47026 , \47959 );
not \g132293/U$3 ( \56481 , \56480 );
not \g132293/U$4 ( \56482 , \47948 );
or \g132293/U$2 ( \56483 , \56481 , \56482 );
or \g132293/U$5 ( \56484 , \47948 , \56480 );
nand \g132293/U$1 ( \56485 , \56483 , \56484 );
and \g132242/U$2 ( \56486 , \47948 , \56485 );
xor \g132164/U$1 ( \56487 , \56479 , \56486 );
xor \g132061/U$1_r1 ( \56488 , \56472 , \56487 );
xor \g131972/U$1_r1 ( \56489 , \56455 , \56488 );
and \g131869/U$3 ( \56490 , \56408 , \56489 );
and \g131869/U$5 ( \56491 , \56399 , \56407 );
or \g131869/U$2 ( \56492 , \56490 , \56491 );
xor \g456145/U$11 ( \56493 , \56336 , \56344 );
xor \g456145/U$11_r1 ( \56494 , \56493 , \56389 );
and \g456145/U$10 ( \56495 , \56492 , \56494 );
and \g456145/U$12 ( \56496 , \56328 , \56492 );
or \g456145/U$7 ( \56497 , \56391 , \56495 , \56496 );
not \g132085/U$3 ( \56498 , \49925 );
and \g132127/U$2 ( \56499 , \53610 , \50160 );
and \g132127/U$3 ( \56500 , \50159 , \53300 );
nor \g132127/U$1 ( \56501 , \56499 , \56500 );
not \g132085/U$4 ( \56502 , \56501 );
or \g132085/U$2 ( \56503 , \56498 , \56502 );
or \g132085/U$5 ( \56504 , \56501 , \49925 );
nand \g132085/U$1 ( \56505 , \56503 , \56504 );
not \g132251/U$3 ( \56506 , \49568 );
and \g132302/U$2 ( \56507 , \53848 , \49812 );
and \g132302/U$3 ( \56508 , \49813 , \54015 );
nor \g132302/U$1 ( \56509 , \56507 , \56508 );
not \g132251/U$4 ( \56510 , \56509 );
or \g132251/U$2 ( \56511 , \56506 , \56510 );
or \g132251/U$5 ( \56512 , \56509 , \49568 );
nand \g132251/U$1 ( \56513 , \56511 , \56512 );
xor \g131746/U$1 ( \56514 , \56505 , \56513 );
not \g131786/U$3 ( \56515 , \50759 );
and \g131816/U$2 ( \56516 , \52620 , \51055 );
and \g131816/U$3 ( \56517 , \51053 , \52352 );
nor \g131816/U$1 ( \56518 , \56516 , \56517 );
not \g131786/U$4 ( \56519 , \56518 );
or \g131786/U$2 ( \56520 , \56515 , \56519 );
or \g131786/U$5 ( \56521 , \56518 , \50759 );
nand \g131786/U$1 ( \56522 , \56520 , \56521 );
xor \g131746/U$1_r1 ( \56523 , \56514 , \56522 );
xor \g131672/U$4 ( \56524 , \56497 , \56523 );
and \g132419/U$2 ( \56525 , \47913 , \56368 );
and \g132419/U$3 ( \56526 , \56370 , \47914 );
nor \g132419/U$1 ( \56527 , \56525 , \56526 );
and \g132336/U$2 ( \56528 , \56527 , \47977 );
not \g132336/U$4 ( \56529 , \56527 );
and \g132336/U$3 ( \56530 , \56529 , \47976 );
nor \g132336/U$1 ( \56531 , \56528 , \56530 );
not \g132224/U$3 ( \56532 , \47948 );
and \g132277/U$2 ( \56533 , \47960 , \56377 );
and \g132277/U$3 ( \56534 , \56379 , \47959 );
nor \g132277/U$1 ( \56535 , \56533 , \56534 );
not \g132224/U$4 ( \56536 , \56535 );
or \g132224/U$2 ( \56537 , \56532 , \56536 );
or \g132224/U$5 ( \56538 , \56535 , \47948 );
nand \g132224/U$1 ( \56539 , \56537 , \56538 );
xor \g132173/U$1 ( \56540 , \56531 , \56539 );
not \g132708/U$3 ( \56541 , \48159 );
and \g132753/U$2 ( \56542 , \48155 , \56357 );
and \g132753/U$3 ( \56543 , \56448 , \48154 );
nor \g132753/U$1 ( \56544 , \56542 , \56543 );
not \g132708/U$4 ( \56545 , \56544 );
or \g132708/U$2 ( \56546 , \56541 , \56545 );
or \g132708/U$5 ( \56547 , \56544 , \48159 );
nand \g132708/U$1 ( \56548 , \56546 , \56547 );
xor \g131971/U$4 ( \56549 , \56540 , \56548 );
xor \g132061/U$4 ( \56550 , \56463 , \56471 );
and \g132061/U$3 ( \56551 , \56550 , \56487 );
and \g132061/U$5 ( \56552 , \56463 , \56471 );
or \g132061/U$2 ( \56553 , \56551 , \56552 );
and \g131971/U$3 ( \56554 , \56549 , \56553 );
and \g131971/U$5 ( \56555 , \56540 , \56548 );
or \g131971/U$2 ( \56556 , \56554 , \56555 );
not \g132805/U$3 ( \56557 , \48323 );
and \g132842/U$2 ( \56558 , \48335 , \56167 );
and \g132842/U$3 ( \56559 , \55884 , \48334 );
nor \g132842/U$1 ( \56560 , \56558 , \56559 );
not \g132805/U$4 ( \56561 , \56560 );
or \g132805/U$2 ( \56562 , \56557 , \56561 );
or \g132805/U$5 ( \56563 , \56560 , \48323 );
nand \g132805/U$1 ( \56564 , \56562 , \56563 );
xor \g456146/U$2 ( \56565 , \56556 , \56564 );
not \g132482/U$3 ( \56566 , \47935 );
and \g132546/U$2 ( \56567 , \47930 , \56347 );
and \g132546/U$3 ( \56568 , \56349 , \47931 );
nor \g132546/U$1 ( \56569 , \56567 , \56568 );
not \g132482/U$4 ( \56570 , \56569 );
or \g132482/U$2 ( \56571 , \56566 , \56570 );
or \g132482/U$5 ( \56572 , \56569 , \47935 );
nand \g132482/U$1 ( \56573 , \56571 , \56572 );
not \g132605/U$3 ( \56574 , \47997 );
and \g132664/U$2 ( \56575 , \48063 , \56357 );
and \g132664/U$3 ( \56576 , \56359 , \48064 );
nor \g132664/U$1 ( \56577 , \56575 , \56576 );
not \g132605/U$4 ( \56578 , \56577 );
or \g132605/U$2 ( \56579 , \56574 , \56578 );
or \g132605/U$5 ( \56580 , \56577 , \47997 );
nand \g132605/U$1 ( \56581 , \56579 , \56580 );
xor \g132067/U$1 ( \56582 , \56573 , \56581 );
and \g132173/U$2 ( \56583 , \56531 , \56539 );
xor \g132067/U$1_r1 ( \56584 , \56582 , \56583 );
xor \g456146/U$1 ( \56585 , \56565 , \56584 );
xor \g456145/U$5 ( \56586 , \56336 , \56344 );
and \g456145/U$4 ( \56587 , \56586 , \56389 );
and \g456145/U$6 ( \56588 , \56336 , \56344 );
or \g456145/U$3 ( \56589 , \56587 , \56588 );
not \g132742/U$3 ( \56590 , \48685 );
and \g132781/U$2 ( \56591 , \54853 , \48858 );
and \g132781/U$3 ( \56592 , \48860 , \55127 );
nor \g132781/U$1 ( \56593 , \56591 , \56592 );
not \g132742/U$4 ( \56594 , \56593 );
or \g132742/U$2 ( \56595 , \56590 , \56594 );
or \g132742/U$5 ( \56596 , \56593 , \48685 );
nand \g132742/U$1 ( \56597 , \56595 , \56596 );
not \g132872/U$3 ( \56598 , \48483 );
and \g132908/U$2 ( \56599 , \55460 , \48478 );
and \g132908/U$3 ( \56600 , \55707 , \48479 );
nor \g132908/U$1 ( \56601 , \56599 , \56600 );
not \g132872/U$4 ( \56602 , \56601 );
or \g132872/U$2 ( \56603 , \56598 , \56602 );
or \g132872/U$5 ( \56604 , \56601 , \48483 );
nand \g132872/U$1 ( \56605 , \56603 , \56604 );
xor \g131872/U$1 ( \56606 , \56597 , \56605 );
not \g132483/U$3 ( \56607 , \47935 );
and \g132547/U$2 ( \56608 , \47930 , \56349 );
and \g132547/U$3 ( \56609 , \56411 , \47931 );
nor \g132547/U$1 ( \56610 , \56608 , \56609 );
not \g132483/U$4 ( \56611 , \56610 );
or \g132483/U$2 ( \56612 , \56607 , \56611 );
or \g132483/U$5 ( \56613 , \56610 , \47935 );
nand \g132483/U$1 ( \56614 , \56612 , \56613 );
not \g132606/U$3 ( \56615 , \47997 );
and \g132653/U$2 ( \56616 , \48064 , \56347 );
and \g132653/U$3 ( \56617 , \56359 , \48063 );
nor \g132653/U$1 ( \56618 , \56616 , \56617 );
not \g132606/U$4 ( \56619 , \56618 );
or \g132606/U$2 ( \56620 , \56615 , \56619 );
or \g132606/U$5 ( \56621 , \56618 , \47997 );
nand \g132606/U$1 ( \56622 , \56620 , \56621 );
xor \g132068/U$4 ( \56623 , \56614 , \56622 );
and \g132164/U$2 ( \56624 , \56479 , \56486 );
and \g132068/U$3 ( \56625 , \56623 , \56624 );
and \g132068/U$5 ( \56626 , \56614 , \56622 );
or \g132068/U$2 ( \56627 , \56625 , \56626 );
not \g132717/U$3 ( \56628 , \48159 );
and \g132758/U$2 ( \56629 , \48154 , \56446 );
and \g132758/U$3 ( \56630 , \56448 , \48155 );
nor \g132758/U$1 ( \56631 , \56629 , \56630 );
not \g132717/U$4 ( \56632 , \56631 );
or \g132717/U$2 ( \56633 , \56628 , \56632 );
or \g132717/U$5 ( \56634 , \56631 , \48159 );
nand \g132717/U$1 ( \56635 , \56633 , \56634 );
xor \g131975/U$1 ( \56636 , \56627 , \56635 );
and \g132416/U$2 ( \56637 , \47913 , \56411 );
and \g132416/U$3 ( \56638 , \56368 , \47914 );
nor \g132416/U$1 ( \56639 , \56637 , \56638 );
and \g132334/U$2 ( \56640 , \56639 , \47977 );
not \g132334/U$4 ( \56641 , \56639 );
and \g132334/U$3 ( \56642 , \56641 , \47976 );
nor \g132334/U$1 ( \56643 , \56640 , \56642 );
not \g135565/U$2 ( \56644 , \56377 );
nor \g135565/U$1 ( \56645 , \56644 , \40060 );
xor \g132137/U$1 ( \56646 , \56643 , \56645 );
not \g132223/U$3 ( \56647 , \47948 );
and \g132276/U$2 ( \56648 , \47959 , \56370 );
and \g132276/U$3 ( \56649 , \56379 , \47960 );
nor \g132276/U$1 ( \56650 , \56648 , \56649 );
not \g132223/U$4 ( \56651 , \56650 );
or \g132223/U$2 ( \56652 , \56647 , \56651 );
or \g132223/U$5 ( \56653 , \56650 , \47948 );
nand \g132223/U$1 ( \56654 , \56652 , \56653 );
xor \g132137/U$1_r1 ( \56655 , \56646 , \56654 );
xor \g131975/U$1_r1 ( \56656 , \56636 , \56655 );
xor \g131872/U$1_r1 ( \56657 , \56606 , \56656 );
xor \g456146/U$1_r1 ( \56658 , \56589 , \56657 );
xor \g456146/U$1_r2 ( \56659 , \56585 , \56658 );
and \g131672/U$3 ( \56660 , \56524 , \56659 );
and \g131672/U$5 ( \56661 , \56497 , \56523 );
or \g131672/U$2 ( \56662 , \56660 , \56661 );
xor \g131972/U$4 ( \56663 , \56444 , \56454 );
and \g131972/U$3 ( \56664 , \56663 , \56488 );
and \g131972/U$5 ( \56665 , \56444 , \56454 );
or \g131972/U$2 ( \56666 , \56664 , \56665 );
not \g132529/U$3 ( \56667 , \49233 );
and \g132570/U$2 ( \56668 , \54251 , \49403 );
and \g132570/U$3 ( \56669 , \49405 , \54529 );
nor \g132570/U$1 ( \56670 , \56668 , \56669 );
not \g132529/U$4 ( \56671 , \56670 );
or \g132529/U$2 ( \56672 , \56667 , \56671 );
or \g132529/U$5 ( \56673 , \56670 , \49233 );
nand \g132529/U$1 ( \56674 , \56672 , \56673 );
xor \g131878/U$1 ( \56675 , \56666 , \56674 );
xor \g131971/U$1 ( \56676 , \56540 , \56548 );
xor \g131971/U$1_r1 ( \56677 , \56676 , \56553 );
xor \g131878/U$1_r1 ( \56678 , \56675 , \56677 );
and \g131638/U$2 ( \56679 , \51604 , \52270 );
and \g131638/U$3 ( \56680 , \52273 , \51854 );
nor \g131638/U$1 ( \56681 , \56679 , \56680 );
and \g131595/U$2 ( \56682 , \56681 , \51513 );
not \g131595/U$4 ( \56683 , \56681 );
and \g131595/U$3 ( \56684 , \56683 , \51120 );
nor \g131595/U$1 ( \56685 , \56682 , \56684 );
xor \g456125/U$5 ( \56686 , \56678 , \56685 );
xor \g132289/U$1 ( \56687 , \56376 , \56385 );
not \g132826/U$3 ( \56688 , \48323 );
and \g132846/U$2 ( \56689 , \48335 , \56357 );
and \g132846/U$3 ( \56690 , \56448 , \48334 );
nor \g132846/U$1 ( \56691 , \56689 , \56690 );
not \g132826/U$4 ( \56692 , \56691 );
or \g132826/U$2 ( \56693 , \56688 , \56692 );
or \g132826/U$5 ( \56694 , \56691 , \48323 );
nand \g132826/U$1 ( \56695 , \56693 , \56694 );
xor \g132094/U$4 ( \56696 , \56687 , \56695 );
and \g132401/U$2 ( \56697 , \47914 , \47026 );
and \g132401/U$3 ( \56698 , \56377 , \47913 );
nor \g132401/U$1 ( \56699 , \56697 , \56698 );
and \g132340/U$2 ( \56700 , \56699 , \47977 );
not \g132340/U$4 ( \56701 , \56699 );
and \g132340/U$3 ( \56702 , \56701 , \47976 );
nor \g132340/U$1 ( \56703 , \56700 , \56702 );
not \g132611/U$3 ( \56704 , \47997 );
and \g132663/U$2 ( \56705 , \48063 , \56411 );
and \g132663/U$3 ( \56706 , \56368 , \48064 );
nor \g132663/U$1 ( \56707 , \56705 , \56706 );
not \g132611/U$4 ( \56708 , \56707 );
or \g132611/U$2 ( \56709 , \56704 , \56708 );
or \g132611/U$5 ( \56710 , \56707 , \47997 );
nand \g132611/U$1 ( \56711 , \56709 , \56710 );
xor \g132187/U$4 ( \56712 , \56703 , \56711 );
xor \g132309/U$1 ( \56713 , \56434 , \56440 );
and \g132187/U$3 ( \56714 , \56712 , \56713 );
and \g132187/U$5 ( \56715 , \56703 , \56711 );
or \g132187/U$2 ( \56716 , \56714 , \56715 );
and \g132094/U$3 ( \56717 , \56696 , \56716 );
and \g132094/U$5 ( \56718 , \56687 , \56695 );
or \g132094/U$2 ( \56719 , \56717 , \56718 );
not \g132895/U$3 ( \56720 , \48483 );
and \g132939/U$2 ( \56721 , \48479 , \56167 );
and \g132939/U$3 ( \56722 , \55884 , \48478 );
nor \g132939/U$1 ( \56723 , \56721 , \56722 );
not \g132895/U$4 ( \56724 , \56723 );
or \g132895/U$2 ( \56725 , \56720 , \56724 );
or \g132895/U$5 ( \56726 , \56723 , \48483 );
nand \g132895/U$1 ( \56727 , \56725 , \56726 );
xor \g131994/U$4 ( \56728 , \56719 , \56727 );
xor \g132175/U$1 ( \56729 , \56355 , \56365 );
xor \g132175/U$1_r1 ( \56730 , \56729 , \56386 );
and \g131994/U$3 ( \56731 , \56728 , \56730 );
and \g131994/U$5 ( \56732 , \56719 , \56727 );
or \g131994/U$2 ( \56733 , \56731 , \56732 );
not \g132342/U$3 ( \56734 , \49568 );
and \g132424/U$2 ( \56735 , \54185 , \49813 );
and \g132424/U$3 ( \56736 , \49812 , \54015 );
nor \g132424/U$1 ( \56737 , \56735 , \56736 );
not \g132342/U$4 ( \56738 , \56737 );
or \g132342/U$2 ( \56739 , \56734 , \56738 );
or \g132342/U$5 ( \56740 , \56737 , \49568 );
nand \g132342/U$1 ( \56741 , \56739 , \56740 );
xor \g131870/U$1 ( \56742 , \56733 , \56741 );
not \g132813/U$3 ( \56743 , \48323 );
and \g132849/U$2 ( \56744 , \48335 , \56446 );
and \g132849/U$3 ( \56745 , \56167 , \48334 );
nor \g132849/U$1 ( \56746 , \56744 , \56745 );
not \g132813/U$4 ( \56747 , \56746 );
or \g132813/U$2 ( \56748 , \56743 , \56747 );
or \g132813/U$5 ( \56749 , \56746 , \48323 );
nand \g132813/U$1 ( \56750 , \56748 , \56749 );
not \g132906/U$3 ( \56751 , \48483 );
and \g132943/U$2 ( \56752 , \48479 , \55884 );
and \g132943/U$3 ( \56753 , \55707 , \48478 );
nor \g132943/U$1 ( \56754 , \56752 , \56753 );
not \g132906/U$4 ( \56755 , \56754 );
or \g132906/U$2 ( \56756 , \56751 , \56755 );
or \g132906/U$5 ( \56757 , \56754 , \48483 );
nand \g132906/U$1 ( \56758 , \56756 , \56757 );
xor \g131973/U$1 ( \56759 , \56750 , \56758 );
xor \g132068/U$1 ( \56760 , \56614 , \56622 );
xor \g132068/U$1_r1 ( \56761 , \56760 , \56624 );
xor \g131973/U$1_r1 ( \56762 , \56759 , \56761 );
xor \g131870/U$1_r1 ( \56763 , \56742 , \56762 );
and \g456125/U$4 ( \56764 , \56686 , \56763 );
and \g456125/U$6 ( \56765 , \56678 , \56685 );
or \g456125/U$3 ( \56766 , \56764 , \56765 );
not \g131850/U$3 ( \56767 , \50759 );
and \g131891/U$2 ( \56768 , \52620 , \51053 );
and \g131891/U$3 ( \56769 , \51055 , \52883 );
nor \g131891/U$1 ( \56770 , \56768 , \56769 );
not \g131850/U$4 ( \56771 , \56770 );
or \g131850/U$2 ( \56772 , \56767 , \56771 );
or \g131850/U$5 ( \56773 , \56770 , \50759 );
nand \g131850/U$1 ( \56774 , \56772 , \56773 );
not \g132006/U$3 ( \56775 , \50362 );
and \g132044/U$2 ( \56776 , \52978 , \50587 );
and \g132044/U$3 ( \56777 , \50588 , \53300 );
nor \g132044/U$1 ( \56778 , \56776 , \56777 );
not \g132006/U$4 ( \56779 , \56778 );
or \g132006/U$2 ( \56780 , \56775 , \56779 );
or \g132006/U$5 ( \56781 , \56778 , \50362 );
nand \g132006/U$1 ( \56782 , \56780 , \56781 );
xor \g131674/U$4 ( \56783 , \56774 , \56782 );
not \g131725/U$3 ( \56784 , \51124 );
and \g131766/U$2 ( \56785 , \52108 , \51517 );
and \g131766/U$3 ( \56786 , \51518 , \52352 );
nor \g131766/U$1 ( \56787 , \56785 , \56786 );
not \g131725/U$4 ( \56788 , \56787 );
or \g131725/U$2 ( \56789 , \56784 , \56788 );
or \g131725/U$5 ( \56790 , \56787 , \51124 );
nand \g131725/U$1 ( \56791 , \56789 , \56790 );
and \g131674/U$3 ( \56792 , \56783 , \56791 );
and \g131674/U$5 ( \56793 , \56774 , \56782 );
or \g131674/U$2 ( \56794 , \56792 , \56793 );
xor \g456117/U$5 ( \56795 , \56766 , \56794 );
not \g131657/U$3 ( \56796 , \51124 );
and \g131698/U$2 ( \56797 , \52108 , \51518 );
and \g131698/U$3 ( \56798 , \51517 , \51854 );
nor \g131698/U$1 ( \56799 , \56797 , \56798 );
not \g131657/U$4 ( \56800 , \56799 );
or \g131657/U$2 ( \56801 , \56796 , \56800 );
or \g131657/U$5 ( \56802 , \56799 , \51124 );
nand \g131657/U$1 ( \56803 , \56801 , \56802 );
not \g131925/U$3 ( \56804 , \50362 );
and \g131960/U$2 ( \56805 , \52978 , \50588 );
and \g131960/U$3 ( \56806 , \50587 , \52883 );
nor \g131960/U$1 ( \56807 , \56805 , \56806 );
not \g131925/U$4 ( \56808 , \56807 );
or \g131925/U$2 ( \56809 , \56804 , \56808 );
or \g131925/U$5 ( \56810 , \56807 , \50362 );
nand \g131925/U$1 ( \56811 , \56809 , \56810 );
xor \g131610/U$1 ( \56812 , \56803 , \56811 );
xor \g131878/U$4 ( \56813 , \56666 , \56674 );
and \g131878/U$3 ( \56814 , \56813 , \56677 );
and \g131878/U$5 ( \56815 , \56666 , \56674 );
or \g131878/U$2 ( \56816 , \56814 , \56815 );
xor \g131610/U$1_r1 ( \56817 , \56812 , \56816 );
and \g456117/U$4 ( \56818 , \56795 , \56817 );
and \g456117/U$6 ( \56819 , \56766 , \56794 );
or \g456117/U$3 ( \56820 , \56818 , \56819 );
xor \g131344/U$4 ( \56821 , \56662 , \56820 );
xor \g456146/U$9 ( \56822 , \56556 , \56564 );
xor \g456146/U$9_r1 ( \56823 , \56822 , \56584 );
and \g456146/U$8 ( \56824 , \56589 , \56823 );
xor \g456146/U$11 ( \56825 , \56556 , \56564 );
xor \g456146/U$11_r1 ( \56826 , \56825 , \56584 );
and \g456146/U$10 ( \56827 , \56657 , \56826 );
and \g456146/U$12 ( \56828 , \56589 , \56657 );
or \g456146/U$7 ( \56829 , \56824 , \56827 , \56828 );
not \g132453/U$3 ( \56830 , \49233 );
and \g132500/U$2 ( \56831 , \54185 , \49403 );
and \g132500/U$3 ( \56832 , \49405 , \54251 );
nor \g132500/U$1 ( \56833 , \56831 , \56832 );
not \g132453/U$4 ( \56834 , \56833 );
or \g132453/U$2 ( \56835 , \56830 , \56834 );
or \g132453/U$5 ( \56836 , \56833 , \49233 );
nand \g132453/U$1 ( \56837 , \56835 , \56836 );
not \g132615/U$3 ( \56838 , \49014 );
and \g132658/U$2 ( \56839 , \54537 , \49075 );
and \g132658/U$3 ( \56840 , \49074 , \54529 );
nor \g132658/U$1 ( \56841 , \56839 , \56840 );
not \g132615/U$4 ( \56842 , \56841 );
or \g132615/U$2 ( \56843 , \56838 , \56842 );
or \g132615/U$5 ( \56844 , \56841 , \49014 );
nand \g132615/U$1 ( \56845 , \56843 , \56844 );
xor \g456127/U$5 ( \56846 , \56837 , \56845 );
xor \g131973/U$4 ( \56847 , \56750 , \56758 );
and \g131973/U$3 ( \56848 , \56847 , \56761 );
and \g131973/U$5 ( \56849 , \56750 , \56758 );
or \g131973/U$2 ( \56850 , \56848 , \56849 );
and \g456127/U$4 ( \56851 , \56846 , \56850 );
and \g456127/U$6 ( \56852 , \56837 , \56845 );
or \g456127/U$3 ( \56853 , \56851 , \56852 );
xor \g131421/U$1 ( \56854 , \56829 , \56853 );
not \g131481/U$3 ( \56855 , \51120 );
and \g131519/U$2 ( \56856 , \51564 , \52273 );
and \g131519/U$3 ( \56857 , \52270 , \51098 );
nor \g131519/U$1 ( \56858 , \56856 , \56857 );
not \g131481/U$4 ( \56859 , \56858 );
or \g131481/U$2 ( \56860 , \56855 , \56859 );
or \g131481/U$5 ( \56861 , \56858 , \51120 );
nand \g131481/U$1 ( \56862 , \56860 , \56861 );
xor \g131421/U$1_r1 ( \56863 , \56854 , \56862 );
and \g131344/U$3 ( \56864 , \56821 , \56863 );
and \g131344/U$5 ( \56865 , \56662 , \56820 );
or \g131344/U$2 ( \56866 , \56864 , \56865 );
xor \g131870/U$4 ( \56867 , \56733 , \56741 );
and \g131870/U$3 ( \56868 , \56867 , \56762 );
and \g131870/U$5 ( \56869 , \56733 , \56741 );
or \g131870/U$2 ( \56870 , \56868 , \56869 );
xor \g456127/U$9 ( \56871 , \56837 , \56845 );
xor \g456127/U$9_r1 ( \56872 , \56871 , \56850 );
and \g456127/U$8 ( \56873 , \56870 , \56872 );
not \g131545/U$3 ( \56874 , \51120 );
and \g131586/U$2 ( \56875 , \51604 , \52273 );
and \g131586/U$3 ( \56876 , \52270 , \51564 );
nor \g131586/U$1 ( \56877 , \56875 , \56876 );
not \g131545/U$4 ( \56878 , \56877 );
or \g131545/U$2 ( \56879 , \56874 , \56878 );
or \g131545/U$5 ( \56880 , \56877 , \51120 );
nand \g131545/U$1 ( \56881 , \56879 , \56880 );
xor \g456127/U$11 ( \56882 , \56837 , \56845 );
xor \g456127/U$11_r1 ( \56883 , \56882 , \56850 );
and \g456127/U$10 ( \56884 , \56881 , \56883 );
and \g456127/U$12 ( \56885 , \56870 , \56881 );
or \g456127/U$7 ( \56886 , \56873 , \56884 , \56885 );
not \g131849/U$3 ( \56887 , \50362 );
and \g131892/U$2 ( \56888 , \52620 , \50587 );
and \g131892/U$3 ( \56889 , \50588 , \52883 );
nor \g131892/U$1 ( \56890 , \56888 , \56889 );
not \g131849/U$4 ( \56891 , \56890 );
or \g131849/U$2 ( \56892 , \56887 , \56891 );
or \g131849/U$5 ( \56893 , \56890 , \50362 );
nand \g131849/U$1 ( \56894 , \56892 , \56893 );
not \g132154/U$3 ( \56895 , \49568 );
and \g132200/U$2 ( \56896 , \53610 , \49812 );
and \g132200/U$3 ( \56897 , \49813 , \53848 );
nor \g132200/U$1 ( \56898 , \56896 , \56897 );
not \g132154/U$4 ( \56899 , \56898 );
or \g132154/U$2 ( \56900 , \56895 , \56899 );
or \g132154/U$5 ( \56901 , \56898 , \49568 );
nand \g132154/U$1 ( \56902 , \56900 , \56901 );
xor \g131673/U$1 ( \56903 , \56894 , \56902 );
not \g131726/U$3 ( \56904 , \50759 );
and \g131758/U$2 ( \56905 , \52108 , \51053 );
and \g131758/U$3 ( \56906 , \51055 , \52352 );
nor \g131758/U$1 ( \56907 , \56905 , \56906 );
not \g131726/U$4 ( \56908 , \56907 );
or \g131726/U$2 ( \56909 , \56904 , \56908 );
or \g131726/U$5 ( \56910 , \56907 , \50759 );
nand \g131726/U$1 ( \56911 , \56909 , \56910 );
xor \g131673/U$1_r1 ( \56912 , \56903 , \56911 );
xor \g456113/U$5 ( \56913 , \56886 , \56912 );
not \g132479/U$3 ( \56914 , \47935 );
and \g132550/U$2 ( \56915 , \47931 , \56347 );
and \g132550/U$3 ( \56916 , \56359 , \47930 );
nor \g132550/U$1 ( \56917 , \56915 , \56916 );
not \g132479/U$4 ( \56918 , \56917 );
or \g132479/U$2 ( \56919 , \56914 , \56918 );
or \g132479/U$5 ( \56920 , \56917 , \47935 );
nand \g132479/U$1 ( \56921 , \56919 , \56920 );
not \g132602/U$3 ( \56922 , \47997 );
and \g132649/U$2 ( \56923 , \48064 , \56357 );
and \g132649/U$3 ( \56924 , \56448 , \48063 );
nor \g132649/U$1 ( \56925 , \56923 , \56924 );
not \g132602/U$4 ( \56926 , \56925 );
or \g132602/U$2 ( \56927 , \56922 , \56926 );
or \g132602/U$5 ( \56928 , \56925 , \47997 );
nand \g132602/U$1 ( \56929 , \56927 , \56928 );
xor \g132028/U$1 ( \56930 , \56921 , \56929 );
xor \g132137/U$4 ( \56931 , \56643 , \56645 );
and \g132137/U$3 ( \56932 , \56931 , \56654 );
and \g132137/U$5 ( \56933 , \56643 , \56645 );
or \g132137/U$2 ( \56934 , \56932 , \56933 );
xor \g132028/U$1_r1 ( \56935 , \56930 , \56934 );
not \g132527/U$3 ( \56936 , \49014 );
and \g132574/U$2 ( \56937 , \54251 , \49074 );
and \g132574/U$3 ( \56938 , \49075 , \54529 );
nor \g132574/U$1 ( \56939 , \56937 , \56938 );
not \g132527/U$4 ( \56940 , \56939 );
or \g132527/U$2 ( \56941 , \56936 , \56940 );
or \g132527/U$5 ( \56942 , \56939 , \49014 );
nand \g132527/U$1 ( \56943 , \56941 , \56942 );
xor \g456131/U$2 ( \56944 , \56935 , \56943 );
xor \g131975/U$4 ( \56945 , \56627 , \56635 );
and \g131975/U$3 ( \56946 , \56945 , \56655 );
and \g131975/U$5 ( \56947 , \56627 , \56635 );
or \g131975/U$2 ( \56948 , \56946 , \56947 );
xor \g456131/U$1 ( \56949 , \56944 , \56948 );
not \g131597/U$3 ( \56950 , \51124 );
and \g131637/U$2 ( \56951 , \51604 , \51517 );
and \g131637/U$3 ( \56952 , \51518 , \51854 );
nor \g131637/U$1 ( \56953 , \56951 , \56952 );
not \g131597/U$4 ( \56954 , \56953 );
or \g131597/U$2 ( \56955 , \56950 , \56954 );
or \g131597/U$5 ( \56956 , \56953 , \51124 );
nand \g131597/U$1 ( \56957 , \56955 , \56956 );
xor \g456146/U$5 ( \56958 , \56556 , \56564 );
and \g456146/U$4 ( \56959 , \56958 , \56584 );
and \g456146/U$6 ( \56960 , \56556 , \56564 );
or \g456146/U$3 ( \56961 , \56959 , \56960 );
not \g132338/U$3 ( \56962 , \49233 );
and \g132421/U$2 ( \56963 , \54185 , \49405 );
and \g132421/U$3 ( \56964 , \49403 , \54015 );
nor \g132421/U$1 ( \56965 , \56963 , \56964 );
not \g132338/U$4 ( \56966 , \56965 );
or \g132338/U$2 ( \56967 , \56962 , \56966 );
or \g132338/U$5 ( \56968 , \56965 , \49233 );
nand \g132338/U$1 ( \56969 , \56967 , \56968 );
xor \g131796/U$1 ( \56970 , \56961 , \56969 );
xor \g132067/U$4 ( \56971 , \56573 , \56581 );
and \g132067/U$3 ( \56972 , \56971 , \56583 );
and \g132067/U$5 ( \56973 , \56573 , \56581 );
or \g132067/U$2 ( \56974 , \56972 , \56973 );
not \g132707/U$3 ( \56975 , \48159 );
and \g132757/U$2 ( \56976 , \48155 , \56446 );
and \g132757/U$3 ( \56977 , \56167 , \48154 );
nor \g132757/U$1 ( \56978 , \56976 , \56977 );
not \g132707/U$4 ( \56979 , \56978 );
or \g132707/U$2 ( \56980 , \56975 , \56979 );
or \g132707/U$5 ( \56981 , \56978 , \48159 );
nand \g132707/U$1 ( \56982 , \56980 , \56981 );
xor \g131970/U$1 ( \56983 , \56974 , \56982 );
and \g132418/U$2 ( \56984 , \47913 , \56349 );
and \g132418/U$3 ( \56985 , \56411 , \47914 );
nor \g132418/U$1 ( \56986 , \56984 , \56985 );
and \g132335/U$2 ( \56987 , \56986 , \47977 );
not \g132335/U$4 ( \56988 , \56986 );
and \g132335/U$3 ( \56989 , \56988 , \47976 );
nor \g132335/U$1 ( \56990 , \56987 , \56989 );
not \g135563/U$2 ( \56991 , \56379 );
nor \g135563/U$1 ( \56992 , \56991 , \40060 );
not \g132222/U$3 ( \56993 , \47948 );
and \g132278/U$2 ( \56994 , \47959 , \56368 );
and \g132278/U$3 ( \56995 , \56370 , \47960 );
nor \g132278/U$1 ( \56996 , \56994 , \56995 );
not \g132222/U$4 ( \56997 , \56996 );
or \g132222/U$2 ( \56998 , \56993 , \56997 );
or \g132222/U$5 ( \56999 , \56996 , \47948 );
nand \g132222/U$1 ( \57000 , \56998 , \56999 );
xor \g132174/U$1 ( \57001 , \56992 , \57000 );
xor \g132108/U$1 ( \57002 , \56990 , \57001 );
xor \g131970/U$1_r1 ( \57003 , \56983 , \57002 );
xor \g131796/U$1_r1 ( \57004 , \56970 , \57003 );
xor \g456131/U$1_r1 ( \57005 , \56957 , \57004 );
xor \g456131/U$1_r2 ( \57006 , \56949 , \57005 );
and \g456113/U$4 ( \57007 , \56913 , \57006 );
and \g456113/U$6 ( \57008 , \56886 , \56912 );
or \g456113/U$3 ( \57009 , \57007 , \57008 );
xor \g131278/U$4 ( \57010 , \56866 , \57009 );
not \g132449/U$3 ( \57011 , \49014 );
and \g132496/U$2 ( \57012 , \54185 , \49074 );
and \g132496/U$3 ( \57013 , \49075 , \54251 );
nor \g132496/U$1 ( \57014 , \57012 , \57013 );
not \g132449/U$4 ( \57015 , \57014 );
or \g132449/U$2 ( \57016 , \57011 , \57015 );
or \g132449/U$5 ( \57017 , \57014 , \49014 );
nand \g132449/U$1 ( \57018 , \57016 , \57017 );
not \g132604/U$3 ( \57019 , \48685 );
and \g132652/U$2 ( \57020 , \54537 , \48860 );
and \g132652/U$3 ( \57021 , \48858 , \54529 );
nor \g132652/U$1 ( \57022 , \57020 , \57021 );
not \g132604/U$4 ( \57023 , \57022 );
or \g132604/U$2 ( \57024 , \57019 , \57023 );
or \g132604/U$5 ( \57025 , \57022 , \48685 );
nand \g132604/U$1 ( \57026 , \57024 , \57025 );
xor \g131879/U$1 ( \57027 , \57018 , \57026 );
xor \g131970/U$4 ( \57028 , \56974 , \56982 );
and \g131970/U$3 ( \57029 , \57028 , \57002 );
and \g131970/U$5 ( \57030 , \56974 , \56982 );
or \g131970/U$2 ( \57031 , \57029 , \57030 );
xor \g131879/U$1_r1 ( \57032 , \57027 , \57031 );
not \g131655/U$3 ( \57033 , \50759 );
and \g131689/U$2 ( \57034 , \52108 , \51055 );
and \g131689/U$3 ( \57035 , \51053 , \51854 );
nor \g131689/U$1 ( \57036 , \57034 , \57035 );
not \g131655/U$4 ( \57037 , \57036 );
or \g131655/U$2 ( \57038 , \57033 , \57037 );
or \g131655/U$5 ( \57039 , \57036 , \50759 );
nand \g131655/U$1 ( \57040 , \57038 , \57039 );
xor \g456115/U$2 ( \57041 , \57032 , \57040 );
not \g131544/U$3 ( \57042 , \51124 );
and \g131585/U$2 ( \57043 , \51604 , \51518 );
and \g131585/U$3 ( \57044 , \51517 , \51564 );
nor \g131585/U$1 ( \57045 , \57043 , \57044 );
not \g131544/U$4 ( \57046 , \57045 );
or \g131544/U$2 ( \57047 , \57042 , \57046 );
or \g131544/U$5 ( \57048 , \57045 , \51124 );
nand \g131544/U$1 ( \57049 , \57047 , \57048 );
xor \g456115/U$1 ( \57050 , \57041 , \57049 );
xor \g456131/U$9 ( \57051 , \56935 , \56943 );
xor \g456131/U$9_r1 ( \57052 , \57051 , \56948 );
and \g456131/U$8 ( \57053 , \56957 , \57052 );
xor \g456131/U$11 ( \57054 , \56935 , \56943 );
xor \g456131/U$11_r1 ( \57055 , \57054 , \56948 );
and \g456131/U$10 ( \57056 , \57004 , \57055 );
and \g456131/U$12 ( \57057 , \56957 , \57004 );
or \g456131/U$7 ( \57058 , \57053 , \57056 , \57057 );
xor \g131421/U$4 ( \57059 , \56829 , \56853 );
and \g131421/U$3 ( \57060 , \57059 , \56862 );
and \g131421/U$5 ( \57061 , \56829 , \56853 );
or \g131421/U$2 ( \57062 , \57060 , \57061 );
xor \g456115/U$1_r1 ( \57063 , \57058 , \57062 );
xor \g456115/U$1_r2 ( \57064 , \57050 , \57063 );
and \g131278/U$3 ( \57065 , \57010 , \57064 );
and \g131278/U$5 ( \57066 , \56866 , \57009 );
or \g131278/U$2 ( \57067 , \57065 , \57066 );
xor \g456131/U$5 ( \57068 , \56935 , \56943 );
and \g456131/U$4 ( \57069 , \57068 , \56948 );
and \g456131/U$6 ( \57070 , \56935 , \56943 );
or \g456131/U$3 ( \57071 , \57069 , \57070 );
not \g131783/U$3 ( \57072 , \50362 );
and \g131815/U$2 ( \57073 , \52620 , \50588 );
and \g131815/U$3 ( \57074 , \50587 , \52352 );
nor \g131815/U$1 ( \57075 , \57073 , \57074 );
not \g131783/U$4 ( \57076 , \57075 );
or \g131783/U$2 ( \57077 , \57072 , \57076 );
or \g131783/U$5 ( \57078 , \57075 , \50362 );
nand \g131783/U$1 ( \57079 , \57077 , \57078 );
xor \g456133/U$5 ( \57080 , \57071 , \57079 );
xor \g131796/U$4 ( \57081 , \56961 , \56969 );
and \g131796/U$3 ( \57082 , \57081 , \57003 );
and \g131796/U$5 ( \57083 , \56961 , \56969 );
or \g131796/U$2 ( \57084 , \57082 , \57083 );
and \g456133/U$4 ( \57085 , \57080 , \57084 );
and \g456133/U$6 ( \57086 , \57071 , \57079 );
or \g456133/U$3 ( \57087 , \57085 , \57086 );
not \g131921/U$3 ( \57088 , \49925 );
and \g131958/U$2 ( \57089 , \52978 , \50160 );
and \g131958/U$3 ( \57090 , \50159 , \52883 );
nor \g131958/U$1 ( \57091 , \57089 , \57090 );
not \g131921/U$4 ( \57092 , \57091 );
or \g131921/U$2 ( \57093 , \57088 , \57092 );
or \g131921/U$5 ( \57094 , \57091 , \49925 );
nand \g131921/U$1 ( \57095 , \57093 , \57094 );
not \g132248/U$3 ( \57096 , \49233 );
and \g132299/U$2 ( \57097 , \53848 , \49403 );
and \g132299/U$3 ( \57098 , \49405 , \54015 );
nor \g132299/U$1 ( \57099 , \57097 , \57098 );
not \g132248/U$4 ( \57100 , \57099 );
or \g132248/U$2 ( \57101 , \57096 , \57100 );
or \g132248/U$5 ( \57102 , \57099 , \49233 );
nand \g132248/U$1 ( \57103 , \57101 , \57102 );
xor \g131828/U$4 ( \57104 , \57095 , \57103 );
not \g132802/U$3 ( \57105 , \48323 );
and \g132840/U$2 ( \57106 , \48334 , \55460 );
and \g132840/U$3 ( \57107 , \55707 , \48335 );
nor \g132840/U$1 ( \57108 , \57106 , \57107 );
not \g132802/U$4 ( \57109 , \57108 );
or \g132802/U$2 ( \57110 , \57105 , \57109 );
or \g132802/U$5 ( \57111 , \57108 , \48323 );
nand \g132802/U$1 ( \57112 , \57110 , \57111 );
not \g132741/U$3 ( \57113 , \48483 );
and \g132780/U$2 ( \57114 , \54853 , \48478 );
and \g132780/U$3 ( \57115 , \55127 , \48479 );
nor \g132780/U$1 ( \57116 , \57114 , \57115 );
not \g132741/U$4 ( \57117 , \57116 );
or \g132741/U$2 ( \57118 , \57113 , \57117 );
or \g132741/U$5 ( \57119 , \57116 , \48483 );
nand \g132741/U$1 ( \57120 , \57118 , \57119 );
xor \g131913/U$1 ( \57121 , \57112 , \57120 );
not \g132480/U$3 ( \57122 , \47935 );
and \g132545/U$2 ( \57123 , \47930 , \56357 );
and \g132545/U$3 ( \57124 , \56359 , \47931 );
nor \g132545/U$1 ( \57125 , \57123 , \57124 );
not \g132480/U$4 ( \57126 , \57125 );
or \g132480/U$2 ( \57127 , \57122 , \57126 );
or \g132480/U$5 ( \57128 , \57125 , \47935 );
nand \g132480/U$1 ( \57129 , \57127 , \57128 );
not \g132603/U$3 ( \57130 , \47997 );
and \g132651/U$2 ( \57131 , \48063 , \56446 );
and \g132651/U$3 ( \57132 , \56448 , \48064 );
nor \g132651/U$1 ( \57133 , \57131 , \57132 );
not \g132603/U$4 ( \57134 , \57133 );
or \g132603/U$2 ( \57135 , \57130 , \57134 );
or \g132603/U$5 ( \57136 , \57133 , \47997 );
nand \g132603/U$1 ( \57137 , \57135 , \57136 );
xor \g132021/U$1 ( \57138 , \57129 , \57137 );
and \g132108/U$2 ( \57139 , \56990 , \57001 );
xor \g132021/U$1_r1 ( \57140 , \57138 , \57139 );
xor \g131913/U$1_r1 ( \57141 , \57121 , \57140 );
and \g131828/U$3 ( \57142 , \57104 , \57141 );
and \g131828/U$5 ( \57143 , \57095 , \57103 );
or \g131828/U$2 ( \57144 , \57142 , \57143 );
xor \g456112/U$2 ( \57145 , \57087 , \57144 );
xor \g456115/U$5 ( \57146 , \57032 , \57040 );
and \g456115/U$4 ( \57147 , \57146 , \57049 );
and \g456115/U$6 ( \57148 , \57032 , \57040 );
or \g456115/U$3 ( \57149 , \57147 , \57148 );
xor \g456112/U$1 ( \57150 , \57145 , \57149 );
xor \g131673/U$4 ( \57151 , \56894 , \56902 );
and \g131673/U$3 ( \57152 , \57151 , \56911 );
and \g131673/U$5 ( \57153 , \56894 , \56902 );
or \g131673/U$2 ( \57154 , \57152 , \57153 );
xor \g456133/U$9 ( \57155 , \57071 , \57079 );
xor \g456133/U$9_r1 ( \57156 , \57155 , \57084 );
and \g456133/U$8 ( \57157 , \57154 , \57156 );
xor \g131828/U$1 ( \57158 , \57095 , \57103 );
xor \g131828/U$1_r1 ( \57159 , \57158 , \57141 );
xor \g456133/U$11 ( \57160 , \57071 , \57079 );
xor \g456133/U$11_r1 ( \57161 , \57160 , \57084 );
and \g456133/U$10 ( \57162 , \57159 , \57161 );
and \g456133/U$12 ( \57163 , \57154 , \57159 );
or \g456133/U$7 ( \57164 , \57157 , \57162 , \57163 );
xor \g131913/U$4 ( \57165 , \57112 , \57120 );
and \g131913/U$3 ( \57166 , \57165 , \57140 );
and \g131913/U$5 ( \57167 , \57112 , \57120 );
or \g131913/U$2 ( \57168 , \57166 , \57167 );
not \g132003/U$3 ( \57169 , \49568 );
and \g132042/U$2 ( \57170 , \52978 , \49812 );
and \g132042/U$3 ( \57171 , \49813 , \53300 );
nor \g132042/U$1 ( \57172 , \57170 , \57171 );
not \g132003/U$4 ( \57173 , \57172 );
or \g132003/U$2 ( \57174 , \57169 , \57173 );
or \g132003/U$5 ( \57175 , \57172 , \49568 );
nand \g132003/U$1 ( \57176 , \57174 , \57175 );
xor \g456142/U$2 ( \57177 , \57168 , \57176 );
not \g132706/U$3 ( \57178 , \48159 );
and \g132766/U$2 ( \57179 , \48155 , \55884 );
and \g132766/U$3 ( \57180 , \55707 , \48154 );
nor \g132766/U$1 ( \57181 , \57179 , \57180 );
not \g132706/U$4 ( \57182 , \57181 );
or \g132706/U$2 ( \57183 , \57178 , \57182 );
or \g132706/U$5 ( \57184 , \57181 , \48159 );
nand \g132706/U$1 ( \57185 , \57183 , \57184 );
not \g132801/U$3 ( \57186 , \48323 );
and \g132839/U$2 ( \57187 , \48334 , \55127 );
and \g132839/U$3 ( \57188 , \55460 , \48335 );
nor \g132839/U$1 ( \57189 , \57187 , \57188 );
not \g132801/U$4 ( \57190 , \57189 );
or \g132801/U$2 ( \57191 , \57186 , \57190 );
or \g132801/U$5 ( \57192 , \57189 , \48323 );
nand \g132801/U$1 ( \57193 , \57191 , \57192 );
xor \g131969/U$1 ( \57194 , \57185 , \57193 );
not \g135562/U$2 ( \57195 , \56370 );
nor \g135562/U$1 ( \57196 , \57195 , \40060 );
not \g132221/U$3 ( \57197 , \47948 );
and \g132275/U$2 ( \57198 , \47959 , \56411 );
and \g132275/U$3 ( \57199 , \56368 , \47960 );
nor \g132275/U$1 ( \57200 , \57198 , \57199 );
not \g132221/U$4 ( \57201 , \57200 );
or \g132221/U$2 ( \57202 , \57197 , \57201 );
or \g132221/U$5 ( \57203 , \57200 , \47948 );
nand \g132221/U$1 ( \57204 , \57202 , \57203 );
and \g132169/U$2 ( \57205 , \57196 , \57204 );
and \g132412/U$2 ( \57206 , \47914 , \56347 );
and \g132412/U$3 ( \57207 , \56359 , \47913 );
nor \g132412/U$1 ( \57208 , \57206 , \57207 );
and \g132331/U$2 ( \57209 , \57208 , \47977 );
not \g132331/U$4 ( \57210 , \57208 );
and \g132331/U$3 ( \57211 , \57210 , \47976 );
nor \g132331/U$1 ( \57212 , \57209 , \57211 );
xor \g132059/U$1 ( \57213 , \57205 , \57212 );
not \g135559/U$2 ( \57214 , \56368 );
nor \g135559/U$1 ( \57215 , \57214 , \40060 );
not \g132220/U$3 ( \57216 , \47948 );
and \g132272/U$2 ( \57217 , \47959 , \56349 );
and \g132272/U$3 ( \57218 , \56411 , \47960 );
nor \g132272/U$1 ( \57219 , \57217 , \57218 );
not \g132220/U$4 ( \57220 , \57219 );
or \g132220/U$2 ( \57221 , \57216 , \57220 );
or \g132220/U$5 ( \57222 , \57219 , \47948 );
nand \g132220/U$1 ( \57223 , \57221 , \57222 );
xor \g132165/U$1 ( \57224 , \57215 , \57223 );
xor \g132059/U$1_r1 ( \57225 , \57213 , \57224 );
xor \g131969/U$1_r1 ( \57226 , \57194 , \57225 );
xor \g456142/U$1 ( \57227 , \57177 , \57226 );
not \g132082/U$3 ( \57228 , \49568 );
and \g132124/U$2 ( \57229 , \53610 , \49813 );
and \g132124/U$3 ( \57230 , \49812 , \53300 );
nor \g132124/U$1 ( \57231 , \57229 , \57230 );
not \g132082/U$4 ( \57232 , \57231 );
or \g132082/U$2 ( \57233 , \57228 , \57232 );
or \g132082/U$5 ( \57234 , \57231 , \49568 );
nand \g132082/U$1 ( \57235 , \57233 , \57234 );
not \g132804/U$3 ( \57236 , \48323 );
and \g132855/U$2 ( \57237 , \48335 , \55884 );
and \g132855/U$3 ( \57238 , \55707 , \48334 );
nor \g132855/U$1 ( \57239 , \57237 , \57238 );
not \g132804/U$4 ( \57240 , \57239 );
or \g132804/U$2 ( \57241 , \57236 , \57240 );
or \g132804/U$5 ( \57242 , \57239 , \48323 );
nand \g132804/U$1 ( \57243 , \57241 , \57242 );
not \g132803/U$3 ( \57244 , \48483 );
and \g132841/U$2 ( \57245 , \55127 , \48478 );
and \g132841/U$3 ( \57246 , \55460 , \48479 );
nor \g132841/U$1 ( \57247 , \57245 , \57246 );
not \g132803/U$4 ( \57248 , \57247 );
or \g132803/U$2 ( \57249 , \57244 , \57248 );
or \g132803/U$5 ( \57250 , \57247 , \48483 );
nand \g132803/U$1 ( \57251 , \57249 , \57250 );
xor \g132623/U$4 ( \57252 , \57243 , \57251 );
not \g132678/U$3 ( \57253 , \48685 );
and \g132722/U$2 ( \57254 , \54853 , \48860 );
and \g132722/U$3 ( \57255 , \48858 , \54537 );
nor \g132722/U$1 ( \57256 , \57254 , \57255 );
not \g132678/U$4 ( \57257 , \57256 );
or \g132678/U$2 ( \57258 , \57253 , \57257 );
or \g132678/U$5 ( \57259 , \57256 , \48685 );
nand \g132678/U$1 ( \57260 , \57258 , \57259 );
and \g132623/U$3 ( \57261 , \57252 , \57260 );
and \g132623/U$5 ( \57262 , \57243 , \57251 );
or \g132623/U$2 ( \57263 , \57261 , \57262 );
xor \g131837/U$4 ( \57264 , \57235 , \57263 );
xor \g132028/U$4 ( \57265 , \56921 , \56929 );
and \g132028/U$3 ( \57266 , \57265 , \56934 );
and \g132028/U$5 ( \57267 , \56921 , \56929 );
or \g132028/U$2 ( \57268 , \57266 , \57267 );
not \g132705/U$3 ( \57269 , \48159 );
and \g132756/U$2 ( \57270 , \48155 , \56167 );
and \g132756/U$3 ( \57271 , \55884 , \48154 );
nor \g132756/U$1 ( \57272 , \57270 , \57271 );
not \g132705/U$4 ( \57273 , \57272 );
or \g132705/U$2 ( \57274 , \57269 , \57273 );
or \g132705/U$5 ( \57275 , \57272 , \48159 );
nand \g132705/U$1 ( \57276 , \57274 , \57275 );
xor \g131933/U$1 ( \57277 , \57268 , \57276 );
and \g132174/U$2 ( \57278 , \56992 , \57000 );
and \g132413/U$2 ( \57279 , \47913 , \56347 );
and \g132413/U$3 ( \57280 , \56349 , \47914 );
nor \g132413/U$1 ( \57281 , \57279 , \57280 );
and \g132349/U$2 ( \57282 , \57281 , \47977 );
not \g132349/U$4 ( \57283 , \57281 );
and \g132349/U$3 ( \57284 , \57283 , \47976 );
nor \g132349/U$1 ( \57285 , \57282 , \57284 );
xor \g132064/U$1 ( \57286 , \57278 , \57285 );
xor \g132169/U$1 ( \57287 , \57196 , \57204 );
xor \g132064/U$1_r1 ( \57288 , \57286 , \57287 );
xor \g131933/U$1_r1 ( \57289 , \57277 , \57288 );
and \g131837/U$3 ( \57290 , \57264 , \57289 );
and \g131837/U$5 ( \57291 , \57235 , \57263 );
or \g131837/U$2 ( \57292 , \57290 , \57291 );
not \g131848/U$3 ( \57293 , \49925 );
and \g131899/U$2 ( \57294 , \52620 , \50159 );
and \g131899/U$3 ( \57295 , \50160 , \52883 );
nor \g131899/U$1 ( \57296 , \57294 , \57295 );
not \g131848/U$4 ( \57297 , \57296 );
or \g131848/U$2 ( \57298 , \57293 , \57297 );
or \g131848/U$5 ( \57299 , \57296 , \49925 );
nand \g131848/U$1 ( \57300 , \57298 , \57299 );
not \g132148/U$3 ( \57301 , \49233 );
and \g132196/U$2 ( \57302 , \53610 , \49403 );
and \g132196/U$3 ( \57303 , \49405 , \53848 );
nor \g132196/U$1 ( \57304 , \57302 , \57303 );
not \g132148/U$4 ( \57305 , \57304 );
or \g132148/U$2 ( \57306 , \57301 , \57305 );
or \g132148/U$5 ( \57307 , \57304 , \49233 );
nand \g132148/U$1 ( \57308 , \57306 , \57307 );
xor \g131795/U$1 ( \57309 , \57300 , \57308 );
xor \g132021/U$4 ( \57310 , \57129 , \57137 );
and \g132021/U$3 ( \57311 , \57310 , \57139 );
and \g132021/U$5 ( \57312 , \57129 , \57137 );
or \g132021/U$2 ( \57313 , \57311 , \57312 );
not \g132675/U$3 ( \57314 , \48483 );
and \g132721/U$2 ( \57315 , \54853 , \48479 );
and \g132721/U$3 ( \57316 , \48478 , \54537 );
nor \g132721/U$1 ( \57317 , \57315 , \57316 );
not \g132675/U$4 ( \57318 , \57317 );
or \g132675/U$2 ( \57319 , \57314 , \57318 );
or \g132675/U$5 ( \57320 , \57317 , \48483 );
nand \g132675/U$1 ( \57321 , \57319 , \57320 );
xor \g131874/U$1 ( \57322 , \57313 , \57321 );
not \g132478/U$3 ( \57323 , \47935 );
and \g132544/U$2 ( \57324 , \47931 , \56357 );
and \g132544/U$3 ( \57325 , \56448 , \47930 );
nor \g132544/U$1 ( \57326 , \57324 , \57325 );
not \g132478/U$4 ( \57327 , \57326 );
or \g132478/U$2 ( \57328 , \57323 , \57327 );
or \g132478/U$5 ( \57329 , \57326 , \47935 );
nand \g132478/U$1 ( \57330 , \57328 , \57329 );
not \g132600/U$3 ( \57331 , \47997 );
and \g132666/U$2 ( \57332 , \48064 , \56446 );
and \g132666/U$3 ( \57333 , \56167 , \48063 );
nor \g132666/U$1 ( \57334 , \57332 , \57333 );
not \g132600/U$4 ( \57335 , \57334 );
or \g132600/U$2 ( \57336 , \57331 , \57335 );
or \g132600/U$5 ( \57337 , \57334 , \47997 );
nand \g132600/U$1 ( \57338 , \57336 , \57337 );
xor \g131987/U$1 ( \57339 , \57330 , \57338 );
xor \g132064/U$4 ( \57340 , \57278 , \57285 );
and \g132064/U$3 ( \57341 , \57340 , \57287 );
and \g132064/U$5 ( \57342 , \57278 , \57285 );
or \g132064/U$2 ( \57343 , \57341 , \57342 );
xor \g131987/U$1_r1 ( \57344 , \57339 , \57343 );
xor \g131874/U$1_r1 ( \57345 , \57322 , \57344 );
xor \g131795/U$1_r1 ( \57346 , \57309 , \57345 );
xor \g456142/U$1_r1 ( \57347 , \57292 , \57346 );
xor \g456142/U$1_r2 ( \57348 , \57227 , \57347 );
xor \g456112/U$1_r1 ( \57349 , \57164 , \57348 );
xor \g456112/U$1_r2 ( \57350 , \57150 , \57349 );
and \g131119/U$2 ( \57351 , \57067 , \57350 );
not \g131131/U$3 ( \57352 , \57067 );
not \g131131/U$4 ( \57353 , \57350 );
and \g131131/U$2 ( \57354 , \57352 , \57353 );
xor \g131610/U$4 ( \57355 , \56803 , \56811 );
and \g131610/U$3 ( \57356 , \57355 , \56816 );
and \g131610/U$5 ( \57357 , \56803 , \56811 );
or \g131610/U$2 ( \57358 , \57356 , \57357 );
xor \g131746/U$4 ( \57359 , \56505 , \56513 );
and \g131746/U$3 ( \57360 , \57359 , \56522 );
and \g131746/U$5 ( \57361 , \56505 , \56513 );
or \g131746/U$2 ( \57362 , \57360 , \57361 );
xor \g131557/U$4 ( \57363 , \57358 , \57362 );
not \g132004/U$3 ( \57364 , \49925 );
and \g132043/U$2 ( \57365 , \52978 , \50159 );
and \g132043/U$3 ( \57366 , \50160 , \53300 );
nor \g132043/U$1 ( \57367 , \57365 , \57366 );
not \g132004/U$4 ( \57368 , \57367 );
or \g132004/U$2 ( \57369 , \57364 , \57368 );
or \g132004/U$5 ( \57370 , \57367 , \49925 );
nand \g132004/U$1 ( \57371 , \57369 , \57370 );
xor \g132623/U$1 ( \57372 , \57243 , \57251 );
xor \g132623/U$1_r1 ( \57373 , \57372 , \57260 );
xor \g131801/U$1 ( \57374 , \57371 , \57373 );
xor \g131872/U$4 ( \57375 , \56597 , \56605 );
and \g131872/U$3 ( \57376 , \57375 , \56656 );
and \g131872/U$5 ( \57377 , \56597 , \56605 );
or \g131872/U$2 ( \57378 , \57376 , \57377 );
xor \g131801/U$1_r1 ( \57379 , \57374 , \57378 );
and \g131557/U$3 ( \57380 , \57363 , \57379 );
and \g131557/U$5 ( \57381 , \57358 , \57362 );
or \g131557/U$2 ( \57382 , \57380 , \57381 );
xor \g131837/U$1 ( \57383 , \57235 , \57263 );
xor \g131837/U$1_r1 ( \57384 , \57383 , \57289 );
xor \g131801/U$4 ( \57385 , \57371 , \57373 );
and \g131801/U$3 ( \57386 , \57385 , \57378 );
and \g131801/U$5 ( \57387 , \57371 , \57373 );
or \g131801/U$2 ( \57388 , \57386 , \57387 );
xor \g456109/U$9 ( \57389 , \57384 , \57388 );
not \g131408/U$3 ( \57390 , \51120 );
and \g131452/U$2 ( \57391 , \51117 , \52270 );
and \g131452/U$3 ( \57392 , \52273 , \51098 );
nor \g131452/U$1 ( \57393 , \57391 , \57392 );
not \g131408/U$4 ( \57394 , \57393 );
or \g131408/U$2 ( \57395 , \57390 , \57394 );
or \g131408/U$5 ( \57396 , \57393 , \51120 );
nand \g131408/U$1 ( \57397 , \57395 , \57396 );
xor \g456109/U$9_r1 ( \57398 , \57389 , \57397 );
and \g456109/U$8 ( \57399 , \57382 , \57398 );
xor \g456133/U$2 ( \57400 , \57071 , \57079 );
xor \g456133/U$1 ( \57401 , \57400 , \57084 );
xor \g456133/U$1_r1 ( \57402 , \57154 , \57159 );
xor \g456133/U$1_r2 ( \57403 , \57401 , \57402 );
xor \g456109/U$11 ( \57404 , \57384 , \57388 );
xor \g456109/U$11_r1 ( \57405 , \57404 , \57397 );
and \g456109/U$10 ( \57406 , \57403 , \57405 );
and \g456109/U$12 ( \57407 , \57382 , \57403 );
or \g456109/U$7 ( \57408 , \57399 , \57406 , \57407 );
xor \g456109/U$5 ( \57409 , \57384 , \57388 );
and \g456109/U$4 ( \57410 , \57409 , \57397 );
and \g456109/U$6 ( \57411 , \57384 , \57388 );
or \g456109/U$3 ( \57412 , \57410 , \57411 );
xor \g131879/U$4 ( \57413 , \57018 , \57026 );
and \g131879/U$3 ( \57414 , \57413 , \57031 );
and \g131879/U$5 ( \57415 , \57018 , \57026 );
or \g131879/U$2 ( \57416 , \57414 , \57415 );
not \g131723/U$3 ( \57417 , \50362 );
and \g131756/U$2 ( \57418 , \52108 , \50587 );
and \g131756/U$3 ( \57419 , \50588 , \52352 );
nor \g131756/U$1 ( \57420 , \57418 , \57419 );
not \g131723/U$4 ( \57421 , \57420 );
or \g131723/U$2 ( \57422 , \57417 , \57421 );
or \g131723/U$5 ( \57423 , \57420 , \50362 );
nand \g131723/U$1 ( \57424 , \57422 , \57423 );
xor \g131427/U$1 ( \57425 , \57416 , \57424 );
not \g131479/U$3 ( \57426 , \51124 );
and \g131518/U$2 ( \57427 , \51564 , \51518 );
and \g131518/U$3 ( \57428 , \51517 , \51098 );
nor \g131518/U$1 ( \57429 , \57427 , \57428 );
not \g131479/U$4 ( \57430 , \57429 );
or \g131479/U$2 ( \57431 , \57426 , \57430 );
or \g131479/U$5 ( \57432 , \57429 , \51124 );
nand \g131479/U$1 ( \57433 , \57431 , \57432 );
xor \g131427/U$1_r1 ( \57434 , \57425 , \57433 );
xor \g131246/U$1 ( \57435 , \57412 , \57434 );
not \g132333/U$3 ( \57436 , \49014 );
and \g132415/U$2 ( \57437 , \54185 , \49075 );
and \g132415/U$3 ( \57438 , \49074 , \54015 );
nor \g132415/U$1 ( \57439 , \57437 , \57438 );
not \g132333/U$4 ( \57440 , \57439 );
or \g132333/U$2 ( \57441 , \57436 , \57440 );
or \g132333/U$5 ( \57442 , \57439 , \49014 );
nand \g132333/U$1 ( \57443 , \57441 , \57442 );
not \g132526/U$3 ( \57444 , \48685 );
and \g132565/U$2 ( \57445 , \54251 , \48858 );
and \g132565/U$3 ( \57446 , \48860 , \54529 );
nor \g132565/U$1 ( \57447 , \57445 , \57446 );
not \g132526/U$4 ( \57448 , \57447 );
or \g132526/U$2 ( \57449 , \57444 , \57448 );
or \g132526/U$5 ( \57450 , \57447 , \48685 );
nand \g132526/U$1 ( \57451 , \57449 , \57450 );
xor \g456111/U$2 ( \57452 , \57443 , \57451 );
xor \g131933/U$4 ( \57453 , \57268 , \57276 );
and \g131933/U$3 ( \57454 , \57453 , \57288 );
and \g131933/U$5 ( \57455 , \57268 , \57276 );
or \g131933/U$2 ( \57456 , \57454 , \57455 );
xor \g456111/U$1 ( \57457 , \57452 , \57456 );
not \g131604/U$3 ( \57458 , \50759 );
and \g131630/U$2 ( \57459 , \51604 , \51053 );
and \g131630/U$3 ( \57460 , \51055 , \51854 );
nor \g131630/U$1 ( \57461 , \57459 , \57460 );
not \g131604/U$4 ( \57462 , \57461 );
or \g131604/U$2 ( \57463 , \57458 , \57462 );
or \g131604/U$5 ( \57464 , \57461 , \50759 );
nand \g131604/U$1 ( \57465 , \57463 , \57464 );
not \g131351/U$3 ( \57466 , \51120 );
and \g131384/U$2 ( \57467 , \51117 , \52273 );
and \g131384/U$3 ( \57468 , \52270 , \50957 );
nor \g131384/U$1 ( \57469 , \57467 , \57468 );
not \g131351/U$4 ( \57470 , \57469 );
or \g131351/U$2 ( \57471 , \57466 , \57470 );
or \g131351/U$5 ( \57472 , \57469 , \51120 );
nand \g131351/U$1 ( \57473 , \57471 , \57472 );
xor \g456111/U$1_r1 ( \57474 , \57465 , \57473 );
xor \g456111/U$1_r2 ( \57475 , \57457 , \57474 );
xor \g131246/U$1_r1 ( \57476 , \57435 , \57475 );
xnor \g131205/U$1 ( \57477 , \57408 , \57476 );
not \g131190/U$3 ( \57478 , \57477 );
xor \g456115/U$9 ( \57479 , \57032 , \57040 );
xor \g456115/U$9_r1 ( \57480 , \57479 , \57049 );
and \g456115/U$8 ( \57481 , \57058 , \57480 );
xor \g456115/U$11 ( \57482 , \57032 , \57040 );
xor \g456115/U$11_r1 ( \57483 , \57482 , \57049 );
and \g456115/U$10 ( \57484 , \57062 , \57483 );
and \g456115/U$12 ( \57485 , \57058 , \57062 );
or \g456115/U$7 ( \57486 , \57481 , \57484 , \57485 );
not \g131190/U$4 ( \57487 , \57486 );
and \g131190/U$2 ( \57488 , \57478 , \57487 );
and \g131190/U$5 ( \57489 , \57477 , \57486 );
nor \g131190/U$1 ( \57490 , \57488 , \57489 );
nor \g131131/U$1 ( \57491 , \57354 , \57490 );
nor \g131119/U$1 ( \57492 , \57351 , \57491 );
not \g133315/U$3 ( \57493 , \49925 );
and \g133366/U$2 ( \57494 , \50159 , \56368 );
and \g133366/U$3 ( \57495 , \56370 , \50160 );
nor \g133366/U$1 ( \57496 , \57494 , \57495 );
not \g133315/U$4 ( \57497 , \57496 );
or \g133315/U$2 ( \57498 , \57493 , \57497 );
or \g133315/U$5 ( \57499 , \57496 , \49925 );
nand \g133315/U$1 ( \57500 , \57498 , \57499 );
not \g133223/U$3 ( \57501 , \49568 );
and \g133268/U$2 ( \57502 , \49813 , \56377 );
and \g133268/U$3 ( \57503 , \56379 , \49812 );
nor \g133268/U$1 ( \57504 , \57502 , \57503 );
not \g133223/U$4 ( \57505 , \57504 );
or \g133223/U$2 ( \57506 , \57501 , \57505 );
or \g133223/U$5 ( \57507 , \57504 , \49568 );
nand \g133223/U$1 ( \57508 , \57506 , \57507 );
and \g133180/U$2 ( \57509 , \57500 , \57508 );
not \g133323/U$3 ( \57510 , \50362 );
and \g133361/U$2 ( \57511 , \56347 , \50587 );
and \g133361/U$3 ( \57512 , \50588 , \56349 );
nor \g133361/U$1 ( \57513 , \57511 , \57512 );
not \g133323/U$4 ( \57514 , \57513 );
or \g133323/U$2 ( \57515 , \57510 , \57514 );
or \g133323/U$5 ( \57516 , \57513 , \50362 );
nand \g133323/U$1 ( \57517 , \57515 , \57516 );
xor \g133032/U$4 ( \57518 , \57509 , \57517 );
not \g133228/U$3 ( \57519 , \49568 );
and \g133265/U$2 ( \57520 , \49812 , \56370 );
and \g133265/U$3 ( \57521 , \56379 , \49813 );
nor \g133265/U$1 ( \57522 , \57520 , \57521 );
not \g133228/U$4 ( \57523 , \57522 );
or \g133228/U$2 ( \57524 , \57519 , \57523 );
or \g133228/U$5 ( \57525 , \57522 , \49568 );
nand \g133228/U$1 ( \57526 , \57524 , \57525 );
not \g135551/U$2 ( \57527 , \49233 );
nor \g133220/U$1 ( \57528 , \49404 , \47025 );
nor \g135551/U$1 ( \57529 , \57527 , \57528 );
xor \g133172/U$1 ( \57530 , \57526 , \57529 );
not \g133320/U$3 ( \57531 , \49925 );
and \g133363/U$2 ( \57532 , \56411 , \50159 );
and \g133363/U$3 ( \57533 , \56368 , \50160 );
nor \g133363/U$1 ( \57534 , \57532 , \57533 );
not \g133320/U$4 ( \57535 , \57534 );
or \g133320/U$2 ( \57536 , \57531 , \57535 );
or \g133320/U$5 ( \57537 , \57534 , \49925 );
nand \g133320/U$1 ( \57538 , \57536 , \57537 );
xor \g133087/U$1 ( \57539 , \57530 , \57538 );
not \g133142/U$3 ( \57540 , \49233 );
and \g133156/U$2 ( \57541 , \49405 , \47026 );
and \g133156/U$3 ( \57542 , \56377 , \49403 );
nor \g133156/U$1 ( \57543 , \57541 , \57542 );
not \g133142/U$4 ( \57544 , \57543 );
or \g133142/U$2 ( \57545 , \57540 , \57544 );
or \g133142/U$5 ( \57546 , \57543 , \49233 );
nand \g133142/U$1 ( \57547 , \57545 , \57546 );
xor \g133087/U$1_r1 ( \57548 , \57539 , \57547 );
and \g133032/U$3 ( \57549 , \57518 , \57548 );
and \g133032/U$5 ( \57550 , \57509 , \57517 );
or \g133032/U$2 ( \57551 , \57549 , \57550 );
not \g133321/U$3 ( \57552 , \49925 );
and \g133364/U$2 ( \57553 , \50159 , \56370 );
and \g133364/U$3 ( \57554 , \56379 , \50160 );
nor \g133364/U$1 ( \57555 , \57553 , \57554 );
not \g133321/U$4 ( \57556 , \57555 );
or \g133321/U$2 ( \57557 , \57552 , \57556 );
or \g133321/U$5 ( \57558 , \57555 , \49925 );
nand \g133321/U$1 ( \57559 , \57557 , \57558 );
nand \g133312/U$1 ( \57560 , \47026 , \49812 );
not \g133283/U$3 ( \57561 , \57560 );
not \g133283/U$4 ( \57562 , \49568 );
or \g133283/U$2 ( \57563 , \57561 , \57562 );
or \g133283/U$5 ( \57564 , \49568 , \57560 );
nand \g133283/U$1 ( \57565 , \57563 , \57564 );
and \g133247/U$2 ( \57566 , \49568 , \57565 );
and \g133201/U$2 ( \57567 , \57559 , \57566 );
not \g133386/U$3 ( \57568 , \50362 );
and \g133444/U$2 ( \57569 , \56349 , \50587 );
and \g133444/U$3 ( \57570 , \50588 , \56411 );
nor \g133444/U$1 ( \57571 , \57569 , \57570 );
not \g133386/U$4 ( \57572 , \57571 );
or \g133386/U$2 ( \57573 , \57568 , \57572 );
or \g133386/U$5 ( \57574 , \57571 , \50362 );
nand \g133386/U$1 ( \57575 , \57573 , \57574 );
xor \g133123/U$4 ( \57576 , \57567 , \57575 );
xor \g133180/U$1 ( \57577 , \57500 , \57508 );
and \g133123/U$3 ( \57578 , \57576 , \57577 );
and \g133123/U$5 ( \57579 , \57567 , \57575 );
or \g133123/U$2 ( \57580 , \57578 , \57579 );
not \g133196/U$3 ( \57581 , \50759 );
and \g133234/U$2 ( \57582 , \56357 , \51053 );
and \g133234/U$3 ( \57583 , \51055 , \56359 );
nor \g133234/U$1 ( \57584 , \57582 , \57583 );
not \g133196/U$4 ( \57585 , \57584 );
or \g133196/U$2 ( \57586 , \57581 , \57585 );
or \g133196/U$5 ( \57587 , \57584 , \50759 );
nand \g133196/U$1 ( \57588 , \57586 , \57587 );
xor \g133047/U$4 ( \57589 , \57580 , \57588 );
not \g133092/U$3 ( \57590 , \51124 );
and \g133121/U$2 ( \57591 , \56446 , \51517 );
and \g133121/U$3 ( \57592 , \51518 , \56448 );
nor \g133121/U$1 ( \57593 , \57591 , \57592 );
not \g133092/U$4 ( \57594 , \57593 );
or \g133092/U$2 ( \57595 , \57590 , \57594 );
or \g133092/U$5 ( \57596 , \57593 , \51124 );
nand \g133092/U$1 ( \57597 , \57595 , \57596 );
and \g133047/U$3 ( \57598 , \57589 , \57597 );
and \g133047/U$5 ( \57599 , \57580 , \57588 );
or \g133047/U$2 ( \57600 , \57598 , \57599 );
xor \g132953/U$1 ( \57601 , \57551 , \57600 );
not \g133143/U$3 ( \57602 , \50759 );
and \g133165/U$2 ( \57603 , \56357 , \51055 );
and \g133165/U$3 ( \57604 , \51053 , \56448 );
nor \g133165/U$1 ( \57605 , \57603 , \57604 );
not \g133143/U$4 ( \57606 , \57605 );
or \g133143/U$2 ( \57607 , \57602 , \57606 );
or \g133143/U$5 ( \57608 , \57605 , \50759 );
nand \g133143/U$1 ( \57609 , \57607 , \57608 );
not \g133255/U$3 ( \57610 , \50362 );
and \g133286/U$2 ( \57611 , \56347 , \50588 );
and \g133286/U$3 ( \57612 , \50587 , \56359 );
nor \g133286/U$1 ( \57613 , \57611 , \57612 );
not \g133255/U$4 ( \57614 , \57613 );
or \g133255/U$2 ( \57615 , \57610 , \57614 );
or \g133255/U$5 ( \57616 , \57613 , \50362 );
nand \g133255/U$1 ( \57617 , \57615 , \57616 );
xor \g133031/U$1 ( \57618 , \57609 , \57617 );
xor \g133087/U$4 ( \57619 , \57530 , \57538 );
and \g133087/U$3 ( \57620 , \57619 , \57547 );
and \g133087/U$5 ( \57621 , \57530 , \57538 );
or \g133087/U$2 ( \57622 , \57620 , \57621 );
xor \g133031/U$1_r1 ( \57623 , \57618 , \57622 );
xor \g132953/U$1_r1 ( \57624 , \57601 , \57623 );
and \g133028/U$2 ( \57625 , \56167 , \52273 );
and \g133028/U$3 ( \57626 , \52270 , \55884 );
nor \g133028/U$1 ( \57627 , \57625 , \57626 );
and \g132995/U$2 ( \57628 , \57627 , \51513 );
not \g132995/U$4 ( \57629 , \57627 );
and \g132995/U$3 ( \57630 , \57629 , \51120 );
nor \g132995/U$1 ( \57631 , \57628 , \57630 );
not \g133230/U$3 ( \57632 , \49568 );
and \g133262/U$2 ( \57633 , \49813 , \47026 );
and \g133262/U$3 ( \57634 , \56377 , \49812 );
nor \g133262/U$1 ( \57635 , \57633 , \57634 );
not \g133230/U$4 ( \57636 , \57635 );
or \g133230/U$2 ( \57637 , \57632 , \57636 );
or \g133230/U$5 ( \57638 , \57635 , \49568 );
nand \g133230/U$1 ( \57639 , \57637 , \57638 );
not \g133435/U$3 ( \57640 , \50362 );
and \g133489/U$2 ( \57641 , \56411 , \50587 );
and \g133489/U$3 ( \57642 , \56368 , \50588 );
nor \g133489/U$1 ( \57643 , \57641 , \57642 );
not \g133435/U$4 ( \57644 , \57643 );
or \g133435/U$2 ( \57645 , \57640 , \57644 );
or \g133435/U$5 ( \57646 , \57643 , \50362 );
nand \g133435/U$1 ( \57647 , \57645 , \57646 );
xor \g133127/U$4 ( \57648 , \57639 , \57647 );
xor \g133201/U$1 ( \57649 , \57559 , \57566 );
and \g133127/U$3 ( \57650 , \57648 , \57649 );
and \g133127/U$5 ( \57651 , \57639 , \57647 );
or \g133127/U$2 ( \57652 , \57650 , \57651 );
not \g133258/U$3 ( \57653 , \50759 );
and \g133287/U$2 ( \57654 , \56347 , \51055 );
and \g133287/U$3 ( \57655 , \51053 , \56359 );
nor \g133287/U$1 ( \57656 , \57654 , \57655 );
not \g133258/U$4 ( \57657 , \57656 );
or \g133258/U$2 ( \57658 , \57653 , \57657 );
or \g133258/U$5 ( \57659 , \57656 , \50759 );
nand \g133258/U$1 ( \57660 , \57658 , \57659 );
xor \g133078/U$4 ( \57661 , \57652 , \57660 );
not \g133144/U$3 ( \57662 , \51124 );
and \g133170/U$2 ( \57663 , \56357 , \51518 );
and \g133170/U$3 ( \57664 , \51517 , \56448 );
nor \g133170/U$1 ( \57665 , \57663 , \57664 );
not \g133144/U$4 ( \57666 , \57665 );
or \g133144/U$2 ( \57667 , \57662 , \57666 );
or \g133144/U$5 ( \57668 , \57665 , \51124 );
nand \g133144/U$1 ( \57669 , \57667 , \57668 );
and \g133078/U$3 ( \57670 , \57661 , \57669 );
and \g133078/U$5 ( \57671 , \57652 , \57660 );
or \g133078/U$2 ( \57672 , \57670 , \57671 );
xor \g132954/U$4 ( \57673 , \57631 , \57672 );
xor \g133032/U$1 ( \57674 , \57509 , \57517 );
xor \g133032/U$1_r1 ( \57675 , \57674 , \57548 );
and \g132954/U$3 ( \57676 , \57673 , \57675 );
and \g132954/U$5 ( \57677 , \57631 , \57672 );
or \g132954/U$2 ( \57678 , \57676 , \57677 );
xor \g456168/U$5 ( \57679 , \57624 , \57678 );
and \g133172/U$2 ( \57680 , \57526 , \57529 );
not \g133317/U$3 ( \57681 , \49925 );
and \g133359/U$2 ( \57682 , \56349 , \50159 );
and \g133359/U$3 ( \57683 , \56411 , \50160 );
nor \g133359/U$1 ( \57684 , \57682 , \57683 );
not \g133317/U$4 ( \57685 , \57684 );
or \g133317/U$2 ( \57686 , \57681 , \57685 );
or \g133317/U$5 ( \57687 , \57684 , \49925 );
nand \g133317/U$1 ( \57688 , \57686 , \57687 );
xor \g456169/U$2 ( \57689 , \57680 , \57688 );
not \g133224/U$3 ( \57690 , \49568 );
and \g133266/U$2 ( \57691 , \49812 , \56368 );
and \g133266/U$3 ( \57692 , \56370 , \49813 );
nor \g133266/U$1 ( \57693 , \57691 , \57692 );
not \g133224/U$4 ( \57694 , \57693 );
or \g133224/U$2 ( \57695 , \57690 , \57694 );
or \g133224/U$5 ( \57696 , \57693 , \49568 );
nand \g133224/U$1 ( \57697 , \57695 , \57696 );
not \g133141/U$3 ( \57698 , \49233 );
and \g133158/U$2 ( \57699 , \49405 , \56377 );
and \g133158/U$3 ( \57700 , \56379 , \49403 );
nor \g133158/U$1 ( \57701 , \57699 , \57700 );
not \g133141/U$4 ( \57702 , \57701 );
or \g133141/U$2 ( \57703 , \57698 , \57702 );
or \g133141/U$5 ( \57704 , \57701 , \49233 );
nand \g133141/U$1 ( \57705 , \57703 , \57704 );
xor \g133112/U$1 ( \57706 , \57697 , \57705 );
xor \g456169/U$1 ( \57707 , \57689 , \57706 );
not \g133042/U$3 ( \57708 , \51124 );
and \g133076/U$2 ( \57709 , \56446 , \51518 );
and \g133076/U$3 ( \57710 , \51517 , \56167 );
nor \g133076/U$1 ( \57711 , \57709 , \57710 );
not \g133042/U$4 ( \57712 , \57711 );
or \g133042/U$2 ( \57713 , \57708 , \57712 );
or \g133042/U$5 ( \57714 , \57711 , \51124 );
nand \g133042/U$1 ( \57715 , \57713 , \57714 );
and \g132969/U$2 ( \57716 , \55884 , \52273 );
and \g132969/U$3 ( \57717 , \52270 , \55707 );
nor \g132969/U$1 ( \57718 , \57716 , \57717 );
and \g132934/U$2 ( \57719 , \57718 , \51513 );
not \g132934/U$4 ( \57720 , \57718 );
and \g132934/U$3 ( \57721 , \57720 , \51120 );
nor \g132934/U$1 ( \57722 , \57719 , \57721 );
xor \g456169/U$1_r1 ( \57723 , \57715 , \57722 );
xor \g456169/U$1_r2 ( \57724 , \57707 , \57723 );
and \g456168/U$4 ( \57725 , \57679 , \57724 );
and \g456168/U$6 ( \57726 , \57624 , \57678 );
or \g456168/U$3 ( \57727 , \57725 , \57726 );
not \g133191/U$3 ( \57728 , \50362 );
and \g133235/U$2 ( \57729 , \56357 , \50587 );
and \g133235/U$3 ( \57730 , \50588 , \56359 );
nor \g133235/U$1 ( \57731 , \57729 , \57730 );
not \g133191/U$4 ( \57732 , \57731 );
or \g133191/U$2 ( \57733 , \57728 , \57732 );
or \g133191/U$5 ( \57734 , \57731 , \50362 );
nand \g133191/U$1 ( \57735 , \57733 , \57734 );
not \g133318/U$3 ( \57736 , \49925 );
and \g133365/U$2 ( \57737 , \56347 , \50159 );
and \g133365/U$3 ( \57738 , \56349 , \50160 );
nor \g133365/U$1 ( \57739 , \57737 , \57738 );
not \g133318/U$4 ( \57740 , \57739 );
or \g133318/U$2 ( \57741 , \57736 , \57740 );
or \g133318/U$5 ( \57742 , \57739 , \49925 );
nand \g133318/U$1 ( \57743 , \57741 , \57742 );
xor \g456170/U$2 ( \57744 , \57735 , \57743 );
and \g133112/U$2 ( \57745 , \57697 , \57705 );
xor \g456170/U$1 ( \57746 , \57744 , \57745 );
xor \g133031/U$4 ( \57747 , \57609 , \57617 );
and \g133031/U$3 ( \57748 , \57747 , \57622 );
and \g133031/U$5 ( \57749 , \57609 , \57617 );
or \g133031/U$2 ( \57750 , \57748 , \57749 );
not \g132994/U$3 ( \57751 , \51124 );
and \g133027/U$2 ( \57752 , \56167 , \51518 );
and \g133027/U$3 ( \57753 , \51517 , \55884 );
nor \g133027/U$1 ( \57754 , \57752 , \57753 );
not \g132994/U$4 ( \57755 , \57754 );
or \g132994/U$2 ( \57756 , \57751 , \57755 );
or \g132994/U$5 ( \57757 , \57754 , \51124 );
nand \g132994/U$1 ( \57758 , \57756 , \57757 );
xor \g456170/U$1_r1 ( \57759 , \57750 , \57758 );
xor \g456170/U$1_r2 ( \57760 , \57746 , \57759 );
xor \g132953/U$4 ( \57761 , \57551 , \57600 );
and \g132953/U$3 ( \57762 , \57761 , \57623 );
and \g132953/U$5 ( \57763 , \57551 , \57600 );
or \g132953/U$2 ( \57764 , \57762 , \57763 );
xor \g456165/U$9 ( \57765 , \57760 , \57764 );
and \g132917/U$2 ( \57766 , \55460 , \52270 );
and \g132917/U$3 ( \57767 , \52273 , \55707 );
nor \g132917/U$1 ( \57768 , \57766 , \57767 );
and \g132879/U$2 ( \57769 , \57768 , \51513 );
not \g132879/U$4 ( \57770 , \57768 );
and \g132879/U$3 ( \57771 , \57770 , \51120 );
nor \g132879/U$1 ( \57772 , \57769 , \57771 );
xor \g456169/U$9 ( \57773 , \57680 , \57688 );
xor \g456169/U$9_r1 ( \57774 , \57773 , \57706 );
and \g456169/U$8 ( \57775 , \57715 , \57774 );
xor \g456169/U$11 ( \57776 , \57680 , \57688 );
xor \g456169/U$11_r1 ( \57777 , \57776 , \57706 );
and \g456169/U$10 ( \57778 , \57722 , \57777 );
and \g456169/U$12 ( \57779 , \57715 , \57722 );
or \g456169/U$7 ( \57780 , \57775 , \57778 , \57779 );
xor \g132827/U$1 ( \57781 , \57772 , \57780 );
xor \g456169/U$5 ( \57782 , \57680 , \57688 );
and \g456169/U$4 ( \57783 , \57782 , \57706 );
and \g456169/U$6 ( \57784 , \57680 , \57688 );
or \g456169/U$3 ( \57785 , \57783 , \57784 );
not \g133088/U$3 ( \57786 , \50759 );
and \g133118/U$2 ( \57787 , \56446 , \51053 );
and \g133118/U$3 ( \57788 , \51055 , \56448 );
nor \g133118/U$1 ( \57789 , \57787 , \57788 );
not \g133088/U$4 ( \57790 , \57789 );
or \g133088/U$2 ( \57791 , \57786 , \57790 );
or \g133088/U$5 ( \57792 , \57789 , \50759 );
nand \g133088/U$1 ( \57793 , \57791 , \57792 );
xor \g132919/U$1 ( \57794 , \57785 , \57793 );
not \g133063/U$3 ( \57795 , \49014 );
and \g133096/U$2 ( \57796 , \49075 , \47026 );
and \g133096/U$3 ( \57797 , \56377 , \49074 );
nor \g133096/U$1 ( \57798 , \57796 , \57797 );
not \g133063/U$4 ( \57799 , \57798 );
or \g133063/U$2 ( \57800 , \57795 , \57799 );
or \g133063/U$5 ( \57801 , \57798 , \49014 );
nand \g133063/U$1 ( \57802 , \57800 , \57801 );
not \g133229/U$3 ( \57803 , \49568 );
and \g133269/U$2 ( \57804 , \49812 , \56411 );
and \g133269/U$3 ( \57805 , \56368 , \49813 );
nor \g133269/U$1 ( \57806 , \57804 , \57805 );
not \g133229/U$4 ( \57807 , \57806 );
or \g133229/U$2 ( \57808 , \57803 , \57807 );
or \g133229/U$5 ( \57809 , \57806 , \49568 );
nand \g133229/U$1 ( \57810 , \57808 , \57809 );
xor \g132974/U$1 ( \57811 , \57802 , \57810 );
not \g133135/U$3 ( \57812 , \49233 );
and \g133163/U$2 ( \57813 , \49403 , \56370 );
and \g133163/U$3 ( \57814 , \56379 , \49405 );
nor \g133163/U$1 ( \57815 , \57813 , \57814 );
not \g133135/U$4 ( \57816 , \57815 );
or \g133135/U$2 ( \57817 , \57812 , \57816 );
or \g133135/U$5 ( \57818 , \57815 , \49233 );
nand \g133135/U$1 ( \57819 , \57817 , \57818 );
nand \g133129/U$1 ( \57820 , \47026 , \49074 );
not \g133115/U$3 ( \57821 , \57820 );
not \g133115/U$4 ( \57822 , \49014 );
or \g133115/U$2 ( \57823 , \57821 , \57822 );
or \g133115/U$5 ( \57824 , \49014 , \57820 );
nand \g133115/U$1 ( \57825 , \57823 , \57824 );
and \g133083/U$2 ( \57826 , \49014 , \57825 );
xor \g133049/U$1 ( \57827 , \57819 , \57826 );
xor \g132974/U$1_r1 ( \57828 , \57811 , \57827 );
xor \g132919/U$1_r1 ( \57829 , \57794 , \57828 );
xor \g132827/U$1_r1 ( \57830 , \57781 , \57829 );
xor \g456165/U$9_r1 ( \57831 , \57765 , \57830 );
and \g456165/U$8 ( \57832 , \57727 , \57831 );
not \g133324/U$3 ( \57833 , \50759 );
and \g133362/U$2 ( \57834 , \56347 , \51053 );
and \g133362/U$3 ( \57835 , \51055 , \56349 );
nor \g133362/U$1 ( \57836 , \57834 , \57835 );
not \g133324/U$4 ( \57837 , \57836 );
or \g133324/U$2 ( \57838 , \57833 , \57837 );
or \g133324/U$5 ( \57839 , \57836 , \50759 );
nand \g133324/U$1 ( \57840 , \57838 , \57839 );
not \g133436/U$3 ( \57841 , \50362 );
and \g133492/U$2 ( \57842 , \56368 , \50587 );
and \g133492/U$3 ( \57843 , \56370 , \50588 );
nor \g133492/U$1 ( \57844 , \57842 , \57843 );
not \g133436/U$4 ( \57845 , \57844 );
or \g133436/U$2 ( \57846 , \57841 , \57845 );
or \g133436/U$5 ( \57847 , \57844 , \50362 );
nand \g133436/U$1 ( \57848 , \57846 , \57847 );
not \g133314/U$3 ( \57849 , \49925 );
and \g133360/U$2 ( \57850 , \50160 , \56377 );
and \g133360/U$3 ( \57851 , \56379 , \50159 );
nor \g133360/U$1 ( \57852 , \57850 , \57851 );
not \g133314/U$4 ( \57853 , \57852 );
or \g133314/U$2 ( \57854 , \57849 , \57853 );
or \g133314/U$5 ( \57855 , \57852 , \49925 );
nand \g133314/U$1 ( \57856 , \57854 , \57855 );
and \g133280/U$2 ( \57857 , \57848 , \57856 );
xor \g456171/U$5 ( \57858 , \57840 , \57857 );
xor \g133127/U$1 ( \57859 , \57639 , \57647 );
xor \g133127/U$1_r1 ( \57860 , \57859 , \57649 );
and \g456171/U$4 ( \57861 , \57858 , \57860 );
and \g456171/U$6 ( \57862 , \57840 , \57857 );
or \g456171/U$3 ( \57863 , \57861 , \57862 );
xor \g133123/U$1 ( \57864 , \57567 , \57575 );
xor \g133123/U$1_r1 ( \57865 , \57864 , \57577 );
xor \g133001/U$4 ( \57866 , \57863 , \57865 );
and \g133077/U$2 ( \57867 , \56446 , \52273 );
and \g133077/U$3 ( \57868 , \52270 , \56167 );
nor \g133077/U$1 ( \57869 , \57867 , \57868 );
and \g133044/U$2 ( \57870 , \57869 , \51513 );
not \g133044/U$4 ( \57871 , \57869 );
and \g133044/U$3 ( \57872 , \57871 , \51120 );
nor \g133044/U$1 ( \57873 , \57870 , \57872 );
and \g133001/U$3 ( \57874 , \57866 , \57873 );
and \g133001/U$5 ( \57875 , \57863 , \57865 );
or \g133001/U$2 ( \57876 , \57874 , \57875 );
xor \g133047/U$1 ( \57877 , \57580 , \57588 );
xor \g133047/U$1_r1 ( \57878 , \57877 , \57597 );
xor \g132869/U$4 ( \57879 , \57876 , \57878 );
xor \g132954/U$1 ( \57880 , \57631 , \57672 );
xor \g132954/U$1_r1 ( \57881 , \57880 , \57675 );
and \g132869/U$3 ( \57882 , \57879 , \57881 );
and \g132869/U$5 ( \57883 , \57876 , \57878 );
or \g132869/U$2 ( \57884 , \57882 , \57883 );
xor \g456168/U$9 ( \57885 , \57624 , \57678 );
xor \g456168/U$9_r1 ( \57886 , \57885 , \57724 );
and \g456168/U$8 ( \57887 , \57884 , \57886 );
not \g133434/U$3 ( \57888 , \50362 );
and \g133490/U$2 ( \57889 , \50587 , \56379 );
and \g133490/U$3 ( \57890 , \56377 , \50588 );
nor \g133490/U$1 ( \57891 , \57889 , \57890 );
not \g133434/U$4 ( \57892 , \57891 );
or \g133434/U$2 ( \57893 , \57888 , \57892 );
or \g133434/U$5 ( \57894 , \57891 , \50362 );
nand \g133434/U$1 ( \57895 , \57893 , \57894 );
nand \g133592/U$1 ( \57896 , \47026 , \50587 );
not \g133527/U$3 ( \57897 , \57896 );
not \g133527/U$4 ( \57898 , \50362 );
or \g133527/U$2 ( \57899 , \57897 , \57898 );
or \g133527/U$5 ( \57900 , \50362 , \57896 );
nand \g133527/U$1 ( \57901 , \57899 , \57900 );
and \g133478/U$2 ( \57902 , \50362 , \57901 );
not \g133438/U$3 ( \57903 , \50362 );
and \g133488/U$2 ( \57904 , \50588 , \47026 );
and \g133488/U$3 ( \57905 , \56377 , \50587 );
nor \g133488/U$1 ( \57906 , \57904 , \57905 );
not \g133438/U$4 ( \57907 , \57906 );
or \g133438/U$2 ( \57908 , \57903 , \57907 );
or \g133438/U$5 ( \57909 , \57906 , \50362 );
nand \g133438/U$1 ( \57910 , \57908 , \57909 );
and \g133384/U$2 ( \57911 , \57902 , \57910 );
xor \g133333/U$1 ( \57912 , \57895 , \57911 );
not \g133596/U$3 ( \57913 , \50759 );
and \g133650/U$2 ( \57914 , \56368 , \51053 );
and \g133650/U$3 ( \57915 , \51055 , \56370 );
nor \g133650/U$1 ( \57916 , \57914 , \57915 );
not \g133596/U$4 ( \57917 , \57916 );
or \g133596/U$2 ( \57918 , \57913 , \57917 );
or \g133596/U$5 ( \57919 , \57916 , \50759 );
nand \g133596/U$1 ( \57920 , \57918 , \57919 );
xor \g133238/U$1 ( \57921 , \57912 , \57920 );
not \g133387/U$3 ( \57922 , \51124 );
and \g133448/U$2 ( \57923 , \56349 , \51517 );
and \g133448/U$3 ( \57924 , \51518 , \56411 );
nor \g133448/U$1 ( \57925 , \57923 , \57924 );
not \g133387/U$4 ( \57926 , \57925 );
or \g133387/U$2 ( \57927 , \57922 , \57926 );
or \g133387/U$5 ( \57928 , \57925 , \51124 );
nand \g133387/U$1 ( \57929 , \57927 , \57928 );
xor \g133238/U$1_r1 ( \57930 , \57921 , \57929 );
xor \g133384/U$1 ( \57931 , \57902 , \57910 );
not \g133595/U$3 ( \57932 , \50759 );
and \g133648/U$2 ( \57933 , \56370 , \51053 );
and \g133648/U$3 ( \57934 , \56379 , \51055 );
nor \g133648/U$1 ( \57935 , \57933 , \57934 );
not \g133595/U$4 ( \57936 , \57935 );
or \g133595/U$2 ( \57937 , \57932 , \57936 );
or \g133595/U$5 ( \57938 , \57935 , \50759 );
nand \g133595/U$1 ( \57939 , \57937 , \57938 );
xor \g456175/U$5 ( \57940 , \57931 , \57939 );
not \g133484/U$3 ( \57941 , \51124 );
and \g133533/U$2 ( \57942 , \56411 , \51517 );
and \g133533/U$3 ( \57943 , \51518 , \56368 );
nor \g133533/U$1 ( \57944 , \57942 , \57943 );
not \g133484/U$4 ( \57945 , \57944 );
or \g133484/U$2 ( \57946 , \57941 , \57945 );
or \g133484/U$5 ( \57947 , \57944 , \51124 );
nand \g133484/U$1 ( \57948 , \57946 , \57947 );
and \g456175/U$4 ( \57949 , \57940 , \57948 );
and \g456175/U$6 ( \57950 , \57931 , \57939 );
or \g456175/U$3 ( \57951 , \57949 , \57950 );
xor \g456173/U$5 ( \57952 , \57930 , \57951 );
and \g133289/U$2 ( \57953 , \56347 , \52273 );
and \g133289/U$3 ( \57954 , \52270 , \56359 );
nor \g133289/U$1 ( \57955 , \57953 , \57954 );
and \g133257/U$2 ( \57956 , \57955 , \51513 );
not \g133257/U$4 ( \57957 , \57955 );
and \g133257/U$3 ( \57958 , \57957 , \51120 );
nor \g133257/U$1 ( \57959 , \57956 , \57958 );
and \g456173/U$4 ( \57960 , \57952 , \57959 );
and \g456173/U$6 ( \57961 , \57930 , \57951 );
or \g456173/U$3 ( \57962 , \57960 , \57961 );
not \g133483/U$3 ( \57963 , \50759 );
and \g133531/U$2 ( \57964 , \56411 , \51053 );
and \g133531/U$3 ( \57965 , \51055 , \56368 );
nor \g133531/U$1 ( \57966 , \57964 , \57965 );
not \g133483/U$4 ( \57967 , \57966 );
or \g133483/U$2 ( \57968 , \57963 , \57967 );
or \g133483/U$5 ( \57969 , \57966 , \50759 );
nand \g133483/U$1 ( \57970 , \57968 , \57969 );
not \g133437/U$3 ( \57971 , \50362 );
and \g133491/U$2 ( \57972 , \56370 , \50587 );
and \g133491/U$3 ( \57973 , \56379 , \50588 );
nor \g133491/U$1 ( \57974 , \57972 , \57973 );
not \g133437/U$4 ( \57975 , \57974 );
or \g133437/U$2 ( \57976 , \57971 , \57975 );
or \g133437/U$5 ( \57977 , \57974 , \50362 );
nand \g133437/U$1 ( \57978 , \57976 , \57977 );
xor \g133199/U$1 ( \57979 , \57970 , \57978 );
nand \g133431/U$1 ( \57980 , \47026 , \50159 );
not \g133391/U$3 ( \57981 , \57980 );
not \g133391/U$4 ( \57982 , \49925 );
or \g133391/U$2 ( \57983 , \57981 , \57982 );
or \g133391/U$5 ( \57984 , \49925 , \57980 );
nand \g133391/U$1 ( \57985 , \57983 , \57984 );
and \g133348/U$2 ( \57986 , \49925 , \57985 );
not \g133316/U$3 ( \57987 , \49925 );
and \g133358/U$2 ( \57988 , \50160 , \47026 );
and \g133358/U$3 ( \57989 , \56377 , \50159 );
nor \g133358/U$1 ( \57990 , \57988 , \57989 );
not \g133316/U$4 ( \57991 , \57990 );
or \g133316/U$2 ( \57992 , \57987 , \57991 );
or \g133316/U$5 ( \57993 , \57990 , \49925 );
nand \g133316/U$1 ( \57994 , \57992 , \57993 );
xor \g133279/U$1 ( \57995 , \57986 , \57994 );
xor \g133199/U$1_r1 ( \57996 , \57979 , \57995 );
xor \g133238/U$4 ( \57997 , \57912 , \57920 );
and \g133238/U$3 ( \57998 , \57997 , \57929 );
and \g133238/U$5 ( \57999 , \57912 , \57920 );
or \g133238/U$2 ( \58000 , \57998 , \57999 );
and \g133333/U$2 ( \58001 , \57895 , \57911 );
xor \g133153/U$1 ( \58002 , \58000 , \58001 );
not \g133322/U$3 ( \58003 , \51124 );
and \g133367/U$2 ( \58004 , \56347 , \51517 );
and \g133367/U$3 ( \58005 , \51518 , \56349 );
nor \g133367/U$1 ( \58006 , \58004 , \58005 );
not \g133322/U$4 ( \58007 , \58006 );
or \g133322/U$2 ( \58008 , \58003 , \58007 );
or \g133322/U$5 ( \58009 , \58006 , \51124 );
nand \g133322/U$1 ( \58010 , \58008 , \58009 );
xor \g133153/U$1_r1 ( \58011 , \58002 , \58010 );
xor \g456172/U$9 ( \58012 , \57996 , \58011 );
and \g133237/U$2 ( \58013 , \56357 , \52270 );
and \g133237/U$3 ( \58014 , \52273 , \56359 );
nor \g133237/U$1 ( \58015 , \58013 , \58014 );
and \g133193/U$2 ( \58016 , \58015 , \51513 );
not \g133193/U$4 ( \58017 , \58015 );
and \g133193/U$3 ( \58018 , \58017 , \51120 );
nor \g133193/U$1 ( \58019 , \58016 , \58018 );
xor \g456172/U$9_r1 ( \58020 , \58012 , \58019 );
and \g456172/U$8 ( \58021 , \57962 , \58020 );
not \g133598/U$3 ( \58022 , \50759 );
and \g133649/U$2 ( \58023 , \56379 , \51053 );
and \g133649/U$3 ( \58024 , \56377 , \51055 );
nor \g133649/U$1 ( \58025 , \58023 , \58024 );
not \g133598/U$4 ( \58026 , \58025 );
or \g133598/U$2 ( \58027 , \58022 , \58026 );
or \g133598/U$5 ( \58028 , \58025 , \50759 );
nand \g133598/U$1 ( \58029 , \58027 , \58028 );
not \g135560/U$2 ( \58030 , \50759 );
nor \g133813/U$1 ( \58031 , \51054 , \47025 );
nor \g135560/U$1 ( \58032 , \58030 , \58031 );
not \g133597/U$3 ( \58033 , \50759 );
and \g133647/U$2 ( \58034 , \51055 , \47026 );
and \g133647/U$3 ( \58035 , \56377 , \51053 );
nor \g133647/U$1 ( \58036 , \58034 , \58035 );
not \g133597/U$4 ( \58037 , \58036 );
or \g133597/U$2 ( \58038 , \58033 , \58037 );
or \g133597/U$5 ( \58039 , \58036 , \50759 );
nand \g133597/U$1 ( \58040 , \58038 , \58039 );
and \g133511/U$2 ( \58041 , \58032 , \58040 );
and \g133453/U$2 ( \58042 , \58029 , \58041 );
xor \g456175/U$9 ( \58043 , \57931 , \57939 );
xor \g456175/U$9_r1 ( \58044 , \58043 , \57948 );
and \g456175/U$8 ( \58045 , \58042 , \58044 );
and \g133368/U$2 ( \58046 , \56347 , \52270 );
and \g133368/U$3 ( \58047 , \52273 , \56349 );
nor \g133368/U$1 ( \58048 , \58046 , \58047 );
and \g133319/U$2 ( \58049 , \58048 , \51513 );
not \g133319/U$4 ( \58050 , \58048 );
and \g133319/U$3 ( \58051 , \58050 , \51120 );
nor \g133319/U$1 ( \58052 , \58049 , \58051 );
xor \g456175/U$11 ( \58053 , \57931 , \57939 );
xor \g456175/U$11_r1 ( \58054 , \58053 , \57948 );
and \g456175/U$10 ( \58055 , \58052 , \58054 );
and \g456175/U$12 ( \58056 , \58042 , \58052 );
or \g456175/U$7 ( \58057 , \58045 , \58055 , \58056 );
xor \g456173/U$9 ( \58058 , \57930 , \57951 );
xor \g456173/U$9_r1 ( \58059 , \58058 , \57959 );
and \g456173/U$8 ( \58060 , \58057 , \58059 );
and \g133836/U$2 ( \58061 , \56377 , \52270 );
and \g133939/U$2 ( \58062 , \56379 , \52270 );
and \g133939/U$3 ( \58063 , \52273 , \56377 );
nor \g133939/U$1 ( \58064 , \58062 , \58063 );
and \g133868/U$2 ( \58065 , \58064 , \51120 );
not \g133868/U$4 ( \58066 , \58064 );
and \g133868/U$3 ( \58067 , \58066 , \51513 );
nor \g133868/U$1 ( \58068 , \58065 , \58067 );
nor \g133836/U$1 ( \58069 , \58061 , \58068 );
not \g135561/U$2 ( \58070 , \58069 );
nor \g135561/U$1 ( \58071 , \58070 , \47026 , \51513 );
nand \g134084/U$1 ( \58072 , \47026 , \51517 );
and \g134061/U$1 ( \58073 , \51124 , \58072 );
not \g133822/U$3 ( \58074 , \51124 );
and \g133873/U$2 ( \58075 , \51518 , \47026 );
and \g133873/U$3 ( \58076 , \51517 , \56377 );
nor \g133873/U$1 ( \58077 , \58075 , \58076 );
not \g133822/U$4 ( \58078 , \58077 );
or \g133822/U$2 ( \58079 , \58074 , \58078 );
or \g133822/U$5 ( \58080 , \58077 , \51124 );
nand \g133822/U$1 ( \58081 , \58079 , \58080 );
xor \g133676/U$1 ( \58082 , \58073 , \58081 );
xor \g133537/U$4 ( \58083 , \58071 , \58082 );
and \g133826/U$2 ( \58084 , \56370 , \52270 );
and \g133826/U$3 ( \58085 , \52273 , \56379 );
nor \g133826/U$1 ( \58086 , \58084 , \58085 );
and \g133697/U$2 ( \58087 , \58086 , \51513 );
not \g133697/U$4 ( \58088 , \58086 );
and \g133697/U$3 ( \58089 , \58088 , \51120 );
nor \g133697/U$1 ( \58090 , \58087 , \58089 );
and \g133537/U$3 ( \58091 , \58083 , \58090 );
and \g133537/U$5 ( \58092 , \58071 , \58082 );
or \g133537/U$2 ( \58093 , \58091 , \58092 );
not \g133821/U$3 ( \58094 , \51124 );
and \g133874/U$2 ( \58095 , \56379 , \51517 );
and \g133874/U$3 ( \58096 , \56377 , \51518 );
nor \g133874/U$1 ( \58097 , \58095 , \58096 );
not \g133821/U$4 ( \58098 , \58097 );
or \g133821/U$2 ( \58099 , \58094 , \58098 );
or \g133821/U$5 ( \58100 , \58097 , \51124 );
nand \g133821/U$1 ( \58101 , \58099 , \58100 );
and \g133676/U$2 ( \58102 , \58073 , \58081 );
xor \g133611/U$1 ( \58103 , \58101 , \58102 );
xor \g133396/U$4 ( \58104 , \58093 , \58103 );
and \g133652/U$2 ( \58105 , \56368 , \52270 );
and \g133652/U$3 ( \58106 , \52273 , \56370 );
nor \g133652/U$1 ( \58107 , \58105 , \58106 );
and \g133599/U$2 ( \58108 , \58107 , \51513 );
not \g133599/U$4 ( \58109 , \58107 );
and \g133599/U$3 ( \58110 , \58109 , \51120 );
nor \g133599/U$1 ( \58111 , \58108 , \58110 );
and \g133396/U$3 ( \58112 , \58104 , \58111 );
and \g133396/U$5 ( \58113 , \58093 , \58103 );
or \g133396/U$2 ( \58114 , \58112 , \58113 );
and \g133611/U$2 ( \58115 , \58101 , \58102 );
xor \g133291/U$4 ( \58116 , \58114 , \58115 );
xor \g133511/U$1 ( \58117 , \58032 , \58040 );
not \g133696/U$3 ( \58118 , \51124 );
and \g133824/U$2 ( \58119 , \56370 , \51517 );
and \g133824/U$3 ( \58120 , \51518 , \56379 );
nor \g133824/U$1 ( \58121 , \58119 , \58120 );
not \g133696/U$4 ( \58122 , \58121 );
or \g133696/U$2 ( \58123 , \58118 , \58122 );
or \g133696/U$5 ( \58124 , \58121 , \51124 );
nand \g133696/U$1 ( \58125 , \58123 , \58124 );
xor \g133382/U$1 ( \58126 , \58117 , \58125 );
and \g133534/U$2 ( \58127 , \56411 , \52270 );
and \g133534/U$3 ( \58128 , \52273 , \56368 );
nor \g133534/U$1 ( \58129 , \58127 , \58128 );
and \g133485/U$2 ( \58130 , \58129 , \51513 );
not \g133485/U$4 ( \58131 , \58129 );
and \g133485/U$3 ( \58132 , \58131 , \51120 );
nor \g133485/U$1 ( \58133 , \58130 , \58132 );
xor \g133382/U$1_r1 ( \58134 , \58126 , \58133 );
and \g133291/U$3 ( \58135 , \58116 , \58134 );
and \g133291/U$5 ( \58136 , \58114 , \58115 );
or \g133291/U$2 ( \58137 , \58135 , \58136 );
xor \g133382/U$4 ( \58138 , \58117 , \58125 );
and \g133382/U$3 ( \58139 , \58138 , \58133 );
and \g133382/U$5 ( \58140 , \58117 , \58125 );
or \g133382/U$2 ( \58141 , \58139 , \58140 );
xor \g133213/U$4 ( \58142 , \58137 , \58141 );
not \g133600/U$3 ( \58143 , \51124 );
and \g133651/U$2 ( \58144 , \56368 , \51517 );
and \g133651/U$3 ( \58145 , \51518 , \56370 );
nor \g133651/U$1 ( \58146 , \58144 , \58145 );
not \g133600/U$4 ( \58147 , \58146 );
or \g133600/U$2 ( \58148 , \58143 , \58147 );
or \g133600/U$5 ( \58149 , \58146 , \51124 );
nand \g133600/U$1 ( \58150 , \58148 , \58149 );
xor \g133453/U$1 ( \58151 , \58029 , \58041 );
xor \g133334/U$1 ( \58152 , \58150 , \58151 );
and \g133449/U$2 ( \58153 , \56349 , \52270 );
and \g133449/U$3 ( \58154 , \52273 , \56411 );
nor \g133449/U$1 ( \58155 , \58153 , \58154 );
and \g133389/U$2 ( \58156 , \58155 , \51513 );
not \g133389/U$4 ( \58157 , \58155 );
and \g133389/U$3 ( \58158 , \58157 , \51120 );
nor \g133389/U$1 ( \58159 , \58156 , \58158 );
xor \g133334/U$1_r1 ( \58160 , \58152 , \58159 );
and \g133213/U$3 ( \58161 , \58142 , \58160 );
and \g133213/U$5 ( \58162 , \58137 , \58141 );
or \g133213/U$2 ( \58163 , \58161 , \58162 );
xor \g133334/U$4 ( \58164 , \58150 , \58151 );
and \g133334/U$3 ( \58165 , \58164 , \58159 );
and \g133334/U$5 ( \58166 , \58150 , \58151 );
or \g133334/U$2 ( \58167 , \58165 , \58166 );
xor \g133128/U$4 ( \58168 , \58163 , \58167 );
xor \g456175/U$2 ( \58169 , \57931 , \57939 );
xor \g456175/U$1 ( \58170 , \58169 , \57948 );
xor \g456175/U$1_r1 ( \58171 , \58042 , \58052 );
xor \g456175/U$1_r2 ( \58172 , \58170 , \58171 );
and \g133128/U$3 ( \58173 , \58168 , \58172 );
and \g133128/U$5 ( \58174 , \58163 , \58167 );
or \g133128/U$2 ( \58175 , \58173 , \58174 );
xor \g456173/U$11 ( \58176 , \57930 , \57951 );
xor \g456173/U$11_r1 ( \58177 , \58176 , \57959 );
and \g456173/U$10 ( \58178 , \58175 , \58177 );
and \g456173/U$12 ( \58179 , \58057 , \58175 );
or \g456173/U$7 ( \58180 , \58060 , \58178 , \58179 );
xor \g456172/U$11 ( \58181 , \57996 , \58011 );
xor \g456172/U$11_r1 ( \58182 , \58181 , \58019 );
and \g456172/U$10 ( \58183 , \58180 , \58182 );
and \g456172/U$12 ( \58184 , \57962 , \58180 );
or \g456172/U$7 ( \58185 , \58021 , \58183 , \58184 );
xor \g456172/U$5 ( \58186 , \57996 , \58011 );
and \g456172/U$4 ( \58187 , \58186 , \58019 );
and \g456172/U$6 ( \58188 , \57996 , \58011 );
or \g456172/U$3 ( \58189 , \58187 , \58188 );
xor \g132976/U$4 ( \58190 , \58185 , \58189 );
and \g133279/U$2 ( \58191 , \57986 , \57994 );
not \g133388/U$3 ( \58192 , \50759 );
and \g133445/U$2 ( \58193 , \56349 , \51053 );
and \g133445/U$3 ( \58194 , \51055 , \56411 );
nor \g133445/U$1 ( \58195 , \58193 , \58194 );
not \g133388/U$4 ( \58196 , \58195 );
or \g133388/U$2 ( \58197 , \58192 , \58196 );
or \g133388/U$5 ( \58198 , \58195 , \50759 );
nand \g133388/U$1 ( \58199 , \58197 , \58198 );
xor \g456174/U$2 ( \58200 , \58191 , \58199 );
xor \g133280/U$1 ( \58201 , \57848 , \57856 );
xor \g456174/U$1 ( \58202 , \58200 , \58201 );
xor \g133153/U$4 ( \58203 , \58000 , \58001 );
and \g133153/U$3 ( \58204 , \58203 , \58010 );
and \g133153/U$5 ( \58205 , \58000 , \58001 );
or \g133153/U$2 ( \58206 , \58204 , \58205 );
not \g133256/U$3 ( \58207 , \51124 );
and \g133288/U$2 ( \58208 , \56347 , \51518 );
and \g133288/U$3 ( \58209 , \51517 , \56359 );
nor \g133288/U$1 ( \58210 , \58208 , \58209 );
not \g133256/U$4 ( \58211 , \58210 );
or \g133256/U$2 ( \58212 , \58207 , \58211 );
or \g133256/U$5 ( \58213 , \58210 , \51124 );
nand \g133256/U$1 ( \58214 , \58212 , \58213 );
xor \g133199/U$4 ( \58215 , \57970 , \57978 );
and \g133199/U$3 ( \58216 , \58215 , \57995 );
and \g133199/U$5 ( \58217 , \57970 , \57978 );
or \g133199/U$2 ( \58218 , \58216 , \58217 );
xor \g133113/U$1 ( \58219 , \58214 , \58218 );
and \g133171/U$2 ( \58220 , \56357 , \52273 );
and \g133171/U$3 ( \58221 , \52270 , \56448 );
nor \g133171/U$1 ( \58222 , \58220 , \58221 );
and \g133145/U$2 ( \58223 , \58222 , \51513 );
not \g133145/U$4 ( \58224 , \58222 );
and \g133145/U$3 ( \58225 , \58224 , \51120 );
nor \g133145/U$1 ( \58226 , \58223 , \58225 );
xor \g133113/U$1_r1 ( \58227 , \58219 , \58226 );
xor \g456174/U$1_r1 ( \58228 , \58206 , \58227 );
xor \g456174/U$1_r2 ( \58229 , \58202 , \58228 );
and \g132976/U$3 ( \58230 , \58190 , \58229 );
and \g132976/U$5 ( \58231 , \58185 , \58189 );
or \g132976/U$2 ( \58232 , \58230 , \58231 );
xor \g456174/U$9 ( \58233 , \58191 , \58199 );
xor \g456174/U$9_r1 ( \58234 , \58233 , \58201 );
and \g456174/U$8 ( \58235 , \58206 , \58234 );
xor \g456174/U$11 ( \58236 , \58191 , \58199 );
xor \g456174/U$11_r1 ( \58237 , \58236 , \58201 );
and \g456174/U$10 ( \58238 , \58227 , \58237 );
and \g456174/U$12 ( \58239 , \58206 , \58227 );
or \g456174/U$7 ( \58240 , \58235 , \58238 , \58239 );
xor \g132920/U$4 ( \58241 , \58232 , \58240 );
xor \g456171/U$2 ( \58242 , \57840 , \57857 );
xor \g456171/U$1 ( \58243 , \58242 , \57860 );
xor \g133113/U$4 ( \58244 , \58214 , \58218 );
and \g133113/U$3 ( \58245 , \58244 , \58226 );
and \g133113/U$5 ( \58246 , \58214 , \58218 );
or \g133113/U$2 ( \58247 , \58245 , \58246 );
not \g133192/U$3 ( \58248 , \51124 );
and \g133236/U$2 ( \58249 , \56357 , \51517 );
and \g133236/U$3 ( \58250 , \51518 , \56359 );
nor \g133236/U$1 ( \58251 , \58249 , \58250 );
not \g133192/U$4 ( \58252 , \58251 );
or \g133192/U$2 ( \58253 , \58248 , \58252 );
or \g133192/U$5 ( \58254 , \58251 , \51124 );
nand \g133192/U$1 ( \58255 , \58253 , \58254 );
xor \g456174/U$5 ( \58256 , \58191 , \58199 );
and \g456174/U$4 ( \58257 , \58256 , \58201 );
and \g456174/U$6 ( \58258 , \58191 , \58199 );
or \g456174/U$3 ( \58259 , \58257 , \58258 );
xor \g133055/U$1 ( \58260 , \58255 , \58259 );
and \g133122/U$2 ( \58261 , \56446 , \52270 );
and \g133122/U$3 ( \58262 , \52273 , \56448 );
nor \g133122/U$1 ( \58263 , \58261 , \58262 );
and \g133093/U$2 ( \58264 , \58263 , \51513 );
not \g133093/U$4 ( \58265 , \58263 );
and \g133093/U$3 ( \58266 , \58265 , \51120 );
nor \g133093/U$1 ( \58267 , \58264 , \58266 );
xor \g133055/U$1_r1 ( \58268 , \58260 , \58267 );
xor \g456171/U$1_r1 ( \58269 , \58247 , \58268 );
xor \g456171/U$1_r2 ( \58270 , \58243 , \58269 );
and \g132920/U$3 ( \58271 , \58241 , \58270 );
and \g132920/U$5 ( \58272 , \58232 , \58240 );
or \g132920/U$2 ( \58273 , \58271 , \58272 );
xor \g456171/U$9 ( \58274 , \57840 , \57857 );
xor \g456171/U$9_r1 ( \58275 , \58274 , \57860 );
and \g456171/U$8 ( \58276 , \58247 , \58275 );
xor \g456171/U$11 ( \58277 , \57840 , \57857 );
xor \g456171/U$11_r1 ( \58278 , \58277 , \57860 );
and \g456171/U$10 ( \58279 , \58268 , \58278 );
and \g456171/U$12 ( \58280 , \58247 , \58268 );
or \g456171/U$7 ( \58281 , \58276 , \58279 , \58280 );
xor \g132864/U$4 ( \58282 , \58273 , \58281 );
xor \g133055/U$4 ( \58283 , \58255 , \58259 );
and \g133055/U$3 ( \58284 , \58283 , \58267 );
and \g133055/U$5 ( \58285 , \58255 , \58259 );
or \g133055/U$2 ( \58286 , \58284 , \58285 );
xor \g133078/U$1 ( \58287 , \57652 , \57660 );
xor \g133078/U$1_r1 ( \58288 , \58287 , \57669 );
xor \g132926/U$1 ( \58289 , \58286 , \58288 );
xor \g133001/U$1 ( \58290 , \57863 , \57865 );
xor \g133001/U$1_r1 ( \58291 , \58290 , \57873 );
xor \g132926/U$1_r1 ( \58292 , \58289 , \58291 );
and \g132864/U$3 ( \58293 , \58282 , \58292 );
and \g132864/U$5 ( \58294 , \58273 , \58281 );
or \g132864/U$2 ( \58295 , \58293 , \58294 );
xor \g132926/U$4 ( \58296 , \58286 , \58288 );
and \g132926/U$3 ( \58297 , \58296 , \58291 );
and \g132926/U$5 ( \58298 , \58286 , \58288 );
or \g132926/U$2 ( \58299 , \58297 , \58298 );
xor \g132790/U$4 ( \58300 , \58295 , \58299 );
xor \g132869/U$1 ( \58301 , \57876 , \57878 );
xor \g132869/U$1_r1 ( \58302 , \58301 , \57881 );
and \g132790/U$3 ( \58303 , \58300 , \58302 );
and \g132790/U$5 ( \58304 , \58295 , \58299 );
or \g132790/U$2 ( \58305 , \58303 , \58304 );
xor \g456168/U$11 ( \58306 , \57624 , \57678 );
xor \g456168/U$11_r1 ( \58307 , \58306 , \57724 );
and \g456168/U$10 ( \58308 , \58305 , \58307 );
and \g456168/U$12 ( \58309 , \57884 , \58305 );
or \g456168/U$7 ( \58310 , \57887 , \58308 , \58309 );
xor \g456165/U$11 ( \58311 , \57760 , \57764 );
xor \g456165/U$11_r1 ( \58312 , \58311 , \57830 );
and \g456165/U$10 ( \58313 , \58310 , \58312 );
and \g456165/U$12 ( \58314 , \57727 , \58310 );
or \g456165/U$7 ( \58315 , \57832 , \58313 , \58314 );
xor \g456165/U$5 ( \58316 , \57760 , \57764 );
and \g456165/U$4 ( \58317 , \58316 , \57830 );
and \g456165/U$6 ( \58318 , \57760 , \57764 );
or \g456165/U$3 ( \58319 , \58317 , \58318 );
xor \g132518/U$4 ( \58320 , \58315 , \58319 );
not \g133136/U$3 ( \58321 , \50362 );
and \g133160/U$2 ( \58322 , \56357 , \50588 );
and \g133160/U$3 ( \58323 , \50587 , \56448 );
nor \g133160/U$1 ( \58324 , \58322 , \58323 );
not \g133136/U$4 ( \58325 , \58324 );
or \g133136/U$2 ( \58326 , \58321 , \58325 );
or \g133136/U$5 ( \58327 , \58324 , \50362 );
nand \g133136/U$1 ( \58328 , \58326 , \58327 );
not \g133254/U$3 ( \58329 , \49925 );
and \g133285/U$2 ( \58330 , \56347 , \50160 );
and \g133285/U$3 ( \58331 , \50159 , \56359 );
nor \g133285/U$1 ( \58332 , \58330 , \58331 );
not \g133254/U$4 ( \58333 , \58332 );
or \g133254/U$2 ( \58334 , \58329 , \58333 );
or \g133254/U$5 ( \58335 , \58332 , \49925 );
nand \g133254/U$1 ( \58336 , \58334 , \58335 );
xor \g132918/U$1 ( \58337 , \58328 , \58336 );
xor \g132974/U$4 ( \58338 , \57802 , \57810 );
and \g132974/U$3 ( \58339 , \58338 , \57827 );
and \g132974/U$5 ( \58340 , \57802 , \57810 );
or \g132974/U$2 ( \58341 , \58339 , \58340 );
xor \g132918/U$1_r1 ( \58342 , \58337 , \58341 );
not \g132932/U$3 ( \58343 , \51124 );
and \g132968/U$2 ( \58344 , \55884 , \51518 );
and \g132968/U$3 ( \58345 , \51517 , \55707 );
nor \g132968/U$1 ( \58346 , \58344 , \58345 );
not \g132932/U$4 ( \58347 , \58346 );
or \g132932/U$2 ( \58348 , \58343 , \58347 );
or \g132932/U$5 ( \58349 , \58346 , \51124 );
nand \g132932/U$1 ( \58350 , \58348 , \58349 );
xor \g456167/U$2 ( \58351 , \58342 , \58350 );
and \g132862/U$2 ( \58352 , \55127 , \52270 );
and \g132862/U$3 ( \58353 , \52273 , \55460 );
nor \g132862/U$1 ( \58354 , \58352 , \58353 );
and \g132812/U$2 ( \58355 , \58354 , \51513 );
not \g132812/U$4 ( \58356 , \58354 );
and \g132812/U$3 ( \58357 , \58356 , \51120 );
nor \g132812/U$1 ( \58358 , \58355 , \58357 );
xor \g456167/U$1 ( \58359 , \58351 , \58358 );
xor \g132827/U$4 ( \58360 , \57772 , \57780 );
and \g132827/U$3 ( \58361 , \58360 , \57829 );
and \g132827/U$5 ( \58362 , \57772 , \57780 );
or \g132827/U$2 ( \58363 , \58361 , \58362 );
xor \g132919/U$4 ( \58364 , \57785 , \57793 );
and \g132919/U$3 ( \58365 , \58364 , \57828 );
and \g132919/U$5 ( \58366 , \57785 , \57793 );
or \g132919/U$2 ( \58367 , \58365 , \58366 );
xor \g456170/U$9 ( \58368 , \57735 , \57743 );
xor \g456170/U$9_r1 ( \58369 , \58368 , \57745 );
and \g456170/U$8 ( \58370 , \57750 , \58369 );
xor \g456170/U$11 ( \58371 , \57735 , \57743 );
xor \g456170/U$11_r1 ( \58372 , \58371 , \57745 );
and \g456170/U$10 ( \58373 , \57758 , \58372 );
and \g456170/U$12 ( \58374 , \57750 , \57758 );
or \g456170/U$7 ( \58375 , \58370 , \58373 , \58374 );
xor \g132829/U$1 ( \58376 , \58367 , \58375 );
not \g133043/U$3 ( \58377 , \50759 );
and \g133073/U$2 ( \58378 , \56446 , \51055 );
and \g133073/U$3 ( \58379 , \51053 , \56167 );
nor \g133073/U$1 ( \58380 , \58378 , \58379 );
not \g133043/U$4 ( \58381 , \58380 );
or \g133043/U$2 ( \58382 , \58377 , \58381 );
or \g133043/U$5 ( \58383 , \58380 , \50759 );
nand \g133043/U$1 ( \58384 , \58382 , \58383 );
xor \g456170/U$5 ( \58385 , \57735 , \57743 );
and \g456170/U$4 ( \58386 , \58385 , \57745 );
and \g456170/U$6 ( \58387 , \57735 , \57743 );
or \g456170/U$3 ( \58388 , \58386 , \58387 );
xor \g132889/U$1 ( \58389 , \58384 , \58388 );
and \g133049/U$2 ( \58390 , \57819 , \57826 );
not \g133227/U$3 ( \58391 , \49568 );
and \g133267/U$2 ( \58392 , \49812 , \56349 );
and \g133267/U$3 ( \58393 , \56411 , \49813 );
nor \g133267/U$1 ( \58394 , \58392 , \58393 );
not \g133227/U$4 ( \58395 , \58394 );
or \g133227/U$2 ( \58396 , \58391 , \58395 );
or \g133227/U$5 ( \58397 , \58394 , \49568 );
nand \g133227/U$1 ( \58398 , \58396 , \58397 );
xor \g132970/U$1 ( \58399 , \58390 , \58398 );
not \g133137/U$3 ( \58400 , \49233 );
and \g133159/U$2 ( \58401 , \49403 , \56368 );
and \g133159/U$3 ( \58402 , \56370 , \49405 );
nor \g133159/U$1 ( \58403 , \58401 , \58402 );
not \g133137/U$4 ( \58404 , \58403 );
or \g133137/U$2 ( \58405 , \58400 , \58404 );
or \g133137/U$5 ( \58406 , \58403 , \49233 );
nand \g133137/U$1 ( \58407 , \58405 , \58406 );
not \g133064/U$3 ( \58408 , \49014 );
and \g133102/U$2 ( \58409 , \49075 , \56377 );
and \g133102/U$3 ( \58410 , \56379 , \49074 );
nor \g133102/U$1 ( \58411 , \58409 , \58410 );
not \g133064/U$4 ( \58412 , \58411 );
or \g133064/U$2 ( \58413 , \58408 , \58412 );
or \g133064/U$5 ( \58414 , \58411 , \49014 );
nand \g133064/U$1 ( \58415 , \58413 , \58414 );
xor \g133036/U$1 ( \58416 , \58407 , \58415 );
xor \g132970/U$1_r1 ( \58417 , \58399 , \58416 );
xor \g132889/U$1_r1 ( \58418 , \58389 , \58417 );
xor \g132829/U$1_r1 ( \58419 , \58376 , \58418 );
xor \g456167/U$1_r1 ( \58420 , \58363 , \58419 );
xor \g456167/U$1_r2 ( \58421 , \58359 , \58420 );
and \g132518/U$3 ( \58422 , \58320 , \58421 );
and \g132518/U$5 ( \58423 , \58315 , \58319 );
or \g132518/U$2 ( \58424 , \58422 , \58423 );
xor \g456167/U$9 ( \58425 , \58342 , \58350 );
xor \g456167/U$9_r1 ( \58426 , \58425 , \58358 );
and \g456167/U$8 ( \58427 , \58363 , \58426 );
xor \g456167/U$11 ( \58428 , \58342 , \58350 );
xor \g456167/U$11_r1 ( \58429 , \58428 , \58358 );
and \g456167/U$10 ( \58430 , \58419 , \58429 );
and \g456167/U$12 ( \58431 , \58363 , \58419 );
or \g456167/U$7 ( \58432 , \58427 , \58430 , \58431 );
xor \g132291/U$4 ( \58433 , \58424 , \58432 );
xor \g456172/U$2 ( \58434 , \57996 , \58011 );
xor \g456172/U$1 ( \58435 , \58434 , \58019 );
xor \g456172/U$1_r1 ( \58436 , \57962 , \58180 );
xor \g456172/U$1_r2 ( \58437 , \58435 , \58436 );
nor \g133834/U$1 ( \58438 , \58068 , \58072 );
xor \g133537/U$1 ( \58439 , \58071 , \58082 );
xor \g133537/U$1_r1 ( \58440 , \58439 , \58090 );
and \g133477/U$2 ( \58441 , \58438 , \58440 );
xor \g133351/U$4 ( \58442 , \58441 , \58031 );
xor \g133396/U$1 ( \58443 , \58093 , \58103 );
xor \g133396/U$1_r1 ( \58444 , \58443 , \58111 );
and \g133351/U$3 ( \58445 , \58442 , \58444 );
and \g133351/U$5 ( \58446 , \58441 , \58031 );
or \g133351/U$2 ( \58447 , \58445 , \58446 );
xor \g133291/U$1 ( \58448 , \58114 , \58115 );
xor \g133291/U$1_r1 ( \58449 , \58448 , \58134 );
and \g133249/U$2 ( \58450 , \58447 , \58449 );
xor \g133478/U$1 ( \58451 , \50362 , \57901 );
xor \g133150/U$4 ( \58452 , \58450 , \58451 );
xor \g133213/U$1 ( \58453 , \58137 , \58141 );
xor \g133213/U$1_r1 ( \58454 , \58453 , \58160 );
and \g133150/U$3 ( \58455 , \58452 , \58454 );
and \g133150/U$5 ( \58456 , \58450 , \58451 );
or \g133150/U$2 ( \58457 , \58455 , \58456 );
xor \g133128/U$1 ( \58458 , \58163 , \58167 );
xor \g133128/U$1_r1 ( \58459 , \58458 , \58172 );
and \g133108/U$2 ( \58460 , \58457 , \58459 );
xor \g133348/U$1 ( \58461 , \49925 , \57985 );
xor \g133030/U$4 ( \58462 , \58460 , \58461 );
xor \g456173/U$2 ( \58463 , \57930 , \57951 );
xor \g456173/U$1 ( \58464 , \58463 , \57959 );
xor \g456173/U$1_r1 ( \58465 , \58057 , \58175 );
xor \g456173/U$1_r2 ( \58466 , \58464 , \58465 );
and \g133030/U$3 ( \58467 , \58462 , \58466 );
and \g133030/U$5 ( \58468 , \58460 , \58461 );
or \g133030/U$2 ( \58469 , \58467 , \58468 );
and \g132977/U$2 ( \58470 , \58437 , \58469 );
xor \g133247/U$1 ( \58471 , \49568 , \57565 );
xor \g132891/U$4 ( \58472 , \58470 , \58471 );
xor \g132976/U$1 ( \58473 , \58185 , \58189 );
xor \g132976/U$1_r1 ( \58474 , \58473 , \58229 );
and \g132891/U$3 ( \58475 , \58472 , \58474 );
and \g132891/U$5 ( \58476 , \58470 , \58471 );
or \g132891/U$2 ( \58477 , \58475 , \58476 );
xor \g132920/U$1 ( \58478 , \58232 , \58240 );
xor \g132920/U$1_r1 ( \58479 , \58478 , \58270 );
and \g132866/U$2 ( \58480 , \58477 , \58479 );
xor \g132770/U$4 ( \58481 , \58480 , \57528 );
xor \g132864/U$1 ( \58482 , \58273 , \58281 );
xor \g132864/U$1_r1 ( \58483 , \58482 , \58292 );
and \g132770/U$3 ( \58484 , \58481 , \58483 );
and \g132770/U$5 ( \58485 , \58480 , \57528 );
or \g132770/U$2 ( \58486 , \58484 , \58485 );
xor \g132790/U$1 ( \58487 , \58295 , \58299 );
xor \g132790/U$1_r1 ( \58488 , \58487 , \58302 );
and \g132698/U$2 ( \58489 , \58486 , \58488 );
xor \g133083/U$1 ( \58490 , \49014 , \57825 );
xor \g132586/U$4 ( \58491 , \58489 , \58490 );
xor \g456168/U$2 ( \58492 , \57624 , \57678 );
xor \g456168/U$1 ( \58493 , \58492 , \57724 );
xor \g456168/U$1_r1 ( \58494 , \57884 , \58305 );
xor \g456168/U$1_r2 ( \58495 , \58493 , \58494 );
and \g132586/U$3 ( \58496 , \58491 , \58495 );
and \g132586/U$5 ( \58497 , \58489 , \58490 );
or \g132586/U$2 ( \58498 , \58496 , \58497 );
xor \g456165/U$2 ( \58499 , \57760 , \57764 );
xor \g456165/U$1 ( \58500 , \58499 , \57830 );
xor \g456165/U$1_r1 ( \58501 , \57727 , \58310 );
xor \g456165/U$1_r2 ( \58502 , \58500 , \58501 );
and \g132556/U$2 ( \58503 , \58498 , \58502 );
nor \g133056/U$1 ( \58504 , \48859 , \47025 );
xor \g132437/U$4 ( \58505 , \58503 , \58504 );
xor \g132518/U$1 ( \58506 , \58315 , \58319 );
xor \g132518/U$1_r1 ( \58507 , \58506 , \58421 );
and \g132437/U$3 ( \58508 , \58505 , \58507 );
and \g132437/U$5 ( \58509 , \58503 , \58504 );
or \g132437/U$2 ( \58510 , \58508 , \58509 );
and \g132291/U$3 ( \58511 , \58433 , \58510 );
and \g132291/U$5 ( \58512 , \58424 , \58432 );
or \g132291/U$2 ( \58513 , \58511 , \58512 );
nand \g132978/U$1 ( \58514 , \47026 , \48478 );
not \g132960/U$3 ( \58515 , \58514 );
not \g132960/U$4 ( \58516 , \48483 );
or \g132960/U$2 ( \58517 , \58515 , \58516 );
or \g132960/U$5 ( \58518 , \48483 , \58514 );
nand \g132960/U$1 ( \58519 , \58517 , \58518 );
xor \g132924/U$1 ( \58520 , \48483 , \58519 );
xor \g132109/U$4 ( \58521 , \58513 , \58520 );
not \g133091/U$3 ( \58522 , \50362 );
and \g133119/U$2 ( \58523 , \56446 , \50587 );
and \g133119/U$3 ( \58524 , \50588 , \56448 );
nor \g133119/U$1 ( \58525 , \58523 , \58524 );
not \g133091/U$4 ( \58526 , \58525 );
or \g133091/U$2 ( \58527 , \58522 , \58526 );
or \g133091/U$5 ( \58528 , \58525 , \50362 );
nand \g133091/U$1 ( \58529 , \58527 , \58528 );
not \g133195/U$3 ( \58530 , \49925 );
and \g133232/U$2 ( \58531 , \56357 , \50159 );
and \g133232/U$3 ( \58532 , \50160 , \56359 );
nor \g133232/U$1 ( \58533 , \58531 , \58532 );
not \g133195/U$4 ( \58534 , \58533 );
or \g133195/U$2 ( \58535 , \58530 , \58534 );
or \g133195/U$5 ( \58536 , \58533 , \49925 );
nand \g133195/U$1 ( \58537 , \58535 , \58536 );
xor \g132888/U$1 ( \58538 , \58529 , \58537 );
xor \g132970/U$4 ( \58539 , \58390 , \58398 );
and \g132970/U$3 ( \58540 , \58539 , \58416 );
and \g132970/U$5 ( \58541 , \58390 , \58398 );
or \g132970/U$2 ( \58542 , \58540 , \58541 );
xor \g132888/U$1_r1 ( \58543 , \58538 , \58542 );
not \g132881/U$3 ( \58544 , \51124 );
and \g132916/U$2 ( \58545 , \55460 , \51517 );
and \g132916/U$3 ( \58546 , \51518 , \55707 );
nor \g132916/U$1 ( \58547 , \58545 , \58546 );
not \g132881/U$4 ( \58548 , \58547 );
or \g132881/U$2 ( \58549 , \58544 , \58548 );
or \g132881/U$5 ( \58550 , \58547 , \51124 );
nand \g132881/U$1 ( \58551 , \58549 , \58550 );
xor \g456164/U$2 ( \58552 , \58543 , \58551 );
and \g132789/U$2 ( \58553 , \54853 , \52270 );
and \g132789/U$3 ( \58554 , \52273 , \55127 );
nor \g132789/U$1 ( \58555 , \58553 , \58554 );
and \g132747/U$2 ( \58556 , \58555 , \51513 );
not \g132747/U$4 ( \58557 , \58555 );
and \g132747/U$3 ( \58558 , \58557 , \51120 );
nor \g132747/U$1 ( \58559 , \58556 , \58558 );
xor \g456164/U$1 ( \58560 , \58552 , \58559 );
xor \g132829/U$4 ( \58561 , \58367 , \58375 );
and \g132829/U$3 ( \58562 , \58561 , \58418 );
and \g132829/U$5 ( \58563 , \58367 , \58375 );
or \g132829/U$2 ( \58564 , \58562 , \58563 );
xor \g456167/U$5 ( \58565 , \58342 , \58350 );
and \g456167/U$4 ( \58566 , \58565 , \58358 );
and \g456167/U$6 ( \58567 , \58342 , \58350 );
or \g456167/U$3 ( \58568 , \58566 , \58567 );
xor \g132889/U$4 ( \58569 , \58384 , \58388 );
and \g132889/U$3 ( \58570 , \58569 , \58417 );
and \g132889/U$5 ( \58571 , \58384 , \58388 );
or \g132889/U$2 ( \58572 , \58570 , \58571 );
xor \g132671/U$1 ( \58573 , \58568 , \58572 );
xor \g132918/U$4 ( \58574 , \58328 , \58336 );
and \g132918/U$3 ( \58575 , \58574 , \58341 );
and \g132918/U$5 ( \58576 , \58328 , \58336 );
or \g132918/U$2 ( \58577 , \58575 , \58576 );
not \g132991/U$3 ( \58578 , \50759 );
and \g133022/U$2 ( \58579 , \56167 , \51055 );
and \g133022/U$3 ( \58580 , \51053 , \55884 );
nor \g133022/U$1 ( \58581 , \58579 , \58580 );
not \g132991/U$4 ( \58582 , \58581 );
or \g132991/U$2 ( \58583 , \58578 , \58582 );
or \g132991/U$5 ( \58584 , \58581 , \50759 );
nand \g132991/U$1 ( \58585 , \58583 , \58584 );
xor \g132774/U$1 ( \58586 , \58577 , \58585 );
and \g133036/U$2 ( \58587 , \58407 , \58415 );
not \g133226/U$3 ( \58588 , \49568 );
and \g133263/U$2 ( \58589 , \56347 , \49812 );
and \g133263/U$3 ( \58590 , \56349 , \49813 );
nor \g133263/U$1 ( \58591 , \58589 , \58590 );
not \g133226/U$4 ( \58592 , \58591 );
or \g133226/U$2 ( \58593 , \58588 , \58592 );
or \g133226/U$5 ( \58594 , \58591 , \49568 );
nand \g133226/U$1 ( \58595 , \58593 , \58594 );
xor \g132863/U$1 ( \58596 , \58587 , \58595 );
not \g133059/U$3 ( \58597 , \49014 );
and \g133097/U$2 ( \58598 , \49074 , \56370 );
and \g133097/U$3 ( \58599 , \56379 , \49075 );
nor \g133097/U$1 ( \58600 , \58598 , \58599 );
not \g133059/U$4 ( \58601 , \58600 );
or \g133059/U$2 ( \58602 , \58597 , \58601 );
or \g133059/U$5 ( \58603 , \58600 , \49014 );
nand \g133059/U$1 ( \58604 , \58602 , \58603 );
not \g135546/U$2 ( \58605 , \48685 );
nor \g135546/U$1 ( \58606 , \58605 , \58504 );
xor \g133029/U$1 ( \58607 , \58604 , \58606 );
not \g133138/U$3 ( \58608 , \49233 );
and \g133157/U$2 ( \58609 , \49403 , \56411 );
and \g133157/U$3 ( \58610 , \56368 , \49405 );
nor \g133157/U$1 ( \58611 , \58609 , \58610 );
not \g133138/U$4 ( \58612 , \58611 );
or \g133138/U$2 ( \58613 , \58608 , \58612 );
or \g133138/U$5 ( \58614 , \58611 , \49233 );
nand \g133138/U$1 ( \58615 , \58613 , \58614 );
xor \g132925/U$1 ( \58616 , \58607 , \58615 );
not \g132992/U$3 ( \58617 , \48685 );
and \g133008/U$2 ( \58618 , \48860 , \47026 );
and \g133008/U$3 ( \58619 , \56377 , \48858 );
nor \g133008/U$1 ( \58620 , \58618 , \58619 );
not \g132992/U$4 ( \58621 , \58620 );
or \g132992/U$2 ( \58622 , \58617 , \58621 );
or \g132992/U$5 ( \58623 , \58620 , \48685 );
nand \g132992/U$1 ( \58624 , \58622 , \58623 );
xor \g132925/U$1_r1 ( \58625 , \58616 , \58624 );
xor \g132863/U$1_r1 ( \58626 , \58596 , \58625 );
xor \g132774/U$1_r1 ( \58627 , \58586 , \58626 );
xor \g132671/U$1_r1 ( \58628 , \58573 , \58627 );
xor \g456164/U$1_r1 ( \58629 , \58564 , \58628 );
xor \g456164/U$1_r2 ( \58630 , \58560 , \58629 );
xor \g132291/U$1 ( \58631 , \58424 , \58432 );
xor \g132291/U$1_r1 ( \58632 , \58631 , \58510 );
and \g132210/U$2 ( \58633 , \58630 , \58632 );
and \g132109/U$3 ( \58634 , \58521 , \58633 );
and \g132109/U$5 ( \58635 , \58513 , \58520 );
or \g132109/U$2 ( \58636 , \58634 , \58635 );
xor \g132774/U$4 ( \58637 , \58577 , \58585 );
and \g132774/U$3 ( \58638 , \58637 , \58626 );
and \g132774/U$5 ( \58639 , \58577 , \58585 );
or \g132774/U$2 ( \58640 , \58638 , \58639 );
xor \g132888/U$4 ( \58641 , \58529 , \58537 );
and \g132888/U$3 ( \58642 , \58641 , \58542 );
and \g132888/U$5 ( \58643 , \58529 , \58537 );
or \g132888/U$2 ( \58644 , \58642 , \58643 );
xor \g132626/U$1 ( \58645 , \58640 , \58644 );
and \g132730/U$2 ( \58646 , \54853 , \52273 );
and \g132730/U$3 ( \58647 , \52270 , \54537 );
nor \g132730/U$1 ( \58648 , \58646 , \58647 );
and \g132685/U$2 ( \58649 , \58648 , \51513 );
not \g132685/U$4 ( \58650 , \58648 );
and \g132685/U$3 ( \58651 , \58650 , \51120 );
nor \g132685/U$1 ( \58652 , \58649 , \58651 );
xor \g132626/U$1_r1 ( \58653 , \58645 , \58652 );
xor \g132671/U$4 ( \58654 , \58568 , \58572 );
and \g132671/U$3 ( \58655 , \58654 , \58627 );
and \g132671/U$5 ( \58656 , \58568 , \58572 );
or \g132671/U$2 ( \58657 , \58655 , \58656 );
xor \g456153/U$5 ( \58658 , \58653 , \58657 );
not \g132933/U$3 ( \58659 , \50759 );
and \g132967/U$2 ( \58660 , \55884 , \51055 );
and \g132967/U$3 ( \58661 , \51053 , \55707 );
nor \g132967/U$1 ( \58662 , \58660 , \58661 );
not \g132933/U$4 ( \58663 , \58662 );
or \g132933/U$2 ( \58664 , \58659 , \58663 );
or \g132933/U$5 ( \58665 , \58662 , \50759 );
nand \g132933/U$1 ( \58666 , \58664 , \58665 );
not \g133045/U$3 ( \58667 , \50362 );
and \g133074/U$2 ( \58668 , \56446 , \50588 );
and \g133074/U$3 ( \58669 , \50587 , \56167 );
nor \g133074/U$1 ( \58670 , \58668 , \58669 );
not \g133045/U$4 ( \58671 , \58670 );
or \g133045/U$2 ( \58672 , \58667 , \58671 );
or \g133045/U$5 ( \58673 , \58670 , \50362 );
nand \g133045/U$1 ( \58674 , \58672 , \58673 );
xor \g456166/U$2 ( \58675 , \58666 , \58674 );
and \g133029/U$2 ( \58676 , \58604 , \58606 );
not \g133140/U$3 ( \58677 , \49233 );
and \g133167/U$2 ( \58678 , \49403 , \56349 );
and \g133167/U$3 ( \58679 , \56411 , \49405 );
nor \g133167/U$1 ( \58680 , \58678 , \58679 );
not \g133140/U$4 ( \58681 , \58680 );
or \g133140/U$2 ( \58682 , \58677 , \58681 );
or \g133140/U$5 ( \58683 , \58680 , \49233 );
nand \g133140/U$1 ( \58684 , \58682 , \58683 );
xor \g132884/U$1 ( \58685 , \58676 , \58684 );
not \g133065/U$3 ( \58686 , \49014 );
and \g133105/U$2 ( \58687 , \49074 , \56368 );
and \g133105/U$3 ( \58688 , \56370 , \49075 );
nor \g133105/U$1 ( \58689 , \58687 , \58688 );
not \g133065/U$4 ( \58690 , \58689 );
or \g133065/U$2 ( \58691 , \58686 , \58690 );
or \g133065/U$5 ( \58692 , \58689 , \49014 );
nand \g133065/U$1 ( \58693 , \58691 , \58692 );
not \g132993/U$3 ( \58694 , \48685 );
and \g133009/U$2 ( \58695 , \48860 , \56377 );
and \g133009/U$3 ( \58696 , \56379 , \48858 );
nor \g133009/U$1 ( \58697 , \58695 , \58696 );
not \g132993/U$4 ( \58698 , \58697 );
or \g132993/U$2 ( \58699 , \58694 , \58698 );
or \g132993/U$5 ( \58700 , \58697 , \48685 );
nand \g132993/U$1 ( \58701 , \58699 , \58700 );
xor \g132958/U$1 ( \58702 , \58693 , \58701 );
xor \g132884/U$1_r1 ( \58703 , \58685 , \58702 );
xor \g456166/U$1 ( \58704 , \58675 , \58703 );
xor \g456164/U$5 ( \58705 , \58543 , \58551 );
and \g456164/U$4 ( \58706 , \58705 , \58559 );
and \g456164/U$6 ( \58707 , \58543 , \58551 );
or \g456164/U$3 ( \58708 , \58706 , \58707 );
xor \g132863/U$4 ( \58709 , \58587 , \58595 );
and \g132863/U$3 ( \58710 , \58709 , \58625 );
and \g132863/U$5 ( \58711 , \58587 , \58595 );
or \g132863/U$2 ( \58712 , \58710 , \58711 );
not \g132824/U$3 ( \58713 , \51124 );
and \g132861/U$2 ( \58714 , \55127 , \51517 );
and \g132861/U$3 ( \58715 , \51518 , \55460 );
nor \g132861/U$1 ( \58716 , \58714 , \58715 );
not \g132824/U$4 ( \58717 , \58716 );
or \g132824/U$2 ( \58718 , \58713 , \58717 );
or \g132824/U$5 ( \58719 , \58716 , \51124 );
nand \g132824/U$1 ( \58720 , \58718 , \58719 );
xor \g132769/U$1 ( \58721 , \58712 , \58720 );
not \g133139/U$3 ( \58722 , \49925 );
and \g133166/U$2 ( \58723 , \56357 , \50160 );
and \g133166/U$3 ( \58724 , \50159 , \56448 );
nor \g133166/U$1 ( \58725 , \58723 , \58724 );
not \g133139/U$4 ( \58726 , \58725 );
or \g133139/U$2 ( \58727 , \58722 , \58726 );
or \g133139/U$5 ( \58728 , \58725 , \49925 );
nand \g133139/U$1 ( \58729 , \58727 , \58728 );
not \g133225/U$3 ( \58730 , \49568 );
and \g133264/U$2 ( \58731 , \49813 , \56347 );
and \g133264/U$3 ( \58732 , \49812 , \56359 );
nor \g133264/U$1 ( \58733 , \58731 , \58732 );
not \g133225/U$4 ( \58734 , \58733 );
or \g133225/U$2 ( \58735 , \58730 , \58734 );
or \g133225/U$5 ( \58736 , \58733 , \49568 );
nand \g133225/U$1 ( \58737 , \58735 , \58736 );
xor \g132865/U$1 ( \58738 , \58729 , \58737 );
xor \g132925/U$4 ( \58739 , \58607 , \58615 );
and \g132925/U$3 ( \58740 , \58739 , \58624 );
and \g132925/U$5 ( \58741 , \58607 , \58615 );
or \g132925/U$2 ( \58742 , \58740 , \58741 );
xor \g132865/U$1_r1 ( \58743 , \58738 , \58742 );
xor \g132769/U$1_r1 ( \58744 , \58721 , \58743 );
xor \g456166/U$1_r1 ( \58745 , \58708 , \58744 );
xor \g456166/U$1_r2 ( \58746 , \58704 , \58745 );
and \g456153/U$4 ( \58747 , \58658 , \58746 );
and \g456153/U$6 ( \58748 , \58653 , \58657 );
or \g456153/U$3 ( \58749 , \58747 , \58748 );
xor \g131912/U$4 ( \58750 , \58636 , \58749 );
xor \g456164/U$9 ( \58751 , \58543 , \58551 );
xor \g456164/U$9_r1 ( \58752 , \58751 , \58559 );
and \g456164/U$8 ( \58753 , \58564 , \58752 );
xor \g456164/U$11 ( \58754 , \58543 , \58551 );
xor \g456164/U$11_r1 ( \58755 , \58754 , \58559 );
and \g456164/U$10 ( \58756 , \58628 , \58755 );
and \g456164/U$12 ( \58757 , \58564 , \58628 );
or \g456164/U$7 ( \58758 , \58753 , \58756 , \58757 );
xor \g456153/U$9 ( \58759 , \58653 , \58657 );
xor \g456153/U$9_r1 ( \58760 , \58759 , \58746 );
and \g456153/U$8 ( \58761 , \58758 , \58760 );
xor \g132109/U$1 ( \58762 , \58513 , \58520 );
xor \g132109/U$1_r1 ( \58763 , \58762 , \58633 );
xor \g456153/U$11 ( \58764 , \58653 , \58657 );
xor \g456153/U$11_r1 ( \58765 , \58764 , \58746 );
and \g456153/U$10 ( \58766 , \58763 , \58765 );
and \g456153/U$12 ( \58767 , \58758 , \58763 );
or \g456153/U$7 ( \58768 , \58761 , \58766 , \58767 );
and \g131912/U$3 ( \58769 , \58750 , \58768 );
and \g131912/U$5 ( \58770 , \58636 , \58749 );
or \g131912/U$2 ( \58771 , \58769 , \58770 );
nand \g132892/U$1 ( \58772 , \47026 , \48334 );
not \g132877/U$3 ( \58773 , \58772 );
not \g132877/U$4 ( \58774 , \48323 );
or \g132877/U$2 ( \58775 , \58773 , \58774 );
or \g132877/U$5 ( \58776 , \48323 , \58772 );
nand \g132877/U$1 ( \58777 , \58775 , \58776 );
xor \g132832/U$1 ( \58778 , \48323 , \58777 );
xor \g131776/U$4 ( \58779 , \58771 , \58778 );
xor \g132769/U$4 ( \58780 , \58712 , \58720 );
and \g132769/U$3 ( \58781 , \58780 , \58743 );
and \g132769/U$5 ( \58782 , \58712 , \58720 );
or \g132769/U$2 ( \58783 , \58781 , \58782 );
xor \g456166/U$5 ( \58784 , \58666 , \58674 );
and \g456166/U$4 ( \58785 , \58784 , \58703 );
and \g456166/U$6 ( \58786 , \58666 , \58674 );
or \g456166/U$3 ( \58787 , \58785 , \58786 );
xor \g456162/U$2 ( \58788 , \58783 , \58787 );
and \g132668/U$2 ( \58789 , \54537 , \52273 );
and \g132668/U$3 ( \58790 , \52270 , \54529 );
nor \g132668/U$1 ( \58791 , \58789 , \58790 );
and \g132619/U$2 ( \58792 , \58791 , \51513 );
not \g132619/U$4 ( \58793 , \58791 );
and \g132619/U$3 ( \58794 , \58793 , \51120 );
nor \g132619/U$1 ( \58795 , \58792 , \58794 );
xor \g456162/U$1 ( \58796 , \58788 , \58795 );
xor \g456166/U$9 ( \58797 , \58666 , \58674 );
xor \g456166/U$9_r1 ( \58798 , \58797 , \58703 );
and \g456166/U$8 ( \58799 , \58708 , \58798 );
xor \g456166/U$11 ( \58800 , \58666 , \58674 );
xor \g456166/U$11_r1 ( \58801 , \58800 , \58703 );
and \g456166/U$10 ( \58802 , \58744 , \58801 );
and \g456166/U$12 ( \58803 , \58708 , \58744 );
or \g456166/U$7 ( \58804 , \58799 , \58802 , \58803 );
not \g132740/U$3 ( \58805 , \51124 );
and \g132788/U$2 ( \58806 , \54853 , \51517 );
and \g132788/U$3 ( \58807 , \51518 , \55127 );
nor \g132788/U$1 ( \58808 , \58806 , \58807 );
not \g132740/U$4 ( \58809 , \58808 );
or \g132740/U$2 ( \58810 , \58805 , \58809 );
or \g132740/U$5 ( \58811 , \58808 , \51124 );
nand \g132740/U$1 ( \58812 , \58810 , \58811 );
not \g132880/U$3 ( \58813 , \50759 );
and \g132913/U$2 ( \58814 , \55460 , \51053 );
and \g132913/U$3 ( \58815 , \51055 , \55707 );
nor \g132913/U$1 ( \58816 , \58814 , \58815 );
not \g132880/U$4 ( \58817 , \58816 );
or \g132880/U$2 ( \58818 , \58813 , \58817 );
or \g132880/U$5 ( \58819 , \58816 , \50759 );
nand \g132880/U$1 ( \58820 , \58818 , \58819 );
xor \g456163/U$2 ( \58821 , \58812 , \58820 );
not \g133094/U$3 ( \58822 , \49925 );
and \g133116/U$2 ( \58823 , \56446 , \50159 );
and \g133116/U$3 ( \58824 , \50160 , \56448 );
nor \g133116/U$1 ( \58825 , \58823 , \58824 );
not \g133094/U$4 ( \58826 , \58825 );
or \g133094/U$2 ( \58827 , \58822 , \58826 );
or \g133094/U$5 ( \58828 , \58825 , \49925 );
nand \g133094/U$1 ( \58829 , \58827 , \58828 );
not \g133194/U$3 ( \58830 , \49568 );
and \g133233/U$2 ( \58831 , \56357 , \49812 );
and \g133233/U$3 ( \58832 , \56359 , \49813 );
nor \g133233/U$1 ( \58833 , \58831 , \58832 );
not \g133194/U$4 ( \58834 , \58833 );
or \g133194/U$2 ( \58835 , \58830 , \58834 );
or \g133194/U$5 ( \58836 , \58833 , \49568 );
nand \g133194/U$1 ( \58837 , \58835 , \58836 );
xor \g132795/U$1 ( \58838 , \58829 , \58837 );
xor \g132884/U$4 ( \58839 , \58676 , \58684 );
and \g132884/U$3 ( \58840 , \58839 , \58702 );
and \g132884/U$5 ( \58841 , \58676 , \58684 );
or \g132884/U$2 ( \58842 , \58840 , \58841 );
xor \g132795/U$1_r1 ( \58843 , \58838 , \58842 );
xor \g456163/U$1 ( \58844 , \58821 , \58843 );
xor \g132626/U$4 ( \58845 , \58640 , \58644 );
and \g132626/U$3 ( \58846 , \58845 , \58652 );
and \g132626/U$5 ( \58847 , \58640 , \58644 );
or \g132626/U$2 ( \58848 , \58846 , \58847 );
xor \g132865/U$4 ( \58849 , \58729 , \58737 );
and \g132865/U$3 ( \58850 , \58849 , \58742 );
and \g132865/U$5 ( \58851 , \58729 , \58737 );
or \g132865/U$2 ( \58852 , \58850 , \58851 );
not \g132998/U$3 ( \58853 , \50362 );
and \g133026/U$2 ( \58854 , \56167 , \50588 );
and \g133026/U$3 ( \58855 , \50587 , \55884 );
nor \g133026/U$1 ( \58856 , \58854 , \58855 );
not \g132998/U$4 ( \58857 , \58856 );
or \g132998/U$2 ( \58858 , \58853 , \58857 );
or \g132998/U$5 ( \58859 , \58856 , \50362 );
nand \g132998/U$1 ( \58860 , \58858 , \58859 );
xor \g132634/U$1 ( \58861 , \58852 , \58860 );
and \g132958/U$2 ( \58862 , \58693 , \58701 );
not \g133146/U$3 ( \58863 , \49233 );
and \g133168/U$2 ( \58864 , \49403 , \56347 );
and \g133168/U$3 ( \58865 , \56349 , \49405 );
nor \g133168/U$1 ( \58866 , \58864 , \58865 );
not \g133146/U$4 ( \58867 , \58866 );
or \g133146/U$2 ( \58868 , \58863 , \58867 );
or \g133146/U$5 ( \58869 , \58866 , \49233 );
nand \g133146/U$1 ( \58870 , \58868 , \58869 );
xor \g132732/U$1 ( \58871 , \58862 , \58870 );
not \g132901/U$3 ( \58872 , \48483 );
and \g132938/U$2 ( \58873 , \48479 , \47026 );
and \g132938/U$3 ( \58874 , \56377 , \48478 );
nor \g132938/U$1 ( \58875 , \58873 , \58874 );
not \g132901/U$4 ( \58876 , \58875 );
or \g132901/U$2 ( \58877 , \58872 , \58876 );
or \g132901/U$5 ( \58878 , \58875 , \48483 );
nand \g132901/U$1 ( \58879 , \58877 , \58878 );
not \g133067/U$3 ( \58880 , \49014 );
and \g133101/U$2 ( \58881 , \49074 , \56411 );
and \g133101/U$3 ( \58882 , \56368 , \49075 );
nor \g133101/U$1 ( \58883 , \58881 , \58882 );
not \g133067/U$4 ( \58884 , \58883 );
or \g133067/U$2 ( \58885 , \58880 , \58884 );
or \g133067/U$5 ( \58886 , \58883 , \49014 );
nand \g133067/U$1 ( \58887 , \58885 , \58886 );
xor \g132797/U$1 ( \58888 , \58879 , \58887 );
not \g132997/U$3 ( \58889 , \48685 );
and \g133020/U$2 ( \58890 , \48858 , \56370 );
and \g133020/U$3 ( \58891 , \56379 , \48860 );
nor \g133020/U$1 ( \58892 , \58890 , \58891 );
not \g132997/U$4 ( \58893 , \58892 );
or \g132997/U$2 ( \58894 , \58889 , \58893 );
or \g132997/U$5 ( \58895 , \58892 , \48685 );
nand \g132997/U$1 ( \58896 , \58894 , \58895 );
and \g132924/U$2 ( \58897 , \48483 , \58519 );
xor \g132883/U$1 ( \58898 , \58896 , \58897 );
xor \g132797/U$1_r1 ( \58899 , \58888 , \58898 );
xor \g132732/U$1_r1 ( \58900 , \58871 , \58899 );
xor \g132634/U$1_r1 ( \58901 , \58861 , \58900 );
xor \g456163/U$1_r1 ( \58902 , \58848 , \58901 );
xor \g456163/U$1_r2 ( \58903 , \58844 , \58902 );
xor \g456162/U$1_r1 ( \58904 , \58804 , \58903 );
xor \g456162/U$1_r2 ( \58905 , \58796 , \58904 );
xor \g131912/U$1 ( \58906 , \58636 , \58749 );
xor \g131912/U$1_r1 ( \58907 , \58906 , \58768 );
and \g131861/U$2 ( \58908 , \58905 , \58907 );
and \g131776/U$3 ( \58909 , \58779 , \58908 );
and \g131776/U$5 ( \58910 , \58771 , \58778 );
or \g131776/U$2 ( \58911 , \58909 , \58910 );
and \g132577/U$2 ( \58912 , \54251 , \52270 );
and \g132577/U$3 ( \58913 , \52273 , \54529 );
nor \g132577/U$1 ( \58914 , \58912 , \58913 );
and \g132534/U$2 ( \58915 , \58914 , \51513 );
not \g132534/U$4 ( \58916 , \58914 );
and \g132534/U$3 ( \58917 , \58916 , \51120 );
nor \g132534/U$1 ( \58918 , \58915 , \58917 );
not \g132935/U$3 ( \58919 , \50362 );
and \g132966/U$2 ( \58920 , \55884 , \50588 );
and \g132966/U$3 ( \58921 , \50587 , \55707 );
nor \g132966/U$1 ( \58922 , \58920 , \58921 );
not \g132935/U$4 ( \58923 , \58922 );
or \g132935/U$2 ( \58924 , \58919 , \58923 );
or \g132935/U$5 ( \58925 , \58922 , \50362 );
nand \g132935/U$1 ( \58926 , \58924 , \58925 );
not \g133039/U$3 ( \58927 , \49925 );
and \g133071/U$2 ( \58928 , \56446 , \50160 );
and \g133071/U$3 ( \58929 , \50159 , \56167 );
nor \g133071/U$1 ( \58930 , \58928 , \58929 );
not \g133039/U$4 ( \58931 , \58930 );
or \g133039/U$2 ( \58932 , \58927 , \58931 );
or \g133039/U$5 ( \58933 , \58930 , \49925 );
nand \g133039/U$1 ( \58934 , \58932 , \58933 );
xor \g132731/U$1 ( \58935 , \58926 , \58934 );
not \g133062/U$3 ( \58936 , \49014 );
and \g133104/U$2 ( \58937 , \49074 , \56349 );
and \g133104/U$3 ( \58938 , \56411 , \49075 );
nor \g133104/U$1 ( \58939 , \58937 , \58938 );
not \g133062/U$4 ( \58940 , \58939 );
or \g133062/U$2 ( \58941 , \58936 , \58940 );
or \g133062/U$5 ( \58942 , \58939 , \49014 );
nand \g133062/U$1 ( \58943 , \58941 , \58942 );
not \g133132/U$3 ( \58944 , \49233 );
and \g133161/U$2 ( \58945 , \49405 , \56347 );
and \g133161/U$3 ( \58946 , \56359 , \49403 );
nor \g133161/U$1 ( \58947 , \58945 , \58946 );
not \g133132/U$4 ( \58948 , \58947 );
or \g133132/U$2 ( \58949 , \58944 , \58948 );
or \g133132/U$5 ( \58950 , \58947 , \49233 );
nand \g133132/U$1 ( \58951 , \58949 , \58950 );
xor \g132796/U$1 ( \58952 , \58943 , \58951 );
and \g132883/U$2 ( \58953 , \58896 , \58897 );
xor \g132796/U$1_r1 ( \58954 , \58952 , \58953 );
xor \g132731/U$1_r1 ( \58955 , \58935 , \58954 );
xor \g132461/U$1 ( \58956 , \58918 , \58955 );
xor \g132732/U$4 ( \58957 , \58862 , \58870 );
and \g132732/U$3 ( \58958 , \58957 , \58899 );
and \g132732/U$5 ( \58959 , \58862 , \58870 );
or \g132732/U$2 ( \58960 , \58958 , \58959 );
xor \g132795/U$4 ( \58961 , \58829 , \58837 );
and \g132795/U$3 ( \58962 , \58961 , \58842 );
and \g132795/U$5 ( \58963 , \58829 , \58837 );
or \g132795/U$2 ( \58964 , \58962 , \58963 );
xor \g132627/U$1 ( \58965 , \58960 , \58964 );
not \g132996/U$3 ( \58966 , \48685 );
and \g133024/U$2 ( \58967 , \48858 , \56368 );
and \g133024/U$3 ( \58968 , \56370 , \48860 );
nor \g133024/U$1 ( \58969 , \58967 , \58968 );
not \g132996/U$4 ( \58970 , \58969 );
or \g132996/U$2 ( \58971 , \58966 , \58970 );
or \g132996/U$5 ( \58972 , \58969 , \48685 );
nand \g132996/U$1 ( \58973 , \58971 , \58972 );
not \g132894/U$3 ( \58974 , \48483 );
and \g132950/U$2 ( \58975 , \48479 , \56377 );
and \g132950/U$3 ( \58976 , \56379 , \48478 );
nor \g132950/U$1 ( \58977 , \58975 , \58976 );
not \g132894/U$4 ( \58978 , \58977 );
or \g132894/U$2 ( \58979 , \58974 , \58978 );
or \g132894/U$5 ( \58980 , \58977 , \48483 );
nand \g132894/U$1 ( \58981 , \58979 , \58980 );
xor \g132870/U$1 ( \58982 , \58973 , \58981 );
not \g133134/U$3 ( \58983 , \49568 );
and \g133169/U$2 ( \58984 , \56357 , \49813 );
and \g133169/U$3 ( \58985 , \49812 , \56448 );
nor \g133169/U$1 ( \58986 , \58984 , \58985 );
not \g133134/U$4 ( \58987 , \58986 );
or \g133134/U$2 ( \58988 , \58983 , \58987 );
or \g133134/U$5 ( \58989 , \58986 , \49568 );
nand \g133134/U$1 ( \58990 , \58988 , \58989 );
xor \g132733/U$1 ( \58991 , \58982 , \58990 );
xor \g132797/U$4 ( \58992 , \58879 , \58887 );
and \g132797/U$3 ( \58993 , \58992 , \58898 );
and \g132797/U$5 ( \58994 , \58879 , \58887 );
or \g132797/U$2 ( \58995 , \58993 , \58994 );
xor \g132733/U$1_r1 ( \58996 , \58991 , \58995 );
xor \g132627/U$1_r1 ( \58997 , \58965 , \58996 );
xor \g132461/U$1_r1 ( \58998 , \58956 , \58997 );
xor \g456163/U$9 ( \58999 , \58812 , \58820 );
xor \g456163/U$9_r1 ( \59000 , \58999 , \58843 );
and \g456163/U$8 ( \59001 , \58848 , \59000 );
xor \g456163/U$11 ( \59002 , \58812 , \58820 );
xor \g456163/U$11_r1 ( \59003 , \59002 , \58843 );
and \g456163/U$10 ( \59004 , \58901 , \59003 );
and \g456163/U$12 ( \59005 , \58848 , \58901 );
or \g456163/U$7 ( \59006 , \59001 , \59004 , \59005 );
xor \g456139/U$5 ( \59007 , \58998 , \59006 );
xor \g456162/U$5 ( \59008 , \58783 , \58787 );
and \g456162/U$4 ( \59009 , \59008 , \58795 );
and \g456162/U$6 ( \59010 , \58783 , \58787 );
or \g456162/U$3 ( \59011 , \59009 , \59010 );
xor \g456163/U$5 ( \59012 , \58812 , \58820 );
and \g456163/U$4 ( \59013 , \59012 , \58843 );
and \g456163/U$6 ( \59014 , \58812 , \58820 );
or \g456163/U$3 ( \59015 , \59013 , \59014 );
xor \g132442/U$1 ( \59016 , \59011 , \59015 );
not \g132686/U$3 ( \59017 , \51124 );
and \g132729/U$2 ( \59018 , \54853 , \51518 );
and \g132729/U$3 ( \59019 , \51517 , \54537 );
nor \g132729/U$1 ( \59020 , \59018 , \59019 );
not \g132686/U$4 ( \59021 , \59020 );
or \g132686/U$2 ( \59022 , \59017 , \59021 );
or \g132686/U$5 ( \59023 , \59020 , \51124 );
nand \g132686/U$1 ( \59024 , \59022 , \59023 );
not \g132825/U$3 ( \59025 , \50759 );
and \g132858/U$2 ( \59026 , \55127 , \51053 );
and \g132858/U$3 ( \59027 , \51055 , \55460 );
nor \g132858/U$1 ( \59028 , \59026 , \59027 );
not \g132825/U$4 ( \59029 , \59028 );
or \g132825/U$2 ( \59030 , \59025 , \59029 );
or \g132825/U$5 ( \59031 , \59028 , \50759 );
nand \g132825/U$1 ( \59032 , \59030 , \59031 );
xor \g132558/U$1 ( \59033 , \59024 , \59032 );
xor \g132634/U$4 ( \59034 , \58852 , \58860 );
and \g132634/U$3 ( \59035 , \59034 , \58900 );
and \g132634/U$5 ( \59036 , \58852 , \58860 );
or \g132634/U$2 ( \59037 , \59035 , \59036 );
xor \g132558/U$1_r1 ( \59038 , \59033 , \59037 );
xor \g132442/U$1_r1 ( \59039 , \59016 , \59038 );
and \g456139/U$4 ( \59040 , \59007 , \59039 );
and \g456139/U$6 ( \59041 , \58998 , \59006 );
or \g456139/U$3 ( \59042 , \59040 , \59041 );
xor \g131614/U$4 ( \59043 , \58911 , \59042 );
xor \g456162/U$9 ( \59044 , \58783 , \58787 );
xor \g456162/U$9_r1 ( \59045 , \59044 , \58795 );
and \g456162/U$8 ( \59046 , \58804 , \59045 );
xor \g456162/U$11 ( \59047 , \58783 , \58787 );
xor \g456162/U$11_r1 ( \59048 , \59047 , \58795 );
and \g456162/U$10 ( \59049 , \58903 , \59048 );
and \g456162/U$12 ( \59050 , \58804 , \58903 );
or \g456162/U$7 ( \59051 , \59046 , \59049 , \59050 );
xor \g456139/U$9 ( \59052 , \58998 , \59006 );
xor \g456139/U$9_r1 ( \59053 , \59052 , \59039 );
and \g456139/U$8 ( \59054 , \59051 , \59053 );
xor \g131776/U$1 ( \59055 , \58771 , \58778 );
xor \g131776/U$1_r1 ( \59056 , \59055 , \58908 );
xor \g456139/U$11 ( \59057 , \58998 , \59006 );
xor \g456139/U$11_r1 ( \59058 , \59057 , \59039 );
and \g456139/U$10 ( \59059 , \59056 , \59058 );
and \g456139/U$12 ( \59060 , \59051 , \59056 );
or \g456139/U$7 ( \59061 , \59054 , \59059 , \59060 );
and \g131614/U$3 ( \59062 , \59043 , \59061 );
and \g131614/U$5 ( \59063 , \58911 , \59042 );
or \g131614/U$2 ( \59064 , \59062 , \59063 );
nand \g132799/U$1 ( \59065 , \47026 , \48154 );
not \g132778/U$3 ( \59066 , \59065 );
not \g132778/U$4 ( \59067 , \48159 );
or \g132778/U$2 ( \59068 , \59066 , \59067 );
or \g132778/U$5 ( \59069 , \48159 , \59065 );
nand \g132778/U$1 ( \59070 , \59068 , \59069 );
xor \g132735/U$1 ( \59071 , \48159 , \59070 );
xor \g131494/U$4 ( \59072 , \59064 , \59071 );
xor \g132461/U$4 ( \59073 , \58918 , \58955 );
and \g132461/U$3 ( \59074 , \59073 , \58997 );
and \g132461/U$5 ( \59075 , \58918 , \58955 );
or \g132461/U$2 ( \59076 , \59074 , \59075 );
xor \g132558/U$4 ( \59077 , \59024 , \59032 );
and \g132558/U$3 ( \59078 , \59077 , \59037 );
and \g132558/U$5 ( \59079 , \59024 , \59032 );
or \g132558/U$2 ( \59080 , \59078 , \59079 );
xor \g456159/U$2 ( \59081 , \59076 , \59080 );
not \g132620/U$3 ( \59082 , \51124 );
and \g132667/U$2 ( \59083 , \54537 , \51518 );
and \g132667/U$3 ( \59084 , \51517 , \54529 );
nor \g132667/U$1 ( \59085 , \59083 , \59084 );
not \g132620/U$4 ( \59086 , \59085 );
or \g132620/U$2 ( \59087 , \59082 , \59086 );
or \g132620/U$5 ( \59088 , \59085 , \51124 );
nand \g132620/U$1 ( \59089 , \59087 , \59088 );
xor \g132731/U$4 ( \59090 , \58926 , \58934 );
and \g132731/U$3 ( \59091 , \59090 , \58954 );
and \g132731/U$5 ( \59092 , \58926 , \58934 );
or \g132731/U$2 ( \59093 , \59091 , \59092 );
xor \g132515/U$1 ( \59094 , \59089 , \59093 );
xor \g132627/U$4 ( \59095 , \58960 , \58964 );
and \g132627/U$3 ( \59096 , \59095 , \58996 );
and \g132627/U$5 ( \59097 , \58960 , \58964 );
or \g132627/U$2 ( \59098 , \59096 , \59097 );
xor \g132515/U$1_r1 ( \59099 , \59094 , \59098 );
xor \g456159/U$1 ( \59100 , \59081 , \59099 );
xor \g132442/U$4 ( \59101 , \59011 , \59015 );
and \g132442/U$3 ( \59102 , \59101 , \59038 );
and \g132442/U$5 ( \59103 , \59011 , \59015 );
or \g132442/U$2 ( \59104 , \59102 , \59103 );
and \g132504/U$2 ( \59105 , \54185 , \52270 );
and \g132504/U$3 ( \59106 , \52273 , \54251 );
nor \g132504/U$1 ( \59107 , \59105 , \59106 );
and \g132457/U$2 ( \59108 , \59107 , \51513 );
not \g132457/U$4 ( \59109 , \59107 );
and \g132457/U$3 ( \59110 , \59109 , \51120 );
nor \g132457/U$1 ( \59111 , \59108 , \59110 );
xor \g132733/U$4 ( \59112 , \58982 , \58990 );
and \g132733/U$3 ( \59113 , \59112 , \58995 );
and \g132733/U$5 ( \59114 , \58982 , \58990 );
or \g132733/U$2 ( \59115 , \59113 , \59114 );
not \g132990/U$3 ( \59116 , \49925 );
and \g133021/U$2 ( \59117 , \56167 , \50160 );
and \g133021/U$3 ( \59118 , \50159 , \55884 );
nor \g133021/U$1 ( \59119 , \59117 , \59118 );
not \g132990/U$4 ( \59120 , \59119 );
or \g132990/U$2 ( \59121 , \59116 , \59120 );
or \g132990/U$5 ( \59122 , \59119 , \49925 );
nand \g132990/U$1 ( \59123 , \59121 , \59122 );
xor \g132631/U$1 ( \59124 , \59115 , \59123 );
not \g133068/U$3 ( \59125 , \49014 );
and \g133103/U$2 ( \59126 , \49074 , \56347 );
and \g133103/U$3 ( \59127 , \56349 , \49075 );
nor \g133103/U$1 ( \59128 , \59126 , \59127 );
not \g133068/U$4 ( \59129 , \59128 );
or \g133068/U$2 ( \59130 , \59125 , \59129 );
or \g133068/U$5 ( \59131 , \59128 , \49014 );
nand \g133068/U$1 ( \59132 , \59130 , \59131 );
not \g133133/U$3 ( \59133 , \49233 );
and \g133162/U$2 ( \59134 , \56357 , \49403 );
and \g133162/U$3 ( \59135 , \56359 , \49405 );
nor \g133162/U$1 ( \59136 , \59134 , \59135 );
not \g133133/U$4 ( \59137 , \59136 );
or \g133133/U$2 ( \59138 , \59133 , \59137 );
or \g133133/U$5 ( \59139 , \59136 , \49233 );
nand \g133133/U$1 ( \59140 , \59138 , \59139 );
xor \g132791/U$1 ( \59141 , \59132 , \59140 );
and \g132870/U$2 ( \59142 , \58973 , \58981 );
xor \g132791/U$1_r1 ( \59143 , \59141 , \59142 );
xor \g132631/U$1_r1 ( \59144 , \59124 , \59143 );
xor \g132360/U$1 ( \59145 , \59111 , \59144 );
not \g132749/U$3 ( \59146 , \50759 );
and \g132786/U$2 ( \59147 , \54853 , \51053 );
and \g132786/U$3 ( \59148 , \51055 , \55127 );
nor \g132786/U$1 ( \59149 , \59147 , \59148 );
not \g132749/U$4 ( \59150 , \59149 );
or \g132749/U$2 ( \59151 , \59146 , \59150 );
or \g132749/U$5 ( \59152 , \59149 , \50759 );
nand \g132749/U$1 ( \59153 , \59151 , \59152 );
not \g132878/U$3 ( \59154 , \50362 );
and \g132912/U$2 ( \59155 , \55460 , \50587 );
and \g132912/U$3 ( \59156 , \50588 , \55707 );
nor \g132912/U$1 ( \59157 , \59155 , \59156 );
not \g132878/U$4 ( \59158 , \59157 );
or \g132878/U$2 ( \59159 , \59154 , \59158 );
or \g132878/U$5 ( \59160 , \59157 , \50362 );
nand \g132878/U$1 ( \59161 , \59159 , \59160 );
xor \g132509/U$1 ( \59162 , \59153 , \59161 );
xor \g132796/U$4 ( \59163 , \58943 , \58951 );
and \g132796/U$3 ( \59164 , \59163 , \58953 );
and \g132796/U$5 ( \59165 , \58943 , \58951 );
or \g132796/U$2 ( \59166 , \59164 , \59165 );
not \g133090/U$3 ( \59167 , \49568 );
and \g133120/U$2 ( \59168 , \56446 , \49812 );
and \g133120/U$3 ( \59169 , \49813 , \56448 );
nor \g133120/U$1 ( \59170 , \59168 , \59169 );
not \g133090/U$4 ( \59171 , \59170 );
or \g133090/U$2 ( \59172 , \59167 , \59171 );
or \g133090/U$5 ( \59173 , \59170 , \49568 );
nand \g133090/U$1 ( \59174 , \59172 , \59173 );
xor \g132587/U$1 ( \59175 , \59166 , \59174 );
not \g132903/U$3 ( \59176 , \48483 );
and \g132947/U$2 ( \59177 , \48478 , \56370 );
and \g132947/U$3 ( \59178 , \56379 , \48479 );
nor \g132947/U$1 ( \59179 , \59177 , \59178 );
not \g132903/U$4 ( \59180 , \59179 );
or \g132903/U$2 ( \59181 , \59176 , \59180 );
or \g132903/U$5 ( \59182 , \59179 , \48483 );
nand \g132903/U$1 ( \59183 , \59181 , \59182 );
not \g132988/U$3 ( \59184 , \48685 );
and \g133018/U$2 ( \59185 , \48858 , \56411 );
and \g133018/U$3 ( \59186 , \56368 , \48860 );
nor \g133018/U$1 ( \59187 , \59185 , \59186 );
not \g132988/U$4 ( \59188 , \59187 );
or \g132988/U$2 ( \59189 , \59184 , \59188 );
or \g132988/U$5 ( \59190 , \59187 , \48685 );
nand \g132988/U$1 ( \59191 , \59189 , \59190 );
xor \g132690/U$1 ( \59192 , \59183 , \59191 );
and \g132832/U$2 ( \59193 , \48323 , \58777 );
not \g132820/U$3 ( \59194 , \48323 );
and \g132837/U$2 ( \59195 , \48335 , \47026 );
and \g132837/U$3 ( \59196 , \56377 , \48334 );
nor \g132837/U$1 ( \59197 , \59195 , \59196 );
not \g132820/U$4 ( \59198 , \59197 );
or \g132820/U$2 ( \59199 , \59194 , \59198 );
or \g132820/U$5 ( \59200 , \59197 , \48323 );
nand \g132820/U$1 ( \59201 , \59199 , \59200 );
xor \g132773/U$1 ( \59202 , \59193 , \59201 );
xor \g132690/U$1_r1 ( \59203 , \59192 , \59202 );
xor \g132587/U$1_r1 ( \59204 , \59175 , \59203 );
xor \g132509/U$1_r1 ( \59205 , \59162 , \59204 );
xor \g132360/U$1_r1 ( \59206 , \59145 , \59205 );
xor \g456159/U$1_r1 ( \59207 , \59104 , \59206 );
xor \g456159/U$1_r2 ( \59208 , \59100 , \59207 );
xor \g131614/U$1 ( \59209 , \58911 , \59042 );
xor \g131614/U$1_r1 ( \59210 , \59209 , \59061 );
and \g131587/U$2 ( \59211 , \59208 , \59210 );
and \g131494/U$3 ( \59212 , \59072 , \59211 );
and \g131494/U$5 ( \59213 , \59064 , \59071 );
or \g131494/U$2 ( \59214 , \59212 , \59213 );
xor \g132515/U$4 ( \59215 , \59089 , \59093 );
and \g132515/U$3 ( \59216 , \59215 , \59098 );
and \g132515/U$5 ( \59217 , \59089 , \59093 );
or \g132515/U$2 ( \59218 , \59216 , \59217 );
not \g132931/U$3 ( \59219 , \49925 );
and \g132965/U$2 ( \59220 , \55884 , \50160 );
and \g132965/U$3 ( \59221 , \50159 , \55707 );
nor \g132965/U$1 ( \59222 , \59220 , \59221 );
not \g132931/U$4 ( \59223 , \59222 );
or \g132931/U$2 ( \59224 , \59219 , \59223 );
or \g132931/U$5 ( \59225 , \59222 , \49925 );
nand \g132931/U$1 ( \59226 , \59224 , \59225 );
not \g133041/U$3 ( \59227 , \49568 );
and \g133075/U$2 ( \59228 , \56446 , \49813 );
and \g133075/U$3 ( \59229 , \49812 , \56167 );
nor \g133075/U$1 ( \59230 , \59228 , \59229 );
not \g133041/U$4 ( \59231 , \59230 );
or \g133041/U$2 ( \59232 , \59227 , \59231 );
or \g133041/U$5 ( \59233 , \59230 , \49568 );
nand \g133041/U$1 ( \59234 , \59232 , \59233 );
xor \g132589/U$1 ( \59235 , \59226 , \59234 );
not \g132987/U$3 ( \59236 , \48685 );
and \g133017/U$2 ( \59237 , \48858 , \56349 );
and \g133017/U$3 ( \59238 , \56411 , \48860 );
nor \g133017/U$1 ( \59239 , \59237 , \59238 );
not \g132987/U$4 ( \59240 , \59239 );
or \g132987/U$2 ( \59241 , \59236 , \59240 );
or \g132987/U$5 ( \59242 , \59239 , \48685 );
nand \g132987/U$1 ( \59243 , \59241 , \59242 );
not \g133061/U$3 ( \59244 , \49014 );
and \g133106/U$2 ( \59245 , \49075 , \56347 );
and \g133106/U$3 ( \59246 , \56359 , \49074 );
nor \g133106/U$1 ( \59247 , \59245 , \59246 );
not \g133061/U$4 ( \59248 , \59247 );
or \g133061/U$2 ( \59249 , \59244 , \59248 );
or \g133061/U$5 ( \59250 , \59247 , \49014 );
nand \g133061/U$1 ( \59251 , \59249 , \59250 );
xor \g132691/U$1 ( \59252 , \59243 , \59251 );
and \g132773/U$2 ( \59253 , \59193 , \59201 );
xor \g132691/U$1_r1 ( \59254 , \59252 , \59253 );
xor \g132589/U$1_r1 ( \59255 , \59235 , \59254 );
not \g132533/U$3 ( \59256 , \51124 );
and \g132576/U$2 ( \59257 , \54251 , \51517 );
and \g132576/U$3 ( \59258 , \51518 , \54529 );
nor \g132576/U$1 ( \59259 , \59257 , \59258 );
not \g132533/U$4 ( \59260 , \59259 );
or \g132533/U$2 ( \59261 , \59256 , \59260 );
or \g132533/U$5 ( \59262 , \59259 , \51124 );
nand \g132533/U$1 ( \59263 , \59261 , \59262 );
xor \g456157/U$9 ( \59264 , \59255 , \59263 );
and \g132436/U$2 ( \59265 , \54185 , \52273 );
and \g132436/U$3 ( \59266 , \52270 , \54015 );
nor \g132436/U$1 ( \59267 , \59265 , \59266 );
and \g132346/U$2 ( \59268 , \59267 , \51513 );
not \g132346/U$4 ( \59269 , \59267 );
and \g132346/U$3 ( \59270 , \59269 , \51120 );
nor \g132346/U$1 ( \59271 , \59268 , \59270 );
xor \g456157/U$9_r1 ( \59272 , \59264 , \59271 );
and \g456157/U$8 ( \59273 , \59218 , \59272 );
xor \g132360/U$4 ( \59274 , \59111 , \59144 );
and \g132360/U$3 ( \59275 , \59274 , \59205 );
and \g132360/U$5 ( \59276 , \59111 , \59144 );
or \g132360/U$2 ( \59277 , \59275 , \59276 );
xor \g456157/U$11 ( \59278 , \59255 , \59263 );
xor \g456157/U$11_r1 ( \59279 , \59278 , \59271 );
and \g456157/U$10 ( \59280 , \59277 , \59279 );
and \g456157/U$12 ( \59281 , \59218 , \59277 );
or \g456157/U$7 ( \59282 , \59273 , \59280 , \59281 );
and \g132308/U$2 ( \59283 , \53848 , \52270 );
and \g132308/U$3 ( \59284 , \52273 , \54015 );
nor \g132308/U$1 ( \59285 , \59283 , \59284 );
and \g132254/U$2 ( \59286 , \59285 , \51513 );
not \g132254/U$4 ( \59287 , \59285 );
and \g132254/U$3 ( \59288 , \59287 , \51120 );
nor \g132254/U$1 ( \59289 , \59286 , \59288 );
xor \g132631/U$4 ( \59290 , \59115 , \59123 );
and \g132631/U$3 ( \59291 , \59290 , \59143 );
and \g132631/U$5 ( \59292 , \59115 , \59123 );
or \g132631/U$2 ( \59293 , \59291 , \59292 );
not \g132823/U$3 ( \59294 , \50362 );
and \g132857/U$2 ( \59295 , \55127 , \50587 );
and \g132857/U$3 ( \59296 , \50588 , \55460 );
nor \g132857/U$1 ( \59297 , \59295 , \59296 );
not \g132823/U$4 ( \59298 , \59297 );
or \g132823/U$2 ( \59299 , \59294 , \59298 );
or \g132823/U$5 ( \59300 , \59297 , \50362 );
nand \g132823/U$1 ( \59301 , \59299 , \59300 );
xor \g456161/U$5 ( \59302 , \59293 , \59301 );
xor \g132587/U$4 ( \59303 , \59166 , \59174 );
and \g132587/U$3 ( \59304 , \59303 , \59203 );
and \g132587/U$5 ( \59305 , \59166 , \59174 );
or \g132587/U$2 ( \59306 , \59304 , \59305 );
and \g456161/U$4 ( \59307 , \59302 , \59306 );
and \g456161/U$6 ( \59308 , \59293 , \59301 );
or \g456161/U$3 ( \59309 , \59307 , \59308 );
xor \g132144/U$1 ( \59310 , \59289 , \59309 );
xor \g456157/U$5 ( \59311 , \59255 , \59263 );
and \g456157/U$4 ( \59312 , \59311 , \59271 );
and \g456157/U$6 ( \59313 , \59255 , \59263 );
or \g456157/U$3 ( \59314 , \59312 , \59313 );
xor \g132144/U$1_r1 ( \59315 , \59310 , \59314 );
xor \g132027/U$1 ( \59316 , \59282 , \59315 );
xor \g132509/U$4 ( \59317 , \59153 , \59161 );
and \g132509/U$3 ( \59318 , \59317 , \59204 );
and \g132509/U$5 ( \59319 , \59153 , \59161 );
or \g132509/U$2 ( \59320 , \59318 , \59319 );
xor \g456161/U$9 ( \59321 , \59293 , \59301 );
xor \g456161/U$9_r1 ( \59322 , \59321 , \59306 );
and \g456161/U$8 ( \59323 , \59320 , \59322 );
not \g132684/U$3 ( \59324 , \50759 );
and \g132727/U$2 ( \59325 , \54853 , \51055 );
and \g132727/U$3 ( \59326 , \51053 , \54537 );
nor \g132727/U$1 ( \59327 , \59325 , \59326 );
not \g132684/U$4 ( \59328 , \59327 );
or \g132684/U$2 ( \59329 , \59324 , \59328 );
or \g132684/U$5 ( \59330 , \59327 , \50759 );
nand \g132684/U$1 ( \59331 , \59329 , \59330 );
xor \g132791/U$4 ( \59332 , \59132 , \59140 );
and \g132791/U$3 ( \59333 , \59332 , \59142 );
and \g132791/U$5 ( \59334 , \59132 , \59140 );
or \g132791/U$2 ( \59335 , \59333 , \59334 );
xor \g132505/U$1 ( \59336 , \59331 , \59335 );
not \g132902/U$3 ( \59337 , \48483 );
and \g132946/U$2 ( \59338 , \48478 , \56368 );
and \g132946/U$3 ( \59339 , \56370 , \48479 );
nor \g132946/U$1 ( \59340 , \59338 , \59339 );
not \g132902/U$4 ( \59341 , \59340 );
or \g132902/U$2 ( \59342 , \59337 , \59341 );
or \g132902/U$5 ( \59343 , \59340 , \48483 );
nand \g132902/U$1 ( \59344 , \59342 , \59343 );
not \g132821/U$3 ( \59345 , \48323 );
and \g132854/U$2 ( \59346 , \48335 , \56377 );
and \g132854/U$3 ( \59347 , \56379 , \48334 );
nor \g132854/U$1 ( \59348 , \59346 , \59347 );
not \g132821/U$4 ( \59349 , \59348 );
or \g132821/U$2 ( \59350 , \59345 , \59349 );
or \g132821/U$5 ( \59351 , \59348 , \48323 );
nand \g132821/U$1 ( \59352 , \59350 , \59351 );
xor \g132776/U$1 ( \59353 , \59344 , \59352 );
not \g133131/U$3 ( \59354 , \49233 );
and \g133164/U$2 ( \59355 , \49405 , \56357 );
and \g133164/U$3 ( \59356 , \49403 , \56448 );
nor \g133164/U$1 ( \59357 , \59355 , \59356 );
not \g133131/U$4 ( \59358 , \59357 );
or \g133131/U$2 ( \59359 , \59354 , \59358 );
or \g133131/U$5 ( \59360 , \59357 , \49233 );
nand \g133131/U$1 ( \59361 , \59359 , \59360 );
xor \g132584/U$1 ( \59362 , \59353 , \59361 );
xor \g132690/U$4 ( \59363 , \59183 , \59191 );
and \g132690/U$3 ( \59364 , \59363 , \59202 );
and \g132690/U$5 ( \59365 , \59183 , \59191 );
or \g132690/U$2 ( \59366 , \59364 , \59365 );
xor \g132584/U$1_r1 ( \59367 , \59362 , \59366 );
xor \g132505/U$1_r1 ( \59368 , \59336 , \59367 );
xor \g456161/U$11 ( \59369 , \59293 , \59301 );
xor \g456161/U$11_r1 ( \59370 , \59369 , \59306 );
and \g456161/U$10 ( \59371 , \59368 , \59370 );
and \g456161/U$12 ( \59372 , \59320 , \59368 );
or \g456161/U$7 ( \59373 , \59323 , \59371 , \59372 );
xor \g132589/U$4 ( \59374 , \59226 , \59234 );
and \g132589/U$3 ( \59375 , \59374 , \59254 );
and \g132589/U$5 ( \59376 , \59226 , \59234 );
or \g132589/U$2 ( \59377 , \59375 , \59376 );
not \g132617/U$3 ( \59378 , \50759 );
and \g132662/U$2 ( \59379 , \54537 , \51055 );
and \g132662/U$3 ( \59380 , \51053 , \54529 );
nor \g132662/U$1 ( \59381 , \59379 , \59380 );
not \g132617/U$4 ( \59382 , \59381 );
or \g132617/U$2 ( \59383 , \59378 , \59382 );
or \g132617/U$5 ( \59384 , \59381 , \50759 );
nand \g132617/U$1 ( \59385 , \59383 , \59384 );
xor \g132392/U$1 ( \59386 , \59377 , \59385 );
xor \g132505/U$4 ( \59387 , \59331 , \59335 );
and \g132505/U$3 ( \59388 , \59387 , \59367 );
and \g132505/U$5 ( \59389 , \59331 , \59335 );
or \g132505/U$2 ( \59390 , \59388 , \59389 );
xor \g132392/U$1_r1 ( \59391 , \59386 , \59390 );
xor \g132143/U$1 ( \59392 , \59373 , \59391 );
not \g132985/U$3 ( \59393 , \48685 );
and \g133025/U$2 ( \59394 , \48858 , \56347 );
and \g133025/U$3 ( \59395 , \56349 , \48860 );
nor \g133025/U$1 ( \59396 , \59394 , \59395 );
not \g132985/U$4 ( \59397 , \59396 );
or \g132985/U$2 ( \59398 , \59393 , \59397 );
or \g132985/U$5 ( \59399 , \59396 , \48685 );
nand \g132985/U$1 ( \59400 , \59398 , \59399 );
not \g133066/U$3 ( \59401 , \49014 );
and \g133099/U$2 ( \59402 , \49074 , \56357 );
and \g133099/U$3 ( \59403 , \56359 , \49075 );
nor \g133099/U$1 ( \59404 , \59402 , \59403 );
not \g133066/U$4 ( \59405 , \59404 );
or \g133066/U$2 ( \59406 , \59401 , \59405 );
or \g133066/U$5 ( \59407 , \59404 , \49014 );
nand \g133066/U$1 ( \59408 , \59406 , \59407 );
xor \g132694/U$1 ( \59409 , \59400 , \59408 );
and \g132776/U$2 ( \59410 , \59344 , \59352 );
xor \g132694/U$1_r1 ( \59411 , \59409 , \59410 );
not \g132986/U$3 ( \59412 , \49568 );
and \g133023/U$2 ( \59413 , \56167 , \49813 );
and \g133023/U$3 ( \59414 , \49812 , \55884 );
nor \g133023/U$1 ( \59415 , \59413 , \59414 );
not \g132986/U$4 ( \59416 , \59415 );
or \g132986/U$2 ( \59417 , \59412 , \59416 );
or \g132986/U$5 ( \59418 , \59415 , \49568 );
nand \g132986/U$1 ( \59419 , \59417 , \59418 );
xor \g456160/U$2 ( \59420 , \59411 , \59419 );
xor \g132584/U$4 ( \59421 , \59353 , \59361 );
and \g132584/U$3 ( \59422 , \59421 , \59366 );
and \g132584/U$5 ( \59423 , \59353 , \59361 );
or \g132584/U$2 ( \59424 , \59422 , \59423 );
xor \g456160/U$1 ( \59425 , \59420 , \59424 );
not \g132456/U$3 ( \59426 , \51124 );
and \g132503/U$2 ( \59427 , \54185 , \51517 );
and \g132503/U$3 ( \59428 , \51518 , \54251 );
nor \g132503/U$1 ( \59429 , \59427 , \59428 );
not \g132456/U$4 ( \59430 , \59429 );
or \g132456/U$2 ( \59431 , \59426 , \59430 );
or \g132456/U$5 ( \59432 , \59429 , \51124 );
nand \g132456/U$1 ( \59433 , \59431 , \59432 );
not \g132745/U$3 ( \59434 , \50362 );
and \g132785/U$2 ( \59435 , \54853 , \50587 );
and \g132785/U$3 ( \59436 , \50588 , \55127 );
nor \g132785/U$1 ( \59437 , \59435 , \59436 );
not \g132745/U$4 ( \59438 , \59437 );
or \g132745/U$2 ( \59439 , \59434 , \59438 );
or \g132745/U$5 ( \59440 , \59437 , \50362 );
nand \g132745/U$1 ( \59441 , \59439 , \59440 );
not \g132876/U$3 ( \59442 , \49925 );
and \g132915/U$2 ( \59443 , \55460 , \50159 );
and \g132915/U$3 ( \59444 , \50160 , \55707 );
nor \g132915/U$1 ( \59445 , \59443 , \59444 );
not \g132876/U$4 ( \59446 , \59445 );
or \g132876/U$2 ( \59447 , \59442 , \59446 );
or \g132876/U$5 ( \59448 , \59445 , \49925 );
nand \g132876/U$1 ( \59449 , \59447 , \59448 );
xor \g132388/U$1 ( \59450 , \59441 , \59449 );
xor \g132691/U$4 ( \59451 , \59243 , \59251 );
and \g132691/U$3 ( \59452 , \59451 , \59253 );
and \g132691/U$5 ( \59453 , \59243 , \59251 );
or \g132691/U$2 ( \59454 , \59452 , \59453 );
not \g133089/U$3 ( \59455 , \49233 );
and \g133117/U$2 ( \59456 , \56446 , \49403 );
and \g133117/U$3 ( \59457 , \56448 , \49405 );
nor \g133117/U$1 ( \59458 , \59456 , \59457 );
not \g133089/U$4 ( \59459 , \59458 );
or \g133089/U$2 ( \59460 , \59455 , \59459 );
or \g133089/U$5 ( \59461 , \59458 , \49233 );
nand \g133089/U$1 ( \59462 , \59460 , \59461 );
xor \g132507/U$1 ( \59463 , \59454 , \59462 );
not \g132716/U$3 ( \59464 , \48159 );
and \g132751/U$2 ( \59465 , \48155 , \47026 );
and \g132751/U$3 ( \59466 , \56377 , \48154 );
nor \g132751/U$1 ( \59467 , \59465 , \59466 );
not \g132716/U$4 ( \59468 , \59467 );
or \g132716/U$2 ( \59469 , \59464 , \59468 );
or \g132716/U$5 ( \59470 , \59467 , \48159 );
nand \g132716/U$1 ( \59471 , \59469 , \59470 );
not \g132900/U$3 ( \59472 , \48483 );
and \g132945/U$2 ( \59473 , \48478 , \56411 );
and \g132945/U$3 ( \59474 , \56368 , \48479 );
nor \g132945/U$1 ( \59475 , \59473 , \59474 );
not \g132900/U$4 ( \59476 , \59475 );
or \g132900/U$2 ( \59477 , \59472 , \59476 );
or \g132900/U$5 ( \59478 , \59475 , \48483 );
nand \g132900/U$1 ( \59479 , \59477 , \59478 );
xor \g132588/U$1 ( \59480 , \59471 , \59479 );
not \g132819/U$3 ( \59481 , \48323 );
and \g132853/U$2 ( \59482 , \48334 , \56370 );
and \g132853/U$3 ( \59483 , \56379 , \48335 );
nor \g132853/U$1 ( \59484 , \59482 , \59483 );
not \g132819/U$4 ( \59485 , \59484 );
or \g132819/U$2 ( \59486 , \59481 , \59485 );
or \g132819/U$5 ( \59487 , \59484 , \48323 );
nand \g132819/U$1 ( \59488 , \59486 , \59487 );
and \g132735/U$2 ( \59489 , \48159 , \59070 );
xor \g132687/U$1 ( \59490 , \59488 , \59489 );
xor \g132588/U$1_r1 ( \59491 , \59480 , \59490 );
xor \g132507/U$1_r1 ( \59492 , \59463 , \59491 );
xor \g132388/U$1_r1 ( \59493 , \59450 , \59492 );
xor \g456160/U$1_r1 ( \59494 , \59433 , \59493 );
xor \g456160/U$1_r2 ( \59495 , \59425 , \59494 );
xor \g132143/U$1_r1 ( \59496 , \59392 , \59495 );
xor \g132027/U$1_r1 ( \59497 , \59316 , \59496 );
xor \g131343/U$4 ( \59498 , \59214 , \59497 );
xor \g456159/U$9 ( \59499 , \59076 , \59080 );
xor \g456159/U$9_r1 ( \59500 , \59499 , \59099 );
and \g456159/U$8 ( \59501 , \59104 , \59500 );
xor \g456159/U$11 ( \59502 , \59076 , \59080 );
xor \g456159/U$11_r1 ( \59503 , \59502 , \59099 );
and \g456159/U$10 ( \59504 , \59206 , \59503 );
and \g456159/U$12 ( \59505 , \59104 , \59206 );
or \g456159/U$7 ( \59506 , \59501 , \59504 , \59505 );
xor \g456161/U$2 ( \59507 , \59293 , \59301 );
xor \g456161/U$1 ( \59508 , \59507 , \59306 );
xor \g456161/U$1_r1 ( \59509 , \59320 , \59368 );
xor \g456161/U$1_r2 ( \59510 , \59508 , \59509 );
xor \g456159/U$5 ( \59511 , \59076 , \59080 );
and \g456159/U$4 ( \59512 , \59511 , \59099 );
and \g456159/U$6 ( \59513 , \59076 , \59080 );
or \g456159/U$3 ( \59514 , \59512 , \59513 );
xor \g456121/U$9 ( \59515 , \59510 , \59514 );
xor \g456157/U$2 ( \59516 , \59255 , \59263 );
xor \g456157/U$1 ( \59517 , \59516 , \59271 );
xor \g456157/U$1_r1 ( \59518 , \59218 , \59277 );
xor \g456157/U$1_r2 ( \59519 , \59517 , \59518 );
xor \g456121/U$9_r1 ( \59520 , \59515 , \59519 );
and \g456121/U$8 ( \59521 , \59506 , \59520 );
xor \g131494/U$1 ( \59522 , \59064 , \59071 );
xor \g131494/U$1_r1 ( \59523 , \59522 , \59211 );
xor \g456121/U$11 ( \59524 , \59510 , \59514 );
xor \g456121/U$11_r1 ( \59525 , \59524 , \59519 );
and \g456121/U$10 ( \59526 , \59523 , \59525 );
and \g456121/U$12 ( \59527 , \59506 , \59523 );
or \g456121/U$7 ( \59528 , \59521 , \59526 , \59527 );
and \g131343/U$3 ( \59529 , \59498 , \59528 );
and \g131343/U$5 ( \59530 , \59214 , \59497 );
or \g131343/U$2 ( \59531 , \59529 , \59530 );
nand \g132700/U$1 ( \59532 , \47026 , \48063 );
not \g132682/U$3 ( \59533 , \59532 );
not \g132682/U$4 ( \59534 , \47997 );
or \g132682/U$2 ( \59535 , \59533 , \59534 );
or \g132682/U$5 ( \59536 , \47997 , \59532 );
nand \g132682/U$1 ( \59537 , \59535 , \59536 );
xor \g132636/U$1 ( \59538 , \47997 , \59537 );
xor \g131225/U$4 ( \59539 , \59531 , \59538 );
xor \g456121/U$5 ( \59540 , \59510 , \59514 );
and \g456121/U$4 ( \59541 , \59540 , \59519 );
and \g456121/U$6 ( \59542 , \59510 , \59514 );
or \g456121/U$3 ( \59543 , \59541 , \59542 );
xor \g131343/U$1 ( \59544 , \59214 , \59497 );
xor \g131343/U$1_r1 ( \59545 , \59544 , \59528 );
and \g131306/U$2 ( \59546 , \59543 , \59545 );
and \g131225/U$3 ( \59547 , \59539 , \59546 );
and \g131225/U$5 ( \59548 , \59531 , \59538 );
or \g131225/U$2 ( \59549 , \59547 , \59548 );
xor \g132143/U$4 ( \59550 , \59373 , \59391 );
and \g132143/U$3 ( \59551 , \59550 , \59495 );
and \g132143/U$5 ( \59552 , \59373 , \59391 );
or \g132143/U$2 ( \59553 , \59551 , \59552 );
xor \g456160/U$5 ( \59554 , \59411 , \59419 );
and \g456160/U$4 ( \59555 , \59554 , \59424 );
and \g456160/U$6 ( \59556 , \59411 , \59419 );
or \g456160/U$3 ( \59557 , \59555 , \59556 );
not \g132531/U$3 ( \59558 , \50759 );
and \g132575/U$2 ( \59559 , \54251 , \51053 );
and \g132575/U$3 ( \59560 , \51055 , \54529 );
nor \g132575/U$1 ( \59561 , \59559 , \59560 );
not \g132531/U$4 ( \59562 , \59561 );
or \g132531/U$2 ( \59563 , \59558 , \59562 );
or \g132531/U$5 ( \59564 , \59561 , \50759 );
nand \g132531/U$1 ( \59565 , \59563 , \59564 );
xor \g456158/U$2 ( \59566 , \59557 , \59565 );
not \g132344/U$3 ( \59567 , \51124 );
and \g132435/U$2 ( \59568 , \54185 , \51518 );
and \g132435/U$3 ( \59569 , \51517 , \54015 );
nor \g132435/U$1 ( \59570 , \59568 , \59569 );
not \g132344/U$4 ( \59571 , \59570 );
or \g132344/U$2 ( \59572 , \59567 , \59571 );
or \g132344/U$5 ( \59573 , \59570 , \51124 );
nand \g132344/U$1 ( \59574 , \59572 , \59573 );
xor \g456158/U$1 ( \59575 , \59566 , \59574 );
xor \g132392/U$4 ( \59576 , \59377 , \59385 );
and \g132392/U$3 ( \59577 , \59576 , \59390 );
and \g132392/U$5 ( \59578 , \59377 , \59385 );
or \g132392/U$2 ( \59579 , \59577 , \59578 );
xor \g132507/U$4 ( \59580 , \59454 , \59462 );
and \g132507/U$3 ( \59581 , \59580 , \59491 );
and \g132507/U$5 ( \59582 , \59454 , \59462 );
or \g132507/U$2 ( \59583 , \59581 , \59582 );
not \g132677/U$3 ( \59584 , \50362 );
and \g132724/U$2 ( \59585 , \54853 , \50588 );
and \g132724/U$3 ( \59586 , \50587 , \54537 );
nor \g132724/U$1 ( \59587 , \59585 , \59586 );
not \g132677/U$4 ( \59588 , \59587 );
or \g132677/U$2 ( \59589 , \59584 , \59588 );
or \g132677/U$5 ( \59590 , \59587 , \50362 );
nand \g132677/U$1 ( \59591 , \59589 , \59590 );
xor \g132389/U$1 ( \59592 , \59583 , \59591 );
xor \g132694/U$4 ( \59593 , \59400 , \59408 );
and \g132694/U$3 ( \59594 , \59593 , \59410 );
and \g132694/U$5 ( \59595 , \59400 , \59408 );
or \g132694/U$2 ( \59596 , \59594 , \59595 );
not \g133038/U$3 ( \59597 , \49233 );
and \g133070/U$2 ( \59598 , \56446 , \49405 );
and \g133070/U$3 ( \59599 , \49403 , \56167 );
nor \g133070/U$1 ( \59600 , \59598 , \59599 );
not \g133038/U$4 ( \59601 , \59600 );
or \g133038/U$2 ( \59602 , \59597 , \59601 );
or \g133038/U$5 ( \59603 , \59600 , \49233 );
nand \g133038/U$1 ( \59604 , \59602 , \59603 );
xor \g132511/U$1 ( \59605 , \59596 , \59604 );
not \g132904/U$3 ( \59606 , \48483 );
and \g132948/U$2 ( \59607 , \48478 , \56349 );
and \g132948/U$3 ( \59608 , \56411 , \48479 );
nor \g132948/U$1 ( \59609 , \59607 , \59608 );
not \g132904/U$4 ( \59610 , \59609 );
or \g132904/U$2 ( \59611 , \59606 , \59610 );
or \g132904/U$5 ( \59612 , \59609 , \48483 );
nand \g132904/U$1 ( \59613 , \59611 , \59612 );
not \g133000/U$3 ( \59614 , \48685 );
and \g133019/U$2 ( \59615 , \48860 , \56347 );
and \g133019/U$3 ( \59616 , \56359 , \48858 );
nor \g133019/U$1 ( \59617 , \59615 , \59616 );
not \g133000/U$4 ( \59618 , \59617 );
or \g133000/U$2 ( \59619 , \59614 , \59618 );
or \g133000/U$5 ( \59620 , \59617 , \48685 );
nand \g133000/U$1 ( \59621 , \59619 , \59620 );
xor \g132585/U$1 ( \59622 , \59613 , \59621 );
and \g132687/U$2 ( \59623 , \59488 , \59489 );
xor \g132585/U$1_r1 ( \59624 , \59622 , \59623 );
xor \g132511/U$1_r1 ( \59625 , \59605 , \59624 );
xor \g132389/U$1_r1 ( \59626 , \59592 , \59625 );
xor \g456158/U$1_r1 ( \59627 , \59579 , \59626 );
xor \g456158/U$1_r2 ( \59628 , \59575 , \59627 );
xor \g456101/U$5 ( \59629 , \59553 , \59628 );
xor \g456160/U$9 ( \59630 , \59411 , \59419 );
xor \g456160/U$9_r1 ( \59631 , \59630 , \59424 );
and \g456160/U$8 ( \59632 , \59433 , \59631 );
xor \g456160/U$11 ( \59633 , \59411 , \59419 );
xor \g456160/U$11_r1 ( \59634 , \59633 , \59424 );
and \g456160/U$10 ( \59635 , \59493 , \59634 );
and \g456160/U$12 ( \59636 , \59433 , \59493 );
or \g456160/U$7 ( \59637 , \59632 , \59635 , \59636 );
xor \g132144/U$4 ( \59638 , \59289 , \59309 );
and \g132144/U$3 ( \59639 , \59638 , \59314 );
and \g132144/U$5 ( \59640 , \59289 , \59309 );
or \g132144/U$2 ( \59641 , \59639 , \59640 );
xor \g131976/U$1 ( \59642 , \59637 , \59641 );
xor \g132388/U$4 ( \59643 , \59441 , \59449 );
and \g132388/U$3 ( \59644 , \59643 , \59492 );
and \g132388/U$5 ( \59645 , \59441 , \59449 );
or \g132388/U$2 ( \59646 , \59644 , \59645 );
and \g132207/U$2 ( \59647 , \53610 , \52270 );
and \g132207/U$3 ( \59648 , \52273 , \53848 );
nor \g132207/U$1 ( \59649 , \59647 , \59648 );
and \g132151/U$2 ( \59650 , \59649 , \51513 );
not \g132151/U$4 ( \59651 , \59649 );
and \g132151/U$3 ( \59652 , \59651 , \51120 );
nor \g132151/U$1 ( \59653 , \59650 , \59652 );
xor \g132096/U$1 ( \59654 , \59646 , \59653 );
not \g132817/U$3 ( \59655 , \49925 );
and \g132851/U$2 ( \59656 , \55127 , \50159 );
and \g132851/U$3 ( \59657 , \50160 , \55460 );
nor \g132851/U$1 ( \59658 , \59656 , \59657 );
not \g132817/U$4 ( \59659 , \59658 );
or \g132817/U$2 ( \59660 , \59655 , \59659 );
or \g132817/U$5 ( \59661 , \59658 , \49925 );
nand \g132817/U$1 ( \59662 , \59660 , \59661 );
not \g132929/U$3 ( \59663 , \49568 );
and \g132963/U$2 ( \59664 , \55884 , \49813 );
and \g132963/U$3 ( \59665 , \49812 , \55707 );
nor \g132963/U$1 ( \59666 , \59664 , \59665 );
not \g132929/U$4 ( \59667 , \59666 );
or \g132929/U$2 ( \59668 , \59663 , \59667 );
or \g132929/U$5 ( \59669 , \59666 , \49568 );
nand \g132929/U$1 ( \59670 , \59668 , \59669 );
xor \g132394/U$1 ( \59671 , \59662 , \59670 );
not \g132818/U$3 ( \59672 , \48323 );
and \g132852/U$2 ( \59673 , \48334 , \56368 );
and \g132852/U$3 ( \59674 , \56370 , \48335 );
nor \g132852/U$1 ( \59675 , \59673 , \59674 );
not \g132818/U$4 ( \59676 , \59675 );
or \g132818/U$2 ( \59677 , \59672 , \59676 );
or \g132818/U$5 ( \59678 , \59675 , \48323 );
nand \g132818/U$1 ( \59679 , \59677 , \59678 );
not \g132715/U$3 ( \59680 , \48159 );
and \g132763/U$2 ( \59681 , \48155 , \56377 );
and \g132763/U$3 ( \59682 , \56379 , \48154 );
nor \g132763/U$1 ( \59683 , \59681 , \59682 );
not \g132715/U$4 ( \59684 , \59683 );
or \g132715/U$2 ( \59685 , \59680 , \59684 );
or \g132715/U$5 ( \59686 , \59683 , \48159 );
nand \g132715/U$1 ( \59687 , \59685 , \59686 );
xor \g132672/U$1 ( \59688 , \59679 , \59687 );
not \g133060/U$3 ( \59689 , \49014 );
and \g133098/U$2 ( \59690 , \49075 , \56357 );
and \g133098/U$3 ( \59691 , \56448 , \49074 );
nor \g133098/U$1 ( \59692 , \59690 , \59691 );
not \g133060/U$4 ( \59693 , \59692 );
or \g133060/U$2 ( \59694 , \59689 , \59693 );
or \g133060/U$5 ( \59695 , \59692 , \49014 );
nand \g133060/U$1 ( \59696 , \59694 , \59695 );
xor \g132508/U$1 ( \59697 , \59688 , \59696 );
xor \g132588/U$4 ( \59698 , \59471 , \59479 );
and \g132588/U$3 ( \59699 , \59698 , \59490 );
and \g132588/U$5 ( \59700 , \59471 , \59479 );
or \g132588/U$2 ( \59701 , \59699 , \59700 );
xor \g132508/U$1_r1 ( \59702 , \59697 , \59701 );
xor \g132394/U$1_r1 ( \59703 , \59671 , \59702 );
xor \g132096/U$1_r1 ( \59704 , \59654 , \59703 );
xor \g131976/U$1_r1 ( \59705 , \59642 , \59704 );
and \g456101/U$4 ( \59706 , \59629 , \59705 );
and \g456101/U$6 ( \59707 , \59553 , \59628 );
or \g456101/U$3 ( \59708 , \59706 , \59707 );
xor \g131041/U$4 ( \59709 , \59549 , \59708 );
xor \g132027/U$4 ( \59710 , \59282 , \59315 );
and \g132027/U$3 ( \59711 , \59710 , \59496 );
and \g132027/U$5 ( \59712 , \59282 , \59315 );
or \g132027/U$2 ( \59713 , \59711 , \59712 );
xor \g456101/U$9 ( \59714 , \59553 , \59628 );
xor \g456101/U$9_r1 ( \59715 , \59714 , \59705 );
and \g456101/U$8 ( \59716 , \59713 , \59715 );
xor \g131225/U$1 ( \59717 , \59531 , \59538 );
xor \g131225/U$1_r1 ( \59718 , \59717 , \59546 );
xor \g456101/U$11 ( \59719 , \59553 , \59628 );
xor \g456101/U$11_r1 ( \59720 , \59719 , \59705 );
and \g456101/U$10 ( \59721 , \59718 , \59720 );
and \g456101/U$12 ( \59722 , \59713 , \59718 );
or \g456101/U$7 ( \59723 , \59716 , \59721 , \59722 );
and \g131041/U$3 ( \59724 , \59709 , \59723 );
and \g131041/U$5 ( \59725 , \59549 , \59708 );
or \g131041/U$2 ( \59726 , \59724 , \59725 );
nand \g132590/U$1 ( \59727 , \47026 , \47930 );
not \g132564/U$3 ( \59728 , \59727 );
not \g132564/U$4 ( \59729 , \47935 );
or \g132564/U$2 ( \59730 , \59728 , \59729 );
or \g132564/U$5 ( \59731 , \47935 , \59727 );
nand \g132564/U$1 ( \59732 , \59730 , \59731 );
xor \g132514/U$1 ( \59733 , \47935 , \59732 );
xor \g130916/U$4 ( \59734 , \59726 , \59733 );
xor \g131976/U$4 ( \59735 , \59637 , \59641 );
and \g131976/U$3 ( \59736 , \59735 , \59704 );
and \g131976/U$5 ( \59737 , \59637 , \59641 );
or \g131976/U$2 ( \59738 , \59736 , \59737 );
xor \g132511/U$4 ( \59739 , \59596 , \59604 );
and \g132511/U$3 ( \59740 , \59739 , \59624 );
and \g132511/U$5 ( \59741 , \59596 , \59604 );
or \g132511/U$2 ( \59742 , \59740 , \59741 );
not \g132616/U$3 ( \59743 , \50362 );
and \g132660/U$2 ( \59744 , \54537 , \50588 );
and \g132660/U$3 ( \59745 , \50587 , \54529 );
nor \g132660/U$1 ( \59746 , \59744 , \59745 );
not \g132616/U$4 ( \59747 , \59746 );
or \g132616/U$2 ( \59748 , \59743 , \59747 );
or \g132616/U$5 ( \59749 , \59746 , \50362 );
nand \g132616/U$1 ( \59750 , \59748 , \59749 );
xor \g456154/U$2 ( \59751 , \59742 , \59750 );
xor \g132394/U$4 ( \59752 , \59662 , \59670 );
and \g132394/U$3 ( \59753 , \59752 , \59702 );
and \g132394/U$5 ( \59754 , \59662 , \59670 );
or \g132394/U$2 ( \59755 , \59753 , \59754 );
xor \g456154/U$1 ( \59756 , \59751 , \59755 );
xor \g456158/U$5 ( \59757 , \59557 , \59565 );
and \g456158/U$4 ( \59758 , \59757 , \59574 );
and \g456158/U$6 ( \59759 , \59557 , \59565 );
or \g456158/U$3 ( \59760 , \59758 , \59759 );
xor \g132096/U$4 ( \59761 , \59646 , \59653 );
and \g132096/U$3 ( \59762 , \59761 , \59703 );
and \g132096/U$5 ( \59763 , \59646 , \59653 );
or \g132096/U$2 ( \59764 , \59762 , \59763 );
xor \g456154/U$1_r1 ( \59765 , \59760 , \59764 );
xor \g456154/U$1_r2 ( \59766 , \59756 , \59765 );
xor \g131806/U$1 ( \59767 , \59738 , \59766 );
xor \g132389/U$4 ( \59768 , \59583 , \59591 );
and \g132389/U$3 ( \59769 , \59768 , \59625 );
and \g132389/U$5 ( \59770 , \59583 , \59591 );
or \g132389/U$2 ( \59771 , \59769 , \59770 );
not \g132253/U$3 ( \59772 , \51124 );
and \g132307/U$2 ( \59773 , \53848 , \51517 );
and \g132307/U$3 ( \59774 , \51518 , \54015 );
nor \g132307/U$1 ( \59775 , \59773 , \59774 );
not \g132253/U$4 ( \59776 , \59775 );
or \g132253/U$2 ( \59777 , \59772 , \59776 );
or \g132253/U$5 ( \59778 , \59775 , \51124 );
nand \g132253/U$1 ( \59779 , \59777 , \59778 );
xor \g456149/U$2 ( \59780 , \59771 , \59779 );
and \g132134/U$2 ( \59781 , \53610 , \52273 );
and \g132134/U$3 ( \59782 , \52270 , \53300 );
nor \g132134/U$1 ( \59783 , \59781 , \59782 );
and \g132087/U$2 ( \59784 , \59783 , \51513 );
not \g132087/U$4 ( \59785 , \59783 );
and \g132087/U$3 ( \59786 , \59785 , \51120 );
nor \g132087/U$1 ( \59787 , \59784 , \59786 );
xor \g456149/U$1 ( \59788 , \59780 , \59787 );
xor \g456158/U$9 ( \59789 , \59557 , \59565 );
xor \g456158/U$9_r1 ( \59790 , \59789 , \59574 );
and \g456158/U$8 ( \59791 , \59579 , \59790 );
xor \g456158/U$11 ( \59792 , \59557 , \59565 );
xor \g456158/U$11_r1 ( \59793 , \59792 , \59574 );
and \g456158/U$10 ( \59794 , \59626 , \59793 );
and \g456158/U$12 ( \59795 , \59579 , \59626 );
or \g456158/U$7 ( \59796 , \59791 , \59794 , \59795 );
xor \g132508/U$4 ( \59797 , \59688 , \59696 );
and \g132508/U$3 ( \59798 , \59797 , \59701 );
and \g132508/U$5 ( \59799 , \59688 , \59696 );
or \g132508/U$2 ( \59800 , \59798 , \59799 );
not \g132989/U$3 ( \59801 , \49233 );
and \g133013/U$2 ( \59802 , \56167 , \49405 );
and \g133013/U$3 ( \59803 , \49403 , \55884 );
nor \g133013/U$1 ( \59804 , \59802 , \59803 );
not \g132989/U$4 ( \59805 , \59804 );
or \g132989/U$2 ( \59806 , \59801 , \59805 );
or \g132989/U$5 ( \59807 , \59804 , \49233 );
nand \g132989/U$1 ( \59808 , \59806 , \59807 );
xor \g456156/U$2 ( \59809 , \59800 , \59808 );
not \g132905/U$3 ( \59810 , \48483 );
and \g132949/U$2 ( \59811 , \48478 , \56347 );
and \g132949/U$3 ( \59812 , \56349 , \48479 );
nor \g132949/U$1 ( \59813 , \59811 , \59812 );
not \g132905/U$4 ( \59814 , \59813 );
or \g132905/U$2 ( \59815 , \59810 , \59814 );
or \g132905/U$5 ( \59816 , \59813 , \48483 );
nand \g132905/U$1 ( \59817 , \59815 , \59816 );
not \g132980/U$3 ( \59818 , \48685 );
and \g133012/U$2 ( \59819 , \48858 , \56357 );
and \g133012/U$3 ( \59820 , \56359 , \48860 );
nor \g133012/U$1 ( \59821 , \59819 , \59820 );
not \g132980/U$4 ( \59822 , \59821 );
or \g132980/U$2 ( \59823 , \59818 , \59822 );
or \g132980/U$5 ( \59824 , \59821 , \48685 );
nand \g132980/U$1 ( \59825 , \59823 , \59824 );
xor \g132581/U$1 ( \59826 , \59817 , \59825 );
and \g132672/U$2 ( \59827 , \59679 , \59687 );
xor \g132581/U$1_r1 ( \59828 , \59826 , \59827 );
xor \g456156/U$1 ( \59829 , \59809 , \59828 );
not \g132455/U$3 ( \59830 , \50759 );
and \g132501/U$2 ( \59831 , \54185 , \51053 );
and \g132501/U$3 ( \59832 , \51055 , \54251 );
nor \g132501/U$1 ( \59833 , \59831 , \59832 );
not \g132455/U$4 ( \59834 , \59833 );
or \g132455/U$2 ( \59835 , \59830 , \59834 );
or \g132455/U$5 ( \59836 , \59833 , \50759 );
nand \g132455/U$1 ( \59837 , \59835 , \59836 );
not \g132746/U$3 ( \59838 , \49925 );
and \g132787/U$2 ( \59839 , \54853 , \50159 );
and \g132787/U$3 ( \59840 , \50160 , \55127 );
nor \g132787/U$1 ( \59841 , \59839 , \59840 );
not \g132746/U$4 ( \59842 , \59841 );
or \g132746/U$2 ( \59843 , \59838 , \59842 );
or \g132746/U$5 ( \59844 , \59841 , \49925 );
nand \g132746/U$1 ( \59845 , \59843 , \59844 );
not \g132882/U$3 ( \59846 , \49568 );
and \g132911/U$2 ( \59847 , \55460 , \49812 );
and \g132911/U$3 ( \59848 , \49813 , \55707 );
nor \g132911/U$1 ( \59849 , \59847 , \59848 );
not \g132882/U$4 ( \59850 , \59849 );
or \g132882/U$2 ( \59851 , \59846 , \59850 );
or \g132882/U$5 ( \59852 , \59849 , \49568 );
nand \g132882/U$1 ( \59853 , \59851 , \59852 );
xor \g132238/U$1 ( \59854 , \59845 , \59853 );
xor \g132585/U$4 ( \59855 , \59613 , \59621 );
and \g132585/U$3 ( \59856 , \59855 , \59623 );
and \g132585/U$5 ( \59857 , \59613 , \59621 );
or \g132585/U$2 ( \59858 , \59856 , \59857 );
not \g133069/U$3 ( \59859 , \49014 );
and \g133100/U$2 ( \59860 , \56446 , \49074 );
and \g133100/U$3 ( \59861 , \56448 , \49075 );
nor \g133100/U$1 ( \59862 , \59860 , \59861 );
not \g133069/U$4 ( \59863 , \59862 );
or \g133069/U$2 ( \59864 , \59859 , \59863 );
or \g133069/U$5 ( \59865 , \59862 , \49014 );
nand \g133069/U$1 ( \59866 , \59864 , \59865 );
xor \g132358/U$1 ( \59867 , \59858 , \59866 );
not \g132614/U$3 ( \59868 , \47997 );
and \g132638/U$2 ( \59869 , \48064 , \47026 );
and \g132638/U$3 ( \59870 , \56377 , \48063 );
nor \g132638/U$1 ( \59871 , \59869 , \59870 );
not \g132614/U$4 ( \59872 , \59871 );
or \g132614/U$2 ( \59873 , \59868 , \59872 );
or \g132614/U$5 ( \59874 , \59871 , \47997 );
nand \g132614/U$1 ( \59875 , \59873 , \59874 );
not \g132816/U$3 ( \59876 , \48323 );
and \g132859/U$2 ( \59877 , \48334 , \56411 );
and \g132859/U$3 ( \59878 , \56368 , \48335 );
nor \g132859/U$1 ( \59879 , \59877 , \59878 );
not \g132816/U$4 ( \59880 , \59879 );
or \g132816/U$2 ( \59881 , \59876 , \59880 );
or \g132816/U$5 ( \59882 , \59879 , \48323 );
nand \g132816/U$1 ( \59883 , \59881 , \59882 );
xor \g132467/U$1 ( \59884 , \59875 , \59883 );
not \g132714/U$3 ( \59885 , \48159 );
and \g132767/U$2 ( \59886 , \48154 , \56370 );
and \g132767/U$3 ( \59887 , \56379 , \48155 );
nor \g132767/U$1 ( \59888 , \59886 , \59887 );
not \g132714/U$4 ( \59889 , \59888 );
or \g132714/U$2 ( \59890 , \59885 , \59889 );
or \g132714/U$5 ( \59891 , \59888 , \48159 );
nand \g132714/U$1 ( \59892 , \59890 , \59891 );
and \g132636/U$2 ( \59893 , \47997 , \59537 );
xor \g132579/U$1 ( \59894 , \59892 , \59893 );
xor \g132467/U$1_r1 ( \59895 , \59884 , \59894 );
xor \g132358/U$1_r1 ( \59896 , \59867 , \59895 );
xor \g132238/U$1_r1 ( \59897 , \59854 , \59896 );
xor \g456156/U$1_r1 ( \59898 , \59837 , \59897 );
xor \g456156/U$1_r2 ( \59899 , \59829 , \59898 );
xor \g456149/U$1_r1 ( \59900 , \59796 , \59899 );
xor \g456149/U$1_r2 ( \59901 , \59788 , \59900 );
xor \g131806/U$1_r1 ( \59902 , \59767 , \59901 );
xor \g131041/U$1 ( \59903 , \59549 , \59708 );
xor \g131041/U$1_r1 ( \59904 , \59903 , \59723 );
and \g130996/U$2 ( \59905 , \59902 , \59904 );
and \g130916/U$3 ( \59906 , \59734 , \59905 );
and \g130916/U$5 ( \59907 , \59726 , \59733 );
or \g130916/U$2 ( \59908 , \59906 , \59907 );
xor \g456156/U$9 ( \59909 , \59800 , \59808 );
xor \g456156/U$9_r1 ( \59910 , \59909 , \59828 );
and \g456156/U$8 ( \59911 , \59837 , \59910 );
xor \g456156/U$11 ( \59912 , \59800 , \59808 );
xor \g456156/U$11_r1 ( \59913 , \59912 , \59828 );
and \g456156/U$10 ( \59914 , \59897 , \59913 );
and \g456156/U$12 ( \59915 , \59837 , \59897 );
or \g456156/U$7 ( \59916 , \59911 , \59914 , \59915 );
xor \g456154/U$5 ( \59917 , \59742 , \59750 );
and \g456154/U$4 ( \59918 , \59917 , \59755 );
and \g456154/U$6 ( \59919 , \59742 , \59750 );
or \g456154/U$3 ( \59920 , \59918 , \59919 );
xor \g131995/U$1 ( \59921 , \59916 , \59920 );
xor \g132238/U$4 ( \59922 , \59845 , \59853 );
and \g132238/U$3 ( \59923 , \59922 , \59896 );
and \g132238/U$5 ( \59924 , \59845 , \59853 );
or \g132238/U$2 ( \59925 , \59923 , \59924 );
not \g132152/U$3 ( \59926 , \51124 );
and \g132206/U$2 ( \59927 , \53610 , \51517 );
and \g132206/U$3 ( \59928 , \51518 , \53848 );
nor \g132206/U$1 ( \59929 , \59927 , \59928 );
not \g132152/U$4 ( \59930 , \59929 );
or \g132152/U$2 ( \59931 , \59926 , \59930 );
or \g132152/U$5 ( \59932 , \59929 , \51124 );
nand \g132152/U$1 ( \59933 , \59931 , \59932 );
xor \g132097/U$1 ( \59934 , \59925 , \59933 );
xor \g132581/U$4 ( \59935 , \59817 , \59825 );
and \g132581/U$3 ( \59936 , \59935 , \59827 );
and \g132581/U$5 ( \59937 , \59817 , \59825 );
or \g132581/U$2 ( \59938 , \59936 , \59937 );
not \g132683/U$3 ( \59939 , \49925 );
and \g132726/U$2 ( \59940 , \54853 , \50160 );
and \g132726/U$3 ( \59941 , \50159 , \54537 );
nor \g132726/U$1 ( \59942 , \59940 , \59941 );
not \g132683/U$4 ( \59943 , \59942 );
or \g132683/U$2 ( \59944 , \59939 , \59943 );
or \g132683/U$5 ( \59945 , \59942 , \49925 );
nand \g132683/U$1 ( \59946 , \59944 , \59945 );
xor \g132237/U$1 ( \59947 , \59938 , \59946 );
not \g132712/U$3 ( \59948 , \48159 );
and \g132765/U$2 ( \59949 , \48154 , \56368 );
and \g132765/U$3 ( \59950 , \56370 , \48155 );
nor \g132765/U$1 ( \59951 , \59949 , \59950 );
not \g132712/U$4 ( \59952 , \59951 );
or \g132712/U$2 ( \59953 , \59948 , \59952 );
or \g132712/U$5 ( \59954 , \59951 , \48159 );
nand \g132712/U$1 ( \59955 , \59953 , \59954 );
not \g132612/U$3 ( \59956 , \47997 );
and \g132656/U$2 ( \59957 , \48064 , \56377 );
and \g132656/U$3 ( \59958 , \56379 , \48063 );
nor \g132656/U$1 ( \59959 , \59957 , \59958 );
not \g132612/U$4 ( \59960 , \59959 );
or \g132612/U$2 ( \59961 , \59956 , \59960 );
or \g132612/U$5 ( \59962 , \59959 , \47997 );
nand \g132612/U$1 ( \59963 , \59961 , \59962 );
xor \g132562/U$1 ( \59964 , \59955 , \59963 );
not \g132999/U$3 ( \59965 , \48685 );
and \g133016/U$2 ( \59966 , \48860 , \56357 );
and \g133016/U$3 ( \59967 , \56448 , \48858 );
nor \g133016/U$1 ( \59968 , \59966 , \59967 );
not \g132999/U$4 ( \59969 , \59968 );
or \g132999/U$2 ( \59970 , \59965 , \59969 );
or \g132999/U$5 ( \59971 , \59968 , \48685 );
nand \g132999/U$1 ( \59972 , \59970 , \59971 );
xor \g132361/U$1 ( \59973 , \59964 , \59972 );
xor \g132467/U$4 ( \59974 , \59875 , \59883 );
and \g132467/U$3 ( \59975 , \59974 , \59894 );
and \g132467/U$5 ( \59976 , \59875 , \59883 );
or \g132467/U$2 ( \59977 , \59975 , \59976 );
xor \g132361/U$1_r1 ( \59978 , \59973 , \59977 );
xor \g132237/U$1_r1 ( \59979 , \59947 , \59978 );
xor \g132097/U$1_r1 ( \59980 , \59934 , \59979 );
xor \g131995/U$1_r1 ( \59981 , \59921 , \59980 );
xor \g456149/U$9 ( \59982 , \59771 , \59779 );
xor \g456149/U$9_r1 ( \59983 , \59982 , \59787 );
and \g456149/U$8 ( \59984 , \59796 , \59983 );
xor \g456149/U$11 ( \59985 , \59771 , \59779 );
xor \g456149/U$11_r1 ( \59986 , \59985 , \59787 );
and \g456149/U$10 ( \59987 , \59899 , \59986 );
and \g456149/U$12 ( \59988 , \59796 , \59899 );
or \g456149/U$7 ( \59989 , \59984 , \59987 , \59988 );
xor \g456091/U$5 ( \59990 , \59981 , \59989 );
xor \g456154/U$9 ( \59991 , \59742 , \59750 );
xor \g456154/U$9_r1 ( \59992 , \59991 , \59755 );
and \g456154/U$8 ( \59993 , \59760 , \59992 );
xor \g456154/U$11 ( \59994 , \59742 , \59750 );
xor \g456154/U$11_r1 ( \59995 , \59994 , \59755 );
and \g456154/U$10 ( \59996 , \59764 , \59995 );
and \g456154/U$12 ( \59997 , \59760 , \59764 );
or \g456154/U$7 ( \59998 , \59993 , \59996 , \59997 );
xor \g456149/U$5 ( \59999 , \59771 , \59779 );
and \g456149/U$4 ( \60000 , \59999 , \59787 );
and \g456149/U$6 ( \60001 , \59771 , \59779 );
or \g456149/U$3 ( \60002 , \60000 , \60001 );
xor \g131838/U$1 ( \60003 , \59998 , \60002 );
and \g132054/U$2 ( \60004 , \52978 , \52270 );
and \g132054/U$3 ( \60005 , \52273 , \53300 );
nor \g132054/U$1 ( \60006 , \60004 , \60005 );
and \g132010/U$2 ( \60007 , \60006 , \51513 );
not \g132010/U$4 ( \60008 , \60006 );
and \g132010/U$3 ( \60009 , \60008 , \51120 );
nor \g132010/U$1 ( \60010 , \60007 , \60009 );
not \g132345/U$3 ( \60011 , \50759 );
and \g132430/U$2 ( \60012 , \54185 , \51055 );
and \g132430/U$3 ( \60013 , \51053 , \54015 );
nor \g132430/U$1 ( \60014 , \60012 , \60013 );
not \g132345/U$4 ( \60015 , \60014 );
or \g132345/U$2 ( \60016 , \60011 , \60015 );
or \g132345/U$5 ( \60017 , \60014 , \50759 );
nand \g132345/U$1 ( \60018 , \60016 , \60017 );
not \g132532/U$3 ( \60019 , \50362 );
and \g132572/U$2 ( \60020 , \54251 , \50587 );
and \g132572/U$3 ( \60021 , \50588 , \54529 );
nor \g132572/U$1 ( \60022 , \60020 , \60021 );
not \g132532/U$4 ( \60023 , \60022 );
or \g132532/U$2 ( \60024 , \60019 , \60023 );
or \g132532/U$5 ( \60025 , \60022 , \50362 );
nand \g132532/U$1 ( \60026 , \60024 , \60025 );
xor \g132258/U$1 ( \60027 , \60018 , \60026 );
xor \g456156/U$5 ( \60028 , \59800 , \59808 );
and \g456156/U$4 ( \60029 , \60028 , \59828 );
and \g456156/U$6 ( \60030 , \59800 , \59808 );
or \g456156/U$3 ( \60031 , \60029 , \60030 );
xor \g132258/U$1_r1 ( \60032 , \60027 , \60031 );
xor \g131935/U$1 ( \60033 , \60010 , \60032 );
xor \g132358/U$4 ( \60034 , \59858 , \59866 );
and \g132358/U$3 ( \60035 , \60034 , \59895 );
and \g132358/U$5 ( \60036 , \59858 , \59866 );
or \g132358/U$2 ( \60037 , \60035 , \60036 );
not \g132822/U$3 ( \60038 , \49568 );
and \g132856/U$2 ( \60039 , \55127 , \49812 );
and \g132856/U$3 ( \60040 , \49813 , \55460 );
nor \g132856/U$1 ( \60041 , \60039 , \60040 );
not \g132822/U$4 ( \60042 , \60041 );
or \g132822/U$2 ( \60043 , \60038 , \60042 );
or \g132822/U$5 ( \60044 , \60041 , \49568 );
nand \g132822/U$1 ( \60045 , \60043 , \60044 );
xor \g132239/U$1 ( \60046 , \60037 , \60045 );
not \g132930/U$3 ( \60047 , \49233 );
and \g132964/U$2 ( \60048 , \55884 , \49405 );
and \g132964/U$3 ( \60049 , \49403 , \55707 );
nor \g132964/U$1 ( \60050 , \60048 , \60049 );
not \g132930/U$4 ( \60051 , \60050 );
or \g132930/U$2 ( \60052 , \60047 , \60051 );
or \g132930/U$5 ( \60053 , \60050 , \49233 );
nand \g132930/U$1 ( \60054 , \60052 , \60053 );
not \g133040/U$3 ( \60055 , \49014 );
and \g133072/U$2 ( \60056 , \49075 , \56446 );
and \g133072/U$3 ( \60057 , \49074 , \56167 );
nor \g133072/U$1 ( \60058 , \60056 , \60057 );
not \g133040/U$4 ( \60059 , \60058 );
or \g133040/U$2 ( \60060 , \60055 , \60059 );
or \g133040/U$5 ( \60061 , \60058 , \49014 );
nand \g133040/U$1 ( \60062 , \60060 , \60061 );
xor \g132359/U$1 ( \60063 , \60054 , \60062 );
not \g132815/U$3 ( \60064 , \48323 );
and \g132838/U$2 ( \60065 , \48334 , \56349 );
and \g132838/U$3 ( \60066 , \56411 , \48335 );
nor \g132838/U$1 ( \60067 , \60065 , \60066 );
not \g132815/U$4 ( \60068 , \60067 );
or \g132815/U$2 ( \60069 , \60064 , \60068 );
or \g132815/U$5 ( \60070 , \60067 , \48323 );
nand \g132815/U$1 ( \60071 , \60069 , \60070 );
not \g132899/U$3 ( \60072 , \48483 );
and \g132944/U$2 ( \60073 , \48479 , \56347 );
and \g132944/U$3 ( \60074 , \56359 , \48478 );
nor \g132944/U$1 ( \60075 , \60073 , \60074 );
not \g132899/U$4 ( \60076 , \60075 );
or \g132899/U$2 ( \60077 , \60072 , \60076 );
or \g132899/U$5 ( \60078 , \60075 , \48483 );
nand \g132899/U$1 ( \60079 , \60077 , \60078 );
xor \g132466/U$1 ( \60080 , \60071 , \60079 );
and \g132579/U$2 ( \60081 , \59892 , \59893 );
xor \g132466/U$1_r1 ( \60082 , \60080 , \60081 );
xor \g132359/U$1_r1 ( \60083 , \60063 , \60082 );
xor \g132239/U$1_r1 ( \60084 , \60046 , \60083 );
xor \g131935/U$1_r1 ( \60085 , \60033 , \60084 );
xor \g131838/U$1_r1 ( \60086 , \60003 , \60085 );
and \g456091/U$4 ( \60087 , \59990 , \60086 );
and \g456091/U$6 ( \60088 , \59981 , \59989 );
or \g456091/U$3 ( \60089 , \60087 , \60088 );
xor \g130779/U$4 ( \60090 , \59908 , \60089 );
xor \g131806/U$4 ( \60091 , \59738 , \59766 );
and \g131806/U$3 ( \60092 , \60091 , \59901 );
and \g131806/U$5 ( \60093 , \59738 , \59766 );
or \g131806/U$2 ( \60094 , \60092 , \60093 );
xor \g456091/U$9 ( \60095 , \59981 , \59989 );
xor \g456091/U$9_r1 ( \60096 , \60095 , \60086 );
and \g456091/U$8 ( \60097 , \60094 , \60096 );
xor \g130916/U$1 ( \60098 , \59726 , \59733 );
xor \g130916/U$1_r1 ( \60099 , \60098 , \59905 );
xor \g456091/U$11 ( \60100 , \59981 , \59989 );
xor \g456091/U$11_r1 ( \60101 , \60100 , \60086 );
and \g456091/U$10 ( \60102 , \60099 , \60101 );
and \g456091/U$12 ( \60103 , \60094 , \60099 );
or \g456091/U$7 ( \60104 , \60097 , \60102 , \60103 );
and \g130779/U$3 ( \60105 , \60090 , \60104 );
and \g130779/U$5 ( \60106 , \59908 , \60089 );
or \g130779/U$2 ( \60107 , \60105 , \60106 );
xor \g132390/U$1 ( \60108 , \47976 , \56439 );
xor \g130668/U$4 ( \60109 , \60107 , \60108 );
not \g132086/U$3 ( \60110 , \51124 );
and \g132133/U$2 ( \60111 , \53610 , \51518 );
and \g132133/U$3 ( \60112 , \51517 , \53300 );
nor \g132133/U$1 ( \60113 , \60111 , \60112 );
not \g132086/U$4 ( \60114 , \60113 );
or \g132086/U$2 ( \60115 , \60110 , \60114 );
or \g132086/U$5 ( \60116 , \60113 , \51124 );
nand \g132086/U$1 ( \60117 , \60115 , \60116 );
not \g132252/U$3 ( \60118 , \50759 );
and \g132297/U$2 ( \60119 , \53848 , \51053 );
and \g132297/U$3 ( \60120 , \51055 , \54015 );
nor \g132297/U$1 ( \60121 , \60119 , \60120 );
not \g132252/U$4 ( \60122 , \60121 );
or \g132252/U$2 ( \60123 , \60118 , \60122 );
or \g132252/U$5 ( \60124 , \60121 , \50759 );
nand \g132252/U$1 ( \60125 , \60123 , \60124 );
xor \g131876/U$1 ( \60126 , \60117 , \60125 );
and \g131968/U$2 ( \60127 , \52978 , \52273 );
and \g131968/U$3 ( \60128 , \52270 , \52883 );
nor \g131968/U$1 ( \60129 , \60127 , \60128 );
and \g131926/U$2 ( \60130 , \60129 , \51513 );
not \g131926/U$4 ( \60131 , \60129 );
and \g131926/U$3 ( \60132 , \60131 , \51120 );
nor \g131926/U$1 ( \60133 , \60130 , \60132 );
xor \g131876/U$1_r1 ( \60134 , \60126 , \60133 );
xor \g132097/U$4 ( \60135 , \59925 , \59933 );
and \g132097/U$3 ( \60136 , \60135 , \59979 );
and \g132097/U$5 ( \60137 , \59925 , \59933 );
or \g132097/U$2 ( \60138 , \60136 , \60137 );
xor \g456140/U$2 ( \60139 , \60134 , \60138 );
xor \g132361/U$4 ( \60140 , \59964 , \59972 );
and \g132361/U$3 ( \60141 , \60140 , \59977 );
and \g132361/U$5 ( \60142 , \59964 , \59972 );
or \g132361/U$2 ( \60143 , \60141 , \60142 );
not \g132984/U$3 ( \60144 , \49014 );
and \g133015/U$2 ( \60145 , \49075 , \56167 );
and \g133015/U$3 ( \60146 , \49074 , \55884 );
nor \g133015/U$1 ( \60147 , \60145 , \60146 );
not \g132984/U$4 ( \60148 , \60147 );
or \g132984/U$2 ( \60149 , \60144 , \60148 );
or \g132984/U$5 ( \60150 , \60147 , \49014 );
nand \g132984/U$1 ( \60151 , \60149 , \60150 );
xor \g456155/U$2 ( \60152 , \60143 , \60151 );
not \g132810/U$3 ( \60153 , \48323 );
and \g132847/U$2 ( \60154 , \48334 , \56347 );
and \g132847/U$3 ( \60155 , \56349 , \48335 );
nor \g132847/U$1 ( \60156 , \60154 , \60155 );
not \g132810/U$4 ( \60157 , \60156 );
or \g132810/U$2 ( \60158 , \60153 , \60157 );
or \g132810/U$5 ( \60159 , \60156 , \48323 );
nand \g132810/U$1 ( \60160 , \60158 , \60159 );
not \g132896/U$3 ( \60161 , \48483 );
and \g132941/U$2 ( \60162 , \48478 , \56357 );
and \g132941/U$3 ( \60163 , \56359 , \48479 );
nor \g132941/U$1 ( \60164 , \60162 , \60163 );
not \g132896/U$4 ( \60165 , \60164 );
or \g132896/U$2 ( \60166 , \60161 , \60165 );
or \g132896/U$5 ( \60167 , \60164 , \48483 );
nand \g132896/U$1 ( \60168 , \60166 , \60167 );
xor \g132460/U$1 ( \60169 , \60160 , \60168 );
and \g132562/U$2 ( \60170 , \59955 , \59963 );
xor \g132460/U$1_r1 ( \60171 , \60169 , \60170 );
xor \g456155/U$1 ( \60172 , \60152 , \60171 );
xor \g132237/U$4 ( \60173 , \59938 , \59946 );
and \g132237/U$3 ( \60174 , \60173 , \59978 );
and \g132237/U$5 ( \60175 , \59938 , \59946 );
or \g132237/U$2 ( \60176 , \60174 , \60175 );
not \g132744/U$3 ( \60177 , \49568 );
and \g132784/U$2 ( \60178 , \54853 , \49812 );
and \g132784/U$3 ( \60179 , \49813 , \55127 );
nor \g132784/U$1 ( \60180 , \60178 , \60179 );
not \g132744/U$4 ( \60181 , \60180 );
or \g132744/U$2 ( \60182 , \60177 , \60181 );
or \g132744/U$5 ( \60183 , \60180 , \49568 );
nand \g132744/U$1 ( \60184 , \60182 , \60183 );
not \g132875/U$3 ( \60185 , \49233 );
and \g132910/U$2 ( \60186 , \55460 , \49403 );
and \g132910/U$3 ( \60187 , \49405 , \55707 );
nor \g132910/U$1 ( \60188 , \60186 , \60187 );
not \g132875/U$4 ( \60189 , \60188 );
or \g132875/U$2 ( \60190 , \60185 , \60189 );
or \g132875/U$5 ( \60191 , \60188 , \49233 );
nand \g132875/U$1 ( \60192 , \60190 , \60191 );
xor \g132107/U$1 ( \60193 , \60184 , \60192 );
xor \g132466/U$4 ( \60194 , \60071 , \60079 );
and \g132466/U$3 ( \60195 , \60194 , \60081 );
and \g132466/U$5 ( \60196 , \60071 , \60079 );
or \g132466/U$2 ( \60197 , \60195 , \60196 );
not \g132983/U$3 ( \60198 , \48685 );
and \g133014/U$2 ( \60199 , \48858 , \56446 );
and \g133014/U$3 ( \60200 , \56448 , \48860 );
nor \g133014/U$1 ( \60201 , \60199 , \60200 );
not \g132983/U$4 ( \60202 , \60201 );
or \g132983/U$2 ( \60203 , \60198 , \60202 );
or \g132983/U$5 ( \60204 , \60201 , \48685 );
nand \g132983/U$1 ( \60205 , \60203 , \60204 );
xor \g132211/U$1 ( \60206 , \60197 , \60205 );
not \g132488/U$3 ( \60207 , \47935 );
and \g132536/U$2 ( \60208 , \47931 , \47026 );
and \g132536/U$3 ( \60209 , \56377 , \47930 );
nor \g132536/U$1 ( \60210 , \60208 , \60209 );
not \g132488/U$4 ( \60211 , \60210 );
or \g132488/U$2 ( \60212 , \60207 , \60211 );
or \g132488/U$5 ( \60213 , \60210 , \47935 );
nand \g132488/U$1 ( \60214 , \60212 , \60213 );
not \g132718/U$3 ( \60215 , \48159 );
and \g132762/U$2 ( \60216 , \48154 , \56411 );
and \g132762/U$3 ( \60217 , \56368 , \48155 );
nor \g132762/U$1 ( \60218 , \60216 , \60217 );
not \g132718/U$4 ( \60219 , \60218 );
or \g132718/U$2 ( \60220 , \60215 , \60219 );
or \g132718/U$5 ( \60221 , \60218 , \48159 );
nand \g132718/U$1 ( \60222 , \60220 , \60221 );
xor \g132316/U$1 ( \60223 , \60214 , \60222 );
not \g132613/U$3 ( \60224 , \47997 );
and \g132657/U$2 ( \60225 , \48063 , \56370 );
and \g132657/U$3 ( \60226 , \56379 , \48064 );
nor \g132657/U$1 ( \60227 , \60225 , \60226 );
not \g132613/U$4 ( \60228 , \60227 );
or \g132613/U$2 ( \60229 , \60224 , \60228 );
or \g132613/U$5 ( \60230 , \60227 , \47997 );
nand \g132613/U$1 ( \60231 , \60229 , \60230 );
and \g132514/U$2 ( \60232 , \47935 , \59732 );
xor \g132462/U$1 ( \60233 , \60231 , \60232 );
xor \g132316/U$1_r1 ( \60234 , \60223 , \60233 );
xor \g132211/U$1_r1 ( \60235 , \60206 , \60234 );
xor \g132107/U$1_r1 ( \60236 , \60193 , \60235 );
xor \g456155/U$1_r1 ( \60237 , \60176 , \60236 );
xor \g456155/U$1_r2 ( \60238 , \60172 , \60237 );
xor \g456140/U$1 ( \60239 , \60139 , \60238 );
xor \g131838/U$4 ( \60240 , \59998 , \60002 );
and \g131838/U$3 ( \60241 , \60240 , \60085 );
and \g131838/U$5 ( \60242 , \59998 , \60002 );
or \g131838/U$2 ( \60243 , \60241 , \60242 );
xor \g132239/U$4 ( \60244 , \60037 , \60045 );
and \g132239/U$3 ( \60245 , \60244 , \60083 );
and \g132239/U$5 ( \60246 , \60037 , \60045 );
or \g132239/U$2 ( \60247 , \60245 , \60246 );
xor \g132258/U$4 ( \60248 , \60018 , \60026 );
and \g132258/U$3 ( \60249 , \60248 , \60031 );
and \g132258/U$5 ( \60250 , \60018 , \60026 );
or \g132258/U$2 ( \60251 , \60249 , \60250 );
xor \g456148/U$2 ( \60252 , \60247 , \60251 );
not \g132454/U$3 ( \60253 , \50362 );
and \g132499/U$2 ( \60254 , \54185 , \50587 );
and \g132499/U$3 ( \60255 , \50588 , \54251 );
nor \g132499/U$1 ( \60256 , \60254 , \60255 );
not \g132454/U$4 ( \60257 , \60256 );
or \g132454/U$2 ( \60258 , \60253 , \60257 );
or \g132454/U$5 ( \60259 , \60256 , \50362 );
nand \g132454/U$1 ( \60260 , \60258 , \60259 );
not \g132621/U$3 ( \60261 , \49925 );
and \g132661/U$2 ( \60262 , \54537 , \50160 );
and \g132661/U$3 ( \60263 , \50159 , \54529 );
nor \g132661/U$1 ( \60264 , \60262 , \60263 );
not \g132621/U$4 ( \60265 , \60264 );
or \g132621/U$2 ( \60266 , \60261 , \60265 );
or \g132621/U$5 ( \60267 , \60264 , \49925 );
nand \g132621/U$1 ( \60268 , \60266 , \60267 );
xor \g132240/U$1 ( \60269 , \60260 , \60268 );
xor \g132359/U$4 ( \60270 , \60054 , \60062 );
and \g132359/U$3 ( \60271 , \60270 , \60082 );
and \g132359/U$5 ( \60272 , \60054 , \60062 );
or \g132359/U$2 ( \60273 , \60271 , \60272 );
xor \g132240/U$1_r1 ( \60274 , \60269 , \60273 );
xor \g456148/U$1 ( \60275 , \60252 , \60274 );
xor \g131935/U$4 ( \60276 , \60010 , \60032 );
and \g131935/U$3 ( \60277 , \60276 , \60084 );
and \g131935/U$5 ( \60278 , \60010 , \60032 );
or \g131935/U$2 ( \60279 , \60277 , \60278 );
xor \g131995/U$4 ( \60280 , \59916 , \59920 );
and \g131995/U$3 ( \60281 , \60280 , \59980 );
and \g131995/U$5 ( \60282 , \59916 , \59920 );
or \g131995/U$2 ( \60283 , \60281 , \60282 );
xor \g456148/U$1_r1 ( \60284 , \60279 , \60283 );
xor \g456148/U$1_r2 ( \60285 , \60275 , \60284 );
xor \g456140/U$1_r1 ( \60286 , \60243 , \60285 );
xor \g456140/U$1_r2 ( \60287 , \60239 , \60286 );
xor \g130779/U$1 ( \60288 , \59908 , \60089 );
xor \g130779/U$1_r1 ( \60289 , \60288 , \60104 );
and \g130744/U$2 ( \60290 , \60287 , \60289 );
and \g130668/U$3 ( \60291 , \60109 , \60290 );
and \g130668/U$5 ( \60292 , \60107 , \60108 );
or \g130668/U$2 ( \60293 , \60291 , \60292 );
xor \g131876/U$4 ( \60294 , \60117 , \60125 );
and \g131876/U$3 ( \60295 , \60294 , \60133 );
and \g131876/U$5 ( \60296 , \60117 , \60125 );
or \g131876/U$2 ( \60297 , \60295 , \60296 );
xor \g456148/U$5 ( \60298 , \60247 , \60251 );
and \g456148/U$4 ( \60299 , \60298 , \60274 );
and \g456148/U$6 ( \60300 , \60247 , \60251 );
or \g456148/U$3 ( \60301 , \60299 , \60300 );
xor \g131807/U$1 ( \60302 , \60297 , \60301 );
xor \g132107/U$4 ( \60303 , \60184 , \60192 );
and \g132107/U$3 ( \60304 , \60303 , \60235 );
and \g132107/U$5 ( \60305 , \60184 , \60192 );
or \g132107/U$2 ( \60306 , \60304 , \60305 );
not \g132007/U$3 ( \60307 , \51124 );
and \g132053/U$2 ( \60308 , \52978 , \51517 );
and \g132053/U$3 ( \60309 , \51518 , \53300 );
nor \g132053/U$1 ( \60310 , \60308 , \60309 );
not \g132007/U$4 ( \60311 , \60310 );
or \g132007/U$2 ( \60312 , \60307 , \60311 );
or \g132007/U$5 ( \60313 , \60310 , \51124 );
nand \g132007/U$1 ( \60314 , \60312 , \60313 );
xor \g131934/U$1 ( \60315 , \60306 , \60314 );
not \g132681/U$3 ( \60316 , \49568 );
and \g132725/U$2 ( \60317 , \54853 , \49813 );
and \g132725/U$3 ( \60318 , \49812 , \54537 );
nor \g132725/U$1 ( \60319 , \60317 , \60318 );
not \g132681/U$4 ( \60320 , \60319 );
or \g132681/U$2 ( \60321 , \60316 , \60320 );
or \g132681/U$5 ( \60322 , \60319 , \49568 );
nand \g132681/U$1 ( \60323 , \60321 , \60322 );
not \g132928/U$3 ( \60324 , \49014 );
and \g132962/U$2 ( \60325 , \55884 , \49075 );
and \g132962/U$3 ( \60326 , \49074 , \55707 );
nor \g132962/U$1 ( \60327 , \60325 , \60326 );
not \g132928/U$4 ( \60328 , \60327 );
or \g132928/U$2 ( \60329 , \60324 , \60328 );
or \g132928/U$5 ( \60330 , \60327 , \49014 );
nand \g132928/U$1 ( \60331 , \60329 , \60330 );
xor \g132105/U$1 ( \60332 , \60323 , \60331 );
not \g132609/U$3 ( \60333 , \47997 );
and \g132659/U$2 ( \60334 , \48063 , \56368 );
and \g132659/U$3 ( \60335 , \56370 , \48064 );
nor \g132659/U$1 ( \60336 , \60334 , \60335 );
not \g132609/U$4 ( \60337 , \60336 );
or \g132609/U$2 ( \60338 , \60333 , \60337 );
or \g132609/U$5 ( \60339 , \60336 , \47997 );
nand \g132609/U$1 ( \60340 , \60338 , \60339 );
not \g132487/U$3 ( \60341 , \47935 );
and \g132549/U$2 ( \60342 , \47931 , \56377 );
and \g132549/U$3 ( \60343 , \56379 , \47930 );
nor \g132549/U$1 ( \60344 , \60342 , \60343 );
not \g132487/U$4 ( \60345 , \60344 );
or \g132487/U$2 ( \60346 , \60341 , \60345 );
or \g132487/U$5 ( \60347 , \60344 , \47935 );
nand \g132487/U$1 ( \60348 , \60346 , \60347 );
xor \g132441/U$1 ( \60349 , \60340 , \60348 );
not \g132897/U$3 ( \60350 , \48483 );
and \g132951/U$2 ( \60351 , \48479 , \56357 );
and \g132951/U$3 ( \60352 , \56448 , \48478 );
nor \g132951/U$1 ( \60353 , \60351 , \60352 );
not \g132897/U$4 ( \60354 , \60353 );
or \g132897/U$2 ( \60355 , \60350 , \60354 );
or \g132897/U$5 ( \60356 , \60353 , \48483 );
nand \g132897/U$1 ( \60357 , \60355 , \60356 );
xor \g132209/U$1 ( \60358 , \60349 , \60357 );
xor \g132316/U$4 ( \60359 , \60214 , \60222 );
and \g132316/U$3 ( \60360 , \60359 , \60233 );
and \g132316/U$5 ( \60361 , \60214 , \60222 );
or \g132316/U$2 ( \60362 , \60360 , \60361 );
xor \g132209/U$1_r1 ( \60363 , \60358 , \60362 );
xor \g132105/U$1_r1 ( \60364 , \60332 , \60363 );
xor \g131934/U$1_r1 ( \60365 , \60315 , \60364 );
xor \g131807/U$1_r1 ( \60366 , \60302 , \60365 );
xor \g456148/U$9 ( \60367 , \60247 , \60251 );
xor \g456148/U$9_r1 ( \60368 , \60367 , \60274 );
and \g456148/U$8 ( \60369 , \60279 , \60368 );
xor \g456148/U$11 ( \60370 , \60247 , \60251 );
xor \g456148/U$11_r1 ( \60371 , \60370 , \60274 );
and \g456148/U$10 ( \60372 , \60283 , \60371 );
and \g456148/U$12 ( \60373 , \60279 , \60283 );
or \g456148/U$7 ( \60374 , \60369 , \60372 , \60373 );
xor \g456077/U$5 ( \60375 , \60366 , \60374 );
xor \g456140/U$5 ( \60376 , \60134 , \60138 );
and \g456140/U$4 ( \60377 , \60376 , \60238 );
and \g456140/U$6 ( \60378 , \60134 , \60138 );
or \g456140/U$3 ( \60379 , \60377 , \60378 );
and \g131902/U$2 ( \60380 , \52620 , \52270 );
and \g131902/U$3 ( \60381 , \52273 , \52883 );
nor \g131902/U$1 ( \60382 , \60380 , \60381 );
and \g131853/U$2 ( \60383 , \60382 , \51513 );
not \g131853/U$4 ( \60384 , \60382 );
and \g131853/U$3 ( \60385 , \60384 , \51120 );
nor \g131853/U$1 ( \60386 , \60383 , \60385 );
not \g132153/U$3 ( \60387 , \50759 );
and \g132195/U$2 ( \60388 , \53610 , \51053 );
and \g132195/U$3 ( \60389 , \51055 , \53848 );
nor \g132195/U$1 ( \60390 , \60388 , \60389 );
not \g132153/U$4 ( \60391 , \60390 );
or \g132153/U$2 ( \60392 , \60387 , \60391 );
or \g132153/U$5 ( \60393 , \60390 , \50759 );
nand \g132153/U$1 ( \60394 , \60392 , \60393 );
xor \g131802/U$1 ( \60395 , \60386 , \60394 );
xor \g132211/U$4 ( \60396 , \60197 , \60205 );
and \g132211/U$3 ( \60397 , \60396 , \60234 );
and \g132211/U$5 ( \60398 , \60197 , \60205 );
or \g132211/U$2 ( \60399 , \60397 , \60398 );
not \g132814/U$3 ( \60400 , \49233 );
and \g132850/U$2 ( \60401 , \55127 , \49403 );
and \g132850/U$3 ( \60402 , \49405 , \55460 );
nor \g132850/U$1 ( \60403 , \60401 , \60402 );
not \g132814/U$4 ( \60404 , \60403 );
or \g132814/U$2 ( \60405 , \60400 , \60404 );
or \g132814/U$5 ( \60406 , \60403 , \49233 );
nand \g132814/U$1 ( \60407 , \60405 , \60406 );
xor \g132106/U$1 ( \60408 , \60399 , \60407 );
xor \g132460/U$4 ( \60409 , \60160 , \60168 );
and \g132460/U$3 ( \60410 , \60409 , \60170 );
and \g132460/U$5 ( \60411 , \60160 , \60168 );
or \g132460/U$2 ( \60412 , \60410 , \60411 );
not \g132981/U$3 ( \60413 , \48685 );
and \g133010/U$2 ( \60414 , \48860 , \56446 );
and \g133010/U$3 ( \60415 , \56167 , \48858 );
nor \g133010/U$1 ( \60416 , \60414 , \60415 );
not \g132981/U$4 ( \60417 , \60416 );
or \g132981/U$2 ( \60418 , \60413 , \60417 );
or \g132981/U$5 ( \60419 , \60416 , \48685 );
nand \g132981/U$1 ( \60420 , \60418 , \60419 );
xor \g132208/U$1 ( \60421 , \60412 , \60420 );
not \g132713/U$3 ( \60422 , \48159 );
and \g132764/U$2 ( \60423 , \48154 , \56349 );
and \g132764/U$3 ( \60424 , \56411 , \48155 );
nor \g132764/U$1 ( \60425 , \60423 , \60424 );
not \g132713/U$4 ( \60426 , \60425 );
or \g132713/U$2 ( \60427 , \60422 , \60426 );
or \g132713/U$5 ( \60428 , \60425 , \48159 );
nand \g132713/U$1 ( \60429 , \60427 , \60428 );
not \g132811/U$3 ( \60430 , \48323 );
and \g132848/U$2 ( \60431 , \48335 , \56347 );
and \g132848/U$3 ( \60432 , \56359 , \48334 );
nor \g132848/U$1 ( \60433 , \60431 , \60432 );
not \g132811/U$4 ( \60434 , \60433 );
or \g132811/U$2 ( \60435 , \60430 , \60434 );
or \g132811/U$5 ( \60436 , \60433 , \48323 );
nand \g132811/U$1 ( \60437 , \60435 , \60436 );
xor \g132317/U$1 ( \60438 , \60429 , \60437 );
and \g132462/U$2 ( \60439 , \60231 , \60232 );
xor \g132317/U$1_r1 ( \60440 , \60438 , \60439 );
xor \g132208/U$1_r1 ( \60441 , \60421 , \60440 );
xor \g132106/U$1_r1 ( \60442 , \60408 , \60441 );
xor \g131802/U$1_r1 ( \60443 , \60395 , \60442 );
xor \g131702/U$1 ( \60444 , \60379 , \60443 );
not \g132343/U$3 ( \60445 , \50362 );
and \g132425/U$2 ( \60446 , \54185 , \50588 );
and \g132425/U$3 ( \60447 , \50587 , \54015 );
nor \g132425/U$1 ( \60448 , \60446 , \60447 );
not \g132343/U$4 ( \60449 , \60448 );
or \g132343/U$2 ( \60450 , \60445 , \60449 );
or \g132343/U$5 ( \60451 , \60448 , \50362 );
nand \g132343/U$1 ( \60452 , \60450 , \60451 );
not \g132530/U$3 ( \60453 , \49925 );
and \g132571/U$2 ( \60454 , \54251 , \50159 );
and \g132571/U$3 ( \60455 , \50160 , \54529 );
nor \g132571/U$1 ( \60456 , \60454 , \60455 );
not \g132530/U$4 ( \60457 , \60456 );
or \g132530/U$2 ( \60458 , \60453 , \60457 );
or \g132530/U$5 ( \60459 , \60456 , \49925 );
nand \g132530/U$1 ( \60460 , \60458 , \60459 );
xor \g456152/U$2 ( \60461 , \60452 , \60460 );
xor \g456155/U$5 ( \60462 , \60143 , \60151 );
and \g456155/U$4 ( \60463 , \60462 , \60171 );
and \g456155/U$6 ( \60464 , \60143 , \60151 );
or \g456155/U$3 ( \60465 , \60463 , \60464 );
xor \g456152/U$1 ( \60466 , \60461 , \60465 );
xor \g132240/U$4 ( \60467 , \60260 , \60268 );
and \g132240/U$3 ( \60468 , \60467 , \60273 );
and \g132240/U$5 ( \60469 , \60260 , \60268 );
or \g132240/U$2 ( \60470 , \60468 , \60469 );
xor \g456155/U$9 ( \60471 , \60143 , \60151 );
xor \g456155/U$9_r1 ( \60472 , \60471 , \60171 );
and \g456155/U$8 ( \60473 , \60176 , \60472 );
xor \g456155/U$11 ( \60474 , \60143 , \60151 );
xor \g456155/U$11_r1 ( \60475 , \60474 , \60171 );
and \g456155/U$10 ( \60476 , \60236 , \60475 );
and \g456155/U$12 ( \60477 , \60176 , \60236 );
or \g456155/U$7 ( \60478 , \60473 , \60476 , \60477 );
xor \g456152/U$1_r1 ( \60479 , \60470 , \60478 );
xor \g456152/U$1_r2 ( \60480 , \60466 , \60479 );
xor \g131702/U$1_r1 ( \60481 , \60444 , \60480 );
and \g456077/U$4 ( \60482 , \60375 , \60481 );
and \g456077/U$6 ( \60483 , \60366 , \60374 );
or \g456077/U$3 ( \60484 , \60482 , \60483 );
xor \g130499/U$4 ( \60485 , \60293 , \60484 );
xor \g456140/U$9 ( \60486 , \60134 , \60138 );
xor \g456140/U$9_r1 ( \60487 , \60486 , \60238 );
and \g456140/U$8 ( \60488 , \60243 , \60487 );
xor \g456140/U$11 ( \60489 , \60134 , \60138 );
xor \g456140/U$11_r1 ( \60490 , \60489 , \60238 );
and \g456140/U$10 ( \60491 , \60285 , \60490 );
and \g456140/U$12 ( \60492 , \60243 , \60285 );
or \g456140/U$7 ( \60493 , \60488 , \60491 , \60492 );
xor \g456077/U$9 ( \60494 , \60366 , \60374 );
xor \g456077/U$9_r1 ( \60495 , \60494 , \60481 );
and \g456077/U$8 ( \60496 , \60493 , \60495 );
xor \g130668/U$1 ( \60497 , \60107 , \60108 );
xor \g130668/U$1_r1 ( \60498 , \60497 , \60290 );
xor \g456077/U$11 ( \60499 , \60366 , \60374 );
xor \g456077/U$11_r1 ( \60500 , \60499 , \60481 );
and \g456077/U$10 ( \60501 , \60498 , \60500 );
and \g456077/U$12 ( \60502 , \60493 , \60498 );
or \g456077/U$7 ( \60503 , \60496 , \60501 , \60502 );
and \g130499/U$3 ( \60504 , \60485 , \60503 );
and \g130499/U$5 ( \60505 , \60293 , \60484 );
or \g130499/U$2 ( \60506 , \60504 , \60505 );
xor \g132242/U$1 ( \60507 , \47948 , \56485 );
xor \g130356/U$4 ( \60508 , \60506 , \60507 );
xor \g131807/U$4 ( \60509 , \60297 , \60301 );
and \g131807/U$3 ( \60510 , \60509 , \60365 );
and \g131807/U$5 ( \60511 , \60297 , \60301 );
or \g131807/U$2 ( \60512 , \60510 , \60511 );
xor \g456152/U$9 ( \60513 , \60452 , \60460 );
xor \g456152/U$9_r1 ( \60514 , \60513 , \60465 );
and \g456152/U$8 ( \60515 , \60470 , \60514 );
xor \g456152/U$11 ( \60516 , \60452 , \60460 );
xor \g456152/U$11_r1 ( \60517 , \60516 , \60465 );
and \g456152/U$10 ( \60518 , \60478 , \60517 );
and \g456152/U$12 ( \60519 , \60470 , \60478 );
or \g456152/U$7 ( \60520 , \60515 , \60518 , \60519 );
xor \g456132/U$2 ( \60521 , \60512 , \60520 );
not \g132084/U$3 ( \60522 , \50759 );
and \g132125/U$2 ( \60523 , \53610 , \51055 );
and \g132125/U$3 ( \60524 , \51053 , \53300 );
nor \g132125/U$1 ( \60525 , \60523 , \60524 );
not \g132084/U$4 ( \60526 , \60525 );
or \g132084/U$2 ( \60527 , \60522 , \60526 );
or \g132084/U$5 ( \60528 , \60525 , \50759 );
nand \g132084/U$1 ( \60529 , \60527 , \60528 );
not \g132452/U$3 ( \60530 , \49925 );
and \g132498/U$2 ( \60531 , \54185 , \50159 );
and \g132498/U$3 ( \60532 , \50160 , \54251 );
nor \g132498/U$1 ( \60533 , \60531 , \60532 );
not \g132452/U$4 ( \60534 , \60533 );
or \g132452/U$2 ( \60535 , \60530 , \60534 );
or \g132452/U$5 ( \60536 , \60533 , \49925 );
nand \g132452/U$1 ( \60537 , \60535 , \60536 );
xor \g456147/U$2 ( \60538 , \60529 , \60537 );
xor \g132105/U$4 ( \60539 , \60323 , \60331 );
and \g132105/U$3 ( \60540 , \60539 , \60363 );
and \g132105/U$5 ( \60541 , \60323 , \60331 );
or \g132105/U$2 ( \60542 , \60540 , \60541 );
xor \g456147/U$1 ( \60543 , \60538 , \60542 );
xor \g456152/U$5 ( \60544 , \60452 , \60460 );
and \g456152/U$4 ( \60545 , \60544 , \60465 );
and \g456152/U$6 ( \60546 , \60452 , \60460 );
or \g456152/U$3 ( \60547 , \60545 , \60546 );
xor \g131934/U$4 ( \60548 , \60306 , \60314 );
and \g131934/U$3 ( \60549 , \60548 , \60364 );
and \g131934/U$5 ( \60550 , \60306 , \60314 );
or \g131934/U$2 ( \60551 , \60549 , \60550 );
xor \g456147/U$1_r1 ( \60552 , \60547 , \60551 );
xor \g456147/U$1_r2 ( \60553 , \60543 , \60552 );
xor \g456132/U$1 ( \60554 , \60521 , \60553 );
xor \g131702/U$4 ( \60555 , \60379 , \60443 );
and \g131702/U$3 ( \60556 , \60555 , \60480 );
and \g131702/U$5 ( \60557 , \60379 , \60443 );
or \g131702/U$2 ( \60558 , \60556 , \60557 );
and \g131826/U$2 ( \60559 , \52620 , \52273 );
and \g131826/U$3 ( \60560 , \52270 , \52352 );
nor \g131826/U$1 ( \60561 , \60559 , \60560 );
and \g131785/U$2 ( \60562 , \60561 , \51513 );
not \g131785/U$4 ( \60563 , \60561 );
and \g131785/U$3 ( \60564 , \60563 , \51120 );
nor \g131785/U$1 ( \60565 , \60562 , \60564 );
xor \g132106/U$4 ( \60566 , \60399 , \60407 );
and \g132106/U$3 ( \60567 , \60566 , \60441 );
and \g132106/U$5 ( \60568 , \60399 , \60407 );
or \g132106/U$2 ( \60569 , \60567 , \60568 );
xor \g456135/U$2 ( \60570 , \60565 , \60569 );
xor \g132208/U$4 ( \60571 , \60412 , \60420 );
and \g132208/U$3 ( \60572 , \60571 , \60440 );
and \g132208/U$5 ( \60573 , \60412 , \60420 );
or \g132208/U$2 ( \60574 , \60572 , \60573 );
not \g132596/U$3 ( \60575 , \49568 );
and \g132640/U$2 ( \60576 , \54537 , \49813 );
and \g132640/U$3 ( \60577 , \49812 , \54529 );
nor \g132640/U$1 ( \60578 , \60576 , \60577 );
not \g132596/U$4 ( \60579 , \60578 );
or \g132596/U$2 ( \60580 , \60575 , \60579 );
or \g132596/U$5 ( \60581 , \60578 , \49568 );
nand \g132596/U$1 ( \60582 , \60580 , \60581 );
xor \g132015/U$1 ( \60583 , \60574 , \60582 );
xor \g132209/U$4 ( \60584 , \60349 , \60357 );
and \g132209/U$3 ( \60585 , \60584 , \60362 );
and \g132209/U$5 ( \60586 , \60349 , \60357 );
or \g132209/U$2 ( \60587 , \60585 , \60586 );
not \g132982/U$3 ( \60588 , \48685 );
and \g133011/U$2 ( \60589 , \48860 , \56167 );
and \g133011/U$3 ( \60590 , \48858 , \55884 );
nor \g133011/U$1 ( \60591 , \60589 , \60590 );
not \g132982/U$4 ( \60592 , \60591 );
or \g132982/U$2 ( \60593 , \60588 , \60592 );
or \g132982/U$5 ( \60594 , \60591 , \48685 );
nand \g132982/U$1 ( \60595 , \60593 , \60594 );
xor \g132104/U$1 ( \60596 , \60587 , \60595 );
not \g132711/U$3 ( \60597 , \48159 );
and \g132761/U$2 ( \60598 , \48154 , \56347 );
and \g132761/U$3 ( \60599 , \56349 , \48155 );
nor \g132761/U$1 ( \60600 , \60598 , \60599 );
not \g132711/U$4 ( \60601 , \60600 );
or \g132711/U$2 ( \60602 , \60597 , \60601 );
or \g132711/U$5 ( \60603 , \60600 , \48159 );
nand \g132711/U$1 ( \60604 , \60602 , \60603 );
not \g132809/U$3 ( \60605 , \48323 );
and \g132845/U$2 ( \60606 , \48334 , \56357 );
and \g132845/U$3 ( \60607 , \56359 , \48335 );
nor \g132845/U$1 ( \60608 , \60606 , \60607 );
not \g132809/U$4 ( \60609 , \60608 );
or \g132809/U$2 ( \60610 , \60605 , \60609 );
or \g132809/U$5 ( \60611 , \60608 , \48323 );
nand \g132809/U$1 ( \60612 , \60610 , \60611 );
xor \g132312/U$1 ( \60613 , \60604 , \60612 );
and \g132441/U$2 ( \60614 , \60340 , \60348 );
xor \g132312/U$1_r1 ( \60615 , \60613 , \60614 );
xor \g132104/U$1_r1 ( \60616 , \60596 , \60615 );
xor \g132015/U$1_r1 ( \60617 , \60583 , \60616 );
xor \g456135/U$1 ( \60618 , \60570 , \60617 );
xor \g131802/U$4 ( \60619 , \60386 , \60394 );
and \g131802/U$3 ( \60620 , \60619 , \60442 );
and \g131802/U$5 ( \60621 , \60386 , \60394 );
or \g131802/U$2 ( \60622 , \60620 , \60621 );
not \g131924/U$3 ( \60623 , \51124 );
and \g131967/U$2 ( \60624 , \52978 , \51518 );
and \g131967/U$3 ( \60625 , \51517 , \52883 );
nor \g131967/U$1 ( \60626 , \60624 , \60625 );
not \g131924/U$4 ( \60627 , \60626 );
or \g131924/U$2 ( \60628 , \60623 , \60627 );
or \g131924/U$5 ( \60629 , \60626 , \51124 );
nand \g131924/U$1 ( \60630 , \60628 , \60629 );
not \g132250/U$3 ( \60631 , \50362 );
and \g132301/U$2 ( \60632 , \53848 , \50587 );
and \g132301/U$3 ( \60633 , \50588 , \54015 );
nor \g132301/U$1 ( \60634 , \60632 , \60633 );
not \g132250/U$4 ( \60635 , \60634 );
or \g132250/U$2 ( \60636 , \60631 , \60635 );
or \g132250/U$5 ( \60637 , \60634 , \50362 );
nand \g132250/U$1 ( \60638 , \60636 , \60637 );
xor \g131860/U$1 ( \60639 , \60630 , \60638 );
not \g132743/U$3 ( \60640 , \49233 );
and \g132783/U$2 ( \60641 , \54853 , \49403 );
and \g132783/U$3 ( \60642 , \49405 , \55127 );
nor \g132783/U$1 ( \60643 , \60641 , \60642 );
not \g132743/U$4 ( \60644 , \60643 );
or \g132743/U$2 ( \60645 , \60640 , \60644 );
or \g132743/U$5 ( \60646 , \60643 , \49233 );
nand \g132743/U$1 ( \60647 , \60645 , \60646 );
not \g132874/U$3 ( \60648 , \49014 );
and \g132909/U$2 ( \60649 , \55460 , \49074 );
and \g132909/U$3 ( \60650 , \49075 , \55707 );
nor \g132909/U$1 ( \60651 , \60649 , \60650 );
not \g132874/U$4 ( \60652 , \60651 );
or \g132874/U$2 ( \60653 , \60648 , \60652 );
or \g132874/U$5 ( \60654 , \60651 , \49014 );
nand \g132874/U$1 ( \60655 , \60653 , \60654 );
xor \g131993/U$1 ( \60656 , \60647 , \60655 );
xor \g132317/U$4 ( \60657 , \60429 , \60437 );
and \g132317/U$3 ( \60658 , \60657 , \60439 );
and \g132317/U$5 ( \60659 , \60429 , \60437 );
or \g132317/U$2 ( \60660 , \60658 , \60659 );
not \g132898/U$3 ( \60661 , \48483 );
and \g132942/U$2 ( \60662 , \48478 , \56446 );
and \g132942/U$3 ( \60663 , \56448 , \48479 );
nor \g132942/U$1 ( \60664 , \60662 , \60663 );
not \g132898/U$4 ( \60665 , \60664 );
or \g132898/U$2 ( \60666 , \60661 , \60665 );
or \g132898/U$5 ( \60667 , \60664 , \48483 );
nand \g132898/U$1 ( \60668 , \60666 , \60667 );
xor \g132095/U$1 ( \60669 , \60660 , \60668 );
xor \g132187/U$1 ( \60670 , \56703 , \56711 );
xor \g132187/U$1_r1 ( \60671 , \60670 , \56713 );
xor \g132095/U$1_r1 ( \60672 , \60669 , \60671 );
xor \g131993/U$1_r1 ( \60673 , \60656 , \60672 );
xor \g131860/U$1_r1 ( \60674 , \60639 , \60673 );
xor \g456135/U$1_r1 ( \60675 , \60622 , \60674 );
xor \g456135/U$1_r2 ( \60676 , \60618 , \60675 );
xor \g456132/U$1_r1 ( \60677 , \60558 , \60676 );
xor \g456132/U$1_r2 ( \60678 , \60554 , \60677 );
xor \g130499/U$1 ( \60679 , \60293 , \60484 );
xor \g130499/U$1_r1 ( \60680 , \60679 , \60503 );
and \g130452/U$2 ( \60681 , \60678 , \60680 );
and \g130356/U$3 ( \60682 , \60508 , \60681 );
and \g130356/U$5 ( \60683 , \60506 , \60507 );
or \g130356/U$2 ( \60684 , \60682 , \60683 );
xor \g132095/U$4 ( \60685 , \60660 , \60668 );
and \g132095/U$3 ( \60686 , \60685 , \60671 );
and \g132095/U$5 ( \60687 , \60660 , \60668 );
or \g132095/U$2 ( \60688 , \60686 , \60687 );
xor \g132104/U$4 ( \60689 , \60587 , \60595 );
and \g132104/U$3 ( \60690 , \60689 , \60615 );
and \g132104/U$5 ( \60691 , \60587 , \60595 );
or \g132104/U$2 ( \60692 , \60690 , \60691 );
xor \g131991/U$4 ( \60693 , \60688 , \60692 );
xor \g132094/U$1 ( \60694 , \56687 , \56695 );
xor \g132094/U$1_r1 ( \60695 , \60694 , \56716 );
and \g131991/U$3 ( \60696 , \60693 , \60695 );
and \g131991/U$5 ( \60697 , \60688 , \60692 );
or \g131991/U$2 ( \60698 , \60696 , \60697 );
not \g131784/U$3 ( \60699 , \51124 );
and \g131825/U$2 ( \60700 , \52620 , \51518 );
and \g131825/U$3 ( \60701 , \51517 , \52352 );
nor \g131825/U$1 ( \60702 , \60700 , \60701 );
not \g131784/U$4 ( \60703 , \60702 );
or \g131784/U$2 ( \60704 , \60699 , \60703 );
or \g131784/U$5 ( \60705 , \60702 , \51124 );
nand \g131784/U$1 ( \60706 , \60704 , \60705 );
xor \g131608/U$1 ( \60707 , \60698 , \60706 );
and \g131699/U$2 ( \60708 , \52108 , \52273 );
and \g131699/U$3 ( \60709 , \52270 , \51854 );
nor \g131699/U$1 ( \60710 , \60708 , \60709 );
and \g131656/U$2 ( \60711 , \60710 , \51513 );
not \g131656/U$4 ( \60712 , \60710 );
and \g131656/U$3 ( \60713 , \60712 , \51120 );
nor \g131656/U$1 ( \60714 , \60711 , \60713 );
xor \g131608/U$1_r1 ( \60715 , \60707 , \60714 );
and \g131767/U$2 ( \60716 , \52108 , \52270 );
and \g131767/U$3 ( \60717 , \52273 , \52352 );
nor \g131767/U$1 ( \60718 , \60716 , \60717 );
and \g131724/U$2 ( \60719 , \60718 , \51513 );
not \g131724/U$4 ( \60720 , \60718 );
and \g131724/U$3 ( \60721 , \60720 , \51120 );
nor \g131724/U$1 ( \60722 , \60719 , \60721 );
xor \g132015/U$4 ( \60723 , \60574 , \60582 );
and \g132015/U$3 ( \60724 , \60723 , \60616 );
and \g132015/U$5 ( \60725 , \60574 , \60582 );
or \g132015/U$2 ( \60726 , \60724 , \60725 );
xor \g131666/U$4 ( \60727 , \60722 , \60726 );
not \g132341/U$3 ( \60728 , \49925 );
and \g132423/U$2 ( \60729 , \54185 , \50160 );
and \g132423/U$3 ( \60730 , \50159 , \54015 );
nor \g132423/U$1 ( \60731 , \60729 , \60730 );
not \g132341/U$4 ( \60732 , \60731 );
or \g132341/U$2 ( \60733 , \60728 , \60732 );
or \g132341/U$5 ( \60734 , \60731 , \49925 );
nand \g132341/U$1 ( \60735 , \60733 , \60734 );
not \g132528/U$3 ( \60736 , \49568 );
and \g132569/U$2 ( \60737 , \54251 , \49812 );
and \g132569/U$3 ( \60738 , \49813 , \54529 );
nor \g132569/U$1 ( \60739 , \60737 , \60738 );
not \g132528/U$4 ( \60740 , \60739 );
or \g132528/U$2 ( \60741 , \60736 , \60740 );
or \g132528/U$5 ( \60742 , \60739 , \49568 );
nand \g132528/U$1 ( \60743 , \60741 , \60742 );
xor \g131992/U$1 ( \60744 , \60735 , \60743 );
xor \g132312/U$4 ( \60745 , \60604 , \60612 );
and \g132312/U$3 ( \60746 , \60745 , \60614 );
and \g132312/U$5 ( \60747 , \60604 , \60612 );
or \g132312/U$2 ( \60748 , \60746 , \60747 );
not \g132907/U$3 ( \60749 , \48483 );
and \g132940/U$2 ( \60750 , \48479 , \56446 );
and \g132940/U$3 ( \60751 , \56167 , \48478 );
nor \g132940/U$1 ( \60752 , \60750 , \60751 );
not \g132907/U$4 ( \60753 , \60752 );
or \g132907/U$2 ( \60754 , \60749 , \60753 );
or \g132907/U$5 ( \60755 , \60752 , \48483 );
nand \g132907/U$1 ( \60756 , \60754 , \60755 );
xor \g132093/U$1 ( \60757 , \60748 , \60756 );
xor \g132186/U$1 ( \60758 , \56417 , \56425 );
xor \g132186/U$1_r1 ( \60759 , \60758 , \56441 );
xor \g132093/U$1_r1 ( \60760 , \60757 , \60759 );
xor \g131992/U$1_r1 ( \60761 , \60744 , \60760 );
and \g131666/U$3 ( \60762 , \60727 , \60761 );
and \g131666/U$5 ( \60763 , \60722 , \60726 );
or \g131666/U$2 ( \60764 , \60762 , \60763 );
xor \g456126/U$2 ( \60765 , \60715 , \60764 );
not \g132005/U$3 ( \60766 , \50759 );
and \g132045/U$2 ( \60767 , \52978 , \51053 );
and \g132045/U$3 ( \60768 , \51055 , \53300 );
nor \g132045/U$1 ( \60769 , \60767 , \60768 );
not \g132005/U$4 ( \60770 , \60769 );
or \g132005/U$2 ( \60771 , \60766 , \60770 );
or \g132005/U$5 ( \60772 , \60769 , \50759 );
nand \g132005/U$1 ( \60773 , \60771 , \60772 );
not \g132806/U$3 ( \60774 , \49014 );
and \g132860/U$2 ( \60775 , \55127 , \49074 );
and \g132860/U$3 ( \60776 , \49075 , \55460 );
nor \g132860/U$1 ( \60777 , \60775 , \60776 );
not \g132806/U$4 ( \60778 , \60777 );
or \g132806/U$2 ( \60779 , \60774 , \60778 );
or \g132806/U$5 ( \60780 , \60777 , \49014 );
nand \g132806/U$1 ( \60781 , \60779 , \60780 );
not \g132936/U$3 ( \60782 , \48685 );
and \g132961/U$2 ( \60783 , \48860 , \55884 );
and \g132961/U$3 ( \60784 , \48858 , \55707 );
nor \g132961/U$1 ( \60785 , \60783 , \60784 );
not \g132936/U$4 ( \60786 , \60785 );
or \g132936/U$2 ( \60787 , \60782 , \60786 );
or \g132936/U$5 ( \60788 , \60785 , \48685 );
nand \g132936/U$1 ( \60789 , \60787 , \60788 );
xor \g132630/U$1 ( \60790 , \60781 , \60789 );
not \g132679/U$3 ( \60791 , \49233 );
and \g132728/U$2 ( \60792 , \54853 , \49405 );
and \g132728/U$3 ( \60793 , \49403 , \54537 );
nor \g132728/U$1 ( \60794 , \60792 , \60793 );
not \g132679/U$4 ( \60795 , \60794 );
or \g132679/U$2 ( \60796 , \60791 , \60795 );
or \g132679/U$5 ( \60797 , \60794 , \49233 );
nand \g132679/U$1 ( \60798 , \60796 , \60797 );
xor \g132630/U$1_r1 ( \60799 , \60790 , \60798 );
xor \g131904/U$4 ( \60800 , \60773 , \60799 );
xor \g131993/U$4 ( \60801 , \60647 , \60655 );
and \g131993/U$3 ( \60802 , \60801 , \60672 );
and \g131993/U$5 ( \60803 , \60647 , \60655 );
or \g131993/U$2 ( \60804 , \60802 , \60803 );
and \g131904/U$3 ( \60805 , \60800 , \60804 );
and \g131904/U$5 ( \60806 , \60773 , \60799 );
or \g131904/U$2 ( \60807 , \60805 , \60806 );
xor \g131992/U$4 ( \60808 , \60735 , \60743 );
and \g131992/U$3 ( \60809 , \60808 , \60760 );
and \g131992/U$5 ( \60810 , \60735 , \60743 );
or \g131992/U$2 ( \60811 , \60809 , \60810 );
xor \g131798/U$1 ( \60812 , \60807 , \60811 );
xor \g132093/U$4 ( \60813 , \60748 , \60756 );
and \g132093/U$3 ( \60814 , \60813 , \60759 );
and \g132093/U$5 ( \60815 , \60748 , \60756 );
or \g132093/U$2 ( \60816 , \60814 , \60815 );
not \g132610/U$3 ( \60817 , \49233 );
and \g132655/U$2 ( \60818 , \54537 , \49405 );
and \g132655/U$3 ( \60819 , \49403 , \54529 );
nor \g132655/U$1 ( \60820 , \60818 , \60819 );
not \g132610/U$4 ( \60821 , \60820 );
or \g132610/U$2 ( \60822 , \60817 , \60821 );
or \g132610/U$5 ( \60823 , \60820 , \49233 );
nand \g132610/U$1 ( \60824 , \60822 , \60823 );
xor \g131903/U$1 ( \60825 , \60816 , \60824 );
xor \g131994/U$1 ( \60826 , \56719 , \56727 );
xor \g131994/U$1_r1 ( \60827 , \60826 , \56730 );
xor \g131903/U$1_r1 ( \60828 , \60825 , \60827 );
xor \g131798/U$1_r1 ( \60829 , \60812 , \60828 );
xor \g456126/U$1 ( \60830 , \60765 , \60829 );
xor \g456135/U$9 ( \60831 , \60565 , \60569 );
xor \g456135/U$9_r1 ( \60832 , \60831 , \60617 );
and \g456135/U$8 ( \60833 , \60622 , \60832 );
xor \g456135/U$11 ( \60834 , \60565 , \60569 );
xor \g456135/U$11_r1 ( \60835 , \60834 , \60617 );
and \g456135/U$10 ( \60836 , \60674 , \60835 );
and \g456135/U$12 ( \60837 , \60622 , \60674 );
or \g456135/U$7 ( \60838 , \60833 , \60836 , \60837 );
xor \g131666/U$1 ( \60839 , \60722 , \60726 );
xor \g131666/U$1_r1 ( \60840 , \60839 , \60761 );
xor \g131561/U$4 ( \60841 , \60838 , \60840 );
xor \g131860/U$4 ( \60842 , \60630 , \60638 );
and \g131860/U$3 ( \60843 , \60842 , \60673 );
and \g131860/U$5 ( \60844 , \60630 , \60638 );
or \g131860/U$2 ( \60845 , \60843 , \60844 );
xor \g456147/U$5 ( \60846 , \60529 , \60537 );
and \g456147/U$4 ( \60847 , \60846 , \60542 );
and \g456147/U$6 ( \60848 , \60529 , \60537 );
or \g456147/U$3 ( \60849 , \60847 , \60848 );
xor \g131775/U$1 ( \60850 , \60845 , \60849 );
xor \g131904/U$1 ( \60851 , \60773 , \60799 );
xor \g131904/U$1_r1 ( \60852 , \60851 , \60804 );
xor \g131775/U$1_r1 ( \60853 , \60850 , \60852 );
and \g131561/U$3 ( \60854 , \60841 , \60853 );
and \g131561/U$5 ( \60855 , \60838 , \60840 );
or \g131561/U$2 ( \60856 , \60854 , \60855 );
xor \g131775/U$4 ( \60857 , \60845 , \60849 );
and \g131775/U$3 ( \60858 , \60857 , \60852 );
and \g131775/U$5 ( \60859 , \60845 , \60849 );
or \g131775/U$2 ( \60860 , \60858 , \60859 );
xor \g456147/U$9 ( \60861 , \60529 , \60537 );
xor \g456147/U$9_r1 ( \60862 , \60861 , \60542 );
and \g456147/U$8 ( \60863 , \60547 , \60862 );
xor \g456147/U$11 ( \60864 , \60529 , \60537 );
xor \g456147/U$11_r1 ( \60865 , \60864 , \60542 );
and \g456147/U$10 ( \60866 , \60551 , \60865 );
and \g456147/U$12 ( \60867 , \60547 , \60551 );
or \g456147/U$7 ( \60868 , \60863 , \60866 , \60867 );
xor \g456135/U$5 ( \60869 , \60565 , \60569 );
and \g456135/U$4 ( \60870 , \60869 , \60617 );
and \g456135/U$6 ( \60871 , \60565 , \60569 );
or \g456135/U$3 ( \60872 , \60870 , \60871 );
xor \g131639/U$4 ( \60873 , \60868 , \60872 );
not \g131851/U$3 ( \60874 , \51124 );
and \g131901/U$2 ( \60875 , \52620 , \51517 );
and \g131901/U$3 ( \60876 , \51518 , \52883 );
nor \g131901/U$1 ( \60877 , \60875 , \60876 );
not \g131851/U$4 ( \60878 , \60877 );
or \g131851/U$2 ( \60879 , \60874 , \60878 );
or \g131851/U$5 ( \60880 , \60877 , \51124 );
nand \g131851/U$1 ( \60881 , \60879 , \60880 );
not \g132150/U$3 ( \60882 , \50362 );
and \g132198/U$2 ( \60883 , \53610 , \50587 );
and \g132198/U$3 ( \60884 , \50588 , \53848 );
nor \g132198/U$1 ( \60885 , \60883 , \60884 );
not \g132150/U$4 ( \60886 , \60885 );
or \g132150/U$2 ( \60887 , \60882 , \60886 );
or \g132150/U$5 ( \60888 , \60885 , \50362 );
nand \g132150/U$1 ( \60889 , \60887 , \60888 );
xor \g131799/U$1 ( \60890 , \60881 , \60889 );
xor \g131991/U$1 ( \60891 , \60688 , \60692 );
xor \g131991/U$1_r1 ( \60892 , \60891 , \60695 );
xor \g131799/U$1_r1 ( \60893 , \60890 , \60892 );
and \g131639/U$3 ( \60894 , \60873 , \60893 );
and \g131639/U$5 ( \60895 , \60868 , \60872 );
or \g131639/U$2 ( \60896 , \60894 , \60895 );
xor \g131560/U$1 ( \60897 , \60860 , \60896 );
xor \g131799/U$4 ( \60898 , \60881 , \60889 );
and \g131799/U$3 ( \60899 , \60898 , \60892 );
and \g131799/U$5 ( \60900 , \60881 , \60889 );
or \g131799/U$2 ( \60901 , \60899 , \60900 );
not \g132450/U$3 ( \60902 , \49568 );
and \g132497/U$2 ( \60903 , \54185 , \49812 );
and \g132497/U$3 ( \60904 , \49813 , \54251 );
nor \g132497/U$1 ( \60905 , \60903 , \60904 );
not \g132450/U$4 ( \60906 , \60905 );
or \g132450/U$2 ( \60907 , \60902 , \60906 );
or \g132450/U$5 ( \60908 , \60905 , \49568 );
nand \g132450/U$1 ( \60909 , \60907 , \60908 );
xor \g132630/U$4 ( \60910 , \60781 , \60789 );
and \g132630/U$3 ( \60911 , \60910 , \60798 );
and \g132630/U$5 ( \60912 , \60781 , \60789 );
or \g132630/U$2 ( \60913 , \60911 , \60912 );
xor \g132185/U$1 ( \60914 , \60909 , \60913 );
not \g132249/U$3 ( \60915 , \49925 );
and \g132300/U$2 ( \60916 , \53848 , \50159 );
and \g132300/U$3 ( \60917 , \50160 , \54015 );
nor \g132300/U$1 ( \60918 , \60916 , \60917 );
not \g132249/U$4 ( \60919 , \60918 );
or \g132249/U$2 ( \60920 , \60915 , \60919 );
or \g132249/U$5 ( \60921 , \60918 , \49925 );
nand \g132249/U$1 ( \60922 , \60920 , \60921 );
xor \g132185/U$1_r1 ( \60923 , \60914 , \60922 );
xor \g131714/U$1 ( \60924 , \60901 , \60923 );
not \g131923/U$3 ( \60925 , \50759 );
and \g131959/U$2 ( \60926 , \52978 , \51055 );
and \g131959/U$3 ( \60927 , \51053 , \52883 );
nor \g131959/U$1 ( \60928 , \60926 , \60927 );
not \g131923/U$4 ( \60929 , \60928 );
or \g131923/U$2 ( \60930 , \60925 , \60929 );
or \g131923/U$5 ( \60931 , \60928 , \50759 );
nand \g131923/U$1 ( \60932 , \60930 , \60931 );
not \g132083/U$3 ( \60933 , \50362 );
and \g132126/U$2 ( \60934 , \53610 , \50588 );
and \g132126/U$3 ( \60935 , \50587 , \53300 );
nor \g132126/U$1 ( \60936 , \60934 , \60935 );
not \g132083/U$4 ( \60937 , \60936 );
or \g132083/U$2 ( \60938 , \60933 , \60937 );
or \g132083/U$5 ( \60939 , \60936 , \50362 );
nand \g132083/U$1 ( \60940 , \60938 , \60939 );
xor \g131797/U$1 ( \60941 , \60932 , \60940 );
xor \g131869/U$1 ( \60942 , \56399 , \56407 );
xor \g131869/U$1_r1 ( \60943 , \60942 , \56489 );
xor \g131797/U$1_r1 ( \60944 , \60941 , \60943 );
xor \g131714/U$1_r1 ( \60945 , \60924 , \60944 );
xor \g131560/U$1_r1 ( \60946 , \60897 , \60945 );
xor \g456126/U$1_r1 ( \60947 , \60856 , \60946 );
xor \g456126/U$1_r2 ( \60948 , \60830 , \60947 );
xor \g130183/U$4 ( \60949 , \60684 , \60948 );
xor \g131639/U$1 ( \60950 , \60868 , \60872 );
xor \g131639/U$1_r1 ( \60951 , \60950 , \60893 );
xor \g131561/U$1 ( \60952 , \60838 , \60840 );
xor \g131561/U$1_r1 ( \60953 , \60952 , \60853 );
xor \g456128/U$1 ( \60954 , \60951 , \60953 );
xor \g456132/U$5 ( \60955 , \60512 , \60520 );
and \g456132/U$4 ( \60956 , \60955 , \60553 );
and \g456132/U$6 ( \60957 , \60512 , \60520 );
or \g456132/U$3 ( \60958 , \60956 , \60957 );
xor \g456128/U$1_r1 ( \60959 , \60954 , \60958 );
xor \g456132/U$9 ( \60960 , \60512 , \60520 );
xor \g456132/U$9_r1 ( \60961 , \60960 , \60553 );
and \g456132/U$8 ( \60962 , \60558 , \60961 );
xor \g456132/U$11 ( \60963 , \60512 , \60520 );
xor \g456132/U$11_r1 ( \60964 , \60963 , \60553 );
and \g456132/U$10 ( \60965 , \60676 , \60964 );
and \g456132/U$12 ( \60966 , \60558 , \60676 );
or \g456132/U$7 ( \60967 , \60962 , \60965 , \60966 );
xor \g130280/U$4 ( \60968 , \60959 , \60967 );
xor \g130356/U$1 ( \60969 , \60506 , \60507 );
xor \g130356/U$1_r1 ( \60970 , \60969 , \60681 );
and \g130280/U$3 ( \60971 , \60968 , \60970 );
and \g130280/U$5 ( \60972 , \60959 , \60967 );
or \g130280/U$2 ( \60973 , \60971 , \60972 );
and \g130183/U$3 ( \60974 , \60949 , \60973 );
and \g130183/U$5 ( \60975 , \60684 , \60948 );
or \g130183/U$2 ( \60976 , \60974 , \60975 );
nand \g132364/U$1 ( \60977 , \47026 , \40061 );
not \g132363/U$1 ( \60978 , \60977 );
and \g130075/U$2 ( \60979 , \60976 , \60978 );
not \g130097/U$3 ( \60980 , \60976 );
not \g130097/U$4 ( \60981 , \60978 );
and \g130097/U$2 ( \60982 , \60980 , \60981 );
xor \g456128/U$4 ( \60983 , \60951 , \60953 );
and \g456128/U$3 ( \60984 , \60983 , \60958 );
and \g456128/U$5 ( \60985 , \60951 , \60953 );
nor \g456128/U$2 ( \60986 , \60984 , \60985 );
not \g130143/U$2 ( \60987 , \60986 );
xor \g130183/U$1 ( \60988 , \60684 , \60948 );
xor \g130183/U$1_r1 ( \60989 , \60988 , \60973 );
nand \g130143/U$1 ( \60990 , \60987 , \60989 );
nor \g130097/U$1 ( \60991 , \60982 , \60990 );
nor \g130075/U$1 ( \60992 , \60979 , \60991 );
not \g129857/U$2 ( \60993 , \60992 );
xor \g456126/U$9 ( \60994 , \60715 , \60764 );
xor \g456126/U$9_r1 ( \60995 , \60994 , \60829 );
and \g456126/U$8 ( \60996 , \60856 , \60995 );
xor \g456126/U$11 ( \60997 , \60715 , \60764 );
xor \g456126/U$11_r1 ( \60998 , \60997 , \60829 );
and \g456126/U$10 ( \60999 , \60946 , \60998 );
and \g456126/U$12 ( \61000 , \60856 , \60946 );
or \g456126/U$7 ( \61001 , \60996 , \60999 , \61000 );
xor \g131608/U$4 ( \61002 , \60698 , \60706 );
and \g131608/U$3 ( \61003 , \61002 , \60714 );
and \g131608/U$5 ( \61004 , \60698 , \60706 );
or \g131608/U$2 ( \61005 , \61003 , \61004 );
xor \g131674/U$1 ( \61006 , \56774 , \56782 );
xor \g131674/U$1_r1 ( \61007 , \61006 , \56791 );
xor \g456122/U$2 ( \61008 , \61005 , \61007 );
xor \g131797/U$4 ( \61009 , \60932 , \60940 );
and \g131797/U$3 ( \61010 , \61009 , \60943 );
and \g131797/U$5 ( \61011 , \60932 , \60940 );
or \g131797/U$2 ( \61012 , \61010 , \61011 );
xor \g456122/U$1 ( \61013 , \61008 , \61012 );
xor \g456126/U$5 ( \61014 , \60715 , \60764 );
and \g456126/U$4 ( \61015 , \61014 , \60829 );
and \g456126/U$6 ( \61016 , \60715 , \60764 );
or \g456126/U$3 ( \61017 , \61015 , \61016 );
xor \g131903/U$4 ( \61018 , \60816 , \60824 );
and \g131903/U$3 ( \61019 , \61018 , \60827 );
and \g131903/U$5 ( \61020 , \60816 , \60824 );
or \g131903/U$2 ( \61021 , \61019 , \61020 );
xor \g132185/U$4 ( \61022 , \60909 , \60913 );
and \g132185/U$3 ( \61023 , \61022 , \60922 );
and \g132185/U$5 ( \61024 , \60909 , \60913 );
or \g132185/U$2 ( \61025 , \61023 , \61024 );
xor \g131715/U$1 ( \61026 , \61021 , \61025 );
xor \g456145/U$2 ( \61027 , \56336 , \56344 );
xor \g456145/U$1 ( \61028 , \61027 , \56389 );
xor \g456145/U$1_r1 ( \61029 , \56328 , \56492 );
xor \g456145/U$1_r2 ( \61030 , \61028 , \61029 );
xor \g131715/U$1_r1 ( \61031 , \61026 , \61030 );
xor \g456122/U$1_r1 ( \61032 , \61017 , \61031 );
xor \g456122/U$1_r2 ( \61033 , \61013 , \61032 );
xor \g131560/U$4 ( \61034 , \60860 , \60896 );
and \g131560/U$3 ( \61035 , \61034 , \60945 );
and \g131560/U$5 ( \61036 , \60860 , \60896 );
or \g131560/U$2 ( \61037 , \61035 , \61036 );
xor \g456037/U$9 ( \61038 , \61033 , \61037 );
xor \g456125/U$2 ( \61039 , \56678 , \56685 );
xor \g456125/U$1 ( \61040 , \61039 , \56763 );
xor \g131798/U$4 ( \61041 , \60807 , \60811 );
and \g131798/U$3 ( \61042 , \61041 , \60828 );
and \g131798/U$5 ( \61043 , \60807 , \60811 );
or \g131798/U$2 ( \61044 , \61042 , \61043 );
xor \g131714/U$4 ( \61045 , \60901 , \60923 );
and \g131714/U$3 ( \61046 , \61045 , \60944 );
and \g131714/U$5 ( \61047 , \60901 , \60923 );
or \g131714/U$2 ( \61048 , \61046 , \61047 );
xor \g456125/U$1_r1 ( \61049 , \61044 , \61048 );
xor \g456125/U$1_r2 ( \61050 , \61040 , \61049 );
xor \g456037/U$9_r1 ( \61051 , \61038 , \61050 );
and \g456037/U$8 ( \61052 , \61001 , \61051 );
not \g130040/U$3 ( \61053 , \60977 );
not \g130058/U$3 ( \61054 , \60976 );
not \g130058/U$4 ( \61055 , \60990 );
or \g130058/U$2 ( \61056 , \61054 , \61055 );
or \g130058/U$5 ( \61057 , \60990 , \60976 );
nand \g130058/U$1 ( \61058 , \61056 , \61057 );
not \g130040/U$4 ( \61059 , \61058 );
or \g130040/U$2 ( \61060 , \61053 , \61059 );
or \g130040/U$5 ( \61061 , \61058 , \60977 );
nand \g130040/U$1 ( \61062 , \61060 , \61061 );
xor \g456037/U$11 ( \61063 , \61033 , \61037 );
xor \g456037/U$11_r1 ( \61064 , \61063 , \61050 );
and \g456037/U$10 ( \61065 , \61062 , \61064 );
and \g456037/U$12 ( \61066 , \61001 , \61062 );
or \g456037/U$7 ( \61067 , \61052 , \61065 , \61066 );
nand \g129857/U$1 ( \61068 , \60993 , \61067 );
not \g129691/U$2 ( \61069 , \61068 );
xor \g456037/U$5 ( \61070 , \61033 , \61037 );
and \g456037/U$4 ( \61071 , \61070 , \61050 );
and \g456037/U$6 ( \61072 , \61033 , \61037 );
or \g456037/U$3 ( \61073 , \61071 , \61072 );
xor \g131715/U$4 ( \61074 , \61021 , \61025 );
and \g131715/U$3 ( \61075 , \61074 , \61030 );
and \g131715/U$5 ( \61076 , \61021 , \61025 );
or \g131715/U$2 ( \61077 , \61075 , \61076 );
xor \g456127/U$2 ( \61078 , \56837 , \56845 );
xor \g456127/U$1 ( \61079 , \61078 , \56850 );
xor \g456127/U$1_r1 ( \61080 , \56870 , \56881 );
xor \g456127/U$1_r2 ( \61081 , \61079 , \61080 );
xor \g131420/U$1 ( \61082 , \61077 , \61081 );
xor \g131672/U$1 ( \61083 , \56497 , \56523 );
xor \g131672/U$1_r1 ( \61084 , \61083 , \56659 );
xor \g131420/U$1_r1 ( \61085 , \61082 , \61084 );
xor \g456122/U$9 ( \61086 , \61005 , \61007 );
xor \g456122/U$9_r1 ( \61087 , \61086 , \61012 );
and \g456122/U$8 ( \61088 , \61017 , \61087 );
xor \g456122/U$11 ( \61089 , \61005 , \61007 );
xor \g456122/U$11_r1 ( \61090 , \61089 , \61012 );
and \g456122/U$10 ( \61091 , \61031 , \61090 );
and \g456122/U$12 ( \61092 , \61017 , \61031 );
or \g456122/U$7 ( \61093 , \61088 , \61091 , \61092 );
xor \g456026/U$9 ( \61094 , \61085 , \61093 );
xor \g456117/U$2 ( \61095 , \56766 , \56794 );
xor \g456117/U$1 ( \61096 , \61095 , \56817 );
xor \g456122/U$5 ( \61097 , \61005 , \61007 );
and \g456122/U$4 ( \61098 , \61097 , \61012 );
and \g456122/U$6 ( \61099 , \61005 , \61007 );
or \g456122/U$3 ( \61100 , \61098 , \61099 );
xor \g456125/U$9 ( \61101 , \56678 , \56685 );
xor \g456125/U$9_r1 ( \61102 , \61101 , \56763 );
and \g456125/U$8 ( \61103 , \61044 , \61102 );
xor \g456125/U$11 ( \61104 , \56678 , \56685 );
xor \g456125/U$11_r1 ( \61105 , \61104 , \56763 );
and \g456125/U$10 ( \61106 , \61048 , \61105 );
and \g456125/U$12 ( \61107 , \61044 , \61048 );
or \g456125/U$7 ( \61108 , \61103 , \61106 , \61107 );
xor \g456117/U$1_r1 ( \61109 , \61100 , \61108 );
xor \g456117/U$1_r2 ( \61110 , \61096 , \61109 );
xor \g456026/U$9_r1 ( \61111 , \61094 , \61110 );
and \g456026/U$8 ( \61112 , \61073 , \61111 );
not \g129844/U$3 ( \61113 , \60992 );
not \g129844/U$4 ( \61114 , \61067 );
or \g129844/U$2 ( \61115 , \61113 , \61114 );
or \g129844/U$5 ( \61116 , \61067 , \60992 );
nand \g129844/U$1 ( \61117 , \61115 , \61116 );
xor \g456026/U$11 ( \61118 , \61085 , \61093 );
xor \g456026/U$11_r1 ( \61119 , \61118 , \61110 );
and \g456026/U$10 ( \61120 , \61117 , \61119 );
and \g456026/U$12 ( \61121 , \61073 , \61117 );
or \g456026/U$7 ( \61122 , \61112 , \61120 , \61121 );
nand \g129691/U$1 ( \61123 , \61069 , \61122 );
not \g129489/U$2 ( \61124 , \61123 );
xor \g131344/U$1 ( \61125 , \56662 , \56820 );
xor \g131344/U$1_r1 ( \61126 , \61125 , \56863 );
xor \g456113/U$2 ( \61127 , \56886 , \56912 );
xor \g456113/U$1 ( \61128 , \61127 , \57006 );
xor \g131557/U$1 ( \61129 , \57358 , \57362 );
xor \g131557/U$1_r1 ( \61130 , \61129 , \57379 );
xor \g131420/U$4 ( \61131 , \61077 , \61081 );
and \g131420/U$3 ( \61132 , \61131 , \61084 );
and \g131420/U$5 ( \61133 , \61077 , \61081 );
or \g131420/U$2 ( \61134 , \61132 , \61133 );
xor \g456113/U$1_r1 ( \61135 , \61130 , \61134 );
xor \g456113/U$1_r2 ( \61136 , \61128 , \61135 );
xor \g456108/U$1 ( \61137 , \61126 , \61136 );
xor \g456117/U$9 ( \61138 , \56766 , \56794 );
xor \g456117/U$9_r1 ( \61139 , \61138 , \56817 );
and \g456117/U$8 ( \61140 , \61100 , \61139 );
xor \g456117/U$11 ( \61141 , \56766 , \56794 );
xor \g456117/U$11_r1 ( \61142 , \61141 , \56817 );
and \g456117/U$10 ( \61143 , \61108 , \61142 );
and \g456117/U$12 ( \61144 , \61100 , \61108 );
or \g456117/U$7 ( \61145 , \61140 , \61143 , \61144 );
xor \g456108/U$1_r1 ( \61146 , \61137 , \61145 );
xor \g456026/U$5 ( \61147 , \61085 , \61093 );
and \g456026/U$4 ( \61148 , \61147 , \61110 );
and \g456026/U$6 ( \61149 , \61085 , \61093 );
or \g456026/U$3 ( \61150 , \61148 , \61149 );
xor \g129524/U$4 ( \61151 , \61146 , \61150 );
not \g129682/U$3 ( \61152 , \61068 );
not \g129682/U$4 ( \61153 , \61122 );
or \g129682/U$2 ( \61154 , \61152 , \61153 );
or \g129682/U$5 ( \61155 , \61122 , \61068 );
nand \g129682/U$1 ( \61156 , \61154 , \61155 );
and \g129524/U$3 ( \61157 , \61151 , \61156 );
and \g129524/U$5 ( \61158 , \61146 , \61150 );
or \g129524/U$2 ( \61159 , \61157 , \61158 );
nand \g129489/U$1 ( \61160 , \61124 , \61159 );
not \g129244/U$3 ( \61161 , \61160 );
not \g129480/U$3 ( \61162 , \61159 );
not \g129480/U$4 ( \61163 , \61123 );
and \g129480/U$2 ( \61164 , \61162 , \61163 );
and \g129480/U$5 ( \61165 , \61159 , \61123 );
nor \g129480/U$1 ( \61166 , \61164 , \61165 );
xor \g456108/U$4 ( \61167 , \61126 , \61136 );
and \g456108/U$3 ( \61168 , \61167 , \61145 );
and \g456108/U$5 ( \61169 , \61126 , \61136 );
nor \g456108/U$2 ( \61170 , \61168 , \61169 );
or \g129286/U$2 ( \61171 , \61166 , \61170 );
xnor \g129387/U$1 ( \61172 , \61170 , \61166 );
not \g129323/U$2 ( \61173 , \61172 );
xor \g456113/U$9 ( \61174 , \56886 , \56912 );
xor \g456113/U$9_r1 ( \61175 , \61174 , \57006 );
and \g456113/U$8 ( \61176 , \61130 , \61175 );
xor \g456113/U$11 ( \61177 , \56886 , \56912 );
xor \g456113/U$11_r1 ( \61178 , \61177 , \57006 );
and \g456113/U$10 ( \61179 , \61134 , \61178 );
and \g456113/U$12 ( \61180 , \61130 , \61134 );
or \g456113/U$7 ( \61181 , \61176 , \61179 , \61180 );
xor \g456109/U$2 ( \61182 , \57384 , \57388 );
xor \g456109/U$1 ( \61183 , \61182 , \57397 );
xor \g456109/U$1_r1 ( \61184 , \57382 , \57403 );
xor \g456109/U$1_r2 ( \61185 , \61183 , \61184 );
xor \g131199/U$1 ( \61186 , \61181 , \61185 );
xor \g131278/U$1 ( \61187 , \56866 , \57009 );
xor \g131278/U$1_r1 ( \61188 , \61187 , \57064 );
xor \g131199/U$1_r1 ( \61189 , \61186 , \61188 );
nand \g129323/U$1 ( \61190 , \61173 , \61189 );
nand \g129286/U$1 ( \61191 , \61171 , \61190 );
not \g129244/U$4 ( \61192 , \61191 );
or \g129244/U$2 ( \61193 , \61161 , \61192 );
or \g129244/U$5 ( \61194 , \61191 , \61160 );
nand \g129244/U$1 ( \61195 , \61193 , \61194 );
xor \g131199/U$4 ( \61196 , \61181 , \61185 );
and \g131199/U$3 ( \61197 , \61196 , \61188 );
and \g131199/U$5 ( \61198 , \61181 , \61185 );
or \g131199/U$2 ( \61199 , \61197 , \61198 );
and \g129063/U$2 ( \61200 , \61195 , \61199 );
not \g131092/U$3 ( \61201 , \57350 );
not \g131118/U$3 ( \61202 , \57490 );
not \g131118/U$4 ( \61203 , \57067 );
and \g131118/U$2 ( \61204 , \61202 , \61203 );
and \g131118/U$5 ( \61205 , \57490 , \57067 );
nor \g131118/U$1 ( \61206 , \61204 , \61205 );
not \g131092/U$4 ( \61207 , \61206 );
or \g131092/U$2 ( \61208 , \61201 , \61207 );
or \g131092/U$5 ( \61209 , \61206 , \57350 );
nand \g131092/U$1 ( \61210 , \61208 , \61209 );
xor \g129173/U$1 ( \61211 , \61199 , \61195 );
and \g129106/U$2 ( \61212 , \61210 , \61211 );
nor \g129063/U$1 ( \61213 , \61200 , \61212 );
not \g129022/U$3 ( \61214 , \61213 );
nor \g129283/U$1 ( \61215 , \61190 , \61160 );
not \g129022/U$4 ( \61216 , \61215 );
and \g129022/U$2 ( \61217 , \61214 , \61216 );
and \g129022/U$5 ( \61218 , \61213 , \61215 );
nor \g129022/U$1 ( \61219 , \61217 , \61218 );
xnor \g128998/U$1 ( \61220 , \57492 , \61219 );
not \g128948/U$2 ( \61221 , \61220 );
not \g131196/U$3 ( \61222 , \57486 );
not \g131196/U$4 ( \61223 , \57476 );
or \g131196/U$2 ( \61224 , \61222 , \61223 );
or \g131203/U$2 ( \61225 , \57476 , \57486 );
nand \g131203/U$1 ( \61226 , \61225 , \57408 );
nand \g131196/U$1 ( \61227 , \61224 , \61226 );
xor \g456112/U$9 ( \61228 , \57087 , \57144 );
xor \g456112/U$9_r1 ( \61229 , \61228 , \57149 );
and \g456112/U$8 ( \61230 , \57164 , \61229 );
xor \g456112/U$11 ( \61231 , \57087 , \57144 );
xor \g456112/U$11_r1 ( \61232 , \61231 , \57149 );
and \g456112/U$10 ( \61233 , \57348 , \61232 );
and \g456112/U$12 ( \61234 , \57164 , \57348 );
or \g456112/U$7 ( \61235 , \61230 , \61233 , \61234 );
xor \g130974/U$1 ( \61236 , \61227 , \61235 );
xor \g456142/U$9 ( \61237 , \57168 , \57176 );
xor \g456142/U$9_r1 ( \61238 , \61237 , \57226 );
and \g456142/U$8 ( \61239 , \57292 , \61238 );
xor \g456142/U$11 ( \61240 , \57168 , \57176 );
xor \g456142/U$11_r1 ( \61241 , \61240 , \57226 );
and \g456142/U$10 ( \61242 , \57346 , \61241 );
and \g456142/U$12 ( \61243 , \57292 , \57346 );
or \g456142/U$7 ( \61244 , \61239 , \61242 , \61243 );
not \g131654/U$3 ( \61245 , \50362 );
and \g131688/U$2 ( \61246 , \52108 , \50588 );
and \g131688/U$3 ( \61247 , \50587 , \51854 );
nor \g131688/U$1 ( \61248 , \61246 , \61247 );
not \g131654/U$4 ( \61249 , \61248 );
or \g131654/U$2 ( \61250 , \61245 , \61249 );
or \g131654/U$5 ( \61251 , \61248 , \50362 );
nand \g131654/U$1 ( \61252 , \61250 , \61251 );
xor \g456111/U$5 ( \61253 , \57443 , \57451 );
and \g456111/U$4 ( \61254 , \61253 , \57456 );
and \g456111/U$6 ( \61255 , \57443 , \57451 );
or \g456111/U$3 ( \61256 , \61254 , \61255 );
xor \g456136/U$1 ( \61257 , \61252 , \61256 );
xor \g131987/U$4 ( \61258 , \57330 , \57338 );
and \g131987/U$3 ( \61259 , \61258 , \57343 );
and \g131987/U$5 ( \61260 , \57330 , \57338 );
or \g131987/U$2 ( \61261 , \61259 , \61260 );
not \g132622/U$3 ( \61262 , \48483 );
and \g132648/U$2 ( \61263 , \54537 , \48479 );
and \g132648/U$3 ( \61264 , \48478 , \54529 );
nor \g132648/U$1 ( \61265 , \61263 , \61264 );
not \g132622/U$4 ( \61266 , \61265 );
or \g132622/U$2 ( \61267 , \61262 , \61266 );
or \g132622/U$5 ( \61268 , \61265 , \48483 );
nand \g132622/U$1 ( \61269 , \61267 , \61268 );
xor \g131882/U$1 ( \61270 , \61261 , \61269 );
and \g132647/U$2 ( \61271 , \48064 , \56167 );
and \g132647/U$3 ( \61272 , \55884 , \48063 );
nor \g132647/U$1 ( \61273 , \61271 , \61272 );
not \g132618/U$3 ( \61274 , \61273 );
not \g132618/U$4 ( \61275 , \47997 );
and \g132618/U$2 ( \61276 , \61274 , \61275 );
and \g132618/U$5 ( \61277 , \61273 , \47997 );
nor \g132618/U$1 ( \61278 , \61276 , \61277 );
not \g131998/U$3 ( \61279 , \61278 );
and \g132543/U$2 ( \61280 , \47930 , \56446 );
and \g132543/U$3 ( \61281 , \56448 , \47931 );
nor \g132543/U$1 ( \61282 , \61280 , \61281 );
not \g132489/U$3 ( \61283 , \61282 );
not \g132489/U$4 ( \61284 , \47935 );
and \g132489/U$2 ( \61285 , \61283 , \61284 );
and \g132489/U$5 ( \61286 , \61282 , \47935 );
nor \g132489/U$1 ( \61287 , \61285 , \61286 );
not \g132023/U$3 ( \61288 , \61287 );
xor \g132059/U$4 ( \61289 , \57205 , \57212 );
and \g132059/U$3 ( \61290 , \61289 , \57224 );
and \g132059/U$5 ( \61291 , \57205 , \57212 );
or \g132059/U$2 ( \61292 , \61290 , \61291 );
not \g132023/U$4 ( \61293 , \61292 );
or \g132023/U$2 ( \61294 , \61288 , \61293 );
or \g132023/U$5 ( \61295 , \61292 , \61287 );
nand \g132023/U$1 ( \61296 , \61294 , \61295 );
not \g131998/U$4 ( \61297 , \61296 );
or \g131998/U$2 ( \61298 , \61279 , \61297 );
or \g131998/U$5 ( \61299 , \61296 , \61278 );
nand \g131998/U$1 ( \61300 , \61298 , \61299 );
xor \g131882/U$1_r1 ( \61301 , \61270 , \61300 );
xor \g456136/U$1_r1 ( \61302 , \61257 , \61301 );
xor \g456100/U$2 ( \61303 , \61244 , \61302 );
not \g131407/U$3 ( \61304 , \51124 );
and \g131451/U$2 ( \61305 , \51117 , \51517 );
and \g131451/U$3 ( \61306 , \51518 , \51098 );
nor \g131451/U$1 ( \61307 , \61305 , \61306 );
not \g131407/U$4 ( \61308 , \61307 );
or \g131407/U$2 ( \61309 , \61304 , \61308 );
or \g131407/U$5 ( \61310 , \61307 , \51124 );
nand \g131407/U$1 ( \61311 , \61309 , \61310 );
not \g132247/U$3 ( \61312 , \49014 );
and \g132298/U$2 ( \61313 , \53848 , \49074 );
and \g132298/U$3 ( \61314 , \49075 , \54015 );
nor \g132298/U$1 ( \61315 , \61313 , \61314 );
not \g132247/U$4 ( \61316 , \61315 );
or \g132247/U$2 ( \61317 , \61312 , \61316 );
or \g132247/U$5 ( \61318 , \61315 , \49014 );
nand \g132247/U$1 ( \61319 , \61317 , \61318 );
not \g132447/U$3 ( \61320 , \48685 );
and \g132495/U$2 ( \61321 , \54185 , \48858 );
and \g132495/U$3 ( \61322 , \48860 , \54251 );
nor \g132495/U$1 ( \61323 , \61321 , \61322 );
not \g132447/U$4 ( \61324 , \61323 );
or \g132447/U$2 ( \61325 , \61320 , \61324 );
or \g132447/U$5 ( \61326 , \61323 , \48685 );
nand \g132447/U$1 ( \61327 , \61325 , \61326 );
xor \g131873/U$1 ( \61328 , \61319 , \61327 );
xor \g131969/U$4 ( \61329 , \57185 , \57193 );
and \g131969/U$3 ( \61330 , \61329 , \57225 );
and \g131969/U$5 ( \61331 , \57185 , \57193 );
or \g131969/U$2 ( \61332 , \61330 , \61331 );
xor \g131873/U$1_r1 ( \61333 , \61328 , \61332 );
xor \g131250/U$1 ( \61334 , \61311 , \61333 );
not \g131292/U$3 ( \61335 , \51120 );
and \g131329/U$2 ( \61336 , \50957 , \52273 );
and \g131329/U$3 ( \61337 , \52270 , \50752 );
nor \g131329/U$1 ( \61338 , \61336 , \61337 );
not \g131292/U$4 ( \61339 , \61338 );
or \g131292/U$2 ( \61340 , \61335 , \61339 );
or \g131292/U$5 ( \61341 , \61338 , \51120 );
nand \g131292/U$1 ( \61342 , \61340 , \61341 );
xor \g131250/U$1_r1 ( \61343 , \61334 , \61342 );
xor \g456100/U$1 ( \61344 , \61303 , \61343 );
xor \g131427/U$4 ( \61345 , \57416 , \57424 );
and \g131427/U$3 ( \61346 , \61345 , \57433 );
and \g131427/U$5 ( \61347 , \57416 , \57424 );
or \g131427/U$2 ( \61348 , \61346 , \61347 );
not \g131919/U$3 ( \61349 , \49568 );
and \g131955/U$2 ( \61350 , \52978 , \49813 );
and \g131955/U$3 ( \61351 , \49812 , \52883 );
nor \g131955/U$1 ( \61352 , \61350 , \61351 );
not \g131919/U$4 ( \61353 , \61352 );
or \g131919/U$2 ( \61354 , \61349 , \61353 );
or \g131919/U$5 ( \61355 , \61352 , \49568 );
nand \g131919/U$1 ( \61356 , \61354 , \61355 );
not \g131782/U$3 ( \61357 , \49925 );
and \g131814/U$2 ( \61358 , \52620 , \50160 );
and \g131814/U$3 ( \61359 , \50159 , \52352 );
nor \g131814/U$1 ( \61360 , \61358 , \61359 );
not \g131782/U$4 ( \61361 , \61360 );
or \g131782/U$2 ( \61362 , \61357 , \61361 );
or \g131782/U$5 ( \61363 , \61360 , \49925 );
nand \g131782/U$1 ( \61364 , \61362 , \61363 );
xor \g456129/U$1 ( \61365 , \61356 , \61364 );
not \g131543/U$3 ( \61366 , \50759 );
and \g131575/U$2 ( \61367 , \51604 , \51055 );
and \g131575/U$3 ( \61368 , \51053 , \51564 );
nor \g131575/U$1 ( \61369 , \61367 , \61368 );
not \g131543/U$4 ( \61370 , \61369 );
or \g131543/U$2 ( \61371 , \61366 , \61370 );
or \g131543/U$5 ( \61372 , \61369 , \50759 );
nand \g131543/U$1 ( \61373 , \61371 , \61372 );
xor \g456129/U$1_r1 ( \61374 , \61365 , \61373 );
xor \g131245/U$1 ( \61375 , \61348 , \61374 );
xor \g456111/U$9 ( \61376 , \57443 , \57451 );
xor \g456111/U$9_r1 ( \61377 , \61376 , \57456 );
and \g456111/U$8 ( \61378 , \57465 , \61377 );
xor \g456111/U$11 ( \61379 , \57443 , \57451 );
xor \g456111/U$11_r1 ( \61380 , \61379 , \57456 );
and \g456111/U$10 ( \61381 , \57473 , \61380 );
and \g456111/U$12 ( \61382 , \57465 , \57473 );
or \g456111/U$7 ( \61383 , \61378 , \61381 , \61382 );
xor \g131245/U$1_r1 ( \61384 , \61375 , \61383 );
xor \g131795/U$4 ( \61385 , \57300 , \57308 );
and \g131795/U$3 ( \61386 , \61385 , \57345 );
and \g131795/U$5 ( \61387 , \57300 , \57308 );
or \g131795/U$2 ( \61388 , \61386 , \61387 );
xor \g456142/U$5 ( \61389 , \57168 , \57176 );
and \g456142/U$4 ( \61390 , \61389 , \57226 );
and \g456142/U$6 ( \61391 , \57168 , \57176 );
or \g456142/U$3 ( \61392 , \61390 , \61391 );
xor \g456106/U$2 ( \61393 , \61388 , \61392 );
not \g132704/U$3 ( \61394 , \48159 );
and \g132754/U$2 ( \61395 , \48154 , \55460 );
and \g132754/U$3 ( \61396 , \55707 , \48155 );
nor \g132754/U$1 ( \61397 , \61395 , \61396 );
not \g132704/U$4 ( \61398 , \61397 );
or \g132704/U$2 ( \61399 , \61394 , \61398 );
or \g132704/U$5 ( \61400 , \61397 , \48159 );
nand \g132704/U$1 ( \61401 , \61399 , \61400 );
not \g132739/U$3 ( \61402 , \48323 );
and \g132779/U$2 ( \61403 , \54853 , \48334 );
and \g132779/U$3 ( \61404 , \55127 , \48335 );
nor \g132779/U$1 ( \61405 , \61403 , \61404 );
not \g132739/U$4 ( \61406 , \61405 );
or \g132739/U$2 ( \61407 , \61402 , \61406 );
or \g132739/U$5 ( \61408 , \61405 , \48323 );
nand \g132739/U$1 ( \61409 , \61407 , \61408 );
xor \g456144/U$2 ( \61410 , \61401 , \61409 );
and \g132165/U$2 ( \61411 , \57215 , \57223 );
and \g132428/U$2 ( \61412 , \47913 , \56357 );
and \g132428/U$3 ( \61413 , \56359 , \47914 );
nor \g132428/U$1 ( \61414 , \61412 , \61413 );
and \g132330/U$2 ( \61415 , \61414 , \47977 );
not \g132330/U$4 ( \61416 , \61414 );
and \g132330/U$3 ( \61417 , \61416 , \47976 );
nor \g132330/U$1 ( \61418 , \61415 , \61417 );
xor \g132060/U$1 ( \61419 , \61411 , \61418 );
not \g135557/U$2 ( \61420 , \56411 );
nor \g135557/U$1 ( \61421 , \61420 , \40060 );
not \g132219/U$3 ( \61422 , \47948 );
and \g132274/U$2 ( \61423 , \47959 , \56347 );
and \g132274/U$3 ( \61424 , \56349 , \47960 );
nor \g132274/U$1 ( \61425 , \61423 , \61424 );
not \g132219/U$4 ( \61426 , \61425 );
or \g132219/U$2 ( \61427 , \61422 , \61426 );
or \g132219/U$5 ( \61428 , \61425 , \47948 );
nand \g132219/U$1 ( \61429 , \61427 , \61428 );
xor \g132166/U$1 ( \61430 , \61421 , \61429 );
xor \g132060/U$1_r1 ( \61431 , \61419 , \61430 );
xor \g456144/U$1 ( \61432 , \61410 , \61431 );
not \g132081/U$3 ( \61433 , \49233 );
and \g132123/U$2 ( \61434 , \53610 , \49405 );
and \g132123/U$3 ( \61435 , \49403 , \53300 );
nor \g132123/U$1 ( \61436 , \61434 , \61435 );
not \g132081/U$4 ( \61437 , \61436 );
or \g132081/U$2 ( \61438 , \61433 , \61437 );
or \g132081/U$5 ( \61439 , \61436 , \49233 );
nand \g132081/U$1 ( \61440 , \61438 , \61439 );
xor \g131874/U$4 ( \61441 , \57313 , \57321 );
and \g131874/U$3 ( \61442 , \61441 , \57344 );
and \g131874/U$5 ( \61443 , \57313 , \57321 );
or \g131874/U$2 ( \61444 , \61442 , \61443 );
xor \g456144/U$1_r1 ( \61445 , \61440 , \61444 );
xor \g456144/U$1_r2 ( \61446 , \61432 , \61445 );
xor \g456106/U$1 ( \61447 , \61393 , \61446 );
xor \g456112/U$5 ( \61448 , \57087 , \57144 );
and \g456112/U$4 ( \61449 , \61448 , \57149 );
and \g456112/U$6 ( \61450 , \57087 , \57144 );
or \g456112/U$3 ( \61451 , \61449 , \61450 );
xor \g131246/U$4 ( \61452 , \57412 , \57434 );
and \g131246/U$3 ( \61453 , \61452 , \57475 );
and \g131246/U$5 ( \61454 , \57412 , \57434 );
or \g131246/U$2 ( \61455 , \61453 , \61454 );
xor \g456106/U$1_r1 ( \61456 , \61451 , \61455 );
xor \g456106/U$1_r2 ( \61457 , \61447 , \61456 );
xor \g456100/U$1_r1 ( \61458 , \61384 , \61457 );
xor \g456100/U$1_r2 ( \61459 , \61344 , \61458 );
xor \g130974/U$1_r1 ( \61460 , \61236 , \61459 );
nand \g128948/U$1 ( \61461 , \61221 , \61460 );
nand \g129062/U$1 ( \61462 , \61215 , \61212 );
nor \g128913/U$1 ( \61463 , \61461 , \61462 );
xor \g456129/U$4 ( \61464 , \61356 , \61364 );
and \g456129/U$3 ( \61465 , \61464 , \61373 );
and \g456129/U$5 ( \61466 , \61356 , \61364 );
nor \g456129/U$2 ( \61467 , \61465 , \61466 );
not \g131255/U$3 ( \61468 , \61467 );
xor \g456136/U$4 ( \61469 , \61252 , \61256 );
and \g456136/U$3 ( \61470 , \61469 , \61301 );
and \g456136/U$5 ( \61471 , \61252 , \61256 );
nor \g456136/U$2 ( \61472 , \61470 , \61471 );
and \g131383/U$2 ( \61473 , \51117 , \51518 );
and \g131383/U$3 ( \61474 , \51517 , \50957 );
nor \g131383/U$1 ( \61475 , \61473 , \61474 );
not \g131350/U$3 ( \61476 , \61475 );
not \g131350/U$4 ( \61477 , \51124 );
and \g131350/U$2 ( \61478 , \61476 , \61477 );
and \g131350/U$5 ( \61479 , \61475 , \51124 );
nor \g131350/U$1 ( \61480 , \61478 , \61479 );
not \g131335/U$3 ( \61481 , \61480 );
and \g131626/U$2 ( \61482 , \51604 , \50587 );
and \g131626/U$3 ( \61483 , \50588 , \51854 );
nor \g131626/U$1 ( \61484 , \61482 , \61483 );
not \g131594/U$3 ( \61485 , \61484 );
not \g131594/U$4 ( \61486 , \50362 );
and \g131594/U$2 ( \61487 , \61485 , \61486 );
and \g131594/U$5 ( \61488 , \61484 , \50362 );
nor \g131594/U$1 ( \61489 , \61487 , \61488 );
and \g132568/U$2 ( \61490 , \54251 , \48478 );
and \g132568/U$3 ( \61491 , \48479 , \54529 );
nor \g132568/U$1 ( \61492 , \61490 , \61491 );
not \g132525/U$3 ( \61493 , \61492 );
not \g132525/U$4 ( \61494 , \48483 );
and \g132525/U$2 ( \61495 , \61493 , \61494 );
and \g132525/U$5 ( \61496 , \61492 , \48483 );
nor \g132525/U$1 ( \61497 , \61495 , \61496 );
not \g132035/U$3 ( \61498 , \61287 );
not \g132035/U$4 ( \61499 , \61278 );
and \g132035/U$2 ( \61500 , \61498 , \61499 );
and \g132038/U$2 ( \61501 , \61287 , \61278 );
not \g132058/U$1 ( \61502 , \61292 );
nor \g132038/U$1 ( \61503 , \61501 , \61502 );
nor \g132035/U$1 ( \61504 , \61500 , \61503 );
xor \g456151/U$1 ( \61505 , \61497 , \61504 );
and \g132414/U$2 ( \61506 , \54185 , \48860 );
and \g132414/U$3 ( \61507 , \48858 , \54015 );
nor \g132414/U$1 ( \61508 , \61506 , \61507 );
not \g132332/U$3 ( \61509 , \61508 );
not \g132332/U$4 ( \61510 , \48685 );
and \g132332/U$2 ( \61511 , \61509 , \61510 );
and \g132332/U$5 ( \61512 , \61508 , \48685 );
nor \g132332/U$1 ( \61513 , \61511 , \61512 );
xor \g456151/U$1_r1 ( \61514 , \61505 , \61513 );
xor \g131568/U$1 ( \61515 , \61489 , \61514 );
not \g131335/U$4 ( \61516 , \61515 );
and \g131335/U$2 ( \61517 , \61481 , \61516 );
and \g131335/U$5 ( \61518 , \61480 , \61515 );
nor \g131335/U$1 ( \61519 , \61517 , \61518 );
xor \g455956/U$1 ( \61520 , \61472 , \61519 );
not \g131255/U$4 ( \61521 , \61520 );
or \g131255/U$2 ( \61522 , \61468 , \61521 );
or \g131255/U$5 ( \61523 , \61520 , \61467 );
nand \g131255/U$1 ( \61524 , \61522 , \61523 );
xor \g131245/U$4 ( \61525 , \61348 , \61374 );
and \g131245/U$3 ( \61526 , \61525 , \61383 );
and \g131245/U$5 ( \61527 , \61348 , \61374 );
or \g131245/U$2 ( \61528 , \61526 , \61527 );
xor \g131120/U$1 ( \61529 , \61524 , \61528 );
and \g132041/U$2 ( \61530 , \52978 , \49403 );
and \g132041/U$3 ( \61531 , \49405 , \53300 );
nor \g132041/U$1 ( \61532 , \61530 , \61531 );
not \g132002/U$3 ( \61533 , \61532 );
not \g132002/U$4 ( \61534 , \49233 );
and \g132002/U$2 ( \61535 , \61533 , \61534 );
and \g132002/U$5 ( \61536 , \61532 , \49233 );
nor \g132002/U$1 ( \61537 , \61535 , \61536 );
not \g131808/U$3 ( \61538 , \61537 );
and \g132752/U$2 ( \61539 , \48154 , \55127 );
and \g132752/U$3 ( \61540 , \55460 , \48155 );
nor \g132752/U$1 ( \61541 , \61539 , \61540 );
not \g132703/U$3 ( \61542 , \61541 );
not \g132703/U$4 ( \61543 , \48159 );
and \g132703/U$2 ( \61544 , \61542 , \61543 );
and \g132703/U$5 ( \61545 , \61541 , \48159 );
nor \g132703/U$1 ( \61546 , \61544 , \61545 );
not \g132025/U$3 ( \61547 , \61546 );
and \g132166/U$2 ( \61548 , \61421 , \61429 );
and \g132411/U$2 ( \61549 , \47914 , \56357 );
and \g132411/U$3 ( \61550 , \56448 , \47913 );
nor \g132411/U$1 ( \61551 , \61549 , \61550 );
and \g132347/U$2 ( \61552 , \61551 , \47977 );
not \g132347/U$4 ( \61553 , \61551 );
and \g132347/U$3 ( \61554 , \61553 , \47976 );
nor \g132347/U$1 ( \61555 , \61552 , \61554 );
xor \g132066/U$1 ( \61556 , \61548 , \61555 );
not \g135556/U$2 ( \61557 , \56349 );
nor \g135556/U$1 ( \61558 , \61557 , \40060 );
not \g132218/U$3 ( \61559 , \47948 );
and \g132273/U$2 ( \61560 , \47960 , \56347 );
and \g132273/U$3 ( \61561 , \56359 , \47959 );
nor \g132273/U$1 ( \61562 , \61560 , \61561 );
not \g132218/U$4 ( \61563 , \61562 );
or \g132218/U$2 ( \61564 , \61559 , \61563 );
or \g132218/U$5 ( \61565 , \61562 , \47948 );
nand \g132218/U$1 ( \61566 , \61564 , \61565 );
xor \g132163/U$1 ( \61567 , \61558 , \61566 );
xor \g132066/U$1_r1 ( \61568 , \61556 , \61567 );
not \g132025/U$4 ( \61569 , \61568 );
or \g132025/U$2 ( \61570 , \61547 , \61569 );
or \g132025/U$5 ( \61571 , \61568 , \61546 );
nand \g132025/U$1 ( \61572 , \61570 , \61571 );
not \g131997/U$3 ( \61573 , \61572 );
and \g132720/U$2 ( \61574 , \48335 , \54853 );
and \g132720/U$3 ( \61575 , \48334 , \54537 );
nor \g132720/U$1 ( \61576 , \61574 , \61575 );
not \g132676/U$3 ( \61577 , \61576 );
not \g132676/U$4 ( \61578 , \48323 );
and \g132676/U$2 ( \61579 , \61577 , \61578 );
and \g132676/U$5 ( \61580 , \61576 , \48323 );
nor \g132676/U$1 ( \61581 , \61579 , \61580 );
not \g131997/U$4 ( \61582 , \61581 );
and \g131997/U$2 ( \61583 , \61573 , \61582 );
and \g131997/U$5 ( \61584 , \61572 , \61581 );
nor \g131997/U$1 ( \61585 , \61583 , \61584 );
not \g131835/U$3 ( \61586 , \61585 );
xor \g131882/U$4 ( \61587 , \61261 , \61269 );
and \g131882/U$3 ( \61588 , \61587 , \61300 );
and \g131882/U$5 ( \61589 , \61261 , \61269 );
or \g131882/U$2 ( \61590 , \61588 , \61589 );
not \g131835/U$4 ( \61591 , \61590 );
or \g131835/U$2 ( \61592 , \61586 , \61591 );
or \g131835/U$5 ( \61593 , \61590 , \61585 );
nand \g131835/U$1 ( \61594 , \61592 , \61593 );
not \g131808/U$4 ( \61595 , \61594 );
or \g131808/U$2 ( \61596 , \61538 , \61595 );
or \g131808/U$5 ( \61597 , \61594 , \61537 );
nand \g131808/U$1 ( \61598 , \61596 , \61597 );
not \g131847/U$3 ( \61599 , \49568 );
and \g131896/U$2 ( \61600 , \52620 , \49812 );
and \g131896/U$3 ( \61601 , \49813 , \52883 );
nor \g131896/U$1 ( \61602 , \61600 , \61601 );
not \g131847/U$4 ( \61603 , \61602 );
or \g131847/U$2 ( \61604 , \61599 , \61603 );
or \g131847/U$5 ( \61605 , \61602 , \49568 );
nand \g131847/U$1 ( \61606 , \61604 , \61605 );
not \g131722/U$3 ( \61607 , \49925 );
and \g131755/U$2 ( \61608 , \52108 , \50159 );
and \g131755/U$3 ( \61609 , \50160 , \52352 );
nor \g131755/U$1 ( \61610 , \61608 , \61609 );
not \g131722/U$4 ( \61611 , \61610 );
or \g131722/U$2 ( \61612 , \61607 , \61611 );
or \g131722/U$5 ( \61613 , \61610 , \49925 );
nand \g131722/U$1 ( \61614 , \61612 , \61613 );
xor \g456123/U$1 ( \61615 , \61606 , \61614 );
not \g131477/U$3 ( \61616 , \50759 );
and \g131507/U$2 ( \61617 , \51564 , \51055 );
and \g131507/U$3 ( \61618 , \51053 , \51098 );
nor \g131507/U$1 ( \61619 , \61617 , \61618 );
not \g131477/U$4 ( \61620 , \61619 );
or \g131477/U$2 ( \61621 , \61616 , \61620 );
or \g131477/U$5 ( \61622 , \61619 , \50759 );
nand \g131477/U$1 ( \61623 , \61621 , \61622 );
xor \g456123/U$1_r1 ( \61624 , \61615 , \61623 );
xor \g131198/U$1 ( \61625 , \61598 , \61624 );
not \g131231/U$3 ( \61626 , \51120 );
and \g131276/U$2 ( \61627 , \50752 , \52273 );
and \g131276/U$3 ( \61628 , \52270 , \50443 );
nor \g131276/U$1 ( \61629 , \61627 , \61628 );
not \g131231/U$4 ( \61630 , \61629 );
or \g131231/U$2 ( \61631 , \61626 , \61630 );
or \g131231/U$5 ( \61632 , \61629 , \51120 );
nand \g131231/U$1 ( \61633 , \61631 , \61632 );
xor \g131198/U$1_r1 ( \61634 , \61625 , \61633 );
xor \g131120/U$1_r1 ( \61635 , \61529 , \61634 );
xor \g456100/U$9 ( \61636 , \61244 , \61302 );
xor \g456100/U$9_r1 ( \61637 , \61636 , \61343 );
and \g456100/U$8 ( \61638 , \61384 , \61637 );
xor \g456100/U$11 ( \61639 , \61244 , \61302 );
xor \g456100/U$11_r1 ( \61640 , \61639 , \61343 );
and \g456100/U$10 ( \61641 , \61457 , \61640 );
and \g456100/U$12 ( \61642 , \61384 , \61457 );
or \g456100/U$7 ( \61643 , \61638 , \61641 , \61642 );
xor \g456097/U$1 ( \61644 , \61635 , \61643 );
xor \g456106/U$9 ( \61645 , \61388 , \61392 );
xor \g456106/U$9_r1 ( \61646 , \61645 , \61446 );
and \g456106/U$8 ( \61647 , \61451 , \61646 );
xor \g456106/U$11 ( \61648 , \61388 , \61392 );
xor \g456106/U$11_r1 ( \61649 , \61648 , \61446 );
and \g456106/U$10 ( \61650 , \61455 , \61649 );
and \g456106/U$12 ( \61651 , \61451 , \61455 );
or \g456106/U$7 ( \61652 , \61647 , \61650 , \61651 );
xor \g456100/U$5 ( \61653 , \61244 , \61302 );
and \g456100/U$4 ( \61654 , \61653 , \61343 );
and \g456100/U$6 ( \61655 , \61244 , \61302 );
or \g456100/U$3 ( \61656 , \61654 , \61655 );
xor \g131075/U$1 ( \61657 , \61652 , \61656 );
xor \g456106/U$5 ( \61658 , \61388 , \61392 );
and \g456106/U$4 ( \61659 , \61658 , \61446 );
and \g456106/U$6 ( \61660 , \61388 , \61392 );
or \g456106/U$3 ( \61661 , \61659 , \61660 );
xor \g456144/U$5 ( \61662 , \61401 , \61409 );
and \g456144/U$4 ( \61663 , \61662 , \61431 );
and \g456144/U$6 ( \61664 , \61401 , \61409 );
or \g456144/U$3 ( \61665 , \61663 , \61664 );
not \g132159/U$3 ( \61666 , \49014 );
and \g132194/U$2 ( \61667 , \53610 , \49074 );
and \g132194/U$3 ( \61668 , \49075 , \53848 );
nor \g132194/U$1 ( \61669 , \61667 , \61668 );
not \g132159/U$4 ( \61670 , \61669 );
or \g132159/U$2 ( \61671 , \61666 , \61670 );
or \g132159/U$5 ( \61672 , \61669 , \49014 );
nand \g132159/U$1 ( \61673 , \61671 , \61672 );
xor \g456141/U$2 ( \61674 , \61665 , \61673 );
not \g132477/U$3 ( \61675 , \47935 );
and \g132542/U$2 ( \61676 , \47931 , \56446 );
and \g132542/U$3 ( \61677 , \56167 , \47930 );
nor \g132542/U$1 ( \61678 , \61676 , \61677 );
not \g132477/U$4 ( \61679 , \61678 );
or \g132477/U$2 ( \61680 , \61675 , \61679 );
or \g132477/U$5 ( \61681 , \61678 , \47935 );
nand \g132477/U$1 ( \61682 , \61680 , \61681 );
not \g132598/U$3 ( \61683 , \47997 );
and \g132645/U$2 ( \61684 , \48064 , \55884 );
and \g132645/U$3 ( \61685 , \55707 , \48063 );
nor \g132645/U$1 ( \61686 , \61684 , \61685 );
not \g132598/U$4 ( \61687 , \61686 );
or \g132598/U$2 ( \61688 , \61683 , \61687 );
or \g132598/U$5 ( \61689 , \61686 , \47997 );
nand \g132598/U$1 ( \61690 , \61688 , \61689 );
xor \g131977/U$1 ( \61691 , \61682 , \61690 );
xor \g132060/U$4 ( \61692 , \61411 , \61418 );
and \g132060/U$3 ( \61693 , \61692 , \61430 );
and \g132060/U$5 ( \61694 , \61411 , \61418 );
or \g132060/U$2 ( \61695 , \61693 , \61694 );
xor \g131977/U$1_r1 ( \61696 , \61691 , \61695 );
xor \g456141/U$1 ( \61697 , \61674 , \61696 );
xor \g131873/U$4 ( \61698 , \61319 , \61327 );
and \g131873/U$3 ( \61699 , \61698 , \61332 );
and \g131873/U$5 ( \61700 , \61319 , \61327 );
or \g131873/U$2 ( \61701 , \61699 , \61700 );
xor \g456144/U$9 ( \61702 , \61401 , \61409 );
xor \g456144/U$9_r1 ( \61703 , \61702 , \61431 );
and \g456144/U$8 ( \61704 , \61440 , \61703 );
xor \g456144/U$11 ( \61705 , \61401 , \61409 );
xor \g456144/U$11_r1 ( \61706 , \61705 , \61431 );
and \g456144/U$10 ( \61707 , \61444 , \61706 );
and \g456144/U$12 ( \61708 , \61440 , \61444 );
or \g456144/U$7 ( \61709 , \61704 , \61707 , \61708 );
xor \g456141/U$1_r1 ( \61710 , \61701 , \61709 );
xor \g456141/U$1_r2 ( \61711 , \61697 , \61710 );
xor \g131192/U$1 ( \61712 , \61661 , \61711 );
xor \g131250/U$4 ( \61713 , \61311 , \61333 );
and \g131250/U$3 ( \61714 , \61713 , \61342 );
and \g131250/U$5 ( \61715 , \61311 , \61333 );
or \g131250/U$2 ( \61716 , \61714 , \61715 );
xor \g131192/U$1_r1 ( \61717 , \61712 , \61716 );
xor \g131075/U$1_r1 ( \61718 , \61657 , \61717 );
xor \g456097/U$1_r1 ( \61719 , \61644 , \61718 );
xor \g130974/U$4 ( \61720 , \61227 , \61235 );
and \g130974/U$3 ( \61721 , \61720 , \61459 );
and \g130974/U$5 ( \61722 , \61227 , \61235 );
or \g130974/U$2 ( \61723 , \61721 , \61722 );
not \g128882/U$3 ( \61724 , \61462 );
or \g128914/U$2 ( \61725 , \61219 , \57492 );
nand \g128914/U$1 ( \61726 , \61725 , \61461 );
not \g128882/U$4 ( \61727 , \61726 );
or \g128882/U$2 ( \61728 , \61724 , \61727 );
or \g128882/U$5 ( \61729 , \61726 , \61462 );
nand \g128882/U$1 ( \61730 , \61728 , \61729 );
xor \g128854/U$1 ( \61731 , \61723 , \61730 );
and \g128830/U$2 ( \61732 , \61719 , \61731 );
nand \g128821/U$1 ( \61733 , \61463 , \61732 );
not \g128814/U$3 ( \61734 , \61733 );
and \g128822/U$2 ( \61735 , \61730 , \61723 );
nor \g128822/U$1 ( \61736 , \61735 , \61732 );
not \g128820/U$3 ( \61737 , \61736 );
not \g128820/U$4 ( \61738 , \61463 );
and \g128820/U$2 ( \61739 , \61737 , \61738 );
and \g128820/U$5 ( \61740 , \61736 , \61463 );
nor \g128820/U$1 ( \61741 , \61739 , \61740 );
xor \g456097/U$4 ( \61742 , \61635 , \61643 );
and \g456097/U$3 ( \61743 , \61742 , \61718 );
and \g456097/U$5 ( \61744 , \61635 , \61643 );
nor \g456097/U$2 ( \61745 , \61743 , \61744 );
or \g128816/U$2 ( \61746 , \61741 , \61745 );
xnor \g128819/U$1 ( \61747 , \61745 , \61741 );
not \g128818/U$2 ( \61748 , \61747 );
xor \g131075/U$4 ( \61749 , \61652 , \61656 );
and \g131075/U$3 ( \61750 , \61749 , \61717 );
and \g131075/U$5 ( \61751 , \61652 , \61656 );
or \g131075/U$2 ( \61752 , \61750 , \61751 );
and \g131819/U$2 ( \61753 , \52620 , \49813 );
and \g131819/U$3 ( \61754 , \49812 , \52352 );
nor \g131819/U$1 ( \61755 , \61753 , \61754 );
not \g131781/U$3 ( \61756 , \61755 );
not \g131781/U$4 ( \61757 , \49568 );
and \g131781/U$2 ( \61758 , \61756 , \61757 );
and \g131781/U$5 ( \61759 , \61755 , \49568 );
nor \g131781/U$1 ( \61760 , \61758 , \61759 );
and \g131956/U$2 ( \61761 , \52978 , \49405 );
and \g131956/U$3 ( \61762 , \49403 , \52883 );
nor \g131956/U$1 ( \61763 , \61761 , \61762 );
not \g131918/U$3 ( \61764 , \61763 );
not \g131918/U$4 ( \61765 , \49233 );
and \g131918/U$2 ( \61766 , \61764 , \61765 );
and \g131918/U$5 ( \61767 , \61763 , \49233 );
nor \g131918/U$1 ( \61768 , \61766 , \61767 );
xor \g456114/U$2 ( \61769 , \61760 , \61768 );
and \g132163/U$2 ( \61770 , \61558 , \61566 );
not \g132117/U$3 ( \61771 , \61770 );
not \g132217/U$3 ( \61772 , \47948 );
and \g132271/U$2 ( \61773 , \47959 , \56357 );
and \g132271/U$3 ( \61774 , \56359 , \47960 );
nor \g132271/U$1 ( \61775 , \61773 , \61774 );
not \g132217/U$4 ( \61776 , \61775 );
or \g132217/U$2 ( \61777 , \61772 , \61776 );
or \g132217/U$5 ( \61778 , \61775 , \47948 );
nand \g132217/U$1 ( \61779 , \61777 , \61778 );
not \g132180/U$3 ( \61780 , \61779 );
nand \g132368/U$1 ( \61781 , \56347 , \40061 );
not \g132180/U$4 ( \61782 , \61781 );
and \g132180/U$2 ( \61783 , \61780 , \61782 );
and \g132180/U$5 ( \61784 , \61779 , \61781 );
nor \g132180/U$1 ( \61785 , \61783 , \61784 );
not \g132117/U$4 ( \61786 , \61785 );
or \g132117/U$2 ( \61787 , \61771 , \61786 );
or \g132117/U$5 ( \61788 , \61785 , \61770 );
nand \g132117/U$1 ( \61789 , \61787 , \61788 );
not \g132100/U$3 ( \61790 , \61789 );
and \g132409/U$2 ( \61791 , \47913 , \56446 );
and \g132409/U$3 ( \61792 , \56448 , \47914 );
nor \g132409/U$1 ( \61793 , \61791 , \61792 );
and \g132327/U$2 ( \61794 , \61793 , \47976 );
not \g132327/U$4 ( \61795 , \61793 );
and \g132327/U$3 ( \61796 , \61795 , \47977 );
nor \g132327/U$1 ( \61797 , \61794 , \61796 );
not \g132100/U$4 ( \61798 , \61797 );
and \g132100/U$2 ( \61799 , \61790 , \61798 );
and \g132100/U$5 ( \61800 , \61789 , \61797 );
nor \g132100/U$1 ( \61801 , \61799 , \61800 );
not \g131922/U$3 ( \61802 , \61801 );
xor \g131977/U$4 ( \61803 , \61682 , \61690 );
and \g131977/U$3 ( \61804 , \61803 , \61695 );
and \g131977/U$5 ( \61805 , \61682 , \61690 );
or \g131977/U$2 ( \61806 , \61804 , \61805 );
not \g131922/U$4 ( \61807 , \61806 );
or \g131922/U$2 ( \61808 , \61802 , \61807 );
or \g131922/U$5 ( \61809 , \61806 , \61801 );
nand \g131922/U$1 ( \61810 , \61808 , \61809 );
not \g131907/U$3 ( \61811 , \61810 );
and \g132644/U$2 ( \61812 , \48063 , \55460 );
and \g132644/U$3 ( \61813 , \55707 , \48064 );
nor \g132644/U$1 ( \61814 , \61812 , \61813 );
not \g132597/U$3 ( \61815 , \61814 );
not \g132597/U$4 ( \61816 , \47997 );
and \g132597/U$2 ( \61817 , \61815 , \61816 );
and \g132597/U$5 ( \61818 , \61814 , \47997 );
nor \g132597/U$1 ( \61819 , \61817 , \61818 );
not \g131907/U$4 ( \61820 , \61819 );
and \g131907/U$2 ( \61821 , \61811 , \61820 );
and \g131907/U$5 ( \61822 , \61810 , \61819 );
nor \g131907/U$1 ( \61823 , \61821 , \61822 );
xor \g456114/U$1 ( \61824 , \61769 , \61823 );
not \g131841/U$3 ( \61825 , \61585 );
not \g131841/U$4 ( \61826 , \61537 );
and \g131841/U$2 ( \61827 , \61825 , \61826 );
and \g131843/U$2 ( \61828 , \61585 , \61537 );
not \g131881/U$1 ( \61829 , \61590 );
nor \g131843/U$1 ( \61830 , \61828 , \61829 );
nor \g131841/U$1 ( \61831 , \61827 , \61830 );
xor \g456123/U$4 ( \61832 , \61606 , \61614 );
and \g456123/U$3 ( \61833 , \61832 , \61623 );
and \g456123/U$5 ( \61834 , \61606 , \61614 );
nor \g456123/U$2 ( \61835 , \61833 , \61834 );
xor \g456114/U$1_r1 ( \61836 , \61831 , \61835 );
xor \g456114/U$1_r2 ( \61837 , \61824 , \61836 );
not \g131116/U$3 ( \61838 , \61837 );
not \g131286/U$3 ( \61839 , \61472 );
not \g131286/U$4 ( \61840 , \61467 );
and \g131286/U$2 ( \61841 , \61839 , \61840 );
and \g131287/U$2 ( \61842 , \61472 , \61467 );
nor \g131287/U$1 ( \61843 , \61842 , \61519 );
nor \g131286/U$1 ( \61844 , \61841 , \61843 );
not \g131132/U$3 ( \61845 , \61844 );
xor \g131192/U$4 ( \61846 , \61661 , \61711 );
and \g131192/U$3 ( \61847 , \61846 , \61716 );
and \g131192/U$5 ( \61848 , \61661 , \61711 );
or \g131192/U$2 ( \61849 , \61847 , \61848 );
not \g131132/U$4 ( \61850 , \61849 );
or \g131132/U$2 ( \61851 , \61845 , \61850 );
or \g131132/U$5 ( \61852 , \61849 , \61844 );
nand \g131132/U$1 ( \61853 , \61851 , \61852 );
not \g131116/U$4 ( \61854 , \61853 );
or \g131116/U$2 ( \61855 , \61838 , \61854 );
or \g131116/U$5 ( \61856 , \61853 , \61837 );
nand \g131116/U$1 ( \61857 , \61855 , \61856 );
xor \g130910/U$1 ( \61858 , \61752 , \61857 );
xor \g456141/U$9 ( \61859 , \61665 , \61673 );
xor \g456141/U$9_r1 ( \61860 , \61859 , \61696 );
and \g456141/U$8 ( \61861 , \61701 , \61860 );
xor \g456141/U$11 ( \61862 , \61665 , \61673 );
xor \g456141/U$11_r1 ( \61863 , \61862 , \61696 );
and \g456141/U$10 ( \61864 , \61709 , \61863 );
and \g456141/U$12 ( \61865 , \61701 , \61709 );
or \g456141/U$7 ( \61866 , \61861 , \61864 , \61865 );
xor \g456151/U$4 ( \61867 , \61497 , \61504 );
and \g456151/U$3 ( \61868 , \61867 , \61513 );
and \g456151/U$5 ( \61869 , \61497 , \61504 );
nor \g456151/U$2 ( \61870 , \61868 , \61869 );
not \g131651/U$3 ( \61871 , \49925 );
and \g131687/U$2 ( \61872 , \52108 , \50160 );
and \g131687/U$3 ( \61873 , \50159 , \51854 );
nor \g131687/U$1 ( \61874 , \61872 , \61873 );
not \g131651/U$4 ( \61875 , \61874 );
or \g131651/U$2 ( \61876 , \61871 , \61875 );
or \g131651/U$5 ( \61877 , \61874 , \49925 );
nand \g131651/U$1 ( \61878 , \61876 , \61877 );
xor \g131495/U$1 ( \61879 , \61870 , \61878 );
not \g131542/U$3 ( \61880 , \50362 );
and \g131574/U$2 ( \61881 , \51604 , \50588 );
and \g131574/U$3 ( \61882 , \50587 , \51564 );
nor \g131574/U$1 ( \61883 , \61881 , \61882 );
not \g131542/U$4 ( \61884 , \61883 );
or \g131542/U$2 ( \61885 , \61880 , \61884 );
or \g131542/U$5 ( \61886 , \61883 , \50362 );
nand \g131542/U$1 ( \61887 , \61885 , \61886 );
xor \g131495/U$1_r1 ( \61888 , \61879 , \61887 );
xor \g131244/U$1 ( \61889 , \61866 , \61888 );
or \g131333/U$2 ( \61890 , \61514 , \61489 );
and \g131341/U$2 ( \61891 , \61514 , \61489 );
nor \g131341/U$1 ( \61892 , \61891 , \61480 );
not \g131340/U$1 ( \61893 , \61892 );
nand \g131333/U$1 ( \61894 , \61890 , \61893 );
xor \g131244/U$1_r1 ( \61895 , \61889 , \61894 );
xor \g131120/U$4 ( \61896 , \61524 , \61528 );
and \g131120/U$3 ( \61897 , \61896 , \61634 );
and \g131120/U$5 ( \61898 , \61524 , \61528 );
or \g131120/U$2 ( \61899 , \61897 , \61898 );
xor \g456096/U$1 ( \61900 , \61895 , \61899 );
xor \g456141/U$5 ( \61901 , \61665 , \61673 );
and \g456141/U$4 ( \61902 , \61901 , \61696 );
and \g456141/U$6 ( \61903 , \61665 , \61673 );
or \g456141/U$3 ( \61904 , \61902 , \61903 );
not \g132080/U$3 ( \61905 , \49014 );
and \g132122/U$2 ( \61906 , \53610 , \49075 );
and \g132122/U$3 ( \61907 , \49074 , \53300 );
nor \g132122/U$1 ( \61908 , \61906 , \61907 );
not \g132080/U$4 ( \61909 , \61908 );
or \g132080/U$2 ( \61910 , \61905 , \61909 );
or \g132080/U$5 ( \61911 , \61908 , \49014 );
nand \g132080/U$1 ( \61912 , \61910 , \61911 );
not \g132246/U$3 ( \61913 , \48685 );
and \g132296/U$2 ( \61914 , \53848 , \48858 );
and \g132296/U$3 ( \61915 , \48860 , \54015 );
nor \g132296/U$1 ( \61916 , \61914 , \61915 );
not \g132246/U$4 ( \61917 , \61916 );
or \g132246/U$2 ( \61918 , \61913 , \61917 );
or \g132246/U$5 ( \61919 , \61916 , \48685 );
nand \g132246/U$1 ( \61920 , \61918 , \61919 );
xor \g131883/U$1 ( \61921 , \61912 , \61920 );
and \g132755/U$2 ( \61922 , \48154 , \54853 );
and \g132755/U$3 ( \61923 , \55127 , \48155 );
nor \g132755/U$1 ( \61924 , \61922 , \61923 );
not \g132702/U$3 ( \61925 , \61924 );
not \g132702/U$4 ( \61926 , \48159 );
and \g132702/U$2 ( \61927 , \61925 , \61926 );
and \g132702/U$5 ( \61928 , \61924 , \48159 );
nor \g132702/U$1 ( \61929 , \61927 , \61928 );
not \g131996/U$3 ( \61930 , \61929 );
and \g132541/U$2 ( \61931 , \47931 , \56167 );
and \g132541/U$3 ( \61932 , \55884 , \47930 );
nor \g132541/U$1 ( \61933 , \61931 , \61932 );
not \g132476/U$3 ( \61934 , \61933 );
not \g132476/U$4 ( \61935 , \47935 );
and \g132476/U$2 ( \61936 , \61934 , \61935 );
and \g132476/U$5 ( \61937 , \61933 , \47935 );
nor \g132476/U$1 ( \61938 , \61936 , \61937 );
not \g132022/U$3 ( \61939 , \61938 );
xor \g132066/U$4 ( \61940 , \61548 , \61555 );
and \g132066/U$3 ( \61941 , \61940 , \61567 );
and \g132066/U$5 ( \61942 , \61548 , \61555 );
or \g132066/U$2 ( \61943 , \61941 , \61942 );
not \g132022/U$4 ( \61944 , \61943 );
or \g132022/U$2 ( \61945 , \61939 , \61944 );
or \g132022/U$5 ( \61946 , \61943 , \61938 );
nand \g132022/U$1 ( \61947 , \61945 , \61946 );
not \g131996/U$4 ( \61948 , \61947 );
or \g131996/U$2 ( \61949 , \61930 , \61948 );
or \g131996/U$5 ( \61950 , \61947 , \61929 );
nand \g131996/U$1 ( \61951 , \61949 , \61950 );
xor \g131883/U$1_r1 ( \61952 , \61921 , \61951 );
xor \g456119/U$1 ( \61953 , \61904 , \61952 );
not \g131406/U$3 ( \61954 , \50759 );
and \g131441/U$2 ( \61955 , \51117 , \51053 );
and \g131441/U$3 ( \61956 , \51055 , \51098 );
nor \g131441/U$1 ( \61957 , \61955 , \61956 );
not \g131406/U$4 ( \61958 , \61957 );
or \g131406/U$2 ( \61959 , \61954 , \61958 );
or \g131406/U$5 ( \61960 , \61957 , \50759 );
nand \g131406/U$1 ( \61961 , \61959 , \61960 );
xor \g456119/U$1_r1 ( \61962 , \61953 , \61961 );
not \g132448/U$3 ( \61963 , \48483 );
and \g132494/U$2 ( \61964 , \54185 , \48478 );
and \g132494/U$3 ( \61965 , \48479 , \54251 );
nor \g132494/U$1 ( \61966 , \61964 , \61965 );
not \g132448/U$4 ( \61967 , \61966 );
or \g132448/U$2 ( \61968 , \61963 , \61967 );
or \g132448/U$5 ( \61969 , \61966 , \48483 );
nand \g132448/U$1 ( \61970 , \61968 , \61969 );
not \g132599/U$3 ( \61971 , \48323 );
and \g132646/U$2 ( \61972 , \48335 , \54537 );
and \g132646/U$3 ( \61973 , \48334 , \54529 );
nor \g132646/U$1 ( \61974 , \61972 , \61973 );
not \g132599/U$4 ( \61975 , \61974 );
or \g132599/U$2 ( \61976 , \61971 , \61975 );
or \g132599/U$5 ( \61977 , \61974 , \48323 );
nand \g132599/U$1 ( \61978 , \61976 , \61977 );
xor \g131871/U$1 ( \61979 , \61970 , \61978 );
or \g132034/U$2 ( \61980 , \61546 , \61581 );
not \g132037/U$3 ( \61981 , \61581 );
not \g132037/U$4 ( \61982 , \61546 );
or \g132037/U$2 ( \61983 , \61981 , \61982 );
nand \g132037/U$1 ( \61984 , \61983 , \61568 );
nand \g132034/U$1 ( \61985 , \61980 , \61984 );
xor \g131871/U$1_r1 ( \61986 , \61979 , \61985 );
not \g131291/U$3 ( \61987 , \51124 );
and \g131328/U$2 ( \61988 , \50957 , \51518 );
and \g131328/U$3 ( \61989 , \51517 , \50752 );
nor \g131328/U$1 ( \61990 , \61988 , \61989 );
not \g131291/U$4 ( \61991 , \61990 );
or \g131291/U$2 ( \61992 , \61987 , \61991 );
or \g131291/U$5 ( \61993 , \61990 , \51124 );
nand \g131291/U$1 ( \61994 , \61992 , \61993 );
xor \g456102/U$1 ( \61995 , \61986 , \61994 );
not \g131178/U$3 ( \61996 , \51120 );
and \g131221/U$2 ( \61997 , \50305 , \52270 );
and \g131221/U$3 ( \61998 , \52273 , \50443 );
nor \g131221/U$1 ( \61999 , \61997 , \61998 );
not \g131178/U$4 ( \62000 , \61999 );
or \g131178/U$2 ( \62001 , \61996 , \62000 );
or \g131178/U$5 ( \62002 , \61999 , \51120 );
nand \g131178/U$1 ( \62003 , \62001 , \62002 );
xor \g456102/U$1_r1 ( \62004 , \61995 , \62003 );
xor \g456099/U$1 ( \62005 , \61962 , \62004 );
xor \g131198/U$4 ( \62006 , \61598 , \61624 );
and \g131198/U$3 ( \62007 , \62006 , \61633 );
and \g131198/U$5 ( \62008 , \61598 , \61624 );
or \g131198/U$2 ( \62009 , \62007 , \62008 );
xor \g456099/U$1_r1 ( \62010 , \62005 , \62009 );
xor \g456096/U$1_r1 ( \62011 , \61900 , \62010 );
xor \g130910/U$1_r1 ( \62012 , \61858 , \62011 );
nand \g128818/U$1 ( \62013 , \61748 , \62012 );
nand \g128816/U$1 ( \62014 , \61746 , \62013 );
not \g128814/U$4 ( \62015 , \62014 );
or \g128814/U$2 ( \62016 , \61734 , \62015 );
or \g128814/U$5 ( \62017 , \62014 , \61733 );
nand \g128814/U$1 ( \62018 , \62016 , \62017 );
xor \g130910/U$4 ( \62019 , \61752 , \61857 );
and \g130910/U$3 ( \62020 , \62019 , \62011 );
and \g130910/U$5 ( \62021 , \61752 , \61857 );
or \g130910/U$2 ( \62022 , \62020 , \62021 );
and \g128809/U$2 ( \62023 , \62018 , \62022 );
not \g131152/U$3 ( \62024 , \61844 );
not \g131152/U$4 ( \62025 , \61837 );
and \g131152/U$2 ( \62026 , \62024 , \62025 );
and \g131167/U$2 ( \62027 , \61844 , \61837 );
not \g131191/U$1 ( \62028 , \61849 );
nor \g131167/U$1 ( \62029 , \62027 , \62028 );
nor \g131152/U$1 ( \62030 , \62026 , \62029 );
xor \g456114/U$9 ( \62031 , \61760 , \61768 );
xor \g456114/U$9_r1 ( \62032 , \62031 , \61823 );
and \g456114/U$8 ( \62033 , \61831 , \62032 );
xor \g456114/U$11 ( \62034 , \61760 , \61768 );
xor \g456114/U$11_r1 ( \62035 , \62034 , \61823 );
and \g456114/U$10 ( \62036 , \61835 , \62035 );
and \g456114/U$12 ( \62037 , \61831 , \61835 );
or \g456114/U$7 ( \62038 , \62033 , \62036 , \62037 );
xor \g456119/U$4 ( \62039 , \61904 , \61952 );
and \g456119/U$3 ( \62040 , \62039 , \61961 );
and \g456119/U$5 ( \62041 , \61904 , \61952 );
nor \g456119/U$2 ( \62042 , \62040 , \62041 );
xor \g131247/U$1 ( \62043 , \62038 , \62042 );
and \g131372/U$2 ( \62044 , \51117 , \51055 );
and \g131372/U$3 ( \62045 , \51053 , \50957 );
nor \g131372/U$1 ( \62046 , \62044 , \62045 );
not \g131349/U$3 ( \62047 , \62046 );
not \g131349/U$4 ( \62048 , \50759 );
and \g131349/U$2 ( \62049 , \62047 , \62048 );
and \g131349/U$5 ( \62050 , \62046 , \50759 );
nor \g131349/U$1 ( \62051 , \62049 , \62050 );
not \g131334/U$3 ( \62052 , \62051 );
and \g132410/U$2 ( \62053 , \54185 , \48479 );
and \g132410/U$3 ( \62054 , \48478 , \54015 );
nor \g132410/U$1 ( \62055 , \62053 , \62054 );
not \g132329/U$3 ( \62056 , \62055 );
not \g132329/U$4 ( \62057 , \48483 );
and \g132329/U$2 ( \62058 , \62056 , \62057 );
and \g132329/U$5 ( \62059 , \62055 , \48483 );
nor \g132329/U$1 ( \62060 , \62058 , \62059 );
not \g132033/U$3 ( \62061 , \61938 );
not \g132033/U$4 ( \62062 , \61929 );
and \g132033/U$2 ( \62063 , \62061 , \62062 );
and \g132036/U$2 ( \62064 , \61938 , \61929 );
not \g132065/U$1 ( \62065 , \61943 );
nor \g132036/U$1 ( \62066 , \62064 , \62065 );
nor \g132033/U$1 ( \62067 , \62063 , \62066 );
xor \g456150/U$1 ( \62068 , \62060 , \62067 );
and \g132046/U$2 ( \62069 , \52978 , \49074 );
and \g132046/U$3 ( \62070 , \49075 , \53300 );
nor \g132046/U$1 ( \62071 , \62069 , \62070 );
not \g132001/U$3 ( \62072 , \62071 );
not \g132001/U$4 ( \62073 , \49014 );
and \g132001/U$2 ( \62074 , \62072 , \62073 );
and \g132001/U$5 ( \62075 , \62071 , \49014 );
nor \g132001/U$1 ( \62076 , \62074 , \62075 );
xor \g456150/U$1_r1 ( \62077 , \62068 , \62076 );
xor \g456114/U$5 ( \62078 , \61760 , \61768 );
and \g456114/U$4 ( \62079 , \62078 , \61823 );
and \g456114/U$6 ( \62080 , \61760 , \61768 );
or \g456114/U$3 ( \62081 , \62079 , \62080 );
xor \g131680/U$1 ( \62082 , \62077 , \62081 );
not \g131334/U$4 ( \62083 , \62082 );
and \g131334/U$2 ( \62084 , \62052 , \62083 );
and \g131334/U$5 ( \62085 , \62051 , \62082 );
nor \g131334/U$1 ( \62086 , \62084 , \62085 );
xor \g131247/U$1_r1 ( \62087 , \62043 , \62086 );
xor \g456090/U$2 ( \62088 , \62030 , \62087 );
xor \g456099/U$4 ( \62089 , \61962 , \62004 );
and \g456099/U$3 ( \62090 , \62089 , \62009 );
and \g456099/U$5 ( \62091 , \61962 , \62004 );
nor \g456099/U$2 ( \62092 , \62090 , \62091 );
xor \g456090/U$1 ( \62093 , \62088 , \62092 );
xor \g456096/U$4 ( \62094 , \61895 , \61899 );
and \g456096/U$3 ( \62095 , \62094 , \62010 );
and \g456096/U$5 ( \62096 , \61895 , \61899 );
nor \g456096/U$2 ( \62097 , \62095 , \62096 );
xor \g131244/U$4 ( \62098 , \61866 , \61888 );
and \g131244/U$3 ( \62099 , \62098 , \61894 );
and \g131244/U$5 ( \62100 , \61866 , \61888 );
or \g131244/U$2 ( \62101 , \62099 , \62100 );
not \g130920/U$3 ( \62102 , \62101 );
not \g131230/U$3 ( \62103 , \51124 );
and \g131275/U$2 ( \62104 , \50752 , \51518 );
and \g131275/U$3 ( \62105 , \51517 , \50443 );
nor \g131275/U$1 ( \62106 , \62104 , \62105 );
not \g131230/U$4 ( \62107 , \62106 );
or \g131230/U$2 ( \62108 , \62103 , \62107 );
or \g131230/U$5 ( \62109 , \62106 , \51124 );
nand \g131230/U$1 ( \62110 , \62108 , \62109 );
xor \g131883/U$4 ( \62111 , \61912 , \61920 );
and \g131883/U$3 ( \62112 , \62111 , \61951 );
and \g131883/U$5 ( \62113 , \61912 , \61920 );
or \g131883/U$2 ( \62114 , \62112 , \62113 );
xor \g131054/U$1 ( \62115 , \62110 , \62114 );
not \g131099/U$3 ( \62116 , \51120 );
and \g131149/U$2 ( \62117 , \50305 , \52273 );
and \g131149/U$3 ( \62118 , \52270 , \50019 );
nor \g131149/U$1 ( \62119 , \62117 , \62118 );
not \g131099/U$4 ( \62120 , \62119 );
or \g131099/U$2 ( \62121 , \62116 , \62120 );
or \g131099/U$5 ( \62122 , \62119 , \51120 );
nand \g131099/U$1 ( \62123 , \62121 , \62122 );
xor \g131054/U$1_r1 ( \62124 , \62115 , \62123 );
not \g131003/U$3 ( \62125 , \62124 );
xor \g456102/U$4 ( \62126 , \61986 , \61994 );
and \g456102/U$3 ( \62127 , \62126 , \62003 );
and \g456102/U$5 ( \62128 , \61986 , \61994 );
nor \g456102/U$2 ( \62129 , \62127 , \62128 );
not \g131003/U$4 ( \62130 , \62129 );
and \g131003/U$2 ( \62131 , \62125 , \62130 );
and \g131003/U$5 ( \62132 , \62124 , \62129 );
nor \g131003/U$1 ( \62133 , \62131 , \62132 );
not \g130978/U$3 ( \62134 , \62133 );
xor \g131871/U$4 ( \62135 , \61970 , \61978 );
and \g131871/U$3 ( \62136 , \62135 , \61985 );
and \g131871/U$5 ( \62137 , \61970 , \61978 );
or \g131871/U$2 ( \62138 , \62136 , \62137 );
or \g132110/U$2 ( \62139 , \61785 , \61797 );
not \g132113/U$3 ( \62140 , \61797 );
not \g132113/U$4 ( \62141 , \61785 );
or \g132113/U$2 ( \62142 , \62140 , \62141 );
nand \g132113/U$1 ( \62143 , \62142 , \61770 );
nand \g132110/U$1 ( \62144 , \62139 , \62143 );
not \g132523/U$3 ( \62145 , \48323 );
and \g132573/U$2 ( \62146 , \54251 , \48334 );
and \g132573/U$3 ( \62147 , \48335 , \54529 );
nor \g132573/U$1 ( \62148 , \62146 , \62147 );
not \g132523/U$4 ( \62149 , \62148 );
or \g132523/U$2 ( \62150 , \62145 , \62149 );
or \g132523/U$5 ( \62151 , \62148 , \48323 );
nand \g132523/U$1 ( \62152 , \62150 , \62151 );
xor \g131985/U$1 ( \62153 , \62144 , \62152 );
not \g132188/U$2 ( \62154 , \61779 );
nor \g132188/U$1 ( \62155 , \62154 , \61781 );
and \g132407/U$2 ( \62156 , \47914 , \56446 );
and \g132407/U$3 ( \62157 , \56167 , \47913 );
nor \g132407/U$1 ( \62158 , \62156 , \62157 );
and \g132325/U$2 ( \62159 , \62158 , \47977 );
not \g132325/U$4 ( \62160 , \62158 );
and \g132325/U$3 ( \62161 , \62160 , \47976 );
nor \g132325/U$1 ( \62162 , \62159 , \62161 );
xor \g132076/U$1 ( \62163 , \62155 , \62162 );
not \g135553/U$2 ( \62164 , \56359 );
nor \g135553/U$1 ( \62165 , \62164 , \40060 );
not \g132216/U$3 ( \62166 , \47948 );
and \g132270/U$2 ( \62167 , \47960 , \56357 );
and \g132270/U$3 ( \62168 , \56448 , \47959 );
nor \g132270/U$1 ( \62169 , \62167 , \62168 );
not \g132216/U$4 ( \62170 , \62169 );
or \g132216/U$2 ( \62171 , \62166 , \62170 );
or \g132216/U$5 ( \62172 , \62169 , \47948 );
nand \g132216/U$1 ( \62173 , \62171 , \62172 );
xor \g132162/U$1 ( \62174 , \62165 , \62173 );
xor \g132076/U$1_r1 ( \62175 , \62163 , \62174 );
xor \g131985/U$1_r1 ( \62176 , \62153 , \62175 );
xor \g131433/U$1 ( \62177 , \62138 , \62176 );
not \g131476/U$3 ( \62178 , \50362 );
and \g131506/U$2 ( \62179 , \51564 , \50588 );
and \g131506/U$3 ( \62180 , \50587 , \51098 );
nor \g131506/U$1 ( \62181 , \62179 , \62180 );
not \g131476/U$4 ( \62182 , \62181 );
or \g131476/U$2 ( \62183 , \62178 , \62182 );
or \g131476/U$5 ( \62184 , \62181 , \50362 );
nand \g131476/U$1 ( \62185 , \62183 , \62184 );
xor \g131433/U$1_r1 ( \62186 , \62177 , \62185 );
not \g130978/U$4 ( \62187 , \62186 );
and \g130978/U$2 ( \62188 , \62134 , \62187 );
and \g130978/U$5 ( \62189 , \62133 , \62186 );
nor \g130978/U$1 ( \62190 , \62188 , \62189 );
not \g130920/U$4 ( \62191 , \62190 );
or \g130920/U$2 ( \62192 , \62102 , \62191 );
or \g130920/U$5 ( \62193 , \62190 , \62101 );
nand \g130920/U$1 ( \62194 , \62192 , \62193 );
not \g130913/U$3 ( \62195 , \62194 );
and \g131888/U$2 ( \62196 , \52620 , \49403 );
and \g131888/U$3 ( \62197 , \49405 , \52883 );
nor \g131888/U$1 ( \62198 , \62196 , \62197 );
not \g131846/U$3 ( \62199 , \62198 );
not \g131846/U$4 ( \62200 , \49233 );
and \g131846/U$2 ( \62201 , \62199 , \62200 );
and \g131846/U$5 ( \62202 , \62198 , \49233 );
nor \g131846/U$1 ( \62203 , \62201 , \62202 );
not \g131809/U$3 ( \62204 , \62203 );
or \g131939/U$2 ( \62205 , \61801 , \61819 );
not \g131943/U$3 ( \62206 , \61819 );
not \g131943/U$4 ( \62207 , \61801 );
or \g131943/U$2 ( \62208 , \62206 , \62207 );
nand \g131943/U$1 ( \62209 , \62208 , \61806 );
nand \g131939/U$1 ( \62210 , \62205 , \62209 );
not \g131809/U$4 ( \62211 , \62210 );
or \g131809/U$2 ( \62212 , \62204 , \62211 );
or \g131809/U$5 ( \62213 , \62210 , \62203 );
nand \g131809/U$1 ( \62214 , \62212 , \62213 );
not \g131588/U$3 ( \62215 , \62214 );
and \g131625/U$2 ( \62216 , \51604 , \50159 );
and \g131625/U$3 ( \62217 , \50160 , \51854 );
nor \g131625/U$1 ( \62218 , \62216 , \62217 );
not \g131596/U$3 ( \62219 , \62218 );
not \g131596/U$4 ( \62220 , \49925 );
and \g131596/U$2 ( \62221 , \62219 , \62220 );
and \g131596/U$5 ( \62222 , \62218 , \49925 );
nor \g131596/U$1 ( \62223 , \62221 , \62222 );
not \g131588/U$4 ( \62224 , \62223 );
and \g131588/U$2 ( \62225 , \62215 , \62224 );
and \g131588/U$5 ( \62226 , \62214 , \62223 );
nor \g131588/U$1 ( \62227 , \62225 , \62226 );
not \g131464/U$3 ( \62228 , \62227 );
xor \g131495/U$4 ( \62229 , \61870 , \61878 );
and \g131495/U$3 ( \62230 , \62229 , \61887 );
and \g131495/U$5 ( \62231 , \61870 , \61878 );
or \g131495/U$2 ( \62232 , \62230 , \62231 );
not \g131464/U$4 ( \62233 , \62232 );
and \g131464/U$2 ( \62234 , \62228 , \62233 );
and \g131464/U$5 ( \62235 , \62227 , \62232 );
nor \g131464/U$1 ( \62236 , \62234 , \62235 );
not \g131434/U$3 ( \62237 , \62236 );
not \g132595/U$3 ( \62238 , \47997 );
and \g132643/U$2 ( \62239 , \48063 , \55127 );
and \g132643/U$3 ( \62240 , \55460 , \48064 );
nor \g132643/U$1 ( \62241 , \62239 , \62240 );
not \g132595/U$4 ( \62242 , \62241 );
or \g132595/U$2 ( \62243 , \62238 , \62242 );
or \g132595/U$5 ( \62244 , \62241 , \47997 );
nand \g132595/U$1 ( \62245 , \62243 , \62244 );
not \g132674/U$3 ( \62246 , \48159 );
and \g132719/U$2 ( \62247 , \48155 , \54853 );
and \g132719/U$3 ( \62248 , \54537 , \48154 );
nor \g132719/U$1 ( \62249 , \62247 , \62248 );
not \g132674/U$4 ( \62250 , \62249 );
or \g132674/U$2 ( \62251 , \62246 , \62250 );
or \g132674/U$5 ( \62252 , \62249 , \48159 );
nand \g132674/U$1 ( \62253 , \62251 , \62252 );
xor \g456138/U$2 ( \62254 , \62245 , \62253 );
not \g132475/U$3 ( \62255 , \47935 );
and \g132551/U$2 ( \62256 , \47931 , \55884 );
and \g132551/U$3 ( \62257 , \55707 , \47930 );
nor \g132551/U$1 ( \62258 , \62256 , \62257 );
not \g132475/U$4 ( \62259 , \62258 );
or \g132475/U$2 ( \62260 , \62255 , \62259 );
or \g132475/U$5 ( \62261 , \62258 , \47935 );
nand \g132475/U$1 ( \62262 , \62260 , \62261 );
xor \g456138/U$1 ( \62263 , \62254 , \62262 );
not \g132147/U$3 ( \62264 , \48685 );
and \g132199/U$2 ( \62265 , \53610 , \48858 );
and \g132199/U$3 ( \62266 , \48860 , \53848 );
nor \g132199/U$1 ( \62267 , \62265 , \62266 );
not \g132147/U$4 ( \62268 , \62267 );
or \g132147/U$2 ( \62269 , \62264 , \62268 );
or \g132147/U$5 ( \62270 , \62267 , \48685 );
nand \g132147/U$1 ( \62271 , \62269 , \62270 );
not \g131721/U$3 ( \62272 , \49568 );
and \g131754/U$2 ( \62273 , \52108 , \49812 );
and \g131754/U$3 ( \62274 , \49813 , \52352 );
nor \g131754/U$1 ( \62275 , \62273 , \62274 );
not \g131721/U$4 ( \62276 , \62275 );
or \g131721/U$2 ( \62277 , \62272 , \62276 );
or \g131721/U$5 ( \62278 , \62275 , \49568 );
nand \g131721/U$1 ( \62279 , \62277 , \62278 );
xor \g456138/U$1_r1 ( \62280 , \62271 , \62279 );
xor \g456138/U$1_r2 ( \62281 , \62263 , \62280 );
not \g131434/U$4 ( \62282 , \62281 );
and \g131434/U$2 ( \62283 , \62237 , \62282 );
and \g131434/U$5 ( \62284 , \62236 , \62281 );
nor \g131434/U$1 ( \62285 , \62283 , \62284 );
not \g130913/U$4 ( \62286 , \62285 );
and \g130913/U$2 ( \62287 , \62195 , \62286 );
and \g130913/U$5 ( \62288 , \62194 , \62285 );
nor \g130913/U$1 ( \62289 , \62287 , \62288 );
xor \g456090/U$1_r1 ( \62290 , \62097 , \62289 );
xor \g456090/U$1_r2 ( \62291 , \62093 , \62290 );
not \g128812/U$2 ( \62292 , \62291 );
xor \g128813/U$1 ( \62293 , \62022 , \62018 );
nand \g128812/U$1 ( \62294 , \62292 , \62293 );
not \g128810/U$1 ( \62295 , \62294 );
nor \g128815/U$1 ( \62296 , \62013 , \61733 );
nor \g128809/U$1 ( \62297 , \62023 , \62295 , \62296 );
xor \g456090/U$9 ( \62298 , \62030 , \62087 );
xor \g456090/U$9_r1 ( \62299 , \62298 , \62092 );
and \g456090/U$8 ( \62300 , \62097 , \62299 );
xor \g456090/U$11 ( \62301 , \62030 , \62087 );
xor \g456090/U$11_r1 ( \62302 , \62301 , \62092 );
and \g456090/U$10 ( \62303 , \62289 , \62302 );
and \g456090/U$12 ( \62304 , \62097 , \62289 );
or \g456090/U$7 ( \62305 , \62300 , \62303 , \62304 );
or \g128805/U$2 ( \62306 , \62297 , \62305 );
xor \g456090/U$5 ( \62307 , \62030 , \62087 );
and \g456090/U$4 ( \62308 , \62307 , \62092 );
and \g456090/U$6 ( \62309 , \62030 , \62087 );
or \g456090/U$3 ( \62310 , \62308 , \62309 );
not \g130783/U$3 ( \62311 , \62310 );
not \g131243/U$1 ( \62312 , \62101 );
or \g130941/U$2 ( \62313 , \62312 , \62285 );
and \g130948/U$2 ( \62314 , \62312 , \62285 );
nor \g130948/U$1 ( \62315 , \62314 , \62190 );
not \g130947/U$1 ( \62316 , \62315 );
nand \g130941/U$1 ( \62317 , \62313 , \62316 );
not \g132079/U$3 ( \62318 , \48685 );
and \g132121/U$2 ( \62319 , \53610 , \48860 );
and \g132121/U$3 ( \62320 , \48858 , \53300 );
nor \g132121/U$1 ( \62321 , \62319 , \62320 );
not \g132079/U$4 ( \62322 , \62321 );
or \g132079/U$2 ( \62323 , \62318 , \62322 );
or \g132079/U$5 ( \62324 , \62321 , \48685 );
nand \g132079/U$1 ( \62325 , \62323 , \62324 );
not \g132245/U$3 ( \62326 , \48483 );
and \g132295/U$2 ( \62327 , \53848 , \48478 );
and \g132295/U$3 ( \62328 , \48479 , \54015 );
nor \g132295/U$1 ( \62329 , \62327 , \62328 );
not \g132245/U$4 ( \62330 , \62329 );
or \g132245/U$2 ( \62331 , \62326 , \62330 );
or \g132245/U$5 ( \62332 , \62329 , \48483 );
nand \g132245/U$1 ( \62333 , \62331 , \62332 );
xor \g131978/U$1 ( \62334 , \62325 , \62333 );
and \g132162/U$2 ( \62335 , \62165 , \62173 );
and \g132406/U$2 ( \62336 , \47914 , \56167 );
and \g132406/U$3 ( \62337 , \55884 , \47913 );
nor \g132406/U$1 ( \62338 , \62336 , \62337 );
and \g132324/U$2 ( \62339 , \62338 , \47977 );
not \g132324/U$4 ( \62340 , \62338 );
and \g132324/U$3 ( \62341 , \62340 , \47976 );
nor \g132324/U$1 ( \62342 , \62339 , \62341 );
xor \g132075/U$1 ( \62343 , \62335 , \62342 );
not \g135552/U$2 ( \62344 , \56357 );
nor \g135552/U$1 ( \62345 , \62344 , \40060 );
not \g132215/U$3 ( \62346 , \47948 );
and \g132269/U$2 ( \62347 , \47959 , \56446 );
and \g132269/U$3 ( \62348 , \56448 , \47960 );
nor \g132269/U$1 ( \62349 , \62347 , \62348 );
not \g132215/U$4 ( \62350 , \62349 );
or \g132215/U$2 ( \62351 , \62346 , \62350 );
or \g132215/U$5 ( \62352 , \62349 , \47948 );
nand \g132215/U$1 ( \62353 , \62351 , \62352 );
xor \g132176/U$1 ( \62354 , \62345 , \62353 );
xor \g132075/U$1_r1 ( \62355 , \62343 , \62354 );
xor \g131978/U$1_r1 ( \62356 , \62334 , \62355 );
xor \g456138/U$9 ( \62357 , \62245 , \62253 );
xor \g456138/U$9_r1 ( \62358 , \62357 , \62262 );
and \g456138/U$8 ( \62359 , \62271 , \62358 );
xor \g456138/U$11 ( \62360 , \62245 , \62253 );
xor \g456138/U$11_r1 ( \62361 , \62360 , \62262 );
and \g456138/U$10 ( \62362 , \62279 , \62361 );
and \g456138/U$12 ( \62363 , \62271 , \62279 );
or \g456138/U$7 ( \62364 , \62359 , \62362 , \62363 );
xor \g456107/U$2 ( \62365 , \62356 , \62364 );
xor \g131985/U$4 ( \62366 , \62144 , \62152 );
and \g131985/U$3 ( \62367 , \62366 , \62175 );
and \g131985/U$5 ( \62368 , \62144 , \62152 );
or \g131985/U$2 ( \62369 , \62367 , \62368 );
not \g131916/U$3 ( \62370 , \49014 );
and \g131954/U$2 ( \62371 , \52978 , \49075 );
and \g131954/U$3 ( \62372 , \49074 , \52883 );
nor \g131954/U$1 ( \62373 , \62371 , \62372 );
not \g131916/U$4 ( \62374 , \62373 );
or \g131916/U$2 ( \62375 , \62370 , \62374 );
or \g131916/U$5 ( \62376 , \62373 , \49014 );
nand \g131916/U$1 ( \62377 , \62375 , \62376 );
xor \g131865/U$1 ( \62378 , \62369 , \62377 );
not \g132474/U$3 ( \62379 , \47935 );
and \g132540/U$2 ( \62380 , \47930 , \55460 );
and \g132540/U$3 ( \62381 , \55707 , \47931 );
nor \g132540/U$1 ( \62382 , \62380 , \62381 );
not \g132474/U$4 ( \62383 , \62382 );
or \g132474/U$2 ( \62384 , \62379 , \62383 );
or \g132474/U$5 ( \62385 , \62382 , \47935 );
nand \g132474/U$1 ( \62386 , \62384 , \62385 );
not \g132593/U$3 ( \62387 , \47997 );
and \g132641/U$2 ( \62388 , \48063 , \54853 );
and \g132641/U$3 ( \62389 , \55127 , \48064 );
nor \g132641/U$1 ( \62390 , \62388 , \62389 );
not \g132593/U$4 ( \62391 , \62390 );
or \g132593/U$2 ( \62392 , \62387 , \62391 );
or \g132593/U$5 ( \62393 , \62390 , \47997 );
nand \g132593/U$1 ( \62394 , \62392 , \62393 );
xor \g131986/U$1 ( \62395 , \62386 , \62394 );
xor \g132076/U$4 ( \62396 , \62155 , \62162 );
and \g132076/U$3 ( \62397 , \62396 , \62174 );
and \g132076/U$5 ( \62398 , \62155 , \62162 );
or \g132076/U$2 ( \62399 , \62397 , \62398 );
xor \g131986/U$1_r1 ( \62400 , \62395 , \62399 );
xor \g131865/U$1_r1 ( \62401 , \62378 , \62400 );
xor \g456107/U$1 ( \62402 , \62365 , \62401 );
not \g131678/U$1 ( \62403 , \62281 );
or \g131471/U$2 ( \62404 , \62227 , \62403 );
not \g131473/U$3 ( \62405 , \62403 );
not \g131473/U$4 ( \62406 , \62227 );
or \g131473/U$2 ( \62407 , \62405 , \62406 );
nand \g131473/U$1 ( \62408 , \62407 , \62232 );
nand \g131471/U$1 ( \62409 , \62404 , \62408 );
or \g131332/U$2 ( \62410 , \62081 , \62077 );
and \g131339/U$2 ( \62411 , \62081 , \62077 );
nor \g131339/U$1 ( \62412 , \62411 , \62051 );
not \g131338/U$1 ( \62413 , \62412 );
nand \g131332/U$1 ( \62414 , \62410 , \62413 );
xor \g456107/U$1_r1 ( \62415 , \62409 , \62414 );
xor \g456107/U$1_r2 ( \62416 , \62402 , \62415 );
xor \g130828/U$1 ( \62417 , \62317 , \62416 );
xor \g131054/U$4 ( \62418 , \62110 , \62114 );
and \g131054/U$3 ( \62419 , \62418 , \62123 );
and \g131054/U$5 ( \62420 , \62110 , \62114 );
or \g131054/U$2 ( \62421 , \62419 , \62420 );
not \g131405/U$3 ( \62422 , \50362 );
and \g131440/U$2 ( \62423 , \51117 , \50587 );
and \g131440/U$3 ( \62424 , \50588 , \51098 );
nor \g131440/U$1 ( \62425 , \62423 , \62424 );
not \g131405/U$4 ( \62426 , \62425 );
or \g131405/U$2 ( \62427 , \62422 , \62426 );
or \g131405/U$5 ( \62428 , \62425 , \50362 );
nand \g131405/U$1 ( \62429 , \62427 , \62428 );
xor \g456150/U$4 ( \62430 , \62060 , \62067 );
and \g456150/U$3 ( \62431 , \62430 , \62076 );
and \g456150/U$5 ( \62432 , \62060 , \62067 );
nor \g456150/U$2 ( \62433 , \62431 , \62432 );
xor \g131130/U$1 ( \62434 , \62429 , \62433 );
not \g131177/U$3 ( \62435 , \51124 );
and \g131220/U$2 ( \62436 , \50305 , \51517 );
and \g131220/U$3 ( \62437 , \51518 , \50443 );
nor \g131220/U$1 ( \62438 , \62436 , \62437 );
not \g131177/U$4 ( \62439 , \62438 );
or \g131177/U$2 ( \62440 , \62435 , \62439 );
or \g131177/U$5 ( \62441 , \62438 , \51124 );
nand \g131177/U$1 ( \62442 , \62440 , \62441 );
xor \g131130/U$1_r1 ( \62443 , \62434 , \62442 );
xor \g130911/U$1 ( \62444 , \62421 , \62443 );
not \g131290/U$3 ( \62445 , \50759 );
and \g131316/U$2 ( \62446 , \50957 , \51055 );
and \g131316/U$3 ( \62447 , \51053 , \50752 );
nor \g131316/U$1 ( \62448 , \62446 , \62447 );
not \g131290/U$4 ( \62449 , \62448 );
or \g131290/U$2 ( \62450 , \62445 , \62449 );
or \g131290/U$5 ( \62451 , \62448 , \50759 );
nand \g131290/U$1 ( \62452 , \62450 , \62451 );
not \g132446/U$3 ( \62453 , \48323 );
and \g132493/U$2 ( \62454 , \54185 , \48334 );
and \g132493/U$3 ( \62455 , \48335 , \54251 );
nor \g132493/U$1 ( \62456 , \62454 , \62455 );
not \g132446/U$4 ( \62457 , \62456 );
or \g132446/U$2 ( \62458 , \62453 , \62457 );
or \g132446/U$5 ( \62459 , \62456 , \48323 );
nand \g132446/U$1 ( \62460 , \62458 , \62459 );
not \g132594/U$3 ( \62461 , \48159 );
and \g132642/U$2 ( \62462 , \48155 , \54537 );
and \g132642/U$3 ( \62463 , \48154 , \54529 );
nor \g132642/U$1 ( \62464 , \62462 , \62463 );
not \g132594/U$4 ( \62465 , \62464 );
or \g132594/U$2 ( \62466 , \62461 , \62465 );
or \g132594/U$5 ( \62467 , \62464 , \48159 );
nand \g132594/U$1 ( \62468 , \62466 , \62467 );
xor \g132259/U$1 ( \62469 , \62460 , \62468 );
xor \g456138/U$5 ( \62470 , \62245 , \62253 );
and \g456138/U$4 ( \62471 , \62470 , \62262 );
and \g456138/U$6 ( \62472 , \62245 , \62253 );
or \g456138/U$3 ( \62473 , \62471 , \62472 );
xor \g132259/U$1_r1 ( \62474 , \62469 , \62473 );
xor \g130977/U$1 ( \62475 , \62452 , \62474 );
not \g131018/U$3 ( \62476 , \51120 );
and \g131074/U$2 ( \62477 , \49888 , \52270 );
and \g131074/U$3 ( \62478 , \52273 , \50019 );
nor \g131074/U$1 ( \62479 , \62477 , \62478 );
not \g131018/U$4 ( \62480 , \62479 );
or \g131018/U$2 ( \62481 , \62476 , \62480 );
or \g131018/U$5 ( \62482 , \62479 , \51120 );
nand \g131018/U$1 ( \62483 , \62481 , \62482 );
xor \g130977/U$1_r1 ( \62484 , \62475 , \62483 );
xor \g130911/U$1_r1 ( \62485 , \62444 , \62484 );
xor \g130828/U$1_r1 ( \62486 , \62417 , \62485 );
not \g130783/U$4 ( \62487 , \62486 );
or \g130783/U$2 ( \62488 , \62311 , \62487 );
or \g130783/U$5 ( \62489 , \62486 , \62310 );
nand \g130783/U$1 ( \62490 , \62488 , \62489 );
not \g130773/U$3 ( \62491 , \62490 );
not \g131432/U$1 ( \62492 , \62186 );
or \g131008/U$2 ( \62493 , \62129 , \62492 );
not \g131013/U$3 ( \62494 , \62492 );
not \g131013/U$4 ( \62495 , \62129 );
or \g131013/U$2 ( \62496 , \62494 , \62495 );
nand \g131013/U$1 ( \62497 , \62496 , \62124 );
nand \g131008/U$1 ( \62498 , \62493 , \62497 );
not \g130919/U$3 ( \62499 , \62498 );
xor \g131247/U$4 ( \62500 , \62038 , \62042 );
and \g131247/U$3 ( \62501 , \62500 , \62086 );
and \g131247/U$5 ( \62502 , \62038 , \62042 );
or \g131247/U$2 ( \62503 , \62501 , \62502 );
not \g130919/U$4 ( \62504 , \62503 );
and \g130919/U$2 ( \62505 , \62499 , \62504 );
and \g130919/U$5 ( \62506 , \62498 , \62503 );
nor \g130919/U$1 ( \62507 , \62505 , \62506 );
not \g130912/U$3 ( \62508 , \62507 );
not \g131653/U$3 ( \62509 , \49568 );
and \g131686/U$2 ( \62510 , \52108 , \49813 );
and \g131686/U$3 ( \62511 , \49812 , \51854 );
nor \g131686/U$1 ( \62512 , \62510 , \62511 );
not \g131653/U$4 ( \62513 , \62512 );
or \g131653/U$2 ( \62514 , \62509 , \62513 );
or \g131653/U$5 ( \62515 , \62512 , \49568 );
nand \g131653/U$1 ( \62516 , \62514 , \62515 );
not \g131780/U$3 ( \62517 , \49233 );
and \g131813/U$2 ( \62518 , \52620 , \49405 );
and \g131813/U$3 ( \62519 , \49403 , \52352 );
nor \g131813/U$1 ( \62520 , \62518 , \62519 );
not \g131780/U$4 ( \62521 , \62520 );
or \g131780/U$2 ( \62522 , \62517 , \62521 );
or \g131780/U$5 ( \62523 , \62520 , \49233 );
nand \g131780/U$1 ( \62524 , \62522 , \62523 );
xor \g456116/U$2 ( \62525 , \62516 , \62524 );
not \g131541/U$3 ( \62526 , \49925 );
and \g131573/U$2 ( \62527 , \51604 , \50160 );
and \g131573/U$3 ( \62528 , \50159 , \51564 );
nor \g131573/U$1 ( \62529 , \62527 , \62528 );
not \g131541/U$4 ( \62530 , \62529 );
or \g131541/U$2 ( \62531 , \62526 , \62530 );
or \g131541/U$5 ( \62532 , \62529 , \49925 );
nand \g131541/U$1 ( \62533 , \62531 , \62532 );
xor \g456116/U$1 ( \62534 , \62525 , \62533 );
or \g131564/U$2 ( \62535 , \62223 , \62203 );
not \g131567/U$3 ( \62536 , \62203 );
not \g131567/U$4 ( \62537 , \62223 );
or \g131567/U$2 ( \62538 , \62536 , \62537 );
nand \g131567/U$1 ( \62539 , \62538 , \62210 );
nand \g131564/U$1 ( \62540 , \62535 , \62539 );
xor \g131433/U$4 ( \62541 , \62138 , \62176 );
and \g131433/U$3 ( \62542 , \62541 , \62185 );
and \g131433/U$5 ( \62543 , \62138 , \62176 );
or \g131433/U$2 ( \62544 , \62542 , \62543 );
xor \g456116/U$1_r1 ( \62545 , \62540 , \62544 );
xor \g456116/U$1_r2 ( \62546 , \62534 , \62545 );
not \g130912/U$4 ( \62547 , \62546 );
and \g130912/U$2 ( \62548 , \62508 , \62547 );
and \g130912/U$5 ( \62549 , \62507 , \62546 );
nor \g130912/U$1 ( \62550 , \62548 , \62549 );
not \g130773/U$4 ( \62551 , \62550 );
and \g130773/U$2 ( \62552 , \62491 , \62551 );
and \g130773/U$5 ( \62553 , \62490 , \62550 );
nor \g130773/U$1 ( \62554 , \62552 , \62553 );
not \g128807/U$2 ( \62555 , \62554 );
xor \g128808/U$1 ( \62556 , \62305 , \62297 );
nand \g128807/U$1 ( \62557 , \62555 , \62556 );
nand \g128805/U$1 ( \62558 , \62306 , \62557 );
or \g130801/U$2 ( \62559 , \62550 , \62310 );
not \g130803/U$3 ( \62560 , \62310 );
not \g130803/U$4 ( \62561 , \62550 );
or \g130803/U$2 ( \62562 , \62560 , \62561 );
nand \g130803/U$1 ( \62563 , \62562 , \62486 );
nand \g130801/U$1 ( \62564 , \62559 , \62563 );
and \g128802/U$2 ( \62565 , \62558 , \62564 );
not \g131363/U$1 ( \62566 , \62546 );
or \g130940/U$2 ( \62567 , \62503 , \62566 );
not \g130946/U$3 ( \62568 , \62566 );
not \g130946/U$4 ( \62569 , \62503 );
or \g130946/U$2 ( \62570 , \62568 , \62569 );
nand \g130946/U$1 ( \62571 , \62570 , \62498 );
nand \g130940/U$1 ( \62572 , \62567 , \62571 );
xor \g131865/U$4 ( \62573 , \62369 , \62377 );
and \g131865/U$3 ( \62574 , \62573 , \62400 );
and \g131865/U$5 ( \62575 , \62369 , \62377 );
or \g131865/U$2 ( \62576 , \62574 , \62575 );
not \g132000/U$3 ( \62577 , \48685 );
and \g132040/U$2 ( \62578 , \52978 , \48858 );
and \g132040/U$3 ( \62579 , \48860 , \53300 );
nor \g132040/U$1 ( \62580 , \62578 , \62579 );
not \g132000/U$4 ( \62581 , \62580 );
or \g132000/U$2 ( \62582 , \62577 , \62581 );
or \g132000/U$5 ( \62583 , \62580 , \48685 );
nand \g132000/U$1 ( \62584 , \62582 , \62583 );
not \g132146/U$3 ( \62585 , \48483 );
and \g132193/U$2 ( \62586 , \53610 , \48478 );
and \g132193/U$3 ( \62587 , \48479 , \53848 );
nor \g132193/U$1 ( \62588 , \62586 , \62587 );
not \g132146/U$4 ( \62589 , \62588 );
or \g132146/U$2 ( \62590 , \62585 , \62589 );
or \g132146/U$5 ( \62591 , \62588 , \48483 );
nand \g132146/U$1 ( \62592 , \62590 , \62591 );
xor \g131875/U$1 ( \62593 , \62584 , \62592 );
xor \g131986/U$4 ( \62594 , \62386 , \62394 );
and \g131986/U$3 ( \62595 , \62594 , \62399 );
and \g131986/U$5 ( \62596 , \62386 , \62394 );
or \g131986/U$2 ( \62597 , \62595 , \62596 );
xor \g131875/U$1_r1 ( \62598 , \62593 , \62597 );
xor \g456110/U$2 ( \62599 , \62576 , \62598 );
xor \g456116/U$5 ( \62600 , \62516 , \62524 );
and \g456116/U$4 ( \62601 , \62600 , \62533 );
and \g456116/U$6 ( \62602 , \62516 , \62524 );
or \g456116/U$3 ( \62603 , \62601 , \62602 );
xor \g456110/U$1 ( \62604 , \62599 , \62603 );
xor \g456107/U$5 ( \62605 , \62356 , \62364 );
and \g456107/U$4 ( \62606 , \62605 , \62401 );
and \g456107/U$6 ( \62607 , \62356 , \62364 );
or \g456107/U$3 ( \62608 , \62606 , \62607 );
xor \g456116/U$9 ( \62609 , \62516 , \62524 );
xor \g456116/U$9_r1 ( \62610 , \62609 , \62533 );
and \g456116/U$8 ( \62611 , \62540 , \62610 );
xor \g456116/U$11 ( \62612 , \62516 , \62524 );
xor \g456116/U$11_r1 ( \62613 , \62612 , \62533 );
and \g456116/U$10 ( \62614 , \62544 , \62613 );
and \g456116/U$12 ( \62615 , \62540 , \62544 );
or \g456116/U$7 ( \62616 , \62611 , \62614 , \62615 );
xor \g456110/U$1_r1 ( \62617 , \62608 , \62616 );
xor \g456110/U$1_r2 ( \62618 , \62604 , \62617 );
xor \g130806/U$1 ( \62619 , \62572 , \62618 );
xor \g130977/U$4 ( \62620 , \62452 , \62474 );
and \g130977/U$3 ( \62621 , \62620 , \62483 );
and \g130977/U$5 ( \62622 , \62452 , \62474 );
or \g130977/U$2 ( \62623 , \62621 , \62622 );
not \g131348/U$3 ( \62624 , \50362 );
and \g131371/U$2 ( \62625 , \51117 , \50588 );
and \g131371/U$3 ( \62626 , \50587 , \50957 );
nor \g131371/U$1 ( \62627 , \62625 , \62626 );
not \g131348/U$4 ( \62628 , \62627 );
or \g131348/U$2 ( \62629 , \62624 , \62628 );
or \g131348/U$5 ( \62630 , \62627 , \50362 );
nand \g131348/U$1 ( \62631 , \62629 , \62630 );
xor \g131978/U$4 ( \62632 , \62325 , \62333 );
and \g131978/U$3 ( \62633 , \62632 , \62355 );
and \g131978/U$5 ( \62634 , \62325 , \62333 );
or \g131978/U$2 ( \62635 , \62633 , \62634 );
xor \g131053/U$1 ( \62636 , \62631 , \62635 );
not \g131098/U$3 ( \62637 , \51124 );
and \g131148/U$2 ( \62638 , \50305 , \51518 );
and \g131148/U$3 ( \62639 , \51517 , \50019 );
nor \g131148/U$1 ( \62640 , \62638 , \62639 );
not \g131098/U$4 ( \62641 , \62640 );
or \g131098/U$2 ( \62642 , \62637 , \62641 );
or \g131098/U$5 ( \62643 , \62640 , \51124 );
nand \g131098/U$1 ( \62644 , \62642 , \62643 );
xor \g131053/U$1_r1 ( \62645 , \62636 , \62644 );
xor \g130858/U$1 ( \62646 , \62623 , \62645 );
not \g131229/U$3 ( \62647 , \50759 );
and \g131263/U$2 ( \62648 , \50752 , \51055 );
and \g131263/U$3 ( \62649 , \51053 , \50443 );
nor \g131263/U$1 ( \62650 , \62648 , \62649 );
not \g131229/U$4 ( \62651 , \62650 );
or \g131229/U$2 ( \62652 , \62647 , \62651 );
or \g131229/U$5 ( \62653 , \62650 , \50759 );
nand \g131229/U$1 ( \62654 , \62652 , \62653 );
not \g132326/U$3 ( \62655 , \48323 );
and \g132408/U$2 ( \62656 , \54185 , \48335 );
and \g132408/U$3 ( \62657 , \48334 , \54015 );
nor \g132408/U$1 ( \62658 , \62656 , \62657 );
not \g132326/U$4 ( \62659 , \62658 );
or \g132326/U$2 ( \62660 , \62655 , \62659 );
or \g132326/U$5 ( \62661 , \62658 , \48323 );
nand \g132326/U$1 ( \62662 , \62660 , \62661 );
not \g132522/U$3 ( \62663 , \48159 );
and \g132566/U$2 ( \62664 , \54251 , \48154 );
and \g132566/U$3 ( \62665 , \54529 , \48155 );
nor \g132566/U$1 ( \62666 , \62664 , \62665 );
not \g132522/U$4 ( \62667 , \62666 );
or \g132522/U$2 ( \62668 , \62663 , \62667 );
or \g132522/U$5 ( \62669 , \62666 , \48159 );
nand \g132522/U$1 ( \62670 , \62668 , \62669 );
xor \g131974/U$1 ( \62671 , \62662 , \62670 );
and \g132176/U$2 ( \62672 , \62345 , \62353 );
and \g132405/U$2 ( \62673 , \47914 , \55884 );
and \g132405/U$3 ( \62674 , \55707 , \47913 );
nor \g132405/U$1 ( \62675 , \62673 , \62674 );
and \g132323/U$2 ( \62676 , \62675 , \47977 );
not \g132323/U$4 ( \62677 , \62675 );
and \g132323/U$3 ( \62678 , \62677 , \47976 );
nor \g132323/U$1 ( \62679 , \62676 , \62678 );
xor \g132074/U$1 ( \62680 , \62672 , \62679 );
not \g135550/U$2 ( \62681 , \56448 );
nor \g135550/U$1 ( \62682 , \62681 , \40060 );
not \g132213/U$3 ( \62683 , \47948 );
and \g132267/U$2 ( \62684 , \47960 , \56446 );
and \g132267/U$3 ( \62685 , \56167 , \47959 );
nor \g132267/U$1 ( \62686 , \62684 , \62685 );
not \g132213/U$4 ( \62687 , \62686 );
or \g132213/U$2 ( \62688 , \62683 , \62687 );
or \g132213/U$5 ( \62689 , \62686 , \47948 );
nand \g132213/U$1 ( \62690 , \62688 , \62689 );
xor \g132177/U$1 ( \62691 , \62682 , \62690 );
xor \g132074/U$1_r1 ( \62692 , \62680 , \62691 );
xor \g131974/U$1_r1 ( \62693 , \62671 , \62692 );
xor \g130915/U$1 ( \62694 , \62654 , \62693 );
not \g130953/U$3 ( \62695 , \51120 );
and \g130995/U$2 ( \62696 , \49888 , \52273 );
and \g130995/U$3 ( \62697 , \52270 , \49714 );
nor \g130995/U$1 ( \62698 , \62696 , \62697 );
not \g130953/U$4 ( \62699 , \62698 );
or \g130953/U$2 ( \62700 , \62695 , \62699 );
or \g130953/U$5 ( \62701 , \62698 , \51120 );
nand \g130953/U$1 ( \62702 , \62700 , \62701 );
xor \g130915/U$1_r1 ( \62703 , \62694 , \62702 );
xor \g130858/U$1_r1 ( \62704 , \62646 , \62703 );
xor \g130806/U$1_r1 ( \62705 , \62619 , \62704 );
not \g130751/U$3 ( \62706 , \62705 );
not \g131593/U$3 ( \62707 , \49568 );
and \g131624/U$2 ( \62708 , \51604 , \49812 );
and \g131624/U$3 ( \62709 , \49813 , \51854 );
nor \g131624/U$1 ( \62710 , \62708 , \62709 );
not \g131593/U$4 ( \62711 , \62710 );
or \g131593/U$2 ( \62712 , \62707 , \62711 );
or \g131593/U$5 ( \62713 , \62710 , \49568 );
nand \g131593/U$1 ( \62714 , \62712 , \62713 );
xor \g132259/U$4 ( \62715 , \62460 , \62468 );
and \g132259/U$3 ( \62716 , \62715 , \62473 );
and \g132259/U$5 ( \62717 , \62460 , \62468 );
or \g132259/U$2 ( \62718 , \62716 , \62717 );
xor \g131431/U$1 ( \62719 , \62714 , \62718 );
not \g131475/U$3 ( \62720 , \49925 );
and \g131505/U$2 ( \62721 , \51564 , \50160 );
and \g131505/U$3 ( \62722 , \50159 , \51098 );
nor \g131505/U$1 ( \62723 , \62721 , \62722 );
not \g131475/U$4 ( \62724 , \62723 );
or \g131475/U$2 ( \62725 , \62720 , \62724 );
or \g131475/U$5 ( \62726 , \62723 , \49925 );
nand \g131475/U$1 ( \62727 , \62725 , \62726 );
xor \g131431/U$1_r1 ( \62728 , \62719 , \62727 );
not \g131720/U$3 ( \62729 , \49233 );
and \g131753/U$2 ( \62730 , \52108 , \49403 );
and \g131753/U$3 ( \62731 , \49405 , \52352 );
nor \g131753/U$1 ( \62732 , \62730 , \62731 );
not \g131720/U$4 ( \62733 , \62732 );
or \g131720/U$2 ( \62734 , \62729 , \62733 );
or \g131720/U$5 ( \62735 , \62732 , \49233 );
nand \g131720/U$1 ( \62736 , \62734 , \62735 );
not \g131845/U$3 ( \62737 , \49014 );
and \g131887/U$2 ( \62738 , \52620 , \49074 );
and \g131887/U$3 ( \62739 , \49075 , \52883 );
nor \g131887/U$1 ( \62740 , \62738 , \62739 );
not \g131845/U$4 ( \62741 , \62740 );
or \g131845/U$2 ( \62742 , \62737 , \62741 );
or \g131845/U$5 ( \62743 , \62740 , \49014 );
nand \g131845/U$1 ( \62744 , \62742 , \62743 );
xor \g131670/U$1 ( \62745 , \62736 , \62744 );
not \g132481/U$3 ( \62746 , \47935 );
and \g132539/U$2 ( \62747 , \47930 , \55127 );
and \g132539/U$3 ( \62748 , \55460 , \47931 );
nor \g132539/U$1 ( \62749 , \62747 , \62748 );
not \g132481/U$4 ( \62750 , \62749 );
or \g132481/U$2 ( \62751 , \62746 , \62750 );
or \g132481/U$5 ( \62752 , \62749 , \47935 );
nand \g132481/U$1 ( \62753 , \62751 , \62752 );
not \g132601/U$3 ( \62754 , \47997 );
and \g132665/U$2 ( \62755 , \48064 , \54853 );
and \g132665/U$3 ( \62756 , \54537 , \48063 );
nor \g132665/U$1 ( \62757 , \62755 , \62756 );
not \g132601/U$4 ( \62758 , \62757 );
or \g132601/U$2 ( \62759 , \62754 , \62758 );
or \g132601/U$5 ( \62760 , \62757 , \47997 );
nand \g132601/U$1 ( \62761 , \62759 , \62760 );
xor \g131984/U$1 ( \62762 , \62753 , \62761 );
xor \g132075/U$4 ( \62763 , \62335 , \62342 );
and \g132075/U$3 ( \62764 , \62763 , \62354 );
and \g132075/U$5 ( \62765 , \62335 , \62342 );
or \g132075/U$2 ( \62766 , \62764 , \62765 );
xor \g131984/U$1_r1 ( \62767 , \62762 , \62766 );
xor \g131670/U$1_r1 ( \62768 , \62745 , \62767 );
xor \g456089/U$2 ( \62769 , \62728 , \62768 );
xor \g131130/U$4 ( \62770 , \62429 , \62433 );
and \g131130/U$3 ( \62771 , \62770 , \62442 );
and \g131130/U$5 ( \62772 , \62429 , \62433 );
or \g131130/U$2 ( \62773 , \62771 , \62772 );
xor \g456089/U$1 ( \62774 , \62769 , \62773 );
xor \g456107/U$9 ( \62775 , \62356 , \62364 );
xor \g456107/U$9_r1 ( \62776 , \62775 , \62401 );
and \g456107/U$8 ( \62777 , \62409 , \62776 );
xor \g456107/U$11 ( \62778 , \62356 , \62364 );
xor \g456107/U$11_r1 ( \62779 , \62778 , \62401 );
and \g456107/U$10 ( \62780 , \62414 , \62779 );
and \g456107/U$12 ( \62781 , \62409 , \62414 );
or \g456107/U$7 ( \62782 , \62777 , \62780 , \62781 );
xor \g130911/U$4 ( \62783 , \62421 , \62443 );
and \g130911/U$3 ( \62784 , \62783 , \62484 );
and \g130911/U$5 ( \62785 , \62421 , \62443 );
or \g130911/U$2 ( \62786 , \62784 , \62785 );
xor \g456089/U$1_r1 ( \62787 , \62782 , \62786 );
xor \g456089/U$1_r2 ( \62788 , \62774 , \62787 );
xor \g130828/U$4 ( \62789 , \62317 , \62416 );
and \g130828/U$3 ( \62790 , \62789 , \62485 );
and \g130828/U$5 ( \62791 , \62317 , \62416 );
or \g130828/U$2 ( \62792 , \62790 , \62791 );
xnor \g130788/U$1 ( \62793 , \62788 , \62792 );
not \g130751/U$4 ( \62794 , \62793 );
or \g130751/U$2 ( \62795 , \62706 , \62794 );
or \g130751/U$5 ( \62796 , \62793 , \62705 );
nand \g130751/U$1 ( \62797 , \62795 , \62796 );
xor \g128804/U$1 ( \62798 , \62564 , \62558 );
and \g128803/U$2 ( \62799 , \62797 , \62798 );
nor \g128802/U$1 ( \62800 , \62565 , \62799 );
or \g130802/U$1 ( \62801 , \62792 , \62788 );
and \g130750/U$2 ( \62802 , \62705 , \62801 );
and \g130750/U$3 ( \62803 , \62788 , \62792 );
nor \g130750/U$1 ( \62804 , \62802 , \62803 );
or \g128798/U$2 ( \62805 , \62800 , \62804 );
xor \g130806/U$4 ( \62806 , \62572 , \62618 );
and \g130806/U$3 ( \62807 , \62806 , \62704 );
and \g130806/U$5 ( \62808 , \62572 , \62618 );
or \g130806/U$2 ( \62809 , \62807 , \62808 );
xor \g456089/U$9 ( \62810 , \62728 , \62768 );
xor \g456089/U$9_r1 ( \62811 , \62810 , \62773 );
and \g456089/U$8 ( \62812 , \62782 , \62811 );
xor \g456089/U$11 ( \62813 , \62728 , \62768 );
xor \g456089/U$11_r1 ( \62814 , \62813 , \62773 );
and \g456089/U$10 ( \62815 , \62786 , \62814 );
and \g456089/U$12 ( \62816 , \62782 , \62786 );
or \g456089/U$7 ( \62817 , \62812 , \62815 , \62816 );
xor \g130604/U$1 ( \62818 , \62809 , \62817 );
and \g132402/U$2 ( \62819 , \47913 , \55460 );
and \g132402/U$3 ( \62820 , \55707 , \47914 );
nor \g132402/U$1 ( \62821 , \62819 , \62820 );
and \g132320/U$2 ( \62822 , \62821 , \47977 );
not \g132320/U$4 ( \62823 , \62821 );
and \g132320/U$3 ( \62824 , \62823 , \47976 );
nor \g132320/U$1 ( \62825 , \62822 , \62824 );
not \g132471/U$3 ( \62826 , \47935 );
and \g132537/U$2 ( \62827 , \47930 , \54853 );
and \g132537/U$3 ( \62828 , \55127 , \47931 );
nor \g132537/U$1 ( \62829 , \62827 , \62828 );
not \g132471/U$4 ( \62830 , \62829 );
or \g132471/U$2 ( \62831 , \62826 , \62830 );
or \g132471/U$5 ( \62832 , \62829 , \47935 );
nand \g132471/U$1 ( \62833 , \62831 , \62832 );
xor \g132073/U$1 ( \62834 , \62825 , \62833 );
and \g132177/U$2 ( \62835 , \62682 , \62690 );
xor \g132073/U$1_r1 ( \62836 , \62834 , \62835 );
not \g131779/U$3 ( \62837 , \49014 );
and \g131812/U$2 ( \62838 , \52620 , \49075 );
and \g131812/U$3 ( \62839 , \49074 , \52352 );
nor \g131812/U$1 ( \62840 , \62838 , \62839 );
not \g131779/U$4 ( \62841 , \62840 );
or \g131779/U$2 ( \62842 , \62837 , \62841 );
or \g131779/U$5 ( \62843 , \62840 , \49014 );
nand \g131779/U$1 ( \62844 , \62842 , \62843 );
xor \g456118/U$2 ( \62845 , \62836 , \62844 );
xor \g131984/U$4 ( \62846 , \62753 , \62761 );
and \g131984/U$3 ( \62847 , \62846 , \62766 );
and \g131984/U$5 ( \62848 , \62753 , \62761 );
or \g131984/U$2 ( \62849 , \62847 , \62848 );
xor \g456118/U$1 ( \62850 , \62845 , \62849 );
not \g132244/U$3 ( \62851 , \48323 );
and \g132294/U$2 ( \62852 , \53848 , \48334 );
and \g132294/U$3 ( \62853 , \48335 , \54015 );
nor \g132294/U$1 ( \62854 , \62852 , \62853 );
not \g132244/U$4 ( \62855 , \62854 );
or \g132244/U$2 ( \62856 , \62851 , \62855 );
or \g132244/U$5 ( \62857 , \62854 , \48323 );
nand \g132244/U$1 ( \62858 , \62856 , \62857 );
not \g132445/U$3 ( \62859 , \48159 );
and \g132492/U$2 ( \62860 , \54185 , \48154 );
and \g132492/U$3 ( \62861 , \54251 , \48155 );
nor \g132492/U$1 ( \62862 , \62860 , \62861 );
not \g132445/U$4 ( \62863 , \62862 );
or \g132445/U$2 ( \62864 , \62859 , \62863 );
or \g132445/U$5 ( \62865 , \62862 , \48159 );
nand \g132445/U$1 ( \62866 , \62864 , \62865 );
xor \g132032/U$1 ( \62867 , \62858 , \62866 );
not \g132078/U$3 ( \62868 , \48483 );
and \g132120/U$2 ( \62869 , \53610 , \48479 );
and \g132120/U$3 ( \62870 , \48478 , \53300 );
nor \g132120/U$1 ( \62871 , \62869 , \62870 );
not \g132078/U$4 ( \62872 , \62871 );
or \g132078/U$2 ( \62873 , \62868 , \62872 );
or \g132078/U$5 ( \62874 , \62871 , \48483 );
nand \g132078/U$1 ( \62875 , \62873 , \62874 );
xor \g132032/U$1_r1 ( \62876 , \62867 , \62875 );
xor \g131431/U$4 ( \62877 , \62714 , \62718 );
and \g131431/U$3 ( \62878 , \62877 , \62727 );
and \g131431/U$5 ( \62879 , \62714 , \62718 );
or \g131431/U$2 ( \62880 , \62878 , \62879 );
xor \g456118/U$1_r1 ( \62881 , \62876 , \62880 );
xor \g456118/U$1_r2 ( \62882 , \62850 , \62881 );
xor \g456110/U$5 ( \62883 , \62576 , \62598 );
and \g456110/U$4 ( \62884 , \62883 , \62603 );
and \g456110/U$6 ( \62885 , \62576 , \62598 );
or \g456110/U$3 ( \62886 , \62884 , \62885 );
xor \g456082/U$2 ( \62887 , \62882 , \62886 );
xor \g456089/U$5 ( \62888 , \62728 , \62768 );
and \g456089/U$4 ( \62889 , \62888 , \62773 );
and \g456089/U$6 ( \62890 , \62728 , \62768 );
or \g456089/U$3 ( \62891 , \62889 , \62890 );
xor \g456082/U$1 ( \62892 , \62887 , \62891 );
xor \g456110/U$9 ( \62893 , \62576 , \62598 );
xor \g456110/U$9_r1 ( \62894 , \62893 , \62603 );
and \g456110/U$8 ( \62895 , \62608 , \62894 );
xor \g456110/U$11 ( \62896 , \62576 , \62598 );
xor \g456110/U$11_r1 ( \62897 , \62896 , \62603 );
and \g456110/U$10 ( \62898 , \62616 , \62897 );
and \g456110/U$12 ( \62899 , \62608 , \62616 );
or \g456110/U$7 ( \62900 , \62895 , \62898 , \62899 );
xor \g130858/U$4 ( \62901 , \62623 , \62645 );
and \g130858/U$3 ( \62902 , \62901 , \62703 );
and \g130858/U$5 ( \62903 , \62623 , \62645 );
or \g130858/U$2 ( \62904 , \62902 , \62903 );
not \g135548/U$2 ( \62905 , \56446 );
nor \g135548/U$1 ( \62906 , \62905 , \40060 );
not \g132214/U$3 ( \62907 , \47948 );
and \g132268/U$2 ( \62908 , \47960 , \56167 );
and \g132268/U$3 ( \62909 , \55884 , \47959 );
nor \g132268/U$1 ( \62910 , \62908 , \62909 );
not \g132214/U$4 ( \62911 , \62910 );
or \g132214/U$2 ( \62912 , \62907 , \62911 );
or \g132214/U$5 ( \62913 , \62910 , \47948 );
nand \g132214/U$1 ( \62914 , \62912 , \62913 );
xor \g132167/U$1 ( \62915 , \62906 , \62914 );
not \g132592/U$3 ( \62916 , \47997 );
and \g132639/U$2 ( \62917 , \48064 , \54537 );
and \g132639/U$3 ( \62918 , \54529 , \48063 );
nor \g132639/U$1 ( \62919 , \62917 , \62918 );
not \g132592/U$4 ( \62920 , \62919 );
or \g132592/U$2 ( \62921 , \62916 , \62920 );
or \g132592/U$5 ( \62922 , \62919 , \47997 );
nand \g132592/U$1 ( \62923 , \62921 , \62922 );
xor \g131983/U$1 ( \62924 , \62915 , \62923 );
xor \g132074/U$4 ( \62925 , \62672 , \62679 );
and \g132074/U$3 ( \62926 , \62925 , \62691 );
and \g132074/U$5 ( \62927 , \62672 , \62679 );
or \g132074/U$2 ( \62928 , \62926 , \62927 );
xor \g131983/U$1_r1 ( \62929 , \62924 , \62928 );
not \g131652/U$3 ( \62930 , \49233 );
and \g131685/U$2 ( \62931 , \52108 , \49405 );
and \g131685/U$3 ( \62932 , \49403 , \51854 );
nor \g131685/U$1 ( \62933 , \62931 , \62932 );
not \g131652/U$4 ( \62934 , \62933 );
or \g131652/U$2 ( \62935 , \62930 , \62934 );
or \g131652/U$5 ( \62936 , \62933 , \49233 );
nand \g131652/U$1 ( \62937 , \62935 , \62936 );
xor \g456094/U$2 ( \62938 , \62929 , \62937 );
not \g131289/U$3 ( \62939 , \50362 );
and \g131315/U$2 ( \62940 , \50957 , \50588 );
and \g131315/U$3 ( \62941 , \50587 , \50752 );
nor \g131315/U$1 ( \62942 , \62940 , \62941 );
not \g131289/U$4 ( \62943 , \62942 );
or \g131289/U$2 ( \62944 , \62939 , \62943 );
or \g131289/U$5 ( \62945 , \62942 , \50362 );
nand \g131289/U$1 ( \62946 , \62944 , \62945 );
xor \g456094/U$1 ( \62947 , \62938 , \62946 );
xor \g131974/U$4 ( \62948 , \62662 , \62670 );
and \g131974/U$3 ( \62949 , \62948 , \62692 );
and \g131974/U$5 ( \62950 , \62662 , \62670 );
or \g131974/U$2 ( \62951 , \62949 , \62950 );
not \g131915/U$3 ( \62952 , \48685 );
and \g131953/U$2 ( \62953 , \52978 , \48860 );
and \g131953/U$3 ( \62954 , \48858 , \52883 );
nor \g131953/U$1 ( \62955 , \62953 , \62954 );
not \g131915/U$4 ( \62956 , \62955 );
or \g131915/U$2 ( \62957 , \62952 , \62956 );
or \g131915/U$5 ( \62958 , \62955 , \48685 );
nand \g131915/U$1 ( \62959 , \62957 , \62958 );
xor \g131500/U$1 ( \62960 , \62951 , \62959 );
not \g131540/U$3 ( \62961 , \49568 );
and \g131572/U$2 ( \62962 , \51604 , \49813 );
and \g131572/U$3 ( \62963 , \49812 , \51564 );
nor \g131572/U$1 ( \62964 , \62962 , \62963 );
not \g131540/U$4 ( \62965 , \62964 );
or \g131540/U$2 ( \62966 , \62961 , \62965 );
or \g131540/U$5 ( \62967 , \62964 , \49568 );
nand \g131540/U$1 ( \62968 , \62966 , \62967 );
xor \g131500/U$1_r1 ( \62969 , \62960 , \62968 );
xor \g131053/U$4 ( \62970 , \62631 , \62635 );
and \g131053/U$3 ( \62971 , \62970 , \62644 );
and \g131053/U$5 ( \62972 , \62631 , \62635 );
or \g131053/U$2 ( \62973 , \62971 , \62972 );
xor \g456094/U$1_r1 ( \62974 , \62969 , \62973 );
xor \g456094/U$1_r2 ( \62975 , \62947 , \62974 );
xor \g130727/U$1 ( \62976 , \62904 , \62975 );
xor \g130915/U$4 ( \62977 , \62654 , \62693 );
and \g130915/U$3 ( \62978 , \62977 , \62702 );
and \g130915/U$5 ( \62979 , \62654 , \62693 );
or \g130915/U$2 ( \62980 , \62978 , \62979 );
not \g131404/U$3 ( \62981 , \49925 );
and \g131438/U$2 ( \62982 , \51117 , \50159 );
and \g131438/U$3 ( \62983 , \50160 , \51098 );
nor \g131438/U$1 ( \62984 , \62982 , \62983 );
not \g131404/U$4 ( \62985 , \62984 );
or \g131404/U$2 ( \62986 , \62981 , \62985 );
or \g131404/U$5 ( \62987 , \62984 , \49925 );
nand \g131404/U$1 ( \62988 , \62986 , \62987 );
xor \g131875/U$4 ( \62989 , \62584 , \62592 );
and \g131875/U$3 ( \62990 , \62989 , \62597 );
and \g131875/U$5 ( \62991 , \62584 , \62592 );
or \g131875/U$2 ( \62992 , \62990 , \62991 );
xor \g131129/U$1 ( \62993 , \62988 , \62992 );
not \g131175/U$3 ( \62994 , \50759 );
and \g131207/U$2 ( \62995 , \50305 , \51053 );
and \g131207/U$3 ( \62996 , \51055 , \50443 );
nor \g131207/U$1 ( \62997 , \62995 , \62996 );
not \g131175/U$4 ( \62998 , \62997 );
or \g131175/U$2 ( \62999 , \62994 , \62998 );
or \g131175/U$5 ( \63000 , \62997 , \50759 );
nand \g131175/U$1 ( \63001 , \62999 , \63000 );
xor \g131129/U$1_r1 ( \63002 , \62993 , \63001 );
xor \g130800/U$1 ( \63003 , \62980 , \63002 );
not \g131017/U$3 ( \63004 , \51124 );
and \g131073/U$2 ( \63005 , \49888 , \51517 );
and \g131073/U$3 ( \63006 , \51518 , \50019 );
nor \g131073/U$1 ( \63007 , \63005 , \63006 );
not \g131017/U$4 ( \63008 , \63007 );
or \g131017/U$2 ( \63009 , \63004 , \63008 );
or \g131017/U$5 ( \63010 , \63007 , \51124 );
nand \g131017/U$1 ( \63011 , \63009 , \63010 );
xor \g131670/U$4 ( \63012 , \62736 , \62744 );
and \g131670/U$3 ( \63013 , \63012 , \62767 );
and \g131670/U$5 ( \63014 , \62736 , \62744 );
or \g131670/U$2 ( \63015 , \63013 , \63014 );
xor \g130861/U$1 ( \63016 , \63011 , \63015 );
not \g130895/U$3 ( \63017 , \51120 );
and \g130939/U$2 ( \63018 , \49512 , \52270 );
and \g130939/U$3 ( \63019 , \52273 , \49714 );
nor \g130939/U$1 ( \63020 , \63018 , \63019 );
not \g130895/U$4 ( \63021 , \63020 );
or \g130895/U$2 ( \63022 , \63017 , \63021 );
or \g130895/U$5 ( \63023 , \63020 , \51120 );
nand \g130895/U$1 ( \63024 , \63022 , \63023 );
xor \g130861/U$1_r1 ( \63025 , \63016 , \63024 );
xor \g130800/U$1_r1 ( \63026 , \63003 , \63025 );
xor \g130727/U$1_r1 ( \63027 , \62976 , \63026 );
xor \g456082/U$1_r1 ( \63028 , \62900 , \63027 );
xor \g456082/U$1_r2 ( \63029 , \62892 , \63028 );
xor \g130604/U$1_r1 ( \63030 , \62818 , \63029 );
xor \g128801/U$1 ( \63031 , \62804 , \62800 );
and \g128800/U$2 ( \63032 , \63030 , \63031 );
not \g128799/U$1 ( \63033 , \63032 );
nand \g128798/U$1 ( \63034 , \62805 , \63033 );
xor \g130604/U$4 ( \63035 , \62809 , \62817 );
and \g130604/U$3 ( \63036 , \63035 , \63029 );
and \g130604/U$5 ( \63037 , \62809 , \62817 );
or \g130604/U$2 ( \63038 , \63036 , \63037 );
and \g128795/U$2 ( \63039 , \63034 , \63038 );
xor \g131500/U$4 ( \63040 , \62951 , \62959 );
and \g131500/U$3 ( \63041 , \63040 , \62968 );
and \g131500/U$5 ( \63042 , \62951 , \62959 );
or \g131500/U$2 ( \63043 , \63041 , \63042 );
not \g131719/U$3 ( \63044 , \49014 );
and \g131752/U$2 ( \63045 , \52108 , \49074 );
and \g131752/U$3 ( \63046 , \49075 , \52352 );
nor \g131752/U$1 ( \63047 , \63045 , \63046 );
not \g131719/U$4 ( \63048 , \63047 );
or \g131719/U$2 ( \63049 , \63044 , \63048 );
or \g131719/U$5 ( \63050 , \63047 , \49014 );
nand \g131719/U$1 ( \63051 , \63049 , \63050 );
not \g131844/U$3 ( \63052 , \48685 );
and \g131889/U$2 ( \63053 , \52620 , \48858 );
and \g131889/U$3 ( \63054 , \48860 , \52883 );
nor \g131889/U$1 ( \63055 , \63053 , \63054 );
not \g131844/U$4 ( \63056 , \63055 );
or \g131844/U$2 ( \63057 , \63052 , \63056 );
or \g131844/U$5 ( \63058 , \63055 , \48685 );
nand \g131844/U$1 ( \63059 , \63057 , \63058 );
xor \g131669/U$1 ( \63060 , \63051 , \63059 );
and \g132403/U$2 ( \63061 , \47913 , \55127 );
and \g132403/U$3 ( \63062 , \55460 , \47914 );
nor \g132403/U$1 ( \63063 , \63061 , \63062 );
and \g132321/U$2 ( \63064 , \63063 , \47977 );
not \g132321/U$4 ( \63065 , \63063 );
and \g132321/U$3 ( \63066 , \63065 , \47976 );
nor \g132321/U$1 ( \63067 , \63064 , \63066 );
not \g132472/U$3 ( \63068 , \47935 );
and \g132552/U$2 ( \63069 , \47931 , \54853 );
and \g132552/U$3 ( \63070 , \54537 , \47930 );
nor \g132552/U$1 ( \63071 , \63069 , \63070 );
not \g132472/U$4 ( \63072 , \63071 );
or \g132472/U$2 ( \63073 , \63068 , \63072 );
or \g132472/U$5 ( \63074 , \63071 , \47935 );
nand \g132472/U$1 ( \63075 , \63073 , \63074 );
xor \g132069/U$1 ( \63076 , \63067 , \63075 );
and \g132167/U$2 ( \63077 , \62906 , \62914 );
xor \g132069/U$1_r1 ( \63078 , \63076 , \63077 );
xor \g131669/U$1_r1 ( \63079 , \63060 , \63078 );
xor \g131222/U$1 ( \63080 , \63043 , \63079 );
xor \g456094/U$5 ( \63081 , \62929 , \62937 );
and \g456094/U$4 ( \63082 , \63081 , \62946 );
and \g456094/U$6 ( \63083 , \62929 , \62937 );
or \g456094/U$3 ( \63084 , \63082 , \63083 );
xor \g131222/U$1_r1 ( \63085 , \63080 , \63084 );
xor \g456118/U$9 ( \63086 , \62836 , \62844 );
xor \g456118/U$9_r1 ( \63087 , \63086 , \62849 );
and \g456118/U$8 ( \63088 , \62876 , \63087 );
xor \g456118/U$11 ( \63089 , \62836 , \62844 );
xor \g456118/U$11_r1 ( \63090 , \63089 , \62849 );
and \g456118/U$10 ( \63091 , \62880 , \63090 );
and \g456118/U$12 ( \63092 , \62876 , \62880 );
or \g456118/U$7 ( \63093 , \63088 , \63091 , \63092 );
xor \g456080/U$2 ( \63094 , \63085 , \63093 );
xor \g456094/U$9 ( \63095 , \62929 , \62937 );
xor \g456094/U$9_r1 ( \63096 , \63095 , \62946 );
and \g456094/U$8 ( \63097 , \62969 , \63096 );
xor \g456094/U$11 ( \63098 , \62929 , \62937 );
xor \g456094/U$11_r1 ( \63099 , \63098 , \62946 );
and \g456094/U$10 ( \63100 , \62973 , \63099 );
and \g456094/U$12 ( \63101 , \62969 , \62973 );
or \g456094/U$7 ( \63102 , \63097 , \63100 , \63101 );
xor \g456080/U$1 ( \63103 , \63094 , \63102 );
xor \g456082/U$5 ( \63104 , \62882 , \62886 );
and \g456082/U$4 ( \63105 , \63104 , \62891 );
and \g456082/U$6 ( \63106 , \62882 , \62886 );
or \g456082/U$3 ( \63107 , \63105 , \63106 );
xor \g130727/U$4 ( \63108 , \62904 , \62975 );
and \g130727/U$3 ( \63109 , \63108 , \63026 );
and \g130727/U$5 ( \63110 , \62904 , \62975 );
or \g130727/U$2 ( \63111 , \63109 , \63110 );
xor \g456080/U$1_r1 ( \63112 , \63107 , \63111 );
xor \g456080/U$1_r2 ( \63113 , \63103 , \63112 );
xor \g130800/U$4 ( \63114 , \62980 , \63002 );
and \g130800/U$3 ( \63115 , \63114 , \63025 );
and \g130800/U$5 ( \63116 , \62980 , \63002 );
or \g130800/U$2 ( \63117 , \63115 , \63116 );
not \g131347/U$3 ( \63118 , \49925 );
and \g131370/U$2 ( \63119 , \51117 , \50160 );
and \g131370/U$3 ( \63120 , \50159 , \50957 );
nor \g131370/U$1 ( \63121 , \63119 , \63120 );
not \g131347/U$4 ( \63122 , \63121 );
or \g131347/U$2 ( \63123 , \63118 , \63122 );
or \g131347/U$5 ( \63124 , \63121 , \49925 );
nand \g131347/U$1 ( \63125 , \63123 , \63124 );
xor \g132172/U$1 ( \63126 , \56169 , \56177 );
not \g132521/U$3 ( \63127 , \47997 );
and \g132567/U$2 ( \63128 , \48063 , \54251 );
and \g132567/U$3 ( \63129 , \54529 , \48064 );
nor \g132567/U$1 ( \63130 , \63128 , \63129 );
not \g132521/U$4 ( \63131 , \63130 );
or \g132521/U$2 ( \63132 , \63127 , \63131 );
or \g132521/U$5 ( \63133 , \63130 , \47997 );
nand \g132521/U$1 ( \63134 , \63132 , \63133 );
xor \g131982/U$1 ( \63135 , \63126 , \63134 );
xor \g132073/U$4 ( \63136 , \62825 , \62833 );
and \g132073/U$3 ( \63137 , \63136 , \62835 );
and \g132073/U$5 ( \63138 , \62825 , \62833 );
or \g132073/U$2 ( \63139 , \63137 , \63138 );
xor \g131982/U$1_r1 ( \63140 , \63135 , \63139 );
xor \g456098/U$2 ( \63141 , \63125 , \63140 );
not \g131228/U$3 ( \63142 , \50362 );
and \g131262/U$2 ( \63143 , \50752 , \50588 );
and \g131262/U$3 ( \63144 , \50587 , \50443 );
nor \g131262/U$1 ( \63145 , \63143 , \63144 );
not \g131228/U$4 ( \63146 , \63145 );
or \g131228/U$2 ( \63147 , \63142 , \63146 );
or \g131228/U$5 ( \63148 , \63145 , \50362 );
nand \g131228/U$1 ( \63149 , \63147 , \63148 );
xor \g456098/U$1 ( \63150 , \63141 , \63149 );
not \g131592/U$3 ( \63151 , \49233 );
and \g131623/U$2 ( \63152 , \51604 , \49403 );
and \g131623/U$3 ( \63153 , \49405 , \51854 );
nor \g131623/U$1 ( \63154 , \63152 , \63153 );
not \g131592/U$4 ( \63155 , \63154 );
or \g131592/U$2 ( \63156 , \63151 , \63155 );
or \g131592/U$5 ( \63157 , \63154 , \49233 );
nand \g131592/U$1 ( \63158 , \63156 , \63157 );
xor \g131983/U$4 ( \63159 , \62915 , \62923 );
and \g131983/U$3 ( \63160 , \63159 , \62928 );
and \g131983/U$5 ( \63161 , \62915 , \62923 );
or \g131983/U$2 ( \63162 , \63160 , \63161 );
xor \g131430/U$1 ( \63163 , \63158 , \63162 );
not \g131474/U$3 ( \63164 , \49568 );
and \g131504/U$2 ( \63165 , \51564 , \49813 );
and \g131504/U$3 ( \63166 , \49812 , \51098 );
nor \g131504/U$1 ( \63167 , \63165 , \63166 );
not \g131474/U$4 ( \63168 , \63167 );
or \g131474/U$2 ( \63169 , \63164 , \63168 );
or \g131474/U$5 ( \63170 , \63167 , \49568 );
nand \g131474/U$1 ( \63171 , \63169 , \63170 );
xor \g131430/U$1_r1 ( \63172 , \63163 , \63171 );
xor \g131129/U$4 ( \63173 , \62988 , \62992 );
and \g131129/U$3 ( \63174 , \63173 , \63001 );
and \g131129/U$5 ( \63175 , \62988 , \62992 );
or \g131129/U$2 ( \63176 , \63174 , \63175 );
xor \g456098/U$1_r1 ( \63177 , \63172 , \63176 );
xor \g456098/U$1_r2 ( \63178 , \63150 , \63177 );
xor \g130669/U$1 ( \63179 , \63117 , \63178 );
xor \g130861/U$4 ( \63180 , \63011 , \63015 );
and \g130861/U$3 ( \63181 , \63180 , \63024 );
and \g130861/U$5 ( \63182 , \63011 , \63015 );
or \g130861/U$2 ( \63183 , \63181 , \63182 );
xor \g456118/U$5 ( \63184 , \62836 , \62844 );
and \g456118/U$4 ( \63185 , \63184 , \62849 );
and \g456118/U$6 ( \63186 , \62836 , \62844 );
or \g456118/U$3 ( \63187 , \63185 , \63186 );
xor \g132032/U$4 ( \63188 , \62858 , \62866 );
and \g132032/U$3 ( \63189 , \63188 , \62875 );
and \g132032/U$5 ( \63190 , \62858 , \62866 );
or \g132032/U$2 ( \63191 , \63189 , \63190 );
xor \g131052/U$1 ( \63192 , \63187 , \63191 );
not \g131097/U$3 ( \63193 , \50759 );
and \g131135/U$2 ( \63194 , \50305 , \51055 );
and \g131135/U$3 ( \63195 , \51053 , \50019 );
nor \g131135/U$1 ( \63196 , \63194 , \63195 );
not \g131097/U$4 ( \63197 , \63196 );
or \g131097/U$2 ( \63198 , \63193 , \63197 );
or \g131097/U$5 ( \63199 , \63196 , \50759 );
nand \g131097/U$1 ( \63200 , \63198 , \63199 );
xor \g131052/U$1_r1 ( \63201 , \63192 , \63200 );
xor \g130746/U$1 ( \63202 , \63183 , \63201 );
not \g130952/U$3 ( \63203 , \51124 );
and \g130994/U$2 ( \63204 , \49888 , \51518 );
and \g130994/U$3 ( \63205 , \51517 , \49714 );
nor \g130994/U$1 ( \63206 , \63204 , \63205 );
not \g130952/U$4 ( \63207 , \63206 );
or \g130952/U$2 ( \63208 , \63203 , \63207 );
or \g130952/U$5 ( \63209 , \63206 , \51124 );
nand \g130952/U$1 ( \63210 , \63208 , \63209 );
not \g132156/U$3 ( \63211 , \48323 );
and \g132192/U$2 ( \63212 , \53610 , \48334 );
and \g132192/U$3 ( \63213 , \48335 , \53848 );
nor \g132192/U$1 ( \63214 , \63212 , \63213 );
not \g132156/U$4 ( \63215 , \63214 );
or \g132156/U$2 ( \63216 , \63211 , \63215 );
or \g132156/U$5 ( \63217 , \63214 , \48323 );
nand \g132156/U$1 ( \63218 , \63216 , \63217 );
not \g132322/U$3 ( \63219 , \48159 );
and \g132404/U$2 ( \63220 , \54185 , \48155 );
and \g132404/U$3 ( \63221 , \48154 , \54015 );
nor \g132404/U$1 ( \63222 , \63220 , \63221 );
not \g132322/U$4 ( \63223 , \63222 );
or \g132322/U$2 ( \63224 , \63219 , \63223 );
or \g132322/U$5 ( \63225 , \63222 , \48159 );
nand \g132322/U$1 ( \63226 , \63224 , \63225 );
xor \g131950/U$1 ( \63227 , \63218 , \63226 );
not \g131999/U$3 ( \63228 , \48483 );
and \g132039/U$2 ( \63229 , \52978 , \48478 );
and \g132039/U$3 ( \63230 , \48479 , \53300 );
nor \g132039/U$1 ( \63231 , \63229 , \63230 );
not \g131999/U$4 ( \63232 , \63231 );
or \g131999/U$2 ( \63233 , \63228 , \63232 );
or \g131999/U$5 ( \63234 , \63231 , \48483 );
nand \g131999/U$1 ( \63235 , \63233 , \63234 );
xor \g131950/U$1_r1 ( \63236 , \63227 , \63235 );
xor \g130805/U$1 ( \63237 , \63210 , \63236 );
not \g130841/U$3 ( \63238 , \51120 );
and \g130881/U$2 ( \63239 , \49512 , \52273 );
and \g130881/U$3 ( \63240 , \52270 , \49282 );
nor \g130881/U$1 ( \63241 , \63239 , \63240 );
not \g130841/U$4 ( \63242 , \63241 );
or \g130841/U$2 ( \63243 , \63238 , \63242 );
or \g130841/U$5 ( \63244 , \63241 , \51120 );
nand \g130841/U$1 ( \63245 , \63243 , \63244 );
xor \g130805/U$1_r1 ( \63246 , \63237 , \63245 );
xor \g130746/U$1_r1 ( \63247 , \63202 , \63246 );
xor \g130669/U$1_r1 ( \63248 , \63179 , \63247 );
xor \g456076/U$1 ( \63249 , \63113 , \63248 );
xor \g456082/U$9 ( \63250 , \62882 , \62886 );
xor \g456082/U$9_r1 ( \63251 , \63250 , \62891 );
and \g456082/U$8 ( \63252 , \62900 , \63251 );
xor \g456082/U$11 ( \63253 , \62882 , \62886 );
xor \g456082/U$11_r1 ( \63254 , \63253 , \62891 );
and \g456082/U$10 ( \63255 , \63027 , \63254 );
and \g456082/U$12 ( \63256 , \62900 , \63027 );
or \g456082/U$7 ( \63257 , \63252 , \63255 , \63256 );
xor \g456076/U$1_r1 ( \63258 , \63249 , \63257 );
xor \g128797/U$1 ( \63259 , \63038 , \63034 );
and \g128796/U$2 ( \63260 , \63258 , \63259 );
nor \g128795/U$1 ( \63261 , \63039 , \63260 );
xor \g456076/U$4 ( \63262 , \63113 , \63248 );
and \g456076/U$3 ( \63263 , \63262 , \63257 );
and \g456076/U$5 ( \63264 , \63113 , \63248 );
nor \g456076/U$2 ( \63265 , \63263 , \63264 );
or \g128790/U$2 ( \63266 , \63261 , \63265 );
xnor \g128794/U$1 ( \63267 , \63265 , \63261 );
not \g128793/U$2 ( \63268 , \63267 );
xor \g130746/U$4 ( \63269 , \63183 , \63201 );
and \g130746/U$3 ( \63270 , \63269 , \63246 );
and \g130746/U$5 ( \63271 , \63183 , \63201 );
or \g130746/U$2 ( \63272 , \63270 , \63271 );
not \g132473/U$3 ( \63273 , \47935 );
and \g132538/U$2 ( \63274 , \47931 , \54537 );
and \g132538/U$3 ( \63275 , \54529 , \47930 );
nor \g132538/U$1 ( \63276 , \63274 , \63275 );
not \g132473/U$4 ( \63277 , \63276 );
or \g132473/U$2 ( \63278 , \63273 , \63277 );
or \g132473/U$5 ( \63279 , \63276 , \47935 );
nand \g132473/U$1 ( \63280 , \63278 , \63279 );
not \g132444/U$3 ( \63281 , \47997 );
and \g132491/U$2 ( \63282 , \54185 , \48063 );
and \g132491/U$3 ( \63283 , \54251 , \48064 );
nor \g132491/U$1 ( \63284 , \63282 , \63283 );
not \g132444/U$4 ( \63285 , \63284 );
or \g132444/U$2 ( \63286 , \63281 , \63285 );
or \g132444/U$5 ( \63287 , \63284 , \47997 );
nand \g132444/U$1 ( \63288 , \63286 , \63287 );
xor \g131980/U$1 ( \63289 , \63280 , \63288 );
xor \g132069/U$4 ( \63290 , \63067 , \63075 );
and \g132069/U$3 ( \63291 , \63290 , \63077 );
and \g132069/U$5 ( \63292 , \63067 , \63075 );
or \g132069/U$2 ( \63293 , \63291 , \63292 );
xor \g131980/U$1_r1 ( \63294 , \63289 , \63293 );
xor \g131950/U$4 ( \63295 , \63218 , \63226 );
and \g131950/U$3 ( \63296 , \63295 , \63235 );
and \g131950/U$5 ( \63297 , \63218 , \63226 );
or \g131950/U$2 ( \63298 , \63296 , \63297 );
xor \g456095/U$2 ( \63299 , \63294 , \63298 );
not \g131174/U$3 ( \63300 , \50362 );
and \g131206/U$2 ( \63301 , \50305 , \50587 );
and \g131206/U$3 ( \63302 , \50588 , \50443 );
nor \g131206/U$1 ( \63303 , \63301 , \63302 );
not \g131174/U$4 ( \63304 , \63303 );
or \g131174/U$2 ( \63305 , \63300 , \63304 );
or \g131174/U$5 ( \63306 , \63303 , \50362 );
nand \g131174/U$1 ( \63307 , \63305 , \63306 );
xor \g456095/U$1 ( \63308 , \63299 , \63307 );
not \g131539/U$3 ( \63309 , \49233 );
and \g131571/U$2 ( \63310 , \51604 , \49405 );
and \g131571/U$3 ( \63311 , \49403 , \51564 );
nor \g131571/U$1 ( \63312 , \63310 , \63311 );
not \g131539/U$4 ( \63313 , \63312 );
or \g131539/U$2 ( \63314 , \63309 , \63313 );
or \g131539/U$5 ( \63315 , \63312 , \49233 );
nand \g131539/U$1 ( \63316 , \63314 , \63315 );
xor \g131982/U$4 ( \63317 , \63126 , \63134 );
and \g131982/U$3 ( \63318 , \63317 , \63139 );
and \g131982/U$5 ( \63319 , \63126 , \63134 );
or \g131982/U$2 ( \63320 , \63318 , \63319 );
xor \g131253/U$1 ( \63321 , \63316 , \63320 );
not \g131288/U$3 ( \63322 , \49925 );
and \g131314/U$2 ( \63323 , \50957 , \50160 );
and \g131314/U$3 ( \63324 , \50159 , \50752 );
nor \g131314/U$1 ( \63325 , \63323 , \63324 );
not \g131288/U$4 ( \63326 , \63325 );
or \g131288/U$2 ( \63327 , \63322 , \63326 );
or \g131288/U$5 ( \63328 , \63325 , \49925 );
nand \g131288/U$1 ( \63329 , \63327 , \63328 );
xor \g131253/U$1_r1 ( \63330 , \63321 , \63329 );
xor \g131052/U$4 ( \63331 , \63187 , \63191 );
and \g131052/U$3 ( \63332 , \63331 , \63200 );
and \g131052/U$5 ( \63333 , \63187 , \63191 );
or \g131052/U$2 ( \63334 , \63332 , \63333 );
xor \g456095/U$1_r1 ( \63335 , \63330 , \63334 );
xor \g456095/U$1_r2 ( \63336 , \63308 , \63335 );
xor \g456068/U$2 ( \63337 , \63272 , \63336 );
xor \g130805/U$4 ( \63338 , \63210 , \63236 );
and \g130805/U$3 ( \63339 , \63338 , \63245 );
and \g130805/U$5 ( \63340 , \63210 , \63236 );
or \g130805/U$2 ( \63341 , \63339 , \63340 );
xor \g131669/U$4 ( \63342 , \63051 , \63059 );
and \g131669/U$3 ( \63343 , \63342 , \63078 );
and \g131669/U$5 ( \63344 , \63051 , \63059 );
or \g131669/U$2 ( \63345 , \63343 , \63344 );
not \g132077/U$3 ( \63346 , \48323 );
and \g132119/U$2 ( \63347 , \53610 , \48335 );
and \g132119/U$3 ( \63348 , \48334 , \53300 );
nor \g132119/U$1 ( \63349 , \63347 , \63348 );
not \g132077/U$4 ( \63350 , \63349 );
or \g132077/U$2 ( \63351 , \63346 , \63350 );
or \g132077/U$5 ( \63352 , \63349 , \48323 );
nand \g132077/U$1 ( \63353 , \63351 , \63352 );
not \g132243/U$3 ( \63354 , \48159 );
and \g132303/U$2 ( \63355 , \53848 , \48154 );
and \g132303/U$3 ( \63356 , \48155 , \54015 );
nor \g132303/U$1 ( \63357 , \63355 , \63356 );
not \g132243/U$4 ( \63358 , \63357 );
or \g132243/U$2 ( \63359 , \63354 , \63358 );
or \g132243/U$5 ( \63360 , \63357 , \48159 );
nand \g132243/U$1 ( \63361 , \63359 , \63360 );
xor \g131748/U$1 ( \63362 , \63353 , \63361 );
not \g131778/U$3 ( \63363 , \48685 );
and \g131811/U$2 ( \63364 , \52620 , \48860 );
and \g131811/U$3 ( \63365 , \48858 , \52352 );
nor \g131811/U$1 ( \63366 , \63364 , \63365 );
not \g131778/U$4 ( \63367 , \63366 );
or \g131778/U$2 ( \63368 , \63363 , \63367 );
or \g131778/U$5 ( \63369 , \63366 , \48685 );
nand \g131778/U$1 ( \63370 , \63368 , \63369 );
xor \g131748/U$1_r1 ( \63371 , \63362 , \63370 );
xor \g130976/U$1 ( \63372 , \63345 , \63371 );
not \g131016/U$3 ( \63373 , \50759 );
and \g131059/U$2 ( \63374 , \49888 , \51053 );
and \g131059/U$3 ( \63375 , \51055 , \50019 );
nor \g131059/U$1 ( \63376 , \63374 , \63375 );
not \g131016/U$4 ( \63377 , \63376 );
or \g131016/U$2 ( \63378 , \63373 , \63377 );
or \g131016/U$5 ( \63379 , \63376 , \50759 );
nand \g131016/U$1 ( \63380 , \63378 , \63379 );
xor \g130976/U$1_r1 ( \63381 , \63372 , \63380 );
xor \g130715/U$1 ( \63382 , \63341 , \63381 );
not \g130894/U$3 ( \63383 , \51124 );
and \g130938/U$2 ( \63384 , \49512 , \51517 );
and \g130938/U$3 ( \63385 , \51518 , \49714 );
nor \g130938/U$1 ( \63386 , \63384 , \63385 );
not \g130894/U$4 ( \63387 , \63386 );
or \g130894/U$2 ( \63388 , \63383 , \63387 );
or \g130894/U$5 ( \63389 , \63386 , \51124 );
nand \g130894/U$1 ( \63390 , \63388 , \63389 );
not \g131403/U$3 ( \63391 , \49568 );
and \g131437/U$2 ( \63392 , \51117 , \49812 );
and \g131437/U$3 ( \63393 , \49813 , \51098 );
nor \g131437/U$1 ( \63394 , \63392 , \63393 );
not \g131403/U$4 ( \63395 , \63394 );
or \g131403/U$2 ( \63396 , \63391 , \63395 );
or \g131403/U$5 ( \63397 , \63394 , \49568 );
nand \g131403/U$1 ( \63398 , \63396 , \63397 );
xor \g130749/U$1 ( \63399 , \63390 , \63398 );
not \g130782/U$3 ( \63400 , \51120 );
and \g130827/U$2 ( \63401 , \49282 , \52273 );
and \g130827/U$3 ( \63402 , \52270 , \49158 );
nor \g130827/U$1 ( \63403 , \63401 , \63402 );
not \g130782/U$4 ( \63404 , \63403 );
or \g130782/U$2 ( \63405 , \63400 , \63404 );
or \g130782/U$5 ( \63406 , \63403 , \51120 );
nand \g130782/U$1 ( \63407 , \63405 , \63406 );
xor \g130749/U$1_r1 ( \63408 , \63399 , \63407 );
xor \g130715/U$1_r1 ( \63409 , \63382 , \63408 );
xor \g456068/U$1 ( \63410 , \63337 , \63409 );
xor \g456080/U$9 ( \63411 , \63085 , \63093 );
xor \g456080/U$9_r1 ( \63412 , \63411 , \63102 );
and \g456080/U$8 ( \63413 , \63107 , \63412 );
xor \g456080/U$11 ( \63414 , \63085 , \63093 );
xor \g456080/U$11_r1 ( \63415 , \63414 , \63102 );
and \g456080/U$10 ( \63416 , \63111 , \63415 );
and \g456080/U$12 ( \63417 , \63107 , \63111 );
or \g456080/U$7 ( \63418 , \63413 , \63416 , \63417 );
xor \g456080/U$5 ( \63419 , \63085 , \63093 );
and \g456080/U$4 ( \63420 , \63419 , \63102 );
and \g456080/U$6 ( \63421 , \63085 , \63093 );
or \g456080/U$3 ( \63422 , \63420 , \63421 );
xor \g131430/U$4 ( \63423 , \63158 , \63162 );
and \g131430/U$3 ( \63424 , \63423 , \63171 );
and \g131430/U$5 ( \63425 , \63158 , \63162 );
or \g131430/U$2 ( \63426 , \63424 , \63425 );
xor \g456134/U$2 ( \63427 , \56164 , \56165 );
xor \g456134/U$1 ( \63428 , \63427 , \56178 );
not \g131914/U$3 ( \63429 , \48483 );
and \g131957/U$2 ( \63430 , \52978 , \48479 );
and \g131957/U$3 ( \63431 , \48478 , \52883 );
nor \g131957/U$1 ( \63432 , \63430 , \63431 );
not \g131914/U$4 ( \63433 , \63432 );
or \g131914/U$2 ( \63434 , \63429 , \63433 );
or \g131914/U$5 ( \63435 , \63432 , \48483 );
nand \g131914/U$1 ( \63436 , \63434 , \63435 );
not \g131650/U$3 ( \63437 , \49014 );
and \g131684/U$2 ( \63438 , \52108 , \49075 );
and \g131684/U$3 ( \63439 , \49074 , \51854 );
nor \g131684/U$1 ( \63440 , \63438 , \63439 );
not \g131650/U$4 ( \63441 , \63440 );
or \g131650/U$2 ( \63442 , \63437 , \63441 );
or \g131650/U$5 ( \63443 , \63440 , \49014 );
nand \g131650/U$1 ( \63444 , \63442 , \63443 );
xor \g456134/U$1_r1 ( \63445 , \63436 , \63444 );
xor \g456134/U$1_r2 ( \63446 , \63428 , \63445 );
xor \g456093/U$2 ( \63447 , \63426 , \63446 );
xor \g456098/U$5 ( \63448 , \63125 , \63140 );
and \g456098/U$4 ( \63449 , \63448 , \63149 );
and \g456098/U$6 ( \63450 , \63125 , \63140 );
or \g456098/U$3 ( \63451 , \63449 , \63450 );
xor \g456093/U$1 ( \63452 , \63447 , \63451 );
xor \g131222/U$4 ( \63453 , \63043 , \63079 );
and \g131222/U$3 ( \63454 , \63453 , \63084 );
and \g131222/U$5 ( \63455 , \63043 , \63079 );
or \g131222/U$2 ( \63456 , \63454 , \63455 );
xor \g456098/U$9 ( \63457 , \63125 , \63140 );
xor \g456098/U$9_r1 ( \63458 , \63457 , \63149 );
and \g456098/U$8 ( \63459 , \63172 , \63458 );
xor \g456098/U$11 ( \63460 , \63125 , \63140 );
xor \g456098/U$11_r1 ( \63461 , \63460 , \63149 );
and \g456098/U$10 ( \63462 , \63176 , \63461 );
and \g456098/U$12 ( \63463 , \63172 , \63176 );
or \g456098/U$7 ( \63464 , \63459 , \63462 , \63463 );
xor \g456093/U$1_r1 ( \63465 , \63456 , \63464 );
xor \g456093/U$1_r2 ( \63466 , \63452 , \63465 );
xor \g130592/U$1 ( \63467 , \63422 , \63466 );
xor \g130669/U$4 ( \63468 , \63117 , \63178 );
and \g130669/U$3 ( \63469 , \63468 , \63247 );
and \g130669/U$5 ( \63470 , \63117 , \63178 );
or \g130669/U$2 ( \63471 , \63469 , \63470 );
xor \g130592/U$1_r1 ( \63472 , \63467 , \63471 );
xor \g456068/U$1_r1 ( \63473 , \63418 , \63472 );
xor \g456068/U$1_r2 ( \63474 , \63410 , \63473 );
nand \g128793/U$1 ( \63475 , \63268 , \63474 );
nand \g128790/U$1 ( \63476 , \63266 , \63475 );
xor \g456068/U$9 ( \63477 , \63272 , \63336 );
xor \g456068/U$9_r1 ( \63478 , \63477 , \63409 );
and \g456068/U$8 ( \63479 , \63418 , \63478 );
xor \g456068/U$11 ( \63480 , \63272 , \63336 );
xor \g456068/U$11_r1 ( \63481 , \63480 , \63409 );
and \g456068/U$10 ( \63482 , \63472 , \63481 );
and \g456068/U$12 ( \63483 , \63418 , \63472 );
or \g456068/U$7 ( \63484 , \63479 , \63482 , \63483 );
and \g128784/U$2 ( \63485 , \63476 , \63484 );
xor \g130976/U$4 ( \63486 , \63345 , \63371 );
and \g130976/U$3 ( \63487 , \63486 , \63380 );
and \g130976/U$5 ( \63488 , \63345 , \63371 );
or \g130976/U$2 ( \63489 , \63487 , \63488 );
not \g131346/U$3 ( \63490 , \49568 );
and \g131369/U$2 ( \63491 , \51117 , \49813 );
and \g131369/U$3 ( \63492 , \49812 , \50957 );
nor \g131369/U$1 ( \63493 , \63491 , \63492 );
not \g131346/U$4 ( \63494 , \63493 );
or \g131346/U$2 ( \63495 , \63490 , \63494 );
or \g131346/U$5 ( \63496 , \63493 , \49568 );
nand \g131346/U$1 ( \63497 , \63495 , \63496 );
xor \g132099/U$1 ( \63498 , \56087 , \56095 );
xor \g132099/U$1_r1 ( \63499 , \63498 , \56104 );
xor \g131049/U$1 ( \63500 , \63497 , \63499 );
not \g131096/U$3 ( \63501 , \50362 );
and \g131134/U$2 ( \63502 , \50305 , \50588 );
and \g131134/U$3 ( \63503 , \50587 , \50019 );
nor \g131134/U$1 ( \63504 , \63502 , \63503 );
not \g131096/U$4 ( \63505 , \63504 );
or \g131096/U$2 ( \63506 , \63501 , \63505 );
or \g131096/U$5 ( \63507 , \63504 , \50362 );
nand \g131096/U$1 ( \63508 , \63506 , \63507 );
xor \g131049/U$1_r1 ( \63509 , \63500 , \63508 );
xor \g130690/U$1 ( \63510 , \63489 , \63509 );
xor \g130749/U$4 ( \63511 , \63390 , \63398 );
and \g130749/U$3 ( \63512 , \63511 , \63407 );
and \g130749/U$5 ( \63513 , \63390 , \63398 );
or \g130749/U$2 ( \63514 , \63512 , \63513 );
xor \g130690/U$1_r1 ( \63515 , \63510 , \63514 );
xor \g130715/U$4 ( \63516 , \63341 , \63381 );
and \g130715/U$3 ( \63517 , \63516 , \63408 );
and \g130715/U$5 ( \63518 , \63341 , \63381 );
or \g130715/U$2 ( \63519 , \63517 , \63518 );
xor \g456066/U$2 ( \63520 , \63515 , \63519 );
xor \g456134/U$9 ( \63521 , \56164 , \56165 );
xor \g456134/U$9_r1 ( \63522 , \63521 , \56178 );
and \g456134/U$8 ( \63523 , \63436 , \63522 );
xor \g456134/U$11 ( \63524 , \56164 , \56165 );
xor \g456134/U$11_r1 ( \63525 , \63524 , \56178 );
and \g456134/U$10 ( \63526 , \63444 , \63525 );
and \g456134/U$12 ( \63527 , \63436 , \63444 );
or \g456134/U$7 ( \63528 , \63523 , \63526 , \63527 );
xor \g131668/U$1 ( \63529 , \56181 , \56189 );
xor \g131668/U$1_r1 ( \63530 , \63529 , \56198 );
xor \g456079/U$2 ( \63531 , \63528 , \63530 );
not \g130951/U$3 ( \63532 , \50759 );
and \g130980/U$2 ( \63533 , \49888 , \51055 );
and \g130980/U$3 ( \63534 , \51053 , \49714 );
nor \g130980/U$1 ( \63535 , \63533 , \63534 );
not \g130951/U$4 ( \63536 , \63535 );
or \g130951/U$2 ( \63537 , \63532 , \63536 );
or \g130951/U$5 ( \63538 , \63535 , \50759 );
nand \g130951/U$1 ( \63539 , \63537 , \63538 );
xor \g456079/U$1 ( \63540 , \63531 , \63539 );
xor \g131980/U$4 ( \63541 , \63280 , \63288 );
and \g131980/U$3 ( \63542 , \63541 , \63293 );
and \g131980/U$5 ( \63543 , \63280 , \63288 );
or \g131980/U$2 ( \63544 , \63542 , \63543 );
xor \g132145/U$1 ( \63545 , \55883 , \55894 );
xor \g132145/U$1_r1 ( \63546 , \63545 , \55903 );
xor \g131201/U$1 ( \63547 , \63544 , \63546 );
not \g131227/U$3 ( \63548 , \49925 );
and \g131261/U$2 ( \63549 , \50752 , \50160 );
and \g131261/U$3 ( \63550 , \50159 , \50443 );
nor \g131261/U$1 ( \63551 , \63549 , \63550 );
not \g131227/U$4 ( \63552 , \63551 );
or \g131227/U$2 ( \63553 , \63548 , \63552 );
or \g131227/U$5 ( \63554 , \63551 , \49925 );
nand \g131227/U$1 ( \63555 , \63553 , \63554 );
xor \g131201/U$1_r1 ( \63556 , \63547 , \63555 );
not \g130840/U$3 ( \63557 , \51124 );
and \g130880/U$2 ( \63558 , \49512 , \51518 );
and \g130880/U$3 ( \63559 , \51517 , \49282 );
nor \g130880/U$1 ( \63560 , \63558 , \63559 );
not \g130840/U$4 ( \63561 , \63560 );
or \g130840/U$2 ( \63562 , \63557 , \63561 );
or \g130840/U$5 ( \63563 , \63560 , \51124 );
nand \g130840/U$1 ( \63564 , \63562 , \63563 );
xor \g131748/U$4 ( \63565 , \63353 , \63361 );
and \g131748/U$3 ( \63566 , \63565 , \63370 );
and \g131748/U$5 ( \63567 , \63353 , \63361 );
or \g131748/U$2 ( \63568 , \63566 , \63567 );
xor \g130696/U$1 ( \63569 , \63564 , \63568 );
not \g130728/U$3 ( \63570 , \51120 );
and \g130769/U$2 ( \63571 , \49102 , \52270 );
and \g130769/U$3 ( \63572 , \52273 , \49158 );
nor \g130769/U$1 ( \63573 , \63571 , \63572 );
not \g130728/U$4 ( \63574 , \63573 );
or \g130728/U$2 ( \63575 , \63570 , \63574 );
or \g130728/U$5 ( \63576 , \63573 , \51120 );
nand \g130728/U$1 ( \63577 , \63575 , \63576 );
xor \g130696/U$1_r1 ( \63578 , \63569 , \63577 );
xor \g456079/U$1_r1 ( \63579 , \63556 , \63578 );
xor \g456079/U$1_r2 ( \63580 , \63540 , \63579 );
xor \g456066/U$1 ( \63581 , \63520 , \63580 );
xor \g130592/U$4 ( \63582 , \63422 , \63466 );
and \g130592/U$3 ( \63583 , \63582 , \63471 );
and \g130592/U$5 ( \63584 , \63422 , \63466 );
or \g130592/U$2 ( \63585 , \63583 , \63584 );
xor \g131253/U$4 ( \63586 , \63316 , \63320 );
and \g131253/U$3 ( \63587 , \63586 , \63329 );
and \g131253/U$5 ( \63588 , \63316 , \63320 );
or \g131253/U$2 ( \63589 , \63587 , \63588 );
xor \g131428/U$1 ( \63590 , \56225 , \56233 );
xor \g131428/U$1_r1 ( \63591 , \63590 , \56242 );
xor \g131036/U$1 ( \63592 , \63589 , \63591 );
xor \g456095/U$5 ( \63593 , \63294 , \63298 );
and \g456095/U$4 ( \63594 , \63593 , \63307 );
and \g456095/U$6 ( \63595 , \63294 , \63298 );
or \g456095/U$3 ( \63596 , \63594 , \63595 );
xor \g131036/U$1_r1 ( \63597 , \63592 , \63596 );
xor \g456093/U$5 ( \63598 , \63426 , \63446 );
and \g456093/U$4 ( \63599 , \63598 , \63451 );
and \g456093/U$6 ( \63600 , \63426 , \63446 );
or \g456093/U$3 ( \63601 , \63599 , \63600 );
xor \g456075/U$2 ( \63602 , \63597 , \63601 );
xor \g456095/U$9 ( \63603 , \63294 , \63298 );
xor \g456095/U$9_r1 ( \63604 , \63603 , \63307 );
and \g456095/U$8 ( \63605 , \63330 , \63604 );
xor \g456095/U$11 ( \63606 , \63294 , \63298 );
xor \g456095/U$11_r1 ( \63607 , \63606 , \63307 );
and \g456095/U$10 ( \63608 , \63334 , \63607 );
and \g456095/U$12 ( \63609 , \63330 , \63334 );
or \g456095/U$7 ( \63610 , \63605 , \63608 , \63609 );
xor \g456075/U$1 ( \63611 , \63602 , \63610 );
xor \g456093/U$9 ( \63612 , \63426 , \63446 );
xor \g456093/U$9_r1 ( \63613 , \63612 , \63451 );
and \g456093/U$8 ( \63614 , \63456 , \63613 );
xor \g456093/U$11 ( \63615 , \63426 , \63446 );
xor \g456093/U$11_r1 ( \63616 , \63615 , \63451 );
and \g456093/U$10 ( \63617 , \63464 , \63616 );
and \g456093/U$12 ( \63618 , \63456 , \63464 );
or \g456093/U$7 ( \63619 , \63614 , \63617 , \63618 );
xor \g456068/U$5 ( \63620 , \63272 , \63336 );
and \g456068/U$4 ( \63621 , \63620 , \63409 );
and \g456068/U$6 ( \63622 , \63272 , \63336 );
or \g456068/U$3 ( \63623 , \63621 , \63622 );
xor \g456075/U$1_r1 ( \63624 , \63619 , \63623 );
xor \g456075/U$1_r2 ( \63625 , \63611 , \63624 );
xor \g456066/U$1_r1 ( \63626 , \63585 , \63625 );
xor \g456066/U$1_r2 ( \63627 , \63581 , \63626 );
xor \g128789/U$1 ( \63628 , \63484 , \63476 );
and \g128784/U$3 ( \63629 , \63627 , \63628 );
nor \g128784/U$1 ( \63630 , \63485 , \63629 );
xor \g456075/U$9 ( \63631 , \63597 , \63601 );
xor \g456075/U$9_r1 ( \63632 , \63631 , \63610 );
and \g456075/U$8 ( \63633 , \63619 , \63632 );
xor \g456075/U$11 ( \63634 , \63597 , \63601 );
xor \g456075/U$11_r1 ( \63635 , \63634 , \63610 );
and \g456075/U$10 ( \63636 , \63623 , \63635 );
and \g456075/U$12 ( \63637 , \63619 , \63623 );
or \g456075/U$7 ( \63638 , \63633 , \63636 , \63637 );
xor \g131201/U$4 ( \63639 , \63544 , \63546 );
and \g131201/U$3 ( \63640 , \63639 , \63555 );
and \g131201/U$5 ( \63641 , \63544 , \63546 );
or \g131201/U$2 ( \63642 , \63640 , \63641 );
xor \g131498/U$1 ( \63643 , \55818 , \55820 );
xor \g131498/U$1_r1 ( \63644 , \63643 , \55829 );
xor \g130968/U$1 ( \63645 , \63642 , \63644 );
xor \g131049/U$4 ( \63646 , \63497 , \63499 );
and \g131049/U$3 ( \63647 , \63646 , \63508 );
and \g131049/U$5 ( \63648 , \63497 , \63499 );
or \g131049/U$2 ( \63649 , \63647 , \63648 );
xor \g130968/U$1_r1 ( \63650 , \63645 , \63649 );
xor \g131036/U$4 ( \63651 , \63589 , \63591 );
and \g131036/U$3 ( \63652 , \63651 , \63596 );
and \g131036/U$5 ( \63653 , \63589 , \63591 );
or \g131036/U$2 ( \63654 , \63652 , \63653 );
xor \g456070/U$2 ( \63655 , \63650 , \63654 );
xor \g130690/U$4 ( \63656 , \63489 , \63509 );
and \g130690/U$3 ( \63657 , \63656 , \63514 );
and \g130690/U$5 ( \63658 , \63489 , \63509 );
or \g130690/U$2 ( \63659 , \63657 , \63658 );
xor \g456070/U$1 ( \63660 , \63655 , \63659 );
xor \g456075/U$5 ( \63661 , \63597 , \63601 );
and \g456075/U$4 ( \63662 , \63661 , \63610 );
and \g456075/U$6 ( \63663 , \63597 , \63601 );
or \g456075/U$3 ( \63664 , \63662 , \63663 );
xor \g456066/U$5 ( \63665 , \63515 , \63519 );
and \g456066/U$4 ( \63666 , \63665 , \63580 );
and \g456066/U$6 ( \63667 , \63515 , \63519 );
or \g456066/U$3 ( \63668 , \63666 , \63667 );
xor \g456070/U$1_r1 ( \63669 , \63664 , \63668 );
xor \g456070/U$1_r2 ( \63670 , \63660 , \63669 );
xnor \g130469/U$1 ( \63671 , \63638 , \63670 );
not \g130428/U$3 ( \63672 , \63671 );
xor \g456079/U$5 ( \63673 , \63528 , \63530 );
and \g456079/U$4 ( \63674 , \63673 , \63539 );
and \g456079/U$6 ( \63675 , \63528 , \63530 );
or \g456079/U$3 ( \63676 , \63674 , \63675 );
xor \g131127/U$1 ( \63677 , \56079 , \56107 );
xor \g131127/U$1_r1 ( \63678 , \63677 , \56116 );
xor \g456069/U$2 ( \63679 , \63676 , \63678 );
xor \g130696/U$4 ( \63680 , \63564 , \63568 );
and \g130696/U$3 ( \63681 , \63680 , \63577 );
and \g130696/U$5 ( \63682 , \63564 , \63568 );
or \g130696/U$2 ( \63683 , \63681 , \63682 );
xor \g456069/U$1 ( \63684 , \63679 , \63683 );
xor \g456079/U$9 ( \63685 , \63528 , \63530 );
xor \g456079/U$9_r1 ( \63686 , \63685 , \63539 );
and \g456079/U$8 ( \63687 , \63556 , \63686 );
xor \g456079/U$11 ( \63688 , \63528 , \63530 );
xor \g456079/U$11_r1 ( \63689 , \63688 , \63539 );
and \g456079/U$10 ( \63690 , \63578 , \63689 );
and \g456079/U$12 ( \63691 , \63556 , \63578 );
or \g456079/U$7 ( \63692 , \63687 , \63690 , \63691 );
xor \g456073/U$2 ( \63693 , \56156 , \56201 );
xor \g456073/U$1 ( \63694 , \63693 , \56210 );
xor \g456092/U$1 ( \63695 , \56217 , \56245 );
xor \g456092/U$1_r1 ( \63696 , \63695 , \56254 );
xor \g130634/U$1 ( \63697 , \56268 , \56276 );
xor \g130634/U$1_r1 ( \63698 , \63697 , \56285 );
xor \g456073/U$1_r1 ( \63699 , \63696 , \63698 );
xor \g456073/U$1_r2 ( \63700 , \63694 , \63699 );
xor \g456069/U$1_r1 ( \63701 , \63692 , \63700 );
xor \g456069/U$1_r2 ( \63702 , \63684 , \63701 );
not \g130428/U$4 ( \63703 , \63702 );
and \g130428/U$2 ( \63704 , \63672 , \63703 );
and \g130428/U$5 ( \63705 , \63671 , \63702 );
nor \g130428/U$1 ( \63706 , \63704 , \63705 );
or \g128780/U$2 ( \63707 , \63630 , \63706 );
xor \g456066/U$9 ( \63708 , \63515 , \63519 );
xor \g456066/U$9_r1 ( \63709 , \63708 , \63580 );
and \g456066/U$8 ( \63710 , \63585 , \63709 );
xor \g456066/U$11 ( \63711 , \63515 , \63519 );
xor \g456066/U$11_r1 ( \63712 , \63711 , \63580 );
and \g456066/U$10 ( \63713 , \63625 , \63712 );
and \g456066/U$12 ( \63714 , \63585 , \63625 );
or \g456066/U$7 ( \63715 , \63710 , \63713 , \63714 );
xor \g128783/U$1 ( \63716 , \63706 , \63630 );
and \g128782/U$2 ( \63717 , \63715 , \63716 );
not \g128781/U$1 ( \63718 , \63717 );
nand \g128780/U$1 ( \63719 , \63707 , \63718 );
not \g130454/U$3 ( \63720 , \63638 );
not \g130454/U$4 ( \63721 , \63702 );
or \g130454/U$2 ( \63722 , \63720 , \63721 );
or \g130466/U$2 ( \63723 , \63702 , \63638 );
nand \g130466/U$1 ( \63724 , \63723 , \63670 );
nand \g130454/U$1 ( \63725 , \63722 , \63724 );
and \g128776/U$2 ( \63726 , \63719 , \63725 );
not \g130570/U$3 ( \63727 , \56214 );
not \g130603/U$3 ( \63728 , \56257 );
not \g130603/U$4 ( \63729 , \56288 );
or \g130603/U$2 ( \63730 , \63728 , \63729 );
or \g130603/U$5 ( \63731 , \56288 , \56257 );
nand \g130603/U$1 ( \63732 , \63730 , \63731 );
not \g130570/U$4 ( \63733 , \63732 );
or \g130570/U$2 ( \63734 , \63727 , \63733 );
or \g130570/U$5 ( \63735 , \63732 , \56214 );
nand \g130570/U$1 ( \63736 , \63734 , \63735 );
xor \g456073/U$9 ( \63737 , \56156 , \56201 );
xor \g456073/U$9_r1 ( \63738 , \63737 , \56210 );
and \g456073/U$8 ( \63739 , \63696 , \63738 );
xor \g456073/U$11 ( \63740 , \56156 , \56201 );
xor \g456073/U$11_r1 ( \63741 , \63740 , \56210 );
and \g456073/U$10 ( \63742 , \63698 , \63741 );
and \g456073/U$12 ( \63743 , \63696 , \63698 );
or \g456073/U$7 ( \63744 , \63739 , \63742 , \63743 );
xor \g130403/U$1 ( \63745 , \63736 , \63744 );
not \g130505/U$3 ( \63746 , \56139 );
not \g130537/U$3 ( \63747 , \56151 );
not \g130537/U$4 ( \63748 , \56141 );
and \g130537/U$2 ( \63749 , \63747 , \63748 );
and \g130537/U$5 ( \63750 , \56151 , \56141 );
nor \g130537/U$1 ( \63751 , \63749 , \63750 );
not \g130505/U$4 ( \63752 , \63751 );
or \g130505/U$2 ( \63753 , \63746 , \63752 );
or \g130505/U$5 ( \63754 , \63751 , \56139 );
nand \g130505/U$1 ( \63755 , \63753 , \63754 );
xor \g130403/U$1_r1 ( \63756 , \63745 , \63755 );
xor \g456070/U$9 ( \63757 , \63650 , \63654 );
xor \g456070/U$9_r1 ( \63758 , \63757 , \63659 );
and \g456070/U$8 ( \63759 , \63664 , \63758 );
xor \g456070/U$11 ( \63760 , \63650 , \63654 );
xor \g456070/U$11_r1 ( \63761 , \63760 , \63659 );
and \g456070/U$10 ( \63762 , \63668 , \63761 );
and \g456070/U$12 ( \63763 , \63664 , \63668 );
or \g456070/U$7 ( \63764 , \63759 , \63762 , \63763 );
xor \g456062/U$1 ( \63765 , \63756 , \63764 );
xor \g130971/U$1 ( \63766 , \56119 , \56121 );
xor \g130971/U$1_r1 ( \63767 , \63766 , \56124 );
xor \g130968/U$4 ( \63768 , \63642 , \63644 );
and \g130968/U$3 ( \63769 , \63768 , \63649 );
and \g130968/U$5 ( \63770 , \63642 , \63644 );
or \g130968/U$2 ( \63771 , \63769 , \63770 );
xor \g456065/U$2 ( \63772 , \63767 , \63771 );
xor \g456069/U$5 ( \63773 , \63676 , \63678 );
and \g456069/U$4 ( \63774 , \63773 , \63683 );
and \g456069/U$6 ( \63775 , \63676 , \63678 );
or \g456069/U$3 ( \63776 , \63774 , \63775 );
xor \g456065/U$1 ( \63777 , \63772 , \63776 );
xor \g456070/U$5 ( \63778 , \63650 , \63654 );
and \g456070/U$4 ( \63779 , \63778 , \63659 );
and \g456070/U$6 ( \63780 , \63650 , \63654 );
or \g456070/U$3 ( \63781 , \63779 , \63780 );
xor \g456069/U$9 ( \63782 , \63676 , \63678 );
xor \g456069/U$9_r1 ( \63783 , \63782 , \63683 );
and \g456069/U$8 ( \63784 , \63692 , \63783 );
xor \g456069/U$11 ( \63785 , \63676 , \63678 );
xor \g456069/U$11_r1 ( \63786 , \63785 , \63683 );
and \g456069/U$10 ( \63787 , \63700 , \63786 );
and \g456069/U$12 ( \63788 , \63692 , \63700 );
or \g456069/U$7 ( \63789 , \63784 , \63787 , \63788 );
xor \g456065/U$1_r1 ( \63790 , \63781 , \63789 );
xor \g456065/U$1_r2 ( \63791 , \63777 , \63790 );
xor \g456062/U$1_r1 ( \63792 , \63765 , \63791 );
xor \g128779/U$1 ( \63793 , \63725 , \63719 );
and \g128776/U$3 ( \63794 , \63792 , \63793 );
nor \g128776/U$1 ( \63795 , \63726 , \63794 );
xor \g456062/U$4 ( \63796 , \63756 , \63764 );
and \g456062/U$3 ( \63797 , \63796 , \63791 );
and \g456062/U$5 ( \63798 , \63756 , \63764 );
nor \g456062/U$2 ( \63799 , \63797 , \63798 );
or \g128772/U$2 ( \63800 , \63795 , \63799 );
xor \g130473/U$1 ( \63801 , \56071 , \56127 );
xor \g130473/U$1_r1 ( \63802 , \63801 , \56130 );
xor \g456065/U$5 ( \63803 , \63767 , \63771 );
and \g456065/U$4 ( \63804 , \63803 , \63776 );
and \g456065/U$6 ( \63805 , \63767 , \63771 );
or \g456065/U$3 ( \63806 , \63804 , \63805 );
xor \g456054/U$2 ( \63807 , \63802 , \63806 );
xor \g130403/U$4 ( \63808 , \63736 , \63744 );
and \g130403/U$3 ( \63809 , \63808 , \63755 );
and \g130403/U$5 ( \63810 , \63736 , \63744 );
or \g130403/U$2 ( \63811 , \63809 , \63810 );
xor \g456054/U$1 ( \63812 , \63807 , \63811 );
xor \g456065/U$9 ( \63813 , \63767 , \63771 );
xor \g456065/U$9_r1 ( \63814 , \63813 , \63776 );
and \g456065/U$8 ( \63815 , \63781 , \63814 );
xor \g456065/U$11 ( \63816 , \63767 , \63771 );
xor \g456065/U$11_r1 ( \63817 , \63816 , \63776 );
and \g456065/U$10 ( \63818 , \63789 , \63817 );
and \g456065/U$12 ( \63819 , \63781 , \63789 );
or \g456065/U$7 ( \63820 , \63815 , \63818 , \63819 );
not \g130354/U$3 ( \63821 , \56291 );
xor \g455953/U$1 ( \63822 , \56153 , \56304 );
not \g130354/U$4 ( \63823 , \63822 );
or \g130354/U$2 ( \63824 , \63821 , \63823 );
or \g130354/U$5 ( \63825 , \63822 , \56291 );
nand \g130354/U$1 ( \63826 , \63824 , \63825 );
xor \g456054/U$1_r1 ( \63827 , \63820 , \63826 );
xor \g456054/U$1_r2 ( \63828 , \63812 , \63827 );
xor \g128775/U$1 ( \63829 , \63799 , \63795 );
and \g128774/U$2 ( \63830 , \63828 , \63829 );
not \g128773/U$1 ( \63831 , \63830 );
nand \g128772/U$1 ( \63832 , \63800 , \63831 );
xor \g456054/U$9 ( \63833 , \63802 , \63806 );
xor \g456054/U$9_r1 ( \63834 , \63833 , \63811 );
and \g456054/U$8 ( \63835 , \63820 , \63834 );
xor \g456054/U$11 ( \63836 , \63802 , \63806 );
xor \g456054/U$11_r1 ( \63837 , \63836 , \63811 );
and \g456054/U$10 ( \63838 , \63826 , \63837 );
and \g456054/U$12 ( \63839 , \63820 , \63826 );
or \g456054/U$7 ( \63840 , \63835 , \63838 , \63839 );
and \g128769/U$2 ( \63841 , \63832 , \63840 );
not \g130286/U$3 ( \63842 , \56061 );
not \g130286/U$4 ( \63843 , \56306 );
or \g130286/U$2 ( \63844 , \63842 , \63843 );
or \g130286/U$5 ( \63845 , \56306 , \56061 );
nand \g130286/U$1 ( \63846 , \63844 , \63845 );
xor \g455952/U$1 ( \63847 , \56133 , \63846 );
xor \g456054/U$5 ( \63848 , \63802 , \63806 );
and \g456054/U$4 ( \63849 , \63848 , \63811 );
and \g456054/U$6 ( \63850 , \63802 , \63806 );
or \g456054/U$3 ( \63851 , \63849 , \63850 );
xor \g130136/U$1 ( \63852 , \63847 , \63851 );
not \g130283/U$3 ( \63853 , \55862 );
not \g130295/U$3 ( \63854 , \55852 );
not \g130295/U$4 ( \63855 , \55869 );
or \g130295/U$2 ( \63856 , \63854 , \63855 );
or \g130295/U$5 ( \63857 , \55869 , \55852 );
nand \g130295/U$1 ( \63858 , \63856 , \63857 );
not \g130283/U$4 ( \63859 , \63858 );
or \g130283/U$2 ( \63860 , \63853 , \63859 );
or \g130283/U$5 ( \63861 , \63858 , \55862 );
nand \g130283/U$1 ( \63862 , \63860 , \63861 );
xor \g130136/U$1_r1 ( \63863 , \63852 , \63862 );
xor \g128771/U$1 ( \63864 , \63840 , \63832 );
and \g128770/U$2 ( \63865 , \63863 , \63864 );
nor \g128769/U$1 ( \63866 , \63841 , \63865 );
not \g130109/U$3 ( \63867 , \56318 );
not \g130109/U$4 ( \63868 , \56308 );
and \g130109/U$2 ( \63869 , \63867 , \63868 );
and \g130109/U$5 ( \63870 , \56318 , \56308 );
nor \g130109/U$1 ( \63871 , \63869 , \63870 );
not \g130087/U$3 ( \63872 , \63871 );
not \g130087/U$4 ( \63873 , \56050 );
and \g130087/U$2 ( \63874 , \63872 , \63873 );
and \g130087/U$5 ( \63875 , \63871 , \56050 );
nor \g130087/U$1 ( \63876 , \63874 , \63875 );
or \g128765/U$2 ( \63877 , \63866 , \63876 );
xor \g130136/U$4 ( \63878 , \63847 , \63851 );
and \g130136/U$3 ( \63879 , \63878 , \63862 );
and \g130136/U$5 ( \63880 , \63847 , \63851 );
or \g130136/U$2 ( \63881 , \63879 , \63880 );
xor \g128768/U$1 ( \63882 , \63876 , \63866 );
and \g128767/U$2 ( \63883 , \63881 , \63882 );
not \g128766/U$1 ( \63884 , \63883 );
nand \g128765/U$1 ( \63885 , \63877 , \63884 );
xor \g128764/U$1 ( \63886 , \56320 , \63885 );
and \g128759/U$2 ( \63887 , \56048 , \63886 );
and \g128759/U$3 ( \63888 , \56320 , \63885 );
not \g128761/U$2 ( \63889 , \63717 );
not \g128785/U$2 ( \63890 , \62296 );
not \g135509/U$2 ( \63891 , \63475 );
nand \g135509/U$1 ( \63892 , \63891 , \63032 , \62799 , \63260 );
nor \g128785/U$1 ( \63893 , \63890 , \63892 , \62557 , \62294 );
nand \g128763/U$1 ( \63894 , \63883 , \63830 , \63893 , \63865 );
nand \g128778/U$1 ( \63895 , \63792 , \63793 );
nand \g128787/U$1 ( \63896 , \63627 , \63628 );
nor \g128761/U$1 ( \63897 , \63889 , \63894 , \63895 , \63896 );
nor \g128759/U$1 ( \63898 , \63887 , \63888 , \63897 );
not \g130081/U$3 ( \63899 , \56043 );
not \g130081/U$4 ( \63900 , \55805 );
and \g130081/U$2 ( \63901 , \63899 , \63900 );
and \g130098/U$2 ( \63902 , \56043 , \55805 );
nor \g130098/U$1 ( \63903 , \63902 , \56041 );
nor \g130081/U$1 ( \63904 , \63901 , \63903 );
or \g128755/U$2 ( \63905 , \63898 , \63904 );
not \g129944/U$3 ( \63906 , \55792 );
xor \g130008/U$1 ( \63907 , \55780 , \55594 );
not \g129944/U$4 ( \63908 , \63907 );
and \g129944/U$2 ( \63909 , \63906 , \63908 );
and \g129944/U$5 ( \63910 , \55792 , \63907 );
nor \g129944/U$1 ( \63911 , \63909 , \63910 );
xnor \g128758/U$1 ( \63912 , \63904 , \63898 );
or \g128755/U$3 ( \63913 , \63911 , \63912 );
nand \g128760/U$1 ( \63914 , \63886 , \63897 , \56048 );
nand \g128755/U$1 ( \63915 , \63905 , \63913 , \63914 );
xor \g128754/U$1 ( \63916 , \55795 , \63915 );
and \g128751/U$2 ( \63917 , \55588 , \63916 );
and \g128751/U$3 ( \63918 , \55795 , \63915 );
nor \g128757/U$1 ( \63919 , \63912 , \63914 , \63911 );
nor \g128751/U$1 ( \63920 , \63917 , \63918 , \63919 );
xnor \g128750/U$1 ( \63921 , \55586 , \63920 );
nand \g128753/U$1 ( \63922 , \63919 , \63916 , \55588 );
or \g129962/U$1 ( \63923 , \55277 , \55211 );
and \g129895/U$2 ( \63924 , \55087 , \63923 );
and \g129895/U$3 ( \63925 , \55211 , \55277 );
nor \g129895/U$1 ( \63926 , \63924 , \63925 );
xor \g129959/U$4 ( \63927 , \54769 , \54989 );
and \g129959/U$3 ( \63928 , \63927 , \55000 );
and \g129959/U$5 ( \63929 , \54769 , \54989 );
or \g129959/U$2 ( \63930 , \63928 , \63929 );
not \g129860/U$3 ( \63931 , \63930 );
xor \g456047/U$9 ( \63932 , \54250 , \54282 );
xor \g456047/U$9_r1 ( \63933 , \63932 , \54291 );
and \g456047/U$8 ( \63934 , \54996 , \63933 );
xor \g456047/U$11 ( \63935 , \54250 , \54282 );
xor \g456047/U$11_r1 ( \63936 , \63935 , \54291 );
and \g456047/U$10 ( \63937 , \54998 , \63936 );
and \g456047/U$12 ( \63938 , \54996 , \54998 );
or \g456047/U$7 ( \63939 , \63934 , \63937 , \63938 );
not \g129966/U$3 ( \63940 , \63939 );
not \g131162/U$3 ( \63941 , \54099 );
xor \g131258/U$1 ( \63942 , \54089 , \54081 );
not \g131162/U$4 ( \63943 , \63942 );
and \g131162/U$2 ( \63944 , \63941 , \63943 );
and \g131162/U$5 ( \63945 , \54099 , \63942 );
nor \g131162/U$1 ( \63946 , \63944 , \63945 );
not \g130321/U$3 ( \63947 , \63946 );
xor \g130357/U$1 ( \63948 , \54133 , \54141 );
xor \g130357/U$1_r1 ( \63949 , \63948 , \54150 );
not \g130321/U$4 ( \63950 , \63949 );
or \g130321/U$2 ( \63951 , \63947 , \63950 );
or \g130321/U$5 ( \63952 , \63949 , \63946 );
nand \g130321/U$1 ( \63953 , \63951 , \63952 );
not \g130292/U$3 ( \63954 , \63953 );
xor \g456067/U$4 ( \63955 , \55231 , \55239 );
and \g456067/U$3 ( \63956 , \63955 , \55248 );
and \g456067/U$5 ( \63957 , \55231 , \55239 );
nor \g456067/U$2 ( \63958 , \63956 , \63957 );
not \g130292/U$4 ( \63959 , \63958 );
and \g130292/U$2 ( \63960 , \63954 , \63959 );
and \g130292/U$5 ( \63961 , \63953 , \63958 );
nor \g130292/U$1 ( \63962 , \63960 , \63961 );
not \g129966/U$4 ( \63963 , \63962 );
and \g129966/U$2 ( \63964 , \63940 , \63963 );
and \g129966/U$5 ( \63965 , \63939 , \63962 );
nor \g129966/U$1 ( \63966 , \63964 , \63965 );
not \g129946/U$3 ( \63967 , \63966 );
or \g130404/U$2 ( \63968 , \55258 , \55222 );
not \g130406/U$3 ( \63969 , \55222 );
not \g130406/U$4 ( \63970 , \55258 );
or \g130406/U$2 ( \63971 , \63969 , \63970 );
nand \g130406/U$1 ( \63972 , \63971 , \55249 );
nand \g130404/U$1 ( \63973 , \63968 , \63972 );
not \g129946/U$4 ( \63974 , \63973 );
and \g129946/U$2 ( \63975 , \63967 , \63974 );
and \g129946/U$5 ( \63976 , \63966 , \63973 );
nor \g129946/U$1 ( \63977 , \63975 , \63976 );
not \g129860/U$4 ( \63978 , \63977 );
or \g129860/U$2 ( \63979 , \63931 , \63978 );
or \g129860/U$5 ( \63980 , \63977 , \63930 );
nand \g129860/U$1 ( \63981 , \63979 , \63980 );
not \g129831/U$3 ( \63982 , \63981 );
not \g130085/U$3 ( \63983 , \55215 );
not \g130085/U$4 ( \63984 , \55262 );
and \g130085/U$2 ( \63985 , \63983 , \63984 );
and \g130102/U$2 ( \63986 , \55215 , \55262 );
not \g130127/U$1 ( \63987 , \55269 );
nor \g130102/U$1 ( \63988 , \63986 , \63987 );
nor \g130085/U$1 ( \63989 , \63985 , \63988 );
not \g129831/U$4 ( \63990 , \63989 );
and \g129831/U$2 ( \63991 , \63982 , \63990 );
and \g129831/U$5 ( \63992 , \63981 , \63989 );
nor \g129831/U$1 ( \63993 , \63991 , \63992 );
xor \g456025/U$1 ( \63994 , \63926 , \63993 );
xor \g130050/U$1 ( \63995 , \54339 , \54368 );
xor \g130050/U$1_r1 ( \63996 , \63995 , \54377 );
not \g130011/U$3 ( \63997 , \63996 );
xor \g131034/U$4 ( \63998 , \55005 , \55011 );
and \g131034/U$3 ( \63999 , \63998 , \55016 );
and \g131034/U$5 ( \64000 , \55005 , \55011 );
or \g131034/U$2 ( \64001 , \63999 , \64000 );
not \g130011/U$4 ( \64002 , \64001 );
and \g130011/U$2 ( \64003 , \63997 , \64002 );
and \g130011/U$5 ( \64004 , \63996 , \64001 );
nor \g130011/U$1 ( \64005 , \64003 , \64004 );
not \g129961/U$3 ( \64006 , \64005 );
xor \g130219/U$1 ( \64007 , \54389 , \54397 );
xor \g130219/U$1_r1 ( \64008 , \64007 , \54406 );
not \g129961/U$4 ( \64009 , \64008 );
and \g129961/U$2 ( \64010 , \64006 , \64009 );
and \g129961/U$5 ( \64011 , \64005 , \64008 );
nor \g129961/U$1 ( \64012 , \64010 , \64011 );
not \g130084/U$3 ( \64013 , \55022 );
not \g130084/U$4 ( \64014 , \55017 );
and \g130084/U$2 ( \64015 , \64013 , \64014 );
and \g130101/U$2 ( \64016 , \55022 , \55017 );
not \g130126/U$1 ( \64017 , \55079 );
nor \g130101/U$1 ( \64018 , \64016 , \64017 );
nor \g130084/U$1 ( \64019 , \64015 , \64018 );
xor \g129806/U$1 ( \64020 , \64012 , \64019 );
xor \g130036/U$1 ( \64021 , \54294 , \54296 );
xor \g130036/U$1_r1 ( \64022 , \64021 , \54325 );
not \g129965/U$3 ( \64023 , \64022 );
xor \g456052/U$4 ( \64024 , \55025 , \55053 );
and \g456052/U$3 ( \64025 , \64024 , \55078 );
and \g456052/U$5 ( \64026 , \55025 , \55053 );
nor \g456052/U$2 ( \64027 , \64025 , \64026 );
not \g129965/U$4 ( \64028 , \64027 );
and \g129965/U$2 ( \64029 , \64023 , \64028 );
and \g129965/U$5 ( \64030 , \64022 , \64027 );
nor \g129965/U$1 ( \64031 , \64029 , \64030 );
not \g129945/U$3 ( \64032 , \64031 );
xor \g130970/U$1 ( \64033 , \54207 , \54209 );
xor \g130970/U$1_r1 ( \64034 , \64033 , \54239 );
not \g129945/U$4 ( \64035 , \64034 );
and \g129945/U$2 ( \64036 , \64032 , \64035 );
and \g129945/U$5 ( \64037 , \64031 , \64034 );
nor \g129945/U$1 ( \64038 , \64036 , \64037 );
xor \g129806/U$1_r1 ( \64039 , \64020 , \64038 );
xor \g456025/U$1_r1 ( \64040 , \63994 , \64039 );
nor \g128749/U$1 ( \64041 , \63921 , \63922 , \64040 );
xor \g456025/U$4 ( \64042 , \63926 , \63993 );
and \g456025/U$3 ( \64043 , \64042 , \64039 );
and \g456025/U$5 ( \64044 , \63926 , \63993 );
nor \g456025/U$2 ( \64045 , \64043 , \64044 );
or \g128747/U$2 ( \64046 , \63921 , \64040 );
or \g128747/U$3 ( \64047 , \55586 , \63920 );
nand \g128747/U$1 ( \64048 , \64046 , \64047 , \63922 );
xor \g128746/U$1 ( \64049 , \64045 , \64048 );
xor \g456028/U$2 ( \64050 , \54166 , \54168 );
xor \g456028/U$1 ( \64051 , \64050 , \54171 );
not \g130969/U$1 ( \64052 , \64034 );
or \g129990/U$2 ( \64053 , \64027 , \64052 );
not \g130006/U$3 ( \64054 , \64052 );
not \g130006/U$4 ( \64055 , \64027 );
or \g130006/U$2 ( \64056 , \64054 , \64055 );
nand \g130006/U$1 ( \64057 , \64056 , \64022 );
nand \g129990/U$1 ( \64058 , \64053 , \64057 );
xor \g456043/U$1 ( \64059 , \54242 , \54328 );
xor \g456043/U$1_r1 ( \64060 , \64059 , \54410 );
xor \g456028/U$1_r1 ( \64061 , \64058 , \64060 );
xor \g456028/U$1_r2 ( \64062 , \64051 , \64061 );
not \g130347/U$1 ( \64063 , \63973 );
or \g129991/U$2 ( \64064 , \63962 , \64063 );
not \g130007/U$3 ( \64065 , \64063 );
not \g130007/U$4 ( \64066 , \63962 );
or \g130007/U$2 ( \64067 , \64065 , \64066 );
nand \g130007/U$1 ( \64068 , \64067 , \63939 );
nand \g129991/U$1 ( \64069 , \64064 , \64068 );
xor \g456034/U$2 ( \64070 , \54153 , \54155 );
xor \g456034/U$1 ( \64071 , \64070 , \54158 );
or \g130323/U$2 ( \64072 , \63958 , \63946 );
not \g130329/U$3 ( \64073 , \63946 );
not \g130329/U$4 ( \64074 , \63958 );
or \g130329/U$2 ( \64075 , \64073 , \64074 );
nand \g130329/U$1 ( \64076 , \64075 , \63949 );
nand \g130323/U$1 ( \64077 , \64072 , \64076 );
not \g130217/U$1 ( \64078 , \64008 );
or \g130014/U$2 ( \64079 , \64078 , \64001 );
not \g130018/U$3 ( \64080 , \64001 );
not \g130018/U$4 ( \64081 , \64078 );
or \g130018/U$2 ( \64082 , \64080 , \64081 );
nand \g130018/U$1 ( \64083 , \64082 , \63996 );
nand \g130014/U$1 ( \64084 , \64079 , \64083 );
xor \g456034/U$1_r1 ( \64085 , \64077 , \64084 );
xor \g456034/U$1_r2 ( \64086 , \64071 , \64085 );
not \g129761/U$3 ( \64087 , \64086 );
xor \g129806/U$4 ( \64088 , \64012 , \64019 );
and \g129806/U$3 ( \64089 , \64088 , \64038 );
and \g129806/U$5 ( \64090 , \64012 , \64019 );
or \g129806/U$2 ( \64091 , \64089 , \64090 );
not \g129761/U$4 ( \64092 , \64091 );
or \g129761/U$2 ( \64093 , \64087 , \64092 );
or \g129761/U$5 ( \64094 , \64091 , \64086 );
nand \g129761/U$1 ( \64095 , \64093 , \64094 );
xor \g455947/U$1 ( \64096 , \64069 , \64095 );
xor \g456016/U$1 ( \64097 , \64062 , \64096 );
or \g129856/U$2 ( \64098 , \63977 , \63989 );
not \g129858/U$3 ( \64099 , \63989 );
not \g129858/U$4 ( \64100 , \63977 );
or \g129858/U$2 ( \64101 , \64099 , \64100 );
nand \g129858/U$1 ( \64102 , \64101 , \63930 );
nand \g129856/U$1 ( \64103 , \64098 , \64102 );
xor \g456016/U$1_r1 ( \64104 , \64097 , \64103 );
nand \g128745/U$1 ( \64105 , \64041 , \64049 , \64104 );
not \g128737/U$3 ( \64106 , \64105 );
and \g128743/U$2 ( \64107 , \64045 , \64048 );
and \g128743/U$3 ( \64108 , \64104 , \64049 );
nor \g128743/U$1 ( \64109 , \64107 , \64108 , \64041 );
xor \g456016/U$4 ( \64110 , \64062 , \64096 );
and \g456016/U$3 ( \64111 , \64110 , \64103 );
and \g456016/U$5 ( \64112 , \64062 , \64096 );
nor \g456016/U$2 ( \64113 , \64111 , \64112 );
or \g128739/U$2 ( \64114 , \64109 , \64113 );
and \g129765/U$2 ( \64115 , \64086 , \64069 );
not \g129767/U$3 ( \64116 , \64086 );
not \g129767/U$4 ( \64117 , \64069 );
and \g129767/U$2 ( \64118 , \64116 , \64117 );
nor \g129767/U$1 ( \64119 , \64118 , \64091 );
nor \g129765/U$1 ( \64120 , \64115 , \64119 );
not \g129594/U$3 ( \64121 , \64120 );
xor \g456029/U$2 ( \64122 , \54049 , \54105 );
xor \g456029/U$1 ( \64123 , \64122 , \54108 );
xor \g456029/U$1_r1 ( \64124 , \54161 , \54174 );
xor \g456029/U$1_r2 ( \64125 , \64123 , \64124 );
xor \g456028/U$9 ( \64126 , \54166 , \54168 );
xor \g456028/U$9_r1 ( \64127 , \64126 , \54171 );
and \g456028/U$8 ( \64128 , \64058 , \64127 );
xor \g456028/U$11 ( \64129 , \54166 , \54168 );
xor \g456028/U$11_r1 ( \64130 , \64129 , \54171 );
and \g456028/U$10 ( \64131 , \64060 , \64130 );
and \g456028/U$12 ( \64132 , \64058 , \64060 );
or \g456028/U$7 ( \64133 , \64128 , \64131 , \64132 );
xor \g456023/U$1 ( \64134 , \64125 , \64133 );
xor \g456034/U$9 ( \64135 , \54153 , \54155 );
xor \g456034/U$9_r1 ( \64136 , \64135 , \54158 );
and \g456034/U$8 ( \64137 , \64077 , \64136 );
xor \g456034/U$11 ( \64138 , \54153 , \54155 );
xor \g456034/U$11_r1 ( \64139 , \64138 , \54158 );
and \g456034/U$10 ( \64140 , \64084 , \64139 );
and \g456034/U$12 ( \64141 , \64077 , \64084 );
or \g456034/U$7 ( \64142 , \64137 , \64140 , \64141 );
xor \g456023/U$1_r1 ( \64143 , \64134 , \64142 );
not \g129594/U$4 ( \64144 , \64143 );
or \g129594/U$2 ( \64145 , \64121 , \64144 );
or \g129594/U$5 ( \64146 , \64143 , \64120 );
nand \g129594/U$1 ( \64147 , \64145 , \64146 );
not \g129561/U$3 ( \64148 , \64147 );
xor \g456021/U$2 ( \64149 , \54417 , \54423 );
xor \g456021/U$1 ( \64150 , \64149 , \54430 );
xor \g456021/U$1_r1 ( \64151 , \54413 , \54438 );
xor \g456021/U$1_r2 ( \64152 , \64150 , \64151 );
not \g129561/U$4 ( \64153 , \64152 );
and \g129561/U$2 ( \64154 , \64148 , \64153 );
and \g129561/U$5 ( \64155 , \64147 , \64152 );
nor \g129561/U$1 ( \64156 , \64154 , \64155 );
not \g128741/U$2 ( \64157 , \64156 );
xor \g128742/U$1 ( \64158 , \64113 , \64109 );
nand \g128741/U$1 ( \64159 , \64157 , \64158 );
nand \g128739/U$1 ( \64160 , \64114 , \64159 );
not \g128737/U$4 ( \64161 , \64160 );
or \g128737/U$2 ( \64162 , \64106 , \64161 );
or \g128737/U$5 ( \64163 , \64160 , \64105 );
nand \g128737/U$1 ( \64164 , \64162 , \64163 );
or \g129588/U$2 ( \64165 , \64152 , \64120 );
not \g129591/U$3 ( \64166 , \64120 );
not \g129591/U$4 ( \64167 , \64152 );
or \g129591/U$2 ( \64168 , \64166 , \64167 );
nand \g129591/U$1 ( \64169 , \64168 , \64143 );
nand \g129588/U$1 ( \64170 , \64165 , \64169 );
and \g128733/U$2 ( \64171 , \64164 , \64170 );
not \g129660/U$3 ( \64172 , \54469 );
not \g129660/U$4 ( \64173 , \54475 );
or \g129660/U$2 ( \64174 , \64172 , \64173 );
or \g129660/U$5 ( \64175 , \54475 , \54469 );
nand \g129660/U$1 ( \64176 , \64174 , \64175 );
not \g129606/U$3 ( \64177 , \64176 );
not \g129606/U$4 ( \64178 , \54465 );
and \g129606/U$2 ( \64179 , \64177 , \64178 );
and \g129606/U$5 ( \64180 , \64176 , \54465 );
nor \g129606/U$1 ( \64181 , \64179 , \64180 );
not \g129446/U$3 ( \64182 , \64181 );
xor \g456023/U$4 ( \64183 , \64125 , \64133 );
and \g456023/U$3 ( \64184 , \64183 , \64142 );
and \g456023/U$5 ( \64185 , \64125 , \64133 );
nor \g456023/U$2 ( \64186 , \64184 , \64185 );
not \g129476/U$3 ( \64187 , \64186 );
not \g129593/U$3 ( \64188 , \54125 );
not \g129593/U$4 ( \64189 , \54443 );
or \g129593/U$2 ( \64190 , \64188 , \64189 );
or \g129593/U$5 ( \64191 , \54443 , \54125 );
nand \g129593/U$1 ( \64192 , \64190 , \64191 );
xor \g455945/U$1 ( \64193 , \54179 , \64192 );
not \g129476/U$4 ( \64194 , \64193 );
or \g129476/U$2 ( \64195 , \64187 , \64194 );
or \g129476/U$5 ( \64196 , \64193 , \64186 );
nand \g129476/U$1 ( \64197 , \64195 , \64196 );
not \g129446/U$4 ( \64198 , \64197 );
or \g129446/U$2 ( \64199 , \64182 , \64198 );
or \g129446/U$5 ( \64200 , \64197 , \64181 );
nand \g129446/U$1 ( \64201 , \64199 , \64200 );
xor \g128736/U$1 ( \64202 , \64170 , \64164 );
and \g128735/U$2 ( \64203 , \64201 , \64202 );
nor \g128738/U$1 ( \64204 , \64159 , \64105 );
nor \g128733/U$1 ( \64205 , \64171 , \64203 , \64204 );
not \g129488/U$3 ( \64206 , \64181 );
not \g129488/U$4 ( \64207 , \64186 );
and \g129488/U$2 ( \64208 , \64206 , \64207 );
and \g129491/U$2 ( \64209 , \64181 , \64186 );
not \g129526/U$1 ( \64210 , \64193 );
nor \g129491/U$1 ( \64211 , \64209 , \64210 );
nor \g129488/U$1 ( \64212 , \64208 , \64211 );
or \g128729/U$2 ( \64213 , \64205 , \64212 );
not \g129386/U$3 ( \64214 , \54479 );
not \g129386/U$4 ( \64215 , \54445 );
and \g129386/U$2 ( \64216 , \64214 , \64215 );
and \g129386/U$5 ( \64217 , \54479 , \54445 );
nor \g129386/U$1 ( \64218 , \64216 , \64217 );
not \g129356/U$3 ( \64219 , \64218 );
not \g129356/U$4 ( \64220 , \53996 );
and \g129356/U$2 ( \64221 , \64219 , \64220 );
and \g129356/U$5 ( \64222 , \64218 , \53996 );
nor \g129356/U$1 ( \64223 , \64221 , \64222 );
xnor \g128732/U$1 ( \64224 , \64212 , \64205 );
or \g128729/U$3 ( \64225 , \64223 , \64224 );
nand \g128734/U$1 ( \64226 , \64204 , \64203 );
nand \g128729/U$1 ( \64227 , \64213 , \64225 , \64226 );
and \g128725/U$2 ( \64228 , \54481 , \64227 );
not \g129459/U$3 ( \64229 , \53443 );
xor \g129492/U$1 ( \64230 , \53424 , \53577 );
not \g129459/U$4 ( \64231 , \64230 );
or \g129459/U$2 ( \64232 , \64229 , \64231 );
or \g129459/U$5 ( \64233 , \64230 , \53443 );
nand \g129459/U$1 ( \64234 , \64232 , \64233 );
xor \g456003/U$9 ( \64235 , \53961 , \53963 );
xor \g456003/U$9_r1 ( \64236 , \64235 , \53976 );
and \g456003/U$8 ( \64237 , \54459 , \64236 );
xor \g456003/U$11 ( \64238 , \53961 , \53963 );
xor \g456003/U$11_r1 ( \64239 , \64238 , \53976 );
and \g456003/U$10 ( \64240 , \54477 , \64239 );
and \g456003/U$12 ( \64241 , \54459 , \54477 );
or \g456003/U$7 ( \64242 , \64237 , \64240 , \64241 );
not \g129221/U$3 ( \64243 , \64242 );
xor \g129279/U$1 ( \64244 , \53836 , \53980 );
xor \g129279/U$1_r1 ( \64245 , \64244 , \53983 );
not \g129221/U$4 ( \64246 , \64245 );
or \g129221/U$2 ( \64247 , \64243 , \64246 );
or \g129221/U$5 ( \64248 , \64245 , \64242 );
nand \g129221/U$1 ( \64249 , \64247 , \64248 );
xor \g455937/U$1 ( \64250 , \64234 , \64249 );
xor \g128728/U$1 ( \64251 , \54481 , \64227 );
and \g128725/U$3 ( \64252 , \64250 , \64251 );
nor \g128731/U$1 ( \64253 , \64224 , \64226 , \64223 );
nor \g128725/U$1 ( \64254 , \64228 , \64252 , \64253 );
and \g129230/U$2 ( \64255 , \64234 , \64242 );
not \g129242/U$3 ( \64256 , \64234 );
not \g129242/U$4 ( \64257 , \64242 );
and \g129242/U$2 ( \64258 , \64256 , \64257 );
nor \g129242/U$1 ( \64259 , \64258 , \64245 );
nor \g129230/U$1 ( \64260 , \64255 , \64259 );
or \g128721/U$2 ( \64261 , \64254 , \64260 );
xor \g455989/U$1 ( \64262 , \53744 , \53986 );
xor \g455989/U$1_r1 ( \64263 , \64262 , \53991 );
xnor \g128724/U$1 ( \64264 , \64260 , \64254 );
or \g128721/U$3 ( \64265 , \64263 , \64264 );
nand \g128727/U$1 ( \64266 , \64253 , \64251 , \64250 );
nand \g128721/U$1 ( \64267 , \64261 , \64265 , \64266 );
xor \g128720/U$1 ( \64268 , \53994 , \64267 );
and \g128717/U$2 ( \64269 , \53734 , \64268 );
and \g128717/U$3 ( \64270 , \53994 , \64267 );
nor \g128723/U$1 ( \64271 , \64264 , \64266 , \64263 );
nor \g128717/U$1 ( \64272 , \64269 , \64270 , \64271 );
xnor \g128716/U$1 ( \64273 , \53724 , \64272 );
nand \g128719/U$1 ( \64274 , \64271 , \64268 , \53734 );
xor \g129055/U$4 ( \64275 , \53681 , \53685 );
and \g129055/U$3 ( \64276 , \64275 , \53721 );
and \g129055/U$5 ( \64277 , \53681 , \53685 );
or \g129055/U$2 ( \64278 , \64276 , \64277 );
not \g128923/U$3 ( \64279 , \64278 );
or \g129266/U$2 ( \64280 , \53717 , \53688 );
not \g129269/U$3 ( \64281 , \53688 );
not \g129269/U$4 ( \64282 , \53717 );
or \g129269/U$2 ( \64283 , \64281 , \64282 );
nand \g129269/U$1 ( \64284 , \64283 , \53704 );
nand \g129266/U$1 ( \64285 , \64280 , \64284 );
not \g129357/U$3 ( \64286 , \52555 );
xnor \g129433/U$1 ( \64287 , \52595 , \52593 );
not \g129357/U$4 ( \64288 , \64287 );
or \g129357/U$2 ( \64289 , \64286 , \64288 );
or \g129357/U$5 ( \64290 , \64287 , \52555 );
nand \g129357/U$1 ( \64291 , \64289 , \64290 );
or \g129440/U$2 ( \64292 , \52877 , \52837 );
and \g129452/U$2 ( \64293 , \52877 , \52837 );
nor \g129452/U$1 ( \64294 , \64293 , \52834 );
not \g129451/U$1 ( \64295 , \64294 );
nand \g129440/U$1 ( \64296 , \64292 , \64295 );
xor \g129194/U$1 ( \64297 , \64291 , \64296 );
xor \g129288/U$4 ( \64298 , \53694 , \53700 );
and \g129288/U$3 ( \64299 , \64298 , \53703 );
and \g129288/U$5 ( \64300 , \53694 , \53700 );
or \g129288/U$2 ( \64301 , \64299 , \64300 );
xor \g129194/U$1_r1 ( \64302 , \64297 , \64301 );
xor \g128958/U$1 ( \64303 , \64285 , \64302 );
not \g129033/U$3 ( \64304 , \52778 );
xor \g455933/U$1 ( \64305 , \52801 , \52806 );
not \g129033/U$4 ( \64306 , \64305 );
or \g129033/U$2 ( \64307 , \64304 , \64306 );
or \g129033/U$5 ( \64308 , \64305 , \52778 );
nand \g129033/U$1 ( \64309 , \64307 , \64308 );
xor \g128958/U$1_r1 ( \64310 , \64303 , \64309 );
not \g128923/U$4 ( \64311 , \64310 );
or \g128923/U$2 ( \64312 , \64279 , \64311 );
or \g128923/U$5 ( \64313 , \64310 , \64278 );
nand \g128923/U$1 ( \64314 , \64312 , \64313 );
not \g128910/U$3 ( \64315 , \64314 );
xor \g129262/U$4 ( \64316 , \52882 , \53049 );
and \g129262/U$3 ( \64317 , \64316 , \53210 );
and \g129262/U$5 ( \64318 , \52882 , \53049 );
or \g129262/U$2 ( \64319 , \64317 , \64318 );
not \g128910/U$4 ( \64320 , \64319 );
and \g128910/U$2 ( \64321 , \64315 , \64320 );
and \g128910/U$5 ( \64322 , \64314 , \64319 );
nor \g128910/U$1 ( \64323 , \64321 , \64322 );
nor \g128715/U$1 ( \64324 , \64273 , \64274 , \64323 );
not \g128708/U$3 ( \64325 , \64324 );
or \g128713/U$2 ( \64326 , \64272 , \53724 );
or \g128713/U$3 ( \64327 , \64323 , \64273 );
nand \g128713/U$1 ( \64328 , \64326 , \64327 , \64274 );
or \g128932/U$2 ( \64329 , \64278 , \64319 );
not \g128933/U$3 ( \64330 , \64319 );
not \g128933/U$4 ( \64331 , \64278 );
or \g128933/U$2 ( \64332 , \64330 , \64331 );
nand \g128933/U$1 ( \64333 , \64332 , \64310 );
nand \g128932/U$1 ( \64334 , \64329 , \64333 );
and \g128710/U$2 ( \64335 , \64328 , \64334 );
xor \g128958/U$4 ( \64336 , \64285 , \64302 );
and \g128958/U$3 ( \64337 , \64336 , \64309 );
and \g128958/U$5 ( \64338 , \64285 , \64302 );
or \g128958/U$2 ( \64339 , \64337 , \64338 );
xor \g129194/U$4 ( \64340 , \64291 , \64296 );
and \g129194/U$3 ( \64341 , \64340 , \64301 );
and \g129194/U$5 ( \64342 , \64291 , \64296 );
or \g129194/U$2 ( \64343 , \64341 , \64342 );
xor \g128869/U$1 ( \64344 , \64339 , \64343 );
not \g128938/U$3 ( \64345 , \52813 );
xor \g128973/U$1 ( \64346 , \52808 , \52820 );
not \g128938/U$4 ( \64347 , \64346 );
or \g128938/U$2 ( \64348 , \64345 , \64347 );
or \g128938/U$5 ( \64349 , \64346 , \52813 );
nand \g128938/U$1 ( \64350 , \64348 , \64349 );
xor \g128869/U$1_r1 ( \64351 , \64344 , \64350 );
xor \g128712/U$1 ( \64352 , \64334 , \64328 );
and \g128711/U$2 ( \64353 , \64351 , \64352 );
nor \g128710/U$1 ( \64354 , \64335 , \64353 );
not \g128708/U$4 ( \64355 , \64354 );
or \g128708/U$2 ( \64356 , \64325 , \64355 );
or \g128708/U$5 ( \64357 , \64354 , \64324 );
nand \g128708/U$1 ( \64358 , \64356 , \64357 );
xor \g128869/U$4 ( \64359 , \64339 , \64343 );
and \g128869/U$3 ( \64360 , \64359 , \64350 );
and \g128869/U$5 ( \64361 , \64339 , \64343 );
or \g128869/U$2 ( \64362 , \64360 , \64361 );
and \g128704/U$2 ( \64363 , \64358 , \64362 );
not \g128862/U$3 ( \64364 , \52771 );
xor \g128880/U$1 ( \64365 , \52822 , \52760 );
not \g128862/U$4 ( \64366 , \64365 );
or \g128862/U$2 ( \64367 , \64364 , \64366 );
or \g128862/U$5 ( \64368 , \64365 , \52771 );
nand \g128862/U$1 ( \64369 , \64367 , \64368 );
xor \g128707/U$1 ( \64370 , \64362 , \64358 );
and \g128706/U$2 ( \64371 , \64369 , \64370 );
and \g128709/U$1 ( \64372 , \64353 , \64324 );
nor \g128704/U$1 ( \64373 , \64363 , \64371 , \64372 );
xnor \g128703/U$1 ( \64374 , \52824 , \64373 );
nand \g128705/U$1 ( \64375 , \64372 , \64371 );
xor \g128918/U$4 ( \64376 , \52549 , \52752 );
and \g128918/U$3 ( \64377 , \64376 , \52759 );
and \g128918/U$5 ( \64378 , \52549 , \52752 );
or \g128918/U$2 ( \64379 , \64377 , \64378 );
xnor \g128999/U$1 ( \64380 , \52400 , \52464 );
not \g128950/U$3 ( \64381 , \64380 );
not \g128950/U$4 ( \64382 , \52016 );
and \g128950/U$2 ( \64383 , \64381 , \64382 );
and \g128950/U$5 ( \64384 , \64380 , \52016 );
nor \g128950/U$1 ( \64385 , \64383 , \64384 );
xnor \g128881/U$1 ( \64386 , \64379 , \64385 );
not \g128852/U$3 ( \64387 , \64386 );
xor \g128928/U$1 ( \64388 , \52502 , \52506 );
xor \g128928/U$1_r1 ( \64389 , \64388 , \52509 );
not \g128852/U$4 ( \64390 , \64389 );
and \g128852/U$2 ( \64391 , \64387 , \64390 );
and \g128852/U$5 ( \64392 , \64386 , \64389 );
nor \g128852/U$1 ( \64393 , \64391 , \64392 );
nor \g128702/U$1 ( \64394 , \64374 , \64375 , \64393 );
not \g455925/U$2 ( \64395 , \64394 );
or \g128850/U$2 ( \64396 , \64385 , \64379 );
not \g128853/U$3 ( \64397 , \64379 );
not \g128853/U$4 ( \64398 , \64385 );
or \g128853/U$2 ( \64399 , \64397 , \64398 );
nand \g128853/U$1 ( \64400 , \64399 , \64389 );
nand \g128850/U$1 ( \64401 , \64396 , \64400 );
or \g128699/U$2 ( \64402 , \64374 , \64393 );
or \g128699/U$3 ( \64403 , \52824 , \64373 );
nand \g128699/U$1 ( \64404 , \64402 , \64403 , \64375 );
xor \g128698/U$1 ( \64405 , \64401 , \64404 );
xor \g455969/U$2 ( \64406 , \52480 , \52482 );
xor \g455969/U$1 ( \64407 , \64406 , \52485 );
xor \g455969/U$1_r1 ( \64408 , \52466 , \52514 );
xor \g455969/U$1_r2 ( \64409 , \64407 , \64408 );
and \g128695/U$2 ( \64410 , \64405 , \64409 );
and \g128695/U$3 ( \64411 , \64401 , \64404 );
nor \g128695/U$1 ( \64412 , \64410 , \64411 );
nand \g455925/U$1 ( \64413 , \64395 , \64412 );
and \g128690/U$2 ( \64414 , \52519 , \64413 );
xor \g455969/U$5 ( \64415 , \52480 , \52482 );
and \g455969/U$4 ( \64416 , \64415 , \52485 );
and \g455969/U$6 ( \64417 , \52480 , \52482 );
or \g455969/U$3 ( \64418 , \64416 , \64417 );
xor \g455971/U$9 ( \64419 , \51908 , \51918 );
xor \g455971/U$9_r1 ( \64420 , \64419 , \51929 );
and \g455971/U$8 ( \64421 , \52497 , \64420 );
xor \g455971/U$11 ( \64422 , \51908 , \51918 );
xor \g455971/U$11_r1 ( \64423 , \64422 , \51929 );
and \g455971/U$10 ( \64424 , \52512 , \64423 );
and \g455971/U$12 ( \64425 , \52497 , \52512 );
or \g455971/U$7 ( \64426 , \64421 , \64424 , \64425 );
xor \g455968/U$1 ( \64427 , \64418 , \64426 );
xor \g128858/U$1 ( \64428 , \51794 , \51932 );
xor \g128858/U$1_r1 ( \64429 , \64428 , \51939 );
xor \g455968/U$1_r1 ( \64430 , \64427 , \64429 );
xor \g128693/U$1 ( \64431 , \52519 , \64413 );
and \g128690/U$3 ( \64432 , \64430 , \64431 );
and \g128697/U$1 ( \64433 , \64405 , \64394 , \64409 );
nor \g128690/U$1 ( \64434 , \64414 , \64432 , \64433 );
xor \g455968/U$4 ( \64435 , \64418 , \64426 );
and \g455968/U$3 ( \64436 , \64435 , \64429 );
and \g455968/U$5 ( \64437 , \64418 , \64426 );
nor \g455968/U$2 ( \64438 , \64436 , \64437 );
or \g128686/U$2 ( \64439 , \64434 , \64438 );
not \g128842/U$3 ( \64440 , \51942 );
not \g128842/U$4 ( \64441 , \51773 );
and \g128842/U$2 ( \64442 , \64440 , \64441 );
and \g128842/U$5 ( \64443 , \51942 , \51773 );
nor \g128842/U$1 ( \64444 , \64442 , \64443 );
not \g128826/U$3 ( \64445 , \64444 );
not \g128826/U$4 ( \64446 , \51779 );
and \g128826/U$2 ( \64447 , \64445 , \64446 );
and \g128826/U$5 ( \64448 , \64444 , \51779 );
nor \g128826/U$1 ( \64449 , \64447 , \64448 );
xnor \g128689/U$1 ( \64450 , \64438 , \64434 );
or \g128686/U$3 ( \64451 , \64449 , \64450 );
nand \g128692/U$1 ( \64452 , \64433 , \64431 , \64430 );
nand \g128686/U$1 ( \64453 , \64439 , \64451 , \64452 );
xor \g128685/U$1 ( \64454 , \51944 , \64453 );
and \g128682/U$2 ( \64455 , \51769 , \64454 );
and \g128682/U$3 ( \64456 , \51944 , \64453 );
nor \g128688/U$1 ( \64457 , \64450 , \64452 , \64449 );
nor \g128682/U$1 ( \64458 , \64455 , \64456 , \64457 );
not \g128838/U$3 ( \64459 , \51279 );
not \g128838/U$4 ( \64460 , \51448 );
or \g128838/U$2 ( \64461 , \64459 , \64460 );
or \g128838/U$5 ( \64462 , \51448 , \51279 );
nand \g128838/U$1 ( \64463 , \64461 , \64462 );
not \g128825/U$3 ( \64464 , \64463 );
not \g128825/U$4 ( \64465 , \51277 );
and \g128825/U$2 ( \64466 , \64464 , \64465 );
and \g128825/U$5 ( \64467 , \64463 , \51277 );
nor \g128825/U$1 ( \64468 , \64466 , \64467 );
or \g128678/U$2 ( \64469 , \64458 , \64468 );
not \g128829/U$3 ( \64470 , \51764 );
not \g128829/U$4 ( \64471 , \51452 );
and \g128829/U$2 ( \64472 , \64470 , \64471 );
and \g128835/U$2 ( \64473 , \51764 , \51452 );
nor \g128835/U$1 ( \64474 , \64473 , \51762 );
nor \g128829/U$1 ( \64475 , \64472 , \64474 );
xnor \g128681/U$1 ( \64476 , \64468 , \64458 );
or \g128678/U$3 ( \64477 , \64475 , \64476 );
nand \g128684/U$1 ( \64478 , \64457 , \64454 , \51769 );
nand \g128678/U$1 ( \64479 , \64469 , \64477 , \64478 );
and \g128674/U$2 ( \64480 , \51450 , \64479 );
not \g128824/U$3 ( \64481 , \51266 );
xor \g128837/U$1 ( \64482 , \51263 , \51271 );
not \g128824/U$4 ( \64483 , \64482 );
or \g128824/U$2 ( \64484 , \64481 , \64483 );
or \g128824/U$5 ( \64485 , \64482 , \51266 );
nand \g128824/U$1 ( \64486 , \64484 , \64485 );
xor \g128677/U$1 ( \64487 , \51450 , \64479 );
and \g128674/U$3 ( \64488 , \64486 , \64487 );
nor \g128679/U$1 ( \64489 , \64476 , \64478 , \64475 );
nor \g128674/U$1 ( \64490 , \64480 , \64488 , \64489 );
xnor \g128673/U$1 ( \64491 , \51273 , \64490 );
not \g128841/U$3 ( \64492 , \51027 );
not \g128841/U$4 ( \64493 , \50817 );
and \g128841/U$2 ( \64494 , \64492 , \64493 );
and \g128841/U$5 ( \64495 , \51027 , \50817 );
nor \g128841/U$1 ( \64496 , \64494 , \64495 );
not \g128832/U$3 ( \64497 , \64496 );
not \g128832/U$4 ( \64498 , \50810 );
and \g128832/U$2 ( \64499 , \64497 , \64498 );
and \g128832/U$5 ( \64500 , \64496 , \50810 );
nor \g128832/U$1 ( \64501 , \64499 , \64500 );
or \g128670/U$2 ( \64502 , \64491 , \64501 );
or \g128670/U$3 ( \64503 , \51273 , \64490 );
nand \g128676/U$1 ( \64504 , \64489 , \64487 , \64486 );
nand \g128670/U$1 ( \64505 , \64502 , \64503 , \64504 );
xor \g128669/U$1 ( \64506 , \51030 , \64505 );
and \g128666/U$2 ( \64507 , \50806 , \64506 );
and \g128666/U$3 ( \64508 , \51030 , \64505 );
nor \g128672/U$1 ( \64509 , \64491 , \64504 , \64501 );
nor \g128666/U$1 ( \64510 , \64507 , \64508 , \64509 );
xnor \g128665/U$1 ( \64511 , \50800 , \64510 );
not \g128902/U$3 ( \64512 , \50408 );
not \g128902/U$4 ( \64513 , \50422 );
or \g128902/U$2 ( \64514 , \64512 , \64513 );
or \g128902/U$5 ( \64515 , \50422 , \50408 );
nand \g128902/U$1 ( \64516 , \64514 , \64515 );
not \g128875/U$3 ( \64517 , \64516 );
not \g128875/U$4 ( \64518 , \50412 );
and \g128875/U$2 ( \64519 , \64517 , \64518 );
and \g128875/U$5 ( \64520 , \64516 , \50412 );
nor \g128875/U$1 ( \64521 , \64519 , \64520 );
or \g128662/U$2 ( \64522 , \64511 , \64521 );
or \g128662/U$3 ( \64523 , \50800 , \64510 );
nand \g128668/U$1 ( \64524 , \64509 , \64506 , \50806 );
nand \g128662/U$1 ( \64525 , \64522 , \64523 , \64524 );
and \g128658/U$2 ( \64526 , \50424 , \64525 );
not \g128876/U$3 ( \64527 , \50059 );
xor \g128903/U$1 ( \64528 , \50185 , \49990 );
not \g128876/U$4 ( \64529 , \64528 );
or \g128876/U$2 ( \64530 , \64527 , \64529 );
or \g128876/U$5 ( \64531 , \64528 , \50059 );
nand \g128876/U$1 ( \64532 , \64530 , \64531 );
xor \g128661/U$1 ( \64533 , \50424 , \64525 );
and \g128658/U$3 ( \64534 , \64532 , \64533 );
nor \g128664/U$1 ( \64535 , \64511 , \64524 , \64521 );
nor \g128658/U$1 ( \64536 , \64526 , \64534 , \64535 );
xnor \g128657/U$1 ( \64537 , \50187 , \64536 );
xor \g455974/U$9 ( \64538 , \49781 , \49825 );
xor \g455974/U$9_r1 ( \64539 , \64538 , \49856 );
and \g455974/U$8 ( \64540 , \49984 , \64539 );
xor \g455974/U$11 ( \64541 , \49781 , \49825 );
xor \g455974/U$11_r1 ( \64542 , \64541 , \49856 );
and \g455974/U$10 ( \64543 , \49988 , \64542 );
and \g455974/U$12 ( \64544 , \49984 , \49988 );
or \g455974/U$7 ( \64545 , \64540 , \64543 , \64544 );
not \g128899/U$3 ( \64546 , \64545 );
not \g128937/U$3 ( \64547 , \49675 );
xor \g128969/U$1 ( \64548 , \49749 , \49762 );
not \g128937/U$4 ( \64549 , \64548 );
or \g128937/U$2 ( \64550 , \64547 , \64549 );
or \g128937/U$5 ( \64551 , \64548 , \49675 );
nand \g128937/U$1 ( \64552 , \64550 , \64551 );
not \g128899/U$4 ( \64553 , \64552 );
or \g128899/U$2 ( \64554 , \64546 , \64553 );
or \g128899/U$5 ( \64555 , \64552 , \64545 );
nand \g128899/U$1 ( \64556 , \64554 , \64555 );
not \g128874/U$3 ( \64557 , \64556 );
xor \g455974/U$5 ( \64558 , \49781 , \49825 );
and \g455974/U$4 ( \64559 , \64558 , \49856 );
and \g455974/U$6 ( \64560 , \49781 , \49825 );
or \g455974/U$3 ( \64561 , \64559 , \64560 );
not \g128874/U$4 ( \64562 , \64561 );
and \g128874/U$2 ( \64563 , \64557 , \64562 );
and \g128874/U$5 ( \64564 , \64556 , \64561 );
nor \g128874/U$1 ( \64565 , \64563 , \64564 );
or \g128654/U$2 ( \64566 , \64537 , \64565 );
or \g128654/U$3 ( \64567 , \50187 , \64536 );
nand \g128660/U$1 ( \64568 , \64535 , \64533 , \64532 );
nand \g128654/U$1 ( \64569 , \64566 , \64567 , \64568 );
and \g128650/U$2 ( \64570 , \49777 , \64569 );
or \g128884/U$2 ( \64571 , \64545 , \64561 );
not \g128894/U$3 ( \64572 , \64561 );
not \g128894/U$4 ( \64573 , \64545 );
or \g128894/U$2 ( \64574 , \64572 , \64573 );
nand \g128894/U$1 ( \64575 , \64574 , \64552 );
nand \g128884/U$1 ( \64576 , \64571 , \64575 );
xor \g128653/U$1 ( \64577 , \49777 , \64569 );
and \g128650/U$3 ( \64578 , \64576 , \64577 );
nor \g128656/U$1 ( \64579 , \64537 , \64568 , \64565 );
nor \g128650/U$1 ( \64580 , \64570 , \64578 , \64579 );
xnor \g128649/U$1 ( \64581 , \49658 , \64580 );
nand \g128651/U$1 ( \64582 , \64579 , \64577 , \64576 );
and \g128889/U$2 ( \64583 , \49769 , \49664 );
not \g128896/U$3 ( \64584 , \49769 );
not \g128896/U$4 ( \64585 , \49664 );
and \g128896/U$2 ( \64586 , \64584 , \64585 );
nor \g128896/U$1 ( \64587 , \64586 , \49764 );
nor \g128889/U$1 ( \64588 , \64583 , \64587 );
nor \g128647/U$1 ( \64589 , \64581 , \64582 , \64588 );
not \g128887/U$3 ( \64590 , \49263 );
not \g128887/U$4 ( \64591 , \49654 );
or \g128887/U$2 ( \64592 , \64590 , \64591 );
or \g128893/U$2 ( \64593 , \49654 , \49263 );
nand \g128893/U$1 ( \64594 , \64593 , \49610 );
nand \g128887/U$1 ( \64595 , \64592 , \64594 );
or \g128646/U$2 ( \64596 , \64581 , \64588 );
or \g128646/U$3 ( \64597 , \49658 , \64580 );
nand \g128646/U$1 ( \64598 , \64596 , \64597 , \64582 );
xor \g128645/U$1 ( \64599 , \64595 , \64598 );
not \g129045/U$3 ( \64600 , \49248 );
not \g129045/U$4 ( \64601 , \49190 );
and \g129045/U$2 ( \64602 , \64600 , \64601 );
and \g129065/U$2 ( \64603 , \49248 , \49190 );
nor \g129065/U$1 ( \64604 , \64603 , \49258 );
nor \g129045/U$1 ( \64605 , \64602 , \64604 );
not \g128873/U$3 ( \64606 , \64605 );
and \g128935/U$2 ( \64607 , \49630 , \49616 );
not \g128949/U$3 ( \64608 , \49630 );
not \g128949/U$4 ( \64609 , \49616 );
and \g128949/U$2 ( \64610 , \64608 , \64609 );
nor \g128949/U$1 ( \64611 , \64610 , \49650 );
nor \g128935/U$1 ( \64612 , \64607 , \64611 );
not \g129074/U$3 ( \64613 , \49123 );
not \g129074/U$4 ( \64614 , \49027 );
or \g129074/U$2 ( \64615 , \64613 , \64614 );
or \g129074/U$5 ( \64616 , \49027 , \49123 );
nand \g129074/U$1 ( \64617 , \64615 , \64616 );
not \g129038/U$3 ( \64618 , \64617 );
not \g129038/U$4 ( \64619 , \49084 );
and \g129038/U$2 ( \64620 , \64618 , \64619 );
and \g129038/U$5 ( \64621 , \64617 , \49084 );
nor \g129038/U$1 ( \64622 , \64620 , \64621 );
not \g128987/U$3 ( \64623 , \64622 );
and \g129226/U$2 ( \64624 , \49620 , \49622 );
not \g129238/U$3 ( \64625 , \49620 );
not \g129238/U$4 ( \64626 , \49622 );
and \g129238/U$2 ( \64627 , \64625 , \64626 );
nor \g129238/U$1 ( \64628 , \64627 , \49625 );
nor \g129226/U$1 ( \64629 , \64624 , \64628 );
xnor \g455939/U$1 ( \64630 , \48946 , \48925 );
not \g129158/U$3 ( \64631 , \64630 );
not \g129158/U$4 ( \64632 , \48922 );
and \g129158/U$2 ( \64633 , \64631 , \64632 );
and \g129158/U$5 ( \64634 , \64630 , \48922 );
nor \g129158/U$1 ( \64635 , \64633 , \64634 );
xor \g129102/U$1 ( \64636 , \64629 , \64635 );
not \g128987/U$4 ( \64637 , \64636 );
and \g128987/U$2 ( \64638 , \64623 , \64637 );
and \g128987/U$5 ( \64639 , \64622 , \64636 );
nor \g128987/U$1 ( \64640 , \64638 , \64639 );
xor \g128898/U$1 ( \64641 , \64612 , \64640 );
not \g128873/U$4 ( \64642 , \64641 );
or \g128873/U$2 ( \64643 , \64606 , \64642 );
or \g128873/U$5 ( \64644 , \64641 , \64605 );
nand \g128873/U$1 ( \64645 , \64643 , \64644 );
nand \g128644/U$1 ( \64646 , \64589 , \64599 , \64645 );
not \g128636/U$3 ( \64647 , \64646 );
and \g128642/U$2 ( \64648 , \64595 , \64598 );
and \g128642/U$3 ( \64649 , \64645 , \64599 );
nor \g128642/U$1 ( \64650 , \64648 , \64649 , \64589 );
not \g128883/U$3 ( \64651 , \64612 );
not \g128883/U$4 ( \64652 , \64605 );
and \g128883/U$2 ( \64653 , \64651 , \64652 );
and \g128892/U$2 ( \64654 , \64612 , \64605 );
nor \g128892/U$1 ( \64655 , \64654 , \64640 );
nor \g128883/U$1 ( \64656 , \64653 , \64655 );
or \g128638/U$2 ( \64657 , \64650 , \64656 );
xor \g128957/U$1 ( \64658 , \48920 , \48948 );
xor \g128957/U$1_r1 ( \64659 , \64658 , \49125 );
or \g128986/U$2 ( \64660 , \64635 , \64629 );
and \g128997/U$2 ( \64661 , \64635 , \64629 );
nor \g128997/U$1 ( \64662 , \64661 , \64622 );
not \g128996/U$1 ( \64663 , \64662 );
nand \g128986/U$1 ( \64664 , \64660 , \64663 );
xnor \g128924/U$1 ( \64665 , \64659 , \64664 );
not \g128911/U$3 ( \64666 , \64665 );
not \g129080/U$3 ( \64667 , \49130 );
not \g129080/U$4 ( \64668 , \49142 );
or \g129080/U$2 ( \64669 , \64667 , \64668 );
or \g129080/U$5 ( \64670 , \49142 , \49130 );
nand \g129080/U$1 ( \64671 , \64669 , \64670 );
xor \g455932/U$1 ( \64672 , \49134 , \64671 );
not \g128911/U$4 ( \64673 , \64672 );
and \g128911/U$2 ( \64674 , \64666 , \64673 );
and \g128911/U$5 ( \64675 , \64665 , \64672 );
nor \g128911/U$1 ( \64676 , \64674 , \64675 );
not \g128640/U$2 ( \64677 , \64676 );
xor \g128641/U$1 ( \64678 , \64656 , \64650 );
nand \g128640/U$1 ( \64679 , \64677 , \64678 );
nand \g128638/U$1 ( \64680 , \64657 , \64679 );
not \g128636/U$4 ( \64681 , \64680 );
or \g128636/U$2 ( \64682 , \64647 , \64681 );
or \g128636/U$5 ( \64683 , \64680 , \64646 );
nand \g128636/U$1 ( \64684 , \64682 , \64683 );
not \g128921/U$3 ( \64685 , \64672 );
not \g128921/U$4 ( \64686 , \64659 );
or \g128921/U$2 ( \64687 , \64685 , \64686 );
or \g128922/U$2 ( \64688 , \64659 , \64672 );
nand \g128922/U$1 ( \64689 , \64688 , \64664 );
nand \g128921/U$1 ( \64690 , \64687 , \64689 );
and \g128632/U$2 ( \64691 , \64684 , \64690 );
not \g128878/U$3 ( \64692 , \49144 );
not \g128905/U$3 ( \64693 , \49128 );
not \g128905/U$4 ( \64694 , \49155 );
or \g128905/U$2 ( \64695 , \64693 , \64694 );
or \g128905/U$5 ( \64696 , \49155 , \49128 );
nand \g128905/U$1 ( \64697 , \64695 , \64696 );
not \g128878/U$4 ( \64698 , \64697 );
or \g128878/U$2 ( \64699 , \64692 , \64698 );
or \g128878/U$5 ( \64700 , \64697 , \49144 );
nand \g128878/U$1 ( \64701 , \64699 , \64700 );
xor \g128635/U$1 ( \64702 , \64690 , \64684 );
and \g128634/U$2 ( \64703 , \64701 , \64702 );
nor \g128637/U$1 ( \64704 , \64679 , \64646 );
nor \g128632/U$1 ( \64705 , \64691 , \64703 , \64704 );
xnor \g128631/U$1 ( \64706 , \49157 , \64705 );
not \g128901/U$3 ( \64707 , \48912 );
not \g128901/U$4 ( \64708 , \48884 );
or \g128901/U$2 ( \64709 , \64707 , \64708 );
or \g128901/U$5 ( \64710 , \48884 , \48912 );
nand \g128901/U$1 ( \64711 , \64709 , \64710 );
not \g128871/U$3 ( \64712 , \64711 );
not \g128871/U$4 ( \64713 , \48886 );
and \g128871/U$2 ( \64714 , \64712 , \64713 );
and \g128871/U$5 ( \64715 , \64711 , \48886 );
nor \g128871/U$1 ( \64716 , \64714 , \64715 );
or \g128628/U$2 ( \64717 , \64706 , \64716 );
or \g128628/U$3 ( \64718 , \49157 , \64705 );
nand \g128633/U$1 ( \64719 , \64704 , \64703 );
nand \g128628/U$1 ( \64720 , \64717 , \64718 , \64719 );
xor \g128627/U$1 ( \64721 , \48914 , \64720 );
and \g128624/U$2 ( \64722 , \48882 , \64721 );
and \g128624/U$3 ( \64723 , \48914 , \64720 );
nor \g128630/U$1 ( \64724 , \64706 , \64719 , \64716 );
nor \g128624/U$1 ( \64725 , \64722 , \64723 , \64724 );
not \g129006/U$1 ( \64726 , \48702 );
and \g128909/U$2 ( \64727 , \48705 , \64726 );
not \g128917/U$3 ( \64728 , \48705 );
not \g128917/U$4 ( \64729 , \64726 );
and \g128917/U$2 ( \64730 , \64728 , \64729 );
nor \g128917/U$1 ( \64731 , \64730 , \48874 );
nor \g128909/U$1 ( \64732 , \64727 , \64731 );
or \g128620/U$2 ( \64733 , \64725 , \64732 );
not \g128972/U$3 ( \64734 , \48556 );
not \g128972/U$4 ( \64735 , \48640 );
or \g128972/U$2 ( \64736 , \64734 , \64735 );
or \g128972/U$5 ( \64737 , \48640 , \48556 );
nand \g128972/U$1 ( \64738 , \64736 , \64737 );
not \g128942/U$3 ( \64739 , \64738 );
not \g128942/U$4 ( \64740 , \48558 );
and \g128942/U$2 ( \64741 , \64739 , \64740 );
and \g128942/U$5 ( \64742 , \64738 , \48558 );
nor \g128942/U$1 ( \64743 , \64741 , \64742 );
xnor \g128623/U$1 ( \64744 , \64732 , \64725 );
or \g128620/U$3 ( \64745 , \64743 , \64744 );
nand \g128626/U$1 ( \64746 , \64724 , \64721 , \48882 );
nand \g128620/U$1 ( \64747 , \64733 , \64745 , \64746 );
and \g128616/U$2 ( \64748 , \48642 , \64747 );
xor \g129116/U$1 ( \64749 , \48424 , \48428 );
xor \g129116/U$1_r1 ( \64750 , \64749 , \48431 );
not \g128946/U$3 ( \64751 , \64750 );
xor \g129018/U$4 ( \64752 , \48493 , \48503 );
and \g129018/U$3 ( \64753 , \64752 , \48555 );
and \g129018/U$5 ( \64754 , \48493 , \48503 );
or \g129018/U$2 ( \64755 , \64753 , \64754 );
not \g129084/U$3 ( \64756 , \48412 );
not \g129084/U$4 ( \64757 , \48342 );
and \g129084/U$2 ( \64758 , \64756 , \64757 );
and \g129084/U$5 ( \64759 , \48412 , \48342 );
nor \g129084/U$1 ( \64760 , \64758 , \64759 );
not \g129035/U$3 ( \64761 , \64760 );
not \g129035/U$4 ( \64762 , \48277 );
and \g129035/U$2 ( \64763 , \64761 , \64762 );
and \g129035/U$5 ( \64764 , \64760 , \48277 );
nor \g129035/U$1 ( \64765 , \64763 , \64764 );
xor \g128976/U$1 ( \64766 , \64755 , \64765 );
not \g128946/U$4 ( \64767 , \64766 );
or \g128946/U$2 ( \64768 , \64751 , \64767 );
or \g128946/U$5 ( \64769 , \64766 , \64750 );
nand \g128946/U$1 ( \64770 , \64768 , \64769 );
xor \g128619/U$1 ( \64771 , \48642 , \64747 );
and \g128616/U$3 ( \64772 , \64770 , \64771 );
nor \g128622/U$1 ( \64773 , \64744 , \64746 , \64743 );
nor \g128616/U$1 ( \64774 , \64748 , \64772 , \64773 );
xnor \g128615/U$1 ( \64775 , \48438 , \64774 );
not \g128952/U$3 ( \64776 , \64755 );
not \g128952/U$4 ( \64777 , \64750 );
and \g128952/U$2 ( \64778 , \64776 , \64777 );
and \g128961/U$2 ( \64779 , \64755 , \64750 );
nor \g128961/U$1 ( \64780 , \64779 , \64765 );
nor \g128952/U$1 ( \64781 , \64778 , \64780 );
or \g128612/U$2 ( \64782 , \64775 , \64781 );
or \g128612/U$3 ( \64783 , \48438 , \64774 );
nand \g128618/U$1 ( \64784 , \64773 , \64771 , \64770 );
nand \g128612/U$1 ( \64785 , \64782 , \64783 , \64784 );
and \g128608/U$2 ( \64786 , \48264 , \64785 );
or \g128981/U$2 ( \64787 , \48268 , \48434 );
not \g128991/U$3 ( \64788 , \48434 );
not \g128991/U$4 ( \64789 , \48268 );
or \g128991/U$2 ( \64790 , \64788 , \64789 );
nand \g128991/U$1 ( \64791 , \64790 , \48415 );
nand \g128981/U$1 ( \64792 , \64787 , \64791 );
xor \g128611/U$1 ( \64793 , \48264 , \64785 );
and \g128608/U$3 ( \64794 , \64792 , \64793 );
nor \g128613/U$1 ( \64795 , \64775 , \64784 , \64781 );
nor \g128608/U$1 ( \64796 , \64786 , \64794 , \64795 );
not \g128983/U$3 ( \64797 , \48221 );
not \g128983/U$4 ( \64798 , \48171 );
and \g128983/U$2 ( \64799 , \64797 , \64798 );
and \g128993/U$2 ( \64800 , \48221 , \48171 );
nor \g128993/U$1 ( \64801 , \64800 , \48259 );
nor \g128983/U$1 ( \64802 , \64799 , \64801 );
or \g128604/U$2 ( \64803 , \64796 , \64802 );
not \g129184/U$3 ( \64804 , \48232 );
not \g129184/U$4 ( \64805 , \48077 );
and \g129184/U$2 ( \64806 , \64804 , \64805 );
and \g129204/U$2 ( \64807 , \48232 , \48077 );
nor \g129204/U$1 ( \64808 , \64807 , \48238 );
nor \g129184/U$1 ( \64809 , \64806 , \64808 );
xor \g129115/U$1 ( \64810 , \48073 , \48083 );
xor \g129115/U$1_r1 ( \64811 , \64810 , \48086 );
xnor \g129081/U$1 ( \64812 , \64809 , \64811 );
not \g128989/U$3 ( \64813 , \64812 );
or \g129090/U$2 ( \64814 , \48223 , \48255 );
not \g129100/U$3 ( \64815 , \48255 );
not \g129100/U$4 ( \64816 , \48223 );
or \g129100/U$2 ( \64817 , \64815 , \64816 );
nand \g129100/U$1 ( \64818 , \64817 , \48246 );
nand \g129090/U$1 ( \64819 , \64814 , \64818 );
not \g128989/U$4 ( \64820 , \64819 );
and \g128989/U$2 ( \64821 , \64813 , \64820 );
and \g128989/U$5 ( \64822 , \64812 , \64819 );
nor \g128989/U$1 ( \64823 , \64821 , \64822 );
xnor \g128607/U$1 ( \64824 , \64802 , \64796 );
or \g128604/U$3 ( \64825 , \64823 , \64824 );
nand \g128609/U$1 ( \64826 , \64795 , \64793 , \64792 );
nand \g128604/U$1 ( \64827 , \64803 , \64825 , \64826 );
and \g128600/U$2 ( \64828 , \48101 , \64827 );
or \g128985/U$2 ( \64829 , \64811 , \64809 );
not \g128994/U$3 ( \64830 , \64809 );
not \g128994/U$4 ( \64831 , \64811 );
or \g128994/U$2 ( \64832 , \64830 , \64831 );
nand \g128994/U$1 ( \64833 , \64832 , \64819 );
nand \g128985/U$1 ( \64834 , \64829 , \64833 );
xor \g128603/U$1 ( \64835 , \48101 , \64827 );
and \g128600/U$3 ( \64836 , \64834 , \64835 );
nor \g128606/U$1 ( \64837 , \64824 , \64826 , \64823 );
nor \g128600/U$1 ( \64838 , \64828 , \64836 , \64837 );
xnor \g128599/U$1 ( \64839 , \48091 , \64838 );
and \g129189/U$2 ( \64840 , \47939 , \47982 );
not \g129207/U$3 ( \64841 , \47939 );
not \g129207/U$4 ( \64842 , \47982 );
and \g129207/U$2 ( \64843 , \64841 , \64842 );
nor \g129207/U$1 ( \64844 , \64843 , \48009 );
nor \g129189/U$1 ( \64845 , \64840 , \64844 );
not \g129082/U$3 ( \64846 , \64845 );
and \g129627/U$2 ( \64847 , \47970 , \47959 );
and \g129627/U$3 ( \64848 , \47960 , \47962 );
nor \g129627/U$1 ( \64849 , \64847 , \64848 );
not \g129580/U$3 ( \64850 , \64849 );
not \g129580/U$4 ( \64851 , \47948 );
and \g129580/U$2 ( \64852 , \64850 , \64851 );
and \g129580/U$5 ( \64853 , \64849 , \47948 );
nor \g129580/U$1 ( \64854 , \64852 , \64853 );
not \g129147/U$3 ( \64855 , \64854 );
not \g129180/U$3 ( \64856 , \47940 );
nand \g129818/U$1 ( \64857 , \40061 , \47950 );
xor \g129265/U$1 ( \64858 , \64857 , \47935 );
and \g129400/U$2 ( \64859 , \47894 , \47913 );
and \g129400/U$3 ( \64860 , \47914 , \47972 );
nor \g129400/U$1 ( \64861 , \64859 , \64860 );
not \g129348/U$3 ( \64862 , \64861 );
not \g129348/U$4 ( \64863 , \47976 );
and \g129348/U$2 ( \64864 , \64862 , \64863 );
and \g129348/U$5 ( \64865 , \64861 , \47976 );
nor \g129348/U$1 ( \64866 , \64864 , \64865 );
xor \g129265/U$1_r1 ( \64867 , \64858 , \64866 );
not \g129180/U$4 ( \64868 , \64867 );
or \g129180/U$2 ( \64869 , \64856 , \64868 );
or \g129180/U$5 ( \64870 , \64867 , \47940 );
nand \g129180/U$1 ( \64871 , \64869 , \64870 );
not \g129147/U$4 ( \64872 , \64871 );
or \g129147/U$2 ( \64873 , \64855 , \64872 );
or \g129147/U$5 ( \64874 , \64871 , \64854 );
nand \g129147/U$1 ( \64875 , \64873 , \64874 );
not \g129082/U$4 ( \64876 , \64875 );
or \g129082/U$2 ( \64877 , \64846 , \64876 );
or \g129082/U$5 ( \64878 , \64875 , \64845 );
nand \g129082/U$1 ( \64879 , \64877 , \64878 );
not \g129043/U$3 ( \64880 , \64879 );
xor \g456000/U$4 ( \64881 , \47944 , \47968 );
and \g456000/U$3 ( \64882 , \64881 , \47981 );
and \g456000/U$5 ( \64883 , \47944 , \47968 );
nor \g456000/U$2 ( \64884 , \64882 , \64883 );
not \g129043/U$4 ( \64885 , \64884 );
and \g129043/U$2 ( \64886 , \64880 , \64885 );
and \g129043/U$5 ( \64887 , \64879 , \64884 );
nor \g129043/U$1 ( \64888 , \64886 , \64887 );
or \g128596/U$2 ( \64889 , \64839 , \64888 );
or \g128596/U$3 ( \64890 , \48091 , \64838 );
nand \g128601/U$1 ( \64891 , \64837 , \64835 , \64834 );
nand \g128596/U$1 ( \64892 , \64889 , \64890 , \64891 );
xor \g129265/U$4 ( \64893 , \64857 , \47935 );
and \g129265/U$3 ( \64894 , \64893 , \64866 );
and \g129265/U$5 ( \64895 , \64857 , \47935 );
or \g129265/U$2 ( \64896 , \64894 , \64895 );
not \g129036/U$3 ( \64897 , \64896 );
not \g129478/U$3 ( \64898 , \47948 );
and \g129519/U$2 ( \64899 , \47970 , \47960 );
and \g129519/U$3 ( \64900 , \47959 , \47972 );
nor \g129519/U$1 ( \64901 , \64899 , \64900 );
not \g129478/U$4 ( \64902 , \64901 );
or \g129478/U$2 ( \64903 , \64898 , \64902 );
or \g129478/U$5 ( \64904 , \64901 , \47948 );
nand \g129478/U$1 ( \64905 , \64903 , \64904 );
not \g135511/U$2 ( \64906 , \47962 );
nor \g135511/U$1 ( \64907 , \64906 , \40060 );
xor \g129281/U$1 ( \64908 , \64905 , \64907 );
and \g129361/U$2 ( \64909 , \47916 , \47977 );
and \g129361/U$3 ( \64910 , \47915 , \47976 );
nor \g129361/U$1 ( \64911 , \64909 , \64910 );
xor \g129281/U$1_r1 ( \64912 , \64908 , \64911 );
not \g129083/U$3 ( \64913 , \64912 );
not \g129190/U$3 ( \64914 , \47939 );
not \g129190/U$4 ( \64915 , \64854 );
and \g129190/U$2 ( \64916 , \64914 , \64915 );
and \g129208/U$2 ( \64917 , \47939 , \64854 );
nor \g129208/U$1 ( \64918 , \64917 , \64867 );
nor \g129190/U$1 ( \64919 , \64916 , \64918 );
not \g129083/U$4 ( \64920 , \64919 );
or \g129083/U$2 ( \64921 , \64913 , \64920 );
or \g129083/U$5 ( \64922 , \64919 , \64912 );
nand \g129083/U$1 ( \64923 , \64921 , \64922 );
not \g129036/U$4 ( \64924 , \64923 );
or \g129036/U$2 ( \64925 , \64897 , \64924 );
or \g129036/U$5 ( \64926 , \64923 , \64896 );
nand \g129036/U$1 ( \64927 , \64925 , \64926 );
and \g128592/U$2 ( \64928 , \64892 , \64927 );
or \g129051/U$2 ( \64929 , \64845 , \64884 );
not \g129070/U$3 ( \64930 , \64884 );
not \g129070/U$4 ( \64931 , \64845 );
or \g129070/U$2 ( \64932 , \64930 , \64931 );
nand \g129070/U$1 ( \64933 , \64932 , \64875 );
nand \g129051/U$1 ( \64934 , \64929 , \64933 );
xor \g128595/U$1 ( \64935 , \64927 , \64892 );
and \g128594/U$2 ( \64936 , \64934 , \64935 );
nor \g128598/U$1 ( \64937 , \64839 , \64891 , \64888 );
nor \g128592/U$1 ( \64938 , \64928 , \64936 , \64937 );
nand \g128591/U$1 ( \64939 , \47916 , \64938 );
not \g129360/U$1 ( \64940 , \64911 );
xor \g129281/U$4 ( \64941 , \64905 , \64907 );
and \g129281/U$3 ( \64942 , \64941 , \64911 );
and \g129281/U$5 ( \64943 , \64905 , \64907 );
or \g129281/U$2 ( \64944 , \64942 , \64943 );
xor \g455991/U$1 ( \64945 , \64940 , \64944 );
nand \g129648/U$1 ( \64946 , \40061 , \47970 );
not \g129270/U$3 ( \64947 , \64946 );
not \g129330/U$3 ( \64948 , \47948 );
and \g129388/U$2 ( \64949 , \47894 , \47959 );
and \g129388/U$3 ( \64950 , \47960 , \47972 );
nor \g129388/U$1 ( \64951 , \64949 , \64950 );
not \g129330/U$4 ( \64952 , \64951 );
or \g129330/U$2 ( \64953 , \64948 , \64952 );
or \g129330/U$5 ( \64954 , \64951 , \47948 );
nand \g129330/U$1 ( \64955 , \64953 , \64954 );
and \g129301/U$2 ( \64956 , \64955 , \64911 );
not \g129301/U$4 ( \64957 , \64955 );
and \g129301/U$3 ( \64958 , \64957 , \64940 );
nor \g129301/U$1 ( \64959 , \64956 , \64958 );
not \g129270/U$4 ( \64960 , \64959 );
or \g129270/U$2 ( \64961 , \64947 , \64960 );
or \g129270/U$5 ( \64962 , \64959 , \64946 );
nand \g129270/U$1 ( \64963 , \64961 , \64962 );
xor \g455991/U$1_r1 ( \64964 , \64945 , \64963 );
not \g128587/U$3 ( \64965 , \64964 );
or \g128590/U$2 ( \64966 , \64938 , \47916 );
nand \g128590/U$1 ( \64967 , \64966 , \64939 );
not \g128587/U$4 ( \64968 , \64967 );
or \g128587/U$2 ( \64969 , \64965 , \64968 );
xnor \g128589/U$1 ( \64970 , \64964 , \64967 );
not \g129264/U$1 ( \64971 , \64896 );
and \g129086/U$2 ( \64972 , \64912 , \64971 );
not \g129097/U$3 ( \64973 , \64912 );
not \g129097/U$4 ( \64974 , \64971 );
and \g129097/U$2 ( \64975 , \64973 , \64974 );
nor \g129097/U$1 ( \64976 , \64975 , \64919 );
nor \g129086/U$1 ( \64977 , \64972 , \64976 );
or \g128587/U$5 ( \64978 , \64970 , \64977 );
nand \g128587/U$1 ( \64979 , \64969 , \64978 );
and \g128586/U$2 ( \64980 , \64939 , \64979 );
not \g128583/U$4 ( \64981 , \64980 );
or \g128583/U$2 ( \64982 , \47896 , \64981 );
or \g128583/U$5 ( \64983 , \64980 , \47895 );
nand \g128583/U$1 ( \64984 , \64982 , \64983 );
not \g128582/U$3 ( \64985 , \64984 );
nand \g129428/U$1 ( \64986 , \47960 , \47894 );
not \g129383/U$3 ( \64987 , \64986 );
not \g129383/U$4 ( \64988 , \47948 );
and \g129383/U$2 ( \64989 , \64987 , \64988 );
and \g129383/U$5 ( \64990 , \64986 , \47948 );
nor \g129383/U$1 ( \64991 , \64989 , \64990 );
or \g129285/U$2 ( \64992 , \64940 , \64946 );
not \g129647/U$1 ( \64993 , \64946 );
or \g129285/U$3 ( \64994 , \64993 , \64911 );
nand \g129285/U$1 ( \64995 , \64992 , \64994 , \64955 );
xor \g455992/U$5 ( \64996 , \64991 , \64995 );
nor \g129608/U$1 ( \64997 , \64946 , \47976 );
not \g455992/U$6 ( \64998 , \64997 );
and \g455992/U$4 ( \64999 , \64996 , \64998 );
and \g455992/U$7 ( \65000 , \64991 , \64995 );
or \g455992/U$3 ( \65001 , \64999 , \65000 );
not \g3/U$1 ( \65002 , \65001 );
not \g128582/U$4 ( \65003 , \65002 );
and \g128582/U$2 ( \65004 , \64985 , \65003 );
and \g128582/U$5 ( \65005 , \64984 , \65002 );
nor \g128582/U$1 ( \65006 , \65004 , \65005 );
not \g128571/U$3 ( \65007 , \65006 );
xor \g128586/U$1 ( \65008 , \64939 , \64979 );
not \g128585/U$2 ( \65009 , \65008 );
nand \g128593/U$1 ( \65010 , \64937 , \64936 );
nand \g128585/U$1 ( \65011 , \65009 , \65010 );
and \g129268/U$2 ( \65012 , \47976 , \64940 );
and \g129268/U$3 ( \65013 , \64946 , \64911 );
nor \g129268/U$1 ( \65014 , \65012 , \65013 , \64997 );
and \g128578/U$2 ( \65015 , \65011 , \65014 );
not \g135510/U$2 ( \65016 , \47972 );
nor \g135510/U$1 ( \65017 , \65016 , \40060 );
not \g128581/U$3 ( \65018 , \65014 );
not \g128584/U$3 ( \65019 , \65008 );
not \g128584/U$4 ( \65020 , \65010 );
and \g128584/U$2 ( \65021 , \65019 , \65020 );
and \g128584/U$5 ( \65022 , \65008 , \65010 );
nor \g128584/U$1 ( \65023 , \65021 , \65022 );
not \g128581/U$4 ( \65024 , \65023 );
or \g128581/U$2 ( \65025 , \65018 , \65024 );
or \g128581/U$5 ( \65026 , \65023 , \65014 );
nand \g128581/U$1 ( \65027 , \65025 , \65026 );
and \g128578/U$3 ( \65028 , \65017 , \65027 );
nor \g128578/U$1 ( \65029 , \65015 , \65028 );
not \g128572/U$3 ( \65030 , \65029 );
not \g128573/U$3 ( \65031 , \47948 );
xor \g455991/U$4 ( \65032 , \64940 , \64944 );
and \g455991/U$3 ( \65033 , \65032 , \64963 );
and \g455991/U$5 ( \65034 , \64940 , \64944 );
nor \g455991/U$2 ( \65035 , \65033 , \65034 );
not \g128575/U$3 ( \65036 , \65035 );
xor \g455992/U$1 ( \65037 , \64991 , \64995 );
not \g455992/U$2 ( \65038 , \64997 );
xor \g455992/U$1_r1 ( \65039 , \65037 , \65038 );
not \g128575/U$4 ( \65040 , \65039 );
and \g128575/U$2 ( \65041 , \65036 , \65040 );
and \g128577/U$2 ( \65042 , \65035 , \65039 );
xnor \g128580/U$1 ( \65043 , \65017 , \65027 );
nor \g128577/U$1 ( \65044 , \65042 , \65043 );
nor \g128575/U$1 ( \65045 , \65041 , \65044 );
not \g128573/U$4 ( \65046 , \65045 );
or \g128573/U$2 ( \65047 , \65031 , \65046 );
or \g128573/U$5 ( \65048 , \65045 , \47948 );
nand \g128573/U$1 ( \65049 , \65047 , \65048 );
not \g128572/U$4 ( \65050 , \65049 );
or \g128572/U$2 ( \65051 , \65030 , \65050 );
or \g128572/U$5 ( \65052 , \65049 , \65029 );
nand \g128572/U$1 ( \65053 , \65051 , \65052 );
not \g128571/U$4 ( \65054 , \65053 );
or \g128571/U$2 ( \65055 , \65007 , \65054 );
or \g128571/U$5 ( \65056 , \65053 , \65006 );
nand \g128571/U$1 ( \65057 , \65055 , \65056 );
not \g128574/U$3 ( \65058 , \65035 );
xor \g455928/U$1 ( \65059 , \65039 , \65043 );
not \g128574/U$4 ( \65060 , \65059 );
or \g128574/U$2 ( \65061 , \65058 , \65060 );
or \g128574/U$5 ( \65062 , \65059 , \65035 );
nand \g128574/U$1 ( \65063 , \65061 , \65062 );
xor \g128588/U$1 ( \65064 , \64977 , \64970 );
xor \g128594/U$1 ( \65065 , \64934 , \64935 );
xor \g128597/U$1 ( \65066 , \64888 , \64839 );
xor \g128602/U$1 ( \65067 , \64834 , \64835 );
xor \g128605/U$1 ( \65068 , \64823 , \64824 );
xor \g128610/U$1 ( \65069 , \64792 , \64793 );
xor \g128614/U$1 ( \65070 , \64781 , \64775 );
xor \g128617/U$1 ( \65071 , \64770 , \64771 );
xor \g128621/U$1 ( \65072 , \64743 , \64744 );
xor \g128625/U$1 ( \65073 , \48882 , \64721 );
xor \g128629/U$1 ( \65074 , \64716 , \64706 );
xor \g128634/U$1 ( \65075 , \64701 , \64702 );
not \g128639/U$3 ( \65076 , \64676 );
not \g128639/U$4 ( \65077 , \64678 );
or \g128639/U$2 ( \65078 , \65076 , \65077 );
or \g128639/U$5 ( \65079 , \64678 , \64676 );
nand \g128639/U$1 ( \65080 , \65078 , \65079 );
xor \g128643/U$1 ( \65081 , \64645 , \64599 );
xor \g128648/U$1 ( \65082 , \64588 , \64581 );
xor \g128652/U$1 ( \65083 , \64576 , \64577 );
xor \g128655/U$1 ( \65084 , \64565 , \64537 );
xor \g128659/U$1 ( \65085 , \64532 , \64533 );
xor \g128663/U$1 ( \65086 , \64521 , \64511 );
xor \g128667/U$1 ( \65087 , \50806 , \64506 );
xor \g128671/U$1 ( \65088 , \64501 , \64491 );
xor \g128675/U$1 ( \65089 , \64486 , \64487 );
xor \g128680/U$1 ( \65090 , \64475 , \64476 );
xor \g128683/U$1 ( \65091 , \51769 , \64454 );
xor \g128687/U$1 ( \65092 , \64449 , \64450 );
xor \g128691/U$1 ( \65093 , \64430 , \64431 );
xor \g128696/U$1 ( \65094 , \64409 , \64405 );
xor \g128700/U$1 ( \65095 , \64393 , \64374 );
xor \g128706/U$1 ( \65096 , \64369 , \64370 );
xor \g128711/U$1 ( \65097 , \64351 , \64352 );
xor \g128714/U$1 ( \65098 , \64323 , \64273 );
xor \g128718/U$1 ( \65099 , \53734 , \64268 );
xor \g128722/U$1 ( \65100 , \64263 , \64264 );
xor \g128726/U$1 ( \65101 , \64250 , \64251 );
xor \g128730/U$1 ( \65102 , \64223 , \64224 );
xor \g128735/U$1 ( \65103 , \64201 , \64202 );
not \g128740/U$3 ( \65104 , \64156 );
not \g128740/U$4 ( \65105 , \64158 );
or \g128740/U$2 ( \65106 , \65104 , \65105 );
or \g128740/U$5 ( \65107 , \64158 , \64156 );
nand \g128740/U$1 ( \65108 , \65106 , \65107 );
xor \g128744/U$1 ( \65109 , \64104 , \64049 );
xor \g128748/U$1 ( \65110 , \64040 , \63921 );
xor \g128752/U$1 ( \65111 , \55588 , \63916 );
xor \g128756/U$1 ( \65112 , \63911 , \63912 );
xor \g128762/U$1 ( \65113 , \56048 , \63886 );
xor \g128767/U$1 ( \65114 , \63881 , \63882 );
xor \g128770/U$1 ( \65115 , \63863 , \63864 );
xor \g128774/U$1 ( \65116 , \63828 , \63829 );
xor \g128777/U$1 ( \65117 , \63792 , \63793 );
xor \g128782/U$1 ( \65118 , \63715 , \63716 );
xor \g128786/U$1 ( \65119 , \63627 , \63628 );
not \g128792/U$3 ( \65120 , \63474 );
not \g128792/U$4 ( \65121 , \63267 );
or \g128792/U$2 ( \65122 , \65120 , \65121 );
or \g128792/U$5 ( \65123 , \63267 , \63474 );
nand \g128792/U$1 ( \65124 , \65122 , \65123 );
xor \g128796/U$1 ( \65125 , \63258 , \63259 );
xor \g128800/U$1 ( \65126 , \63030 , \63031 );
xor \g128803/U$1 ( \65127 , \62797 , \62798 );
not \g128806/U$3 ( \65128 , \62554 );
not \g128806/U$4 ( \65129 , \62556 );
or \g128806/U$2 ( \65130 , \65128 , \65129 );
or \g128806/U$5 ( \65131 , \62556 , \62554 );
nand \g128806/U$1 ( \65132 , \65130 , \65131 );
not \g128811/U$3 ( \65133 , \62291 );
not \g128811/U$4 ( \65134 , \62293 );
or \g128811/U$2 ( \65135 , \65133 , \65134 );
or \g128811/U$5 ( \65136 , \62293 , \62291 );
nand \g128811/U$1 ( \65137 , \65135 , \65136 );
not \g128817/U$3 ( \65138 , \62012 );
not \g128817/U$4 ( \65139 , \61747 );
or \g128817/U$2 ( \65140 , \65138 , \65139 );
or \g128817/U$5 ( \65141 , \61747 , \62012 );
nand \g128817/U$1 ( \65142 , \65140 , \65141 );
xor \g128830/U$1 ( \65143 , \61719 , \61731 );
not \g128934/U$3 ( \65144 , \61460 );
not \g128934/U$4 ( \65145 , \61220 );
or \g128934/U$2 ( \65146 , \65144 , \65145 );
or \g128934/U$5 ( \65147 , \61220 , \61460 );
nand \g128934/U$1 ( \65148 , \65146 , \65147 );
xor \g129106/U$1 ( \65149 , \61210 , \61211 );
not \g129316/U$3 ( \65150 , \61189 );
not \g129316/U$4 ( \65151 , \61172 );
or \g129316/U$2 ( \65152 , \65150 , \65151 );
or \g129316/U$5 ( \65153 , \61172 , \61189 );
nand \g129316/U$1 ( \65154 , \65152 , \65153 );
not \g129380/U$3 ( \65155 , \52389 );
not \g129380/U$4 ( \65156 , \51120 );
xor \g129524/U$1 ( \65157 , \61146 , \61150 );
xor \g129524/U$1_r1 ( \65158 , \65157 , \61156 );
not \g130133/U$3 ( \65159 , \60986 );
not \g130133/U$4 ( \65160 , \60989 );
or \g130133/U$2 ( \65161 , \65159 , \65160 );
or \g130133/U$5 ( \65162 , \60989 , \60986 );
nand \g130133/U$1 ( \65163 , \65161 , \65162 );
xor \g130280/U$1 ( \65164 , \60959 , \60967 );
xor \g130280/U$1_r1 ( \65165 , \65164 , \60970 );
xor \g130452/U$1 ( \65166 , \60678 , \60680 );
xor \g130744/U$1 ( \65167 , \60287 , \60289 );
xor \g130996/U$1 ( \65168 , \59902 , \59904 );
xor \g131306/U$1 ( \65169 , \59543 , \59545 );
xor \g131587/U$1 ( \65170 , \59208 , \59210 );
xor \g131861/U$1 ( \65171 , \58905 , \58907 );
xor \g132210/U$1 ( \65172 , \58630 , \58632 );
xor \g132437/U$1 ( \65173 , \58503 , \58504 );
xor \g132437/U$1_r1 ( \65174 , \65173 , \58507 );
xor \g132556/U$1 ( \65175 , \58498 , \58502 );
xor \g132586/U$1 ( \65176 , \58489 , \58490 );
xor \g132586/U$1_r1 ( \65177 , \65176 , \58495 );
xor \g132698/U$1 ( \65178 , \58486 , \58488 );
xor \g132770/U$1 ( \65179 , \58480 , \57528 );
xor \g132770/U$1_r1 ( \65180 , \65179 , \58483 );
xor \g132866/U$1 ( \65181 , \58477 , \58479 );
xor \g132891/U$1 ( \65182 , \58470 , \58471 );
xor \g132891/U$1_r1 ( \65183 , \65182 , \58474 );
xor \g132977/U$1 ( \65184 , \58437 , \58469 );
xor \g133030/U$1 ( \65185 , \58460 , \58461 );
xor \g133030/U$1_r1 ( \65186 , \65185 , \58466 );
xor \g133108/U$1 ( \65187 , \58457 , \58459 );
xor \g133150/U$1 ( \65188 , \58450 , \58451 );
xor \g133150/U$1_r1 ( \65189 , \65188 , \58454 );
xor \g133249/U$1 ( \65190 , \58447 , \58449 );
xor \g133351/U$1 ( \65191 , \58441 , \58031 );
xor \g133351/U$1_r1 ( \65192 , \65191 , \58444 );
xor \g133477/U$1 ( \65193 , \58438 , \58440 );
xor \g456026/U$2 ( \65194 , \61085 , \61093 );
xor \g456026/U$1 ( \65195 , \65194 , \61110 );
xor \g456026/U$1_r1 ( \65196 , \61073 , \61117 );
xor \g456026/U$1_r2 ( \65197 , \65195 , \65196 );
xor \g456037/U$2 ( \65198 , \61033 , \61037 );
xor \g456037/U$1 ( \65199 , \65198 , \61050 );
xor \g456037/U$1_r1 ( \65200 , \61001 , \61062 );
xor \g456037/U$1_r2 ( \65201 , \65199 , \65200 );
xor \g456077/U$2 ( \65202 , \60366 , \60374 );
xor \g456077/U$1 ( \65203 , \65202 , \60481 );
xor \g456077/U$1_r1 ( \65204 , \60493 , \60498 );
xor \g456077/U$1_r2 ( \65205 , \65203 , \65204 );
xor \g456091/U$2 ( \65206 , \59981 , \59989 );
xor \g456091/U$1 ( \65207 , \65206 , \60086 );
xor \g456091/U$1_r1 ( \65208 , \60094 , \60099 );
xor \g456091/U$1_r2 ( \65209 , \65207 , \65208 );
xor \g456101/U$2 ( \65210 , \59553 , \59628 );
xor \g456101/U$1 ( \65211 , \65210 , \59705 );
xor \g456101/U$1_r1 ( \65212 , \59713 , \59718 );
xor \g456101/U$1_r2 ( \65213 , \65211 , \65212 );
xor \g456121/U$2 ( \65214 , \59510 , \59514 );
xor \g456121/U$1 ( \65215 , \65214 , \59519 );
xor \g456121/U$1_r1 ( \65216 , \59506 , \59523 );
xor \g456121/U$1_r2 ( \65217 , \65215 , \65216 );
xor \g456139/U$2 ( \65218 , \58998 , \59006 );
xor \g456139/U$1 ( \65219 , \65218 , \59039 );
xor \g456139/U$1_r1 ( \65220 , \59051 , \59056 );
xor \g456139/U$1_r2 ( \65221 , \65219 , \65220 );
xor \g456153/U$2 ( \65222 , \58653 , \58657 );
xor \g456153/U$1 ( \65223 , \65222 , \58746 );
xor \g456153/U$1_r1 ( \65224 , \58758 , \58763 );
xor \g456153/U$1_r2 ( \65225 , \65223 , \65224 );
endmodule

