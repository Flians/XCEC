//
// Conformal-LEC Version 20.10-d214 (03-Sep-2020)
//
module top(RIb54a900_11,RIb54a888_10,RIb54a810_9,RIb54a798_8,RIb54a720_7,RIb54a6a8_6,RIb54a630_5,RIb54a5b8_4,RIb54a540_3,
        RIb54a4c8_2,RIb54a450_1,RIb5517a0_247,RIb551980_251,RIb54ab58_16,RIb54abd0_17,RIb54aae0_15,RIb54aa68_14,RIb54a9f0_13,RIb551908_250,
        RIb551b60_255,RIb551ae8_254,RIb551f98_264,RIb551f20_263,RIb551cc8_258,RIb551c50_257,RIb551bd8_256,RIb551890_249,RIb551818_248,RIb551ea8_262,
        RIb551e30_261,RIb551db8_260,RIb551d40_259,RIb5519f8_252,RIb551a70_253,RIb54ad38_20,RIb54acc0_19,RIb54af18_24,RIb54aea0_23,RIb54b350_33,
        RIb54b2d8_32,RIb54af90_25,RIb54b008_26,RIb54b080_27,RIb54ac48_18,RIb54a978_12,RIb54b260_31,RIb54b1e8_30,RIb54b170_29,RIb54b0f8_28,
        RIb54adb0_21,RIb54ae28_22,RIb54b968_46,RIb54b8f0_45,RIb54b710_41,RIb54b698_40,RIb54bb48_50,RIb54bad0_49,RIb54b788_42,RIb54b620_39,
        RIb54b878_44,RIb54b800_43,RIb54b3c8_34,RIb54b4b8_36,RIb54b440_35,RIb54ba58_48,RIb54b9e0_47,RIb54b5a8_38,RIb54b530_37,RIb54bf08_58,
        RIb54be90_57,RIb54c160_63,RIb54bda0_55,RIb54bd28_54,RIb54bc38_52,RIb54be18_56,RIb54bcb0_53,RIb54c340_67,RIb54c0e8_62,RIb54bbc0_51,
        RIb54c250_65,RIb54c1d8_64,RIb54c070_61,RIb54bff8_60,RIb54c2c8_66,RIb54bf80_59,RIb54c8e0_79,RIb54c700_75,RIb54c778_76,RIb54c610_73,
        RIb54c520_71,RIb54c430_69,RIb54c598_72,RIb54c4a8_70,RIb54c868_78,RIb54c7f0_77,RIb54c3b8_68,RIb54cb38_84,RIb54cac0_83,RIb54ca48_82,
        RIb54c9d0_81,RIb54c958_80,RIb54c688_74,RIb54cca0_87,RIb54cc28_86,RIb54cef8_92,RIb54ce80_91,RIb54cd90_89,RIb54cfe8_94,RIb54d240_99,
        RIb54ce08_90,RIb54d330_101,RIb54d2b8_100,RIb54cbb0_85,RIb54d150_97,RIb54d1c8_98,RIb54d0d8_96,RIb54d060_95,RIb54cf70_93,RIb54cd18_88,
        RIb54d498_104,RIb54d420_103,RIb54d6f0_109,RIb54d678_108,RIb54db28_118,RIb54dab0_117,RIb54d768_110,RIb54d510_105,RIb54d858_112,RIb54d7e0_111,
        RIb54d3a8_102,RIb54da38_116,RIb54d9c0_115,RIb54d948_114,RIb54d8d0_113,RIb54d588_106,RIb54d600_107,RIb54dee8_126,RIb54de70_125,RIb54e050_129,
        RIb54dfd8_128,RIb54e140_131,RIb54e0c8_130,RIb54df60_127,RIb54dd08_122,RIb54e230_133,RIb54e1b8_132,RIb54dba0_119,RIb54dc90_121,RIb54dc18_120,
        RIb54e320_135,RIb54e2a8_134,RIb54dd80_123,RIb54ddf8_124,RIb54e500_139,RIb54e488_138,RIb54e6e0_143,RIb54e668_142,RIb54eb18_152,RIb54eaa0_151,
        RIb54e758_144,RIb54e7d0_145,RIb54e848_146,RIb54e410_137,RIb54e398_136,RIb54ea28_150,RIb54e9b0_149,RIb54e938_148,RIb54e8c0_147,RIb54e578_140,
        RIb54e5f0_141,RIb54eed8_160,RIb54ee60_159,RIb54f040_163,RIb54efc8_162,RIb54f220_167,RIb54f1a8_166,RIb54ef50_161,RIb54ede8_158,RIb54f130_165,
        RIb54f0b8_164,RIb54eb90_153,RIb54ec80_155,RIb54ec08_154,RIb54f310_169,RIb54f298_168,RIb54ed70_157,RIb54ecf8_156,RIb54f6d0_177,RIb54f658_176,
        RIb54f838_180,RIb54f7c0_179,RIb54f478_172,RIb54f400_171,RIb54fa18_184,RIb54f9a0_183,RIb54f928_182,RIb54f8b0_181,RIb54f388_170,RIb54f748_178,
        RIb54f5e0_175,RIb54fb08_186,RIb54fa90_185,RIb54f568_174,RIb54f4f0_173,RIb54ff40_195,RIb54fdd8_192,RIb54fc70_189,RIb54fbf8_188,RIb550300_203,
        RIb550288_202,RIb54fd60_191,RIb54fce8_190,RIb54fec8_194,RIb54fe50_193,RIb54fb80_187,RIb550120_199,RIb5500a8_198,RIb550030_197,RIb54ffb8_196,
        RIb550210_201,RIb550198_200,RIb550990_217,RIb550918_216,RIb550738_212,RIb5506c0_211,RIb550b70_221,RIb550af8_220,RIb5505d0_209,RIb550558_208,
        RIb5504e0_207,RIb550468_206,RIb5503f0_205,RIb550a80_219,RIb550a08_218,RIb5508a0_215,RIb550828_214,RIb5507b0_213,RIb550648_210,RIb550378_204,
        RIb550e40_227,RIb550eb8_228,RIb550f30_229,RIb550fa8_230,RIb550c60_223,RIb550cd8_224,RIb550d50_225,RIb550dc8_226,RIb5515c0_243,RIb551728_246,
        RIb551458_240,RIb5513e0_239,RIb5516b0_245,RIb551548_242,RIb5514d0_241,RIb550be8_222,RIb551200_235,RIb551368_238,RIb5512f0_237,RIb551188_234,
        RIb551110_233,RIb551638_244,RIb551020_231,RIb551278_236,RIb551098_232,RIb552448_274,RIb5526a0_279,RIb552628_278,RIb552010_265,RIb552268_270,
        RIb5525b0_277,RIb552538_276,RIb5521f0_269,RIb552178_268,RIb552718_280,RIb5524c0_275,RIb552358_272,RIb5522e0_271,RIb552100_267,RIb552088_266,
        RIb552790_281,RIb5523d0_273,RIb552c40_291,RIb552e98_296,RIb552e20_295,RIb552808_282,RIb552a60_287,RIb552da8_294,RIb552d30_293,RIb5529e8_286,
        RIb552970_285,RIb552f10_297,RIb552cb8_292,RIb552b50_289,RIb552ad8_288,RIb5528f8_284,RIb552880_283,RIb552f88_298,RIb552bc8_290,RIb553c30_325,
        RIb553e88_330,RIb553e10_329,RIb5537f8_316,RIb553a50_321,RIb553d98_328,RIb553d20_327,RIb5539d8_320,RIb553960_319,RIb553f00_331,RIb553ca8_326,
        RIb553b40_323,RIb553ac8_322,RIb5538e8_318,RIb553870_317,RIb553f78_332,RIb553bb8_324,RIb553618_312,RIb553780_315,RIb5534b0_309,RIb553438_308,
        RIb553708_314,RIb5535a0_311,RIb553528_310,RIb553000_299,RIb553258_304,RIb5533c0_307,RIb553348_306,RIb5531e0_303,RIb553168_302,RIb553690_313,
        RIb553078_300,RIb5532d0_305,RIb5530f0_301,RIb554068_334,RIb554680_347,RIb554608_346,RIb553ff0_333,RIb554248_338,RIb554590_345,RIb554518_344,
        RIb5541d0_337,RIb554158_336,RIb5542c0_339,RIb5540e0_335,RIb5543b0_341,RIb554338_340,RIb5544a0_343,RIb554428_342,RIb554770_349,RIb5546f8_348,
        RIb554ba8_358,RIb554d88_362,RIb554e00_363,RIb5549c8_354,RIb554950_353,RIb554d10_361,RIb554c98_360,RIb5547e8_350,RIb554ef0_365,RIb554e78_364,
        RIb554c20_359,RIb554ab8_356,RIb554a40_355,RIb5548d8_352,RIb554860_351,RIb554f68_366,RIb554b30_357,RIb555058_368,RIb555670_381,RIb5555f8_380,
        RIb554fe0_367,RIb555238_372,RIb555580_379,RIb555508_378,RIb5551c0_371,RIb555148_370,RIb5552b0_373,RIb5550d0_369,RIb5553a0_375,RIb555328_374,
        RIb555490_377,RIb555418_376,RIb555760_383,RIb5556e8_382,RIb5565e8_414,RIb556750_417,RIb556480_411,RIb556408_410,RIb5566d8_416,RIb556570_413,
        RIb5564f8_412,RIb555fd0_401,RIb556228_406,RIb556390_409,RIb556318_408,RIb5561b0_405,RIb556138_404,RIb556660_415,RIb556048_402,RIb5562a0_407,
        RIb5560c0_403,RIb555940_387,RIb555ee0_399,RIb555e68_398,RIb555aa8_390,RIb555a30_389,RIb5558c8_386,RIb555850_385,RIb5557d8_384,RIb555df0_397,
        RIb555b20_391,RIb5559b8_388,RIb555b98_392,RIb555c10_393,RIb555d00_395,RIb555c88_394,RIb555f58_400,RIb555d78_396,RIb557308_442,RIb557560_447,
        RIb5575d8_448,RIb5571a0_439,RIb557128_438,RIb5574e8_446,RIb557470_445,RIb556fc0_435,RIb557650_449,RIb557380_443,RIb5573f8_444,RIb557290_441,
        RIb557218_440,RIb5570b0_437,RIb557038_436,RIb557740_451,RIb5576c8_450,RIb556c00_427,RIb556ed0_433,RIb556e58_432,RIb5569a8_422,RIb556930_421,
        RIb5567c8_418,RIb556a20_423,RIb556d68_430,RIb556de0_431,RIb556cf0_429,RIb556c78_428,RIb556b10_425,RIb556a98_424,RIb5568b8_420,RIb556840_419,
        RIb556f48_434,RIb556b88_426,RIb557fb0_469,RIb5580a0_471,RIb5585c8_482,RIb558028_470,RIb558370_477,RIb5582f8_476,RIb558280_475,RIb558208_474,
        RIb558730_485,RIb558640_483,RIb558550_481,RIb558190_473,RIb558118_472,RIb558460_479,RIb5583e8_478,RIb5586b8_484,RIb5584d8_480,RIb557b00_459,
        RIb557830_453,RIb557ce0_463,RIb557bf0_461,RIb557b78_460,RIb557c68_462,RIb557a88_458,RIb557a10_457,RIb557f38_468,RIb557d58_464,RIb557dd0_465,
        RIb557998_456,RIb557920_455,RIb5577b8_452,RIb5578a8_454,RIb557ec0_467,RIb557e48_466,RIb559180_507,RIb5591f8_508,RIb558fa0_503,RIb559018_504,
        RIb559108_506,RIb559090_505,RIb559540_515,RIb5595b8_516,RIb559720_519,RIb5596a8_518,RIb559630_517,RIb559360_511,RIb5593d8_512,RIb5594c8_514,
        RIb559450_513,RIb5592e8_510,RIb559270_509,RIb558a00_491,RIb558988_490,RIb558910_489,RIb5587a8_486,RIb558cd0_497,RIb558c58_496,RIb558be0_495,
        RIb558898_488,RIb558820_487,RIb558d48_498,RIb558dc0_499,RIb558e38_500,RIb558a78_492,RIb558b68_494,RIb558af0_493,RIb558f28_502,RIb558eb0_501,
        RIb55a4b8_548,RIb55a440_547,RIb55a080_539,RIb55a008_538,RIb55a350_545,RIb55a3c8_546,RIb559f90_537,RIb55a2d8_544,RIb55a710_553,RIb55a698_552,
        RIb55a0f8_540,RIb55a170_541,RIb55a1e8_542,RIb55a530_549,RIb55a260_543,RIb55a620_551,RIb55a5a8_550,RIb559d38_532,RIb559db0_533,RIb559978_524,
        RIb5599f0_525,RIb559ae0_527,RIb559a68_526,RIb559cc0_531,RIb559c48_530,RIb559f18_536,RIb559b58_528,RIb559bd0_529,RIb559900_523,RIb559888_522,
        RIb559798_520,RIb559810_521,RIb559ea0_535,RIb559e28_534,RIb55ab48_562,RIb55aad0_561,RIb55a968_558,RIb55a8f0_557,RIb55aa58_560,RIb55a9e0_559,
        RIb55a878_556,RIb55a800_555,RIb55af08_570,RIb55ad28_566,RIb55ada0_567,RIb55a788_554,RIb55abc0_563,RIb55acb0_565,RIb55ac38_564,RIb55ae90_569,
        RIb55ae18_568,RIb55af80_571,RIb55aff8_572,RIb55b160_575,RIb55b1d8_576,RIb55b2c8_578,RIb55b250_577,RIb55b4a8_582,RIb55b430_581,RIb55b700_587,
        RIb55b340_579,RIb55b3b8_580,RIb55b520_583,RIb55b598_584,RIb55b0e8_574,RIb55b070_573,RIb55b688_586,RIb55b610_585,RIb55b778_588,RIb55bca0_599,
        RIb55bc28_598,RIb55bbb0_597,RIb55bb38_596,RIb55bac0_595,RIb55ba48_594,RIb55b9d0_593,RIb55b958_592,RIb55b8e0_591,RIb55b868_590,RIb55b7f0_589,
        RIb55c3a8_614,RIb55be80_603,RIb55bef8_604,RIb55be08_602,RIb55bd90_601,RIb55bd18_600,RIb55bf70_605,RIb55bfe8_606,RIb55c060_607,RIb55c0d8_608,
        RIb55c150_609,RIb55c1c8_610,RIb55c240_611,RIb55c2b8_612,RIb55c330_613,R_267_b942f48,R_268_b942ff0,R_269_b943098,R_26a_b943140,R_26b_b9431e8,
        R_26c_b943290,R_26d_b943338,R_26e_b9433e0,R_26f_b943488,R_270_b943530,R_271_b9435d8,R_272_b943680,R_273_b943728,R_274_b9437d0,R_275_b943878,
        R_276_b943920,R_277_b9439c8,R_278_b943a70,R_279_b943b18,R_27a_b943bc0,R_27b_b943c68,R_27c_b943d10,R_27d_b943db8,R_27e_b943e60,R_27f_b943f08,
        R_280_b943fb0,R_281_b944058,R_289_b944598,R_28a_b944640,R_28b_b9446e8,R_28c_b944790,R_28d_b944838,R_28e_b9448e0,R_28f_b944988,R_290_b944a30,
        R_291_b944ad8,R_292_b944b80,R_293_b944c28,R_294_b944cd0,R_295_b944d78,R_296_b944e20,R_297_b944ec8,R_298_b944f70,R_299_b945018,R_29a_b9450c0,
        R_29b_b945168,R_29c_b945210,R_29d_b9452b8,R_29e_b945360,R_29f_b945408,R_2a0_b9454b0,R_2a1_b945558,R_2a2_b945600,R_2a3_b9456a8);
input RIb54a900_11,RIb54a888_10,RIb54a810_9,RIb54a798_8,RIb54a720_7,RIb54a6a8_6,RIb54a630_5,RIb54a5b8_4,RIb54a540_3,
        RIb54a4c8_2,RIb54a450_1,RIb5517a0_247,RIb551980_251,RIb54ab58_16,RIb54abd0_17,RIb54aae0_15,RIb54aa68_14,RIb54a9f0_13,RIb551908_250,
        RIb551b60_255,RIb551ae8_254,RIb551f98_264,RIb551f20_263,RIb551cc8_258,RIb551c50_257,RIb551bd8_256,RIb551890_249,RIb551818_248,RIb551ea8_262,
        RIb551e30_261,RIb551db8_260,RIb551d40_259,RIb5519f8_252,RIb551a70_253,RIb54ad38_20,RIb54acc0_19,RIb54af18_24,RIb54aea0_23,RIb54b350_33,
        RIb54b2d8_32,RIb54af90_25,RIb54b008_26,RIb54b080_27,RIb54ac48_18,RIb54a978_12,RIb54b260_31,RIb54b1e8_30,RIb54b170_29,RIb54b0f8_28,
        RIb54adb0_21,RIb54ae28_22,RIb54b968_46,RIb54b8f0_45,RIb54b710_41,RIb54b698_40,RIb54bb48_50,RIb54bad0_49,RIb54b788_42,RIb54b620_39,
        RIb54b878_44,RIb54b800_43,RIb54b3c8_34,RIb54b4b8_36,RIb54b440_35,RIb54ba58_48,RIb54b9e0_47,RIb54b5a8_38,RIb54b530_37,RIb54bf08_58,
        RIb54be90_57,RIb54c160_63,RIb54bda0_55,RIb54bd28_54,RIb54bc38_52,RIb54be18_56,RIb54bcb0_53,RIb54c340_67,RIb54c0e8_62,RIb54bbc0_51,
        RIb54c250_65,RIb54c1d8_64,RIb54c070_61,RIb54bff8_60,RIb54c2c8_66,RIb54bf80_59,RIb54c8e0_79,RIb54c700_75,RIb54c778_76,RIb54c610_73,
        RIb54c520_71,RIb54c430_69,RIb54c598_72,RIb54c4a8_70,RIb54c868_78,RIb54c7f0_77,RIb54c3b8_68,RIb54cb38_84,RIb54cac0_83,RIb54ca48_82,
        RIb54c9d0_81,RIb54c958_80,RIb54c688_74,RIb54cca0_87,RIb54cc28_86,RIb54cef8_92,RIb54ce80_91,RIb54cd90_89,RIb54cfe8_94,RIb54d240_99,
        RIb54ce08_90,RIb54d330_101,RIb54d2b8_100,RIb54cbb0_85,RIb54d150_97,RIb54d1c8_98,RIb54d0d8_96,RIb54d060_95,RIb54cf70_93,RIb54cd18_88,
        RIb54d498_104,RIb54d420_103,RIb54d6f0_109,RIb54d678_108,RIb54db28_118,RIb54dab0_117,RIb54d768_110,RIb54d510_105,RIb54d858_112,RIb54d7e0_111,
        RIb54d3a8_102,RIb54da38_116,RIb54d9c0_115,RIb54d948_114,RIb54d8d0_113,RIb54d588_106,RIb54d600_107,RIb54dee8_126,RIb54de70_125,RIb54e050_129,
        RIb54dfd8_128,RIb54e140_131,RIb54e0c8_130,RIb54df60_127,RIb54dd08_122,RIb54e230_133,RIb54e1b8_132,RIb54dba0_119,RIb54dc90_121,RIb54dc18_120,
        RIb54e320_135,RIb54e2a8_134,RIb54dd80_123,RIb54ddf8_124,RIb54e500_139,RIb54e488_138,RIb54e6e0_143,RIb54e668_142,RIb54eb18_152,RIb54eaa0_151,
        RIb54e758_144,RIb54e7d0_145,RIb54e848_146,RIb54e410_137,RIb54e398_136,RIb54ea28_150,RIb54e9b0_149,RIb54e938_148,RIb54e8c0_147,RIb54e578_140,
        RIb54e5f0_141,RIb54eed8_160,RIb54ee60_159,RIb54f040_163,RIb54efc8_162,RIb54f220_167,RIb54f1a8_166,RIb54ef50_161,RIb54ede8_158,RIb54f130_165,
        RIb54f0b8_164,RIb54eb90_153,RIb54ec80_155,RIb54ec08_154,RIb54f310_169,RIb54f298_168,RIb54ed70_157,RIb54ecf8_156,RIb54f6d0_177,RIb54f658_176,
        RIb54f838_180,RIb54f7c0_179,RIb54f478_172,RIb54f400_171,RIb54fa18_184,RIb54f9a0_183,RIb54f928_182,RIb54f8b0_181,RIb54f388_170,RIb54f748_178,
        RIb54f5e0_175,RIb54fb08_186,RIb54fa90_185,RIb54f568_174,RIb54f4f0_173,RIb54ff40_195,RIb54fdd8_192,RIb54fc70_189,RIb54fbf8_188,RIb550300_203,
        RIb550288_202,RIb54fd60_191,RIb54fce8_190,RIb54fec8_194,RIb54fe50_193,RIb54fb80_187,RIb550120_199,RIb5500a8_198,RIb550030_197,RIb54ffb8_196,
        RIb550210_201,RIb550198_200,RIb550990_217,RIb550918_216,RIb550738_212,RIb5506c0_211,RIb550b70_221,RIb550af8_220,RIb5505d0_209,RIb550558_208,
        RIb5504e0_207,RIb550468_206,RIb5503f0_205,RIb550a80_219,RIb550a08_218,RIb5508a0_215,RIb550828_214,RIb5507b0_213,RIb550648_210,RIb550378_204,
        RIb550e40_227,RIb550eb8_228,RIb550f30_229,RIb550fa8_230,RIb550c60_223,RIb550cd8_224,RIb550d50_225,RIb550dc8_226,RIb5515c0_243,RIb551728_246,
        RIb551458_240,RIb5513e0_239,RIb5516b0_245,RIb551548_242,RIb5514d0_241,RIb550be8_222,RIb551200_235,RIb551368_238,RIb5512f0_237,RIb551188_234,
        RIb551110_233,RIb551638_244,RIb551020_231,RIb551278_236,RIb551098_232,RIb552448_274,RIb5526a0_279,RIb552628_278,RIb552010_265,RIb552268_270,
        RIb5525b0_277,RIb552538_276,RIb5521f0_269,RIb552178_268,RIb552718_280,RIb5524c0_275,RIb552358_272,RIb5522e0_271,RIb552100_267,RIb552088_266,
        RIb552790_281,RIb5523d0_273,RIb552c40_291,RIb552e98_296,RIb552e20_295,RIb552808_282,RIb552a60_287,RIb552da8_294,RIb552d30_293,RIb5529e8_286,
        RIb552970_285,RIb552f10_297,RIb552cb8_292,RIb552b50_289,RIb552ad8_288,RIb5528f8_284,RIb552880_283,RIb552f88_298,RIb552bc8_290,RIb553c30_325,
        RIb553e88_330,RIb553e10_329,RIb5537f8_316,RIb553a50_321,RIb553d98_328,RIb553d20_327,RIb5539d8_320,RIb553960_319,RIb553f00_331,RIb553ca8_326,
        RIb553b40_323,RIb553ac8_322,RIb5538e8_318,RIb553870_317,RIb553f78_332,RIb553bb8_324,RIb553618_312,RIb553780_315,RIb5534b0_309,RIb553438_308,
        RIb553708_314,RIb5535a0_311,RIb553528_310,RIb553000_299,RIb553258_304,RIb5533c0_307,RIb553348_306,RIb5531e0_303,RIb553168_302,RIb553690_313,
        RIb553078_300,RIb5532d0_305,RIb5530f0_301,RIb554068_334,RIb554680_347,RIb554608_346,RIb553ff0_333,RIb554248_338,RIb554590_345,RIb554518_344,
        RIb5541d0_337,RIb554158_336,RIb5542c0_339,RIb5540e0_335,RIb5543b0_341,RIb554338_340,RIb5544a0_343,RIb554428_342,RIb554770_349,RIb5546f8_348,
        RIb554ba8_358,RIb554d88_362,RIb554e00_363,RIb5549c8_354,RIb554950_353,RIb554d10_361,RIb554c98_360,RIb5547e8_350,RIb554ef0_365,RIb554e78_364,
        RIb554c20_359,RIb554ab8_356,RIb554a40_355,RIb5548d8_352,RIb554860_351,RIb554f68_366,RIb554b30_357,RIb555058_368,RIb555670_381,RIb5555f8_380,
        RIb554fe0_367,RIb555238_372,RIb555580_379,RIb555508_378,RIb5551c0_371,RIb555148_370,RIb5552b0_373,RIb5550d0_369,RIb5553a0_375,RIb555328_374,
        RIb555490_377,RIb555418_376,RIb555760_383,RIb5556e8_382,RIb5565e8_414,RIb556750_417,RIb556480_411,RIb556408_410,RIb5566d8_416,RIb556570_413,
        RIb5564f8_412,RIb555fd0_401,RIb556228_406,RIb556390_409,RIb556318_408,RIb5561b0_405,RIb556138_404,RIb556660_415,RIb556048_402,RIb5562a0_407,
        RIb5560c0_403,RIb555940_387,RIb555ee0_399,RIb555e68_398,RIb555aa8_390,RIb555a30_389,RIb5558c8_386,RIb555850_385,RIb5557d8_384,RIb555df0_397,
        RIb555b20_391,RIb5559b8_388,RIb555b98_392,RIb555c10_393,RIb555d00_395,RIb555c88_394,RIb555f58_400,RIb555d78_396,RIb557308_442,RIb557560_447,
        RIb5575d8_448,RIb5571a0_439,RIb557128_438,RIb5574e8_446,RIb557470_445,RIb556fc0_435,RIb557650_449,RIb557380_443,RIb5573f8_444,RIb557290_441,
        RIb557218_440,RIb5570b0_437,RIb557038_436,RIb557740_451,RIb5576c8_450,RIb556c00_427,RIb556ed0_433,RIb556e58_432,RIb5569a8_422,RIb556930_421,
        RIb5567c8_418,RIb556a20_423,RIb556d68_430,RIb556de0_431,RIb556cf0_429,RIb556c78_428,RIb556b10_425,RIb556a98_424,RIb5568b8_420,RIb556840_419,
        RIb556f48_434,RIb556b88_426,RIb557fb0_469,RIb5580a0_471,RIb5585c8_482,RIb558028_470,RIb558370_477,RIb5582f8_476,RIb558280_475,RIb558208_474,
        RIb558730_485,RIb558640_483,RIb558550_481,RIb558190_473,RIb558118_472,RIb558460_479,RIb5583e8_478,RIb5586b8_484,RIb5584d8_480,RIb557b00_459,
        RIb557830_453,RIb557ce0_463,RIb557bf0_461,RIb557b78_460,RIb557c68_462,RIb557a88_458,RIb557a10_457,RIb557f38_468,RIb557d58_464,RIb557dd0_465,
        RIb557998_456,RIb557920_455,RIb5577b8_452,RIb5578a8_454,RIb557ec0_467,RIb557e48_466,RIb559180_507,RIb5591f8_508,RIb558fa0_503,RIb559018_504,
        RIb559108_506,RIb559090_505,RIb559540_515,RIb5595b8_516,RIb559720_519,RIb5596a8_518,RIb559630_517,RIb559360_511,RIb5593d8_512,RIb5594c8_514,
        RIb559450_513,RIb5592e8_510,RIb559270_509,RIb558a00_491,RIb558988_490,RIb558910_489,RIb5587a8_486,RIb558cd0_497,RIb558c58_496,RIb558be0_495,
        RIb558898_488,RIb558820_487,RIb558d48_498,RIb558dc0_499,RIb558e38_500,RIb558a78_492,RIb558b68_494,RIb558af0_493,RIb558f28_502,RIb558eb0_501,
        RIb55a4b8_548,RIb55a440_547,RIb55a080_539,RIb55a008_538,RIb55a350_545,RIb55a3c8_546,RIb559f90_537,RIb55a2d8_544,RIb55a710_553,RIb55a698_552,
        RIb55a0f8_540,RIb55a170_541,RIb55a1e8_542,RIb55a530_549,RIb55a260_543,RIb55a620_551,RIb55a5a8_550,RIb559d38_532,RIb559db0_533,RIb559978_524,
        RIb5599f0_525,RIb559ae0_527,RIb559a68_526,RIb559cc0_531,RIb559c48_530,RIb559f18_536,RIb559b58_528,RIb559bd0_529,RIb559900_523,RIb559888_522,
        RIb559798_520,RIb559810_521,RIb559ea0_535,RIb559e28_534,RIb55ab48_562,RIb55aad0_561,RIb55a968_558,RIb55a8f0_557,RIb55aa58_560,RIb55a9e0_559,
        RIb55a878_556,RIb55a800_555,RIb55af08_570,RIb55ad28_566,RIb55ada0_567,RIb55a788_554,RIb55abc0_563,RIb55acb0_565,RIb55ac38_564,RIb55ae90_569,
        RIb55ae18_568,RIb55af80_571,RIb55aff8_572,RIb55b160_575,RIb55b1d8_576,RIb55b2c8_578,RIb55b250_577,RIb55b4a8_582,RIb55b430_581,RIb55b700_587,
        RIb55b340_579,RIb55b3b8_580,RIb55b520_583,RIb55b598_584,RIb55b0e8_574,RIb55b070_573,RIb55b688_586,RIb55b610_585,RIb55b778_588,RIb55bca0_599,
        RIb55bc28_598,RIb55bbb0_597,RIb55bb38_596,RIb55bac0_595,RIb55ba48_594,RIb55b9d0_593,RIb55b958_592,RIb55b8e0_591,RIb55b868_590,RIb55b7f0_589,
        RIb55c3a8_614,RIb55be80_603,RIb55bef8_604,RIb55be08_602,RIb55bd90_601,RIb55bd18_600,RIb55bf70_605,RIb55bfe8_606,RIb55c060_607,RIb55c0d8_608,
        RIb55c150_609,RIb55c1c8_610,RIb55c240_611,RIb55c2b8_612,RIb55c330_613;
output R_267_b942f48,R_268_b942ff0,R_269_b943098,R_26a_b943140,R_26b_b9431e8,R_26c_b943290,R_26d_b943338,R_26e_b9433e0,R_26f_b943488,
        R_270_b943530,R_271_b9435d8,R_272_b943680,R_273_b943728,R_274_b9437d0,R_275_b943878,R_276_b943920,R_277_b9439c8,R_278_b943a70,R_279_b943b18,
        R_27a_b943bc0,R_27b_b943c68,R_27c_b943d10,R_27d_b943db8,R_27e_b943e60,R_27f_b943f08,R_280_b943fb0,R_281_b944058,R_289_b944598,R_28a_b944640,
        R_28b_b9446e8,R_28c_b944790,R_28d_b944838,R_28e_b9448e0,R_28f_b944988,R_290_b944a30,R_291_b944ad8,R_292_b944b80,R_293_b944c28,R_294_b944cd0,
        R_295_b944d78,R_296_b944e20,R_297_b944ec8,R_298_b944f70,R_299_b945018,R_29a_b9450c0,R_29b_b945168,R_29c_b945210,R_29d_b9452b8,R_29e_b945360,
        R_29f_b945408,R_2a0_b9454b0,R_2a1_b945558,R_2a2_b945600,R_2a3_b9456a8;


wire \649_ZERO , \650_ONE , \651 , \652 , \653 , \654 , \655 , \656 , \657 ,
         \658 , \659 , \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 ,
         \668 , \669 , \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677 ,
         \678 , \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 ,
         \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 ,
         \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 ,
         \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 ,
         \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 ,
         \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 ,
         \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 ,
         \748 , \749 , \750 , \751 , \752_nG11dc , \753 , \754 , \755 , \756 , \757 ,
         \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 ,
         \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 ,
         \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 ,
         \788_nGff1 , \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 ,
         \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 ,
         \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 ,
         \818 , \819 , \820 , \821 , \822 , \823 , \824_nGfef , \825 , \826 , \827 ,
         \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 ,
         \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 ,
         \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 ,
         \858 , \859 , \860_nGe41 , \861 , \862 , \863 , \864 , \865 , \866 , \867 ,
         \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 ,
         \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 ,
         \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 ,
         \898_nGe3f , \899 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 ,
         \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 ,
         \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 ,
         \928 , \929 , \930 , \931 , \932 , \933 , \934_nGcc4 , \935 , \936 , \937 ,
         \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 ,
         \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 ,
         \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 ,
         \968 , \969 , \970 , \971 , \972_nGcc2 , \973 , \974 , \975 , \976 , \977 ,
         \978 , \979 , \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 ,
         \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 ,
         \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 ,
         \1008_nGb97 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 ,
         \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 ,
         \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 ,
         \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044_nGb95 , \1045 , \1046 , \1047 ,
         \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 ,
         \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 ,
         \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076_nGac0 , \1077 ,
         \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 ,
         \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 ,
         \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 ,
         \1108_nGac2 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 ,
         \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 ,
         \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 ,
         \1138 , \1139_nG95e , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 ,
         \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 ,
         \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 ,
         \1168 , \1169 , \1170 , \1171 , \1172_nG95c , \1173 , \1174 , \1175 , \1176 , \1177 ,
         \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 ,
         \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 ,
         \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 ,
         \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 ,
         \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 ,
         \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 ,
         \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244_nG1807 , \1245 , \1246 , \1247 ,
         \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 ,
         \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 ,
         \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 ,
         \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 ,
         \1288 , \1289 , \1290_nG191a , \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 ,
         \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 ,
         \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 ,
         \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 ,
         \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 ,
         \1338_nG1711 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 ,
         \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 ,
         \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 ,
         \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 ,
         \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 ,
         \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 ,
         \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 ,
         \1408 , \1409 , \1410 , \1411_nG15f9 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 ,
         \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 ,
         \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 ,
         \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 ,
         \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 ,
         \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 ,
         \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 ,
         \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 ,
         \1488 , \1489 , \1490 , \1491 , \1492 , \1493_nG14ed , \1494 , \1495 , \1496 , \1497 ,
         \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 ,
         \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 ,
         \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 ,
         \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 ,
         \1538_nG13f2 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 ,
         \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 ,
         \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 ,
         \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 ,
         \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 ,
         \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 ,
         \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 ,
         \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 ,
         \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 ,
         \1628_nG1300 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 ,
         \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 ,
         \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 ,
         \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 ,
         \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 ,
         \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 ,
         \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 ,
         \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707_nG11f7 ,
         \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 ,
         \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 ,
         \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 ,
         \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 ,
         \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 ,
         \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 ,
         \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 ,
         \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 ,
         \1788 , \1789_nG1116 , \1790 , \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 ,
         \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 ,
         \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 ,
         \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 ,
         \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 ,
         \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 ,
         \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 ,
         \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 ,
         \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 ,
         \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 ,
         \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 ,
         \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 ,
         \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 ,
         \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 ,
         \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 ,
         \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 ,
         \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 ,
         \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 ,
         \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 ,
         \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 ,
         \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 ,
         \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 ,
         \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 ,
         \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 , \2025_nG100c , \2026 , \2027 ,
         \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 ,
         \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 ,
         \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 ,
         \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 ,
         \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 ,
         \2078 , \2079 , \2080 , \2081_nGf30 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 ,
         \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 ,
         \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 ,
         \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 ,
         \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 ,
         \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 ,
         \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 ,
         \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 ,
         \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 ,
         \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 ,
         \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 ,
         \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 ,
         \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 ,
         \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 ,
         \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 ,
         \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 ,
         \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 ,
         \2248 , \2249 , \2250 , \2251 , \2252_nGe5c , \2253 , \2254 , \2255 , \2256 , \2257 ,
         \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 ,
         \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 ,
         \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 ,
         \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 ,
         \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 ,
         \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 ,
         \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 ,
         \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 ,
         \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 ,
         \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 ,
         \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365_nGda9 , \2366 , \2367 ,
         \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 ,
         \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 ,
         \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 ,
         \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407_nGcdf ,
         \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 ,
         \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 ,
         \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 ,
         \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 ,
         \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 ,
         \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 ,
         \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 ,
         \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 ,
         \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 ,
         \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 ,
         \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 ,
         \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 ,
         \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 ,
         \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 ,
         \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 ,
         \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 ,
         \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 ,
         \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 ,
         \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 ,
         \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 ,
         \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 ,
         \2618 , \2619 , \2620 , \2621_nGc52 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 ,
         \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 ,
         \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 ,
         \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 ,
         \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 ,
         \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 ,
         \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 ,
         \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 ,
         \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 ,
         \2708_nGbb2 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 ,
         \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 ,
         \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 ,
         \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 ,
         \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 ,
         \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 ,
         \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 ,
         \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 ,
         \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 ,
         \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 ,
         \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 ,
         \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 ,
         \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 ,
         \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 ,
         \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 , \2856_nGb3b , \2857 ,
         \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 ,
         \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 ,
         \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 ,
         \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 ,
         \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 ,
         \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 ,
         \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 ,
         \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 ,
         \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 ,
         \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 ,
         \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 ,
         \2968 , \2969_nGabe , \2970 , \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 ,
         \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 ,
         \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 ,
         \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 ,
         \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 ,
         \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 ,
         \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 ,
         \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 ,
         \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 ,
         \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 ,
         \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 ,
         \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 ,
         \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 ,
         \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 ,
         \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 ,
         \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124_nGa6e , \3125 , \3126 , \3127 ,
         \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 ,
         \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 ,
         \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 ,
         \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 ,
         \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 ,
         \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 ,
         \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 ,
         \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 , \3206_nG959 , \3207 ,
         \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 ,
         \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 ,
         \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 ,
         \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 ,
         \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 ,
         \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 ,
         \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 ,
         \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 ,
         \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 ,
         \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 ,
         \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 ,
         \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 ,
         \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 ,
         \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 ,
         \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 ,
         \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 ,
         \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 ,
         \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 ,
         \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 ,
         \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 ,
         \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 ,
         \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 ,
         \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 ,
         \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 ,
         \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 ,
         \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 ,
         \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 ,
         \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 ,
         \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 ,
         \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 ,
         \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 ,
         \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 ,
         \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 ,
         \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 ,
         \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 ,
         \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 ,
         \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 ,
         \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 ,
         \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 ,
         \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 ,
         \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 ,
         \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 ,
         \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 ,
         \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 ,
         \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 ,
         \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 ,
         \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 ,
         \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 ,
         \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 ,
         \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 ,
         \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 ,
         \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 ,
         \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 ,
         \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 ,
         \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 ,
         \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 ,
         \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 ,
         \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 ,
         \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 ,
         \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 ,
         \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 ,
         \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 ,
         \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 ,
         \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 ,
         \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 ,
         \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 ,
         \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 ,
         \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 ,
         \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 ,
         \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 ,
         \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 ,
         \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 ,
         \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 ,
         \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 ,
         \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 ,
         \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 ,
         \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 ,
         \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 ,
         \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 ,
         \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 ,
         \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 ,
         \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 ,
         \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 ,
         \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 ,
         \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 ,
         \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 ,
         \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 ,
         \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 ,
         \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 ,
         \4098 , \4099 , \4100 , \4101_nG11f9 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 ,
         \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 ,
         \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 ,
         \4128 , \4129 , \4130_nG1010 , \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 ,
         \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 ,
         \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 ,
         \4158 , \4159_nG100e , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 ,
         \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 ,
         \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187_nGe60 ,
         \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 ,
         \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 ,
         \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 , \4216_nGe5e , \4217 ,
         \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 ,
         \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 ,
         \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245_nGce3 , \4246 , \4247 ,
         \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 ,
         \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 ,
         \4268 , \4269 , \4270 , \4271 , \4272 , \4273_nGce1 , \4274 , \4275 , \4276 , \4277 ,
         \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 ,
         \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 ,
         \4298 , \4299 , \4300 , \4301 , \4302_nGbb6 , \4303 , \4304 , \4305 , \4306 , \4307 ,
         \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 ,
         \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 ,
         \4328 , \4329 , \4330 , \4331_nGbb4 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 ,
         \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 ,
         \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 ,
         \4358 , \4359 , \4360_nGade , \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 ,
         \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 ,
         \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 ,
         \4388 , \4389_nGae0 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 ,
         \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 ,
         \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 ,
         \4418_nG97f , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 ,
         \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 ,
         \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 , \4445 , \4446_nG97d , \4447 ,
         \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 ,
         \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 ,
         \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 ,
         \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 ,
         \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 ,
         \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 ,
         \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514_nG1821 , \4515 , \4516 , \4517 ,
         \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 ,
         \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 ,
         \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 ,
         \4548 , \4549 , \4550 , \4551 , \4552_nG1933 , \4553 , \4554 , \4555 , \4556 , \4557 ,
         \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 ,
         \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 ,
         \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 ,
         \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 ,
         \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 , \4605 , \4606_nG172a , \4607 ,
         \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 ,
         \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 ,
         \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 ,
         \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 ,
         \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 ,
         \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 ,
         \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 ,
         \4678 , \4679 , \4680 , \4681 , \4682 , \4683_nG1613 , \4684 , \4685 , \4686 , \4687 ,
         \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 ,
         \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 ,
         \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 ,
         \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 ,
         \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 ,
         \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 ,
         \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 ,
         \4758 , \4759 , \4760 , \4761 , \4762_nG1506 , \4763 , \4764 , \4765 , \4766 , \4767 ,
         \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 ,
         \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 ,
         \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 ,
         \4798 , \4799 , \4800_nG140b , \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 ,
         \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 ,
         \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 ,
         \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 ,
         \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 ,
         \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 ,
         \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 ,
         \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 , \4875 , \4876_nG1212 , \4877 ,
         \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 ,
         \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 ,
         \4898 , \4899 , \4900 , \4901 , \4902 , \4903_nG1319 , \4904 , \4905 , \4906 , \4907 ,
         \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 ,
         \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 ,
         \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 ,
         \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 ,
         \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 ,
         \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 ,
         \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 ,
         \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 ,
         \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 ,
         \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 ,
         \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 ,
         \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 ,
         \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 ,
         \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 ,
         \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 ,
         \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 , \5065_nG112f , \5066 , \5067 ,
         \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 ,
         \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 ,
         \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 ,
         \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 ,
         \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 ,
         \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 ,
         \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 ,
         \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 ,
         \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 ,
         \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 ,
         \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 ,
         \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 ,
         \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 ,
         \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 ,
         \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 ,
         \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 ,
         \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 ,
         \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 ,
         \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 ,
         \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 ,
         \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 ,
         \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 ,
         \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 ,
         \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 ,
         \5308 , \5309 , \5310 , \5311_nG1029 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 ,
         \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 ,
         \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 ,
         \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 ,
         \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 ,
         \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 ,
         \5368 , \5369 , \5370 , \5371_nGf4a , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 ,
         \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 ,
         \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 ,
         \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 ,
         \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 ,
         \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 ,
         \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 ,
         \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 ,
         \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 ,
         \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 ,
         \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 ,
         \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 ,
         \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 ,
         \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 ,
         \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 ,
         \5518 , \5519 , \5520_nGe7a , \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 ,
         \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 ,
         \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547_nGdc3 ,
         \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 ,
         \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 ,
         \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 ,
         \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 ,
         \5588_nGcfd , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 ,
         \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 ,
         \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 ,
         \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 ,
         \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 ,
         \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 ,
         \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 ,
         \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 ,
         \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 ,
         \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 ,
         \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 ,
         \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 ,
         \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 ,
         \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 ,
         \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 ,
         \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 ,
         \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 ,
         \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 ,
         \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 ,
         \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 ,
         \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 ,
         \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 ,
         \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 ,
         \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 ,
         \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 ,
         \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 ,
         \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 ,
         \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 ,
         \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 ,
         \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 ,
         \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 ,
         \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 ,
         \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 ,
         \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927_nGc6b ,
         \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 ,
         \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 ,
         \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 ,
         \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 ,
         \5968_nGbd0 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 ,
         \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 ,
         \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 ,
         \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 ,
         \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 ,
         \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 ,
         \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 ,
         \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 ,
         \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 ,
         \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 ,
         \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 ,
         \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 ,
         \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 ,
         \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 ,
         \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 ,
         \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 ,
         \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 ,
         \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 ,
         \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 ,
         \6158 , \6159 , \6160 , \6161 , \6162 , \6163_nGb55 , \6164 , \6165 , \6166 , \6167 ,
         \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 ,
         \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 ,
         \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 ,
         \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 ,
         \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 ,
         \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 ,
         \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 ,
         \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 ,
         \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 ,
         \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 ,
         \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 ,
         \6278 , \6279_nGadc , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 ,
         \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 ,
         \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 ,
         \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 ,
         \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 ,
         \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 ,
         \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 ,
         \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 ,
         \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 ,
         \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 ,
         \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 ,
         \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 ,
         \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 ,
         \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 ,
         \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 ,
         \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 ,
         \6438 , \6439 , \6440 , \6441 , \6442 , \6443_nGa88 , \6444 , \6445 , \6446 , \6447 ,
         \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 ,
         \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 ,
         \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 ,
         \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 ,
         \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 ,
         \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 ,
         \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 ,
         \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 ,
         \6528 , \6529 , \6530_nG97a , \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 ,
         \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 ,
         \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 ,
         \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 ,
         \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 ,
         \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 ,
         \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 ,
         \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 ,
         \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 ,
         \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 ,
         \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 ,
         \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 ,
         \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 ,
         \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 ,
         \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 ,
         \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 ,
         \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 ,
         \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 ,
         \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 ,
         \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 ,
         \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 ,
         \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 ,
         \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 ,
         \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 ,
         \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 ,
         \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 ,
         \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 ,
         \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 ,
         \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 ,
         \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 ,
         \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 ,
         \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 ,
         \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 ,
         \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 ,
         \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 ,
         \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 ,
         \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 ,
         \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 ,
         \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 ,
         \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 ,
         \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 ,
         \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 ,
         \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 ,
         \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 ,
         \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 ,
         \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 ,
         \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 ,
         \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 ,
         \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 ,
         \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 ,
         \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 ,
         \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 ,
         \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 ,
         \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 ,
         \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 ,
         \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 ,
         \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 ,
         \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 ,
         \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 ,
         \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 ,
         \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 ,
         \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 ,
         \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 ,
         \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 ,
         \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 ,
         \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 ,
         \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 ,
         \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 ,
         \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 ,
         \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 ,
         \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 ,
         \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 ,
         \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 ,
         \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 ,
         \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 ,
         \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 ,
         \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 ,
         \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 ,
         \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 ,
         \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 ,
         \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 ,
         \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 ,
         \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 ,
         \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 ,
         \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 ,
         \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 ,
         \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 ,
         \7398 , \7399 , \7400 , \7401 , \7402 , \7403_nG476 , \7404 , \7405 , \7406 , \7407_nG473 ,
         \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 ,
         \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 ,
         \7428_nG2fa , \7429 , \7430 , \7431 , \7432 , \7433_nG317 , \7434 , \7435_nG334 , \7436 , \7437 ,
         \7438 , \7439 , \7440 , \7441 , \7442_nG3a6 , \7443 , \7444 , \7445 , \7446 , \7447 ,
         \7448 , \7449 , \7450 , \7451 , \7452_nG3c3 , \7453 , \7454 , \7455_nG3e0 , \7456 , \7457 ,
         \7458 , \7459 , \7460 , \7461_nG41a , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 ,
         \7468_nG437 , \7469 , \7470 , \7471_nG453 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 ,
         \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 , \7485_nG3fd , \7486 , \7487 ,
         \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 ,
         \7498 , \7499 , \7500 , \7501 , \7502 , \7503_nG38a , \7504 , \7505 , \7506 , \7507 ,
         \7508 , \7509 , \7510 , \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 ,
         \7518_nG36d , \7519 , \7520 , \7521 , \7522_nG350 , \7523 , \7524 , \7525 , \7526 , \7527 ,
         \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 ,
         \7538 , \7539 , \7540 , \7541 , \7542_nG495 , \7543 , \7544_nG5cd , \7545 , \7546 , \7547 ,
         \7548_nG5cf , \7549 , \7550 , \7551 , \7552_nG5ee , \7553 , \7554 , \7555_nG5f0 , \7556 , \7557 ,
         \7558 , \7559 , \7560_nG5b0 , \7561 , \7562 , \7563_nG5ae , \7564 , \7565 , \7566 , \7567 ,
         \7568 , \7569_nG591 , \7570 , \7571 , \7572 , \7573 , \7574 , \7575_nG58f , \7576 , \7577 ,
         \7578 , \7579_nG570 , \7580 , \7581 , \7582 , \7583 , \7584 , \7585_nG572 , \7586 , \7587 ,
         \7588 , \7589_nG553 , \7590 , \7591 , \7592 , \7593 , \7594 , \7595_nG551 , \7596 , \7597 ,
         \7598 , \7599_nG534 , \7600 , \7601 , \7602_nG532 , \7603 , \7604 , \7605 , \7606 , \7607 ,
         \7608_nG513 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614_nG511 , \7615 , \7616 , \7617 ,
         \7618_nG4f4 , \7619 , \7620 , \7621_nG4f2 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627_nG4d3 ,
         \7628 , \7629 , \7630 , \7631 , \7632 , \7633_nG4d1 , \7634 , \7635 , \7636 , \7637_nG4b4 ,
         \7638 , \7639 , \7640_nG4b2 , \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 ,
         \7648 , \7649 , \7650 , \7651 , \7652_nG493 , \7653 , \7654 , \7655 , \7656 , \7657 ,
         \7658 , \7659_nG2231 , \7660 , \7661 , \7662 , \7663 , \7664 , \7665_nG21f6 , \7666 , \7667 ,
         \7668 , \7669 , \7670 , \7671 , \7672_nG21c6 , \7673 , \7674 , \7675 , \7676 , \7677 ,
         \7678 , \7679 , \7680 , \7681_nG2179 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 ,
         \7688 , \7689 , \7690 , \7691 , \7692_nG2115 , \7693 , \7694 , \7695 , \7696 , \7697 ,
         \7698_nG209c , \7699 , \7700 , \7701 , \7702 , \7703 , \7704_nG2013 , \7705 , \7706 , \7707 ,
         \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 , \7715_nG1f8e , \7716 , \7717 ,
         \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 , \7725 , \7726_nG1eef , \7727 ,
         \7728 , \7729 , \7730 , \7731 , \7732 , \7733 , \7734 , \7735 , \7736_nG1e25 , \7737 ,
         \7738 , \7739 , \7740 , \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747_nG1d58 ,
         \7748 , \7749 , \7750 , \7751 , \7752 , \7753_nG1c7b , \7754 , \7755 , \7756 , \7757 ,
         \7758 , \7759_nG1baa , \7760 , \7761 , \7762 , \7763 , \7764 , \7765_nG1ad8 , \7766 , \7767 ,
         \7768 , \7769 , \7770 , \7771_nG19f9 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777_nG18ff ,
         \7778 , \7779 , \7780 , \7781 , \7782 , \7783_nG17ec , \7784 , \7785 , \7786 , \7787 ,
         \7788 , \7789_nG16f6 , \7790 , \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797_nG15de ,
         \7798 , \7799 , \7800 , \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 ,
         \7808 , \7809 , \7810 , \7811 , \7812 , \7813_nG14d2 , \7814 , \7815 , \7816 , \7817 ,
         \7818 , \7819_nG13d7 , \7820 , \7821 , \7822 , \7823 , \7824 , \7825_nG12e5 , \7826 , \7827 ,
         \7828 , \7829 , \7830 , \7831_nG11da , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 ,
         \7838 , \7839 , \7840 , \7841_nG10fb , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 ,
         \7848 , \7849 , \7850 , \7851 , \7852_nGfed , \7853 , \7854 , \7855 , \7856 , \7857 ,
         \7858_nGf15 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864_nGe3d , \7865 , \7866 , \7867 ,
         \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 ,
         \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 ,
         \7888 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 ,
         \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 ,
         \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 ,
         \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 ,
         \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 ,
         \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 ,
         \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 ,
         \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964_nG2ace , \7965 , \7966 , \7967 ,
         \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 ,
         \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 ,
         \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 ,
         \7998 , \7999 , \8000_nG28f2 , \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 ,
         \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 ,
         \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 ,
         \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 ,
         \8038_nG28f0 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 ,
         \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 ,
         \8058 , \8059 , \8060 , \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 ,
         \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 , \8075 , \8076_nG273d , \8077 ,
         \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 ,
         \8088 , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 ,
         \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 ,
         \8108 , \8109 , \8110 , \8111 , \8112_nG273b , \8113 , \8114 , \8115 , \8116 , \8117 ,
         \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 ,
         \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 ,
         \8138 , \8139 , \8140 , \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 ,
         \8148 , \8149 , \8150_nG25c7 , \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 ,
         \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 ,
         \8168 , \8169 , \8170 , \8171 , \8172 , \8173 , \8174 , \8175 , \8176 , \8177 ,
         \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 ,
         \8188_nG25c5 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 ,
         \8198 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 ,
         \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 ,
         \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 , \8225 , \8226_nG2497 , \8227 ,
         \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 ,
         \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 ,
         \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 ,
         \8258 , \8259 , \8260 , \8261 , \8262_nG2495 , \8263 , \8264 , \8265 , \8266 , \8267 ,
         \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 ,
         \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 ,
         \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 ,
         \8298 , \8299 , \8300_nG23c0 , \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 ,
         \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 ,
         \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 ,
         \8328 , \8329 , \8330 , \8331 , \8332_nG23c2 , \8333 , \8334 , \8335 , \8336 , \8337 ,
         \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 ,
         \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 ,
         \8358 , \8359 , \8360 , \8361 , \8362 , \8363_nG2255 , \8364 , \8365 , \8366 , \8367 ,
         \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 ,
         \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 ,
         \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394_nG2253 , \8395 , \8396 , \8397 ,
         \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 ,
         \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 ,
         \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 ,
         \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 ,
         \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 ,
         \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 ,
         \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 ,
         \8468_nG310a , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 ,
         \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 ,
         \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 ,
         \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 ,
         \8508_nG3222 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 ,
         \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 ,
         \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 ,
         \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 ,
         \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 ,
         \8558 , \8559 , \8560 , \8561 , \8562 , \8563_nG3003 , \8564 , \8565 , \8566 , \8567 ,
         \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 ,
         \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 ,
         \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 ,
         \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 ,
         \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 ,
         \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 ,
         \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 ,
         \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 ,
         \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 ,
         \8658_nG2ee1 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 ,
         \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 ,
         \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 ,
         \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 ,
         \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 ,
         \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 ,
         \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 ,
         \8728 , \8729 , \8730_nG2df7 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 ,
         \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 ,
         \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 ,
         \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 ,
         \8768 , \8769 , \8770_nG2cf7 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 ,
         \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 ,
         \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 ,
         \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 ,
         \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 ,
         \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 ,
         \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 ,
         \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 ,
         \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857_nG2bf3 ,
         \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 ,
         \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 ,
         \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 ,
         \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 ,
         \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 ,
         \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 ,
         \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924_nG2ae9 , \8925 , \8926 , \8927 ,
         \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 ,
         \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 ,
         \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 ,
         \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 ,
         \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 ,
         \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 ,
         \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 ,
         \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 ,
         \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 ,
         \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 ,
         \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 , \9035_nG2a09 , \9036 , \9037 ,
         \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 ,
         \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 ,
         \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 ,
         \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 ,
         \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 ,
         \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 ,
         \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 ,
         \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 ,
         \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 , \9125 , \9126 , \9127 ,
         \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 ,
         \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 ,
         \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 ,
         \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 ,
         \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177 ,
         \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 ,
         \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 ,
         \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 ,
         \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 ,
         \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 ,
         \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 ,
         \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 ,
         \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 ,
         \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 ,
         \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 ,
         \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 ,
         \9288 , \9289_nG290d , \9290 , \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 ,
         \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 ,
         \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 ,
         \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 ,
         \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 ,
         \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 , \9345_nG282e , \9346 , \9347 ,
         \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 , \9355 , \9356 , \9357 ,
         \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 ,
         \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 ,
         \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 ,
         \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 ,
         \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 ,
         \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 ,
         \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 ,
         \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 ,
         \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 ,
         \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 ,
         \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 ,
         \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 , \9475 , \9476_nG2758 , \9477 ,
         \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 ,
         \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 ,
         \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 ,
         \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 ,
         \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 ,
         \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 ,
         \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 ,
         \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 ,
         \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 ,
         \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 ,
         \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 ,
         \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 ,
         \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 ,
         \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 ,
         \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 ,
         \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637_nG26ac ,
         \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 ,
         \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 ,
         \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 ,
         \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 ,
         \9678 , \9679_nG25e2 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 ,
         \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 ,
         \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 ,
         \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 ,
         \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 ,
         \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 ,
         \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 ,
         \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 ,
         \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 ,
         \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 ,
         \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 ,
         \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 ,
         \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 ,
         \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 ,
         \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 ,
         \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 ,
         \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 ,
         \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 ,
         \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 ,
         \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 ,
         \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886_nG2554 , \9887 ,
         \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 ,
         \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 ,
         \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 ,
         \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 ,
         \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 ,
         \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 ,
         \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 ,
         \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 ,
         \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974_nG24b2 , \9975 , \9976 , \9977 ,
         \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 ,
         \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 ,
         \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 ,
         \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 ,
         \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 ,
         \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 ,
         \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 ,
         \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 ,
         \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 ,
         \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 ,
         \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 ,
         \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 ,
         \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 ,
         \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 ,
         \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 ,
         \10128_nG2440 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 ,
         \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 ,
         \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 ,
         \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 ,
         \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 ,
         \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 ,
         \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 ,
         \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 ,
         \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 ,
         \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 ,
         \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 ,
         \10238_nG23be , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 ,
         \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 ,
         \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 ,
         \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 ,
         \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 ,
         \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 ,
         \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 ,
         \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 ,
         \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 ,
         \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 ,
         \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 ,
         \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 ,
         \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 ,
         \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 ,
         \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 ,
         \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 ,
         \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407_nG236e ,
         \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 ,
         \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 ,
         \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 ,
         \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 ,
         \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 ,
         \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 ,
         \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 ,
         \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 ,
         \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 ,
         \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504_nG2250 , \10505 , \10506 , \10507 ,
         \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 ,
         \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 ,
         \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 ,
         \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 ,
         \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 ,
         \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 ,
         \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 ,
         \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 ,
         \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 ,
         \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 ,
         \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 ,
         \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 ,
         \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 ,
         \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 ,
         \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 ,
         \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 ,
         \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 ,
         \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 ,
         \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 ,
         \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 ,
         \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 ,
         \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 ,
         \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 ,
         \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 ,
         \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 ,
         \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 ,
         \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 ,
         \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 ,
         \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 ,
         \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 ,
         \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 ,
         \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 ,
         \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 ,
         \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 ,
         \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 ,
         \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 ,
         \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 ,
         \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 ,
         \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 ,
         \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 ,
         \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 ,
         \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 ,
         \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 ,
         \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 ,
         \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 ,
         \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 ,
         \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 ,
         \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 ,
         \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 ,
         \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 ,
         \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 ,
         \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 ,
         \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 ,
         \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 ,
         \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 ,
         \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 ,
         \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 ,
         \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 ,
         \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 ,
         \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 ,
         \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 ,
         \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 ,
         \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 ,
         \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 ,
         \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 ,
         \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 ,
         \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 ,
         \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 ,
         \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 ,
         \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 ,
         \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 ,
         \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 ,
         \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 ,
         \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 ,
         \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 ,
         \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 ,
         \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 ,
         \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 ,
         \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 ,
         \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 ,
         \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 ,
         \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 ,
         \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 ,
         \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 ,
         \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 ,
         \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 ,
         \11368 , \11369 , \11370_nG2aeb , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 ,
         \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 ,
         \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 ,
         \11398 , \11399_nG2911 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 ,
         \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 ,
         \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 ,
         \11428_nG290f , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 ,
         \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 ,
         \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457_nG275c ,
         \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 ,
         \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 ,
         \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486_nG275a , \11487 ,
         \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 ,
         \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 ,
         \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515_nG25e6 , \11516 , \11517 ,
         \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 ,
         \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 ,
         \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544_nG25e4 , \11545 , \11546 , \11547 ,
         \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 ,
         \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 ,
         \11568 , \11569 , \11570 , \11571 , \11572 , \11573_nG24b6 , \11574 , \11575 , \11576 , \11577 ,
         \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 ,
         \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 ,
         \11598 , \11599 , \11600 , \11601 , \11602_nG24b4 , \11603 , \11604 , \11605 , \11606 , \11607 ,
         \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 ,
         \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 ,
         \11628 , \11629 , \11630 , \11631_nG23de , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 ,
         \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 ,
         \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 ,
         \11658 , \11659 , \11660_nG23e0 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 ,
         \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 ,
         \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 ,
         \11688 , \11689_nG2277 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 ,
         \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 ,
         \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 ,
         \11718_nG2275 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 ,
         \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 ,
         \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 ,
         \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 ,
         \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 ,
         \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 ,
         \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787_nG3124 ,
         \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 ,
         \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 ,
         \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 ,
         \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 ,
         \11828 , \11829 , \11830 , \11831 , \11832_nG323c , \11833 , \11834 , \11835 , \11836 , \11837 ,
         \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 ,
         \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 ,
         \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 ,
         \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 ,
         \11878 , \11879_nG301d , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 ,
         \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 ,
         \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 ,
         \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 ,
         \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 ,
         \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 ,
         \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 ,
         \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 ,
         \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 ,
         \11968 , \11969 , \11970 , \11971 , \11972_nG2efb , \11973 , \11974 , \11975 , \11976 , \11977 ,
         \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 ,
         \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 ,
         \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 ,
         \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 ,
         \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 ,
         \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 ,
         \12038_nG2e11 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 ,
         \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 ,
         \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 ,
         \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 ,
         \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 ,
         \12088 , \12089_nG2d11 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 ,
         \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 ,
         \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 ,
         \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 ,
         \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 ,
         \12138 , \12139 , \12140 , \12141 , \12142_nG2c0d , \12143 , \12144 , \12145 , \12146 , \12147 ,
         \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 ,
         \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 ,
         \12168 , \12169_nG2b05 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 ,
         \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 ,
         \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 ,
         \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 ,
         \12208 , \12209 , \12210_nG2a23 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 ,
         \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 ,
         \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 ,
         \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 ,
         \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 ,
         \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 ,
         \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 ,
         \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 ,
         \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 ,
         \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 ,
         \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 ,
         \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 ,
         \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 ,
         \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 ,
         \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 ,
         \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 ,
         \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 ,
         \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 ,
         \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 ,
         \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 ,
         \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 ,
         \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 ,
         \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 ,
         \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 ,
         \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 ,
         \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 ,
         \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 ,
         \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 ,
         \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 ,
         \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 ,
         \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 ,
         \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 ,
         \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 ,
         \12538 , \12539 , \12540 , \12541 , \12542 , \12543_nG292b , \12544 , \12545 , \12546 , \12547 ,
         \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 ,
         \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 ,
         \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 ,
         \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 ,
         \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 ,
         \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 ,
         \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 ,
         \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 ,
         \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 ,
         \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 ,
         \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 ,
         \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 ,
         \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 ,
         \12678 , \12679 , \12680 , \12681 , \12682_nG2848 , \12683 , \12684 , \12685 , \12686 , \12687 ,
         \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 ,
         \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 ,
         \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 ,
         \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 ,
         \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 ,
         \12738 , \12739 , \12740 , \12741_nG2776 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 ,
         \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 ,
         \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 ,
         \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 ,
         \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 ,
         \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 ,
         \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 ,
         \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 ,
         \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 ,
         \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 ,
         \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 ,
         \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 ,
         \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 ,
         \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 ,
         \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 ,
         \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 ,
         \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 ,
         \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 ,
         \12918_nG26c6 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 ,
         \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 ,
         \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 ,
         \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 ,
         \12958 , \12959_nG2600 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 ,
         \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 ,
         \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 ,
         \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 ,
         \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 ,
         \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 ,
         \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 ,
         \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 ,
         \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 ,
         \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 ,
         \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 ,
         \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 ,
         \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 ,
         \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 ,
         \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 ,
         \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 ,
         \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 ,
         \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 ,
         \13138 , \13139_nG256e , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 ,
         \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 ,
         \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 ,
         \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 ,
         \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 ,
         \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 ,
         \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 ,
         \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 ,
         \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 ,
         \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 ,
         \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 ,
         \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 ,
         \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 ,
         \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 ,
         \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 ,
         \13288 , \13289 , \13290 , \13291_nG24d0 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 ,
         \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 ,
         \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 ,
         \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 ,
         \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 ,
         \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 ,
         \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 ,
         \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 ,
         \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 ,
         \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 ,
         \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 ,
         \13398 , \13399 , \13400 , \13401 , \13402 , \13403_nG245a , \13404 , \13405 , \13406 , \13407 ,
         \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 ,
         \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 ,
         \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 ,
         \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 ,
         \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 ,
         \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 ,
         \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 ,
         \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 ,
         \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 ,
         \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 ,
         \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 ,
         \13518 , \13519 , \13520 , \13521 , \13522 , \13523_nG23dc , \13524 , \13525 , \13526 , \13527 ,
         \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 ,
         \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 ,
         \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 ,
         \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 ,
         \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 ,
         \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 ,
         \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 ,
         \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 ,
         \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 ,
         \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 ,
         \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 ,
         \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 ,
         \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 ,
         \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 ,
         \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 ,
         \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685_nG2388 , \13686 , \13687 ,
         \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 ,
         \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 ,
         \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 ,
         \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 ,
         \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 ,
         \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 ,
         \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 ,
         \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 ,
         \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775_nG2272 , \13776 , \13777 ,
         \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 ,
         \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 ,
         \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 ,
         \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 ,
         \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 ,
         \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 ,
         \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 ,
         \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 ,
         \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 ,
         \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 ,
         \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 ,
         \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 ,
         \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 ,
         \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 ,
         \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 ,
         \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 ,
         \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 ,
         \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 ,
         \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 ,
         \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 ,
         \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 ,
         \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 ,
         \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 ,
         \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 ,
         \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 ,
         \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 ,
         \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 ,
         \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 ,
         \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 ,
         \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 ,
         \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 ,
         \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 ,
         \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 ,
         \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 ,
         \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 ,
         \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 ,
         \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 ,
         \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 ,
         \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 ,
         \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 ,
         \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 ,
         \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 ,
         \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 ,
         \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 ,
         \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 ,
         \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 ,
         \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 ,
         \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 ,
         \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 ,
         \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 ,
         \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 ,
         \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 ,
         \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 ,
         \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 ,
         \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 ,
         \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 ,
         \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 ,
         \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 ,
         \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 ,
         \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 ,
         \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 ,
         \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 ,
         \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 ,
         \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 ,
         \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 ,
         \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 ,
         \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 ,
         \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 ,
         \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 ,
         \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 ,
         \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 ,
         \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 ,
         \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 ,
         \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 ,
         \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 ,
         \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 ,
         \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 ,
         \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 ,
         \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 ,
         \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 ,
         \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 ,
         \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 ,
         \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 ,
         \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 ,
         \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 ,
         \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 ,
         \14638_nG7bc , \14639 , \14640 , \14641 , \14642_nG7b9 , \14643 , \14644 , \14645_nG91b , \14646 , \14647 ,
         \14648 , \14649_nG91d , \14650 , \14651 , \14652 , \14653_nG93a , \14654 , \14655 , \14656_nG93c , \14657 ,
         \14658 , \14659 , \14660 , \14661_nG8fe , \14662 , \14663 , \14664 , \14665_nG8fc , \14666 , \14667 ,
         \14668 , \14669 , \14670_nG8df , \14671 , \14672 , \14673_nG8dd , \14674 , \14675 , \14676 , \14677 ,
         \14678 , \14679 , \14680_nG8bc , \14681 , \14682 , \14683 , \14684 , \14685 , \14686_nG8be , \14687 ,
         \14688 , \14689 , \14690_nG89f , \14691 , \14692 , \14693 , \14694 , \14695 , \14696_nG89d , \14697 ,
         \14698 , \14699 , \14700_nG87c , \14701 , \14702 , \14703 , \14704 , \14705 , \14706_nG87e , \14707 ,
         \14708 , \14709 , \14710_nG85d , \14711 , \14712 , \14713 , \14714 , \14715 , \14716_nG85b , \14717 ,
         \14718 , \14719 , \14720_nG83c , \14721 , \14722 , \14723_nG83a , \14724 , \14725 , \14726 , \14727 ,
         \14728 , \14729_nG81d , \14730 , \14731 , \14732 , \14733 , \14734 , \14735_nG81b , \14736 , \14737 ,
         \14738 , \14739_nG7fa , \14740 , \14741 , \14742 , \14743 , \14744 , \14745_nG7fc , \14746 , \14747 ,
         \14748 , \14749_nG7db , \14750 , \14751 , \14752 , \14753 , \14754 , \14755_nG7d9 , \14756 , \14757 ,
         \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 ,
         \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 ,
         \14778 , \14779_nG63b , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786_nG658 , \14787 ,
         \14788 , \14789 , \14790 , \14791 , \14792 , \14793_nG692 , \14794 , \14795 , \14796 , \14797 ,
         \14798 , \14799 , \14800 , \14801 , \14802 , \14803_nG6cc , \14804 , \14805_nG6e9 , \14806 , \14807 ,
         \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817_nG723 ,
         \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 ,
         \14828_nG740 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 ,
         \14838 , \14839_nG75d , \14840 , \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 ,
         \14848 , \14849 , \14850_nG77a , \14851 , \14852 , \14853 , \14854 , \14855 , \14856_nG797 , \14857 ,
         \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865_nG706 , \14866 , \14867 ,
         \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875_nG6af , \14876 , \14877 ,
         \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 ,
         \14888 , \14889 , \14890 , \14891 , \14892_nG675 , \14893 , \14894 , \14895 , \14896 , \14897 ,
         \14898 , \14899 , \14900 , \14901_nG3b42 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 ,
         \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 ,
         \14918 , \14919 , \14920_nG3b06 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 ,
         \14928 , \14929 , \14930 , \14931_nG3ac7 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 ,
         \14938_nG3a68 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 ,
         \14948 , \14949_nG39fa , \14950 , \14951 , \14952 , \14953 , \14954 , \14955_nG397d , \14956 , \14957 ,
         \14958 , \14959 , \14960 , \14961_nG38f4 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967_nG386b ,
         \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 ,
         \14978_nG37d3 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 , \14985_nG3717 , \14986 , \14987 ,
         \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995 , \14996_nG365e , \14997 ,
         \14998 , \14999 , \15000 , \15001 , \15002_nG358f , \15003 , \15004 , \15005 , \15006 , \15007 ,
         \15008_nG34be , \15009 , \15010 , \15011 , \15012 , \15013 , \15014_nG33ea , \15015 , \15016 , \15017 ,
         \15018 , \15019 , \15020_nG3309 , \15021 , \15022 , \15023 , \15024 , \15025 , \15026_nG3207 , \15027 ,
         \15028 , \15029 , \15030 , \15031 , \15032 , \15033_nG30ef , \15034 , \15035 , \15036 , \15037 ,
         \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 , \15045_nG2fe8 , \15046 , \15047 ,
         \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057_nG2ec6 ,
         \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 ,
         \15068 , \15069 , \15070 , \15071 , \15072 , \15073_nG2ddc , \15074 , \15075 , \15076 , \15077 ,
         \15078 , \15079_nG2cdc , \15080 , \15081 , \15082 , \15083 , \15084 , \15085_nG2bd8 , \15086 , \15087 ,
         \15088 , \15089 , \15090 , \15091_nG2acc , \15092 , \15093 , \15094 , \15095 , \15096 , \15097_nG29ee ,
         \15098 , \15099 , \15100 , \15101 , \15102 , \15103_nG28ee , \15104 , \15105 , \15106 , \15107 ,
         \15108 , \15109_nG2813 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115_nG2739 , \15116 ;
buf \U$labajz1583 ( R_267_b942f48, \7660 );
buf \U$labajz1584 ( R_268_b942ff0, \7666 );
buf \U$labajz1585 ( R_269_b943098, \7673 );
buf \U$labajz1586 ( R_26a_b943140, \7682 );
buf \U$labajz1587 ( R_26b_b9431e8, \7693 );
buf \U$labajz1588 ( R_26c_b943290, \7699 );
buf \U$labajz1589 ( R_26d_b943338, \7705 );
buf \U$labajz1590 ( R_26e_b9433e0, \7716 );
buf \U$labajz1591 ( R_26f_b943488, \7727 );
buf \U$labajz1592 ( R_270_b943530, \7737 );
buf \U$labajz1593 ( R_271_b9435d8, \7748 );
buf \U$labajz1594 ( R_272_b943680, \7754 );
buf \U$labajz1595 ( R_273_b943728, \7760 );
buf \U$labajz1596 ( R_274_b9437d0, \7766 );
buf \U$labajz1597 ( R_275_b943878, \7772 );
buf \U$labajz1598 ( R_276_b943920, \7778 );
buf \U$labajz1599 ( R_277_b9439c8, \7784 );
buf \U$labajz1600 ( R_278_b943a70, \7790 );
buf \U$labajz1601 ( R_279_b943b18, \7798 );
buf \U$labajz1602 ( R_27a_b943bc0, \7814 );
buf \U$labajz1603 ( R_27b_b943c68, \7820 );
buf \U$labajz1604 ( R_27c_b943d10, \7826 );
buf \U$labajz1605 ( R_27d_b943db8, \7832 );
buf \U$labajz1606 ( R_27e_b943e60, \7842 );
buf \U$labajz1607 ( R_27f_b943f08, \7853 );
buf \U$labajz1608 ( R_280_b943fb0, \7859 );
buf \U$labajz1609 ( R_281_b944058, \7865 );
buf \U$labajz1610 ( R_289_b944598, \14902 );
buf \U$labajz1611 ( R_28a_b944640, \14921 );
buf \U$labajz1612 ( R_28b_b9446e8, \14932 );
buf \U$labajz1613 ( R_28c_b944790, \14939 );
buf \U$labajz1614 ( R_28d_b944838, \14950 );
buf \U$labajz1615 ( R_28e_b9448e0, \14956 );
buf \U$labajz1616 ( R_28f_b944988, \14962 );
buf \U$labajz1617 ( R_290_b944a30, \14968 );
buf \U$labajz1618 ( R_291_b944ad8, \14979 );
buf \U$labajz1619 ( R_292_b944b80, \14986 );
buf \U$labajz1620 ( R_293_b944c28, \14997 );
buf \U$labajz1621 ( R_294_b944cd0, \15003 );
buf \U$labajz1622 ( R_295_b944d78, \15009 );
buf \U$labajz1623 ( R_296_b944e20, \15015 );
buf \U$labajz1624 ( R_297_b944ec8, \15021 );
buf \U$labajz1625 ( R_298_b944f70, \15027 );
buf \U$labajz1626 ( R_299_b945018, \15034 );
buf \U$labajz1627 ( R_29a_b9450c0, \15046 );
buf \U$labajz1628 ( R_29b_b945168, \15058 );
buf \U$labajz1629 ( R_29c_b945210, \15074 );
buf \U$labajz1630 ( R_29d_b9452b8, \15080 );
buf \U$labajz1631 ( R_29e_b945360, \15086 );
buf \U$labajz1632 ( R_29f_b945408, \15092 );
buf \U$labajz1633 ( R_2a0_b9454b0, \15098 );
buf \U$labajz1634 ( R_2a1_b945558, \15104 );
buf \U$labajz1635 ( R_2a2_b945600, \15110 );
buf \U$labajz1636 ( R_2a3_b9456a8, \15116 );
and \U$1 ( \651 , RIb54a888_10, RIb54a900_11);
nand \U$2 ( \652 , RIb54a810_9, \651 );
not \U$3 ( \653 , \652 );
nand \U$4 ( \654 , \653 , RIb54a798_8);
not \U$5 ( \655 , \654 );
nand \U$6 ( \656 , \655 , RIb54a720_7);
not \U$7 ( \657 , \656 );
nand \U$8 ( \658 , \657 , RIb54a6a8_6);
not \U$9 ( \659 , \658 );
nand \U$10 ( \660 , \659 , RIb54a630_5);
not \U$11 ( \661 , \660 );
nand \U$12 ( \662 , \661 , RIb54a5b8_4);
not \U$13 ( \663 , \662 );
nand \U$14 ( \664 , \663 , RIb54a540_3);
not \U$15 ( \665 , \664 );
nand \U$16 ( \666 , \665 , RIb54a4c8_2);
not \U$17 ( \667 , \666 );
nand \U$18 ( \668 , \667 , RIb54a450_1);
not \U$19 ( \669 , \668 );
not \U$20 ( \670 , RIb5517a0_247);
and \U$21 ( \671 , \669 , \670 );
and \U$22 ( \672 , \668 , RIb5517a0_247);
nor \U$23 ( \673 , \671 , \672 );
nor \U$24 ( \674 , RIb550dc8_226, RIb550e40_227);
not \U$25 ( \675 , \674 );
or \U$26 ( \676 , RIb550cd8_224, RIb550d50_225, RIb550eb8_228, RIb550f30_229);
nor \U$27 ( \677 , \675 , \676 , RIb550c60_223, RIb550fa8_230);
not \U$28 ( \678 , \677 );
nor \U$29 ( \679 , \678 , RIb54abd0_17);
nand \U$30 ( \680 , RIb54a9f0_13, \679 );
and \U$31 ( \681 , RIb54aa68_14, RIb54ab58_16);
nand \U$32 ( \682 , RIb54aae0_15, \681 );
nor \U$33 ( \683 , \680 , \682 );
and \U$34 ( \684 , RIb551890_249, \683 );
not \U$35 ( \685 , RIb54a9f0_13);
nand \U$36 ( \686 , \685 , \679 );
nor \U$37 ( \687 , \686 , RIb54aae0_15);
not \U$38 ( \688 , RIb54ab58_16);
nor \U$39 ( \689 , \688 , RIb54aa68_14);
and \U$40 ( \690 , \687 , \689 );
and \U$41 ( \691 , RIb551bd8_256, \690 );
not \U$42 ( \692 , RIb54aae0_15);
nor \U$43 ( \693 , \686 , \692 );
nor \U$44 ( \694 , RIb54aa68_14, RIb54ab58_16);
and \U$45 ( \695 , \693 , \694 );
and \U$46 ( \696 , \695 , RIb551db8_260);
nor \U$47 ( \697 , \680 , \692 );
and \U$48 ( \698 , \697 , \694 );
and \U$49 ( \699 , RIb551d40_259, \698 );
nor \U$50 ( \700 , \696 , \699 );
not \U$51 ( \701 , RIb54aa68_14);
nor \U$52 ( \702 , \701 , RIb54ab58_16);
and \U$53 ( \703 , \693 , \702 );
and \U$54 ( \704 , \703 , RIb551cc8_258);
and \U$55 ( \705 , \697 , \702 );
and \U$56 ( \706 , RIb551c50_257, \705 );
nor \U$57 ( \707 , \704 , \706 );
not \U$58 ( \708 , \686 );
and \U$59 ( \709 , \694 , \692 );
and \U$60 ( \710 , \708 , \709 );
and \U$61 ( \711 , \710 , RIb551f98_264);
not \U$62 ( \712 , \680 );
and \U$63 ( \713 , \712 , \709 );
and \U$64 ( \714 , RIb551f20_263, \713 );
nor \U$65 ( \715 , \711 , \714 );
and \U$66 ( \716 , \687 , \702 );
and \U$67 ( \717 , \716 , RIb551ea8_262);
nor \U$68 ( \718 , \680 , RIb54aae0_15);
and \U$69 ( \719 , \718 , \702 );
and \U$70 ( \720 , RIb551e30_261, \719 );
nor \U$71 ( \721 , \717 , \720 );
nand \U$72 ( \722 , \700 , \707 , \715 , \721 );
nor \U$73 ( \723 , \684 , \691 , \722 );
and \U$74 ( \724 , \687 , \681 );
and \U$75 ( \725 , \724 , RIb551ae8_254);
and \U$76 ( \726 , \718 , \689 );
and \U$77 ( \727 , RIb551b60_255, \726 );
nor \U$78 ( \728 , \725 , \727 );
not \U$79 ( \729 , RIb54a9f0_13);
nand \U$80 ( \730 , \729 , \709 );
not \U$81 ( \731 , \730 );
and \U$82 ( \732 , \731 , \677 , RIb54abd0_17);
nand \U$83 ( \733 , RIb551818_248, \732 );
and \U$84 ( \734 , \697 , \689 );
and \U$85 ( \735 , RIb551980_251, \734 );
nor \U$86 ( \736 , \686 , \682 );
and \U$87 ( \737 , RIb551908_250, \736 );
and \U$88 ( \738 , \693 , \689 );
and \U$89 ( \739 , \738 , RIb5519f8_252);
and \U$90 ( \740 , \718 , \681 );
and \U$91 ( \741 , RIb551a70_253, \740 );
nor \U$92 ( \742 , \739 , \741 );
not \U$93 ( \743 , \742 );
nor \U$94 ( \744 , \735 , \737 , \743 );
nand \U$95 ( \745 , \723 , \728 , \733 , \744 );
buf \U$96 ( \746 , \745 );
not \U$97 ( \747 , RIb54abd0_17);
not \U$98 ( \748 , \730 );
or \U$99 ( \749 , \747 , \748 );
nand \U$100 ( \750 , \749 , \677 );
buf \U$101 ( \751 , \750 );
_DC g11dc ( \752_nG11dc , \746 , \751 );
xor \U$102 ( \753 , \673 , \752_nG11dc );
not \U$103 ( \754 , \666 );
not \U$104 ( \755 , RIb54a450_1);
and \U$105 ( \756 , \754 , \755 );
and \U$106 ( \757 , \666 , RIb54a450_1);
nor \U$107 ( \758 , \756 , \757 );
and \U$108 ( \759 , RIb54b008_26, \705 );
and \U$109 ( \760 , RIb54b350_33, \710 );
and \U$110 ( \761 , \690 , RIb54af90_25);
and \U$111 ( \762 , RIb54ad38_20, \734 );
nor \U$112 ( \763 , \761 , \762 );
and \U$113 ( \764 , \724 , RIb54aea0_23);
and \U$114 ( \765 , RIb54af18_24, \726 );
nor \U$115 ( \766 , \764 , \765 );
and \U$116 ( \767 , \736 , RIb54acc0_19);
and \U$117 ( \768 , RIb54ac48_18, \683 );
nor \U$118 ( \769 , \767 , \768 );
and \U$119 ( \770 , \738 , RIb54adb0_21);
and \U$120 ( \771 , RIb54ae28_22, \740 );
nor \U$121 ( \772 , \770 , \771 );
nand \U$122 ( \773 , \763 , \766 , \769 , \772 );
nor \U$123 ( \774 , \759 , \760 , \773 );
and \U$124 ( \775 , \716 , RIb54b260_31);
and \U$125 ( \776 , RIb54b2d8_32, \713 );
nor \U$126 ( \777 , \775 , \776 );
nand \U$127 ( \778 , RIb54a978_12, \732 );
and \U$128 ( \779 , RIb54b170_29, \695 );
and \U$129 ( \780 , RIb54b1e8_30, \719 );
and \U$130 ( \781 , \703 , RIb54b080_27);
and \U$131 ( \782 , RIb54b0f8_28, \698 );
nor \U$132 ( \783 , \781 , \782 );
not \U$133 ( \784 , \783 );
nor \U$134 ( \785 , \779 , \780 , \784 );
nand \U$135 ( \786 , \774 , \777 , \778 , \785 );
buf \U$136 ( \787 , \786 );
_DC gff1 ( \788_nGff1 , \787 , \751 );
xor \U$137 ( \789 , \758 , \788_nGff1 );
not \U$138 ( \790 , \664 );
not \U$139 ( \791 , RIb54a4c8_2);
and \U$140 ( \792 , \790 , \791 );
and \U$141 ( \793 , \664 , RIb54a4c8_2);
nor \U$142 ( \794 , \792 , \793 );
and \U$143 ( \795 , RIb54b698_40, \724 );
and \U$144 ( \796 , RIb54bb48_50, \710 );
and \U$145 ( \797 , \703 , RIb54b878_44);
and \U$146 ( \798 , RIb54b8f0_45, \698 );
nor \U$147 ( \799 , \797 , \798 );
and \U$148 ( \800 , \719 , RIb54b9e0_47);
and \U$149 ( \801 , RIb54b620_39, \740 );
nor \U$150 ( \802 , \800 , \801 );
and \U$151 ( \803 , \734 , RIb54b530_37);
and \U$152 ( \804 , RIb54b4b8_36, \736 );
nor \U$153 ( \805 , \803 , \804 );
and \U$154 ( \806 , \738 , RIb54b5a8_38);
and \U$155 ( \807 , RIb54b440_35, \683 );
nor \U$156 ( \808 , \806 , \807 );
nand \U$157 ( \809 , \799 , \802 , \805 , \808 );
nor \U$158 ( \810 , \795 , \796 , \809 );
and \U$159 ( \811 , \716 , RIb54ba58_48);
and \U$160 ( \812 , RIb54bad0_49, \713 );
nor \U$161 ( \813 , \811 , \812 );
nand \U$162 ( \814 , RIb54b3c8_34, \732 );
and \U$163 ( \815 , RIb54b788_42, \690 );
and \U$164 ( \816 , RIb54b710_41, \726 );
and \U$165 ( \817 , \695 , RIb54b968_46);
and \U$166 ( \818 , RIb54b800_43, \705 );
nor \U$167 ( \819 , \817 , \818 );
not \U$168 ( \820 , \819 );
nor \U$169 ( \821 , \815 , \816 , \820 );
nand \U$170 ( \822 , \810 , \813 , \814 , \821 );
buf \U$171 ( \823 , \822 );
_DC gfef ( \824_nGfef , \823 , \751 );
xor \U$172 ( \825 , \794 , \824_nGfef );
and \U$173 ( \826 , \662 , RIb54a540_3);
not \U$174 ( \827 , \662 );
not \U$175 ( \828 , RIb54a540_3);
and \U$176 ( \829 , \827 , \828 );
nor \U$177 ( \830 , \826 , \829 );
and \U$178 ( \831 , \683 , RIb54bc38_52);
and \U$179 ( \832 , RIb54be90_57, \724 );
and \U$180 ( \833 , \740 , RIb54be18_56);
and \U$181 ( \834 , RIb54c0e8_62, \698 );
nor \U$182 ( \835 , \832 , \833 , \834 );
and \U$183 ( \836 , \703 , RIb54c070_61);
and \U$184 ( \837 , RIb54bff8_60, \705 );
nor \U$185 ( \838 , \836 , \837 );
and \U$186 ( \839 , \710 , RIb54c340_67);
and \U$187 ( \840 , RIb54c2c8_66, \713 );
nor \U$188 ( \841 , \839 , \840 );
and \U$189 ( \842 , \690 , RIb54bf80_59);
and \U$190 ( \843 , RIb54bf08_58, \726 );
nor \U$191 ( \844 , \842 , \843 );
nand \U$192 ( \845 , \835 , \838 , \841 , \844 );
nand \U$193 ( \846 , RIb54bbc0_51, \732 );
not \U$194 ( \847 , \846 );
nor \U$195 ( \848 , \831 , \845 , \847 );
and \U$196 ( \849 , \716 , RIb54c250_65);
and \U$197 ( \850 , RIb54c1d8_64, \719 );
nor \U$198 ( \851 , \849 , \850 );
and \U$199 ( \852 , \734 , RIb54bd28_54);
and \U$200 ( \853 , RIb54bcb0_53, \736 );
nor \U$201 ( \854 , \852 , \853 );
and \U$202 ( \855 , \695 , RIb54c160_63);
and \U$203 ( \856 , RIb54bda0_55, \738 );
nor \U$204 ( \857 , \855 , \856 );
nand \U$205 ( \858 , \848 , \851 , \854 , \857 );
buf \U$206 ( \859 , \858 );
_DC ge41 ( \860_nGe41 , \859 , \751 );
xor \U$207 ( \861 , \830 , \860_nGe41 );
not \U$208 ( \862 , \660 );
not \U$209 ( \863 , RIb54a5b8_4);
and \U$210 ( \864 , \862 , \863 );
and \U$211 ( \865 , \660 , RIb54a5b8_4);
nor \U$212 ( \866 , \864 , \865 );
and \U$213 ( \867 , \736 , RIb54c4a8_70);
and \U$214 ( \868 , \724 , RIb54c688_74);
and \U$215 ( \869 , RIb54c700_75, \726 );
nor \U$216 ( \870 , \868 , \869 );
and \U$217 ( \871 , \738 , RIb54c598_72);
and \U$218 ( \872 , RIb54c610_73, \740 );
nor \U$219 ( \873 , \871 , \872 );
and \U$220 ( \874 , \710 , RIb54cb38_84);
and \U$221 ( \875 , RIb54cac0_83, \713 );
nor \U$222 ( \876 , \874 , \875 );
and \U$223 ( \877 , \690 , RIb54c778_76);
and \U$224 ( \878 , RIb54c7f0_77, \705 );
nor \U$225 ( \879 , \877 , \878 );
nand \U$226 ( \880 , \870 , \873 , \876 , \879 );
not \U$227 ( \881 , RIb54c520_71);
not \U$228 ( \882 , \734 );
or \U$229 ( \883 , \881 , \882 );
nand \U$230 ( \884 , RIb54c3b8_68, \732 );
nand \U$231 ( \885 , \883 , \884 );
nor \U$232 ( \886 , \867 , \880 , \885 );
and \U$233 ( \887 , \695 , RIb54c958_80);
and \U$234 ( \888 , RIb54c9d0_81, \719 );
nor \U$235 ( \889 , \887 , \888 );
and \U$236 ( \890 , \703 , RIb54c868_78);
and \U$237 ( \891 , RIb54c8e0_79, \698 );
nor \U$238 ( \892 , \890 , \891 );
and \U$239 ( \893 , \716 , RIb54ca48_82);
and \U$240 ( \894 , RIb54c430_69, \683 );
nor \U$241 ( \895 , \893 , \894 );
nand \U$242 ( \896 , \886 , \889 , \892 , \895 );
buf \U$243 ( \897 , \896 );
_DC ge3f ( \898_nGe3f , \897 , \751 );
xor \U$244 ( \899 , \866 , \898_nGe3f );
and \U$245 ( \900 , \658 , RIb54a630_5);
not \U$246 ( \901 , \658 );
not \U$247 ( \902 , RIb54a630_5);
and \U$248 ( \903 , \901 , \902 );
nor \U$249 ( \904 , \900 , \903 );
and \U$250 ( \905 , \683 , RIb54cc28_86);
and \U$251 ( \906 , RIb54ce80_91, \724 );
and \U$252 ( \907 , \740 , RIb54ce08_90);
and \U$253 ( \908 , RIb54d0d8_96, \698 );
nor \U$254 ( \909 , \906 , \907 , \908 );
and \U$255 ( \910 , \703 , RIb54d060_95);
and \U$256 ( \911 , RIb54cfe8_94, \705 );
nor \U$257 ( \912 , \910 , \911 );
and \U$258 ( \913 , \710 , RIb54d330_101);
and \U$259 ( \914 , RIb54d2b8_100, \713 );
nor \U$260 ( \915 , \913 , \914 );
and \U$261 ( \916 , \690 , RIb54cf70_93);
and \U$262 ( \917 , RIb54cef8_92, \726 );
nor \U$263 ( \918 , \916 , \917 );
nand \U$264 ( \919 , \909 , \912 , \915 , \918 );
nand \U$265 ( \920 , RIb54cbb0_85, \732 );
not \U$266 ( \921 , \920 );
nor \U$267 ( \922 , \905 , \919 , \921 );
and \U$268 ( \923 , \716 , RIb54d240_99);
and \U$269 ( \924 , RIb54d1c8_98, \719 );
nor \U$270 ( \925 , \923 , \924 );
and \U$271 ( \926 , \734 , RIb54cd18_88);
and \U$272 ( \927 , RIb54cca0_87, \736 );
nor \U$273 ( \928 , \926 , \927 );
and \U$274 ( \929 , \695 , RIb54d150_97);
and \U$275 ( \930 , RIb54cd90_89, \738 );
nor \U$276 ( \931 , \929 , \930 );
nand \U$277 ( \932 , \922 , \925 , \928 , \931 );
buf \U$278 ( \933 , \932 );
_DC gcc4 ( \934_nGcc4 , \933 , \751 );
xor \U$279 ( \935 , \904 , \934_nGcc4 );
and \U$280 ( \936 , \656 , RIb54a6a8_6);
not \U$281 ( \937 , \656 );
not \U$282 ( \938 , RIb54a6a8_6);
and \U$283 ( \939 , \937 , \938 );
nor \U$284 ( \940 , \936 , \939 );
and \U$285 ( \941 , \736 , RIb54d498_104);
and \U$286 ( \942 , \716 , RIb54da38_116);
and \U$287 ( \943 , RIb54dab0_117, \713 );
nor \U$288 ( \944 , \942 , \943 );
and \U$289 ( \945 , \695 , RIb54d948_114);
nand \U$290 ( \946 , RIb54d3a8_102, \732 );
not \U$291 ( \947 , \946 );
nor \U$292 ( \948 , \945 , \947 );
and \U$293 ( \949 , \719 , RIb54d9c0_115);
and \U$294 ( \950 , RIb54d420_103, \683 );
nor \U$295 ( \951 , \949 , \950 );
and \U$296 ( \952 , \703 , RIb54d858_112);
and \U$297 ( \953 , RIb54d8d0_113, \698 );
nor \U$298 ( \954 , \952 , \953 );
nand \U$299 ( \955 , \944 , \948 , \951 , \954 );
and \U$300 ( \956 , \738 , RIb54d588_106);
and \U$301 ( \957 , RIb54d510_105, \734 );
nor \U$302 ( \958 , \956 , \957 );
not \U$303 ( \959 , \958 );
nor \U$304 ( \960 , \941 , \955 , \959 );
and \U$305 ( \961 , \690 , RIb54d768_110);
and \U$306 ( \962 , RIb54d7e0_111, \705 );
nor \U$307 ( \963 , \961 , \962 );
and \U$308 ( \964 , \710 , RIb54db28_118);
and \U$309 ( \965 , RIb54d600_107, \740 );
nor \U$310 ( \966 , \964 , \965 );
and \U$311 ( \967 , \724 , RIb54d678_108);
and \U$312 ( \968 , RIb54d6f0_109, \726 );
nor \U$313 ( \969 , \967 , \968 );
nand \U$314 ( \970 , \960 , \963 , \966 , \969 );
buf \U$315 ( \971 , \970 );
_DC gcc2 ( \972_nGcc2 , \971 , \751 );
xor \U$316 ( \973 , \940 , \972_nGcc2 );
not \U$317 ( \974 , \654 );
not \U$318 ( \975 , RIb54a720_7);
and \U$319 ( \976 , \974 , \975 );
and \U$320 ( \977 , \654 , RIb54a720_7);
nor \U$321 ( \978 , \976 , \977 );
and \U$322 ( \979 , \683 , RIb54dc18_120);
and \U$323 ( \980 , RIb54dfd8_128, \705 );
and \U$324 ( \981 , \734 , RIb54dd08_122);
and \U$325 ( \982 , RIb54dc90_121, \736 );
nor \U$326 ( \983 , \980 , \981 , \982 );
and \U$327 ( \984 , \710 , RIb54e320_135);
and \U$328 ( \985 , RIb54dd80_123, \738 );
nor \U$329 ( \986 , \984 , \985 );
and \U$330 ( \987 , \690 , RIb54df60_127);
and \U$331 ( \988 , RIb54dee8_126, \726 );
nor \U$332 ( \989 , \987 , \988 );
and \U$333 ( \990 , \724 , RIb54de70_125);
and \U$334 ( \991 , RIb54ddf8_124, \740 );
nor \U$335 ( \992 , \990 , \991 );
nand \U$336 ( \993 , \983 , \986 , \989 , \992 );
and \U$337 ( \994 , \703 , RIb54e050_129);
and \U$338 ( \995 , RIb54e0c8_130, \698 );
nor \U$339 ( \996 , \994 , \995 );
not \U$340 ( \997 , \996 );
nor \U$341 ( \998 , \979 , \993 , \997 );
and \U$342 ( \999 , \716 , RIb54e230_133);
and \U$343 ( \1000 , RIb54e2a8_134, \713 );
nor \U$344 ( \1001 , \999 , \1000 );
nand \U$345 ( \1002 , RIb54dba0_119, \732 );
and \U$346 ( \1003 , \695 , RIb54e140_131);
and \U$347 ( \1004 , RIb54e1b8_132, \719 );
nor \U$348 ( \1005 , \1003 , \1004 );
nand \U$349 ( \1006 , \998 , \1001 , \1002 , \1005 );
buf \U$350 ( \1007 , \1006 );
_DC gb97 ( \1008_nGb97 , \1007 , \751 );
xor \U$351 ( \1009 , \978 , \1008_nGb97 );
not \U$352 ( \1010 , \652 );
not \U$353 ( \1011 , RIb54a798_8);
and \U$354 ( \1012 , \1010 , \1011 );
and \U$355 ( \1013 , \652 , RIb54a798_8);
nor \U$356 ( \1014 , \1012 , \1013 );
and \U$357 ( \1015 , RIb54e578_140, \738 );
and \U$358 ( \1016 , RIb54eb18_152, \710 );
and \U$359 ( \1017 , \695 , RIb54e938_148);
and \U$360 ( \1018 , RIb54e410_137, \683 );
nor \U$361 ( \1019 , \1017 , \1018 );
and \U$362 ( \1020 , \690 , RIb54e758_144);
and \U$363 ( \1021 , RIb54e7d0_145, \705 );
nor \U$364 ( \1022 , \1020 , \1021 );
and \U$365 ( \1023 , \734 , RIb54e500_139);
and \U$366 ( \1024 , RIb54e488_138, \736 );
nor \U$367 ( \1025 , \1023 , \1024 );
and \U$368 ( \1026 , \703 , RIb54e848_146);
and \U$369 ( \1027 , RIb54e8c0_147, \698 );
nor \U$370 ( \1028 , \1026 , \1027 );
nand \U$371 ( \1029 , \1019 , \1022 , \1025 , \1028 );
nor \U$372 ( \1030 , \1015 , \1016 , \1029 );
and \U$373 ( \1031 , \716 , RIb54ea28_150);
and \U$374 ( \1032 , RIb54eaa0_151, \713 );
nor \U$375 ( \1033 , \1031 , \1032 );
nand \U$376 ( \1034 , RIb54e398_136, \732 );
and \U$377 ( \1035 , RIb54e9b0_149, \719 );
and \U$378 ( \1036 , RIb54e6e0_143, \726 );
and \U$379 ( \1037 , \724 , RIb54e668_142);
and \U$380 ( \1038 , RIb54e5f0_141, \740 );
nor \U$381 ( \1039 , \1037 , \1038 );
not \U$382 ( \1040 , \1039 );
nor \U$383 ( \1041 , \1035 , \1036 , \1040 );
nand \U$384 ( \1042 , \1030 , \1033 , \1034 , \1041 );
buf \U$385 ( \1043 , \1042 );
_DC gb95 ( \1044_nGb95 , \1043 , \751 );
xor \U$386 ( \1045 , \1014 , \1044_nGb95 );
xnor \U$387 ( \1046 , RIb54a810_9, \651 );
and \U$388 ( \1047 , RIb54ec08_154, \683 );
and \U$389 ( \1048 , RIb54f130_165, \695 );
and \U$390 ( \1049 , \724 , RIb54ee60_159);
and \U$391 ( \1050 , RIb54eed8_160, \726 );
nor \U$392 ( \1051 , \1049 , \1050 );
and \U$393 ( \1052 , \738 , RIb54ed70_157);
and \U$394 ( \1053 , RIb54ede8_158, \740 );
nor \U$395 ( \1054 , \1052 , \1053 );
and \U$396 ( \1055 , \710 , RIb54f310_169);
and \U$397 ( \1056 , RIb54f298_168, \713 );
nor \U$398 ( \1057 , \1055 , \1056 );
and \U$399 ( \1058 , \716 , RIb54f220_167);
and \U$400 ( \1059 , RIb54f1a8_166, \719 );
nor \U$401 ( \1060 , \1058 , \1059 );
nand \U$402 ( \1061 , \1051 , \1054 , \1057 , \1060 );
nor \U$403 ( \1062 , \1047 , \1048 , \1061 );
and \U$404 ( \1063 , \703 , RIb54f040_163);
and \U$405 ( \1064 , RIb54f0b8_164, \698 );
nor \U$406 ( \1065 , \1063 , \1064 );
nand \U$407 ( \1066 , RIb54eb90_153, \732 );
and \U$408 ( \1067 , RIb54ef50_161, \690 );
and \U$409 ( \1068 , RIb54efc8_162, \705 );
and \U$410 ( \1069 , \734 , RIb54ecf8_156);
and \U$411 ( \1070 , RIb54ec80_155, \736 );
nor \U$412 ( \1071 , \1069 , \1070 );
not \U$413 ( \1072 , \1071 );
nor \U$414 ( \1073 , \1067 , \1068 , \1072 );
nand \U$415 ( \1074 , \1062 , \1065 , \1066 , \1073 );
buf \U$416 ( \1075 , \1074 );
_DC gac0 ( \1076_nGac0 , \1075 , \751 );
xor \U$417 ( \1077 , \1046 , \1076_nGac0 );
xnor \U$418 ( \1078 , RIb54a888_10, RIb54a900_11);
and \U$419 ( \1079 , RIb54f400_171, \683 );
and \U$420 ( \1080 , RIb54f928_182, \695 );
and \U$421 ( \1081 , \724 , RIb54f658_176);
and \U$422 ( \1082 , RIb54f6d0_177, \726 );
nor \U$423 ( \1083 , \1081 , \1082 );
and \U$424 ( \1084 , \738 , RIb54f568_174);
and \U$425 ( \1085 , RIb54f5e0_175, \740 );
nor \U$426 ( \1086 , \1084 , \1085 );
and \U$427 ( \1087 , \710 , RIb54fb08_186);
and \U$428 ( \1088 , RIb54fa90_185, \713 );
nor \U$429 ( \1089 , \1087 , \1088 );
and \U$430 ( \1090 , \716 , RIb54fa18_184);
and \U$431 ( \1091 , RIb54f9a0_183, \719 );
nor \U$432 ( \1092 , \1090 , \1091 );
nand \U$433 ( \1093 , \1083 , \1086 , \1089 , \1092 );
nor \U$434 ( \1094 , \1079 , \1080 , \1093 );
and \U$435 ( \1095 , \703 , RIb54f838_180);
and \U$436 ( \1096 , RIb54f8b0_181, \698 );
nor \U$437 ( \1097 , \1095 , \1096 );
nand \U$438 ( \1098 , RIb54f388_170, \732 );
and \U$439 ( \1099 , RIb54f748_178, \690 );
and \U$440 ( \1100 , RIb54f7c0_179, \705 );
and \U$441 ( \1101 , \734 , RIb54f4f0_173);
and \U$442 ( \1102 , RIb54f478_172, \736 );
nor \U$443 ( \1103 , \1101 , \1102 );
not \U$444 ( \1104 , \1103 );
nor \U$445 ( \1105 , \1099 , \1100 , \1104 );
nand \U$446 ( \1106 , \1094 , \1097 , \1098 , \1105 );
buf \U$447 ( \1107 , \1106 );
_DC gac2 ( \1108_nGac2 , \1107 , \751 );
xor \U$448 ( \1109 , \1078 , \1108_nGac2 );
and \U$449 ( \1110 , RIb54fbf8_188, \683 );
and \U$450 ( \1111 , RIb54ff40_195, \690 );
and \U$451 ( \1112 , \695 , RIb550120_199);
and \U$452 ( \1113 , RIb5500a8_198, \698 );
nor \U$453 ( \1114 , \1112 , \1113 );
and \U$454 ( \1115 , \703 , RIb550030_197);
and \U$455 ( \1116 , RIb54ffb8_196, \705 );
nor \U$456 ( \1117 , \1115 , \1116 );
and \U$457 ( \1118 , \710 , RIb550300_203);
and \U$458 ( \1119 , RIb550288_202, \713 );
nor \U$459 ( \1120 , \1118 , \1119 );
and \U$460 ( \1121 , \716 , RIb550210_201);
and \U$461 ( \1122 , RIb550198_200, \719 );
nor \U$462 ( \1123 , \1121 , \1122 );
nand \U$463 ( \1124 , \1114 , \1117 , \1120 , \1123 );
nor \U$464 ( \1125 , \1110 , \1111 , \1124 );
and \U$465 ( \1126 , \724 , RIb54fe50_193);
and \U$466 ( \1127 , RIb54fec8_194, \726 );
nor \U$467 ( \1128 , \1126 , \1127 );
nand \U$468 ( \1129 , RIb54fb80_187, \732 );
and \U$469 ( \1130 , RIb54fce8_190, \734 );
and \U$470 ( \1131 , RIb54fc70_189, \736 );
and \U$471 ( \1132 , \738 , RIb54fd60_191);
and \U$472 ( \1133 , RIb54fdd8_192, \740 );
nor \U$473 ( \1134 , \1132 , \1133 );
not \U$474 ( \1135 , \1134 );
nor \U$475 ( \1136 , \1130 , \1131 , \1135 );
nand \U$476 ( \1137 , \1125 , \1128 , \1129 , \1136 );
buf \U$477 ( \1138 , \1137 );
_DC g95e ( \1139_nG95e , \1138 , \751 );
xor \U$478 ( \1140 , RIb54a900_11, \1139_nG95e );
and \U$479 ( \1141 , \736 , RIb5504e0_207);
and \U$480 ( \1142 , \724 , RIb5506c0_211);
and \U$481 ( \1143 , RIb550648_210, \740 );
nor \U$482 ( \1144 , \1142 , \1143 );
and \U$483 ( \1145 , \726 , RIb550738_212);
nand \U$484 ( \1146 , RIb5503f0_205, \732 );
not \U$485 ( \1147 , \1146 );
nor \U$486 ( \1148 , \1145 , \1147 );
and \U$487 ( \1149 , \698 , RIb550918_216);
and \U$488 ( \1150 , RIb550468_206, \683 );
nor \U$489 ( \1151 , \1149 , \1150 );
and \U$490 ( \1152 , \716 , RIb550a80_219);
and \U$491 ( \1153 , RIb550af8_220, \713 );
nor \U$492 ( \1154 , \1152 , \1153 );
nand \U$493 ( \1155 , \1144 , \1148 , \1151 , \1154 );
and \U$494 ( \1156 , \695 , RIb550990_217);
and \U$495 ( \1157 , RIb550a08_218, \719 );
nor \U$496 ( \1158 , \1156 , \1157 );
not \U$497 ( \1159 , \1158 );
nor \U$498 ( \1160 , \1141 , \1155 , \1159 );
and \U$499 ( \1161 , \703 , RIb5508a0_215);
and \U$500 ( \1162 , RIb550828_214, \705 );
nor \U$501 ( \1163 , \1161 , \1162 );
and \U$502 ( \1164 , \710 , RIb550b70_221);
and \U$503 ( \1165 , RIb550558_208, \734 );
nor \U$504 ( \1166 , \1164 , \1165 );
and \U$505 ( \1167 , \690 , RIb5507b0_213);
and \U$506 ( \1168 , RIb5505d0_209, \738 );
nor \U$507 ( \1169 , \1167 , \1168 );
nand \U$508 ( \1170 , \1160 , \1163 , \1166 , \1169 );
buf \U$509 ( \1171 , \1170 );
_DC g95c ( \1172_nG95c , \1171 , \751 );
not \U$510 ( \1173 , RIb550378_204);
nand \U$511 ( \1174 , \1172_nG95c , \1173 );
not \U$512 ( \1175 , \1174 );
and \U$513 ( \1176 , \1140 , \1175 );
and \U$514 ( \1177 , RIb54a900_11, \1139_nG95e );
or \U$515 ( \1178 , \1176 , \1177 );
and \U$516 ( \1179 , \1109 , \1178 );
and \U$517 ( \1180 , \1078 , \1108_nGac2 );
or \U$518 ( \1181 , \1179 , \1180 );
and \U$519 ( \1182 , \1077 , \1181 );
and \U$520 ( \1183 , \1046 , \1076_nGac0 );
or \U$521 ( \1184 , \1182 , \1183 );
and \U$522 ( \1185 , \1045 , \1184 );
and \U$523 ( \1186 , \1014 , \1044_nGb95 );
or \U$524 ( \1187 , \1185 , \1186 );
and \U$525 ( \1188 , \1009 , \1187 );
and \U$526 ( \1189 , \978 , \1008_nGb97 );
or \U$527 ( \1190 , \1188 , \1189 );
and \U$528 ( \1191 , \973 , \1190 );
and \U$529 ( \1192 , \940 , \972_nGcc2 );
or \U$530 ( \1193 , \1191 , \1192 );
and \U$531 ( \1194 , \935 , \1193 );
and \U$532 ( \1195 , \904 , \934_nGcc4 );
or \U$533 ( \1196 , \1194 , \1195 );
and \U$534 ( \1197 , \899 , \1196 );
and \U$535 ( \1198 , \866 , \898_nGe3f );
or \U$536 ( \1199 , \1197 , \1198 );
and \U$537 ( \1200 , \861 , \1199 );
and \U$538 ( \1201 , \830 , \860_nGe41 );
or \U$539 ( \1202 , \1200 , \1201 );
and \U$540 ( \1203 , \825 , \1202 );
and \U$541 ( \1204 , \794 , \824_nGfef );
or \U$542 ( \1205 , \1203 , \1204 );
and \U$543 ( \1206 , \789 , \1205 );
and \U$544 ( \1207 , \758 , \788_nGff1 );
or \U$545 ( \1208 , \1206 , \1207 );
and \U$546 ( \1209 , \753 , \1208 );
and \U$547 ( \1210 , \673 , \752_nG11dc );
or \U$548 ( \1211 , \1209 , \1210 );
not \U$549 ( \1212 , \668 );
nand \U$550 ( \1213 , \1212 , RIb5517a0_247);
nor \U$551 ( \1214 , \1211 , \1213 );
not \U$552 ( \1215 , \1214 );
and \U$553 ( \1216 , RIb551020_231, \736 );
and \U$554 ( \1217 , RIb5512f0_237, \690 );
and \U$555 ( \1218 , \738 , RIb551110_233);
and \U$556 ( \1219 , RIb551098_232, \734 );
nor \U$557 ( \1220 , \1218 , \1219 );
and \U$558 ( \1221 , \695 , RIb5514d0_241);
and \U$559 ( \1222 , RIb551548_242, \719 );
nor \U$560 ( \1223 , \1221 , \1222 );
or \U$561 ( \1224 , \683 , \732 );
and \U$562 ( \1225 , \1224 , RIb550be8_222);
and \U$563 ( \1226 , RIb551458_240, \698 );
nor \U$564 ( \1227 , \1225 , \1226 );
and \U$565 ( \1228 , \724 , RIb551200_235);
and \U$566 ( \1229 , RIb551188_234, \740 );
nor \U$567 ( \1230 , \1228 , \1229 );
nand \U$568 ( \1231 , \1220 , \1223 , \1227 , \1230 );
nor \U$569 ( \1232 , \1216 , \1217 , \1231 );
and \U$570 ( \1233 , \710 , RIb5516b0_245);
and \U$571 ( \1234 , RIb5515c0_243, \716 );
nor \U$572 ( \1235 , \1233 , \1234 );
and \U$573 ( \1236 , \713 , RIb551638_244);
and \U$574 ( \1237 , RIb551278_236, \726 );
nor \U$575 ( \1238 , \1236 , \1237 );
and \U$576 ( \1239 , \703 , RIb5513e0_239);
and \U$577 ( \1240 , RIb551368_238, \705 );
nor \U$578 ( \1241 , \1239 , \1240 );
nand \U$579 ( \1242 , \1232 , \1235 , \1238 , \1241 );
buf \U$580 ( \1243 , \750 );
_DC g1807 ( \1244_nG1807 , \1242 , \1243 );
not \U$581 ( \1245 , \1244_nG1807 );
nor \U$582 ( \1246 , \1215 , \1245 );
xor \U$583 ( \1247 , \673 , \752_nG11dc );
xor \U$584 ( \1248 , \1247 , \1208 );
not \U$585 ( \1249 , \1248 );
xor \U$586 ( \1250 , \758 , \788_nGff1 );
xor \U$587 ( \1251 , \1250 , \1205 );
not \U$588 ( \1252 , \1251 );
and \U$589 ( \1253 , \1249 , \1252 );
and \U$590 ( \1254 , \1211 , \1213 );
nor \U$591 ( \1255 , \1254 , \1214 );
nor \U$592 ( \1256 , \1253 , \1255 );
not \U$593 ( \1257 , \1256 );
and \U$594 ( \1258 , \1255 , \1248 );
nor \U$595 ( \1259 , \1255 , \1248 );
xnor \U$596 ( \1260 , \1251 , \1248 );
not \U$597 ( \1261 , \1260 );
nor \U$598 ( \1262 , \1258 , \1259 , \1261 );
nand \U$599 ( \1263 , \1257 , \1262 );
and \U$600 ( \1264 , RIb552088_266, \736 );
and \U$601 ( \1265 , RIb552448_274, \703 );
and \U$602 ( \1266 , \738 , RIb552178_268);
and \U$603 ( \1267 , RIb552100_267, \734 );
nor \U$604 ( \1268 , \1266 , \1267 );
and \U$605 ( \1269 , \695 , RIb552538_276);
and \U$606 ( \1270 , RIb5525b0_277, \719 );
nor \U$607 ( \1271 , \1269 , \1270 );
and \U$608 ( \1272 , \1224 , RIb552010_265);
and \U$609 ( \1273 , RIb5524c0_275, \698 );
nor \U$610 ( \1274 , \1272 , \1273 );
and \U$611 ( \1275 , \724 , RIb552268_270);
and \U$612 ( \1276 , RIb5521f0_269, \740 );
nor \U$613 ( \1277 , \1275 , \1276 );
nand \U$614 ( \1278 , \1268 , \1271 , \1274 , \1277 );
nor \U$615 ( \1279 , \1264 , \1265 , \1278 );
and \U$616 ( \1280 , \690 , RIb552358_272);
and \U$617 ( \1281 , RIb5523d0_273, \705 );
nor \U$618 ( \1282 , \1280 , \1281 );
and \U$619 ( \1283 , \710 , RIb552718_280);
and \U$620 ( \1284 , RIb5522e0_271, \726 );
nor \U$621 ( \1285 , \1283 , \1284 );
and \U$622 ( \1286 , \716 , RIb552628_278);
and \U$623 ( \1287 , RIb5526a0_279, \713 );
nor \U$624 ( \1288 , \1286 , \1287 );
nand \U$625 ( \1289 , \1279 , \1282 , \1285 , \1288 );
_DC g191a ( \1290_nG191a , \1289 , \1243 );
not \U$626 ( \1291 , \1290_nG191a );
or \U$627 ( \1292 , \1263 , \1291 );
or \U$628 ( \1293 , \1290_nG191a , \1257 );
or \U$629 ( \1294 , \1257 , \1262 );
nand \U$630 ( \1295 , \1292 , \1293 , \1294 );
xnor \U$631 ( \1296 , \1246 , \1295 );
nand \U$632 ( \1297 , \1261 , \1257 );
or \U$633 ( \1298 , \1297 , \1291 );
or \U$634 ( \1299 , \1245 , \1263 );
or \U$635 ( \1300 , \1260 , \1291 );
or \U$636 ( \1301 , \1257 , \1244_nG1807 );
nand \U$637 ( \1302 , \1301 , \1294 );
nand \U$638 ( \1303 , \1300 , \1302 );
nand \U$639 ( \1304 , \1298 , \1299 , \1303 );
xor \U$640 ( \1305 , \794 , \824_nGfef );
xor \U$641 ( \1306 , \1305 , \1202 );
xor \U$642 ( \1307 , \830 , \860_nGe41 );
xor \U$643 ( \1308 , \1307 , \1199 );
nor \U$644 ( \1309 , \1306 , \1308 );
or \U$645 ( \1310 , \1251 , \1309 );
and \U$646 ( \1311 , \1304 , \1310 );
and \U$647 ( \1312 , RIb552880_283, \736 );
and \U$648 ( \1313 , RIb552b50_289, \690 );
and \U$649 ( \1314 , \724 , RIb552a60_287);
and \U$650 ( \1315 , RIb5529e8_286, \740 );
nor \U$651 ( \1316 , \1314 , \1315 );
and \U$652 ( \1317 , \738 , RIb552970_285);
and \U$653 ( \1318 , RIb552cb8_292, \698 );
nor \U$654 ( \1319 , \1317 , \1318 );
and \U$655 ( \1320 , \1224 , RIb552808_282);
and \U$656 ( \1321 , RIb5528f8_284, \734 );
nor \U$657 ( \1322 , \1320 , \1321 );
and \U$658 ( \1323 , \695 , RIb552d30_293);
and \U$659 ( \1324 , RIb552da8_294, \719 );
nor \U$660 ( \1325 , \1323 , \1324 );
nand \U$661 ( \1326 , \1316 , \1319 , \1322 , \1325 );
nor \U$662 ( \1327 , \1312 , \1313 , \1326 );
and \U$663 ( \1328 , \703 , RIb552c40_291);
and \U$664 ( \1329 , RIb552ad8_288, \726 );
nor \U$665 ( \1330 , \1328 , \1329 );
and \U$666 ( \1331 , \710 , RIb552f10_297);
and \U$667 ( \1332 , RIb552bc8_290, \705 );
nor \U$668 ( \1333 , \1331 , \1332 );
and \U$669 ( \1334 , \716 , RIb552e20_295);
and \U$670 ( \1335 , RIb552e98_296, \713 );
nor \U$671 ( \1336 , \1334 , \1335 );
nand \U$672 ( \1337 , \1327 , \1330 , \1333 , \1336 );
_DC g1711 ( \1338_nG1711 , \1337 , \1243 );
not \U$673 ( \1339 , \1338_nG1711 );
nor \U$674 ( \1340 , \1215 , \1339 );
nor \U$675 ( \1341 , \1311 , \1340 );
xor \U$676 ( \1342 , \1296 , \1341 );
not \U$677 ( \1343 , \1342 );
not \U$678 ( \1344 , \1306 );
not \U$679 ( \1345 , \1251 );
or \U$680 ( \1346 , \1344 , \1345 );
or \U$681 ( \1347 , \1251 , \1306 );
nand \U$682 ( \1348 , \1346 , \1347 );
xor \U$683 ( \1349 , \1308 , \1306 );
nor \U$684 ( \1350 , \1348 , \1349 );
not \U$685 ( \1351 , \1350 );
not \U$686 ( \1352 , \1310 );
nor \U$687 ( \1353 , \1351 , \1352 );
not \U$688 ( \1354 , \1353 );
or \U$689 ( \1355 , \1354 , \1291 );
or \U$690 ( \1356 , \1351 , \1291 );
nand \U$691 ( \1357 , \1356 , \1352 );
nand \U$692 ( \1358 , \1355 , \1357 );
or \U$693 ( \1359 , \1297 , \1245 );
or \U$694 ( \1360 , \1339 , \1263 );
or \U$695 ( \1361 , \1260 , \1245 );
or \U$696 ( \1362 , \1257 , \1338_nG1711 );
nand \U$697 ( \1363 , \1362 , \1294 );
nand \U$698 ( \1364 , \1361 , \1363 );
nand \U$699 ( \1365 , \1359 , \1360 , \1364 );
and \U$700 ( \1366 , \1358 , \1365 );
and \U$701 ( \1367 , \1304 , \1310 );
not \U$702 ( \1368 , \1304 );
and \U$703 ( \1369 , \1368 , \1352 );
nor \U$704 ( \1370 , \1367 , \1369 );
xor \U$705 ( \1371 , \1340 , \1370 );
and \U$706 ( \1372 , \1366 , \1371 );
xor \U$707 ( \1373 , \1343 , \1372 );
nand \U$708 ( \1374 , \1244_nG1807 , \1350 );
or \U$709 ( \1375 , \1310 , \1290_nG191a );
or \U$710 ( \1376 , \1310 , \1349 );
nand \U$711 ( \1377 , \1375 , \1376 );
and \U$712 ( \1378 , \1374 , \1377 );
and \U$713 ( \1379 , \1310 , \1349 );
and \U$714 ( \1380 , \1379 , \1290_nG191a );
and \U$715 ( \1381 , \1244_nG1807 , \1353 );
nor \U$716 ( \1382 , \1378 , \1380 , \1381 );
not \U$717 ( \1383 , \1297 );
and \U$718 ( \1384 , \1338_nG1711 , \1383 );
and \U$719 ( \1385 , RIb553ca8_326, \698 );
and \U$720 ( \1386 , RIb5538e8_318, \734 );
and \U$721 ( \1387 , \703 , RIb553c30_325);
and \U$722 ( \1388 , RIb553bb8_324, \705 );
nor \U$723 ( \1389 , \1387 , \1388 );
and \U$724 ( \1390 , \716 , RIb553e10_329);
and \U$725 ( \1391 , RIb553870_317, \736 );
nor \U$726 ( \1392 , \1390 , \1391 );
and \U$727 ( \1393 , \710 , RIb553f00_331);
and \U$728 ( \1394 , RIb553e88_330, \713 );
nor \U$729 ( \1395 , \1393 , \1394 );
and \U$730 ( \1396 , \690 , RIb553b40_323);
and \U$731 ( \1397 , RIb553ac8_322, \726 );
nor \U$732 ( \1398 , \1396 , \1397 );
nand \U$733 ( \1399 , \1389 , \1392 , \1395 , \1398 );
nor \U$734 ( \1400 , \1385 , \1386 , \1399 );
and \U$735 ( \1401 , \1224 , RIb5537f8_316);
and \U$736 ( \1402 , RIb553a50_321, \724 );
nor \U$737 ( \1403 , \1401 , \1402 );
and \U$738 ( \1404 , \719 , RIb553d98_328);
and \U$739 ( \1405 , RIb5539d8_320, \740 );
nor \U$740 ( \1406 , \1404 , \1405 );
and \U$741 ( \1407 , \695 , RIb553d20_327);
and \U$742 ( \1408 , RIb553960_319, \738 );
nor \U$743 ( \1409 , \1407 , \1408 );
nand \U$744 ( \1410 , \1400 , \1403 , \1406 , \1409 );
_DC g15f9 ( \1411_nG15f9 , \1410 , \1243 );
or \U$745 ( \1412 , \1257 , \1411_nG15f9 );
nand \U$746 ( \1413 , \1412 , \1294 );
nand \U$747 ( \1414 , \1338_nG1711 , \1261 );
and \U$748 ( \1415 , \1413 , \1414 );
not \U$749 ( \1416 , \1263 );
and \U$750 ( \1417 , \1411_nG15f9 , \1416 );
nor \U$751 ( \1418 , \1384 , \1415 , \1417 );
nand \U$752 ( \1419 , \1382 , \1418 );
xor \U$753 ( \1420 , \866 , \898_nGe3f );
xor \U$754 ( \1421 , \1420 , \1196 );
xor \U$755 ( \1422 , \904 , \934_nGcc4 );
xor \U$756 ( \1423 , \1422 , \1193 );
nor \U$757 ( \1424 , \1421 , \1423 );
or \U$758 ( \1425 , \1308 , \1424 );
and \U$759 ( \1426 , \1419 , \1425 );
nor \U$760 ( \1427 , \1418 , \1382 );
nor \U$761 ( \1428 , \1426 , \1427 );
xor \U$762 ( \1429 , \1358 , \1365 );
not \U$763 ( \1430 , \1429 );
nand \U$764 ( \1431 , \1411_nG15f9 , \1214 );
not \U$765 ( \1432 , \1431 );
and \U$766 ( \1433 , \1430 , \1432 );
and \U$767 ( \1434 , \1429 , \1431 );
nor \U$768 ( \1435 , \1433 , \1434 );
nand \U$769 ( \1436 , \1428 , \1435 );
xor \U$770 ( \1437 , \1366 , \1371 );
and \U$771 ( \1438 , \1436 , \1437 );
and \U$772 ( \1439 , \1373 , \1438 );
not \U$773 ( \1440 , \1439 );
and \U$774 ( \1441 , \1343 , \1372 );
or \U$775 ( \1442 , \1441 , \1256 );
and \U$776 ( \1443 , \1295 , \1246 );
and \U$777 ( \1444 , \1256 , \1441 );
nor \U$778 ( \1445 , \1443 , \1444 );
nand \U$779 ( \1446 , \1442 , \1445 );
not \U$780 ( \1447 , \1446 );
and \U$781 ( \1448 , \1214 , \1290_nG191a );
and \U$782 ( \1449 , \1296 , \1341 );
nor \U$783 ( \1450 , \1448 , \1449 );
not \U$784 ( \1451 , \1450 );
and \U$785 ( \1452 , \1447 , \1451 );
and \U$786 ( \1453 , \1446 , \1450 );
nor \U$787 ( \1454 , \1452 , \1453 );
not \U$788 ( \1455 , \1454 );
or \U$789 ( \1456 , \1440 , \1455 );
or \U$790 ( \1457 , \1454 , \1439 );
nand \U$791 ( \1458 , \1456 , \1457 );
not \U$792 ( \1459 , \1458 );
xor \U$793 ( \1460 , \1436 , \1437 );
not \U$794 ( \1461 , \1429 );
nor \U$795 ( \1462 , \1461 , \1431 );
xor \U$796 ( \1463 , \1460 , \1462 );
or \U$797 ( \1464 , \1435 , \1428 );
nand \U$798 ( \1465 , \1464 , \1436 );
not \U$799 ( \1466 , \1465 );
and \U$800 ( \1467 , RIb553078_300, \736 );
and \U$801 ( \1468 , RIb553438_308, \703 );
and \U$802 ( \1469 , \738 , RIb553168_302);
and \U$803 ( \1470 , RIb5530f0_301, \734 );
nor \U$804 ( \1471 , \1469 , \1470 );
and \U$805 ( \1472 , \695 , RIb553528_310);
and \U$806 ( \1473 , RIb5535a0_311, \719 );
nor \U$807 ( \1474 , \1472 , \1473 );
and \U$808 ( \1475 , \1224 , RIb553000_299);
and \U$809 ( \1476 , RIb5534b0_309, \698 );
nor \U$810 ( \1477 , \1475 , \1476 );
and \U$811 ( \1478 , \724 , RIb553258_304);
and \U$812 ( \1479 , RIb5531e0_303, \740 );
nor \U$813 ( \1480 , \1478 , \1479 );
nand \U$814 ( \1481 , \1471 , \1474 , \1477 , \1480 );
nor \U$815 ( \1482 , \1467 , \1468 , \1481 );
and \U$816 ( \1483 , \690 , RIb553348_306);
and \U$817 ( \1484 , RIb5533c0_307, \705 );
nor \U$818 ( \1485 , \1483 , \1484 );
and \U$819 ( \1486 , \710 , RIb553708_314);
and \U$820 ( \1487 , RIb5532d0_305, \726 );
nor \U$821 ( \1488 , \1486 , \1487 );
and \U$822 ( \1489 , \716 , RIb553618_312);
and \U$823 ( \1490 , RIb553690_313, \713 );
nor \U$824 ( \1491 , \1489 , \1490 );
nand \U$825 ( \1492 , \1482 , \1485 , \1488 , \1491 );
_DC g14ed ( \1493_nG14ed , \1492 , \1243 );
not \U$826 ( \1494 , \1493_nG14ed );
nor \U$827 ( \1495 , \1215 , \1494 );
not \U$828 ( \1496 , \1425 );
not \U$829 ( \1497 , \1427 );
nand \U$830 ( \1498 , \1497 , \1419 );
not \U$831 ( \1499 , \1498 );
or \U$832 ( \1500 , \1496 , \1499 );
or \U$833 ( \1501 , \1498 , \1425 );
nand \U$834 ( \1502 , \1500 , \1501 );
xnor \U$835 ( \1503 , \1495 , \1502 );
not \U$836 ( \1504 , \1503 );
and \U$837 ( \1505 , \1411_nG15f9 , \1383 );
or \U$838 ( \1506 , \1257 , \1493_nG14ed );
nand \U$839 ( \1507 , \1506 , \1294 );
nand \U$840 ( \1508 , \1411_nG15f9 , \1261 );
and \U$841 ( \1509 , \1507 , \1508 );
and \U$842 ( \1510 , \1493_nG14ed , \1416 );
nor \U$843 ( \1511 , \1505 , \1509 , \1510 );
and \U$844 ( \1512 , RIb5541d0_337, \740 );
and \U$845 ( \1513 , RIb5544a0_343, \698 );
and \U$846 ( \1514 , \703 , RIb554428_342);
and \U$847 ( \1515 , RIb5543b0_341, \705 );
nor \U$848 ( \1516 , \1514 , \1515 );
and \U$849 ( \1517 , \710 , RIb5546f8_348);
and \U$850 ( \1518 , RIb554338_340, \690 );
nor \U$851 ( \1519 , \1517 , \1518 );
and \U$852 ( \1520 , \726 , RIb5542c0_339);
and \U$853 ( \1521 , RIb554068_334, \736 );
nor \U$854 ( \1522 , \1520 , \1521 );
and \U$855 ( \1523 , \716 , RIb554608_346);
and \U$856 ( \1524 , RIb554680_347, \713 );
nor \U$857 ( \1525 , \1523 , \1524 );
nand \U$858 ( \1526 , \1516 , \1519 , \1522 , \1525 );
nor \U$859 ( \1527 , \1512 , \1513 , \1526 );
and \U$860 ( \1528 , \1224 , RIb553ff0_333);
and \U$861 ( \1529 , RIb554158_336, \738 );
nor \U$862 ( \1530 , \1528 , \1529 );
and \U$863 ( \1531 , \719 , RIb554590_345);
and \U$864 ( \1532 , RIb5540e0_335, \734 );
nor \U$865 ( \1533 , \1531 , \1532 );
and \U$866 ( \1534 , \695 , RIb554518_344);
and \U$867 ( \1535 , RIb554248_338, \724 );
nor \U$868 ( \1536 , \1534 , \1535 );
nand \U$869 ( \1537 , \1527 , \1530 , \1533 , \1536 );
_DC g13f2 ( \1538_nG13f2 , \1537 , \1243 );
nand \U$870 ( \1539 , \1538_nG13f2 , \1214 );
or \U$871 ( \1540 , \1511 , \1539 );
and \U$872 ( \1541 , \1308 , \1421 );
nor \U$873 ( \1542 , \1308 , \1421 );
xor \U$874 ( \1543 , \1421 , \1423 );
nor \U$875 ( \1544 , \1541 , \1542 , \1543 );
and \U$876 ( \1545 , \1544 , \1425 );
and \U$877 ( \1546 , \1290_nG191a , \1545 );
not \U$878 ( \1547 , \1425 );
and \U$879 ( \1548 , \1291 , \1547 );
or \U$880 ( \1549 , \1544 , \1425 );
not \U$881 ( \1550 , \1549 );
nor \U$882 ( \1551 , \1546 , \1548 , \1550 );
nand \U$883 ( \1552 , \1338_nG1711 , \1350 );
or \U$884 ( \1553 , \1310 , \1244_nG1807 );
nand \U$885 ( \1554 , \1553 , \1376 );
and \U$886 ( \1555 , \1552 , \1554 );
and \U$887 ( \1556 , \1379 , \1244_nG1807 );
and \U$888 ( \1557 , \1338_nG1711 , \1353 );
nor \U$889 ( \1558 , \1555 , \1556 , \1557 );
or \U$890 ( \1559 , \1551 , \1558 );
nand \U$891 ( \1560 , \1540 , \1559 );
nand \U$892 ( \1561 , \1504 , \1560 );
nor \U$893 ( \1562 , \1466 , \1561 );
and \U$894 ( \1563 , \1463 , \1562 );
and \U$895 ( \1564 , \1460 , \1462 );
or \U$896 ( \1565 , \1563 , \1564 );
xor \U$897 ( \1566 , \1373 , \1438 );
xor \U$898 ( \1567 , \1565 , \1566 );
xor \U$899 ( \1568 , \1460 , \1462 );
xor \U$900 ( \1569 , \1568 , \1562 );
and \U$901 ( \1570 , \1502 , \1495 );
xor \U$902 ( \1571 , \940 , \972_nGcc2 );
xor \U$903 ( \1572 , \1571 , \1190 );
xor \U$904 ( \1573 , \978 , \1008_nGb97 );
xor \U$905 ( \1574 , \1573 , \1187 );
nor \U$906 ( \1575 , \1572 , \1574 );
or \U$907 ( \1576 , \1423 , \1575 );
not \U$908 ( \1577 , \1576 );
nand \U$909 ( \1578 , \1411_nG15f9 , \1350 );
or \U$910 ( \1579 , \1310 , \1338_nG1711 );
nand \U$911 ( \1580 , \1579 , \1376 );
and \U$912 ( \1581 , \1578 , \1580 );
and \U$913 ( \1582 , \1379 , \1338_nG1711 );
and \U$914 ( \1583 , \1411_nG15f9 , \1353 );
nor \U$915 ( \1584 , \1581 , \1582 , \1583 );
nand \U$916 ( \1585 , \1290_nG191a , \1543 );
or \U$917 ( \1586 , \1425 , \1244_nG1807 );
nand \U$918 ( \1587 , \1586 , \1549 );
and \U$919 ( \1588 , \1585 , \1587 );
and \U$920 ( \1589 , \1545 , \1244_nG1807 );
not \U$921 ( \1590 , \1543 );
nor \U$922 ( \1591 , \1547 , \1590 );
and \U$923 ( \1592 , \1290_nG191a , \1591 );
nor \U$924 ( \1593 , \1588 , \1589 , \1592 );
nor \U$925 ( \1594 , \1584 , \1593 );
not \U$926 ( \1595 , \1594 );
nand \U$927 ( \1596 , \1593 , \1584 );
nand \U$928 ( \1597 , \1595 , \1596 );
not \U$929 ( \1598 , \1597 );
or \U$930 ( \1599 , \1577 , \1598 );
or \U$931 ( \1600 , \1597 , \1576 );
nand \U$932 ( \1601 , \1599 , \1600 );
and \U$933 ( \1602 , RIb555238_372, \724 );
and \U$934 ( \1603 , RIb5550d0_369, \734 );
and \U$935 ( \1604 , \713 , RIb555670_381);
and \U$936 ( \1605 , RIb555418_376, \703 );
nor \U$937 ( \1606 , \1604 , \1605 );
and \U$938 ( \1607 , \705 , RIb5553a0_375);
and \U$939 ( \1608 , RIb555058_368, \736 );
nor \U$940 ( \1609 , \1607 , \1608 );
and \U$941 ( \1610 , \710 , RIb5556e8_382);
and \U$942 ( \1611 , RIb555490_377, \698 );
nor \U$943 ( \1612 , \1610 , \1611 );
and \U$944 ( \1613 , \716 , RIb5555f8_380);
and \U$945 ( \1614 , RIb555580_379, \719 );
nor \U$946 ( \1615 , \1613 , \1614 );
nand \U$947 ( \1616 , \1606 , \1609 , \1612 , \1615 );
nor \U$948 ( \1617 , \1602 , \1603 , \1616 );
and \U$949 ( \1618 , \738 , RIb555148_370);
and \U$950 ( \1619 , RIb5551c0_371, \740 );
nor \U$951 ( \1620 , \1618 , \1619 );
and \U$952 ( \1621 , \695 , RIb555508_378);
and \U$953 ( \1622 , RIb5552b0_373, \726 );
nor \U$954 ( \1623 , \1621 , \1622 );
and \U$955 ( \1624 , \1224 , RIb554fe0_367);
and \U$956 ( \1625 , RIb555328_374, \690 );
nor \U$957 ( \1626 , \1624 , \1625 );
nand \U$958 ( \1627 , \1617 , \1620 , \1623 , \1626 );
_DC g1300 ( \1628_nG1300 , \1627 , \1243 );
not \U$959 ( \1629 , \1628_nG1300 );
nor \U$960 ( \1630 , \1215 , \1629 );
or \U$961 ( \1631 , \1297 , \1494 );
not \U$962 ( \1632 , \1538_nG13f2 );
or \U$963 ( \1633 , \1632 , \1263 );
or \U$964 ( \1634 , \1260 , \1494 );
or \U$965 ( \1635 , \1257 , \1538_nG13f2 );
nand \U$966 ( \1636 , \1635 , \1294 );
nand \U$967 ( \1637 , \1634 , \1636 );
nand \U$968 ( \1638 , \1631 , \1633 , \1637 );
xor \U$969 ( \1639 , \1630 , \1638 );
and \U$970 ( \1640 , \1601 , \1639 );
not \U$971 ( \1641 , \1572 );
not \U$972 ( \1642 , \1423 );
or \U$973 ( \1643 , \1641 , \1642 );
or \U$974 ( \1644 , \1423 , \1572 );
nand \U$975 ( \1645 , \1643 , \1644 );
xor \U$976 ( \1646 , \1574 , \1572 );
nor \U$977 ( \1647 , \1645 , \1646 );
not \U$978 ( \1648 , \1647 );
not \U$979 ( \1649 , \1576 );
nor \U$980 ( \1650 , \1648 , \1649 );
not \U$981 ( \1651 , \1650 );
or \U$982 ( \1652 , \1651 , \1291 );
or \U$983 ( \1653 , \1648 , \1291 );
nand \U$984 ( \1654 , \1653 , \1649 );
nand \U$985 ( \1655 , \1652 , \1654 );
not \U$986 ( \1656 , \1591 );
or \U$987 ( \1657 , \1656 , \1245 );
not \U$988 ( \1658 , \1545 );
or \U$989 ( \1659 , \1339 , \1658 );
or \U$990 ( \1660 , \1590 , \1245 );
or \U$991 ( \1661 , \1425 , \1338_nG1711 );
nand \U$992 ( \1662 , \1661 , \1549 );
nand \U$993 ( \1663 , \1660 , \1662 );
nand \U$994 ( \1664 , \1657 , \1659 , \1663 );
and \U$995 ( \1665 , \1655 , \1664 );
and \U$996 ( \1666 , \1538_nG13f2 , \1383 );
or \U$997 ( \1667 , \1257 , \1628_nG1300 );
nand \U$998 ( \1668 , \1667 , \1294 );
nand \U$999 ( \1669 , \1538_nG13f2 , \1261 );
and \U$1000 ( \1670 , \1668 , \1669 );
and \U$1001 ( \1671 , \1628_nG1300 , \1416 );
nor \U$1002 ( \1672 , \1666 , \1670 , \1671 );
nand \U$1003 ( \1673 , \1493_nG14ed , \1350 );
or \U$1004 ( \1674 , \1310 , \1411_nG15f9 );
nand \U$1005 ( \1675 , \1674 , \1376 );
and \U$1006 ( \1676 , \1673 , \1675 );
and \U$1007 ( \1677 , \1379 , \1411_nG15f9 );
and \U$1008 ( \1678 , \1493_nG14ed , \1353 );
nor \U$1009 ( \1679 , \1676 , \1677 , \1678 );
and \U$1010 ( \1680 , \1672 , \1679 );
and \U$1011 ( \1681 , RIb5548d8_352, \734 );
and \U$1012 ( \1682 , RIb554b30_357, \690 );
and \U$1013 ( \1683 , \695 , RIb554d10_361);
and \U$1014 ( \1684 , RIb554e78_364, \713 );
nor \U$1015 ( \1685 , \1683 , \1684 );
and \U$1016 ( \1686 , \698 , RIb554c98_360);
and \U$1017 ( \1687 , RIb554860_351, \736 );
nor \U$1018 ( \1688 , \1686 , \1687 );
and \U$1019 ( \1689 , \710 , RIb554ef0_365);
and \U$1020 ( \1690 , RIb554d88_362, \719 );
nor \U$1021 ( \1691 , \1689 , \1690 );
and \U$1022 ( \1692 , \716 , RIb554e00_363);
and \U$1023 ( \1693 , RIb554ab8_356, \726 );
nor \U$1024 ( \1694 , \1692 , \1693 );
nand \U$1025 ( \1695 , \1685 , \1688 , \1691 , \1694 );
nor \U$1026 ( \1696 , \1681 , \1682 , \1695 );
and \U$1027 ( \1697 , \738 , RIb554950_353);
and \U$1028 ( \1698 , RIb5549c8_354, \740 );
nor \U$1029 ( \1699 , \1697 , \1698 );
and \U$1030 ( \1700 , \724 , RIb554a40_355);
and \U$1031 ( \1701 , RIb554ba8_358, \705 );
nor \U$1032 ( \1702 , \1700 , \1701 );
and \U$1033 ( \1703 , \1224 , RIb5547e8_350);
and \U$1034 ( \1704 , RIb554c20_359, \703 );
nor \U$1035 ( \1705 , \1703 , \1704 );
nand \U$1036 ( \1706 , \1696 , \1699 , \1702 , \1705 );
_DC g11f7 ( \1707_nG11f7 , \1706 , \1243 );
nand \U$1037 ( \1708 , \1707_nG11f7 , \1214 );
or \U$1038 ( \1709 , \1680 , \1708 );
or \U$1039 ( \1710 , \1672 , \1679 );
nand \U$1040 ( \1711 , \1709 , \1710 );
and \U$1041 ( \1712 , \1665 , \1711 );
and \U$1042 ( \1713 , \1640 , \1712 );
and \U$1043 ( \1714 , \1596 , \1576 );
and \U$1044 ( \1715 , \1630 , \1638 );
nor \U$1045 ( \1716 , \1714 , \1715 , \1594 );
xnor \U$1046 ( \1717 , \1539 , \1511 );
not \U$1047 ( \1718 , \1717 );
xor \U$1048 ( \1719 , \1551 , \1558 );
not \U$1049 ( \1720 , \1719 );
and \U$1050 ( \1721 , \1718 , \1720 );
and \U$1051 ( \1722 , \1717 , \1719 );
nor \U$1052 ( \1723 , \1721 , \1722 );
nand \U$1053 ( \1724 , \1716 , \1723 );
xor \U$1054 ( \1725 , \1713 , \1724 );
not \U$1055 ( \1726 , \1560 );
not \U$1056 ( \1727 , \1503 );
or \U$1057 ( \1728 , \1726 , \1727 );
or \U$1058 ( \1729 , \1503 , \1560 );
nand \U$1059 ( \1730 , \1728 , \1729 );
and \U$1060 ( \1731 , \1725 , \1730 );
and \U$1061 ( \1732 , \1713 , \1724 );
or \U$1062 ( \1733 , \1731 , \1732 );
nor \U$1063 ( \1734 , \1570 , \1733 );
not \U$1064 ( \1735 , \1465 );
not \U$1065 ( \1736 , \1561 );
and \U$1066 ( \1737 , \1735 , \1736 );
and \U$1067 ( \1738 , \1465 , \1561 );
nor \U$1068 ( \1739 , \1737 , \1738 );
nor \U$1069 ( \1740 , \1734 , \1739 );
xor \U$1070 ( \1741 , \1569 , \1740 );
and \U$1071 ( \1742 , \1734 , \1739 );
nor \U$1072 ( \1743 , \1742 , \1740 );
xor \U$1073 ( \1744 , \1601 , \1639 );
xor \U$1074 ( \1745 , \1665 , \1711 );
and \U$1075 ( \1746 , \1744 , \1745 );
and \U$1076 ( \1747 , \1628_nG1300 , \1383 );
or \U$1077 ( \1748 , \1257 , \1707_nG11f7 );
nand \U$1078 ( \1749 , \1748 , \1294 );
nand \U$1079 ( \1750 , \1628_nG1300 , \1261 );
and \U$1080 ( \1751 , \1749 , \1750 );
and \U$1081 ( \1752 , \1707_nG11f7 , \1416 );
nor \U$1082 ( \1753 , \1747 , \1751 , \1752 );
nand \U$1083 ( \1754 , \1538_nG13f2 , \1350 );
or \U$1084 ( \1755 , \1310 , \1493_nG14ed );
nand \U$1085 ( \1756 , \1755 , \1376 );
and \U$1086 ( \1757 , \1754 , \1756 );
and \U$1087 ( \1758 , \1379 , \1493_nG14ed );
and \U$1088 ( \1759 , \1538_nG13f2 , \1353 );
nor \U$1089 ( \1760 , \1757 , \1758 , \1759 );
and \U$1090 ( \1761 , \1753 , \1760 );
not \U$1091 ( \1762 , \1761 );
and \U$1092 ( \1763 , RIb556048_402, \736 );
and \U$1093 ( \1764 , RIb556480_411, \698 );
and \U$1094 ( \1765 , \1224 , RIb555fd0_401);
and \U$1095 ( \1766 , RIb556228_406, \724 );
nor \U$1096 ( \1767 , \1765 , \1766 );
and \U$1097 ( \1768 , \695 , RIb5564f8_412);
and \U$1098 ( \1769 , RIb556570_413, \719 );
nor \U$1099 ( \1770 , \1768 , \1769 );
and \U$1100 ( \1771 , \726 , RIb5562a0_407);
and \U$1101 ( \1772 , RIb5561b0_405, \740 );
nor \U$1102 ( \1773 , \1771 , \1772 );
and \U$1103 ( \1774 , \738 , RIb556138_404);
and \U$1104 ( \1775 , RIb5560c0_403, \734 );
nor \U$1105 ( \1776 , \1774 , \1775 );
nand \U$1106 ( \1777 , \1767 , \1770 , \1773 , \1776 );
nor \U$1107 ( \1778 , \1763 , \1764 , \1777 );
and \U$1108 ( \1779 , \710 , RIb5566d8_416);
and \U$1109 ( \1780 , RIb5565e8_414, \716 );
nor \U$1110 ( \1781 , \1779 , \1780 );
and \U$1111 ( \1782 , \713 , RIb556660_415);
and \U$1112 ( \1783 , RIb556408_410, \703 );
nor \U$1113 ( \1784 , \1782 , \1783 );
and \U$1114 ( \1785 , \690 , RIb556318_408);
and \U$1115 ( \1786 , RIb556390_409, \705 );
nor \U$1116 ( \1787 , \1785 , \1786 );
nand \U$1117 ( \1788 , \1778 , \1781 , \1784 , \1787 );
_DC g1116 ( \1789_nG1116 , \1788 , \1243 );
nand \U$1118 ( \1790 , \1789_nG1116 , \1214 );
not \U$1119 ( \1791 , \1790 );
and \U$1120 ( \1792 , \1762 , \1791 );
nor \U$1121 ( \1793 , \1753 , \1760 );
nor \U$1122 ( \1794 , \1792 , \1793 );
and \U$1123 ( \1795 , \1244_nG1807 , \1650 );
nand \U$1124 ( \1796 , \1244_nG1807 , \1647 );
or \U$1125 ( \1797 , \1576 , \1290_nG191a );
or \U$1126 ( \1798 , \1576 , \1646 );
nand \U$1127 ( \1799 , \1797 , \1798 );
and \U$1128 ( \1800 , \1796 , \1799 );
and \U$1129 ( \1801 , \1576 , \1646 );
and \U$1130 ( \1802 , \1290_nG191a , \1801 );
nor \U$1131 ( \1803 , \1795 , \1800 , \1802 );
not \U$1132 ( \1804 , \1803 );
xor \U$1133 ( \1805 , \1014 , \1044_nGb95 );
xor \U$1134 ( \1806 , \1805 , \1184 );
xor \U$1135 ( \1807 , \1046 , \1076_nGac0 );
xor \U$1136 ( \1808 , \1807 , \1181 );
nor \U$1137 ( \1809 , \1806 , \1808 );
or \U$1138 ( \1810 , \1574 , \1809 );
not \U$1139 ( \1811 , \1810 );
not \U$1140 ( \1812 , \1811 );
and \U$1141 ( \1813 , \1804 , \1812 );
and \U$1142 ( \1814 , \1803 , \1811 );
nand \U$1143 ( \1815 , \1338_nG1711 , \1543 );
or \U$1144 ( \1816 , \1425 , \1411_nG15f9 );
nand \U$1145 ( \1817 , \1816 , \1549 );
and \U$1146 ( \1818 , \1815 , \1817 );
and \U$1147 ( \1819 , \1545 , \1411_nG15f9 );
and \U$1148 ( \1820 , \1338_nG1711 , \1591 );
nor \U$1149 ( \1821 , \1818 , \1819 , \1820 );
nor \U$1150 ( \1822 , \1814 , \1821 );
nor \U$1151 ( \1823 , \1813 , \1822 );
nor \U$1152 ( \1824 , \1794 , \1823 );
xor \U$1153 ( \1825 , \1655 , \1664 );
not \U$1154 ( \1826 , \1825 );
not \U$1155 ( \1827 , \1710 );
nor \U$1156 ( \1828 , \1827 , \1680 );
not \U$1157 ( \1829 , \1828 );
not \U$1158 ( \1830 , \1708 );
and \U$1159 ( \1831 , \1829 , \1830 );
and \U$1160 ( \1832 , \1828 , \1708 );
nor \U$1161 ( \1833 , \1831 , \1832 );
nor \U$1162 ( \1834 , \1826 , \1833 );
and \U$1163 ( \1835 , \1824 , \1834 );
xor \U$1164 ( \1836 , \1746 , \1835 );
or \U$1165 ( \1837 , \1723 , \1716 );
nand \U$1166 ( \1838 , \1837 , \1724 );
and \U$1167 ( \1839 , \1836 , \1838 );
and \U$1168 ( \1840 , \1746 , \1835 );
or \U$1169 ( \1841 , \1839 , \1840 );
not \U$1170 ( \1842 , \1719 );
nor \U$1171 ( \1843 , \1842 , \1717 );
xor \U$1172 ( \1844 , \1841 , \1843 );
xor \U$1173 ( \1845 , \1713 , \1724 );
xor \U$1174 ( \1846 , \1845 , \1730 );
and \U$1175 ( \1847 , \1844 , \1846 );
and \U$1176 ( \1848 , \1841 , \1843 );
or \U$1177 ( \1849 , \1847 , \1848 );
xor \U$1178 ( \1850 , \1743 , \1849 );
xnor \U$1179 ( \1851 , \1823 , \1794 );
not \U$1180 ( \1852 , \1833 );
not \U$1181 ( \1853 , \1825 );
and \U$1182 ( \1854 , \1852 , \1853 );
and \U$1183 ( \1855 , \1833 , \1825 );
nor \U$1184 ( \1856 , \1854 , \1855 );
nand \U$1185 ( \1857 , \1851 , \1856 );
not \U$1186 ( \1858 , \1806 );
not \U$1187 ( \1859 , \1574 );
or \U$1188 ( \1860 , \1858 , \1859 );
or \U$1189 ( \1861 , \1574 , \1806 );
nand \U$1190 ( \1862 , \1860 , \1861 );
xor \U$1191 ( \1863 , \1808 , \1806 );
nor \U$1192 ( \1864 , \1862 , \1863 );
not \U$1193 ( \1865 , \1864 );
nor \U$1194 ( \1866 , \1865 , \1811 );
not \U$1195 ( \1867 , \1866 );
or \U$1196 ( \1868 , \1867 , \1291 );
or \U$1197 ( \1869 , \1865 , \1291 );
nand \U$1198 ( \1870 , \1869 , \1811 );
nand \U$1199 ( \1871 , \1868 , \1870 );
or \U$1200 ( \1872 , \1651 , \1339 );
not \U$1201 ( \1873 , \1801 );
or \U$1202 ( \1874 , \1245 , \1873 );
or \U$1203 ( \1875 , \1648 , \1339 );
or \U$1204 ( \1876 , \1576 , \1244_nG1807 );
nand \U$1205 ( \1877 , \1876 , \1798 );
nand \U$1206 ( \1878 , \1875 , \1877 );
nand \U$1207 ( \1879 , \1872 , \1874 , \1878 );
and \U$1208 ( \1880 , \1871 , \1879 );
nand \U$1209 ( \1881 , \1628_nG1300 , \1350 );
or \U$1210 ( \1882 , \1310 , \1538_nG13f2 );
nand \U$1211 ( \1883 , \1882 , \1376 );
and \U$1212 ( \1884 , \1881 , \1883 );
and \U$1213 ( \1885 , \1379 , \1538_nG13f2 );
and \U$1214 ( \1886 , \1628_nG1300 , \1353 );
nor \U$1215 ( \1887 , \1884 , \1885 , \1886 );
nand \U$1216 ( \1888 , \1411_nG15f9 , \1543 );
or \U$1217 ( \1889 , \1425 , \1493_nG14ed );
nand \U$1218 ( \1890 , \1889 , \1549 );
and \U$1219 ( \1891 , \1888 , \1890 );
and \U$1220 ( \1892 , \1545 , \1493_nG14ed );
and \U$1221 ( \1893 , \1411_nG15f9 , \1591 );
nor \U$1222 ( \1894 , \1891 , \1892 , \1893 );
xor \U$1223 ( \1895 , \1887 , \1894 );
and \U$1224 ( \1896 , \1707_nG11f7 , \1383 );
or \U$1225 ( \1897 , \1257 , \1789_nG1116 );
nand \U$1226 ( \1898 , \1897 , \1294 );
nand \U$1227 ( \1899 , \1707_nG11f7 , \1261 );
and \U$1228 ( \1900 , \1898 , \1899 );
and \U$1229 ( \1901 , \1789_nG1116 , \1416 );
nor \U$1230 ( \1902 , \1896 , \1900 , \1901 );
and \U$1231 ( \1903 , \1895 , \1902 );
and \U$1232 ( \1904 , \1887 , \1894 );
or \U$1233 ( \1905 , \1903 , \1904 );
not \U$1234 ( \1906 , \1905 );
and \U$1235 ( \1907 , \1880 , \1906 );
not \U$1236 ( \1908 , \1803 );
or \U$1237 ( \1909 , \1821 , \1810 );
nand \U$1238 ( \1910 , \1810 , \1821 );
nand \U$1239 ( \1911 , \1909 , \1910 );
not \U$1240 ( \1912 , \1911 );
or \U$1241 ( \1913 , \1908 , \1912 );
or \U$1242 ( \1914 , \1911 , \1803 );
nand \U$1243 ( \1915 , \1913 , \1914 );
not \U$1244 ( \1916 , \1790 );
nor \U$1245 ( \1917 , \1761 , \1793 );
not \U$1246 ( \1918 , \1917 );
or \U$1247 ( \1919 , \1916 , \1918 );
or \U$1248 ( \1920 , \1917 , \1790 );
nand \U$1249 ( \1921 , \1919 , \1920 );
and \U$1250 ( \1922 , \1915 , \1921 );
and \U$1251 ( \1923 , \1907 , \1922 );
xor \U$1252 ( \1924 , \1857 , \1923 );
xor \U$1253 ( \1925 , \1744 , \1745 );
and \U$1254 ( \1926 , \1924 , \1925 );
and \U$1255 ( \1927 , \1857 , \1923 );
or \U$1256 ( \1928 , \1926 , \1927 );
xor \U$1257 ( \1929 , \1640 , \1712 );
xor \U$1258 ( \1930 , \1928 , \1929 );
xor \U$1259 ( \1931 , \1746 , \1835 );
xor \U$1260 ( \1932 , \1931 , \1838 );
and \U$1261 ( \1933 , \1930 , \1932 );
and \U$1262 ( \1934 , \1928 , \1929 );
or \U$1263 ( \1935 , \1933 , \1934 );
xor \U$1264 ( \1936 , \1841 , \1843 );
xor \U$1265 ( \1937 , \1936 , \1846 );
xor \U$1266 ( \1938 , \1935 , \1937 );
xor \U$1267 ( \1939 , \1928 , \1929 );
xor \U$1268 ( \1940 , \1939 , \1932 );
xor \U$1269 ( \1941 , \1824 , \1834 );
xor \U$1270 ( \1942 , \1857 , \1923 );
xor \U$1271 ( \1943 , \1942 , \1925 );
and \U$1272 ( \1944 , \1941 , \1943 );
xor \U$1273 ( \1945 , \1880 , \1906 );
xor \U$1274 ( \1946 , \1915 , \1921 );
and \U$1275 ( \1947 , \1945 , \1946 );
xor \U$1276 ( \1948 , \1871 , \1879 );
xor \U$1277 ( \1949 , \1887 , \1894 );
xor \U$1278 ( \1950 , \1949 , \1902 );
not \U$1279 ( \1951 , \1950 );
and \U$1280 ( \1952 , \1948 , \1951 );
or \U$1281 ( \1953 , \1867 , \1245 );
and \U$1282 ( \1954 , \1810 , \1863 );
not \U$1283 ( \1955 , \1954 );
or \U$1284 ( \1956 , \1291 , \1955 );
or \U$1285 ( \1957 , \1865 , \1245 );
or \U$1286 ( \1958 , \1810 , \1290_nG191a );
or \U$1287 ( \1959 , \1810 , \1863 );
nand \U$1288 ( \1960 , \1958 , \1959 );
nand \U$1289 ( \1961 , \1957 , \1960 );
nand \U$1290 ( \1962 , \1953 , \1956 , \1961 );
xor \U$1291 ( \1963 , RIb54a900_11, \1139_nG95e );
xor \U$1292 ( \1964 , \1963 , \1175 );
not \U$1293 ( \1965 , \1964 );
xor \U$1294 ( \1966 , \1078 , \1108_nGac2 );
xor \U$1295 ( \1967 , \1966 , \1178 );
not \U$1296 ( \1968 , \1967 );
and \U$1297 ( \1969 , \1965 , \1968 );
or \U$1298 ( \1970 , \1808 , \1969 );
xor \U$1299 ( \1971 , \1962 , \1970 );
not \U$1300 ( \1972 , \1411_nG15f9 );
or \U$1301 ( \1973 , \1651 , \1972 );
or \U$1302 ( \1974 , \1339 , \1873 );
or \U$1303 ( \1975 , \1648 , \1972 );
or \U$1304 ( \1976 , \1576 , \1338_nG1711 );
nand \U$1305 ( \1977 , \1976 , \1798 );
nand \U$1306 ( \1978 , \1975 , \1977 );
nand \U$1307 ( \1979 , \1973 , \1974 , \1978 );
and \U$1308 ( \1980 , \1971 , \1979 );
and \U$1309 ( \1981 , \1962 , \1970 );
or \U$1310 ( \1982 , \1980 , \1981 );
nand \U$1311 ( \1983 , \1707_nG11f7 , \1350 );
or \U$1312 ( \1984 , \1310 , \1628_nG1300 );
nand \U$1313 ( \1985 , \1984 , \1376 );
and \U$1314 ( \1986 , \1983 , \1985 );
and \U$1315 ( \1987 , \1379 , \1628_nG1300 );
and \U$1316 ( \1988 , \1707_nG11f7 , \1353 );
nor \U$1317 ( \1989 , \1986 , \1987 , \1988 );
nand \U$1318 ( \1990 , \1493_nG14ed , \1543 );
or \U$1319 ( \1991 , \1425 , \1538_nG13f2 );
nand \U$1320 ( \1992 , \1991 , \1549 );
and \U$1321 ( \1993 , \1990 , \1992 );
and \U$1322 ( \1994 , \1545 , \1538_nG13f2 );
and \U$1323 ( \1995 , \1493_nG14ed , \1591 );
nor \U$1324 ( \1996 , \1993 , \1994 , \1995 );
xor \U$1325 ( \1997 , \1989 , \1996 );
and \U$1326 ( \1998 , \1789_nG1116 , \1383 );
and \U$1327 ( \1999 , RIb555c88_394, \698 );
and \U$1328 ( \2000 , RIb5558c8_386, \734 );
and \U$1329 ( \2001 , \703 , RIb555c10_393);
and \U$1330 ( \2002 , RIb555b98_392, \705 );
nor \U$1331 ( \2003 , \2001 , \2002 );
and \U$1332 ( \2004 , \710 , RIb555ee0_399);
and \U$1333 ( \2005 , RIb555b20_391, \690 );
nor \U$1334 ( \2006 , \2004 , \2005 );
and \U$1335 ( \2007 , \726 , RIb555aa8_390);
and \U$1336 ( \2008 , RIb555850_385, \736 );
nor \U$1337 ( \2009 , \2007 , \2008 );
and \U$1338 ( \2010 , \716 , RIb555df0_397);
and \U$1339 ( \2011 , RIb555e68_398, \713 );
nor \U$1340 ( \2012 , \2010 , \2011 );
nand \U$1341 ( \2013 , \2003 , \2006 , \2009 , \2012 );
nor \U$1342 ( \2014 , \1999 , \2000 , \2013 );
and \U$1343 ( \2015 , \738 , RIb555940_387);
and \U$1344 ( \2016 , RIb5559b8_388, \740 );
nor \U$1345 ( \2017 , \2015 , \2016 );
and \U$1346 ( \2018 , \1224 , RIb5557d8_384);
and \U$1347 ( \2019 , RIb555d78_396, \719 );
nor \U$1348 ( \2020 , \2018 , \2019 );
and \U$1349 ( \2021 , \695 , RIb555d00_395);
and \U$1350 ( \2022 , RIb555a30_389, \724 );
nor \U$1351 ( \2023 , \2021 , \2022 );
nand \U$1352 ( \2024 , \2014 , \2017 , \2020 , \2023 );
_DC g100c ( \2025_nG100c , \2024 , \1243 );
or \U$1353 ( \2026 , \1257 , \2025_nG100c );
nand \U$1354 ( \2027 , \2026 , \1294 );
nand \U$1355 ( \2028 , \1789_nG1116 , \1261 );
and \U$1356 ( \2029 , \2027 , \2028 );
and \U$1357 ( \2030 , \2025_nG100c , \1416 );
nor \U$1358 ( \2031 , \1998 , \2029 , \2030 );
and \U$1359 ( \2032 , \1997 , \2031 );
and \U$1360 ( \2033 , \1989 , \1996 );
or \U$1361 ( \2034 , \2032 , \2033 );
not \U$1362 ( \2035 , \2034 );
and \U$1363 ( \2036 , \1982 , \2035 );
and \U$1364 ( \2037 , \1952 , \2036 );
xor \U$1365 ( \2038 , \1947 , \2037 );
or \U$1366 ( \2039 , \1856 , \1851 );
nand \U$1367 ( \2040 , \2039 , \1857 );
and \U$1368 ( \2041 , \2038 , \2040 );
and \U$1369 ( \2042 , \1947 , \2037 );
or \U$1370 ( \2043 , \2041 , \2042 );
xor \U$1371 ( \2044 , \1857 , \1923 );
xor \U$1372 ( \2045 , \2044 , \1925 );
and \U$1373 ( \2046 , \2043 , \2045 );
and \U$1374 ( \2047 , \1941 , \2043 );
or \U$1375 ( \2048 , \1944 , \2046 , \2047 );
xor \U$1376 ( \2049 , \1940 , \2048 );
xor \U$1377 ( \2050 , \1948 , \1951 );
nand \U$1378 ( \2051 , \2025_nG100c , \1214 );
and \U$1379 ( \2052 , \2050 , \2051 );
xor \U$1380 ( \2053 , \1982 , \2035 );
nor \U$1381 ( \2054 , \2052 , \2053 );
and \U$1382 ( \2055 , RIb5570b0_437, \734 );
and \U$1383 ( \2056 , RIb557290_441, \726 );
and \U$1384 ( \2057 , \724 , RIb557218_440);
and \U$1385 ( \2058 , RIb557560_447, \719 );
nor \U$1386 ( \2059 , \2057 , \2058 );
and \U$1387 ( \2060 , \703 , RIb5573f8_444);
and \U$1388 ( \2061 , RIb557470_445, \698 );
nor \U$1389 ( \2062 , \2060 , \2061 );
and \U$1390 ( \2063 , \710 , RIb5576c8_450);
and \U$1391 ( \2064 , RIb557650_449, \713 );
nor \U$1392 ( \2065 , \2063 , \2064 );
and \U$1393 ( \2066 , \695 , RIb5574e8_446);
and \U$1394 ( \2067 , RIb557038_436, \736 );
nor \U$1395 ( \2068 , \2066 , \2067 );
nand \U$1396 ( \2069 , \2059 , \2062 , \2065 , \2068 );
nor \U$1397 ( \2070 , \2055 , \2056 , \2069 );
and \U$1398 ( \2071 , \1224 , RIb556fc0_435);
and \U$1399 ( \2072 , RIb5575d8_448, \716 );
nor \U$1400 ( \2073 , \2071 , \2072 );
and \U$1401 ( \2074 , \740 , RIb5571a0_439);
and \U$1402 ( \2075 , RIb557380_443, \705 );
nor \U$1403 ( \2076 , \2074 , \2075 );
and \U$1404 ( \2077 , \690 , RIb557308_442);
and \U$1405 ( \2078 , RIb557128_438, \738 );
nor \U$1406 ( \2079 , \2077 , \2078 );
nand \U$1407 ( \2080 , \2070 , \2073 , \2076 , \2079 );
_DC gf30 ( \2081_nGf30 , \2080 , \1243 );
nand \U$1408 ( \2082 , \2081_nGf30 , \1214 );
not \U$1409 ( \2083 , \2082 );
xor \U$1410 ( \2084 , \1962 , \1970 );
xor \U$1411 ( \2085 , \2084 , \1979 );
xor \U$1412 ( \2086 , \1989 , \1996 );
xor \U$1413 ( \2087 , \2086 , \2031 );
not \U$1414 ( \2088 , \2087 );
and \U$1415 ( \2089 , \2085 , \2088 );
nor \U$1416 ( \2090 , \2083 , \2089 );
not \U$1417 ( \2091 , \2090 );
not \U$1418 ( \2092 , \1967 );
not \U$1419 ( \2093 , \1808 );
or \U$1420 ( \2094 , \2092 , \2093 );
or \U$1421 ( \2095 , \1808 , \1967 );
nand \U$1422 ( \2096 , \2094 , \2095 );
xor \U$1423 ( \2097 , \1965 , \1968 );
nor \U$1424 ( \2098 , \2096 , \2097 );
nand \U$1425 ( \2099 , \1970 , \2098 );
or \U$1426 ( \2100 , \2099 , \1291 );
not \U$1427 ( \2101 , \2098 );
or \U$1428 ( \2102 , \2101 , \1291 );
not \U$1429 ( \2103 , \1970 );
nand \U$1430 ( \2104 , \2102 , \2103 );
nand \U$1431 ( \2105 , \2100 , \2104 );
not \U$1432 ( \2106 , \2105 );
nand \U$1433 ( \2107 , \1338_nG1711 , \1864 );
or \U$1434 ( \2108 , \1810 , \1244_nG1807 );
nand \U$1435 ( \2109 , \2108 , \1959 );
and \U$1436 ( \2110 , \2107 , \2109 );
and \U$1437 ( \2111 , \1954 , \1244_nG1807 );
and \U$1438 ( \2112 , \1338_nG1711 , \1866 );
nor \U$1439 ( \2113 , \2110 , \2111 , \2112 );
nor \U$1440 ( \2114 , \2106 , \2113 );
not \U$1441 ( \2115 , \2114 );
nand \U$1442 ( \2116 , \1538_nG13f2 , \1543 );
or \U$1443 ( \2117 , \1425 , \1628_nG1300 );
nand \U$1444 ( \2118 , \2117 , \1549 );
and \U$1445 ( \2119 , \2116 , \2118 );
and \U$1446 ( \2120 , \1545 , \1628_nG1300 );
and \U$1447 ( \2121 , \1538_nG13f2 , \1591 );
nor \U$1448 ( \2122 , \2119 , \2120 , \2121 );
and \U$1449 ( \2123 , \1493_nG14ed , \1650 );
nand \U$1450 ( \2124 , \1493_nG14ed , \1647 );
or \U$1451 ( \2125 , \1576 , \1411_nG15f9 );
nand \U$1452 ( \2126 , \2125 , \1798 );
and \U$1453 ( \2127 , \2124 , \2126 );
and \U$1454 ( \2128 , \1411_nG15f9 , \1801 );
nor \U$1455 ( \2129 , \2123 , \2127 , \2128 );
xor \U$1456 ( \2130 , \2122 , \2129 );
nand \U$1457 ( \2131 , \1789_nG1116 , \1350 );
or \U$1458 ( \2132 , \1310 , \1707_nG11f7 );
nand \U$1459 ( \2133 , \2132 , \1376 );
and \U$1460 ( \2134 , \2131 , \2133 );
and \U$1461 ( \2135 , \1379 , \1707_nG11f7 );
and \U$1462 ( \2136 , \1789_nG1116 , \1353 );
nor \U$1463 ( \2137 , \2134 , \2135 , \2136 );
and \U$1464 ( \2138 , \2130 , \2137 );
and \U$1465 ( \2139 , \2122 , \2129 );
or \U$1466 ( \2140 , \2138 , \2139 );
nor \U$1467 ( \2141 , \2115 , \2140 );
nand \U$1468 ( \2142 , \2091 , \2141 );
or \U$1469 ( \2143 , \2054 , \2142 );
not \U$1470 ( \2144 , \2142 );
not \U$1471 ( \2145 , \2054 );
or \U$1472 ( \2146 , \2144 , \2145 );
xor \U$1473 ( \2147 , \1945 , \1946 );
nand \U$1474 ( \2148 , \2146 , \2147 );
nand \U$1475 ( \2149 , \2143 , \2148 );
xor \U$1476 ( \2150 , \1907 , \1922 );
xor \U$1477 ( \2151 , \2149 , \2150 );
xor \U$1478 ( \2152 , \1947 , \2037 );
xor \U$1479 ( \2153 , \2152 , \2040 );
and \U$1480 ( \2154 , \2151 , \2153 );
and \U$1481 ( \2155 , \2149 , \2150 );
or \U$1482 ( \2156 , \2154 , \2155 );
xor \U$1483 ( \2157 , \1857 , \1923 );
xor \U$1484 ( \2158 , \2157 , \1925 );
xor \U$1485 ( \2159 , \1941 , \2043 );
xor \U$1486 ( \2160 , \2158 , \2159 );
xor \U$1487 ( \2161 , \2156 , \2160 );
xor \U$1488 ( \2162 , \2149 , \2150 );
xor \U$1489 ( \2163 , \2162 , \2153 );
not \U$1490 ( \2164 , \2053 );
xnor \U$1491 ( \2165 , \2051 , \2050 );
not \U$1492 ( \2166 , \2165 );
or \U$1493 ( \2167 , \2164 , \2166 );
or \U$1494 ( \2168 , \2165 , \2053 );
nand \U$1495 ( \2169 , \2167 , \2168 );
nand \U$1496 ( \2170 , \1628_nG1300 , \1543 );
or \U$1497 ( \2171 , \1425 , \1707_nG11f7 );
nand \U$1498 ( \2172 , \2171 , \1549 );
and \U$1499 ( \2173 , \2170 , \2172 );
and \U$1500 ( \2174 , \1545 , \1707_nG11f7 );
and \U$1501 ( \2175 , \1628_nG1300 , \1591 );
nor \U$1502 ( \2176 , \2173 , \2174 , \2175 );
and \U$1503 ( \2177 , \1538_nG13f2 , \1650 );
nand \U$1504 ( \2178 , \1538_nG13f2 , \1647 );
or \U$1505 ( \2179 , \1576 , \1493_nG14ed );
nand \U$1506 ( \2180 , \2179 , \1798 );
and \U$1507 ( \2181 , \2178 , \2180 );
and \U$1508 ( \2182 , \1493_nG14ed , \1801 );
nor \U$1509 ( \2183 , \2177 , \2181 , \2182 );
xor \U$1510 ( \2184 , \2176 , \2183 );
nand \U$1511 ( \2185 , \2025_nG100c , \1350 );
or \U$1512 ( \2186 , \1310 , \1789_nG1116 );
nand \U$1513 ( \2187 , \2186 , \1376 );
and \U$1514 ( \2188 , \2185 , \2187 );
and \U$1515 ( \2189 , \1379 , \1789_nG1116 );
and \U$1516 ( \2190 , \2025_nG100c , \1353 );
nor \U$1517 ( \2191 , \2188 , \2189 , \2190 );
and \U$1518 ( \2192 , \2184 , \2191 );
and \U$1519 ( \2193 , \2176 , \2183 );
or \U$1520 ( \2194 , \2192 , \2193 );
nand \U$1521 ( \2195 , \1244_nG1807 , \2098 );
or \U$1522 ( \2196 , \1970 , \1290_nG191a );
or \U$1523 ( \2197 , \1970 , \2097 );
nand \U$1524 ( \2198 , \2196 , \2197 );
and \U$1525 ( \2199 , \2195 , \2198 );
nand \U$1526 ( \2200 , \2097 , \1970 );
not \U$1527 ( \2201 , \2200 );
and \U$1528 ( \2202 , \2201 , \1290_nG191a );
not \U$1529 ( \2203 , \2099 );
and \U$1530 ( \2204 , \1244_nG1807 , \2203 );
nor \U$1531 ( \2205 , \2199 , \2202 , \2204 );
nand \U$1532 ( \2206 , \1411_nG15f9 , \1864 );
or \U$1533 ( \2207 , \1810 , \1338_nG1711 );
nand \U$1534 ( \2208 , \2207 , \1959 );
and \U$1535 ( \2209 , \2206 , \2208 );
and \U$1536 ( \2210 , \1954 , \1338_nG1711 );
and \U$1537 ( \2211 , \1411_nG15f9 , \1866 );
nor \U$1538 ( \2212 , \2209 , \2210 , \2211 );
nand \U$1539 ( \2213 , \2205 , \2212 );
and \U$1540 ( \2214 , \2213 , \1964 );
nor \U$1541 ( \2215 , \2212 , \2205 );
nor \U$1542 ( \2216 , \2214 , \2215 );
nor \U$1543 ( \2217 , \2194 , \2216 );
not \U$1544 ( \2218 , \2113 );
not \U$1545 ( \2219 , \2105 );
and \U$1546 ( \2220 , \2218 , \2219 );
and \U$1547 ( \2221 , \2113 , \2105 );
nor \U$1548 ( \2222 , \2220 , \2221 );
xor \U$1549 ( \2223 , \2122 , \2129 );
xor \U$1550 ( \2224 , \2223 , \2137 );
and \U$1551 ( \2225 , \2222 , \2224 );
and \U$1552 ( \2226 , RIb556e58_432, \713 );
and \U$1553 ( \2227 , RIb556840_419, \736 );
and \U$1554 ( \2228 , \738 , RIb556930_421);
and \U$1555 ( \2229 , RIb5569a8_422, \740 );
nor \U$1556 ( \2230 , \2228 , \2229 );
and \U$1557 ( \2231 , \719 , RIb556d68_430);
and \U$1558 ( \2232 , RIb556b88_426, \705 );
nor \U$1559 ( \2233 , \2231 , \2232 );
and \U$1560 ( \2234 , \1224 , RIb5567c8_418);
and \U$1561 ( \2235 , RIb5568b8_420, \734 );
nor \U$1562 ( \2236 , \2234 , \2235 );
and \U$1563 ( \2237 , \703 , RIb556c00_427);
and \U$1564 ( \2238 , RIb556c78_428, \698 );
nor \U$1565 ( \2239 , \2237 , \2238 );
nand \U$1566 ( \2240 , \2230 , \2233 , \2236 , \2239 );
nor \U$1567 ( \2241 , \2226 , \2227 , \2240 );
and \U$1568 ( \2242 , \724 , RIb556a20_423);
and \U$1569 ( \2243 , RIb556a98_424, \726 );
nor \U$1570 ( \2244 , \2242 , \2243 );
and \U$1571 ( \2245 , \710 , RIb556ed0_433);
and \U$1572 ( \2246 , RIb556cf0_429, \695 );
nor \U$1573 ( \2247 , \2245 , \2246 );
and \U$1574 ( \2248 , \716 , RIb556de0_431);
and \U$1575 ( \2249 , RIb556b10_425, \690 );
nor \U$1576 ( \2250 , \2248 , \2249 );
nand \U$1577 ( \2251 , \2241 , \2244 , \2247 , \2250 );
_DC ge5c ( \2252_nGe5c , \2251 , \1243 );
nand \U$1578 ( \2253 , \2252_nGe5c , \1214 );
and \U$1579 ( \2254 , \2025_nG100c , \1383 );
or \U$1580 ( \2255 , \1257 , \2081_nGf30 );
nand \U$1581 ( \2256 , \2255 , \1294 );
nand \U$1582 ( \2257 , \2025_nG100c , \1261 );
and \U$1583 ( \2258 , \2256 , \2257 );
and \U$1584 ( \2259 , \2081_nGf30 , \1416 );
nor \U$1585 ( \2260 , \2254 , \2258 , \2259 );
xnor \U$1586 ( \2261 , \2253 , \2260 );
xor \U$1587 ( \2262 , \2122 , \2129 );
xor \U$1588 ( \2263 , \2262 , \2137 );
and \U$1589 ( \2264 , \2261 , \2263 );
and \U$1590 ( \2265 , \2222 , \2261 );
or \U$1591 ( \2266 , \2225 , \2264 , \2265 );
not \U$1592 ( \2267 , \2266 );
and \U$1593 ( \2268 , \2217 , \2267 );
nor \U$1594 ( \2269 , \2169 , \2268 );
xor \U$1595 ( \2270 , \2085 , \2088 );
not \U$1596 ( \2271 , \2270 );
not \U$1597 ( \2272 , \2082 );
and \U$1598 ( \2273 , \2271 , \2272 );
and \U$1599 ( \2274 , \2270 , \2082 );
nor \U$1600 ( \2275 , \2273 , \2274 );
not \U$1601 ( \2276 , \2275 );
or \U$1602 ( \2277 , \2140 , \2114 );
or \U$1603 ( \2278 , \2253 , \2260 );
nand \U$1604 ( \2279 , \2114 , \2140 );
nand \U$1605 ( \2280 , \2277 , \2278 , \2279 );
nand \U$1606 ( \2281 , \2276 , \2280 );
or \U$1607 ( \2282 , \2269 , \2281 );
nand \U$1608 ( \2283 , \2268 , \2169 );
nand \U$1609 ( \2284 , \2282 , \2283 );
not \U$1610 ( \2285 , \1952 );
not \U$1611 ( \2286 , \2051 );
nor \U$1612 ( \2287 , \2286 , \2036 );
not \U$1613 ( \2288 , \2287 );
or \U$1614 ( \2289 , \2285 , \2288 );
or \U$1615 ( \2290 , \1952 , \2287 );
nand \U$1616 ( \2291 , \2289 , \2290 );
nor \U$1617 ( \2292 , \2284 , \2291 );
xnor \U$1618 ( \2293 , \2142 , \2054 );
not \U$1619 ( \2294 , \2293 );
not \U$1620 ( \2295 , \2147 );
and \U$1621 ( \2296 , \2294 , \2295 );
and \U$1622 ( \2297 , \2293 , \2147 );
nor \U$1623 ( \2298 , \2296 , \2297 );
or \U$1624 ( \2299 , \2292 , \2298 );
nand \U$1625 ( \2300 , \2291 , \2284 );
nand \U$1626 ( \2301 , \2299 , \2300 );
xor \U$1627 ( \2302 , \2163 , \2301 );
not \U$1628 ( \2303 , \2280 );
not \U$1629 ( \2304 , \2275 );
or \U$1630 ( \2305 , \2303 , \2304 );
or \U$1631 ( \2306 , \2275 , \2280 );
nand \U$1632 ( \2307 , \2305 , \2306 );
xor \U$1633 ( \2308 , \2217 , \2267 );
and \U$1634 ( \2309 , \2307 , \2308 );
not \U$1635 ( \2310 , \2307 );
not \U$1636 ( \2311 , \2308 );
and \U$1637 ( \2312 , \2310 , \2311 );
and \U$1638 ( \2313 , \1628_nG1300 , \1650 );
nand \U$1639 ( \2314 , \1628_nG1300 , \1647 );
or \U$1640 ( \2315 , \1576 , \1538_nG13f2 );
nand \U$1641 ( \2316 , \2315 , \1798 );
and \U$1642 ( \2317 , \2314 , \2316 );
and \U$1643 ( \2318 , \1538_nG13f2 , \1801 );
nor \U$1644 ( \2319 , \2313 , \2317 , \2318 );
nand \U$1645 ( \2320 , \1493_nG14ed , \1864 );
or \U$1646 ( \2321 , \1810 , \1411_nG15f9 );
nand \U$1647 ( \2322 , \2321 , \1959 );
and \U$1648 ( \2323 , \2320 , \2322 );
and \U$1649 ( \2324 , \1954 , \1411_nG15f9 );
and \U$1650 ( \2325 , \1493_nG14ed , \1866 );
nor \U$1651 ( \2326 , \2323 , \2324 , \2325 );
xor \U$1652 ( \2327 , \2319 , \2326 );
nand \U$1653 ( \2328 , \1707_nG11f7 , \1543 );
or \U$1654 ( \2329 , \1425 , \1789_nG1116 );
nand \U$1655 ( \2330 , \2329 , \1549 );
and \U$1656 ( \2331 , \2328 , \2330 );
and \U$1657 ( \2332 , \1545 , \1789_nG1116 );
and \U$1658 ( \2333 , \1707_nG11f7 , \1591 );
nor \U$1659 ( \2334 , \2331 , \2332 , \2333 );
and \U$1660 ( \2335 , \2327 , \2334 );
and \U$1661 ( \2336 , \2319 , \2326 );
or \U$1662 ( \2337 , \2335 , \2336 );
and \U$1663 ( \2338 , \2252_nGe5c , \1383 );
and \U$1664 ( \2339 , RIb558028_470, \736 );
and \U$1665 ( \2340 , RIb558460_479, \698 );
and \U$1666 ( \2341 , \724 , RIb558208_474);
and \U$1667 ( \2342 , RIb558190_473, \740 );
nor \U$1668 ( \2343 , \2341 , \2342 );
and \U$1669 ( \2344 , \710 , RIb5586b8_484);
and \U$1670 ( \2345 , RIb5582f8_476, \690 );
nor \U$1671 ( \2346 , \2344 , \2345 );
and \U$1672 ( \2347 , \713 , RIb558640_483);
and \U$1673 ( \2348 , RIb558280_475, \726 );
nor \U$1674 ( \2349 , \2347 , \2348 );
and \U$1675 ( \2350 , \703 , RIb5583e8_478);
and \U$1676 ( \2351 , RIb558370_477, \705 );
nor \U$1677 ( \2352 , \2350 , \2351 );
nand \U$1678 ( \2353 , \2343 , \2346 , \2349 , \2352 );
nor \U$1679 ( \2354 , \2339 , \2340 , \2353 );
and \U$1680 ( \2355 , \716 , RIb5585c8_482);
and \U$1681 ( \2356 , RIb5580a0_471, \734 );
nor \U$1682 ( \2357 , \2355 , \2356 );
and \U$1683 ( \2358 , \695 , RIb5584d8_480);
and \U$1684 ( \2359 , RIb558550_481, \719 );
nor \U$1685 ( \2360 , \2358 , \2359 );
and \U$1686 ( \2361 , \1224 , RIb557fb0_469);
and \U$1687 ( \2362 , RIb558118_472, \738 );
nor \U$1688 ( \2363 , \2361 , \2362 );
nand \U$1689 ( \2364 , \2354 , \2357 , \2360 , \2363 );
_DC gda9 ( \2365_nGda9 , \2364 , \1243 );
or \U$1690 ( \2366 , \1257 , \2365_nGda9 );
nand \U$1691 ( \2367 , \2366 , \1294 );
nand \U$1692 ( \2368 , \2252_nGe5c , \1261 );
and \U$1693 ( \2369 , \2367 , \2368 );
and \U$1694 ( \2370 , \2365_nGda9 , \1416 );
nor \U$1695 ( \2371 , \2338 , \2369 , \2370 );
nand \U$1696 ( \2372 , \2081_nGf30 , \1350 );
or \U$1697 ( \2373 , \1310 , \2025_nG100c );
nand \U$1698 ( \2374 , \2373 , \1376 );
and \U$1699 ( \2375 , \2372 , \2374 );
and \U$1700 ( \2376 , \1379 , \2025_nG100c );
and \U$1701 ( \2377 , \2081_nGf30 , \1353 );
nor \U$1702 ( \2378 , \2375 , \2376 , \2377 );
and \U$1703 ( \2379 , \2371 , \2378 );
not \U$1704 ( \2380 , \2379 );
and \U$1705 ( \2381 , RIb557e48_466, \713 );
and \U$1706 ( \2382 , RIb557998_456, \740 );
and \U$1707 ( \2383 , \703 , RIb557bf0_461);
and \U$1708 ( \2384 , RIb557b78_460, \705 );
nor \U$1709 ( \2385 , \2383 , \2384 );
and \U$1710 ( \2386 , \719 , RIb557d58_464);
and \U$1711 ( \2387 , RIb5578a8_454, \734 );
nor \U$1712 ( \2388 , \2386 , \2387 );
and \U$1713 ( \2389 , \1224 , RIb5577b8_452);
and \U$1714 ( \2390 , RIb557830_453, \736 );
nor \U$1715 ( \2391 , \2389 , \2390 );
and \U$1716 ( \2392 , \695 , RIb557ce0_463);
and \U$1717 ( \2393 , RIb557c68_462, \698 );
nor \U$1718 ( \2394 , \2392 , \2393 );
nand \U$1719 ( \2395 , \2385 , \2388 , \2391 , \2394 );
nor \U$1720 ( \2396 , \2381 , \2382 , \2395 );
and \U$1721 ( \2397 , \724 , RIb557a10_457);
and \U$1722 ( \2398 , RIb557a88_458, \726 );
nor \U$1723 ( \2399 , \2397 , \2398 );
and \U$1724 ( \2400 , \710 , RIb557ec0_467);
and \U$1725 ( \2401 , RIb557dd0_465, \716 );
nor \U$1726 ( \2402 , \2400 , \2401 );
and \U$1727 ( \2403 , \690 , RIb557b00_459);
and \U$1728 ( \2404 , RIb557920_455, \738 );
nor \U$1729 ( \2405 , \2403 , \2404 );
nand \U$1730 ( \2406 , \2396 , \2399 , \2402 , \2405 );
_DC gcdf ( \2407_nGcdf , \2406 , \1243 );
nand \U$1731 ( \2408 , \2407_nGcdf , \1214 );
not \U$1732 ( \2409 , \2408 );
and \U$1733 ( \2410 , \2380 , \2409 );
nor \U$1734 ( \2411 , \2371 , \2378 );
nor \U$1735 ( \2412 , \2410 , \2411 );
nand \U$1736 ( \2413 , \2337 , \2412 );
or \U$1737 ( \2414 , \1964 , \1290_nG191a );
or \U$1738 ( \2415 , \1173 , \1172_nG95c );
nand \U$1739 ( \2416 , \2415 , \1174 );
nor \U$1740 ( \2417 , \1964 , \2416 );
not \U$1741 ( \2418 , \2417 );
nand \U$1742 ( \2419 , \1965 , \2418 );
nand \U$1743 ( \2420 , \2414 , \2419 );
or \U$1744 ( \2421 , \2099 , \1339 );
or \U$1745 ( \2422 , \1245 , \2200 );
or \U$1746 ( \2423 , \2101 , \1339 );
or \U$1747 ( \2424 , \1970 , \1244_nG1807 );
nand \U$1748 ( \2425 , \2424 , \2197 );
nand \U$1749 ( \2426 , \2423 , \2425 );
nand \U$1750 ( \2427 , \2421 , \2422 , \2426 );
and \U$1751 ( \2428 , \2420 , \2427 );
and \U$1752 ( \2429 , \2413 , \2428 );
nor \U$1753 ( \2430 , \2412 , \2337 );
nor \U$1754 ( \2431 , \2429 , \2430 );
nand \U$1755 ( \2432 , \2365_nGda9 , \1214 );
and \U$1756 ( \2433 , \2081_nGf30 , \1383 );
or \U$1757 ( \2434 , \1257 , \2252_nGe5c );
nand \U$1758 ( \2435 , \2434 , \1294 );
nand \U$1759 ( \2436 , \2081_nGf30 , \1261 );
and \U$1760 ( \2437 , \2435 , \2436 );
and \U$1761 ( \2438 , \2252_nGe5c , \1416 );
nor \U$1762 ( \2439 , \2433 , \2437 , \2438 );
xnor \U$1763 ( \2440 , \2432 , \2439 );
xor \U$1764 ( \2441 , \2431 , \2440 );
xor \U$1765 ( \2442 , \2122 , \2129 );
xor \U$1766 ( \2443 , \2442 , \2137 );
xor \U$1767 ( \2444 , \2222 , \2261 );
xor \U$1768 ( \2445 , \2443 , \2444 );
and \U$1769 ( \2446 , \2441 , \2445 );
and \U$1770 ( \2447 , \2431 , \2440 );
or \U$1771 ( \2448 , \2446 , \2447 );
nor \U$1772 ( \2449 , \2312 , \2448 );
nor \U$1773 ( \2450 , \2309 , \2449 );
not \U$1774 ( \2451 , \2090 );
not \U$1775 ( \2452 , \2141 );
and \U$1776 ( \2453 , \2451 , \2452 );
and \U$1777 ( \2454 , \2090 , \2141 );
nor \U$1778 ( \2455 , \2453 , \2454 );
nor \U$1779 ( \2456 , \2450 , \2455 );
and \U$1780 ( \2457 , \2450 , \2455 );
or \U$1781 ( \2458 , \2456 , \2457 );
not \U$1782 ( \2459 , \2458 );
not \U$1783 ( \2460 , \2283 );
nor \U$1784 ( \2461 , \2460 , \2269 );
not \U$1785 ( \2462 , \2461 );
not \U$1786 ( \2463 , \2281 );
and \U$1787 ( \2464 , \2462 , \2463 );
and \U$1788 ( \2465 , \2461 , \2281 );
nor \U$1789 ( \2466 , \2464 , \2465 );
not \U$1790 ( \2467 , \2466 );
and \U$1791 ( \2468 , \2459 , \2467 );
and \U$1792 ( \2469 , \2458 , \2466 );
nor \U$1793 ( \2470 , \2468 , \2469 );
not \U$1794 ( \2471 , \2216 );
or \U$1795 ( \2472 , \2194 , \2471 );
not \U$1796 ( \2473 , \2194 );
or \U$1797 ( \2474 , \2216 , \2473 );
or \U$1798 ( \2475 , \2432 , \2439 );
nand \U$1799 ( \2476 , \2472 , \2474 , \2475 );
xor \U$1800 ( \2477 , \2431 , \2440 );
xor \U$1801 ( \2478 , \2477 , \2445 );
not \U$1802 ( \2479 , \2478 );
and \U$1803 ( \2480 , \2476 , \2479 );
not \U$1804 ( \2481 , \1964 );
not \U$1805 ( \2482 , \2215 );
nand \U$1806 ( \2483 , \2482 , \2213 );
not \U$1807 ( \2484 , \2483 );
or \U$1808 ( \2485 , \2481 , \2484 );
or \U$1809 ( \2486 , \2483 , \1964 );
nand \U$1810 ( \2487 , \2485 , \2486 );
xor \U$1811 ( \2488 , \2440 , \2487 );
not \U$1812 ( \2489 , \2428 );
not \U$1813 ( \2490 , \2430 );
nand \U$1814 ( \2491 , \2490 , \2413 );
not \U$1815 ( \2492 , \2491 );
or \U$1816 ( \2493 , \2489 , \2492 );
or \U$1817 ( \2494 , \2491 , \2428 );
nand \U$1818 ( \2495 , \2493 , \2494 );
and \U$1819 ( \2496 , \2488 , \2495 );
and \U$1820 ( \2497 , \2440 , \2487 );
or \U$1821 ( \2498 , \2496 , \2497 );
not \U$1822 ( \2499 , \2498 );
nand \U$1823 ( \2500 , \1789_nG1116 , \1543 );
or \U$1824 ( \2501 , \1425 , \2025_nG100c );
nand \U$1825 ( \2502 , \2501 , \1549 );
and \U$1826 ( \2503 , \2500 , \2502 );
and \U$1827 ( \2504 , \1545 , \2025_nG100c );
and \U$1828 ( \2505 , \1789_nG1116 , \1591 );
nor \U$1829 ( \2506 , \2503 , \2504 , \2505 );
and \U$1830 ( \2507 , \1707_nG11f7 , \1650 );
nand \U$1831 ( \2508 , \1707_nG11f7 , \1647 );
or \U$1832 ( \2509 , \1576 , \1628_nG1300 );
nand \U$1833 ( \2510 , \2509 , \1798 );
and \U$1834 ( \2511 , \2508 , \2510 );
and \U$1835 ( \2512 , \1628_nG1300 , \1801 );
nor \U$1836 ( \2513 , \2507 , \2511 , \2512 );
xor \U$1837 ( \2514 , \2506 , \2513 );
nand \U$1838 ( \2515 , \2252_nGe5c , \1350 );
or \U$1839 ( \2516 , \1310 , \2081_nGf30 );
nand \U$1840 ( \2517 , \2516 , \1376 );
and \U$1841 ( \2518 , \2515 , \2517 );
and \U$1842 ( \2519 , \1379 , \2081_nGf30 );
and \U$1843 ( \2520 , \2252_nGe5c , \1353 );
nor \U$1844 ( \2521 , \2518 , \2519 , \2520 );
and \U$1845 ( \2522 , \2514 , \2521 );
and \U$1846 ( \2523 , \2506 , \2513 );
or \U$1847 ( \2524 , \2522 , \2523 );
nand \U$1848 ( \2525 , \1411_nG15f9 , \2098 );
or \U$1849 ( \2526 , \1970 , \1338_nG1711 );
nand \U$1850 ( \2527 , \2526 , \2197 );
and \U$1851 ( \2528 , \2525 , \2527 );
and \U$1852 ( \2529 , \2201 , \1338_nG1711 );
and \U$1853 ( \2530 , \1411_nG15f9 , \2203 );
nor \U$1854 ( \2531 , \2528 , \2529 , \2530 );
not \U$1855 ( \2532 , \2419 );
and \U$1856 ( \2533 , \1291 , \2532 );
and \U$1857 ( \2534 , \2417 , \1245 );
nand \U$1858 ( \2535 , \2416 , \1964 );
not \U$1859 ( \2536 , \2535 );
and \U$1860 ( \2537 , \1290_nG191a , \2536 );
nor \U$1861 ( \2538 , \2533 , \2534 , \2537 );
xor \U$1862 ( \2539 , \2531 , \2538 );
nand \U$1863 ( \2540 , \1538_nG13f2 , \1864 );
or \U$1864 ( \2541 , \1810 , \1493_nG14ed );
nand \U$1865 ( \2542 , \2541 , \1959 );
and \U$1866 ( \2543 , \2540 , \2542 );
and \U$1867 ( \2544 , \1954 , \1493_nG14ed );
and \U$1868 ( \2545 , \1538_nG13f2 , \1866 );
nor \U$1869 ( \2546 , \2543 , \2544 , \2545 );
and \U$1870 ( \2547 , \2539 , \2546 );
and \U$1871 ( \2548 , \2531 , \2538 );
or \U$1872 ( \2549 , \2547 , \2548 );
nor \U$1873 ( \2550 , \2524 , \2549 );
xor \U$1874 ( \2551 , \2176 , \2183 );
xor \U$1875 ( \2552 , \2551 , \2191 );
not \U$1876 ( \2553 , \2552 );
and \U$1877 ( \2554 , \2550 , \2553 );
not \U$1878 ( \2555 , \2550 );
nand \U$1879 ( \2556 , \2555 , \2552 );
xor \U$1880 ( \2557 , \2319 , \2326 );
xor \U$1881 ( \2558 , \2557 , \2334 );
not \U$1882 ( \2559 , \2558 );
not \U$1883 ( \2560 , \2408 );
nor \U$1884 ( \2561 , \2379 , \2411 );
not \U$1885 ( \2562 , \2561 );
or \U$1886 ( \2563 , \2560 , \2562 );
or \U$1887 ( \2564 , \2561 , \2408 );
nand \U$1888 ( \2565 , \2563 , \2564 );
and \U$1889 ( \2566 , \2559 , \2565 );
and \U$1890 ( \2567 , \2556 , \2566 );
nor \U$1891 ( \2568 , \2554 , \2567 );
nand \U$1892 ( \2569 , \2499 , \2568 );
xor \U$1893 ( \2570 , \2480 , \2569 );
not \U$1894 ( \2571 , \2307 );
not \U$1895 ( \2572 , \2448 );
not \U$1896 ( \2573 , \2308 );
and \U$1897 ( \2574 , \2572 , \2573 );
and \U$1898 ( \2575 , \2448 , \2308 );
nor \U$1899 ( \2576 , \2574 , \2575 );
not \U$1900 ( \2577 , \2576 );
or \U$1901 ( \2578 , \2571 , \2577 );
or \U$1902 ( \2579 , \2576 , \2307 );
nand \U$1903 ( \2580 , \2578 , \2579 );
and \U$1904 ( \2581 , \2570 , \2580 );
and \U$1905 ( \2582 , \2480 , \2569 );
or \U$1906 ( \2583 , \2581 , \2582 );
xor \U$1907 ( \2584 , \2470 , \2583 );
xor \U$1908 ( \2585 , \2476 , \2479 );
not \U$1909 ( \2586 , \2498 );
not \U$1910 ( \2587 , \2568 );
and \U$1911 ( \2588 , \2586 , \2587 );
and \U$1912 ( \2589 , \2498 , \2568 );
nor \U$1913 ( \2590 , \2588 , \2589 );
xor \U$1914 ( \2591 , \2585 , \2590 );
xor \U$1915 ( \2592 , \2506 , \2513 );
xor \U$1916 ( \2593 , \2592 , \2521 );
not \U$1917 ( \2594 , \2593 );
and \U$1918 ( \2595 , RIb559018_504, \736 );
and \U$1919 ( \2596 , RIb559450_513, \698 );
and \U$1920 ( \2597 , \724 , RIb5591f8_508);
and \U$1921 ( \2598 , RIb559180_507, \740 );
nor \U$1922 ( \2599 , \2597 , \2598 );
and \U$1923 ( \2600 , \710 , RIb5596a8_518);
and \U$1924 ( \2601 , RIb5592e8_510, \690 );
nor \U$1925 ( \2602 , \2600 , \2601 );
and \U$1926 ( \2603 , \713 , RIb559630_517);
and \U$1927 ( \2604 , RIb559270_509, \726 );
nor \U$1928 ( \2605 , \2603 , \2604 );
and \U$1929 ( \2606 , \703 , RIb5593d8_512);
and \U$1930 ( \2607 , RIb559360_511, \705 );
nor \U$1931 ( \2608 , \2606 , \2607 );
nand \U$1932 ( \2609 , \2599 , \2602 , \2605 , \2608 );
nor \U$1933 ( \2610 , \2595 , \2596 , \2609 );
and \U$1934 ( \2611 , \716 , RIb5595b8_516);
and \U$1935 ( \2612 , RIb559090_505, \734 );
nor \U$1936 ( \2613 , \2611 , \2612 );
and \U$1937 ( \2614 , \695 , RIb5594c8_514);
and \U$1938 ( \2615 , RIb559540_515, \719 );
nor \U$1939 ( \2616 , \2614 , \2615 );
and \U$1940 ( \2617 , \1224 , RIb558fa0_503);
and \U$1941 ( \2618 , RIb559108_506, \738 );
nor \U$1942 ( \2619 , \2617 , \2618 );
nand \U$1943 ( \2620 , \2610 , \2613 , \2616 , \2619 );
_DC gc52 ( \2621_nGc52 , \2620 , \1243 );
nand \U$1944 ( \2622 , \2621_nGc52 , \1214 );
and \U$1945 ( \2623 , \2365_nGda9 , \1383 );
or \U$1946 ( \2624 , \1257 , \2407_nGcdf );
nand \U$1947 ( \2625 , \2624 , \1294 );
nand \U$1948 ( \2626 , \2365_nGda9 , \1261 );
and \U$1949 ( \2627 , \2625 , \2626 );
and \U$1950 ( \2628 , \2407_nGcdf , \1416 );
nor \U$1951 ( \2629 , \2623 , \2627 , \2628 );
xor \U$1952 ( \2630 , \2622 , \2629 );
and \U$1953 ( \2631 , \2594 , \2630 );
xor \U$1954 ( \2632 , \2420 , \2427 );
xor \U$1955 ( \2633 , \2631 , \2632 );
and \U$1956 ( \2634 , \1789_nG1116 , \1650 );
nand \U$1957 ( \2635 , \1789_nG1116 , \1647 );
or \U$1958 ( \2636 , \1576 , \1707_nG11f7 );
nand \U$1959 ( \2637 , \2636 , \1798 );
and \U$1960 ( \2638 , \2635 , \2637 );
and \U$1961 ( \2639 , \1707_nG11f7 , \1801 );
nor \U$1962 ( \2640 , \2634 , \2638 , \2639 );
nand \U$1963 ( \2641 , \1628_nG1300 , \1864 );
or \U$1964 ( \2642 , \1810 , \1538_nG13f2 );
nand \U$1965 ( \2643 , \2642 , \1959 );
and \U$1966 ( \2644 , \2641 , \2643 );
and \U$1967 ( \2645 , \1954 , \1538_nG13f2 );
and \U$1968 ( \2646 , \1628_nG1300 , \1866 );
nor \U$1969 ( \2647 , \2644 , \2645 , \2646 );
xor \U$1970 ( \2648 , \2640 , \2647 );
nand \U$1971 ( \2649 , \2025_nG100c , \1543 );
or \U$1972 ( \2650 , \1425 , \2081_nGf30 );
nand \U$1973 ( \2651 , \2650 , \1549 );
and \U$1974 ( \2652 , \2649 , \2651 );
and \U$1975 ( \2653 , \1545 , \2081_nGf30 );
and \U$1976 ( \2654 , \2025_nG100c , \1591 );
nor \U$1977 ( \2655 , \2652 , \2653 , \2654 );
and \U$1978 ( \2656 , \2648 , \2655 );
and \U$1979 ( \2657 , \2640 , \2647 );
or \U$1980 ( \2658 , \2656 , \2657 );
not \U$1981 ( \2659 , \2658 );
or \U$1982 ( \2660 , \2535 , \1245 );
or \U$1983 ( \2661 , \1244_nG1807 , \2419 );
or \U$1984 ( \2662 , \1338_nG1711 , \2418 );
nand \U$1985 ( \2663 , \2660 , \2661 , \2662 );
or \U$1986 ( \2664 , \2099 , \1494 );
or \U$1987 ( \2665 , \1972 , \2200 );
or \U$1988 ( \2666 , \2101 , \1494 );
or \U$1989 ( \2667 , \1970 , \1411_nG15f9 );
nand \U$1990 ( \2668 , \2667 , \2197 );
nand \U$1991 ( \2669 , \2666 , \2668 );
nand \U$1992 ( \2670 , \2664 , \2665 , \2669 );
and \U$1993 ( \2671 , \2663 , \2670 );
xor \U$1994 ( \2672 , \2659 , \2671 );
not \U$1995 ( \2673 , \2365_nGda9 );
or \U$1996 ( \2674 , \1354 , \2673 );
or \U$1997 ( \2675 , \1310 , \2252_nGe5c );
nand \U$1998 ( \2676 , \2675 , \1376 );
nand \U$1999 ( \2677 , \2365_nGda9 , \1350 );
and \U$2000 ( \2678 , \2676 , \2677 );
and \U$2001 ( \2679 , \2252_nGe5c , \1379 );
nor \U$2002 ( \2680 , \2678 , \2679 );
nand \U$2003 ( \2681 , \2674 , \2680 );
and \U$2004 ( \2682 , RIb558a00_491, \724 );
and \U$2005 ( \2683 , RIb558a78_492, \726 );
and \U$2006 ( \2684 , \703 , RIb558be0_495);
and \U$2007 ( \2685 , RIb558c58_496, \698 );
nor \U$2008 ( \2686 , \2684 , \2685 );
and \U$2009 ( \2687 , \738 , RIb558910_489);
and \U$2010 ( \2688 , RIb558898_488, \734 );
nor \U$2011 ( \2689 , \2687 , \2688 );
and \U$2012 ( \2690 , \1224 , RIb5587a8_486);
and \U$2013 ( \2691 , RIb558820_487, \736 );
nor \U$2014 ( \2692 , \2690 , \2691 );
and \U$2015 ( \2693 , \695 , RIb558cd0_497);
and \U$2016 ( \2694 , RIb558d48_498, \719 );
nor \U$2017 ( \2695 , \2693 , \2694 );
nand \U$2018 ( \2696 , \2686 , \2689 , \2692 , \2695 );
nor \U$2019 ( \2697 , \2682 , \2683 , \2696 );
and \U$2020 ( \2698 , \716 , RIb558dc0_499);
and \U$2021 ( \2699 , RIb558e38_500, \713 );
nor \U$2022 ( \2700 , \2698 , \2699 );
and \U$2023 ( \2701 , \710 , RIb558eb0_501);
and \U$2024 ( \2702 , RIb558988_490, \740 );
nor \U$2025 ( \2703 , \2701 , \2702 );
and \U$2026 ( \2704 , \690 , RIb558af0_493);
and \U$2027 ( \2705 , RIb558b68_494, \705 );
nor \U$2028 ( \2706 , \2704 , \2705 );
nand \U$2029 ( \2707 , \2697 , \2700 , \2703 , \2706 );
_DC gbb2 ( \2708_nGbb2 , \2707 , \1243 );
not \U$2030 ( \2709 , \2708_nGbb2 );
nor \U$2031 ( \2710 , \1215 , \2709 );
xor \U$2032 ( \2711 , \2681 , \2710 );
not \U$2033 ( \2712 , \2407_nGcdf );
or \U$2034 ( \2713 , \1297 , \2712 );
not \U$2035 ( \2714 , \2621_nGc52 );
or \U$2036 ( \2715 , \2714 , \1263 );
or \U$2037 ( \2716 , \1260 , \2712 );
or \U$2038 ( \2717 , \1257 , \2621_nGc52 );
nand \U$2039 ( \2718 , \2717 , \1294 );
nand \U$2040 ( \2719 , \2716 , \2718 );
nand \U$2041 ( \2720 , \2713 , \2715 , \2719 );
and \U$2042 ( \2721 , \2711 , \2720 );
and \U$2043 ( \2722 , \2681 , \2710 );
or \U$2044 ( \2723 , \2721 , \2722 );
and \U$2045 ( \2724 , \2672 , \2723 );
and \U$2046 ( \2725 , \2659 , \2671 );
or \U$2047 ( \2726 , \2724 , \2725 );
and \U$2048 ( \2727 , \2633 , \2726 );
and \U$2049 ( \2728 , \2631 , \2632 );
or \U$2050 ( \2729 , \2727 , \2728 );
not \U$2051 ( \2730 , \2524 );
or \U$2052 ( \2731 , \2730 , \2549 );
not \U$2053 ( \2732 , \2549 );
or \U$2054 ( \2733 , \2732 , \2524 );
or \U$2055 ( \2734 , \2622 , \2629 );
nand \U$2056 ( \2735 , \2731 , \2733 , \2734 );
xor \U$2057 ( \2736 , \2559 , \2565 );
and \U$2058 ( \2737 , \2735 , \2736 );
xor \U$2059 ( \2738 , \2729 , \2737 );
xor \U$2060 ( \2739 , \2440 , \2487 );
xor \U$2061 ( \2740 , \2739 , \2495 );
and \U$2062 ( \2741 , \2738 , \2740 );
and \U$2063 ( \2742 , \2729 , \2737 );
or \U$2064 ( \2743 , \2741 , \2742 );
and \U$2065 ( \2744 , \2591 , \2743 );
and \U$2066 ( \2745 , \2585 , \2590 );
or \U$2067 ( \2746 , \2744 , \2745 );
xor \U$2068 ( \2747 , \2480 , \2569 );
xor \U$2069 ( \2748 , \2747 , \2580 );
xor \U$2070 ( \2749 , \2746 , \2748 );
xor \U$2071 ( \2750 , \2735 , \2736 );
xor \U$2072 ( \2751 , \2531 , \2538 );
xor \U$2073 ( \2752 , \2751 , \2546 );
not \U$2074 ( \2753 , \2752 );
nand \U$2075 ( \2754 , \2081_nGf30 , \1543 );
or \U$2076 ( \2755 , \1425 , \2252_nGe5c );
nand \U$2077 ( \2756 , \2755 , \1549 );
and \U$2078 ( \2757 , \2754 , \2756 );
and \U$2079 ( \2758 , \1545 , \2252_nGe5c );
and \U$2080 ( \2759 , \2081_nGf30 , \1591 );
nor \U$2081 ( \2760 , \2757 , \2758 , \2759 );
and \U$2082 ( \2761 , \2025_nG100c , \1650 );
nand \U$2083 ( \2762 , \2025_nG100c , \1647 );
or \U$2084 ( \2763 , \1576 , \1789_nG1116 );
nand \U$2085 ( \2764 , \2763 , \1798 );
and \U$2086 ( \2765 , \2762 , \2764 );
and \U$2087 ( \2766 , \1789_nG1116 , \1801 );
nor \U$2088 ( \2767 , \2761 , \2765 , \2766 );
xor \U$2089 ( \2768 , \2760 , \2767 );
nand \U$2090 ( \2769 , \2407_nGcdf , \1350 );
or \U$2091 ( \2770 , \1310 , \2365_nGda9 );
nand \U$2092 ( \2771 , \2770 , \1376 );
and \U$2093 ( \2772 , \2769 , \2771 );
and \U$2094 ( \2773 , \1379 , \2365_nGda9 );
and \U$2095 ( \2774 , \2407_nGcdf , \1353 );
nor \U$2096 ( \2775 , \2772 , \2773 , \2774 );
and \U$2097 ( \2776 , \2768 , \2775 );
and \U$2098 ( \2777 , \2760 , \2767 );
or \U$2099 ( \2778 , \2776 , \2777 );
nand \U$2100 ( \2779 , \1538_nG13f2 , \2098 );
or \U$2101 ( \2780 , \1970 , \1493_nG14ed );
nand \U$2102 ( \2781 , \2780 , \2197 );
and \U$2103 ( \2782 , \2779 , \2781 );
and \U$2104 ( \2783 , \2201 , \1493_nG14ed );
and \U$2105 ( \2784 , \1538_nG13f2 , \2203 );
nor \U$2106 ( \2785 , \2782 , \2783 , \2784 );
and \U$2107 ( \2786 , \1339 , \2532 );
and \U$2108 ( \2787 , \2417 , \1972 );
and \U$2109 ( \2788 , \1338_nG1711 , \2536 );
nor \U$2110 ( \2789 , \2786 , \2787 , \2788 );
xor \U$2111 ( \2790 , \2785 , \2789 );
nand \U$2112 ( \2791 , \1707_nG11f7 , \1864 );
or \U$2113 ( \2792 , \1810 , \1628_nG1300 );
nand \U$2114 ( \2793 , \2792 , \1959 );
and \U$2115 ( \2794 , \2791 , \2793 );
and \U$2116 ( \2795 , \1954 , \1628_nG1300 );
and \U$2117 ( \2796 , \1707_nG11f7 , \1866 );
nor \U$2118 ( \2797 , \2794 , \2795 , \2796 );
and \U$2119 ( \2798 , \2790 , \2797 );
and \U$2120 ( \2799 , \2785 , \2789 );
or \U$2121 ( \2800 , \2798 , \2799 );
nor \U$2122 ( \2801 , \2778 , \2800 );
and \U$2123 ( \2802 , \2753 , \2801 );
xor \U$2124 ( \2803 , \2750 , \2802 );
xor \U$2125 ( \2804 , \2631 , \2632 );
xor \U$2126 ( \2805 , \2804 , \2726 );
and \U$2127 ( \2806 , \2803 , \2805 );
and \U$2128 ( \2807 , \2750 , \2802 );
or \U$2129 ( \2808 , \2806 , \2807 );
not \U$2130 ( \2809 , \2552 );
xor \U$2131 ( \2810 , \2550 , \2566 );
not \U$2132 ( \2811 , \2810 );
or \U$2133 ( \2812 , \2809 , \2811 );
or \U$2134 ( \2813 , \2810 , \2552 );
nand \U$2135 ( \2814 , \2812 , \2813 );
xor \U$2136 ( \2815 , \2808 , \2814 );
xor \U$2137 ( \2816 , \2729 , \2737 );
xor \U$2138 ( \2817 , \2816 , \2740 );
and \U$2139 ( \2818 , \2815 , \2817 );
and \U$2140 ( \2819 , \2808 , \2814 );
or \U$2141 ( \2820 , \2818 , \2819 );
xor \U$2142 ( \2821 , \2585 , \2590 );
xor \U$2143 ( \2822 , \2821 , \2743 );
xor \U$2144 ( \2823 , \2820 , \2822 );
xor \U$2145 ( \2824 , \2808 , \2814 );
xor \U$2146 ( \2825 , \2824 , \2817 );
not \U$2147 ( \2826 , \2778 );
or \U$2148 ( \2827 , \2826 , \2800 );
not \U$2149 ( \2828 , \2800 );
or \U$2150 ( \2829 , \2828 , \2778 );
and \U$2151 ( \2830 , RIb55a1e8_542, \724 );
and \U$2152 ( \2831 , RIb55a2d8_544, \690 );
and \U$2153 ( \2832 , \738 , RIb55a0f8_540);
and \U$2154 ( \2833 , RIb55a080_539, \734 );
nor \U$2155 ( \2834 , \2832 , \2833 );
and \U$2156 ( \2835 , \695 , RIb55a4b8_548);
and \U$2157 ( \2836 , RIb55a440_547, \698 );
nor \U$2158 ( \2837 , \2835 , \2836 );
and \U$2159 ( \2838 , \1224 , RIb559f90_537);
and \U$2160 ( \2839 , RIb55a008_538, \736 );
nor \U$2161 ( \2840 , \2838 , \2839 );
and \U$2162 ( \2841 , \716 , RIb55a5a8_550);
and \U$2163 ( \2842 , RIb55a530_549, \719 );
nor \U$2164 ( \2843 , \2841 , \2842 );
nand \U$2165 ( \2844 , \2834 , \2837 , \2840 , \2843 );
nor \U$2166 ( \2845 , \2830 , \2831 , \2844 );
and \U$2167 ( \2846 , \710 , RIb55a698_552);
and \U$2168 ( \2847 , RIb55a260_543, \726 );
nor \U$2169 ( \2848 , \2846 , \2847 );
and \U$2170 ( \2849 , \713 , RIb55a620_551);
and \U$2171 ( \2850 , RIb55a170_541, \740 );
nor \U$2172 ( \2851 , \2849 , \2850 );
and \U$2173 ( \2852 , \703 , RIb55a3c8_546);
and \U$2174 ( \2853 , RIb55a350_545, \705 );
nor \U$2175 ( \2854 , \2852 , \2853 );
nand \U$2176 ( \2855 , \2845 , \2848 , \2851 , \2854 );
_DC gb3b ( \2856_nGb3b , \2855 , \1243 );
nand \U$2177 ( \2857 , \2856_nGb3b , \1214 );
and \U$2178 ( \2858 , \2621_nGc52 , \1383 );
or \U$2179 ( \2859 , \1257 , \2708_nGbb2 );
nand \U$2180 ( \2860 , \2859 , \1294 );
nand \U$2181 ( \2861 , \2621_nGc52 , \1261 );
and \U$2182 ( \2862 , \2860 , \2861 );
and \U$2183 ( \2863 , \2708_nGbb2 , \1416 );
nor \U$2184 ( \2864 , \2858 , \2862 , \2863 );
or \U$2185 ( \2865 , \2857 , \2864 );
nand \U$2186 ( \2866 , \2827 , \2829 , \2865 );
xor \U$2187 ( \2867 , \2663 , \2670 );
xor \U$2188 ( \2868 , \2866 , \2867 );
xor \U$2189 ( \2869 , \2681 , \2710 );
xor \U$2190 ( \2870 , \2869 , \2720 );
and \U$2191 ( \2871 , \2868 , \2870 );
and \U$2192 ( \2872 , \2866 , \2867 );
or \U$2193 ( \2873 , \2871 , \2872 );
xor \U$2194 ( \2874 , \2594 , \2630 );
xor \U$2195 ( \2875 , \2873 , \2874 );
xor \U$2196 ( \2876 , \2760 , \2767 );
xor \U$2197 ( \2877 , \2876 , \2775 );
xor \U$2198 ( \2878 , \2785 , \2789 );
xor \U$2199 ( \2879 , \2878 , \2797 );
xor \U$2200 ( \2880 , \2877 , \2879 );
xnor \U$2201 ( \2881 , \2857 , \2864 );
and \U$2202 ( \2882 , \2880 , \2881 );
and \U$2203 ( \2883 , \2877 , \2879 );
or \U$2204 ( \2884 , \2882 , \2883 );
xor \U$2205 ( \2885 , \2640 , \2647 );
xor \U$2206 ( \2886 , \2885 , \2655 );
xor \U$2207 ( \2887 , \2884 , \2886 );
and \U$2208 ( \2888 , \2081_nGf30 , \1650 );
nand \U$2209 ( \2889 , \2081_nGf30 , \1647 );
or \U$2210 ( \2890 , \1576 , \2025_nG100c );
nand \U$2211 ( \2891 , \2890 , \1798 );
and \U$2212 ( \2892 , \2889 , \2891 );
and \U$2213 ( \2893 , \2025_nG100c , \1801 );
nor \U$2214 ( \2894 , \2888 , \2892 , \2893 );
nand \U$2215 ( \2895 , \1789_nG1116 , \1864 );
or \U$2216 ( \2896 , \1810 , \1707_nG11f7 );
nand \U$2217 ( \2897 , \2896 , \1959 );
and \U$2218 ( \2898 , \2895 , \2897 );
and \U$2219 ( \2899 , \1954 , \1707_nG11f7 );
and \U$2220 ( \2900 , \1789_nG1116 , \1866 );
nor \U$2221 ( \2901 , \2898 , \2899 , \2900 );
xor \U$2222 ( \2902 , \2894 , \2901 );
nand \U$2223 ( \2903 , \2252_nGe5c , \1543 );
or \U$2224 ( \2904 , \1425 , \2365_nGda9 );
nand \U$2225 ( \2905 , \2904 , \1549 );
and \U$2226 ( \2906 , \2903 , \2905 );
and \U$2227 ( \2907 , \1545 , \2365_nGda9 );
and \U$2228 ( \2908 , \2252_nGe5c , \1591 );
nor \U$2229 ( \2909 , \2906 , \2907 , \2908 );
and \U$2230 ( \2910 , \2902 , \2909 );
and \U$2231 ( \2911 , \2894 , \2901 );
or \U$2232 ( \2912 , \2910 , \2911 );
nand \U$2233 ( \2913 , \1628_nG1300 , \2098 );
or \U$2234 ( \2914 , \1970 , \1538_nG13f2 );
nand \U$2235 ( \2915 , \2914 , \2197 );
and \U$2236 ( \2916 , \2913 , \2915 );
and \U$2237 ( \2917 , \2201 , \1538_nG13f2 );
and \U$2238 ( \2918 , \1628_nG1300 , \2203 );
nor \U$2239 ( \2919 , \2916 , \2917 , \2918 );
not \U$2240 ( \2920 , \2919 );
or \U$2241 ( \2921 , \2535 , \1972 );
or \U$2242 ( \2922 , \1411_nG15f9 , \2419 );
or \U$2243 ( \2923 , \1493_nG14ed , \2418 );
nand \U$2244 ( \2924 , \2921 , \2922 , \2923 );
nand \U$2245 ( \2925 , \2920 , \2924 );
xor \U$2246 ( \2926 , \2912 , \2925 );
and \U$2247 ( \2927 , \2708_nGbb2 , \1383 );
or \U$2248 ( \2928 , \1257 , \2856_nGb3b );
nand \U$2249 ( \2929 , \2928 , \1294 );
nand \U$2250 ( \2930 , \2708_nGbb2 , \1261 );
and \U$2251 ( \2931 , \2929 , \2930 );
and \U$2252 ( \2932 , \2856_nGb3b , \1416 );
nor \U$2253 ( \2933 , \2927 , \2931 , \2932 );
nand \U$2254 ( \2934 , \2621_nGc52 , \1350 );
or \U$2255 ( \2935 , \1310 , \2407_nGcdf );
nand \U$2256 ( \2936 , \2935 , \1376 );
and \U$2257 ( \2937 , \2934 , \2936 );
and \U$2258 ( \2938 , \1379 , \2407_nGcdf );
and \U$2259 ( \2939 , \2621_nGc52 , \1353 );
nor \U$2260 ( \2940 , \2937 , \2938 , \2939 );
and \U$2261 ( \2941 , \2933 , \2940 );
not \U$2262 ( \2942 , \2941 );
and \U$2263 ( \2943 , RIb559810_521, \736 );
and \U$2264 ( \2944 , RIb559888_522, \734 );
and \U$2265 ( \2945 , \703 , RIb559bd0_529);
and \U$2266 ( \2946 , RIb559b58_528, \705 );
nor \U$2267 ( \2947 , \2945 , \2946 );
and \U$2268 ( \2948 , \710 , RIb559ea0_535);
and \U$2269 ( \2949 , RIb559ae0_527, \690 );
nor \U$2270 ( \2950 , \2948 , \2949 );
and \U$2271 ( \2951 , \713 , RIb559e28_534);
and \U$2272 ( \2952 , RIb559a68_526, \726 );
nor \U$2273 ( \2953 , \2951 , \2952 );
and \U$2274 ( \2954 , \724 , RIb5599f0_525);
and \U$2275 ( \2955 , RIb559978_524, \740 );
nor \U$2276 ( \2956 , \2954 , \2955 );
nand \U$2277 ( \2957 , \2947 , \2950 , \2953 , \2956 );
nor \U$2278 ( \2958 , \2943 , \2944 , \2957 );
and \U$2279 ( \2959 , \738 , RIb559900_523);
and \U$2280 ( \2960 , RIb559c48_530, \698 );
nor \U$2281 ( \2961 , \2959 , \2960 );
and \U$2282 ( \2962 , \695 , RIb559cc0_531);
and \U$2283 ( \2963 , RIb559d38_532, \719 );
nor \U$2284 ( \2964 , \2962 , \2963 );
and \U$2285 ( \2965 , \1224 , RIb559798_520);
and \U$2286 ( \2966 , RIb559db0_533, \716 );
nor \U$2287 ( \2967 , \2965 , \2966 );
nand \U$2288 ( \2968 , \2958 , \2961 , \2964 , \2967 );
_DC gabe ( \2969_nGabe , \2968 , \1243 );
nand \U$2289 ( \2970 , \2969_nGabe , \1214 );
not \U$2290 ( \2971 , \2970 );
and \U$2291 ( \2972 , \2942 , \2971 );
nor \U$2292 ( \2973 , \2933 , \2940 );
nor \U$2293 ( \2974 , \2972 , \2973 );
and \U$2294 ( \2975 , \2926 , \2974 );
and \U$2295 ( \2976 , \2912 , \2925 );
or \U$2296 ( \2977 , \2975 , \2976 );
and \U$2297 ( \2978 , \2887 , \2977 );
and \U$2298 ( \2979 , \2884 , \2886 );
or \U$2299 ( \2980 , \2978 , \2979 );
not \U$2300 ( \2981 , \2980 );
and \U$2301 ( \2982 , \2875 , \2981 );
and \U$2302 ( \2983 , \2873 , \2874 );
or \U$2303 ( \2984 , \2982 , \2983 );
xor \U$2304 ( \2985 , \2753 , \2801 );
xor \U$2305 ( \2986 , \2659 , \2671 );
xor \U$2306 ( \2987 , \2986 , \2723 );
and \U$2307 ( \2988 , \2985 , \2987 );
xor \U$2308 ( \2989 , \2984 , \2988 );
xor \U$2309 ( \2990 , \2750 , \2802 );
xor \U$2310 ( \2991 , \2990 , \2805 );
and \U$2311 ( \2992 , \2989 , \2991 );
and \U$2312 ( \2993 , \2984 , \2988 );
or \U$2313 ( \2994 , \2992 , \2993 );
xor \U$2314 ( \2995 , \2825 , \2994 );
xor \U$2315 ( \2996 , \2984 , \2988 );
xor \U$2316 ( \2997 , \2996 , \2991 );
xor \U$2317 ( \2998 , \2884 , \2886 );
xor \U$2318 ( \2999 , \2998 , \2977 );
xor \U$2319 ( \3000 , \2877 , \2879 );
xor \U$2320 ( \3001 , \3000 , \2881 );
nand \U$2321 ( \3002 , \2365_nGda9 , \1543 );
or \U$2322 ( \3003 , \1425 , \2407_nGcdf );
nand \U$2323 ( \3004 , \3003 , \1549 );
and \U$2324 ( \3005 , \3002 , \3004 );
and \U$2325 ( \3006 , \1545 , \2407_nGcdf );
and \U$2326 ( \3007 , \2365_nGda9 , \1591 );
nor \U$2327 ( \3008 , \3005 , \3006 , \3007 );
and \U$2328 ( \3009 , \2252_nGe5c , \1650 );
nand \U$2329 ( \3010 , \2252_nGe5c , \1647 );
or \U$2330 ( \3011 , \1576 , \2081_nGf30 );
nand \U$2331 ( \3012 , \3011 , \1798 );
and \U$2332 ( \3013 , \3010 , \3012 );
and \U$2333 ( \3014 , \2081_nGf30 , \1801 );
nor \U$2334 ( \3015 , \3009 , \3013 , \3014 );
xor \U$2335 ( \3016 , \3008 , \3015 );
nand \U$2336 ( \3017 , \2708_nGbb2 , \1350 );
or \U$2337 ( \3018 , \1310 , \2621_nGc52 );
nand \U$2338 ( \3019 , \3018 , \1376 );
and \U$2339 ( \3020 , \3017 , \3019 );
and \U$2340 ( \3021 , \1379 , \2621_nGc52 );
and \U$2341 ( \3022 , \2708_nGbb2 , \1353 );
nor \U$2342 ( \3023 , \3020 , \3021 , \3022 );
and \U$2343 ( \3024 , \3016 , \3023 );
and \U$2344 ( \3025 , \3008 , \3015 );
or \U$2345 ( \3026 , \3024 , \3025 );
nand \U$2346 ( \3027 , \1707_nG11f7 , \2098 );
or \U$2347 ( \3028 , \1970 , \1628_nG1300 );
nand \U$2348 ( \3029 , \3028 , \2197 );
and \U$2349 ( \3030 , \3027 , \3029 );
and \U$2350 ( \3031 , \2201 , \1628_nG1300 );
and \U$2351 ( \3032 , \1707_nG11f7 , \2203 );
nor \U$2352 ( \3033 , \3030 , \3031 , \3032 );
and \U$2353 ( \3034 , \1494 , \2532 );
and \U$2354 ( \3035 , \2417 , \1632 );
and \U$2355 ( \3036 , \1493_nG14ed , \2536 );
nor \U$2356 ( \3037 , \3034 , \3035 , \3036 );
xor \U$2357 ( \3038 , \3033 , \3037 );
nand \U$2358 ( \3039 , \2025_nG100c , \1864 );
or \U$2359 ( \3040 , \1810 , \1789_nG1116 );
nand \U$2360 ( \3041 , \3040 , \1959 );
and \U$2361 ( \3042 , \3039 , \3041 );
and \U$2362 ( \3043 , \1954 , \1789_nG1116 );
and \U$2363 ( \3044 , \2025_nG100c , \1866 );
nor \U$2364 ( \3045 , \3042 , \3043 , \3044 );
and \U$2365 ( \3046 , \3038 , \3045 );
and \U$2366 ( \3047 , \3033 , \3037 );
or \U$2367 ( \3048 , \3046 , \3047 );
nor \U$2368 ( \3049 , \3026 , \3048 );
not \U$2369 ( \3050 , \3049 );
or \U$2370 ( \3051 , \3001 , \3050 );
xor \U$2371 ( \3052 , \2894 , \2901 );
xor \U$2372 ( \3053 , \3052 , \2909 );
not \U$2373 ( \3054 , \3053 );
not \U$2374 ( \3055 , \2970 );
nor \U$2375 ( \3056 , \2941 , \2973 );
not \U$2376 ( \3057 , \3056 );
or \U$2377 ( \3058 , \3055 , \3057 );
or \U$2378 ( \3059 , \3056 , \2970 );
nand \U$2379 ( \3060 , \3058 , \3059 );
nand \U$2380 ( \3061 , \3054 , \3060 );
and \U$2381 ( \3062 , \3001 , \3050 );
or \U$2382 ( \3063 , \3061 , \3062 );
nand \U$2383 ( \3064 , \3051 , \3063 );
xor \U$2384 ( \3065 , \2866 , \2867 );
xor \U$2385 ( \3066 , \3065 , \2870 );
nor \U$2386 ( \3067 , \3064 , \3066 );
or \U$2387 ( \3068 , \2999 , \3067 );
nand \U$2388 ( \3069 , \3066 , \3064 );
nand \U$2389 ( \3070 , \3068 , \3069 );
xor \U$2390 ( \3071 , \2985 , \2987 );
xor \U$2391 ( \3072 , \3070 , \3071 );
xor \U$2392 ( \3073 , \2873 , \2874 );
xor \U$2393 ( \3074 , \3073 , \2981 );
and \U$2394 ( \3075 , \3072 , \3074 );
and \U$2395 ( \3076 , \3070 , \3071 );
or \U$2396 ( \3077 , \3075 , \3076 );
xor \U$2397 ( \3078 , \2997 , \3077 );
xor \U$2398 ( \3079 , \3070 , \3071 );
xor \U$2399 ( \3080 , \3079 , \3074 );
not \U$2400 ( \3081 , \3069 );
nor \U$2401 ( \3082 , \3081 , \3067 );
not \U$2402 ( \3083 , \3082 );
not \U$2403 ( \3084 , \2999 );
and \U$2404 ( \3085 , \3083 , \3084 );
and \U$2405 ( \3086 , \3082 , \2999 );
nor \U$2406 ( \3087 , \3085 , \3086 );
not \U$2407 ( \3088 , \3060 );
not \U$2408 ( \3089 , \3053 );
and \U$2409 ( \3090 , \3088 , \3089 );
and \U$2410 ( \3091 , \3060 , \3053 );
nor \U$2411 ( \3092 , \3090 , \3091 );
not \U$2412 ( \3093 , \3092 );
not \U$2413 ( \3094 , \3048 );
or \U$2414 ( \3095 , \3026 , \3094 );
not \U$2415 ( \3096 , \3026 );
or \U$2416 ( \3097 , \3048 , \3096 );
and \U$2417 ( \3098 , RIb55a968_558, \740 );
and \U$2418 ( \3099 , RIb55ae90_569, \710 );
and \U$2419 ( \3100 , \738 , RIb55a8f0_557);
and \U$2420 ( \3101 , RIb55a878_556, \734 );
nor \U$2421 ( \3102 , \3100 , \3101 );
and \U$2422 ( \3103 , \716 , RIb55ada0_567);
and \U$2423 ( \3104 , RIb55ad28_566, \719 );
nor \U$2424 ( \3105 , \3103 , \3104 );
and \U$2425 ( \3106 , \1224 , RIb55a788_554);
and \U$2426 ( \3107 , RIb55a800_555, \736 );
nor \U$2427 ( \3108 , \3106 , \3107 );
and \U$2428 ( \3109 , \695 , RIb55acb0_565);
and \U$2429 ( \3110 , RIb55ac38_564, \698 );
nor \U$2430 ( \3111 , \3109 , \3110 );
nand \U$2431 ( \3112 , \3102 , \3105 , \3108 , \3111 );
nor \U$2432 ( \3113 , \3098 , \3099 , \3112 );
and \U$2433 ( \3114 , \724 , RIb55a9e0_559);
and \U$2434 ( \3115 , RIb55aa58_560, \726 );
nor \U$2435 ( \3116 , \3114 , \3115 );
and \U$2436 ( \3117 , \713 , RIb55ae18_568);
and \U$2437 ( \3118 , RIb55ab48_562, \705 );
nor \U$2438 ( \3119 , \3117 , \3118 );
and \U$2439 ( \3120 , \690 , RIb55aad0_561);
and \U$2440 ( \3121 , RIb55abc0_563, \703 );
nor \U$2441 ( \3122 , \3120 , \3121 );
nand \U$2442 ( \3123 , \3113 , \3116 , \3119 , \3122 );
_DC ga6e ( \3124_nGa6e , \3123 , \1243 );
nand \U$2443 ( \3125 , \3124_nGa6e , \1214 );
and \U$2444 ( \3126 , \2856_nGb3b , \1383 );
or \U$2445 ( \3127 , \1257 , \2969_nGabe );
nand \U$2446 ( \3128 , \3127 , \1294 );
nand \U$2447 ( \3129 , \2856_nGb3b , \1261 );
and \U$2448 ( \3130 , \3128 , \3129 );
and \U$2449 ( \3131 , \2969_nGabe , \1416 );
nor \U$2450 ( \3132 , \3126 , \3130 , \3131 );
or \U$2451 ( \3133 , \3125 , \3132 );
nand \U$2452 ( \3134 , \3095 , \3097 , \3133 );
nand \U$2453 ( \3135 , \3093 , \3134 );
xor \U$2454 ( \3136 , \2912 , \2925 );
xor \U$2455 ( \3137 , \3136 , \2974 );
xor \U$2456 ( \3138 , \3135 , \3137 );
xor \U$2457 ( \3139 , \3008 , \3015 );
xor \U$2458 ( \3140 , \3139 , \3023 );
xor \U$2459 ( \3141 , \3033 , \3037 );
xor \U$2460 ( \3142 , \3141 , \3045 );
xor \U$2461 ( \3143 , \3140 , \3142 );
xnor \U$2462 ( \3144 , \3125 , \3132 );
and \U$2463 ( \3145 , \3143 , \3144 );
and \U$2464 ( \3146 , \3140 , \3142 );
or \U$2465 ( \3147 , \3145 , \3146 );
and \U$2466 ( \3148 , \2365_nGda9 , \1650 );
nand \U$2467 ( \3149 , \2365_nGda9 , \1647 );
or \U$2468 ( \3150 , \1576 , \2252_nGe5c );
nand \U$2469 ( \3151 , \3150 , \1798 );
and \U$2470 ( \3152 , \3149 , \3151 );
and \U$2471 ( \3153 , \2252_nGe5c , \1801 );
nor \U$2472 ( \3154 , \3148 , \3152 , \3153 );
nand \U$2473 ( \3155 , \2081_nGf30 , \1864 );
or \U$2474 ( \3156 , \1810 , \2025_nG100c );
nand \U$2475 ( \3157 , \3156 , \1959 );
and \U$2476 ( \3158 , \3155 , \3157 );
and \U$2477 ( \3159 , \1954 , \2025_nG100c );
and \U$2478 ( \3160 , \2081_nGf30 , \1866 );
nor \U$2479 ( \3161 , \3158 , \3159 , \3160 );
xor \U$2480 ( \3162 , \3154 , \3161 );
nand \U$2481 ( \3163 , \2407_nGcdf , \1543 );
or \U$2482 ( \3164 , \1425 , \2621_nGc52 );
nand \U$2483 ( \3165 , \3164 , \1549 );
and \U$2484 ( \3166 , \3163 , \3165 );
and \U$2485 ( \3167 , \1545 , \2621_nGc52 );
and \U$2486 ( \3168 , \2407_nGcdf , \1591 );
nor \U$2487 ( \3169 , \3166 , \3167 , \3168 );
and \U$2488 ( \3170 , \3162 , \3169 );
and \U$2489 ( \3171 , \3154 , \3161 );
or \U$2490 ( \3172 , \3170 , \3171 );
nand \U$2491 ( \3173 , \2856_nGb3b , \1350 );
or \U$2492 ( \3174 , \1310 , \2708_nGbb2 );
nand \U$2493 ( \3175 , \3174 , \1376 );
and \U$2494 ( \3176 , \3173 , \3175 );
and \U$2495 ( \3177 , \1379 , \2708_nGbb2 );
and \U$2496 ( \3178 , \2856_nGb3b , \1353 );
nor \U$2497 ( \3179 , \3176 , \3177 , \3178 );
and \U$2498 ( \3180 , RIb55b610_585, \713 );
and \U$2499 ( \3181 , RIb55b160_575, \740 );
and \U$2500 ( \3182 , \695 , RIb55b4a8_582);
and \U$2501 ( \3183 , RIb55b430_581, \698 );
nor \U$2502 ( \3184 , \3182 , \3183 );
and \U$2503 ( \3185 , \738 , RIb55b0e8_574);
and \U$2504 ( \3186 , RIb55b070_573, \734 );
nor \U$2505 ( \3187 , \3185 , \3186 );
and \U$2506 ( \3188 , \1224 , RIb55af80_571);
and \U$2507 ( \3189 , RIb55aff8_572, \736 );
nor \U$2508 ( \3190 , \3188 , \3189 );
and \U$2509 ( \3191 , \716 , RIb55b598_584);
and \U$2510 ( \3192 , RIb55b520_583, \719 );
nor \U$2511 ( \3193 , \3191 , \3192 );
nand \U$2512 ( \3194 , \3184 , \3187 , \3190 , \3193 );
nor \U$2513 ( \3195 , \3180 , \3181 , \3194 );
and \U$2514 ( \3196 , \703 , RIb55b3b8_580);
and \U$2515 ( \3197 , RIb55b250_577, \726 );
nor \U$2516 ( \3198 , \3196 , \3197 );
and \U$2517 ( \3199 , \710 , RIb55b688_586);
and \U$2518 ( \3200 , RIb55b340_579, \705 );
nor \U$2519 ( \3201 , \3199 , \3200 );
and \U$2520 ( \3202 , \690 , RIb55b2c8_578);
and \U$2521 ( \3203 , RIb55b1d8_576, \724 );
nor \U$2522 ( \3204 , \3202 , \3203 );
nand \U$2523 ( \3205 , \3195 , \3198 , \3201 , \3204 );
_DC g959 ( \3206_nG959 , \3205 , \1243 );
nand \U$2524 ( \3207 , \3206_nG959 , \1214 );
xor \U$2525 ( \3208 , \3179 , \3207 );
and \U$2526 ( \3209 , \2969_nGabe , \1383 );
or \U$2527 ( \3210 , \1257 , \3124_nGa6e );
nand \U$2528 ( \3211 , \3210 , \1294 );
nand \U$2529 ( \3212 , \2969_nGabe , \1261 );
and \U$2530 ( \3213 , \3211 , \3212 );
and \U$2531 ( \3214 , \3124_nGa6e , \1416 );
nor \U$2532 ( \3215 , \3209 , \3213 , \3214 );
and \U$2533 ( \3216 , \3208 , \3215 );
and \U$2534 ( \3217 , \3179 , \3207 );
or \U$2535 ( \3218 , \3216 , \3217 );
nand \U$2536 ( \3219 , \3172 , \3218 );
or \U$2537 ( \3220 , \2535 , \1632 );
or \U$2538 ( \3221 , \1538_nG13f2 , \2419 );
or \U$2539 ( \3222 , \1628_nG1300 , \2418 );
nand \U$2540 ( \3223 , \3220 , \3221 , \3222 );
not \U$2541 ( \3224 , \1789_nG1116 );
or \U$2542 ( \3225 , \2099 , \3224 );
not \U$2543 ( \3226 , \1707_nG11f7 );
or \U$2544 ( \3227 , \3226 , \2200 );
or \U$2545 ( \3228 , \2101 , \3224 );
or \U$2546 ( \3229 , \1970 , \1707_nG11f7 );
nand \U$2547 ( \3230 , \3229 , \2197 );
nand \U$2548 ( \3231 , \3228 , \3230 );
nand \U$2549 ( \3232 , \3225 , \3227 , \3231 );
and \U$2550 ( \3233 , \3223 , \3232 );
and \U$2551 ( \3234 , \3219 , \3233 );
nor \U$2552 ( \3235 , \3218 , \3172 );
nor \U$2553 ( \3236 , \3234 , \3235 );
nand \U$2554 ( \3237 , \3147 , \3236 );
not \U$2555 ( \3238 , \2924 );
not \U$2556 ( \3239 , \2919 );
or \U$2557 ( \3240 , \3238 , \3239 );
or \U$2558 ( \3241 , \2919 , \2924 );
nand \U$2559 ( \3242 , \3240 , \3241 );
and \U$2560 ( \3243 , \3237 , \3242 );
nor \U$2561 ( \3244 , \3236 , \3147 );
nor \U$2562 ( \3245 , \3243 , \3244 );
and \U$2563 ( \3246 , \3138 , \3245 );
and \U$2564 ( \3247 , \3135 , \3137 );
or \U$2565 ( \3248 , \3246 , \3247 );
nor \U$2566 ( \3249 , \3087 , \3248 );
xor \U$2567 ( \3250 , \3080 , \3249 );
and \U$2568 ( \3251 , \3087 , \3248 );
nor \U$2569 ( \3252 , \3251 , \3249 );
xor \U$2570 ( \3253 , \3135 , \3137 );
xor \U$2571 ( \3254 , \3253 , \3245 );
not \U$2572 ( \3255 , \3049 );
not \U$2573 ( \3256 , \3061 );
or \U$2574 ( \3257 , \3255 , \3256 );
or \U$2575 ( \3258 , \3061 , \3049 );
nand \U$2576 ( \3259 , \3257 , \3258 );
not \U$2577 ( \3260 , \3259 );
not \U$2578 ( \3261 , \3001 );
and \U$2579 ( \3262 , \3260 , \3261 );
and \U$2580 ( \3263 , \3259 , \3001 );
nor \U$2581 ( \3264 , \3262 , \3263 );
nor \U$2582 ( \3265 , \3254 , \3264 );
xor \U$2583 ( \3266 , \3252 , \3265 );
and \U$2584 ( \3267 , \3254 , \3264 );
nor \U$2585 ( \3268 , \3267 , \3265 );
xor \U$2586 ( \3269 , \3140 , \3142 );
xor \U$2587 ( \3270 , \3269 , \3144 );
not \U$2588 ( \3271 , \3270 );
xor \U$2589 ( \3272 , \3223 , \3232 );
not \U$2590 ( \3273 , \3272 );
xor \U$2591 ( \3274 , \3154 , \3161 );
xor \U$2592 ( \3275 , \3274 , \3169 );
nor \U$2593 ( \3276 , \3273 , \3275 );
xor \U$2594 ( \3277 , \3271 , \3276 );
nand \U$2595 ( \3278 , \2621_nGc52 , \1543 );
or \U$2596 ( \3279 , \1425 , \2708_nGbb2 );
nand \U$2597 ( \3280 , \3279 , \1549 );
and \U$2598 ( \3281 , \3278 , \3280 );
and \U$2599 ( \3282 , \1545 , \2708_nGbb2 );
and \U$2600 ( \3283 , \2621_nGc52 , \1591 );
nor \U$2601 ( \3284 , \3281 , \3282 , \3283 );
and \U$2602 ( \3285 , \2407_nGcdf , \1650 );
nand \U$2603 ( \3286 , \2407_nGcdf , \1647 );
or \U$2604 ( \3287 , \1576 , \2365_nGda9 );
nand \U$2605 ( \3288 , \3287 , \1798 );
and \U$2606 ( \3289 , \3286 , \3288 );
and \U$2607 ( \3290 , \2365_nGda9 , \1801 );
nor \U$2608 ( \3291 , \3285 , \3289 , \3290 );
xor \U$2609 ( \3292 , \3284 , \3291 );
nand \U$2610 ( \3293 , \2969_nGabe , \1350 );
or \U$2611 ( \3294 , \1310 , \2856_nGb3b );
nand \U$2612 ( \3295 , \3294 , \1376 );
and \U$2613 ( \3296 , \3293 , \3295 );
and \U$2614 ( \3297 , \1379 , \2856_nGb3b );
and \U$2615 ( \3298 , \2969_nGabe , \1353 );
nor \U$2616 ( \3299 , \3296 , \3297 , \3298 );
and \U$2617 ( \3300 , \3292 , \3299 );
and \U$2618 ( \3301 , \3284 , \3291 );
or \U$2619 ( \3302 , \3300 , \3301 );
nand \U$2620 ( \3303 , \2025_nG100c , \2098 );
or \U$2621 ( \3304 , \1970 , \1789_nG1116 );
nand \U$2622 ( \3305 , \3304 , \2197 );
and \U$2623 ( \3306 , \3303 , \3305 );
and \U$2624 ( \3307 , \2201 , \1789_nG1116 );
and \U$2625 ( \3308 , \2025_nG100c , \2203 );
nor \U$2626 ( \3309 , \3306 , \3307 , \3308 );
and \U$2627 ( \3310 , \1629 , \2532 );
and \U$2628 ( \3311 , \2417 , \3226 );
and \U$2629 ( \3312 , \1628_nG1300 , \2536 );
nor \U$2630 ( \3313 , \3310 , \3311 , \3312 );
xor \U$2631 ( \3314 , \3309 , \3313 );
nand \U$2632 ( \3315 , \2252_nGe5c , \1864 );
or \U$2633 ( \3316 , \1810 , \2081_nGf30 );
nand \U$2634 ( \3317 , \3316 , \1959 );
and \U$2635 ( \3318 , \3315 , \3317 );
and \U$2636 ( \3319 , \1954 , \2081_nGf30 );
and \U$2637 ( \3320 , \2252_nGe5c , \1866 );
nor \U$2638 ( \3321 , \3318 , \3319 , \3320 );
and \U$2639 ( \3322 , \3314 , \3321 );
and \U$2640 ( \3323 , \3309 , \3313 );
or \U$2641 ( \3324 , \3322 , \3323 );
xor \U$2642 ( \3325 , \3302 , \3324 );
xor \U$2643 ( \3326 , \3179 , \3207 );
xor \U$2644 ( \3327 , \3326 , \3215 );
and \U$2645 ( \3328 , \3325 , \3327 );
and \U$2646 ( \3329 , \3302 , \3324 );
or \U$2647 ( \3330 , \3328 , \3329 );
not \U$2648 ( \3331 , \3330 );
and \U$2649 ( \3332 , \3277 , \3331 );
and \U$2650 ( \3333 , \3271 , \3276 );
or \U$2651 ( \3334 , \3332 , \3333 );
not \U$2652 ( \3335 , \3134 );
not \U$2653 ( \3336 , \3092 );
or \U$2654 ( \3337 , \3335 , \3336 );
or \U$2655 ( \3338 , \3092 , \3134 );
nand \U$2656 ( \3339 , \3337 , \3338 );
xor \U$2657 ( \3340 , \3334 , \3339 );
not \U$2658 ( \3341 , \3242 );
not \U$2659 ( \3342 , \3244 );
nand \U$2660 ( \3343 , \3342 , \3237 );
not \U$2661 ( \3344 , \3343 );
or \U$2662 ( \3345 , \3341 , \3344 );
or \U$2663 ( \3346 , \3343 , \3242 );
nand \U$2664 ( \3347 , \3345 , \3346 );
and \U$2665 ( \3348 , \3340 , \3347 );
and \U$2666 ( \3349 , \3334 , \3339 );
or \U$2667 ( \3350 , \3348 , \3349 );
xor \U$2668 ( \3351 , \3268 , \3350 );
xor \U$2669 ( \3352 , \3334 , \3339 );
xor \U$2670 ( \3353 , \3352 , \3347 );
xor \U$2671 ( \3354 , \3271 , \3276 );
xor \U$2672 ( \3355 , \3354 , \3331 );
not \U$2673 ( \3356 , \3233 );
not \U$2674 ( \3357 , \3235 );
nand \U$2675 ( \3358 , \3357 , \3219 );
not \U$2676 ( \3359 , \3358 );
or \U$2677 ( \3360 , \3356 , \3359 );
or \U$2678 ( \3361 , \3358 , \3233 );
nand \U$2679 ( \3362 , \3360 , \3361 );
nor \U$2680 ( \3363 , \3355 , \3362 );
nand \U$2681 ( \3364 , \2081_nGf30 , \2098 );
or \U$2682 ( \3365 , \1970 , \2025_nG100c );
nand \U$2683 ( \3366 , \3365 , \2197 );
and \U$2684 ( \3367 , \3364 , \3366 );
and \U$2685 ( \3368 , \2201 , \2025_nG100c );
and \U$2686 ( \3369 , \2081_nGf30 , \2203 );
nor \U$2687 ( \3370 , \3367 , \3368 , \3369 );
and \U$2688 ( \3371 , \3226 , \2532 );
and \U$2689 ( \3372 , \2417 , \3224 );
and \U$2690 ( \3373 , \1707_nG11f7 , \2536 );
nor \U$2691 ( \3374 , \3371 , \3372 , \3373 );
xor \U$2692 ( \3375 , \3370 , \3374 );
and \U$2693 ( \3376 , \3375 , \1257 );
and \U$2694 ( \3377 , \3370 , \3374 );
or \U$2695 ( \3378 , \3376 , \3377 );
and \U$2696 ( \3379 , \2621_nGc52 , \1650 );
nand \U$2697 ( \3380 , \2621_nGc52 , \1647 );
or \U$2698 ( \3381 , \1576 , \2407_nGcdf );
nand \U$2699 ( \3382 , \3381 , \1798 );
and \U$2700 ( \3383 , \3380 , \3382 );
and \U$2701 ( \3384 , \2407_nGcdf , \1801 );
nor \U$2702 ( \3385 , \3379 , \3383 , \3384 );
nand \U$2703 ( \3386 , \2365_nGda9 , \1864 );
or \U$2704 ( \3387 , \1810 , \2252_nGe5c );
nand \U$2705 ( \3388 , \3387 , \1959 );
and \U$2706 ( \3389 , \3386 , \3388 );
and \U$2707 ( \3390 , \1954 , \2252_nGe5c );
and \U$2708 ( \3391 , \2365_nGda9 , \1866 );
nor \U$2709 ( \3392 , \3389 , \3390 , \3391 );
xor \U$2710 ( \3393 , \3385 , \3392 );
nand \U$2711 ( \3394 , \2708_nGbb2 , \1543 );
or \U$2712 ( \3395 , \1425 , \2856_nGb3b );
nand \U$2713 ( \3396 , \3395 , \1549 );
and \U$2714 ( \3397 , \3394 , \3396 );
and \U$2715 ( \3398 , \1545 , \2856_nGb3b );
and \U$2716 ( \3399 , \2708_nGbb2 , \1591 );
nor \U$2717 ( \3400 , \3397 , \3398 , \3399 );
and \U$2718 ( \3401 , \3393 , \3400 );
and \U$2719 ( \3402 , \3385 , \3392 );
or \U$2720 ( \3403 , \3401 , \3402 );
xor \U$2721 ( \3404 , \3378 , \3403 );
and \U$2722 ( \3405 , \3124_nGa6e , \1383 );
or \U$2723 ( \3406 , \1257 , \3206_nG959 );
nand \U$2724 ( \3407 , \3406 , \1294 );
nand \U$2725 ( \3408 , \3124_nGa6e , \1261 );
and \U$2726 ( \3409 , \3407 , \3408 );
and \U$2727 ( \3410 , \3206_nG959 , \1416 );
nor \U$2728 ( \3411 , \3405 , \3409 , \3410 );
and \U$2729 ( \3412 , \3404 , \3411 );
and \U$2730 ( \3413 , \3378 , \3403 );
or \U$2731 ( \3414 , \3412 , \3413 );
not \U$2732 ( \3415 , \3275 );
not \U$2733 ( \3416 , \3272 );
and \U$2734 ( \3417 , \3415 , \3416 );
and \U$2735 ( \3418 , \3275 , \3272 );
nor \U$2736 ( \3419 , \3417 , \3418 );
xor \U$2737 ( \3420 , \3414 , \3419 );
xor \U$2738 ( \3421 , \3302 , \3324 );
xor \U$2739 ( \3422 , \3421 , \3327 );
and \U$2740 ( \3423 , \3420 , \3422 );
and \U$2741 ( \3424 , \3414 , \3419 );
or \U$2742 ( \3425 , \3423 , \3424 );
or \U$2743 ( \3426 , \3363 , \3425 );
nand \U$2744 ( \3427 , \3362 , \3355 );
nand \U$2745 ( \3428 , \3426 , \3427 );
xor \U$2746 ( \3429 , \3353 , \3428 );
not \U$2747 ( \3430 , \3425 );
not \U$2748 ( \3431 , \3363 );
nand \U$2749 ( \3432 , \3431 , \3427 );
not \U$2750 ( \3433 , \3432 );
or \U$2751 ( \3434 , \3430 , \3433 );
or \U$2752 ( \3435 , \3432 , \3425 );
nand \U$2753 ( \3436 , \3434 , \3435 );
xor \U$2754 ( \3437 , \3378 , \3403 );
xor \U$2755 ( \3438 , \3437 , \3411 );
xor \U$2756 ( \3439 , \3309 , \3313 );
xor \U$2757 ( \3440 , \3439 , \3321 );
or \U$2758 ( \3441 , \3438 , \3440 );
nand \U$2759 ( \3442 , \3124_nGa6e , \1350 );
or \U$2760 ( \3443 , \1310 , \2969_nGabe );
nand \U$2761 ( \3444 , \3443 , \1376 );
and \U$2762 ( \3445 , \3442 , \3444 );
and \U$2763 ( \3446 , \1379 , \2969_nGabe );
and \U$2764 ( \3447 , \3124_nGa6e , \1353 );
nor \U$2765 ( \3448 , \3445 , \3446 , \3447 );
nand \U$2766 ( \3449 , \2252_nGe5c , \2098 );
or \U$2767 ( \3450 , \1970 , \2081_nGf30 );
nand \U$2768 ( \3451 , \3450 , \2197 );
and \U$2769 ( \3452 , \3449 , \3451 );
and \U$2770 ( \3453 , \2201 , \2081_nGf30 );
and \U$2771 ( \3454 , \2252_nGe5c , \2203 );
nor \U$2772 ( \3455 , \3452 , \3453 , \3454 );
and \U$2773 ( \3456 , \3224 , \2532 );
not \U$2774 ( \3457 , \2025_nG100c );
and \U$2775 ( \3458 , \2417 , \3457 );
and \U$2776 ( \3459 , \1789_nG1116 , \2536 );
nor \U$2777 ( \3460 , \3456 , \3458 , \3459 );
xor \U$2778 ( \3461 , \3455 , \3460 );
nand \U$2779 ( \3462 , \2407_nGcdf , \1864 );
or \U$2780 ( \3463 , \1810 , \2365_nGda9 );
nand \U$2781 ( \3464 , \3463 , \1959 );
and \U$2782 ( \3465 , \3462 , \3464 );
and \U$2783 ( \3466 , \1954 , \2365_nGda9 );
and \U$2784 ( \3467 , \2407_nGcdf , \1866 );
nor \U$2785 ( \3468 , \3465 , \3466 , \3467 );
and \U$2786 ( \3469 , \3461 , \3468 );
and \U$2787 ( \3470 , \3455 , \3460 );
or \U$2788 ( \3471 , \3469 , \3470 );
xor \U$2789 ( \3472 , \3448 , \3471 );
nand \U$2790 ( \3473 , \2856_nGb3b , \1543 );
or \U$2791 ( \3474 , \1425 , \2969_nGabe );
nand \U$2792 ( \3475 , \3474 , \1549 );
and \U$2793 ( \3476 , \3473 , \3475 );
and \U$2794 ( \3477 , \1545 , \2969_nGabe );
and \U$2795 ( \3478 , \2856_nGb3b , \1591 );
nor \U$2796 ( \3479 , \3476 , \3477 , \3478 );
and \U$2797 ( \3480 , \2708_nGbb2 , \1650 );
nand \U$2798 ( \3481 , \2708_nGbb2 , \1647 );
or \U$2799 ( \3482 , \1576 , \2621_nGc52 );
nand \U$2800 ( \3483 , \3482 , \1798 );
and \U$2801 ( \3484 , \3481 , \3483 );
and \U$2802 ( \3485 , \2621_nGc52 , \1801 );
nor \U$2803 ( \3486 , \3480 , \3484 , \3485 );
xor \U$2804 ( \3487 , \3479 , \3486 );
nand \U$2805 ( \3488 , \3206_nG959 , \1350 );
or \U$2806 ( \3489 , \1310 , \3124_nGa6e );
nand \U$2807 ( \3490 , \3489 , \1376 );
and \U$2808 ( \3491 , \3488 , \3490 );
and \U$2809 ( \3492 , \1379 , \3124_nGa6e );
and \U$2810 ( \3493 , \3206_nG959 , \1353 );
nor \U$2811 ( \3494 , \3491 , \3492 , \3493 );
and \U$2812 ( \3495 , \3487 , \3494 );
and \U$2813 ( \3496 , \3479 , \3486 );
or \U$2814 ( \3497 , \3495 , \3496 );
and \U$2815 ( \3498 , \3472 , \3497 );
and \U$2816 ( \3499 , \3448 , \3471 );
or \U$2817 ( \3500 , \3498 , \3499 );
xor \U$2818 ( \3501 , \3284 , \3291 );
xor \U$2819 ( \3502 , \3501 , \3299 );
xor \U$2820 ( \3503 , \3500 , \3502 );
xor \U$2821 ( \3504 , \3385 , \3392 );
xor \U$2822 ( \3505 , \3504 , \3400 );
xor \U$2823 ( \3506 , \3370 , \3374 );
xor \U$2824 ( \3507 , \3506 , \1257 );
and \U$2825 ( \3508 , \3505 , \3507 );
nand \U$2826 ( \3509 , \3206_nG959 , \1261 );
and \U$2827 ( \3510 , \1256 , \3509 );
and \U$2828 ( \3511 , \3206_nG959 , \1383 );
nor \U$2829 ( \3512 , \3510 , \3511 );
xor \U$2830 ( \3513 , \3370 , \3374 );
xor \U$2831 ( \3514 , \3513 , \1257 );
and \U$2832 ( \3515 , \3512 , \3514 );
and \U$2833 ( \3516 , \3505 , \3512 );
or \U$2834 ( \3517 , \3508 , \3515 , \3516 );
and \U$2835 ( \3518 , \3503 , \3517 );
and \U$2836 ( \3519 , \3500 , \3502 );
or \U$2837 ( \3520 , \3518 , \3519 );
xor \U$2838 ( \3521 , \3441 , \3520 );
xor \U$2839 ( \3522 , \3414 , \3419 );
xor \U$2840 ( \3523 , \3522 , \3422 );
and \U$2841 ( \3524 , \3521 , \3523 );
and \U$2842 ( \3525 , \3441 , \3520 );
or \U$2843 ( \3526 , \3524 , \3525 );
xor \U$2844 ( \3527 , \3436 , \3526 );
and \U$2845 ( \3528 , \2856_nGb3b , \1650 );
nand \U$2846 ( \3529 , \2856_nGb3b , \1647 );
or \U$2847 ( \3530 , \1576 , \2708_nGbb2 );
nand \U$2848 ( \3531 , \3530 , \1798 );
and \U$2849 ( \3532 , \3529 , \3531 );
and \U$2850 ( \3533 , \2708_nGbb2 , \1801 );
nor \U$2851 ( \3534 , \3528 , \3532 , \3533 );
nand \U$2852 ( \3535 , \2621_nGc52 , \1864 );
or \U$2853 ( \3536 , \1810 , \2407_nGcdf );
nand \U$2854 ( \3537 , \3536 , \1959 );
and \U$2855 ( \3538 , \3535 , \3537 );
and \U$2856 ( \3539 , \1954 , \2407_nGcdf );
and \U$2857 ( \3540 , \2621_nGc52 , \1866 );
nor \U$2858 ( \3541 , \3538 , \3539 , \3540 );
xor \U$2859 ( \3542 , \3534 , \3541 );
nand \U$2860 ( \3543 , \2969_nGabe , \1543 );
or \U$2861 ( \3544 , \1425 , \3124_nGa6e );
nand \U$2862 ( \3545 , \3544 , \1549 );
and \U$2863 ( \3546 , \3543 , \3545 );
and \U$2864 ( \3547 , \1545 , \3124_nGa6e );
and \U$2865 ( \3548 , \2969_nGabe , \1591 );
nor \U$2866 ( \3549 , \3546 , \3547 , \3548 );
and \U$2867 ( \3550 , \3542 , \3549 );
and \U$2868 ( \3551 , \3534 , \3541 );
or \U$2869 ( \3552 , \3550 , \3551 );
nand \U$2870 ( \3553 , \2365_nGda9 , \2098 );
or \U$2871 ( \3554 , \1970 , \2252_nGe5c );
nand \U$2872 ( \3555 , \3554 , \2197 );
and \U$2873 ( \3556 , \3553 , \3555 );
and \U$2874 ( \3557 , \2201 , \2252_nGe5c );
and \U$2875 ( \3558 , \2365_nGda9 , \2203 );
nor \U$2876 ( \3559 , \3556 , \3557 , \3558 );
and \U$2877 ( \3560 , \3457 , \2532 );
not \U$2878 ( \3561 , \2081_nGf30 );
and \U$2879 ( \3562 , \2417 , \3561 );
and \U$2880 ( \3563 , \2025_nG100c , \2536 );
nor \U$2881 ( \3564 , \3560 , \3562 , \3563 );
xor \U$2882 ( \3565 , \3559 , \3564 );
and \U$2883 ( \3566 , \3565 , \1310 );
and \U$2884 ( \3567 , \3559 , \3564 );
or \U$2885 ( \3568 , \3566 , \3567 );
xor \U$2886 ( \3569 , \3552 , \3568 );
xor \U$2887 ( \3570 , \3479 , \3486 );
xor \U$2888 ( \3571 , \3570 , \3494 );
and \U$2889 ( \3572 , \3569 , \3571 );
and \U$2890 ( \3573 , \3552 , \3568 );
or \U$2891 ( \3574 , \3572 , \3573 );
xor \U$2892 ( \3575 , \3448 , \3471 );
xor \U$2893 ( \3576 , \3575 , \3497 );
xor \U$2894 ( \3577 , \3574 , \3576 );
xor \U$2895 ( \3578 , \3370 , \3374 );
xor \U$2896 ( \3579 , \3578 , \1257 );
xor \U$2897 ( \3580 , \3505 , \3512 );
xor \U$2898 ( \3581 , \3579 , \3580 );
and \U$2899 ( \3582 , \3577 , \3581 );
and \U$2900 ( \3583 , \3574 , \3576 );
or \U$2901 ( \3584 , \3582 , \3583 );
xor \U$2902 ( \3585 , \3500 , \3502 );
xor \U$2903 ( \3586 , \3585 , \3517 );
xor \U$2904 ( \3587 , \3584 , \3586 );
xnor \U$2905 ( \3588 , \3440 , \3438 );
xor \U$2906 ( \3589 , \3587 , \3588 );
not \U$2907 ( \3590 , \3589 );
xor \U$2908 ( \3591 , \3574 , \3576 );
xor \U$2909 ( \3592 , \3591 , \3581 );
nand \U$2910 ( \3593 , \2407_nGcdf , \2098 );
or \U$2911 ( \3594 , \1970 , \2365_nGda9 );
nand \U$2912 ( \3595 , \3594 , \2197 );
and \U$2913 ( \3596 , \3593 , \3595 );
and \U$2914 ( \3597 , \2201 , \2365_nGda9 );
and \U$2915 ( \3598 , \2407_nGcdf , \2203 );
nor \U$2916 ( \3599 , \3596 , \3597 , \3598 );
and \U$2917 ( \3600 , \3561 , \2532 );
not \U$2918 ( \3601 , \2252_nGe5c );
and \U$2919 ( \3602 , \2417 , \3601 );
and \U$2920 ( \3603 , \2081_nGf30 , \2536 );
nor \U$2921 ( \3604 , \3600 , \3602 , \3603 );
xor \U$2922 ( \3605 , \3599 , \3604 );
nand \U$2923 ( \3606 , \2708_nGbb2 , \1864 );
or \U$2924 ( \3607 , \1810 , \2621_nGc52 );
nand \U$2925 ( \3608 , \3607 , \1959 );
and \U$2926 ( \3609 , \3606 , \3608 );
and \U$2927 ( \3610 , \1954 , \2621_nGc52 );
and \U$2928 ( \3611 , \2708_nGbb2 , \1866 );
nor \U$2929 ( \3612 , \3609 , \3610 , \3611 );
and \U$2930 ( \3613 , \3605 , \3612 );
and \U$2931 ( \3614 , \3599 , \3604 );
or \U$2932 ( \3615 , \3613 , \3614 );
xor \U$2933 ( \3616 , \3534 , \3541 );
xor \U$2934 ( \3617 , \3616 , \3549 );
and \U$2935 ( \3618 , \3615 , \3617 );
and \U$2936 ( \3619 , \3206_nG959 , \1379 );
not \U$2937 ( \3620 , \3206_nG959 );
and \U$2938 ( \3621 , \3620 , \1352 );
not \U$2939 ( \3622 , \1376 );
nor \U$2940 ( \3623 , \3619 , \3621 , \3622 );
xor \U$2941 ( \3624 , \3534 , \3541 );
xor \U$2942 ( \3625 , \3624 , \3549 );
and \U$2943 ( \3626 , \3623 , \3625 );
and \U$2944 ( \3627 , \3615 , \3623 );
or \U$2945 ( \3628 , \3618 , \3626 , \3627 );
xor \U$2946 ( \3629 , \3455 , \3460 );
xor \U$2947 ( \3630 , \3629 , \3468 );
xor \U$2948 ( \3631 , \3628 , \3630 );
xor \U$2949 ( \3632 , \3552 , \3568 );
xor \U$2950 ( \3633 , \3632 , \3571 );
and \U$2951 ( \3634 , \3631 , \3633 );
and \U$2952 ( \3635 , \3628 , \3630 );
or \U$2953 ( \3636 , \3634 , \3635 );
nor \U$2954 ( \3637 , \3592 , \3636 );
xor \U$2955 ( \3638 , \3590 , \3637 );
and \U$2956 ( \3639 , \3592 , \3636 );
nor \U$2957 ( \3640 , \3639 , \3637 );
xor \U$2958 ( \3641 , \3628 , \3630 );
xor \U$2959 ( \3642 , \3641 , \3633 );
and \U$2960 ( \3643 , \2969_nGabe , \1650 );
nand \U$2961 ( \3644 , \2969_nGabe , \1647 );
or \U$2962 ( \3645 , \1576 , \2856_nGb3b );
nand \U$2963 ( \3646 , \3645 , \1798 );
and \U$2964 ( \3647 , \3644 , \3646 );
and \U$2965 ( \3648 , \2856_nGb3b , \1801 );
nor \U$2966 ( \3649 , \3643 , \3647 , \3648 );
nand \U$2967 ( \3650 , \2621_nGc52 , \2098 );
or \U$2968 ( \3651 , \1970 , \2407_nGcdf );
nand \U$2969 ( \3652 , \3651 , \2197 );
and \U$2970 ( \3653 , \3650 , \3652 );
and \U$2971 ( \3654 , \2201 , \2407_nGcdf );
and \U$2972 ( \3655 , \2621_nGc52 , \2203 );
nor \U$2973 ( \3656 , \3653 , \3654 , \3655 );
and \U$2974 ( \3657 , \3601 , \2532 );
and \U$2975 ( \3658 , \2417 , \2673 );
and \U$2976 ( \3659 , \2252_nGe5c , \2536 );
nor \U$2977 ( \3660 , \3657 , \3658 , \3659 );
xor \U$2978 ( \3661 , \3656 , \3660 );
and \U$2979 ( \3662 , \3661 , \1425 );
and \U$2980 ( \3663 , \3656 , \3660 );
or \U$2981 ( \3664 , \3662 , \3663 );
xor \U$2982 ( \3665 , \3649 , \3664 );
and \U$2983 ( \3666 , \3124_nGa6e , \1650 );
nand \U$2984 ( \3667 , \3124_nGa6e , \1647 );
or \U$2985 ( \3668 , \1576 , \2969_nGabe );
nand \U$2986 ( \3669 , \3668 , \1798 );
and \U$2987 ( \3670 , \3667 , \3669 );
and \U$2988 ( \3671 , \2969_nGabe , \1801 );
nor \U$2989 ( \3672 , \3666 , \3670 , \3671 );
nand \U$2990 ( \3673 , \2856_nGb3b , \1864 );
or \U$2991 ( \3674 , \1810 , \2708_nGbb2 );
nand \U$2992 ( \3675 , \3674 , \1959 );
and \U$2993 ( \3676 , \3673 , \3675 );
and \U$2994 ( \3677 , \1954 , \2708_nGbb2 );
and \U$2995 ( \3678 , \2856_nGb3b , \1866 );
nor \U$2996 ( \3679 , \3676 , \3677 , \3678 );
xor \U$2997 ( \3680 , \3672 , \3679 );
and \U$2998 ( \3681 , \1591 , \3206_nG959 );
nand \U$2999 ( \3682 , \3206_nG959 , \1543 );
and \U$3000 ( \3683 , \3682 , \1547 );
nor \U$3001 ( \3684 , \3681 , \3683 );
and \U$3002 ( \3685 , \3680 , \3684 );
and \U$3003 ( \3686 , \3672 , \3679 );
or \U$3004 ( \3687 , \3685 , \3686 );
and \U$3005 ( \3688 , \3665 , \3687 );
and \U$3006 ( \3689 , \3649 , \3664 );
or \U$3007 ( \3690 , \3688 , \3689 );
xor \U$3008 ( \3691 , \3559 , \3564 );
xor \U$3009 ( \3692 , \3691 , \1310 );
nand \U$3010 ( \3693 , \3690 , \3692 );
not \U$3011 ( \3694 , \3124_nGa6e );
or \U$3012 ( \3695 , \1656 , \3694 );
or \U$3013 ( \3696 , \3620 , \1658 );
or \U$3014 ( \3697 , \1590 , \3694 );
or \U$3015 ( \3698 , \1425 , \3206_nG959 );
nand \U$3016 ( \3699 , \3698 , \1549 );
nand \U$3017 ( \3700 , \3697 , \3699 );
nand \U$3018 ( \3701 , \3695 , \3696 , \3700 );
not \U$3019 ( \3702 , \3701 );
xor \U$3020 ( \3703 , \3599 , \3604 );
xor \U$3021 ( \3704 , \3703 , \3612 );
nor \U$3022 ( \3705 , \3702 , \3704 );
and \U$3023 ( \3706 , \3693 , \3705 );
nor \U$3024 ( \3707 , \3692 , \3690 );
nor \U$3025 ( \3708 , \3706 , \3707 );
nor \U$3026 ( \3709 , \3642 , \3708 );
xor \U$3027 ( \3710 , \3640 , \3709 );
nand \U$3028 ( \3711 , \2708_nGbb2 , \2098 );
or \U$3029 ( \3712 , \1970 , \2621_nGc52 );
nand \U$3030 ( \3713 , \3712 , \2197 );
and \U$3031 ( \3714 , \3711 , \3713 );
and \U$3032 ( \3715 , \2201 , \2621_nGc52 );
and \U$3033 ( \3716 , \2708_nGbb2 , \2203 );
nor \U$3034 ( \3717 , \3714 , \3715 , \3716 );
and \U$3035 ( \3718 , \2673 , \2532 );
and \U$3036 ( \3719 , \2417 , \2712 );
and \U$3037 ( \3720 , \2365_nGda9 , \2536 );
nor \U$3038 ( \3721 , \3718 , \3719 , \3720 );
xor \U$3039 ( \3722 , \3717 , \3721 );
nand \U$3040 ( \3723 , \2969_nGabe , \1864 );
or \U$3041 ( \3724 , \1810 , \2856_nGb3b );
nand \U$3042 ( \3725 , \3724 , \1959 );
and \U$3043 ( \3726 , \3723 , \3725 );
and \U$3044 ( \3727 , \1954 , \2856_nGb3b );
and \U$3045 ( \3728 , \2969_nGabe , \1866 );
nor \U$3046 ( \3729 , \3726 , \3727 , \3728 );
xor \U$3047 ( \3730 , \3722 , \3729 );
not \U$3048 ( \3731 , \3730 );
or \U$3049 ( \3732 , \1867 , \3694 );
not \U$3050 ( \3733 , \2969_nGabe );
or \U$3051 ( \3734 , \3733 , \1955 );
or \U$3052 ( \3735 , \1865 , \3694 );
or \U$3053 ( \3736 , \1810 , \2969_nGabe );
nand \U$3054 ( \3737 , \3736 , \1959 );
nand \U$3055 ( \3738 , \3735 , \3737 );
nand \U$3056 ( \3739 , \3732 , \3734 , \3738 );
or \U$3057 ( \3740 , \1873 , \3620 );
or \U$3058 ( \3741 , \3206_nG959 , \1576 );
nand \U$3059 ( \3742 , \3740 , \3741 , \1798 );
and \U$3060 ( \3743 , \3739 , \3742 );
not \U$3061 ( \3744 , \3743 );
and \U$3062 ( \3745 , \3206_nG959 , \1650 );
nand \U$3063 ( \3746 , \3206_nG959 , \1647 );
or \U$3064 ( \3747 , \1576 , \3124_nGa6e );
nand \U$3065 ( \3748 , \3747 , \1798 );
and \U$3066 ( \3749 , \3746 , \3748 );
and \U$3067 ( \3750 , \3124_nGa6e , \1801 );
nor \U$3068 ( \3751 , \3745 , \3749 , \3750 );
or \U$3069 ( \3752 , \2535 , \2712 );
or \U$3070 ( \3753 , \2407_nGcdf , \2419 );
or \U$3071 ( \3754 , \2621_nGc52 , \2418 );
nand \U$3072 ( \3755 , \3752 , \3753 , \3754 );
not \U$3073 ( \3756 , \3755 );
nand \U$3074 ( \3757 , \2856_nGb3b , \2098 );
or \U$3075 ( \3758 , \1970 , \2708_nGbb2 );
nand \U$3076 ( \3759 , \3758 , \2197 );
and \U$3077 ( \3760 , \3757 , \3759 );
and \U$3078 ( \3761 , \2201 , \2708_nGbb2 );
and \U$3079 ( \3762 , \2856_nGb3b , \2203 );
nor \U$3080 ( \3763 , \3760 , \3761 , \3762 );
nand \U$3081 ( \3764 , \3756 , \3763 );
and \U$3082 ( \3765 , \1649 , \3764 );
not \U$3083 ( \3766 , \3763 );
and \U$3084 ( \3767 , \3755 , \3766 );
nor \U$3085 ( \3768 , \3765 , \3767 );
nor \U$3086 ( \3769 , \3751 , \3768 );
not \U$3087 ( \3770 , \3769 );
nand \U$3088 ( \3771 , \3768 , \3751 );
nand \U$3089 ( \3772 , \3770 , \3771 );
not \U$3090 ( \3773 , \3772 );
or \U$3091 ( \3774 , \3744 , \3773 );
or \U$3092 ( \3775 , \3772 , \3743 );
nand \U$3093 ( \3776 , \3774 , \3775 );
xor \U$3094 ( \3777 , \3731 , \3776 );
not \U$3095 ( \3778 , \3755 );
and \U$3096 ( \3779 , \3763 , \1649 );
not \U$3097 ( \3780 , \3763 );
and \U$3098 ( \3781 , \3780 , \1576 );
nor \U$3099 ( \3782 , \3779 , \3781 );
not \U$3100 ( \3783 , \3782 );
or \U$3101 ( \3784 , \3778 , \3783 );
or \U$3102 ( \3785 , \3782 , \3755 );
nand \U$3103 ( \3786 , \3784 , \3785 );
nand \U$3104 ( \3787 , \2969_nGabe , \2098 );
or \U$3105 ( \3788 , \1970 , \2856_nGb3b );
nand \U$3106 ( \3789 , \3788 , \2197 );
and \U$3107 ( \3790 , \3787 , \3789 );
and \U$3108 ( \3791 , \2201 , \2856_nGb3b );
and \U$3109 ( \3792 , \2969_nGabe , \2203 );
nor \U$3110 ( \3793 , \3790 , \3791 , \3792 );
and \U$3111 ( \3794 , \2714 , \2532 );
and \U$3112 ( \3795 , \2417 , \2709 );
and \U$3113 ( \3796 , \2621_nGc52 , \2536 );
nor \U$3114 ( \3797 , \3794 , \3795 , \3796 );
xor \U$3115 ( \3798 , \3793 , \3797 );
nand \U$3116 ( \3799 , \3206_nG959 , \1864 );
or \U$3117 ( \3800 , \1810 , \3124_nGa6e );
nand \U$3118 ( \3801 , \3800 , \1959 );
and \U$3119 ( \3802 , \3799 , \3801 );
and \U$3120 ( \3803 , \1954 , \3124_nGa6e );
and \U$3121 ( \3804 , \3206_nG959 , \1866 );
nor \U$3122 ( \3805 , \3802 , \3803 , \3804 );
and \U$3123 ( \3806 , \3798 , \3805 );
and \U$3124 ( \3807 , \3793 , \3797 );
or \U$3125 ( \3808 , \3806 , \3807 );
not \U$3126 ( \3809 , \3808 );
xor \U$3127 ( \3810 , \3786 , \3809 );
xor \U$3128 ( \3811 , \3739 , \3742 );
and \U$3129 ( \3812 , \3810 , \3811 );
and \U$3130 ( \3813 , \3786 , \3809 );
or \U$3131 ( \3814 , \3812 , \3813 );
xor \U$3132 ( \3815 , \3777 , \3814 );
or \U$3133 ( \3816 , \2535 , \3733 );
or \U$3134 ( \3817 , \2969_nGabe , \2419 );
or \U$3135 ( \3818 , \3124_nGa6e , \2418 );
nand \U$3136 ( \3819 , \3816 , \3817 , \3818 );
xor \U$3137 ( \3820 , \3819 , \2103 );
and \U$3138 ( \3821 , \3694 , \2532 );
and \U$3139 ( \3822 , \2417 , \3620 );
and \U$3140 ( \3823 , \3124_nGa6e , \2536 );
nor \U$3141 ( \3824 , \3821 , \3822 , \3823 );
nand \U$3142 ( \3825 , \3206_nG959 , \2418 );
nand \U$3143 ( \3826 , \1965 , \3825 );
nor \U$3144 ( \3827 , \3824 , \3826 );
xor \U$3145 ( \3828 , \3820 , \3827 );
or \U$3146 ( \3829 , \2200 , \3620 );
or \U$3147 ( \3830 , \3206_nG959 , \1970 );
nand \U$3148 ( \3831 , \3829 , \3830 , \2197 );
and \U$3149 ( \3832 , \3828 , \3831 );
and \U$3150 ( \3833 , \3820 , \3827 );
or \U$3151 ( \3834 , \3832 , \3833 );
and \U$3152 ( \3835 , \3819 , \2103 );
xor \U$3153 ( \3836 , \3834 , \3835 );
nand \U$3154 ( \3837 , \3206_nG959 , \2098 );
or \U$3155 ( \3838 , \1970 , \3124_nGa6e );
nand \U$3156 ( \3839 , \3838 , \2197 );
and \U$3157 ( \3840 , \3837 , \3839 );
and \U$3158 ( \3841 , \2201 , \3124_nGa6e );
and \U$3159 ( \3842 , \3206_nG959 , \2203 );
nor \U$3160 ( \3843 , \3840 , \3841 , \3842 );
not \U$3161 ( \3844 , \2856_nGb3b );
and \U$3162 ( \3845 , \3844 , \2532 );
and \U$3163 ( \3846 , \2417 , \3733 );
and \U$3164 ( \3847 , \2856_nGb3b , \2536 );
nor \U$3165 ( \3848 , \3845 , \3846 , \3847 );
and \U$3166 ( \3849 , \3843 , \3848 );
nor \U$3167 ( \3850 , \3843 , \3848 );
nor \U$3168 ( \3851 , \3849 , \3850 );
and \U$3169 ( \3852 , \3836 , \3851 );
and \U$3170 ( \3853 , \3834 , \3835 );
or \U$3171 ( \3854 , \3852 , \3853 );
xor \U$3172 ( \3855 , \3854 , \3850 );
and \U$3173 ( \3856 , \3206_nG959 , \1954 );
and \U$3174 ( \3857 , \3620 , \1811 );
not \U$3175 ( \3858 , \1959 );
nor \U$3176 ( \3859 , \3856 , \3857 , \3858 );
and \U$3177 ( \3860 , \2709 , \2532 );
and \U$3178 ( \3861 , \2417 , \3844 );
and \U$3179 ( \3862 , \2708_nGbb2 , \2536 );
nor \U$3180 ( \3863 , \3860 , \3861 , \3862 );
xor \U$3181 ( \3864 , \1810 , \3863 );
nand \U$3182 ( \3865 , \3124_nGa6e , \2098 );
or \U$3183 ( \3866 , \1970 , \2969_nGabe );
nand \U$3184 ( \3867 , \3866 , \2197 );
and \U$3185 ( \3868 , \3865 , \3867 );
and \U$3186 ( \3869 , \2201 , \2969_nGabe );
and \U$3187 ( \3870 , \3124_nGa6e , \2203 );
nor \U$3188 ( \3871 , \3868 , \3869 , \3870 );
xor \U$3189 ( \3872 , \3864 , \3871 );
and \U$3190 ( \3873 , \3859 , \3872 );
nor \U$3191 ( \3874 , \3859 , \3872 );
nor \U$3192 ( \3875 , \3873 , \3874 );
and \U$3193 ( \3876 , \3855 , \3875 );
and \U$3194 ( \3877 , \3854 , \3850 );
or \U$3195 ( \3878 , \3876 , \3877 );
xor \U$3196 ( \3879 , \3878 , \3874 );
xor \U$3197 ( \3880 , \3793 , \3797 );
xor \U$3198 ( \3881 , \3880 , \3805 );
xor \U$3199 ( \3882 , \1810 , \3863 );
and \U$3200 ( \3883 , \3882 , \3871 );
and \U$3201 ( \3884 , \1810 , \3863 );
or \U$3202 ( \3885 , \3883 , \3884 );
and \U$3203 ( \3886 , \3881 , \3885 );
nor \U$3204 ( \3887 , \3881 , \3885 );
nor \U$3205 ( \3888 , \3886 , \3887 );
and \U$3206 ( \3889 , \3879 , \3888 );
and \U$3207 ( \3890 , \3878 , \3874 );
or \U$3208 ( \3891 , \3889 , \3890 );
xor \U$3209 ( \3892 , \3891 , \3887 );
xor \U$3210 ( \3893 , \3786 , \3809 );
xor \U$3211 ( \3894 , \3893 , \3811 );
and \U$3212 ( \3895 , \3892 , \3894 );
and \U$3213 ( \3896 , \3891 , \3887 );
or \U$3214 ( \3897 , \3895 , \3896 );
and \U$3215 ( \3898 , \3815 , \3897 );
and \U$3216 ( \3899 , \3777 , \3814 );
or \U$3217 ( \3900 , \3898 , \3899 );
and \U$3218 ( \3901 , \3731 , \3776 );
xor \U$3219 ( \3902 , \3900 , \3901 );
xor \U$3220 ( \3903 , \3656 , \3660 );
xor \U$3221 ( \3904 , \3903 , \1425 );
xor \U$3222 ( \3905 , \3717 , \3721 );
and \U$3223 ( \3906 , \3905 , \3729 );
and \U$3224 ( \3907 , \3717 , \3721 );
or \U$3225 ( \3908 , \3906 , \3907 );
xor \U$3226 ( \3909 , \3672 , \3679 );
xor \U$3227 ( \3910 , \3909 , \3684 );
xor \U$3228 ( \3911 , \3908 , \3910 );
xor \U$3229 ( \3912 , \3904 , \3911 );
and \U$3230 ( \3913 , \3771 , \3743 );
nor \U$3231 ( \3914 , \3913 , \3769 );
and \U$3232 ( \3915 , \3912 , \3914 );
nor \U$3233 ( \3916 , \3912 , \3914 );
nor \U$3234 ( \3917 , \3915 , \3916 );
and \U$3235 ( \3918 , \3902 , \3917 );
and \U$3236 ( \3919 , \3900 , \3901 );
or \U$3237 ( \3920 , \3918 , \3919 );
not \U$3238 ( \3921 , \3916 );
xor \U$3239 ( \3922 , \3649 , \3664 );
xor \U$3240 ( \3923 , \3922 , \3687 );
not \U$3241 ( \3924 , \3701 );
not \U$3242 ( \3925 , \3704 );
and \U$3243 ( \3926 , \3924 , \3925 );
and \U$3244 ( \3927 , \3701 , \3704 );
nor \U$3245 ( \3928 , \3926 , \3927 );
xor \U$3246 ( \3929 , \3656 , \3660 );
xor \U$3247 ( \3930 , \3929 , \1425 );
and \U$3248 ( \3931 , \3908 , \3930 );
xor \U$3249 ( \3932 , \3656 , \3660 );
xor \U$3250 ( \3933 , \3932 , \1425 );
and \U$3251 ( \3934 , \3910 , \3933 );
and \U$3252 ( \3935 , \3908 , \3910 );
or \U$3253 ( \3936 , \3931 , \3934 , \3935 );
xor \U$3254 ( \3937 , \3928 , \3936 );
xor \U$3255 ( \3938 , \3923 , \3937 );
nor \U$3256 ( \3939 , \3921 , \3938 );
or \U$3257 ( \3940 , \3920 , \3939 );
not \U$3258 ( \3941 , \3916 );
nand \U$3259 ( \3942 , \3941 , \3938 );
nand \U$3260 ( \3943 , \3940 , \3942 );
not \U$3261 ( \3944 , \3943 );
xor \U$3262 ( \3945 , \3534 , \3541 );
xor \U$3263 ( \3946 , \3945 , \3549 );
xor \U$3264 ( \3947 , \3615 , \3623 );
xor \U$3265 ( \3948 , \3946 , \3947 );
not \U$3266 ( \3949 , \3948 );
not \U$3267 ( \3950 , \3705 );
not \U$3268 ( \3951 , \3707 );
nand \U$3269 ( \3952 , \3951 , \3693 );
not \U$3270 ( \3953 , \3952 );
or \U$3271 ( \3954 , \3950 , \3953 );
or \U$3272 ( \3955 , \3952 , \3705 );
nand \U$3273 ( \3956 , \3954 , \3955 );
not \U$3274 ( \3957 , \3956 );
and \U$3275 ( \3958 , \3949 , \3957 );
and \U$3276 ( \3959 , \3948 , \3956 );
nor \U$3277 ( \3960 , \3958 , \3959 );
xor \U$3278 ( \3961 , \3649 , \3664 );
xor \U$3279 ( \3962 , \3961 , \3687 );
and \U$3280 ( \3963 , \3928 , \3962 );
xor \U$3281 ( \3964 , \3649 , \3664 );
xor \U$3282 ( \3965 , \3964 , \3687 );
and \U$3283 ( \3966 , \3936 , \3965 );
and \U$3284 ( \3967 , \3928 , \3936 );
or \U$3285 ( \3968 , \3963 , \3966 , \3967 );
and \U$3286 ( \3969 , \3960 , \3968 );
not \U$3287 ( \3970 , \3969 );
and \U$3288 ( \3971 , \3944 , \3970 );
nor \U$3289 ( \3972 , \3960 , \3968 );
nor \U$3290 ( \3973 , \3971 , \3972 );
not \U$3291 ( \3974 , \3973 );
not \U$3292 ( \3975 , \3956 );
nor \U$3293 ( \3976 , \3975 , \3948 );
xor \U$3294 ( \3977 , \3974 , \3976 );
and \U$3295 ( \3978 , \3642 , \3708 );
nor \U$3296 ( \3979 , \3978 , \3709 );
and \U$3297 ( \3980 , \3977 , \3979 );
and \U$3298 ( \3981 , \3974 , \3976 );
or \U$3299 ( \3982 , \3980 , \3981 );
and \U$3300 ( \3983 , \3710 , \3982 );
and \U$3301 ( \3984 , \3640 , \3709 );
or \U$3302 ( \3985 , \3983 , \3984 );
and \U$3303 ( \3986 , \3638 , \3985 );
and \U$3304 ( \3987 , \3590 , \3637 );
or \U$3305 ( \3988 , \3986 , \3987 );
xor \U$3306 ( \3989 , \3584 , \3586 );
and \U$3307 ( \3990 , \3989 , \3588 );
and \U$3308 ( \3991 , \3584 , \3586 );
or \U$3309 ( \3992 , \3990 , \3991 );
xor \U$3310 ( \3993 , \3441 , \3520 );
xor \U$3311 ( \3994 , \3993 , \3523 );
nand \U$3312 ( \3995 , \3992 , \3994 );
and \U$3313 ( \3996 , \3988 , \3995 );
nor \U$3314 ( \3997 , \3994 , \3992 );
nor \U$3315 ( \3998 , \3996 , \3997 );
and \U$3316 ( \3999 , \3527 , \3998 );
and \U$3317 ( \4000 , \3436 , \3526 );
or \U$3318 ( \4001 , \3999 , \4000 );
not \U$3319 ( \4002 , \4001 );
and \U$3320 ( \4003 , \3429 , \4002 );
and \U$3321 ( \4004 , \3353 , \3428 );
or \U$3322 ( \4005 , \4003 , \4004 );
and \U$3323 ( \4006 , \3351 , \4005 );
and \U$3324 ( \4007 , \3268 , \3350 );
or \U$3325 ( \4008 , \4006 , \4007 );
and \U$3326 ( \4009 , \3266 , \4008 );
and \U$3327 ( \4010 , \3252 , \3265 );
or \U$3328 ( \4011 , \4009 , \4010 );
and \U$3329 ( \4012 , \3250 , \4011 );
and \U$3330 ( \4013 , \3080 , \3249 );
or \U$3331 ( \4014 , \4012 , \4013 );
and \U$3332 ( \4015 , \3078 , \4014 );
and \U$3333 ( \4016 , \2997 , \3077 );
or \U$3334 ( \4017 , \4015 , \4016 );
and \U$3335 ( \4018 , \2995 , \4017 );
and \U$3336 ( \4019 , \2825 , \2994 );
or \U$3337 ( \4020 , \4018 , \4019 );
and \U$3338 ( \4021 , \2823 , \4020 );
and \U$3339 ( \4022 , \2820 , \2822 );
or \U$3340 ( \4023 , \4021 , \4022 );
and \U$3341 ( \4024 , \2749 , \4023 );
and \U$3342 ( \4025 , \2746 , \2748 );
or \U$3343 ( \4026 , \4024 , \4025 );
and \U$3344 ( \4027 , \2584 , \4026 );
and \U$3345 ( \4028 , \2470 , \2583 );
or \U$3346 ( \4029 , \4027 , \4028 );
not \U$3347 ( \4030 , \2457 );
not \U$3348 ( \4031 , \2466 );
and \U$3349 ( \4032 , \4030 , \4031 );
nor \U$3350 ( \4033 , \4032 , \2456 );
not \U$3351 ( \4034 , \2298 );
not \U$3352 ( \4035 , \2292 );
nand \U$3353 ( \4036 , \4035 , \2300 );
not \U$3354 ( \4037 , \4036 );
or \U$3355 ( \4038 , \4034 , \4037 );
or \U$3356 ( \4039 , \4036 , \2298 );
nand \U$3357 ( \4040 , \4038 , \4039 );
nand \U$3358 ( \4041 , \4033 , \4040 );
and \U$3359 ( \4042 , \4029 , \4041 );
nor \U$3360 ( \4043 , \4040 , \4033 );
nor \U$3361 ( \4044 , \4042 , \4043 );
not \U$3362 ( \4045 , \4044 );
and \U$3363 ( \4046 , \2302 , \4045 );
and \U$3364 ( \4047 , \2163 , \2301 );
or \U$3365 ( \4048 , \4046 , \4047 );
and \U$3366 ( \4049 , \2161 , \4048 );
and \U$3367 ( \4050 , \2156 , \2160 );
or \U$3368 ( \4051 , \4049 , \4050 );
and \U$3369 ( \4052 , \2049 , \4051 );
and \U$3370 ( \4053 , \1940 , \2048 );
or \U$3371 ( \4054 , \4052 , \4053 );
and \U$3372 ( \4055 , \1938 , \4054 );
and \U$3373 ( \4056 , \1935 , \1937 );
or \U$3374 ( \4057 , \4055 , \4056 );
and \U$3375 ( \4058 , \1850 , \4057 );
and \U$3376 ( \4059 , \1743 , \1849 );
or \U$3377 ( \4060 , \4058 , \4059 );
and \U$3378 ( \4061 , \1741 , \4060 );
and \U$3379 ( \4062 , \1569 , \1740 );
or \U$3380 ( \4063 , \4061 , \4062 );
and \U$3381 ( \4064 , \1567 , \4063 );
and \U$3382 ( \4065 , \1565 , \1566 );
or \U$3383 ( \4066 , \4064 , \4065 );
not \U$3384 ( \4067 , \4066 );
or \U$3385 ( \4068 , \1459 , \4067 );
or \U$3386 ( \4069 , \4066 , \1458 );
nand \U$3387 ( \4070 , \4068 , \4069 );
and \U$3388 ( \4071 , \734 , RIb551908_250);
and \U$3389 ( \4072 , \703 , RIb551c50_257);
and \U$3390 ( \4073 , RIb551bd8_256, \705 );
nor \U$3391 ( \4074 , \4072 , \4073 );
and \U$3392 ( \4075 , \716 , RIb551e30_261);
and \U$3393 ( \4076 , RIb551ea8_262, \713 );
nor \U$3394 ( \4077 , \4075 , \4076 );
and \U$3395 ( \4078 , \710 , RIb551f20_263);
and \U$3396 ( \4079 , RIb551cc8_258, \698 );
nor \U$3397 ( \4080 , \4078 , \4079 );
and \U$3398 ( \4081 , \690 , RIb551b60_255);
and \U$3399 ( \4082 , RIb551ae8_254, \726 );
nor \U$3400 ( \4083 , \4081 , \4082 );
nand \U$3401 ( \4084 , \4074 , \4077 , \4080 , \4083 );
not \U$3402 ( \4085 , \733 );
nor \U$3403 ( \4086 , \4071 , \4084 , \4085 );
and \U$3404 ( \4087 , \738 , RIb551980_251);
and \U$3405 ( \4088 , RIb5519f8_252, \740 );
nor \U$3406 ( \4089 , \4087 , \4088 );
and \U$3407 ( \4090 , \695 , RIb551d40_259);
and \U$3408 ( \4091 , RIb551db8_260, \719 );
nor \U$3409 ( \4092 , \4090 , \4091 );
and \U$3410 ( \4093 , \724 , RIb551a70_253);
not \U$3411 ( \4094 , \679 );
nor \U$3412 ( \4095 , \4094 , \682 );
and \U$3413 ( \4096 , RIb551890_249, \4095 );
nor \U$3414 ( \4097 , \4093 , \4096 );
nand \U$3415 ( \4098 , \4086 , \4089 , \4092 , \4097 );
buf \U$3416 ( \4099 , \4098 );
buf \U$3417 ( \4100 , \750 );
_DC g11f9 ( \4101_nG11f9 , \4099 , \4100 );
xor \U$3418 ( \4102 , \673 , \4101_nG11f9 );
and \U$3419 ( \4103 , \724 , RIb54ae28_22);
and \U$3420 ( \4104 , \716 , RIb54b1e8_30);
and \U$3421 ( \4105 , RIb54ad38_20, \738 );
nor \U$3422 ( \4106 , \4104 , \4105 );
and \U$3423 ( \4107 , \740 , RIb54adb0_21);
and \U$3424 ( \4108 , RIb54acc0_19, \734 );
nor \U$3425 ( \4109 , \4107 , \4108 );
and \U$3426 ( \4110 , \710 , RIb54b2d8_32);
and \U$3427 ( \4111 , RIb54b260_31, \713 );
nor \U$3428 ( \4112 , \4110 , \4111 );
and \U$3429 ( \4113 , \690 , RIb54af18_24);
and \U$3430 ( \4114 , RIb54aea0_23, \726 );
nor \U$3431 ( \4115 , \4113 , \4114 );
nand \U$3432 ( \4116 , \4106 , \4109 , \4112 , \4115 );
not \U$3433 ( \4117 , \778 );
nor \U$3434 ( \4118 , \4103 , \4116 , \4117 );
and \U$3435 ( \4119 , \695 , RIb54b0f8_28);
and \U$3436 ( \4120 , RIb54b170_29, \719 );
nor \U$3437 ( \4121 , \4119 , \4120 );
and \U$3438 ( \4122 , \698 , RIb54b080_27);
and \U$3439 ( \4123 , RIb54ac48_18, \4095 );
nor \U$3440 ( \4124 , \4122 , \4123 );
and \U$3441 ( \4125 , \703 , RIb54b008_26);
and \U$3442 ( \4126 , RIb54af90_25, \705 );
nor \U$3443 ( \4127 , \4125 , \4126 );
nand \U$3444 ( \4128 , \4118 , \4121 , \4124 , \4127 );
buf \U$3445 ( \4129 , \4128 );
_DC g1010 ( \4130_nG1010 , \4129 , \4100 );
xor \U$3446 ( \4131 , \758 , \4130_nG1010 );
and \U$3447 ( \4132 , \690 , RIb54b710_41);
and \U$3448 ( \4133 , \738 , RIb54b530_37);
and \U$3449 ( \4134 , RIb54b5a8_38, \740 );
nor \U$3450 ( \4135 , \4133 , \4134 );
and \U$3451 ( \4136 , \716 , RIb54b9e0_47);
and \U$3452 ( \4137 , RIb54b4b8_36, \734 );
nor \U$3453 ( \4138 , \4136 , \4137 );
and \U$3454 ( \4139 , \710 , RIb54bad0_49);
and \U$3455 ( \4140 , RIb54ba58_48, \713 );
nor \U$3456 ( \4141 , \4139 , \4140 );
and \U$3457 ( \4142 , \724 , RIb54b620_39);
and \U$3458 ( \4143 , RIb54b698_40, \726 );
nor \U$3459 ( \4144 , \4142 , \4143 );
nand \U$3460 ( \4145 , \4135 , \4138 , \4141 , \4144 );
not \U$3461 ( \4146 , \814 );
nor \U$3462 ( \4147 , \4132 , \4145 , \4146 );
and \U$3463 ( \4148 , \695 , RIb54b8f0_45);
and \U$3464 ( \4149 , RIb54b968_46, \719 );
nor \U$3465 ( \4150 , \4148 , \4149 );
and \U$3466 ( \4151 , \698 , RIb54b878_44);
and \U$3467 ( \4152 , RIb54b440_35, \4095 );
nor \U$3468 ( \4153 , \4151 , \4152 );
and \U$3469 ( \4154 , \703 , RIb54b800_43);
and \U$3470 ( \4155 , RIb54b788_42, \705 );
nor \U$3471 ( \4156 , \4154 , \4155 );
nand \U$3472 ( \4157 , \4147 , \4150 , \4153 , \4156 );
buf \U$3473 ( \4158 , \4157 );
_DC g100e ( \4159_nG100e , \4158 , \4100 );
xor \U$3474 ( \4160 , \794 , \4159_nG100e );
and \U$3475 ( \4161 , RIb54c250_65, \713 );
and \U$3476 ( \4162 , RIb54bd28_54, \738 );
and \U$3477 ( \4163 , \726 , RIb54be90_57);
and \U$3478 ( \4164 , RIb54bcb0_53, \734 );
nor \U$3479 ( \4165 , \4163 , \4164 );
and \U$3480 ( \4166 , RIb54be18_56, \724 );
and \U$3481 ( \4167 , \740 , RIb54bda0_55);
and \U$3482 ( \4168 , RIb54bf08_58, \690 );
nor \U$3483 ( \4169 , \4166 , \4167 , \4168 );
and \U$3484 ( \4170 , \710 , RIb54c2c8_66);
and \U$3485 ( \4171 , RIb54bc38_52, \4095 );
nor \U$3486 ( \4172 , \4170 , \4171 );
nand \U$3487 ( \4173 , \4165 , \4169 , \4172 );
nor \U$3488 ( \4174 , \4161 , \4162 , \4173 );
and \U$3489 ( \4175 , \716 , RIb54c1d8_64);
and \U$3490 ( \4176 , RIb54c160_63, \719 );
nor \U$3491 ( \4177 , \4175 , \4176 );
and \U$3492 ( \4178 , RIb54c0e8_62, \695 );
and \U$3493 ( \4179 , RIb54c070_61, \698 );
and \U$3494 ( \4180 , \703 , RIb54bff8_60);
and \U$3495 ( \4181 , RIb54bf80_59, \705 );
nor \U$3496 ( \4182 , \4180 , \4181 );
not \U$3497 ( \4183 , \4182 );
nor \U$3498 ( \4184 , \4178 , \4179 , \4183 );
nand \U$3499 ( \4185 , \4174 , \4177 , \846 , \4184 );
buf \U$3500 ( \4186 , \4185 );
_DC ge60 ( \4187_nGe60 , \4186 , \4100 );
xor \U$3501 ( \4188 , \830 , \4187_nGe60 );
and \U$3502 ( \4189 , \4095 , RIb54c430_69);
and \U$3503 ( \4190 , \703 , RIb54c7f0_77);
and \U$3504 ( \4191 , RIb54c778_76, \705 );
nor \U$3505 ( \4192 , \4190 , \4191 );
and \U$3506 ( \4193 , \690 , RIb54c700_75);
and \U$3507 ( \4194 , RIb54c688_74, \726 );
nor \U$3508 ( \4195 , \4193 , \4194 );
and \U$3509 ( \4196 , \710 , RIb54cac0_83);
and \U$3510 ( \4197 , RIb54c868_78, \698 );
nor \U$3511 ( \4198 , \4196 , \4197 );
and \U$3512 ( \4199 , \716 , RIb54c9d0_81);
and \U$3513 ( \4200 , RIb54ca48_82, \713 );
nor \U$3514 ( \4201 , \4199 , \4200 );
nand \U$3515 ( \4202 , \4192 , \4195 , \4198 , \4201 );
and \U$3516 ( \4203 , \738 , RIb54c520_71);
and \U$3517 ( \4204 , RIb54c4a8_70, \734 );
nor \U$3518 ( \4205 , \4203 , \4204 );
not \U$3519 ( \4206 , \4205 );
nor \U$3520 ( \4207 , \4189 , \4202 , \4206 );
and \U$3521 ( \4208 , \695 , RIb54c8e0_79);
and \U$3522 ( \4209 , RIb54c958_80, \719 );
nor \U$3523 ( \4210 , \4208 , \4209 );
and \U$3524 ( \4211 , \724 , RIb54c610_73);
and \U$3525 ( \4212 , RIb54c598_72, \740 );
nor \U$3526 ( \4213 , \4211 , \4212 );
nand \U$3527 ( \4214 , \4207 , \4210 , \884 , \4213 );
buf \U$3528 ( \4215 , \4214 );
_DC ge5e ( \4216_nGe5e , \4215 , \4100 );
xor \U$3529 ( \4217 , \866 , \4216_nGe5e );
and \U$3530 ( \4218 , \4095 , RIb54cc28_86);
and \U$3531 ( \4219 , \703 , RIb54cfe8_94);
and \U$3532 ( \4220 , RIb54d060_95, \698 );
nor \U$3533 ( \4221 , \4219 , \4220 );
and \U$3534 ( \4222 , \695 , RIb54d0d8_96);
and \U$3535 ( \4223 , RIb54d150_97, \719 );
nor \U$3536 ( \4224 , \4222 , \4223 );
and \U$3537 ( \4225 , \716 , RIb54d1c8_98);
and \U$3538 ( \4226 , RIb54d240_99, \713 );
nor \U$3539 ( \4227 , \4225 , \4226 );
and \U$3540 ( \4228 , \690 , RIb54cef8_92);
and \U$3541 ( \4229 , RIb54cf70_93, \705 );
nor \U$3542 ( \4230 , \4228 , \4229 );
nand \U$3543 ( \4231 , \4221 , \4224 , \4227 , \4230 );
and \U$3544 ( \4232 , \738 , RIb54cd18_88);
and \U$3545 ( \4233 , RIb54cca0_87, \734 );
nor \U$3546 ( \4234 , \4232 , \4233 );
not \U$3547 ( \4235 , \4234 );
nor \U$3548 ( \4236 , \4218 , \4231 , \4235 );
and \U$3549 ( \4237 , \710 , RIb54d2b8_100);
and \U$3550 ( \4238 , RIb54ce80_91, \726 );
nor \U$3551 ( \4239 , \4237 , \4238 );
and \U$3552 ( \4240 , \724 , RIb54ce08_90);
and \U$3553 ( \4241 , RIb54cd90_89, \740 );
nor \U$3554 ( \4242 , \4240 , \4241 );
nand \U$3555 ( \4243 , \4236 , \4239 , \920 , \4242 );
buf \U$3556 ( \4244 , \4243 );
_DC gce3 ( \4245_nGce3 , \4244 , \4100 );
xor \U$3557 ( \4246 , \904 , \4245_nGce3 );
and \U$3558 ( \4247 , RIb54da38_116, \713 );
and \U$3559 ( \4248 , RIb54d6f0_109, \690 );
and \U$3560 ( \4249 , \724 , RIb54d600_107);
and \U$3561 ( \4250 , RIb54d588_106, \740 );
nor \U$3562 ( \4251 , \4249 , \4250 );
and \U$3563 ( \4252 , RIb54d510_105, \738 );
and \U$3564 ( \4253 , \734 , RIb54d498_104);
and \U$3565 ( \4254 , RIb54d678_108, \726 );
nor \U$3566 ( \4255 , \4252 , \4253 , \4254 );
and \U$3567 ( \4256 , \710 , RIb54dab0_117);
and \U$3568 ( \4257 , RIb54d420_103, \4095 );
nor \U$3569 ( \4258 , \4256 , \4257 );
nand \U$3570 ( \4259 , \4251 , \4255 , \4258 );
nor \U$3571 ( \4260 , \4247 , \4248 , \4259 );
and \U$3572 ( \4261 , \716 , RIb54d9c0_115);
and \U$3573 ( \4262 , RIb54d948_114, \719 );
nor \U$3574 ( \4263 , \4261 , \4262 );
and \U$3575 ( \4264 , RIb54d8d0_113, \695 );
and \U$3576 ( \4265 , RIb54d858_112, \698 );
and \U$3577 ( \4266 , \703 , RIb54d7e0_111);
and \U$3578 ( \4267 , RIb54d768_110, \705 );
nor \U$3579 ( \4268 , \4266 , \4267 );
not \U$3580 ( \4269 , \4268 );
nor \U$3581 ( \4270 , \4264 , \4265 , \4269 );
nand \U$3582 ( \4271 , \4260 , \4263 , \946 , \4270 );
buf \U$3583 ( \4272 , \4271 );
_DC gce1 ( \4273_nGce1 , \4272 , \4100 );
xor \U$3584 ( \4274 , \940 , \4273_nGce1 );
and \U$3585 ( \4275 , RIb54dc18_120, \4095 );
and \U$3586 ( \4276 , RIb54e2a8_134, \710 );
and \U$3587 ( \4277 , \703 , RIb54dfd8_128);
and \U$3588 ( \4278 , RIb54e050_129, \698 );
nor \U$3589 ( \4279 , \4277 , \4278 );
and \U$3590 ( \4280 , \695 , RIb54e0c8_130);
and \U$3591 ( \4281 , RIb54e140_131, \719 );
nor \U$3592 ( \4282 , \4280 , \4281 );
and \U$3593 ( \4283 , \716 , RIb54e1b8_132);
and \U$3594 ( \4284 , RIb54e230_133, \713 );
nor \U$3595 ( \4285 , \4283 , \4284 );
and \U$3596 ( \4286 , \690 , RIb54dee8_126);
and \U$3597 ( \4287 , RIb54df60_127, \705 );
nor \U$3598 ( \4288 , \4286 , \4287 );
nand \U$3599 ( \4289 , \4279 , \4282 , \4285 , \4288 );
nor \U$3600 ( \4290 , \4275 , \4276 , \4289 );
and \U$3601 ( \4291 , \738 , RIb54dd08_122);
and \U$3602 ( \4292 , RIb54dc90_121, \734 );
nor \U$3603 ( \4293 , \4291 , \4292 );
and \U$3604 ( \4294 , \726 , RIb54de70_125);
not \U$3605 ( \4295 , \1002 );
nor \U$3606 ( \4296 , \4294 , \4295 );
and \U$3607 ( \4297 , \724 , RIb54ddf8_124);
and \U$3608 ( \4298 , RIb54dd80_123, \740 );
nor \U$3609 ( \4299 , \4297 , \4298 );
nand \U$3610 ( \4300 , \4290 , \4293 , \4296 , \4299 );
buf \U$3611 ( \4301 , \4300 );
_DC gbb6 ( \4302_nGbb6 , \4301 , \4100 );
xor \U$3612 ( \4303 , \978 , \4302_nGbb6 );
and \U$3613 ( \4304 , \734 , RIb54e488_138);
and \U$3614 ( \4305 , \703 , RIb54e7d0_145);
and \U$3615 ( \4306 , RIb54e758_144, \705 );
nor \U$3616 ( \4307 , \4305 , \4306 );
and \U$3617 ( \4308 , \716 , RIb54e9b0_149);
and \U$3618 ( \4309 , RIb54e848_146, \698 );
nor \U$3619 ( \4310 , \4308 , \4309 );
and \U$3620 ( \4311 , \710 , RIb54eaa0_151);
and \U$3621 ( \4312 , RIb54ea28_150, \713 );
nor \U$3622 ( \4313 , \4311 , \4312 );
and \U$3623 ( \4314 , \690 , RIb54e6e0_143);
and \U$3624 ( \4315 , RIb54e668_142, \726 );
nor \U$3625 ( \4316 , \4314 , \4315 );
nand \U$3626 ( \4317 , \4307 , \4310 , \4313 , \4316 );
not \U$3627 ( \4318 , \1034 );
nor \U$3628 ( \4319 , \4304 , \4317 , \4318 );
and \U$3629 ( \4320 , \738 , RIb54e500_139);
and \U$3630 ( \4321 , RIb54e578_140, \740 );
nor \U$3631 ( \4322 , \4320 , \4321 );
and \U$3632 ( \4323 , \695 , RIb54e8c0_147);
and \U$3633 ( \4324 , RIb54e938_148, \719 );
nor \U$3634 ( \4325 , \4323 , \4324 );
and \U$3635 ( \4326 , \724 , RIb54e5f0_141);
and \U$3636 ( \4327 , RIb54e410_137, \4095 );
nor \U$3637 ( \4328 , \4326 , \4327 );
nand \U$3638 ( \4329 , \4319 , \4322 , \4325 , \4328 );
buf \U$3639 ( \4330 , \4329 );
_DC gbb4 ( \4331_nGbb4 , \4330 , \4100 );
xor \U$3640 ( \4332 , \1014 , \4331_nGbb4 );
and \U$3641 ( \4333 , \734 , RIb54ec80_155);
and \U$3642 ( \4334 , \703 , RIb54efc8_162);
and \U$3643 ( \4335 , RIb54ef50_161, \705 );
nor \U$3644 ( \4336 , \4334 , \4335 );
and \U$3645 ( \4337 , \716 , RIb54f1a8_166);
and \U$3646 ( \4338 , RIb54f220_167, \713 );
nor \U$3647 ( \4339 , \4337 , \4338 );
and \U$3648 ( \4340 , \710 , RIb54f298_168);
and \U$3649 ( \4341 , RIb54f040_163, \698 );
nor \U$3650 ( \4342 , \4340 , \4341 );
and \U$3651 ( \4343 , \690 , RIb54eed8_160);
and \U$3652 ( \4344 , RIb54ee60_159, \726 );
nor \U$3653 ( \4345 , \4343 , \4344 );
nand \U$3654 ( \4346 , \4336 , \4339 , \4342 , \4345 );
not \U$3655 ( \4347 , \1066 );
nor \U$3656 ( \4348 , \4333 , \4346 , \4347 );
and \U$3657 ( \4349 , \738 , RIb54ecf8_156);
and \U$3658 ( \4350 , RIb54ed70_157, \740 );
nor \U$3659 ( \4351 , \4349 , \4350 );
and \U$3660 ( \4352 , \695 , RIb54f0b8_164);
and \U$3661 ( \4353 , RIb54f130_165, \719 );
nor \U$3662 ( \4354 , \4352 , \4353 );
and \U$3663 ( \4355 , \724 , RIb54ede8_158);
and \U$3664 ( \4356 , RIb54ec08_154, \4095 );
nor \U$3665 ( \4357 , \4355 , \4356 );
nand \U$3666 ( \4358 , \4348 , \4351 , \4354 , \4357 );
buf \U$3667 ( \4359 , \4358 );
_DC gade ( \4360_nGade , \4359 , \4100 );
xor \U$3668 ( \4361 , \1046 , \4360_nGade );
and \U$3669 ( \4362 , \734 , RIb54f478_172);
and \U$3670 ( \4363 , \703 , RIb54f7c0_179);
and \U$3671 ( \4364 , RIb54f748_178, \705 );
nor \U$3672 ( \4365 , \4363 , \4364 );
and \U$3673 ( \4366 , \716 , RIb54f9a0_183);
and \U$3674 ( \4367 , RIb54fa18_184, \713 );
nor \U$3675 ( \4368 , \4366 , \4367 );
and \U$3676 ( \4369 , \710 , RIb54fa90_185);
and \U$3677 ( \4370 , RIb54f838_180, \698 );
nor \U$3678 ( \4371 , \4369 , \4370 );
and \U$3679 ( \4372 , \690 , RIb54f6d0_177);
and \U$3680 ( \4373 , RIb54f658_176, \726 );
nor \U$3681 ( \4374 , \4372 , \4373 );
nand \U$3682 ( \4375 , \4365 , \4368 , \4371 , \4374 );
not \U$3683 ( \4376 , \1098 );
nor \U$3684 ( \4377 , \4362 , \4375 , \4376 );
and \U$3685 ( \4378 , \738 , RIb54f4f0_173);
and \U$3686 ( \4379 , RIb54f568_174, \740 );
nor \U$3687 ( \4380 , \4378 , \4379 );
and \U$3688 ( \4381 , \695 , RIb54f8b0_181);
and \U$3689 ( \4382 , RIb54f928_182, \719 );
nor \U$3690 ( \4383 , \4381 , \4382 );
and \U$3691 ( \4384 , \724 , RIb54f5e0_175);
and \U$3692 ( \4385 , RIb54f400_171, \4095 );
nor \U$3693 ( \4386 , \4384 , \4385 );
nand \U$3694 ( \4387 , \4377 , \4380 , \4383 , \4386 );
buf \U$3695 ( \4388 , \4387 );
_DC gae0 ( \4389_nGae0 , \4388 , \4100 );
xor \U$3696 ( \4390 , \1078 , \4389_nGae0 );
and \U$3697 ( \4391 , \734 , RIb54fc70_189);
and \U$3698 ( \4392 , \703 , RIb54ffb8_196);
and \U$3699 ( \4393 , RIb54ff40_195, \705 );
nor \U$3700 ( \4394 , \4392 , \4393 );
and \U$3701 ( \4395 , \690 , RIb54fec8_194);
and \U$3702 ( \4396 , RIb54fe50_193, \726 );
nor \U$3703 ( \4397 , \4395 , \4396 );
and \U$3704 ( \4398 , \710 , RIb550288_202);
and \U$3705 ( \4399 , RIb550030_197, \698 );
nor \U$3706 ( \4400 , \4398 , \4399 );
and \U$3707 ( \4401 , \716 , RIb550198_200);
and \U$3708 ( \4402 , RIb550210_201, \713 );
nor \U$3709 ( \4403 , \4401 , \4402 );
nand \U$3710 ( \4404 , \4394 , \4397 , \4400 , \4403 );
not \U$3711 ( \4405 , \1129 );
nor \U$3712 ( \4406 , \4391 , \4404 , \4405 );
and \U$3713 ( \4407 , \738 , RIb54fce8_190);
and \U$3714 ( \4408 , RIb54fd60_191, \740 );
nor \U$3715 ( \4409 , \4407 , \4408 );
and \U$3716 ( \4410 , \695 , RIb5500a8_198);
and \U$3717 ( \4411 , RIb550120_199, \719 );
nor \U$3718 ( \4412 , \4410 , \4411 );
and \U$3719 ( \4413 , \724 , RIb54fdd8_192);
and \U$3720 ( \4414 , RIb54fbf8_188, \4095 );
nor \U$3721 ( \4415 , \4413 , \4414 );
nand \U$3722 ( \4416 , \4406 , \4409 , \4412 , \4415 );
buf \U$3723 ( \4417 , \4416 );
_DC g97f ( \4418_nG97f , \4417 , \4100 );
xor \U$3724 ( \4419 , RIb54a900_11, \4418_nG97f );
and \U$3725 ( \4420 , RIb550a80_219, \713 );
and \U$3726 ( \4421 , RIb550738_212, \690 );
and \U$3727 ( \4422 , \724 , RIb550648_210);
and \U$3728 ( \4423 , RIb5505d0_209, \740 );
nor \U$3729 ( \4424 , \4422 , \4423 );
and \U$3730 ( \4425 , RIb550558_208, \738 );
and \U$3731 ( \4426 , \734 , RIb5504e0_207);
and \U$3732 ( \4427 , RIb5506c0_211, \726 );
nor \U$3733 ( \4428 , \4425 , \4426 , \4427 );
and \U$3734 ( \4429 , \710 , RIb550af8_220);
and \U$3735 ( \4430 , RIb550468_206, \4095 );
nor \U$3736 ( \4431 , \4429 , \4430 );
nand \U$3737 ( \4432 , \4424 , \4428 , \4431 );
nor \U$3738 ( \4433 , \4420 , \4421 , \4432 );
and \U$3739 ( \4434 , \716 , RIb550a08_218);
and \U$3740 ( \4435 , RIb550990_217, \719 );
nor \U$3741 ( \4436 , \4434 , \4435 );
and \U$3742 ( \4437 , RIb550918_216, \695 );
and \U$3743 ( \4438 , RIb5508a0_215, \698 );
and \U$3744 ( \4439 , \703 , RIb550828_214);
and \U$3745 ( \4440 , RIb5507b0_213, \705 );
nor \U$3746 ( \4441 , \4439 , \4440 );
not \U$3747 ( \4442 , \4441 );
nor \U$3748 ( \4443 , \4437 , \4438 , \4442 );
nand \U$3749 ( \4444 , \4433 , \4436 , \1146 , \4443 );
buf \U$3750 ( \4445 , \4444 );
_DC g97d ( \4446_nG97d , \4445 , \4100 );
nand \U$3751 ( \4447 , \4446_nG97d , \1173 );
not \U$3752 ( \4448 , \4447 );
and \U$3753 ( \4449 , \4419 , \4448 );
and \U$3754 ( \4450 , RIb54a900_11, \4418_nG97f );
or \U$3755 ( \4451 , \4449 , \4450 );
and \U$3756 ( \4452 , \4390 , \4451 );
and \U$3757 ( \4453 , \1078 , \4389_nGae0 );
or \U$3758 ( \4454 , \4452 , \4453 );
and \U$3759 ( \4455 , \4361 , \4454 );
and \U$3760 ( \4456 , \1046 , \4360_nGade );
or \U$3761 ( \4457 , \4455 , \4456 );
and \U$3762 ( \4458 , \4332 , \4457 );
and \U$3763 ( \4459 , \1014 , \4331_nGbb4 );
or \U$3764 ( \4460 , \4458 , \4459 );
and \U$3765 ( \4461 , \4303 , \4460 );
and \U$3766 ( \4462 , \978 , \4302_nGbb6 );
or \U$3767 ( \4463 , \4461 , \4462 );
and \U$3768 ( \4464 , \4274 , \4463 );
and \U$3769 ( \4465 , \940 , \4273_nGce1 );
or \U$3770 ( \4466 , \4464 , \4465 );
and \U$3771 ( \4467 , \4246 , \4466 );
and \U$3772 ( \4468 , \904 , \4245_nGce3 );
or \U$3773 ( \4469 , \4467 , \4468 );
and \U$3774 ( \4470 , \4217 , \4469 );
and \U$3775 ( \4471 , \866 , \4216_nGe5e );
or \U$3776 ( \4472 , \4470 , \4471 );
and \U$3777 ( \4473 , \4188 , \4472 );
and \U$3778 ( \4474 , \830 , \4187_nGe60 );
or \U$3779 ( \4475 , \4473 , \4474 );
and \U$3780 ( \4476 , \4160 , \4475 );
and \U$3781 ( \4477 , \794 , \4159_nG100e );
or \U$3782 ( \4478 , \4476 , \4477 );
and \U$3783 ( \4479 , \4131 , \4478 );
and \U$3784 ( \4480 , \758 , \4130_nG1010 );
or \U$3785 ( \4481 , \4479 , \4480 );
and \U$3786 ( \4482 , \4102 , \4481 );
and \U$3787 ( \4483 , \673 , \4101_nG11f9 );
or \U$3788 ( \4484 , \4482 , \4483 );
nor \U$3789 ( \4485 , \4484 , \1213 );
not \U$3790 ( \4486 , \4485 );
and \U$3791 ( \4487 , \738 , RIb551098_232);
and \U$3792 ( \4488 , \724 , RIb551188_234);
and \U$3793 ( \4489 , RIb551200_235, \726 );
nor \U$3794 ( \4490 , \4488 , \4489 );
and \U$3795 ( \4491 , \710 , RIb551638_244);
and \U$3796 ( \4492 , RIb551278_236, \690 );
nor \U$3797 ( \4493 , \4491 , \4492 );
and \U$3798 ( \4494 , \716 , RIb551548_242);
and \U$3799 ( \4495 , RIb5515c0_243, \713 );
nor \U$3800 ( \4496 , \4494 , \4495 );
and \U$3801 ( \4497 , \695 , RIb551458_240);
and \U$3802 ( \4498 , RIb5514d0_241, \719 );
nor \U$3803 ( \4499 , \4497 , \4498 );
nand \U$3804 ( \4500 , \4490 , \4493 , \4496 , \4499 );
nor \U$3805 ( \4501 , \4487 , \4500 );
and \U$3806 ( \4502 , \740 , RIb551110_233);
and \U$3807 ( \4503 , RIb551020_231, \734 );
nor \U$3808 ( \4504 , \4502 , \4503 );
or \U$3809 ( \4505 , \732 , \4095 );
and \U$3810 ( \4506 , \4505 , RIb550be8_222);
and \U$3811 ( \4507 , RIb5513e0_239, \698 );
nor \U$3812 ( \4508 , \4506 , \4507 );
and \U$3813 ( \4509 , \703 , RIb551368_238);
and \U$3814 ( \4510 , RIb5512f0_237, \705 );
nor \U$3815 ( \4511 , \4509 , \4510 );
nand \U$3816 ( \4512 , \4501 , \4504 , \4508 , \4511 );
buf \U$3817 ( \4513 , \750 );
_DC g1821 ( \4514_nG1821 , \4512 , \4513 );
not \U$3818 ( \4515 , \4514_nG1821 );
nor \U$3819 ( \4516 , \4486 , \4515 );
xor \U$3820 ( \4517 , \673 , \4101_nG11f9 );
xor \U$3821 ( \4518 , \4517 , \4481 );
not \U$3822 ( \4519 , \4518 );
xor \U$3823 ( \4520 , \758 , \4130_nG1010 );
xor \U$3824 ( \4521 , \4520 , \4478 );
not \U$3825 ( \4522 , \4521 );
and \U$3826 ( \4523 , \4519 , \4522 );
and \U$3827 ( \4524 , \4484 , \1213 );
nor \U$3828 ( \4525 , \4524 , \4485 );
nor \U$3829 ( \4526 , \4523 , \4525 );
not \U$3830 ( \4527 , \4526 );
and \U$3831 ( \4528 , RIb5521f0_269, \724 );
and \U$3832 ( \4529 , RIb5526a0_279, \710 );
and \U$3833 ( \4530 , \703 , RIb5523d0_273);
and \U$3834 ( \4531 , RIb552358_272, \705 );
nor \U$3835 ( \4532 , \4530 , \4531 );
and \U$3836 ( \4533 , RIb552010_265, \4505 );
and \U$3837 ( \4534 , \734 , RIb552088_266);
and \U$3838 ( \4535 , RIb552448_274, \698 );
nor \U$3839 ( \4536 , \4533 , \4534 , \4535 );
and \U$3840 ( \4537 , \738 , RIb552100_267);
and \U$3841 ( \4538 , RIb552178_268, \740 );
nor \U$3842 ( \4539 , \4537 , \4538 );
nand \U$3843 ( \4540 , \4532 , \4536 , \4539 );
nor \U$3844 ( \4541 , \4528 , \4529 , \4540 );
and \U$3845 ( \4542 , \716 , RIb5525b0_277);
and \U$3846 ( \4543 , RIb552538_276, \719 );
nor \U$3847 ( \4544 , \4542 , \4543 );
and \U$3848 ( \4545 , \690 , RIb5522e0_271);
and \U$3849 ( \4546 , RIb552628_278, \713 );
nor \U$3850 ( \4547 , \4545 , \4546 );
and \U$3851 ( \4548 , \695 , RIb5524c0_275);
and \U$3852 ( \4549 , RIb552268_270, \726 );
nor \U$3853 ( \4550 , \4548 , \4549 );
nand \U$3854 ( \4551 , \4541 , \4544 , \4547 , \4550 );
_DC g1933 ( \4552_nG1933 , \4551 , \4513 );
or \U$3855 ( \4553 , \4527 , \4552_nG1933 );
not \U$3856 ( \4554 , \4552_nG1933 );
and \U$3857 ( \4555 , \4525 , \4518 );
nor \U$3858 ( \4556 , \4525 , \4518 );
xor \U$3859 ( \4557 , \4518 , \4521 );
nor \U$3860 ( \4558 , \4555 , \4556 , \4557 );
and \U$3861 ( \4559 , \4558 , \4527 );
not \U$3862 ( \4560 , \4559 );
or \U$3863 ( \4561 , \4554 , \4560 );
or \U$3864 ( \4562 , \4558 , \4527 );
nand \U$3865 ( \4563 , \4553 , \4561 , \4562 );
xnor \U$3866 ( \4564 , \4516 , \4563 );
not \U$3867 ( \4565 , \4557 );
nor \U$3868 ( \4566 , \4526 , \4565 );
not \U$3869 ( \4567 , \4566 );
or \U$3870 ( \4568 , \4567 , \4554 );
or \U$3871 ( \4569 , \4515 , \4560 );
or \U$3872 ( \4570 , \4565 , \4554 );
or \U$3873 ( \4571 , \4527 , \4514_nG1821 );
nand \U$3874 ( \4572 , \4571 , \4562 );
nand \U$3875 ( \4573 , \4570 , \4572 );
nand \U$3876 ( \4574 , \4568 , \4569 , \4573 );
xor \U$3877 ( \4575 , \794 , \4159_nG100e );
xor \U$3878 ( \4576 , \4575 , \4475 );
xor \U$3879 ( \4577 , \830 , \4187_nGe60 );
xor \U$3880 ( \4578 , \4577 , \4472 );
nor \U$3881 ( \4579 , \4576 , \4578 );
or \U$3882 ( \4580 , \4521 , \4579 );
and \U$3883 ( \4581 , \4574 , \4580 );
and \U$3884 ( \4582 , RIb552cb8_292, \695 );
and \U$3885 ( \4583 , RIb552a60_287, \726 );
and \U$3886 ( \4584 , \703 , RIb552bc8_290);
and \U$3887 ( \4585 , RIb552b50_289, \705 );
nor \U$3888 ( \4586 , \4584 , \4585 );
and \U$3889 ( \4587 , RIb552808_282, \4505 );
and \U$3890 ( \4588 , \734 , RIb552880_283);
and \U$3891 ( \4589 , RIb552c40_291, \698 );
nor \U$3892 ( \4590 , \4587 , \4588 , \4589 );
and \U$3893 ( \4591 , \738 , RIb5528f8_284);
and \U$3894 ( \4592 , RIb552970_285, \740 );
nor \U$3895 ( \4593 , \4591 , \4592 );
nand \U$3896 ( \4594 , \4586 , \4590 , \4593 );
nor \U$3897 ( \4595 , \4582 , \4583 , \4594 );
and \U$3898 ( \4596 , \690 , RIb552ad8_288);
and \U$3899 ( \4597 , RIb552e20_295, \713 );
nor \U$3900 ( \4598 , \4596 , \4597 );
and \U$3901 ( \4599 , \710 , RIb552e98_296);
and \U$3902 ( \4600 , RIb5529e8_286, \724 );
nor \U$3903 ( \4601 , \4599 , \4600 );
and \U$3904 ( \4602 , \716 , RIb552da8_294);
and \U$3905 ( \4603 , RIb552d30_293, \719 );
nor \U$3906 ( \4604 , \4602 , \4603 );
nand \U$3907 ( \4605 , \4595 , \4598 , \4601 , \4604 );
_DC g172a ( \4606_nG172a , \4605 , \4513 );
nand \U$3908 ( \4607 , \4606_nG172a , \4485 );
not \U$3909 ( \4608 , \4607 );
nor \U$3910 ( \4609 , \4581 , \4608 );
xor \U$3911 ( \4610 , \4564 , \4609 );
not \U$3912 ( \4611 , \4610 );
not \U$3913 ( \4612 , \4576 );
not \U$3914 ( \4613 , \4521 );
or \U$3915 ( \4614 , \4612 , \4613 );
or \U$3916 ( \4615 , \4521 , \4576 );
nand \U$3917 ( \4616 , \4614 , \4615 );
xor \U$3918 ( \4617 , \4578 , \4576 );
nor \U$3919 ( \4618 , \4616 , \4617 );
not \U$3920 ( \4619 , \4618 );
not \U$3921 ( \4620 , \4580 );
nor \U$3922 ( \4621 , \4619 , \4620 );
not \U$3923 ( \4622 , \4621 );
or \U$3924 ( \4623 , \4622 , \4554 );
or \U$3925 ( \4624 , \4619 , \4554 );
nand \U$3926 ( \4625 , \4624 , \4620 );
nand \U$3927 ( \4626 , \4623 , \4625 );
or \U$3928 ( \4627 , \4567 , \4515 );
not \U$3929 ( \4628 , \4606_nG172a );
or \U$3930 ( \4629 , \4628 , \4560 );
or \U$3931 ( \4630 , \4565 , \4515 );
or \U$3932 ( \4631 , \4527 , \4606_nG172a );
nand \U$3933 ( \4632 , \4631 , \4562 );
nand \U$3934 ( \4633 , \4630 , \4632 );
nand \U$3935 ( \4634 , \4627 , \4629 , \4633 );
and \U$3936 ( \4635 , \4626 , \4634 );
not \U$3937 ( \4636 , \4607 );
and \U$3938 ( \4637 , \4574 , \4580 );
not \U$3939 ( \4638 , \4574 );
and \U$3940 ( \4639 , \4638 , \4620 );
nor \U$3941 ( \4640 , \4637 , \4639 );
not \U$3942 ( \4641 , \4640 );
or \U$3943 ( \4642 , \4636 , \4641 );
or \U$3944 ( \4643 , \4640 , \4607 );
nand \U$3945 ( \4644 , \4642 , \4643 );
and \U$3946 ( \4645 , \4635 , \4644 );
xor \U$3947 ( \4646 , \4611 , \4645 );
xor \U$3948 ( \4647 , \4635 , \4644 );
nand \U$3949 ( \4648 , \4514_nG1821 , \4618 );
or \U$3950 ( \4649 , \4580 , \4552_nG1933 );
or \U$3951 ( \4650 , \4580 , \4617 );
nand \U$3952 ( \4651 , \4649 , \4650 );
and \U$3953 ( \4652 , \4648 , \4651 );
and \U$3954 ( \4653 , \4580 , \4617 );
and \U$3955 ( \4654 , \4653 , \4552_nG1933 );
and \U$3956 ( \4655 , \4514_nG1821 , \4621 );
nor \U$3957 ( \4656 , \4652 , \4654 , \4655 );
and \U$3958 ( \4657 , \4606_nG172a , \4566 );
and \U$3959 ( \4658 , \4505 , RIb5537f8_316);
and \U$3960 ( \4659 , \695 , RIb553ca8_326);
and \U$3961 ( \4660 , RIb553d20_327, \719 );
nor \U$3962 ( \4661 , \4659 , \4660 );
and \U$3963 ( \4662 , \724 , RIb5539d8_320);
and \U$3964 ( \4663 , RIb553a50_321, \726 );
nor \U$3965 ( \4664 , \4662 , \4663 );
and \U$3966 ( \4665 , \710 , RIb553e88_330);
and \U$3967 ( \4666 , RIb553ac8_322, \690 );
nor \U$3968 ( \4667 , \4665 , \4666 );
and \U$3969 ( \4668 , \716 , RIb553d98_328);
and \U$3970 ( \4669 , RIb553e10_329, \713 );
nor \U$3971 ( \4670 , \4668 , \4669 );
nand \U$3972 ( \4671 , \4661 , \4664 , \4667 , \4670 );
nor \U$3973 ( \4672 , \4658 , \4671 );
and \U$3974 ( \4673 , \703 , RIb553bb8_324);
and \U$3975 ( \4674 , RIb553c30_325, \698 );
nor \U$3976 ( \4675 , \4673 , \4674 );
and \U$3977 ( \4676 , \740 , RIb553960_319);
and \U$3978 ( \4677 , RIb553870_317, \734 );
nor \U$3979 ( \4678 , \4676 , \4677 );
and \U$3980 ( \4679 , \738 , RIb5538e8_318);
and \U$3981 ( \4680 , RIb553b40_323, \705 );
nor \U$3982 ( \4681 , \4679 , \4680 );
nand \U$3983 ( \4682 , \4672 , \4675 , \4678 , \4681 );
_DC g1613 ( \4683_nG1613 , \4682 , \4513 );
and \U$3984 ( \4684 , \4559 , \4683_nG1613 );
nand \U$3985 ( \4685 , \4606_nG172a , \4557 );
or \U$3986 ( \4686 , \4527 , \4683_nG1613 );
nand \U$3987 ( \4687 , \4686 , \4562 );
and \U$3988 ( \4688 , \4685 , \4687 );
nor \U$3989 ( \4689 , \4657 , \4684 , \4688 );
nand \U$3990 ( \4690 , \4656 , \4689 );
xor \U$3991 ( \4691 , \866 , \4216_nGe5e );
xor \U$3992 ( \4692 , \4691 , \4469 );
xor \U$3993 ( \4693 , \904 , \4245_nGce3 );
xor \U$3994 ( \4694 , \4693 , \4466 );
nor \U$3995 ( \4695 , \4692 , \4694 );
or \U$3996 ( \4696 , \4578 , \4695 );
and \U$3997 ( \4697 , \4690 , \4696 );
nor \U$3998 ( \4698 , \4689 , \4656 );
nor \U$3999 ( \4699 , \4697 , \4698 );
xor \U$4000 ( \4700 , \4626 , \4634 );
not \U$4001 ( \4701 , \4700 );
nand \U$4002 ( \4702 , \4683_nG1613 , \4485 );
not \U$4003 ( \4703 , \4702 );
and \U$4004 ( \4704 , \4701 , \4703 );
and \U$4005 ( \4705 , \4700 , \4702 );
nor \U$4006 ( \4706 , \4704 , \4705 );
nand \U$4007 ( \4707 , \4699 , \4706 );
and \U$4008 ( \4708 , \4647 , \4707 );
and \U$4009 ( \4709 , \4646 , \4708 );
not \U$4010 ( \4710 , \4709 );
and \U$4011 ( \4711 , \4611 , \4645 );
or \U$4012 ( \4712 , \4711 , \4526 );
and \U$4013 ( \4713 , \4563 , \4516 );
and \U$4014 ( \4714 , \4526 , \4711 );
nor \U$4015 ( \4715 , \4713 , \4714 );
nand \U$4016 ( \4716 , \4712 , \4715 );
not \U$4017 ( \4717 , \4716 );
and \U$4018 ( \4718 , \4485 , \4552_nG1933 );
and \U$4019 ( \4719 , \4564 , \4609 );
nor \U$4020 ( \4720 , \4718 , \4719 );
not \U$4021 ( \4721 , \4720 );
and \U$4022 ( \4722 , \4717 , \4721 );
and \U$4023 ( \4723 , \4716 , \4720 );
nor \U$4024 ( \4724 , \4722 , \4723 );
not \U$4025 ( \4725 , \4724 );
or \U$4026 ( \4726 , \4710 , \4725 );
or \U$4027 ( \4727 , \4724 , \4709 );
nand \U$4028 ( \4728 , \4726 , \4727 );
not \U$4029 ( \4729 , \4728 );
not \U$4030 ( \4730 , \4696 );
not \U$4031 ( \4731 , \4698 );
nand \U$4032 ( \4732 , \4731 , \4690 );
not \U$4033 ( \4733 , \4732 );
or \U$4034 ( \4734 , \4730 , \4733 );
or \U$4035 ( \4735 , \4732 , \4696 );
nand \U$4036 ( \4736 , \4734 , \4735 );
not \U$4037 ( \4737 , \4736 );
and \U$4038 ( \4738 , RIb5534b0_309, \695 );
and \U$4039 ( \4739 , RIb553258_304, \726 );
and \U$4040 ( \4740 , \703 , RIb5533c0_307);
and \U$4041 ( \4741 , RIb553348_306, \705 );
nor \U$4042 ( \4742 , \4740 , \4741 );
and \U$4043 ( \4743 , RIb553000_299, \4505 );
and \U$4044 ( \4744 , \734 , RIb553078_300);
and \U$4045 ( \4745 , RIb553438_308, \698 );
nor \U$4046 ( \4746 , \4743 , \4744 , \4745 );
and \U$4047 ( \4747 , \738 , RIb5530f0_301);
and \U$4048 ( \4748 , RIb553168_302, \740 );
nor \U$4049 ( \4749 , \4747 , \4748 );
nand \U$4050 ( \4750 , \4742 , \4746 , \4749 );
nor \U$4051 ( \4751 , \4738 , \4739 , \4750 );
and \U$4052 ( \4752 , \690 , RIb5532d0_305);
and \U$4053 ( \4753 , RIb553618_312, \713 );
nor \U$4054 ( \4754 , \4752 , \4753 );
and \U$4055 ( \4755 , \710 , RIb553690_313);
and \U$4056 ( \4756 , RIb5531e0_303, \724 );
nor \U$4057 ( \4757 , \4755 , \4756 );
and \U$4058 ( \4758 , \716 , RIb5535a0_311);
and \U$4059 ( \4759 , RIb553528_310, \719 );
nor \U$4060 ( \4760 , \4758 , \4759 );
nand \U$4061 ( \4761 , \4751 , \4754 , \4757 , \4760 );
_DC g1506 ( \4762_nG1506 , \4761 , \4513 );
nand \U$4062 ( \4763 , \4762_nG1506 , \4485 );
not \U$4063 ( \4764 , \4763 );
and \U$4064 ( \4765 , \4737 , \4764 );
and \U$4065 ( \4766 , \4736 , \4763 );
nor \U$4066 ( \4767 , \4765 , \4766 );
not \U$4067 ( \4768 , \4767 );
and \U$4068 ( \4769 , \4683_nG1613 , \4566 );
and \U$4069 ( \4770 , \4559 , \4762_nG1506 );
nand \U$4070 ( \4771 , \4683_nG1613 , \4557 );
or \U$4071 ( \4772 , \4527 , \4762_nG1506 );
nand \U$4072 ( \4773 , \4772 , \4562 );
and \U$4073 ( \4774 , \4771 , \4773 );
nor \U$4074 ( \4775 , \4769 , \4770 , \4774 );
and \U$4075 ( \4776 , RIb5541d0_337, \724 );
and \U$4076 ( \4777 , RIb554518_344, \719 );
and \U$4077 ( \4778 , \703 , RIb5543b0_341);
and \U$4078 ( \4779 , RIb554338_340, \705 );
nor \U$4079 ( \4780 , \4778 , \4779 );
and \U$4080 ( \4781 , RIb553ff0_333, \4505 );
and \U$4081 ( \4782 , \734 , RIb554068_334);
and \U$4082 ( \4783 , RIb554428_342, \698 );
nor \U$4083 ( \4784 , \4781 , \4782 , \4783 );
and \U$4084 ( \4785 , \738 , RIb5540e0_335);
and \U$4085 ( \4786 , RIb554158_336, \740 );
nor \U$4086 ( \4787 , \4785 , \4786 );
nand \U$4087 ( \4788 , \4780 , \4784 , \4787 );
nor \U$4088 ( \4789 , \4776 , \4777 , \4788 );
and \U$4089 ( \4790 , \710 , RIb554680_347);
and \U$4090 ( \4791 , RIb554590_345, \716 );
nor \U$4091 ( \4792 , \4790 , \4791 );
and \U$4092 ( \4793 , \695 , RIb5544a0_343);
and \U$4093 ( \4794 , RIb554608_346, \713 );
nor \U$4094 ( \4795 , \4793 , \4794 );
and \U$4095 ( \4796 , \690 , RIb5542c0_339);
and \U$4096 ( \4797 , RIb554248_338, \726 );
nor \U$4097 ( \4798 , \4796 , \4797 );
nand \U$4098 ( \4799 , \4789 , \4792 , \4795 , \4798 );
_DC g140b ( \4800_nG140b , \4799 , \4513 );
nand \U$4099 ( \4801 , \4800_nG140b , \4485 );
or \U$4100 ( \4802 , \4775 , \4801 );
and \U$4101 ( \4803 , \4578 , \4692 );
nor \U$4102 ( \4804 , \4578 , \4692 );
xor \U$4103 ( \4805 , \4692 , \4694 );
nor \U$4104 ( \4806 , \4803 , \4804 , \4805 );
and \U$4105 ( \4807 , \4806 , \4696 );
and \U$4106 ( \4808 , \4552_nG1933 , \4807 );
not \U$4107 ( \4809 , \4696 );
and \U$4108 ( \4810 , \4554 , \4809 );
or \U$4109 ( \4811 , \4806 , \4696 );
not \U$4110 ( \4812 , \4811 );
nor \U$4111 ( \4813 , \4808 , \4810 , \4812 );
nand \U$4112 ( \4814 , \4606_nG172a , \4618 );
or \U$4113 ( \4815 , \4580 , \4514_nG1821 );
nand \U$4114 ( \4816 , \4815 , \4650 );
and \U$4115 ( \4817 , \4814 , \4816 );
and \U$4116 ( \4818 , \4653 , \4514_nG1821 );
and \U$4117 ( \4819 , \4606_nG172a , \4621 );
nor \U$4118 ( \4820 , \4817 , \4818 , \4819 );
or \U$4119 ( \4821 , \4813 , \4820 );
nand \U$4120 ( \4822 , \4802 , \4821 );
nand \U$4121 ( \4823 , \4768 , \4822 );
not \U$4122 ( \4824 , \4823 );
or \U$4123 ( \4825 , \4706 , \4699 );
nand \U$4124 ( \4826 , \4825 , \4707 );
nand \U$4125 ( \4827 , \4824 , \4826 );
xor \U$4126 ( \4828 , \4647 , \4707 );
not \U$4127 ( \4829 , \4700 );
nor \U$4128 ( \4830 , \4829 , \4702 );
nor \U$4129 ( \4831 , \4828 , \4830 );
or \U$4130 ( \4832 , \4827 , \4831 );
nand \U$4131 ( \4833 , \4830 , \4828 );
nand \U$4132 ( \4834 , \4832 , \4833 );
xor \U$4133 ( \4835 , \4646 , \4708 );
xor \U$4134 ( \4836 , \4834 , \4835 );
not \U$4135 ( \4837 , \4826 );
not \U$4136 ( \4838 , \4823 );
and \U$4137 ( \4839 , \4837 , \4838 );
and \U$4138 ( \4840 , \4826 , \4823 );
nor \U$4139 ( \4841 , \4839 , \4840 );
not \U$4140 ( \4842 , \4763 );
nand \U$4141 ( \4843 , \4842 , \4736 );
xor \U$4142 ( \4844 , \4841 , \4843 );
nand \U$4143 ( \4845 , \4762_nG1506 , \4618 );
or \U$4144 ( \4846 , \4580 , \4683_nG1613 );
nand \U$4145 ( \4847 , \4846 , \4650 );
and \U$4146 ( \4848 , \4845 , \4847 );
and \U$4147 ( \4849 , \4653 , \4683_nG1613 );
and \U$4148 ( \4850 , \4762_nG1506 , \4621 );
nor \U$4149 ( \4851 , \4848 , \4849 , \4850 );
and \U$4150 ( \4852 , RIb554c98_360, \695 );
and \U$4151 ( \4853 , RIb554a40_355, \726 );
and \U$4152 ( \4854 , \703 , RIb554ba8_358);
and \U$4153 ( \4855 , RIb554b30_357, \705 );
nor \U$4154 ( \4856 , \4854 , \4855 );
and \U$4155 ( \4857 , RIb5547e8_350, \4505 );
and \U$4156 ( \4858 , \734 , RIb554860_351);
and \U$4157 ( \4859 , RIb554c20_359, \698 );
nor \U$4158 ( \4860 , \4857 , \4858 , \4859 );
and \U$4159 ( \4861 , \738 , RIb5548d8_352);
and \U$4160 ( \4862 , RIb554950_353, \740 );
nor \U$4161 ( \4863 , \4861 , \4862 );
nand \U$4162 ( \4864 , \4856 , \4860 , \4863 );
nor \U$4163 ( \4865 , \4852 , \4853 , \4864 );
and \U$4164 ( \4866 , \690 , RIb554ab8_356);
and \U$4165 ( \4867 , RIb554e00_363, \713 );
nor \U$4166 ( \4868 , \4866 , \4867 );
and \U$4167 ( \4869 , \710 , RIb554e78_364);
and \U$4168 ( \4870 , RIb5549c8_354, \724 );
nor \U$4169 ( \4871 , \4869 , \4870 );
and \U$4170 ( \4872 , \716 , RIb554d88_362);
and \U$4171 ( \4873 , RIb554d10_361, \719 );
nor \U$4172 ( \4874 , \4872 , \4873 );
nand \U$4173 ( \4875 , \4865 , \4868 , \4871 , \4874 );
_DC g1212 ( \4876_nG1212 , \4875 , \4513 );
nand \U$4174 ( \4877 , \4876_nG1212 , \4485 );
xor \U$4175 ( \4878 , \4851 , \4877 );
and \U$4176 ( \4879 , RIb555490_377, \695 );
and \U$4177 ( \4880 , RIb555238_372, \726 );
and \U$4178 ( \4881 , \703 , RIb5553a0_375);
and \U$4179 ( \4882 , RIb555328_374, \705 );
nor \U$4180 ( \4883 , \4881 , \4882 );
and \U$4181 ( \4884 , RIb554fe0_367, \4505 );
and \U$4182 ( \4885 , \734 , RIb555058_368);
and \U$4183 ( \4886 , RIb555418_376, \698 );
nor \U$4184 ( \4887 , \4884 , \4885 , \4886 );
and \U$4185 ( \4888 , \738 , RIb5550d0_369);
and \U$4186 ( \4889 , RIb555148_370, \740 );
nor \U$4187 ( \4890 , \4888 , \4889 );
nand \U$4188 ( \4891 , \4883 , \4887 , \4890 );
nor \U$4189 ( \4892 , \4879 , \4880 , \4891 );
and \U$4190 ( \4893 , \690 , RIb5552b0_373);
and \U$4191 ( \4894 , RIb5555f8_380, \713 );
nor \U$4192 ( \4895 , \4893 , \4894 );
and \U$4193 ( \4896 , \710 , RIb555670_381);
and \U$4194 ( \4897 , RIb5551c0_371, \724 );
nor \U$4195 ( \4898 , \4896 , \4897 );
and \U$4196 ( \4899 , \716 , RIb555580_379);
and \U$4197 ( \4900 , RIb555508_378, \719 );
nor \U$4198 ( \4901 , \4899 , \4900 );
nand \U$4199 ( \4902 , \4892 , \4895 , \4898 , \4901 );
_DC g1319 ( \4903_nG1319 , \4902 , \4513 );
and \U$4200 ( \4904 , \4903_nG1319 , \4559 );
or \U$4201 ( \4905 , \4527 , \4903_nG1319 );
nand \U$4202 ( \4906 , \4905 , \4562 );
nand \U$4203 ( \4907 , \4800_nG140b , \4557 );
and \U$4204 ( \4908 , \4906 , \4907 );
and \U$4205 ( \4909 , \4800_nG140b , \4566 );
nor \U$4206 ( \4910 , \4904 , \4908 , \4909 );
and \U$4207 ( \4911 , \4878 , \4910 );
and \U$4208 ( \4912 , \4851 , \4877 );
or \U$4209 ( \4913 , \4911 , \4912 );
not \U$4210 ( \4914 , \4913 );
xor \U$4211 ( \4915 , \940 , \4273_nGce1 );
xor \U$4212 ( \4916 , \4915 , \4463 );
not \U$4213 ( \4917 , \4916 );
not \U$4214 ( \4918 , \4694 );
or \U$4215 ( \4919 , \4917 , \4918 );
or \U$4216 ( \4920 , \4694 , \4916 );
nand \U$4217 ( \4921 , \4919 , \4920 );
xor \U$4218 ( \4922 , \978 , \4302_nGbb6 );
xor \U$4219 ( \4923 , \4922 , \4460 );
xor \U$4220 ( \4924 , \4923 , \4916 );
nor \U$4221 ( \4925 , \4921 , \4924 );
not \U$4222 ( \4926 , \4925 );
nor \U$4223 ( \4927 , \4916 , \4923 );
or \U$4224 ( \4928 , \4927 , \4694 );
not \U$4225 ( \4929 , \4928 );
nor \U$4226 ( \4930 , \4926 , \4929 );
not \U$4227 ( \4931 , \4930 );
or \U$4228 ( \4932 , \4931 , \4554 );
or \U$4229 ( \4933 , \4926 , \4554 );
nand \U$4230 ( \4934 , \4933 , \4929 );
nand \U$4231 ( \4935 , \4932 , \4934 );
not \U$4232 ( \4936 , \4805 );
nor \U$4233 ( \4937 , \4809 , \4936 );
not \U$4234 ( \4938 , \4937 );
or \U$4235 ( \4939 , \4938 , \4515 );
not \U$4236 ( \4940 , \4807 );
or \U$4237 ( \4941 , \4628 , \4940 );
or \U$4238 ( \4942 , \4936 , \4515 );
or \U$4239 ( \4943 , \4696 , \4606_nG172a );
nand \U$4240 ( \4944 , \4943 , \4811 );
nand \U$4241 ( \4945 , \4942 , \4944 );
nand \U$4242 ( \4946 , \4939 , \4941 , \4945 );
and \U$4243 ( \4947 , \4935 , \4946 );
nand \U$4244 ( \4948 , \4914 , \4947 );
not \U$4245 ( \4949 , \4948 );
nand \U$4246 ( \4950 , \4552_nG1933 , \4805 );
or \U$4247 ( \4951 , \4696 , \4514_nG1821 );
nand \U$4248 ( \4952 , \4951 , \4811 );
and \U$4249 ( \4953 , \4950 , \4952 );
and \U$4250 ( \4954 , \4807 , \4514_nG1821 );
and \U$4251 ( \4955 , \4552_nG1933 , \4937 );
nor \U$4252 ( \4956 , \4953 , \4954 , \4955 );
not \U$4253 ( \4957 , \4956 );
nand \U$4254 ( \4958 , \4683_nG1613 , \4618 );
or \U$4255 ( \4959 , \4580 , \4606_nG172a );
nand \U$4256 ( \4960 , \4959 , \4650 );
and \U$4257 ( \4961 , \4958 , \4960 );
and \U$4258 ( \4962 , \4653 , \4606_nG172a );
and \U$4259 ( \4963 , \4683_nG1613 , \4621 );
nor \U$4260 ( \4964 , \4961 , \4962 , \4963 );
or \U$4261 ( \4965 , \4964 , \4928 );
nand \U$4262 ( \4966 , \4928 , \4964 );
nand \U$4263 ( \4967 , \4965 , \4966 );
not \U$4264 ( \4968 , \4967 );
or \U$4265 ( \4969 , \4957 , \4968 );
or \U$4266 ( \4970 , \4967 , \4956 );
nand \U$4267 ( \4971 , \4969 , \4970 );
nand \U$4268 ( \4972 , \4903_nG1319 , \4485 );
and \U$4269 ( \4973 , \4762_nG1506 , \4566 );
and \U$4270 ( \4974 , \4559 , \4800_nG140b );
nand \U$4271 ( \4975 , \4762_nG1506 , \4557 );
or \U$4272 ( \4976 , \4527 , \4800_nG140b );
nand \U$4273 ( \4977 , \4976 , \4562 );
and \U$4274 ( \4978 , \4975 , \4977 );
nor \U$4275 ( \4979 , \4973 , \4974 , \4978 );
xor \U$4276 ( \4980 , \4972 , \4979 );
and \U$4277 ( \4981 , \4971 , \4980 );
nand \U$4278 ( \4982 , \4949 , \4981 );
xor \U$4279 ( \4983 , \4813 , \4820 );
not \U$4280 ( \4984 , \4983 );
xnor \U$4281 ( \4985 , \4801 , \4775 );
not \U$4282 ( \4986 , \4985 );
or \U$4283 ( \4987 , \4984 , \4986 );
or \U$4284 ( \4988 , \4985 , \4983 );
nand \U$4285 ( \4989 , \4987 , \4988 );
or \U$4286 ( \4990 , \4979 , \4972 );
not \U$4287 ( \4991 , \4956 );
not \U$4288 ( \4992 , \4929 );
and \U$4289 ( \4993 , \4991 , \4992 );
and \U$4290 ( \4994 , \4956 , \4929 );
nor \U$4291 ( \4995 , \4994 , \4964 );
nor \U$4292 ( \4996 , \4993 , \4995 );
nand \U$4293 ( \4997 , \4990 , \4996 );
nor \U$4294 ( \4998 , \4989 , \4997 );
xor \U$4295 ( \4999 , \4982 , \4998 );
not \U$4296 ( \5000 , \4767 );
not \U$4297 ( \5001 , \4822 );
and \U$4298 ( \5002 , \5000 , \5001 );
and \U$4299 ( \5003 , \4767 , \4822 );
nor \U$4300 ( \5004 , \5002 , \5003 );
and \U$4301 ( \5005 , \4999 , \5004 );
and \U$4302 ( \5006 , \4982 , \4998 );
or \U$4303 ( \5007 , \5005 , \5006 );
and \U$4304 ( \5008 , \4844 , \5007 );
and \U$4305 ( \5009 , \4841 , \4843 );
or \U$4306 ( \5010 , \5008 , \5009 );
not \U$4307 ( \5011 , \4827 );
not \U$4308 ( \5012 , \4831 );
nand \U$4309 ( \5013 , \5012 , \4833 );
not \U$4310 ( \5014 , \5013 );
or \U$4311 ( \5015 , \5011 , \5014 );
or \U$4312 ( \5016 , \5013 , \4827 );
nand \U$4313 ( \5017 , \5015 , \5016 );
xor \U$4314 ( \5018 , \5010 , \5017 );
xor \U$4315 ( \5019 , \4851 , \4877 );
xor \U$4316 ( \5020 , \5019 , \4910 );
not \U$4317 ( \5021 , \5020 );
xor \U$4318 ( \5022 , \4935 , \4946 );
nand \U$4319 ( \5023 , \5021 , \5022 );
not \U$4320 ( \5024 , \5023 );
and \U$4321 ( \5025 , \4903_nG1319 , \4566 );
and \U$4322 ( \5026 , \4559 , \4876_nG1212 );
nand \U$4323 ( \5027 , \4903_nG1319 , \4557 );
or \U$4324 ( \5028 , \4527 , \4876_nG1212 );
nand \U$4325 ( \5029 , \5028 , \4562 );
and \U$4326 ( \5030 , \5027 , \5029 );
nor \U$4327 ( \5031 , \5025 , \5026 , \5030 );
nand \U$4328 ( \5032 , \4800_nG140b , \4618 );
or \U$4329 ( \5033 , \4580 , \4762_nG1506 );
nand \U$4330 ( \5034 , \5033 , \4650 );
and \U$4331 ( \5035 , \5032 , \5034 );
and \U$4332 ( \5036 , \4653 , \4762_nG1506 );
and \U$4333 ( \5037 , \4800_nG140b , \4621 );
nor \U$4334 ( \5038 , \5035 , \5036 , \5037 );
and \U$4335 ( \5039 , \5031 , \5038 );
not \U$4336 ( \5040 , \5039 );
and \U$4337 ( \5041 , RIb5561b0_405, \724 );
and \U$4338 ( \5042 , RIb5564f8_412, \719 );
and \U$4339 ( \5043 , \703 , RIb556390_409);
and \U$4340 ( \5044 , RIb556318_408, \705 );
nor \U$4341 ( \5045 , \5043 , \5044 );
and \U$4342 ( \5046 , RIb555fd0_401, \4505 );
and \U$4343 ( \5047 , \734 , RIb556048_402);
and \U$4344 ( \5048 , RIb556408_410, \698 );
nor \U$4345 ( \5049 , \5046 , \5047 , \5048 );
and \U$4346 ( \5050 , \738 , RIb5560c0_403);
and \U$4347 ( \5051 , RIb556138_404, \740 );
nor \U$4348 ( \5052 , \5050 , \5051 );
nand \U$4349 ( \5053 , \5045 , \5049 , \5052 );
nor \U$4350 ( \5054 , \5041 , \5042 , \5053 );
and \U$4351 ( \5055 , \710 , RIb556660_415);
and \U$4352 ( \5056 , RIb556570_413, \716 );
nor \U$4353 ( \5057 , \5055 , \5056 );
and \U$4354 ( \5058 , \695 , RIb556480_411);
and \U$4355 ( \5059 , RIb5565e8_414, \713 );
nor \U$4356 ( \5060 , \5058 , \5059 );
and \U$4357 ( \5061 , \690 , RIb5562a0_407);
and \U$4358 ( \5062 , RIb556228_406, \726 );
nor \U$4359 ( \5063 , \5061 , \5062 );
nand \U$4360 ( \5064 , \5054 , \5057 , \5060 , \5063 );
_DC g112f ( \5065_nG112f , \5064 , \4513 );
nand \U$4361 ( \5066 , \5065_nG112f , \4485 );
not \U$4362 ( \5067 , \5066 );
and \U$4363 ( \5068 , \5040 , \5067 );
nor \U$4364 ( \5069 , \5031 , \5038 );
nor \U$4365 ( \5070 , \5068 , \5069 );
and \U$4366 ( \5071 , \4928 , \4924 );
and \U$4367 ( \5072 , \4552_nG1933 , \5071 );
or \U$4368 ( \5073 , \4928 , \4552_nG1933 );
or \U$4369 ( \5074 , \4928 , \4924 );
nand \U$4370 ( \5075 , \5073 , \5074 );
nand \U$4371 ( \5076 , \4514_nG1821 , \4925 );
and \U$4372 ( \5077 , \5075 , \5076 );
and \U$4373 ( \5078 , \4514_nG1821 , \4930 );
nor \U$4374 ( \5079 , \5072 , \5077 , \5078 );
nand \U$4375 ( \5080 , \4606_nG172a , \4805 );
or \U$4376 ( \5081 , \4696 , \4683_nG1613 );
nand \U$4377 ( \5082 , \5081 , \4811 );
and \U$4378 ( \5083 , \5080 , \5082 );
and \U$4379 ( \5084 , \4807 , \4683_nG1613 );
and \U$4380 ( \5085 , \4606_nG172a , \4937 );
nor \U$4381 ( \5086 , \5083 , \5084 , \5085 );
nand \U$4382 ( \5087 , \5079 , \5086 );
xor \U$4383 ( \5088 , \1014 , \4331_nGbb4 );
xor \U$4384 ( \5089 , \5088 , \4457 );
xor \U$4385 ( \5090 , \1046 , \4360_nGade );
xor \U$4386 ( \5091 , \5090 , \4454 );
nor \U$4387 ( \5092 , \5089 , \5091 );
or \U$4388 ( \5093 , \4923 , \5092 );
and \U$4389 ( \5094 , \5087 , \5093 );
nor \U$4390 ( \5095 , \5086 , \5079 );
nor \U$4391 ( \5096 , \5094 , \5095 );
nor \U$4392 ( \5097 , \5070 , \5096 );
nand \U$4393 ( \5098 , \5024 , \5097 );
not \U$4394 ( \5099 , \4913 );
not \U$4395 ( \5100 , \4947 );
and \U$4396 ( \5101 , \5099 , \5100 );
and \U$4397 ( \5102 , \4913 , \4947 );
nor \U$4398 ( \5103 , \5101 , \5102 );
not \U$4399 ( \5104 , \5103 );
xor \U$4400 ( \5105 , \4971 , \4980 );
nand \U$4401 ( \5106 , \5104 , \5105 );
xor \U$4402 ( \5107 , \5098 , \5106 );
and \U$4403 ( \5108 , \4989 , \4997 );
nor \U$4404 ( \5109 , \5108 , \4998 );
and \U$4405 ( \5110 , \5107 , \5109 );
and \U$4406 ( \5111 , \5098 , \5106 );
or \U$4407 ( \5112 , \5110 , \5111 );
not \U$4408 ( \5113 , \4985 );
nand \U$4409 ( \5114 , \5113 , \4983 );
xor \U$4410 ( \5115 , \5112 , \5114 );
xor \U$4411 ( \5116 , \4982 , \4998 );
xor \U$4412 ( \5117 , \5116 , \5004 );
and \U$4413 ( \5118 , \5115 , \5117 );
and \U$4414 ( \5119 , \5112 , \5114 );
or \U$4415 ( \5120 , \5118 , \5119 );
xor \U$4416 ( \5121 , \4841 , \4843 );
xor \U$4417 ( \5122 , \5121 , \5007 );
and \U$4418 ( \5123 , \5120 , \5122 );
not \U$4419 ( \5124 , \4948 );
not \U$4420 ( \5125 , \4981 );
or \U$4421 ( \5126 , \5124 , \5125 );
or \U$4422 ( \5127 , \4981 , \4948 );
nand \U$4423 ( \5128 , \5126 , \5127 );
not \U$4424 ( \5129 , \5105 );
not \U$4425 ( \5130 , \5103 );
or \U$4426 ( \5131 , \5129 , \5130 );
or \U$4427 ( \5132 , \5103 , \5105 );
nand \U$4428 ( \5133 , \5131 , \5132 );
not \U$4429 ( \5134 , \5089 );
not \U$4430 ( \5135 , \4923 );
or \U$4431 ( \5136 , \5134 , \5135 );
or \U$4432 ( \5137 , \4923 , \5089 );
nand \U$4433 ( \5138 , \5136 , \5137 );
xor \U$4434 ( \5139 , \5091 , \5089 );
nor \U$4435 ( \5140 , \5138 , \5139 );
not \U$4436 ( \5141 , \5140 );
not \U$4437 ( \5142 , \5093 );
nor \U$4438 ( \5143 , \5141 , \5142 );
not \U$4439 ( \5144 , \5143 );
or \U$4440 ( \5145 , \5144 , \4554 );
or \U$4441 ( \5146 , \5141 , \4554 );
nand \U$4442 ( \5147 , \5146 , \5142 );
nand \U$4443 ( \5148 , \5145 , \5147 );
not \U$4444 ( \5149 , \5071 );
or \U$4445 ( \5150 , \5149 , \4515 );
or \U$4446 ( \5151 , \4628 , \4931 );
or \U$4447 ( \5152 , \4926 , \4628 );
or \U$4448 ( \5153 , \4928 , \4514_nG1821 );
nand \U$4449 ( \5154 , \5153 , \5074 );
nand \U$4450 ( \5155 , \5152 , \5154 );
nand \U$4451 ( \5156 , \5150 , \5151 , \5155 );
and \U$4452 ( \5157 , \5148 , \5156 );
not \U$4453 ( \5158 , \5157 );
nand \U$4454 ( \5159 , \4903_nG1319 , \4618 );
or \U$4455 ( \5160 , \4580 , \4800_nG140b );
nand \U$4456 ( \5161 , \5160 , \4650 );
and \U$4457 ( \5162 , \5159 , \5161 );
and \U$4458 ( \5163 , \4653 , \4800_nG140b );
and \U$4459 ( \5164 , \4903_nG1319 , \4621 );
nor \U$4460 ( \5165 , \5162 , \5163 , \5164 );
nand \U$4461 ( \5166 , \4683_nG1613 , \4805 );
or \U$4462 ( \5167 , \4696 , \4762_nG1506 );
nand \U$4463 ( \5168 , \5167 , \4811 );
and \U$4464 ( \5169 , \5166 , \5168 );
and \U$4465 ( \5170 , \4807 , \4762_nG1506 );
and \U$4466 ( \5171 , \4683_nG1613 , \4937 );
nor \U$4467 ( \5172 , \5169 , \5170 , \5171 );
xor \U$4468 ( \5173 , \5165 , \5172 );
and \U$4469 ( \5174 , \5065_nG112f , \4559 );
or \U$4470 ( \5175 , \4527 , \5065_nG112f );
nand \U$4471 ( \5176 , \5175 , \4562 );
nand \U$4472 ( \5177 , \4876_nG1212 , \4557 );
and \U$4473 ( \5178 , \5176 , \5177 );
and \U$4474 ( \5179 , \4876_nG1212 , \4566 );
nor \U$4475 ( \5180 , \5174 , \5178 , \5179 );
and \U$4476 ( \5181 , \5173 , \5180 );
and \U$4477 ( \5182 , \5165 , \5172 );
or \U$4478 ( \5183 , \5181 , \5182 );
nor \U$4479 ( \5184 , \5158 , \5183 );
not \U$4480 ( \5185 , \5093 );
not \U$4481 ( \5186 , \5095 );
nand \U$4482 ( \5187 , \5186 , \5087 );
not \U$4483 ( \5188 , \5187 );
or \U$4484 ( \5189 , \5185 , \5188 );
or \U$4485 ( \5190 , \5187 , \5093 );
nand \U$4486 ( \5191 , \5189 , \5190 );
not \U$4487 ( \5192 , \5066 );
nor \U$4488 ( \5193 , \5039 , \5069 );
not \U$4489 ( \5194 , \5193 );
or \U$4490 ( \5195 , \5192 , \5194 );
or \U$4491 ( \5196 , \5193 , \5066 );
nand \U$4492 ( \5197 , \5195 , \5196 );
and \U$4493 ( \5198 , \5191 , \5197 );
and \U$4494 ( \5199 , \5184 , \5198 );
xor \U$4495 ( \5200 , \5133 , \5199 );
xnor \U$4496 ( \5201 , \5096 , \5070 );
not \U$4497 ( \5202 , \5020 );
not \U$4498 ( \5203 , \5022 );
and \U$4499 ( \5204 , \5202 , \5203 );
and \U$4500 ( \5205 , \5020 , \5022 );
nor \U$4501 ( \5206 , \5204 , \5205 );
nand \U$4502 ( \5207 , \5201 , \5206 );
and \U$4503 ( \5208 , \5200 , \5207 );
and \U$4504 ( \5209 , \5133 , \5199 );
or \U$4505 ( \5210 , \5208 , \5209 );
nand \U$4506 ( \5211 , \5128 , \5210 );
or \U$4507 ( \5212 , \5210 , \5128 );
nand \U$4508 ( \5213 , \5211 , \5212 );
not \U$4509 ( \5214 , \5213 );
xor \U$4510 ( \5215 , \5098 , \5106 );
xor \U$4511 ( \5216 , \5215 , \5109 );
not \U$4512 ( \5217 , \5216 );
and \U$4513 ( \5218 , \5214 , \5217 );
and \U$4514 ( \5219 , \5213 , \5216 );
nor \U$4515 ( \5220 , \5218 , \5219 );
not \U$4516 ( \5221 , \5097 );
not \U$4517 ( \5222 , \5023 );
or \U$4518 ( \5223 , \5221 , \5222 );
or \U$4519 ( \5224 , \5023 , \5097 );
nand \U$4520 ( \5225 , \5223 , \5224 );
xor \U$4521 ( \5226 , \5133 , \5199 );
xor \U$4522 ( \5227 , \5226 , \5207 );
and \U$4523 ( \5228 , \5225 , \5227 );
xor \U$4524 ( \5229 , \5191 , \5197 );
not \U$4525 ( \5230 , \5229 );
not \U$4526 ( \5231 , \5183 );
not \U$4527 ( \5232 , \5157 );
and \U$4528 ( \5233 , \5231 , \5232 );
and \U$4529 ( \5234 , \5183 , \5157 );
nor \U$4530 ( \5235 , \5233 , \5234 );
nor \U$4531 ( \5236 , \5230 , \5235 );
xor \U$4532 ( \5237 , \5148 , \5156 );
xor \U$4533 ( \5238 , \5165 , \5172 );
xor \U$4534 ( \5239 , \5238 , \5180 );
not \U$4535 ( \5240 , \5239 );
and \U$4536 ( \5241 , \5237 , \5240 );
or \U$4537 ( \5242 , \5144 , \4515 );
and \U$4538 ( \5243 , \5093 , \5139 );
not \U$4539 ( \5244 , \5243 );
or \U$4540 ( \5245 , \4554 , \5244 );
or \U$4541 ( \5246 , \5141 , \4515 );
or \U$4542 ( \5247 , \5093 , \4552_nG1933 );
or \U$4543 ( \5248 , \5093 , \5139 );
nand \U$4544 ( \5249 , \5247 , \5248 );
nand \U$4545 ( \5250 , \5246 , \5249 );
nand \U$4546 ( \5251 , \5242 , \5245 , \5250 );
xor \U$4547 ( \5252 , RIb54a900_11, \4418_nG97f );
xor \U$4548 ( \5253 , \5252 , \4448 );
not \U$4549 ( \5254 , \5253 );
xor \U$4550 ( \5255 , \1078 , \4389_nGae0 );
xor \U$4551 ( \5256 , \5255 , \4451 );
not \U$4552 ( \5257 , \5256 );
and \U$4553 ( \5258 , \5254 , \5257 );
or \U$4554 ( \5259 , \5091 , \5258 );
xor \U$4555 ( \5260 , \5251 , \5259 );
or \U$4556 ( \5261 , \5149 , \4628 );
not \U$4557 ( \5262 , \4683_nG1613 );
or \U$4558 ( \5263 , \5262 , \4931 );
or \U$4559 ( \5264 , \4926 , \5262 );
or \U$4560 ( \5265 , \4928 , \4606_nG172a );
nand \U$4561 ( \5266 , \5265 , \5074 );
nand \U$4562 ( \5267 , \5264 , \5266 );
nand \U$4563 ( \5268 , \5261 , \5263 , \5267 );
and \U$4564 ( \5269 , \5260 , \5268 );
and \U$4565 ( \5270 , \5251 , \5259 );
or \U$4566 ( \5271 , \5269 , \5270 );
nand \U$4567 ( \5272 , \4876_nG1212 , \4618 );
or \U$4568 ( \5273 , \4580 , \4903_nG1319 );
nand \U$4569 ( \5274 , \5273 , \4650 );
and \U$4570 ( \5275 , \5272 , \5274 );
and \U$4571 ( \5276 , \4653 , \4903_nG1319 );
and \U$4572 ( \5277 , \4876_nG1212 , \4621 );
nor \U$4573 ( \5278 , \5275 , \5276 , \5277 );
nand \U$4574 ( \5279 , \4762_nG1506 , \4805 );
or \U$4575 ( \5280 , \4696 , \4800_nG140b );
nand \U$4576 ( \5281 , \5280 , \4811 );
and \U$4577 ( \5282 , \5279 , \5281 );
and \U$4578 ( \5283 , \4807 , \4800_nG140b );
and \U$4579 ( \5284 , \4762_nG1506 , \4937 );
nor \U$4580 ( \5285 , \5282 , \5283 , \5284 );
xor \U$4581 ( \5286 , \5278 , \5285 );
and \U$4582 ( \5287 , RIb555df0_397, \713 );
and \U$4583 ( \5288 , RIb5559b8_388, \724 );
and \U$4584 ( \5289 , \703 , RIb555b98_392);
and \U$4585 ( \5290 , RIb555b20_391, \705 );
nor \U$4586 ( \5291 , \5289 , \5290 );
and \U$4587 ( \5292 , RIb5557d8_384, \4505 );
and \U$4588 ( \5293 , \734 , RIb555850_385);
and \U$4589 ( \5294 , RIb555c10_393, \698 );
nor \U$4590 ( \5295 , \5292 , \5293 , \5294 );
and \U$4591 ( \5296 , \738 , RIb5558c8_386);
and \U$4592 ( \5297 , RIb555940_387, \740 );
nor \U$4593 ( \5298 , \5296 , \5297 );
nand \U$4594 ( \5299 , \5291 , \5295 , \5298 );
nor \U$4595 ( \5300 , \5287 , \5288 , \5299 );
and \U$4596 ( \5301 , \690 , RIb555aa8_390);
and \U$4597 ( \5302 , RIb555d00_395, \719 );
nor \U$4598 ( \5303 , \5301 , \5302 );
and \U$4599 ( \5304 , \710 , RIb555e68_398);
and \U$4600 ( \5305 , RIb555d78_396, \716 );
nor \U$4601 ( \5306 , \5304 , \5305 );
and \U$4602 ( \5307 , \695 , RIb555c88_394);
and \U$4603 ( \5308 , RIb555a30_389, \726 );
nor \U$4604 ( \5309 , \5307 , \5308 );
nand \U$4605 ( \5310 , \5300 , \5303 , \5306 , \5309 );
_DC g1029 ( \5311_nG1029 , \5310 , \4513 );
and \U$4606 ( \5312 , \5311_nG1029 , \4559 );
or \U$4607 ( \5313 , \4527 , \5311_nG1029 );
nand \U$4608 ( \5314 , \5313 , \4562 );
nand \U$4609 ( \5315 , \5065_nG112f , \4557 );
and \U$4610 ( \5316 , \5314 , \5315 );
and \U$4611 ( \5317 , \5065_nG112f , \4566 );
nor \U$4612 ( \5318 , \5312 , \5316 , \5317 );
and \U$4613 ( \5319 , \5286 , \5318 );
and \U$4614 ( \5320 , \5278 , \5285 );
or \U$4615 ( \5321 , \5319 , \5320 );
not \U$4616 ( \5322 , \5321 );
and \U$4617 ( \5323 , \5271 , \5322 );
and \U$4618 ( \5324 , \5241 , \5323 );
xor \U$4619 ( \5325 , \5236 , \5324 );
or \U$4620 ( \5326 , \5206 , \5201 );
nand \U$4621 ( \5327 , \5326 , \5207 );
and \U$4622 ( \5328 , \5325 , \5327 );
and \U$4623 ( \5329 , \5236 , \5324 );
or \U$4624 ( \5330 , \5328 , \5329 );
xor \U$4625 ( \5331 , \5133 , \5199 );
xor \U$4626 ( \5332 , \5331 , \5207 );
and \U$4627 ( \5333 , \5330 , \5332 );
and \U$4628 ( \5334 , \5225 , \5330 );
or \U$4629 ( \5335 , \5228 , \5333 , \5334 );
xor \U$4630 ( \5336 , \5220 , \5335 );
xor \U$4631 ( \5337 , \5236 , \5324 );
xor \U$4632 ( \5338 , \5337 , \5327 );
xor \U$4633 ( \5339 , \5184 , \5198 );
nor \U$4634 ( \5340 , \5338 , \5339 );
not \U$4635 ( \5341 , \5229 );
not \U$4636 ( \5342 , \5235 );
and \U$4637 ( \5343 , \5341 , \5342 );
and \U$4638 ( \5344 , \5229 , \5235 );
nor \U$4639 ( \5345 , \5343 , \5344 );
and \U$4640 ( \5346 , \738 , RIb5570b0_437);
and \U$4641 ( \5347 , \695 , RIb557470_445);
and \U$4642 ( \5348 , RIb5574e8_446, \719 );
nor \U$4643 ( \5349 , \5347 , \5348 );
and \U$4644 ( \5350 , \724 , RIb5571a0_439);
and \U$4645 ( \5351 , RIb557218_440, \726 );
nor \U$4646 ( \5352 , \5350 , \5351 );
and \U$4647 ( \5353 , \710 , RIb557650_449);
and \U$4648 ( \5354 , RIb557290_441, \690 );
nor \U$4649 ( \5355 , \5353 , \5354 );
and \U$4650 ( \5356 , \716 , RIb557560_447);
and \U$4651 ( \5357 , RIb5575d8_448, \713 );
nor \U$4652 ( \5358 , \5356 , \5357 );
nand \U$4653 ( \5359 , \5349 , \5352 , \5355 , \5358 );
nor \U$4654 ( \5360 , \5346 , \5359 );
and \U$4655 ( \5361 , \740 , RIb557128_438);
and \U$4656 ( \5362 , RIb557038_436, \734 );
nor \U$4657 ( \5363 , \5361 , \5362 );
and \U$4658 ( \5364 , \4505 , RIb556fc0_435);
and \U$4659 ( \5365 , RIb5573f8_444, \698 );
nor \U$4660 ( \5366 , \5364 , \5365 );
and \U$4661 ( \5367 , \703 , RIb557380_443);
and \U$4662 ( \5368 , RIb557308_442, \705 );
nor \U$4663 ( \5369 , \5367 , \5368 );
nand \U$4664 ( \5370 , \5360 , \5363 , \5366 , \5369 );
_DC gf4a ( \5371_nGf4a , \5370 , \4513 );
nand \U$4665 ( \5372 , \5371_nGf4a , \4485 );
not \U$4666 ( \5373 , \5372 );
xor \U$4667 ( \5374 , \5251 , \5259 );
xor \U$4668 ( \5375 , \5374 , \5268 );
xor \U$4669 ( \5376 , \5278 , \5285 );
xor \U$4670 ( \5377 , \5376 , \5318 );
not \U$4671 ( \5378 , \5377 );
and \U$4672 ( \5379 , \5375 , \5378 );
nor \U$4673 ( \5380 , \5373 , \5379 );
not \U$4674 ( \5381 , \5380 );
not \U$4675 ( \5382 , \5256 );
not \U$4676 ( \5383 , \5091 );
or \U$4677 ( \5384 , \5382 , \5383 );
or \U$4678 ( \5385 , \5091 , \5256 );
nand \U$4679 ( \5386 , \5384 , \5385 );
xor \U$4680 ( \5387 , \5254 , \5257 );
nor \U$4681 ( \5388 , \5386 , \5387 );
not \U$4682 ( \5389 , \5388 );
not \U$4683 ( \5390 , \5259 );
nor \U$4684 ( \5391 , \5389 , \5390 );
not \U$4685 ( \5392 , \5391 );
or \U$4686 ( \5393 , \5392 , \4554 );
or \U$4687 ( \5394 , \5389 , \4554 );
nand \U$4688 ( \5395 , \5394 , \5390 );
nand \U$4689 ( \5396 , \5393 , \5395 );
not \U$4690 ( \5397 , \5396 );
nand \U$4691 ( \5398 , \4606_nG172a , \5140 );
or \U$4692 ( \5399 , \5093 , \4514_nG1821 );
nand \U$4693 ( \5400 , \5399 , \5248 );
and \U$4694 ( \5401 , \5398 , \5400 );
and \U$4695 ( \5402 , \5243 , \4514_nG1821 );
and \U$4696 ( \5403 , \4606_nG172a , \5143 );
nor \U$4697 ( \5404 , \5401 , \5402 , \5403 );
nor \U$4698 ( \5405 , \5397 , \5404 );
not \U$4699 ( \5406 , \5405 );
nand \U$4700 ( \5407 , \4800_nG140b , \4805 );
or \U$4701 ( \5408 , \4696 , \4903_nG1319 );
nand \U$4702 ( \5409 , \5408 , \4811 );
and \U$4703 ( \5410 , \5407 , \5409 );
and \U$4704 ( \5411 , \4807 , \4903_nG1319 );
and \U$4705 ( \5412 , \4800_nG140b , \4937 );
nor \U$4706 ( \5413 , \5410 , \5411 , \5412 );
and \U$4707 ( \5414 , \4683_nG1613 , \5071 );
or \U$4708 ( \5415 , \4928 , \4683_nG1613 );
nand \U$4709 ( \5416 , \5415 , \5074 );
nand \U$4710 ( \5417 , \4762_nG1506 , \4925 );
and \U$4711 ( \5418 , \5416 , \5417 );
and \U$4712 ( \5419 , \4762_nG1506 , \4930 );
nor \U$4713 ( \5420 , \5414 , \5418 , \5419 );
xor \U$4714 ( \5421 , \5413 , \5420 );
nand \U$4715 ( \5422 , \5065_nG112f , \4618 );
or \U$4716 ( \5423 , \4580 , \4876_nG1212 );
nand \U$4717 ( \5424 , \5423 , \4650 );
and \U$4718 ( \5425 , \5422 , \5424 );
and \U$4719 ( \5426 , \4653 , \4876_nG1212 );
and \U$4720 ( \5427 , \5065_nG112f , \4621 );
nor \U$4721 ( \5428 , \5425 , \5426 , \5427 );
and \U$4722 ( \5429 , \5421 , \5428 );
and \U$4723 ( \5430 , \5413 , \5420 );
or \U$4724 ( \5431 , \5429 , \5430 );
nor \U$4725 ( \5432 , \5406 , \5431 );
nand \U$4726 ( \5433 , \5381 , \5432 );
xor \U$4727 ( \5434 , \5345 , \5433 );
xor \U$4728 ( \5435 , \5237 , \5240 );
nand \U$4729 ( \5436 , \5311_nG1029 , \4485 );
and \U$4730 ( \5437 , \5435 , \5436 );
xor \U$4731 ( \5438 , \5271 , \5322 );
nor \U$4732 ( \5439 , \5437 , \5438 );
and \U$4733 ( \5440 , \5434 , \5439 );
and \U$4734 ( \5441 , \5345 , \5433 );
or \U$4735 ( \5442 , \5440 , \5441 );
or \U$4736 ( \5443 , \5340 , \5442 );
nand \U$4737 ( \5444 , \5339 , \5338 );
nand \U$4738 ( \5445 , \5443 , \5444 );
xor \U$4739 ( \5446 , \5133 , \5199 );
xor \U$4740 ( \5447 , \5446 , \5207 );
xor \U$4741 ( \5448 , \5225 , \5330 );
xor \U$4742 ( \5449 , \5447 , \5448 );
xor \U$4743 ( \5450 , \5445 , \5449 );
and \U$4744 ( \5451 , \4800_nG140b , \5071 );
or \U$4745 ( \5452 , \4928 , \4800_nG140b );
nand \U$4746 ( \5453 , \5452 , \5074 );
nand \U$4747 ( \5454 , \4903_nG1319 , \4925 );
and \U$4748 ( \5455 , \5453 , \5454 );
and \U$4749 ( \5456 , \4903_nG1319 , \4930 );
nor \U$4750 ( \5457 , \5451 , \5455 , \5456 );
and \U$4751 ( \5458 , \4762_nG1506 , \5143 );
or \U$4752 ( \5459 , \5093 , \4683_nG1613 );
nand \U$4753 ( \5460 , \5459 , \5248 );
nand \U$4754 ( \5461 , \4762_nG1506 , \5140 );
and \U$4755 ( \5462 , \5460 , \5461 );
and \U$4756 ( \5463 , \4683_nG1613 , \5243 );
nor \U$4757 ( \5464 , \5458 , \5462 , \5463 );
xor \U$4758 ( \5465 , \5457 , \5464 );
nand \U$4759 ( \5466 , \4876_nG1212 , \4805 );
or \U$4760 ( \5467 , \4696 , \5065_nG112f );
nand \U$4761 ( \5468 , \5467 , \4811 );
and \U$4762 ( \5469 , \5466 , \5468 );
and \U$4763 ( \5470 , \4807 , \5065_nG112f );
and \U$4764 ( \5471 , \4876_nG1212 , \4937 );
nor \U$4765 ( \5472 , \5469 , \5470 , \5471 );
and \U$4766 ( \5473 , \5465 , \5472 );
and \U$4767 ( \5474 , \5457 , \5464 );
or \U$4768 ( \5475 , \5473 , \5474 );
nand \U$4769 ( \5476 , \4606_nG172a , \5388 );
or \U$4770 ( \5477 , \5259 , \4514_nG1821 );
or \U$4771 ( \5478 , \5259 , \5387 );
nand \U$4772 ( \5479 , \5477 , \5478 );
and \U$4773 ( \5480 , \5476 , \5479 );
and \U$4774 ( \5481 , \5259 , \5387 );
and \U$4775 ( \5482 , \5481 , \4514_nG1821 );
and \U$4776 ( \5483 , \4606_nG172a , \5391 );
nor \U$4777 ( \5484 , \5480 , \5482 , \5483 );
not \U$4778 ( \5485 , \5484 );
or \U$4779 ( \5486 , \5253 , \4552_nG1933 );
or \U$4780 ( \5487 , \1173 , \4446_nG97d );
nand \U$4781 ( \5488 , \5487 , \4447 );
nor \U$4782 ( \5489 , \5253 , \5488 );
not \U$4783 ( \5490 , \5489 );
nand \U$4784 ( \5491 , \5254 , \5490 );
nand \U$4785 ( \5492 , \5486 , \5491 );
nand \U$4786 ( \5493 , \5485 , \5492 );
xor \U$4787 ( \5494 , \5475 , \5493 );
and \U$4788 ( \5495 , \4505 , RIb5567c8_418);
and \U$4789 ( \5496 , \695 , RIb556c78_428);
and \U$4790 ( \5497 , RIb556cf0_429, \719 );
nor \U$4791 ( \5498 , \5496 , \5497 );
and \U$4792 ( \5499 , \724 , RIb5569a8_422);
and \U$4793 ( \5500 , RIb556a20_423, \726 );
nor \U$4794 ( \5501 , \5499 , \5500 );
and \U$4795 ( \5502 , \710 , RIb556e58_432);
and \U$4796 ( \5503 , RIb556a98_424, \690 );
nor \U$4797 ( \5504 , \5502 , \5503 );
and \U$4798 ( \5505 , \716 , RIb556d68_430);
and \U$4799 ( \5506 , RIb556de0_431, \713 );
nor \U$4800 ( \5507 , \5505 , \5506 );
nand \U$4801 ( \5508 , \5498 , \5501 , \5504 , \5507 );
nor \U$4802 ( \5509 , \5495 , \5508 );
and \U$4803 ( \5510 , \703 , RIb556b88_426);
and \U$4804 ( \5511 , RIb556c00_427, \698 );
nor \U$4805 ( \5512 , \5510 , \5511 );
and \U$4806 ( \5513 , \740 , RIb556930_421);
and \U$4807 ( \5514 , RIb556840_419, \734 );
nor \U$4808 ( \5515 , \5513 , \5514 );
and \U$4809 ( \5516 , \738 , RIb5568b8_420);
and \U$4810 ( \5517 , RIb556b10_425, \705 );
nor \U$4811 ( \5518 , \5516 , \5517 );
nand \U$4812 ( \5519 , \5509 , \5512 , \5515 , \5518 );
_DC ge7a ( \5520_nGe7a , \5519 , \4513 );
and \U$4813 ( \5521 , \5520_nGe7a , \4566 );
and \U$4814 ( \5522 , \738 , RIb5580a0_471);
and \U$4815 ( \5523 , \724 , RIb558190_473);
and \U$4816 ( \5524 , RIb558208_474, \726 );
nor \U$4817 ( \5525 , \5523 , \5524 );
and \U$4818 ( \5526 , \710 , RIb558640_483);
and \U$4819 ( \5527 , RIb558280_475, \690 );
nor \U$4820 ( \5528 , \5526 , \5527 );
and \U$4821 ( \5529 , \716 , RIb558550_481);
and \U$4822 ( \5530 , RIb5585c8_482, \713 );
nor \U$4823 ( \5531 , \5529 , \5530 );
and \U$4824 ( \5532 , \695 , RIb558460_479);
and \U$4825 ( \5533 , RIb5584d8_480, \719 );
nor \U$4826 ( \5534 , \5532 , \5533 );
nand \U$4827 ( \5535 , \5525 , \5528 , \5531 , \5534 );
nor \U$4828 ( \5536 , \5522 , \5535 );
and \U$4829 ( \5537 , \740 , RIb558118_472);
and \U$4830 ( \5538 , RIb558028_470, \734 );
nor \U$4831 ( \5539 , \5537 , \5538 );
and \U$4832 ( \5540 , \4505 , RIb557fb0_469);
and \U$4833 ( \5541 , RIb5583e8_478, \698 );
nor \U$4834 ( \5542 , \5540 , \5541 );
and \U$4835 ( \5543 , \703 , RIb558370_477);
and \U$4836 ( \5544 , RIb5582f8_476, \705 );
nor \U$4837 ( \5545 , \5543 , \5544 );
nand \U$4838 ( \5546 , \5536 , \5539 , \5542 , \5545 );
_DC gdc3 ( \5547_nGdc3 , \5546 , \4513 );
and \U$4839 ( \5548 , \4559 , \5547_nGdc3 );
nand \U$4840 ( \5549 , \5520_nGe7a , \4557 );
or \U$4841 ( \5550 , \4527 , \5547_nGdc3 );
nand \U$4842 ( \5551 , \5550 , \4562 );
and \U$4843 ( \5552 , \5549 , \5551 );
nor \U$4844 ( \5553 , \5521 , \5548 , \5552 );
nand \U$4845 ( \5554 , \5371_nGf4a , \4618 );
or \U$4846 ( \5555 , \4580 , \5311_nG1029 );
nand \U$4847 ( \5556 , \5555 , \4650 );
and \U$4848 ( \5557 , \5554 , \5556 );
and \U$4849 ( \5558 , \4653 , \5311_nG1029 );
and \U$4850 ( \5559 , \5371_nGf4a , \4621 );
nor \U$4851 ( \5560 , \5557 , \5558 , \5559 );
and \U$4852 ( \5561 , \5553 , \5560 );
not \U$4853 ( \5562 , \5561 );
and \U$4854 ( \5563 , \726 , RIb557a10_457);
and \U$4855 ( \5564 , \695 , RIb557c68_462);
and \U$4856 ( \5565 , RIb557bf0_461, \698 );
nor \U$4857 ( \5566 , \5564 , \5565 );
and \U$4858 ( \5567 , \738 , RIb5578a8_454);
and \U$4859 ( \5568 , RIb557830_453, \734 );
nor \U$4860 ( \5569 , \5567 , \5568 );
and \U$4861 ( \5570 , \710 , RIb557e48_466);
and \U$4862 ( \5571 , RIb557dd0_465, \713 );
nor \U$4863 ( \5572 , \5570 , \5571 );
and \U$4864 ( \5573 , \716 , RIb557d58_464);
and \U$4865 ( \5574 , RIb557ce0_463, \719 );
nor \U$4866 ( \5575 , \5573 , \5574 );
nand \U$4867 ( \5576 , \5566 , \5569 , \5572 , \5575 );
nor \U$4868 ( \5577 , \5563 , \5576 );
and \U$4869 ( \5578 , \4505 , RIb5577b8_452);
and \U$4870 ( \5579 , RIb557b78_460, \703 );
nor \U$4871 ( \5580 , \5578 , \5579 );
and \U$4872 ( \5581 , \690 , RIb557a88_458);
and \U$4873 ( \5582 , RIb557b00_459, \705 );
nor \U$4874 ( \5583 , \5581 , \5582 );
and \U$4875 ( \5584 , \724 , RIb557998_456);
and \U$4876 ( \5585 , RIb557920_455, \740 );
nor \U$4877 ( \5586 , \5584 , \5585 );
nand \U$4878 ( \5587 , \5577 , \5580 , \5583 , \5586 );
_DC gcfd ( \5588_nGcfd , \5587 , \4513 );
nand \U$4879 ( \5589 , \5588_nGcfd , \4485 );
not \U$4880 ( \5590 , \5589 );
and \U$4881 ( \5591 , \5562 , \5590 );
nor \U$4882 ( \5592 , \5553 , \5560 );
nor \U$4883 ( \5593 , \5591 , \5592 );
and \U$4884 ( \5594 , \5494 , \5593 );
and \U$4885 ( \5595 , \5475 , \5493 );
or \U$4886 ( \5596 , \5594 , \5595 );
nand \U$4887 ( \5597 , \5547_nGdc3 , \4485 );
and \U$4888 ( \5598 , \5371_nGf4a , \4566 );
and \U$4889 ( \5599 , \4559 , \5520_nGe7a );
nand \U$4890 ( \5600 , \5371_nGf4a , \4557 );
or \U$4891 ( \5601 , \4527 , \5520_nGe7a );
nand \U$4892 ( \5602 , \5601 , \4562 );
and \U$4893 ( \5603 , \5600 , \5602 );
nor \U$4894 ( \5604 , \5598 , \5599 , \5603 );
xnor \U$4895 ( \5605 , \5597 , \5604 );
xor \U$4896 ( \5606 , \5596 , \5605 );
xor \U$4897 ( \5607 , \5413 , \5420 );
xor \U$4898 ( \5608 , \5607 , \5428 );
not \U$4899 ( \5609 , \5404 );
not \U$4900 ( \5610 , \5396 );
and \U$4901 ( \5611 , \5609 , \5610 );
and \U$4902 ( \5612 , \5404 , \5396 );
nor \U$4903 ( \5613 , \5611 , \5612 );
nand \U$4904 ( \5614 , \5520_nGe7a , \4485 );
and \U$4905 ( \5615 , \5311_nG1029 , \4566 );
and \U$4906 ( \5616 , \4559 , \5371_nGf4a );
nand \U$4907 ( \5617 , \5311_nG1029 , \4557 );
or \U$4908 ( \5618 , \4527 , \5371_nGf4a );
nand \U$4909 ( \5619 , \5618 , \4562 );
and \U$4910 ( \5620 , \5617 , \5619 );
nor \U$4911 ( \5621 , \5615 , \5616 , \5620 );
xnor \U$4912 ( \5622 , \5614 , \5621 );
xor \U$4913 ( \5623 , \5613 , \5622 );
xor \U$4914 ( \5624 , \5608 , \5623 );
and \U$4915 ( \5625 , \5606 , \5624 );
and \U$4916 ( \5626 , \5596 , \5605 );
or \U$4917 ( \5627 , \5625 , \5626 );
xor \U$4918 ( \5628 , \5413 , \5420 );
xor \U$4919 ( \5629 , \5628 , \5428 );
and \U$4920 ( \5630 , \5613 , \5629 );
xor \U$4921 ( \5631 , \5413 , \5420 );
xor \U$4922 ( \5632 , \5631 , \5428 );
and \U$4923 ( \5633 , \5622 , \5632 );
and \U$4924 ( \5634 , \5613 , \5622 );
or \U$4925 ( \5635 , \5630 , \5633 , \5634 );
not \U$4926 ( \5636 , \5635 );
nand \U$4927 ( \5637 , \4514_nG1821 , \5388 );
or \U$4928 ( \5638 , \5259 , \4552_nG1933 );
nand \U$4929 ( \5639 , \5638 , \5478 );
and \U$4930 ( \5640 , \5637 , \5639 );
and \U$4931 ( \5641 , \5481 , \4552_nG1933 );
and \U$4932 ( \5642 , \4514_nG1821 , \5391 );
nor \U$4933 ( \5643 , \5640 , \5641 , \5642 );
or \U$4934 ( \5644 , \5643 , \5254 );
and \U$4935 ( \5645 , \5643 , \5254 );
and \U$4936 ( \5646 , \4683_nG1613 , \5143 );
or \U$4937 ( \5647 , \5093 , \4606_nG172a );
nand \U$4938 ( \5648 , \5647 , \5248 );
nand \U$4939 ( \5649 , \4683_nG1613 , \5140 );
and \U$4940 ( \5650 , \5648 , \5649 );
and \U$4941 ( \5651 , \4606_nG172a , \5243 );
nor \U$4942 ( \5652 , \5646 , \5650 , \5651 );
nor \U$4943 ( \5653 , \5645 , \5652 );
not \U$4944 ( \5654 , \5653 );
nand \U$4945 ( \5655 , \5644 , \5654 );
not \U$4946 ( \5656 , \5655 );
nand \U$4947 ( \5657 , \4903_nG1319 , \4805 );
or \U$4948 ( \5658 , \4696 , \4876_nG1212 );
nand \U$4949 ( \5659 , \5658 , \4811 );
and \U$4950 ( \5660 , \5657 , \5659 );
and \U$4951 ( \5661 , \4807 , \4876_nG1212 );
and \U$4952 ( \5662 , \4903_nG1319 , \4937 );
nor \U$4953 ( \5663 , \5660 , \5661 , \5662 );
and \U$4954 ( \5664 , \4762_nG1506 , \5071 );
or \U$4955 ( \5665 , \4928 , \4762_nG1506 );
nand \U$4956 ( \5666 , \5665 , \5074 );
nand \U$4957 ( \5667 , \4800_nG140b , \4925 );
and \U$4958 ( \5668 , \5666 , \5667 );
and \U$4959 ( \5669 , \4800_nG140b , \4930 );
nor \U$4960 ( \5670 , \5664 , \5668 , \5669 );
xor \U$4961 ( \5671 , \5663 , \5670 );
nand \U$4962 ( \5672 , \5311_nG1029 , \4618 );
or \U$4963 ( \5673 , \4580 , \5065_nG112f );
nand \U$4964 ( \5674 , \5673 , \4650 );
and \U$4965 ( \5675 , \5672 , \5674 );
and \U$4966 ( \5676 , \4653 , \5065_nG112f );
and \U$4967 ( \5677 , \5311_nG1029 , \4621 );
nor \U$4968 ( \5678 , \5675 , \5676 , \5677 );
and \U$4969 ( \5679 , \5671 , \5678 );
and \U$4970 ( \5680 , \5663 , \5670 );
or \U$4971 ( \5681 , \5679 , \5680 );
nor \U$4972 ( \5682 , \5656 , \5681 );
not \U$4973 ( \5683 , \5682 );
and \U$4974 ( \5684 , \5636 , \5683 );
and \U$4975 ( \5685 , \5635 , \5682 );
nor \U$4976 ( \5686 , \5684 , \5685 );
xor \U$4977 ( \5687 , \5627 , \5686 );
xor \U$4978 ( \5688 , \5375 , \5378 );
not \U$4979 ( \5689 , \5688 );
not \U$4980 ( \5690 , \5372 );
and \U$4981 ( \5691 , \5689 , \5690 );
and \U$4982 ( \5692 , \5688 , \5372 );
nor \U$4983 ( \5693 , \5691 , \5692 );
not \U$4984 ( \5694 , \5693 );
or \U$4985 ( \5695 , \5431 , \5405 );
or \U$4986 ( \5696 , \5614 , \5621 );
nand \U$4987 ( \5697 , \5405 , \5431 );
nand \U$4988 ( \5698 , \5695 , \5696 , \5697 );
not \U$4989 ( \5699 , \5698 );
and \U$4990 ( \5700 , \5694 , \5699 );
and \U$4991 ( \5701 , \5693 , \5698 );
nor \U$4992 ( \5702 , \5700 , \5701 );
and \U$4993 ( \5703 , \5687 , \5702 );
and \U$4994 ( \5704 , \5627 , \5686 );
or \U$4995 ( \5705 , \5703 , \5704 );
not \U$4996 ( \5706 , \5682 );
nor \U$4997 ( \5707 , \5706 , \5635 );
not \U$4998 ( \5708 , \5438 );
xnor \U$4999 ( \5709 , \5436 , \5435 );
not \U$5000 ( \5710 , \5709 );
or \U$5001 ( \5711 , \5708 , \5710 );
or \U$5002 ( \5712 , \5709 , \5438 );
nand \U$5003 ( \5713 , \5711 , \5712 );
nand \U$5004 ( \5714 , \5707 , \5713 );
not \U$5005 ( \5715 , \5714 );
nor \U$5006 ( \5716 , \5713 , \5707 );
nor \U$5007 ( \5717 , \5715 , \5716 );
not \U$5008 ( \5718 , \5717 );
not \U$5009 ( \5719 , \5693 );
nand \U$5010 ( \5720 , \5719 , \5698 );
not \U$5011 ( \5721 , \5720 );
and \U$5012 ( \5722 , \5718 , \5721 );
and \U$5013 ( \5723 , \5717 , \5720 );
nor \U$5014 ( \5724 , \5722 , \5723 );
nand \U$5015 ( \5725 , \5705 , \5724 );
not \U$5016 ( \5726 , \5432 );
not \U$5017 ( \5727 , \5380 );
or \U$5018 ( \5728 , \5726 , \5727 );
or \U$5019 ( \5729 , \5380 , \5432 );
nand \U$5020 ( \5730 , \5728 , \5729 );
and \U$5021 ( \5731 , \5725 , \5730 );
nor \U$5022 ( \5732 , \5724 , \5705 );
nor \U$5023 ( \5733 , \5731 , \5732 );
not \U$5024 ( \5734 , \5733 );
not \U$5025 ( \5735 , \5241 );
not \U$5026 ( \5736 , \5436 );
nor \U$5027 ( \5737 , \5736 , \5323 );
not \U$5028 ( \5738 , \5737 );
and \U$5029 ( \5739 , \5735 , \5738 );
and \U$5030 ( \5740 , \5241 , \5737 );
nor \U$5031 ( \5741 , \5739 , \5740 );
xor \U$5032 ( \5742 , \5345 , \5433 );
xor \U$5033 ( \5743 , \5742 , \5439 );
nand \U$5034 ( \5744 , \5741 , \5743 );
not \U$5035 ( \5745 , \5744 );
nor \U$5036 ( \5746 , \5743 , \5741 );
nor \U$5037 ( \5747 , \5745 , \5746 );
not \U$5038 ( \5748 , \5747 );
or \U$5039 ( \5749 , \5716 , \5720 );
nand \U$5040 ( \5750 , \5749 , \5714 );
not \U$5041 ( \5751 , \5750 );
and \U$5042 ( \5752 , \5748 , \5751 );
and \U$5043 ( \5753 , \5747 , \5750 );
nor \U$5044 ( \5754 , \5752 , \5753 );
xor \U$5045 ( \5755 , \5734 , \5754 );
not \U$5046 ( \5756 , \5725 );
nor \U$5047 ( \5757 , \5756 , \5732 );
not \U$5048 ( \5758 , \5757 );
not \U$5049 ( \5759 , \5730 );
and \U$5050 ( \5760 , \5758 , \5759 );
and \U$5051 ( \5761 , \5757 , \5730 );
nor \U$5052 ( \5762 , \5760 , \5761 );
xor \U$5053 ( \5763 , \5627 , \5686 );
xor \U$5054 ( \5764 , \5763 , \5702 );
xor \U$5055 ( \5765 , \5596 , \5605 );
xor \U$5056 ( \5766 , \5765 , \5624 );
not \U$5057 ( \5767 , \5766 );
or \U$5058 ( \5768 , \5681 , \5655 );
or \U$5059 ( \5769 , \5597 , \5604 );
nand \U$5060 ( \5770 , \5655 , \5681 );
nand \U$5061 ( \5771 , \5768 , \5769 , \5770 );
nand \U$5062 ( \5772 , \5767 , \5771 );
or \U$5063 ( \5773 , \5764 , \5772 );
not \U$5064 ( \5774 , \5772 );
not \U$5065 ( \5775 , \5764 );
or \U$5066 ( \5776 , \5774 , \5775 );
nand \U$5067 ( \5777 , \5065_nG112f , \4805 );
or \U$5068 ( \5778 , \4696 , \5311_nG1029 );
nand \U$5069 ( \5779 , \5778 , \4811 );
and \U$5070 ( \5780 , \5777 , \5779 );
and \U$5071 ( \5781 , \4807 , \5311_nG1029 );
and \U$5072 ( \5782 , \5065_nG112f , \4937 );
nor \U$5073 ( \5783 , \5780 , \5781 , \5782 );
and \U$5074 ( \5784 , \4903_nG1319 , \5071 );
or \U$5075 ( \5785 , \4928 , \4903_nG1319 );
nand \U$5076 ( \5786 , \5785 , \5074 );
nand \U$5077 ( \5787 , \4876_nG1212 , \4925 );
and \U$5078 ( \5788 , \5786 , \5787 );
and \U$5079 ( \5789 , \4876_nG1212 , \4930 );
nor \U$5080 ( \5790 , \5784 , \5788 , \5789 );
xor \U$5081 ( \5791 , \5783 , \5790 );
nand \U$5082 ( \5792 , \5520_nGe7a , \4618 );
or \U$5083 ( \5793 , \4580 , \5371_nGf4a );
nand \U$5084 ( \5794 , \5793 , \4650 );
and \U$5085 ( \5795 , \5792 , \5794 );
and \U$5086 ( \5796 , \4653 , \5371_nGf4a );
and \U$5087 ( \5797 , \5520_nGe7a , \4621 );
nor \U$5088 ( \5798 , \5795 , \5796 , \5797 );
and \U$5089 ( \5799 , \5791 , \5798 );
and \U$5090 ( \5800 , \5783 , \5790 );
or \U$5091 ( \5801 , \5799 , \5800 );
nand \U$5092 ( \5802 , \4683_nG1613 , \5388 );
or \U$5093 ( \5803 , \5259 , \4606_nG172a );
nand \U$5094 ( \5804 , \5803 , \5478 );
and \U$5095 ( \5805 , \5802 , \5804 );
and \U$5096 ( \5806 , \5481 , \4606_nG172a );
and \U$5097 ( \5807 , \4683_nG1613 , \5391 );
nor \U$5098 ( \5808 , \5805 , \5806 , \5807 );
not \U$5099 ( \5809 , \5808 );
not \U$5100 ( \5810 , \5491 );
and \U$5101 ( \5811 , \4554 , \5810 );
and \U$5102 ( \5812 , \5489 , \4515 );
nand \U$5103 ( \5813 , \5488 , \5253 );
not \U$5104 ( \5814 , \5813 );
and \U$5105 ( \5815 , \4552_nG1933 , \5814 );
nor \U$5106 ( \5816 , \5811 , \5812 , \5815 );
not \U$5107 ( \5817 , \5816 );
and \U$5108 ( \5818 , \5809 , \5817 );
and \U$5109 ( \5819 , \5808 , \5816 );
nand \U$5110 ( \5820 , \4800_nG140b , \5140 );
or \U$5111 ( \5821 , \5093 , \4762_nG1506 );
nand \U$5112 ( \5822 , \5821 , \5248 );
and \U$5113 ( \5823 , \5820 , \5822 );
and \U$5114 ( \5824 , \5243 , \4762_nG1506 );
and \U$5115 ( \5825 , \4800_nG140b , \5143 );
nor \U$5116 ( \5826 , \5823 , \5824 , \5825 );
nor \U$5117 ( \5827 , \5819 , \5826 );
nor \U$5118 ( \5828 , \5818 , \5827 );
nor \U$5119 ( \5829 , \5801 , \5828 );
xor \U$5120 ( \5830 , \5663 , \5670 );
xor \U$5121 ( \5831 , \5830 , \5678 );
not \U$5122 ( \5832 , \5831 );
xor \U$5123 ( \5833 , \5829 , \5832 );
not \U$5124 ( \5834 , \5589 );
nor \U$5125 ( \5835 , \5561 , \5592 );
not \U$5126 ( \5836 , \5835 );
or \U$5127 ( \5837 , \5834 , \5836 );
or \U$5128 ( \5838 , \5835 , \5589 );
nand \U$5129 ( \5839 , \5837 , \5838 );
not \U$5130 ( \5840 , \5839 );
xor \U$5131 ( \5841 , \5457 , \5464 );
xor \U$5132 ( \5842 , \5841 , \5472 );
nor \U$5133 ( \5843 , \5840 , \5842 );
and \U$5134 ( \5844 , \5833 , \5843 );
and \U$5135 ( \5845 , \5829 , \5832 );
or \U$5136 ( \5846 , \5844 , \5845 );
not \U$5137 ( \5847 , \5846 );
not \U$5138 ( \5848 , \5605 );
or \U$5139 ( \5849 , \5652 , \5253 );
nand \U$5140 ( \5850 , \5253 , \5652 );
nand \U$5141 ( \5851 , \5849 , \5850 );
not \U$5142 ( \5852 , \5851 );
not \U$5143 ( \5853 , \5643 );
and \U$5144 ( \5854 , \5852 , \5853 );
and \U$5145 ( \5855 , \5851 , \5643 );
nor \U$5146 ( \5856 , \5854 , \5855 );
xor \U$5147 ( \5857 , \5848 , \5856 );
xor \U$5148 ( \5858 , \5475 , \5493 );
xor \U$5149 ( \5859 , \5858 , \5593 );
and \U$5150 ( \5860 , \5857 , \5859 );
and \U$5151 ( \5861 , \5848 , \5856 );
or \U$5152 ( \5862 , \5860 , \5861 );
nand \U$5153 ( \5863 , \5847 , \5862 );
nand \U$5154 ( \5864 , \5776 , \5863 );
nand \U$5155 ( \5865 , \5773 , \5864 );
and \U$5156 ( \5866 , \5762 , \5865 );
not \U$5157 ( \5867 , \5762 );
not \U$5158 ( \5868 , \5865 );
and \U$5159 ( \5869 , \5867 , \5868 );
xor \U$5160 ( \5870 , \5848 , \5856 );
xor \U$5161 ( \5871 , \5870 , \5859 );
not \U$5162 ( \5872 , \5484 );
not \U$5163 ( \5873 , \5492 );
and \U$5164 ( \5874 , \5872 , \5873 );
and \U$5165 ( \5875 , \5484 , \5492 );
nor \U$5166 ( \5876 , \5874 , \5875 );
and \U$5167 ( \5877 , \4876_nG1212 , \5071 );
or \U$5168 ( \5878 , \4928 , \4876_nG1212 );
nand \U$5169 ( \5879 , \5878 , \5074 );
nand \U$5170 ( \5880 , \5065_nG112f , \4925 );
and \U$5171 ( \5881 , \5879 , \5880 );
and \U$5172 ( \5882 , \5065_nG112f , \4930 );
nor \U$5173 ( \5883 , \5877 , \5881 , \5882 );
and \U$5174 ( \5884 , \4903_nG1319 , \5143 );
or \U$5175 ( \5885 , \5093 , \4800_nG140b );
nand \U$5176 ( \5886 , \5885 , \5248 );
nand \U$5177 ( \5887 , \4903_nG1319 , \5140 );
and \U$5178 ( \5888 , \5886 , \5887 );
and \U$5179 ( \5889 , \4800_nG140b , \5243 );
nor \U$5180 ( \5890 , \5884 , \5888 , \5889 );
xor \U$5181 ( \5891 , \5883 , \5890 );
nand \U$5182 ( \5892 , \5311_nG1029 , \4805 );
or \U$5183 ( \5893 , \4696 , \5371_nGf4a );
nand \U$5184 ( \5894 , \5893 , \4811 );
and \U$5185 ( \5895 , \5892 , \5894 );
and \U$5186 ( \5896 , \4807 , \5371_nGf4a );
and \U$5187 ( \5897 , \5311_nG1029 , \4937 );
nor \U$5188 ( \5898 , \5895 , \5896 , \5897 );
and \U$5189 ( \5899 , \5891 , \5898 );
and \U$5190 ( \5900 , \5883 , \5890 );
or \U$5191 ( \5901 , \5899 , \5900 );
and \U$5192 ( \5902 , \5588_nGcfd , \4566 );
and \U$5193 ( \5903 , RIb559450_513, \695 );
and \U$5194 ( \5904 , RIb559630_517, \710 );
and \U$5195 ( \5905 , \703 , RIb559360_511);
and \U$5196 ( \5906 , RIb5592e8_510, \705 );
nor \U$5197 ( \5907 , \5905 , \5906 );
and \U$5198 ( \5908 , RIb558fa0_503, \4505 );
and \U$5199 ( \5909 , \734 , RIb559018_504);
and \U$5200 ( \5910 , RIb5593d8_512, \698 );
nor \U$5201 ( \5911 , \5908 , \5909 , \5910 );
and \U$5202 ( \5912 , \738 , RIb559090_505);
and \U$5203 ( \5913 , RIb559108_506, \740 );
nor \U$5204 ( \5914 , \5912 , \5913 );
nand \U$5205 ( \5915 , \5907 , \5911 , \5914 );
nor \U$5206 ( \5916 , \5903 , \5904 , \5915 );
and \U$5207 ( \5917 , \716 , RIb559540_515);
and \U$5208 ( \5918 , RIb5594c8_514, \719 );
nor \U$5209 ( \5919 , \5917 , \5918 );
and \U$5210 ( \5920 , \690 , RIb559270_509);
and \U$5211 ( \5921 , RIb5591f8_508, \726 );
nor \U$5212 ( \5922 , \5920 , \5921 );
and \U$5213 ( \5923 , \713 , RIb5595b8_516);
and \U$5214 ( \5924 , RIb559180_507, \724 );
nor \U$5215 ( \5925 , \5923 , \5924 );
nand \U$5216 ( \5926 , \5916 , \5919 , \5922 , \5925 );
_DC gc6b ( \5927_nGc6b , \5926 , \4513 );
and \U$5217 ( \5928 , \4559 , \5927_nGc6b );
nand \U$5218 ( \5929 , \5588_nGcfd , \4557 );
or \U$5219 ( \5930 , \4527 , \5927_nGc6b );
nand \U$5220 ( \5931 , \5930 , \4562 );
and \U$5221 ( \5932 , \5929 , \5931 );
nor \U$5222 ( \5933 , \5902 , \5928 , \5932 );
nand \U$5223 ( \5934 , \5547_nGdc3 , \4618 );
or \U$5224 ( \5935 , \4580 , \5520_nGe7a );
nand \U$5225 ( \5936 , \5935 , \4650 );
and \U$5226 ( \5937 , \5934 , \5936 );
and \U$5227 ( \5938 , \4653 , \5520_nGe7a );
and \U$5228 ( \5939 , \5547_nGdc3 , \4621 );
nor \U$5229 ( \5940 , \5937 , \5938 , \5939 );
and \U$5230 ( \5941 , \5933 , \5940 );
not \U$5231 ( \5942 , \5941 );
and \U$5232 ( \5943 , \4505 , RIb5587a8_486);
and \U$5233 ( \5944 , \695 , RIb558c58_496);
and \U$5234 ( \5945 , RIb558cd0_497, \719 );
nor \U$5235 ( \5946 , \5944 , \5945 );
and \U$5236 ( \5947 , \724 , RIb558988_490);
and \U$5237 ( \5948 , RIb558a00_491, \726 );
nor \U$5238 ( \5949 , \5947 , \5948 );
and \U$5239 ( \5950 , \710 , RIb558e38_500);
and \U$5240 ( \5951 , RIb558a78_492, \690 );
nor \U$5241 ( \5952 , \5950 , \5951 );
and \U$5242 ( \5953 , \716 , RIb558d48_498);
and \U$5243 ( \5954 , RIb558dc0_499, \713 );
nor \U$5244 ( \5955 , \5953 , \5954 );
nand \U$5245 ( \5956 , \5946 , \5949 , \5952 , \5955 );
nor \U$5246 ( \5957 , \5943 , \5956 );
and \U$5247 ( \5958 , \703 , RIb558b68_494);
and \U$5248 ( \5959 , RIb558be0_495, \698 );
nor \U$5249 ( \5960 , \5958 , \5959 );
and \U$5250 ( \5961 , \740 , RIb558910_489);
and \U$5251 ( \5962 , RIb558820_487, \734 );
nor \U$5252 ( \5963 , \5961 , \5962 );
and \U$5253 ( \5964 , \738 , RIb558898_488);
and \U$5254 ( \5965 , RIb558af0_493, \705 );
nor \U$5255 ( \5966 , \5964 , \5965 );
nand \U$5256 ( \5967 , \5957 , \5960 , \5963 , \5966 );
_DC gbd0 ( \5968_nGbd0 , \5967 , \4513 );
nand \U$5257 ( \5969 , \5968_nGbd0 , \4485 );
not \U$5258 ( \5970 , \5969 );
and \U$5259 ( \5971 , \5942 , \5970 );
nor \U$5260 ( \5972 , \5933 , \5940 );
nor \U$5261 ( \5973 , \5971 , \5972 );
nand \U$5262 ( \5974 , \5901 , \5973 );
or \U$5263 ( \5975 , \5813 , \4515 );
or \U$5264 ( \5976 , \4514_nG1821 , \5491 );
or \U$5265 ( \5977 , \4606_nG172a , \5490 );
nand \U$5266 ( \5978 , \5975 , \5976 , \5977 );
not \U$5267 ( \5979 , \4762_nG1506 );
or \U$5268 ( \5980 , \5392 , \5979 );
not \U$5269 ( \5981 , \5481 );
or \U$5270 ( \5982 , \5262 , \5981 );
or \U$5271 ( \5983 , \5389 , \5979 );
or \U$5272 ( \5984 , \5259 , \4683_nG1613 );
nand \U$5273 ( \5985 , \5984 , \5478 );
nand \U$5274 ( \5986 , \5983 , \5985 );
nand \U$5275 ( \5987 , \5980 , \5982 , \5986 );
and \U$5276 ( \5988 , \5978 , \5987 );
and \U$5277 ( \5989 , \5974 , \5988 );
nor \U$5278 ( \5990 , \5973 , \5901 );
nor \U$5279 ( \5991 , \5989 , \5990 );
nand \U$5280 ( \5992 , \5876 , \5991 );
xor \U$5281 ( \5993 , \5783 , \5790 );
xor \U$5282 ( \5994 , \5993 , \5798 );
not \U$5283 ( \5995 , \5994 );
nand \U$5284 ( \5996 , \5927_nGc6b , \4485 );
and \U$5285 ( \5997 , \5547_nGdc3 , \4566 );
and \U$5286 ( \5998 , \4559 , \5588_nGcfd );
nand \U$5287 ( \5999 , \5547_nGdc3 , \4557 );
or \U$5288 ( \6000 , \4527 , \5588_nGcfd );
nand \U$5289 ( \6001 , \6000 , \4562 );
and \U$5290 ( \6002 , \5999 , \6001 );
nor \U$5291 ( \6003 , \5997 , \5998 , \6002 );
xor \U$5292 ( \6004 , \5996 , \6003 );
and \U$5293 ( \6005 , \5995 , \6004 );
and \U$5294 ( \6006 , \5992 , \6005 );
nor \U$5295 ( \6007 , \5991 , \5876 );
nor \U$5296 ( \6008 , \6006 , \6007 );
and \U$5297 ( \6009 , \5871 , \6008 );
not \U$5298 ( \6010 , \6009 );
not \U$5299 ( \6011 , \5839 );
not \U$5300 ( \6012 , \5842 );
and \U$5301 ( \6013 , \6011 , \6012 );
and \U$5302 ( \6014 , \5839 , \5842 );
nor \U$5303 ( \6015 , \6013 , \6014 );
not \U$5304 ( \6016 , \6015 );
not \U$5305 ( \6017 , \5828 );
or \U$5306 ( \6018 , \5801 , \6017 );
not \U$5307 ( \6019 , \5801 );
or \U$5308 ( \6020 , \5828 , \6019 );
or \U$5309 ( \6021 , \5996 , \6003 );
nand \U$5310 ( \6022 , \6018 , \6020 , \6021 );
nand \U$5311 ( \6023 , \6016 , \6022 );
not \U$5312 ( \6024 , \6023 );
and \U$5313 ( \6025 , \6010 , \6024 );
nor \U$5314 ( \6026 , \5871 , \6008 );
nor \U$5315 ( \6027 , \6025 , \6026 );
not \U$5316 ( \6028 , \5766 );
not \U$5317 ( \6029 , \5771 );
and \U$5318 ( \6030 , \6028 , \6029 );
and \U$5319 ( \6031 , \5766 , \5771 );
nor \U$5320 ( \6032 , \6030 , \6031 );
nor \U$5321 ( \6033 , \6027 , \6032 );
and \U$5322 ( \6034 , \6027 , \6032 );
or \U$5323 ( \6035 , \6033 , \6034 );
not \U$5324 ( \6036 , \6035 );
not \U$5325 ( \6037 , \5846 );
not \U$5326 ( \6038 , \5862 );
or \U$5327 ( \6039 , \6037 , \6038 );
or \U$5328 ( \6040 , \5862 , \5846 );
nand \U$5329 ( \6041 , \6039 , \6040 );
not \U$5330 ( \6042 , \6041 );
and \U$5331 ( \6043 , \6036 , \6042 );
and \U$5332 ( \6044 , \6035 , \6041 );
nor \U$5333 ( \6045 , \6043 , \6044 );
not \U$5334 ( \6046 , \6022 );
not \U$5335 ( \6047 , \6015 );
or \U$5336 ( \6048 , \6046 , \6047 );
or \U$5337 ( \6049 , \6015 , \6022 );
nand \U$5338 ( \6050 , \6048 , \6049 );
not \U$5339 ( \6051 , \5808 );
xor \U$5340 ( \6052 , \5816 , \5826 );
not \U$5341 ( \6053 , \6052 );
or \U$5342 ( \6054 , \6051 , \6053 );
or \U$5343 ( \6055 , \6052 , \5808 );
nand \U$5344 ( \6056 , \6054 , \6055 );
nand \U$5345 ( \6057 , \5371_nGf4a , \4805 );
or \U$5346 ( \6058 , \4696 , \5520_nGe7a );
nand \U$5347 ( \6059 , \6058 , \4811 );
and \U$5348 ( \6060 , \6057 , \6059 );
and \U$5349 ( \6061 , \4807 , \5520_nGe7a );
and \U$5350 ( \6062 , \5371_nGf4a , \4937 );
nor \U$5351 ( \6063 , \6060 , \6061 , \6062 );
and \U$5352 ( \6064 , \5065_nG112f , \5071 );
or \U$5353 ( \6065 , \4928 , \5065_nG112f );
nand \U$5354 ( \6066 , \6065 , \5074 );
nand \U$5355 ( \6067 , \5311_nG1029 , \4925 );
and \U$5356 ( \6068 , \6066 , \6067 );
and \U$5357 ( \6069 , \5311_nG1029 , \4930 );
nor \U$5358 ( \6070 , \6064 , \6068 , \6069 );
xor \U$5359 ( \6071 , \6063 , \6070 );
nand \U$5360 ( \6072 , \5588_nGcfd , \4618 );
or \U$5361 ( \6073 , \4580 , \5547_nGdc3 );
nand \U$5362 ( \6074 , \6073 , \4650 );
and \U$5363 ( \6075 , \6072 , \6074 );
and \U$5364 ( \6076 , \4653 , \5547_nGdc3 );
and \U$5365 ( \6077 , \5588_nGcfd , \4621 );
nor \U$5366 ( \6078 , \6075 , \6076 , \6077 );
and \U$5367 ( \6079 , \6071 , \6078 );
and \U$5368 ( \6080 , \6063 , \6070 );
or \U$5369 ( \6081 , \6079 , \6080 );
nand \U$5370 ( \6082 , \4800_nG140b , \5388 );
or \U$5371 ( \6083 , \5259 , \4762_nG1506 );
nand \U$5372 ( \6084 , \6083 , \5478 );
and \U$5373 ( \6085 , \6082 , \6084 );
and \U$5374 ( \6086 , \5481 , \4762_nG1506 );
and \U$5375 ( \6087 , \4800_nG140b , \5391 );
nor \U$5376 ( \6088 , \6085 , \6086 , \6087 );
and \U$5377 ( \6089 , \4628 , \5810 );
and \U$5378 ( \6090 , \5489 , \5262 );
and \U$5379 ( \6091 , \4606_nG172a , \5814 );
nor \U$5380 ( \6092 , \6089 , \6090 , \6091 );
xor \U$5381 ( \6093 , \6088 , \6092 );
nand \U$5382 ( \6094 , \4876_nG1212 , \5140 );
or \U$5383 ( \6095 , \5093 , \4903_nG1319 );
nand \U$5384 ( \6096 , \6095 , \5248 );
and \U$5385 ( \6097 , \6094 , \6096 );
and \U$5386 ( \6098 , \5243 , \4903_nG1319 );
and \U$5387 ( \6099 , \4876_nG1212 , \5143 );
nor \U$5388 ( \6100 , \6097 , \6098 , \6099 );
and \U$5389 ( \6101 , \6093 , \6100 );
and \U$5390 ( \6102 , \6088 , \6092 );
or \U$5391 ( \6103 , \6101 , \6102 );
nor \U$5392 ( \6104 , \6081 , \6103 );
and \U$5393 ( \6105 , \6056 , \6104 );
xor \U$5394 ( \6106 , \6050 , \6105 );
not \U$5395 ( \6107 , \6005 );
not \U$5396 ( \6108 , \6007 );
nand \U$5397 ( \6109 , \6108 , \5992 );
not \U$5398 ( \6110 , \6109 );
or \U$5399 ( \6111 , \6107 , \6110 );
or \U$5400 ( \6112 , \6109 , \6005 );
nand \U$5401 ( \6113 , \6111 , \6112 );
and \U$5402 ( \6114 , \6106 , \6113 );
and \U$5403 ( \6115 , \6050 , \6105 );
or \U$5404 ( \6116 , \6114 , \6115 );
xor \U$5405 ( \6117 , \5829 , \5832 );
xor \U$5406 ( \6118 , \6117 , \5843 );
xor \U$5407 ( \6119 , \6116 , \6118 );
not \U$5408 ( \6120 , \6023 );
nor \U$5409 ( \6121 , \6026 , \6009 );
not \U$5410 ( \6122 , \6121 );
or \U$5411 ( \6123 , \6120 , \6122 );
or \U$5412 ( \6124 , \6121 , \6023 );
nand \U$5413 ( \6125 , \6123 , \6124 );
and \U$5414 ( \6126 , \6119 , \6125 );
and \U$5415 ( \6127 , \6116 , \6118 );
or \U$5416 ( \6128 , \6126 , \6127 );
xor \U$5417 ( \6129 , \6045 , \6128 );
xor \U$5418 ( \6130 , \6116 , \6118 );
xor \U$5419 ( \6131 , \6130 , \6125 );
xor \U$5420 ( \6132 , \5978 , \5987 );
not \U$5421 ( \6133 , \6132 );
not \U$5422 ( \6134 , \6103 );
or \U$5423 ( \6135 , \6081 , \6134 );
not \U$5424 ( \6136 , \6081 );
or \U$5425 ( \6137 , \6103 , \6136 );
and \U$5426 ( \6138 , \4505 , RIb559f90_537);
and \U$5427 ( \6139 , \724 , RIb55a170_541);
and \U$5428 ( \6140 , RIb55a1e8_542, \726 );
nor \U$5429 ( \6141 , \6139 , \6140 );
and \U$5430 ( \6142 , \710 , RIb55a620_551);
and \U$5431 ( \6143 , RIb55a260_543, \690 );
nor \U$5432 ( \6144 , \6142 , \6143 );
and \U$5433 ( \6145 , \716 , RIb55a530_549);
and \U$5434 ( \6146 , RIb55a5a8_550, \713 );
nor \U$5435 ( \6147 , \6145 , \6146 );
and \U$5436 ( \6148 , \695 , RIb55a440_547);
and \U$5437 ( \6149 , RIb55a4b8_548, \719 );
nor \U$5438 ( \6150 , \6148 , \6149 );
nand \U$5439 ( \6151 , \6141 , \6144 , \6147 , \6150 );
nor \U$5440 ( \6152 , \6138 , \6151 );
and \U$5441 ( \6153 , \703 , RIb55a350_545);
and \U$5442 ( \6154 , RIb55a3c8_546, \698 );
nor \U$5443 ( \6155 , \6153 , \6154 );
and \U$5444 ( \6156 , \740 , RIb55a0f8_540);
and \U$5445 ( \6157 , RIb55a008_538, \734 );
nor \U$5446 ( \6158 , \6156 , \6157 );
and \U$5447 ( \6159 , \738 , RIb55a080_539);
and \U$5448 ( \6160 , RIb55a2d8_544, \705 );
nor \U$5449 ( \6161 , \6159 , \6160 );
nand \U$5450 ( \6162 , \6152 , \6155 , \6158 , \6161 );
_DC gb55 ( \6163_nGb55 , \6162 , \4513 );
nand \U$5451 ( \6164 , \6163_nGb55 , \4485 );
and \U$5452 ( \6165 , \5927_nGc6b , \4566 );
and \U$5453 ( \6166 , \4559 , \5968_nGbd0 );
nand \U$5454 ( \6167 , \5927_nGc6b , \4557 );
or \U$5455 ( \6168 , \4527 , \5968_nGbd0 );
nand \U$5456 ( \6169 , \6168 , \4562 );
and \U$5457 ( \6170 , \6167 , \6169 );
nor \U$5458 ( \6171 , \6165 , \6166 , \6170 );
or \U$5459 ( \6172 , \6164 , \6171 );
nand \U$5460 ( \6173 , \6135 , \6137 , \6172 );
not \U$5461 ( \6174 , \6173 );
or \U$5462 ( \6175 , \6133 , \6174 );
or \U$5463 ( \6176 , \6173 , \6132 );
not \U$5464 ( \6177 , \5969 );
nor \U$5465 ( \6178 , \5941 , \5972 );
not \U$5466 ( \6179 , \6178 );
or \U$5467 ( \6180 , \6177 , \6179 );
or \U$5468 ( \6181 , \6178 , \5969 );
nand \U$5469 ( \6182 , \6180 , \6181 );
nand \U$5470 ( \6183 , \6176 , \6182 );
nand \U$5471 ( \6184 , \6175 , \6183 );
xor \U$5472 ( \6185 , \5995 , \6004 );
xor \U$5473 ( \6186 , \6184 , \6185 );
xor \U$5474 ( \6187 , \5883 , \5890 );
xor \U$5475 ( \6188 , \6187 , \5898 );
xor \U$5476 ( \6189 , \6063 , \6070 );
xor \U$5477 ( \6190 , \6189 , \6078 );
xor \U$5478 ( \6191 , \6088 , \6092 );
xor \U$5479 ( \6192 , \6191 , \6100 );
xor \U$5480 ( \6193 , \6190 , \6192 );
xnor \U$5481 ( \6194 , \6164 , \6171 );
and \U$5482 ( \6195 , \6193 , \6194 );
and \U$5483 ( \6196 , \6190 , \6192 );
or \U$5484 ( \6197 , \6195 , \6196 );
xor \U$5485 ( \6198 , \6188 , \6197 );
and \U$5486 ( \6199 , \5311_nG1029 , \5071 );
or \U$5487 ( \6200 , \4928 , \5311_nG1029 );
nand \U$5488 ( \6201 , \6200 , \5074 );
nand \U$5489 ( \6202 , \5371_nGf4a , \4925 );
and \U$5490 ( \6203 , \6201 , \6202 );
and \U$5491 ( \6204 , \5371_nGf4a , \4930 );
nor \U$5492 ( \6205 , \6199 , \6203 , \6204 );
and \U$5493 ( \6206 , \5065_nG112f , \5143 );
or \U$5494 ( \6207 , \5093 , \4876_nG1212 );
nand \U$5495 ( \6208 , \6207 , \5248 );
nand \U$5496 ( \6209 , \5065_nG112f , \5140 );
and \U$5497 ( \6210 , \6208 , \6209 );
and \U$5498 ( \6211 , \4876_nG1212 , \5243 );
nor \U$5499 ( \6212 , \6206 , \6210 , \6211 );
xor \U$5500 ( \6213 , \6205 , \6212 );
nand \U$5501 ( \6214 , \5520_nGe7a , \4805 );
or \U$5502 ( \6215 , \4696 , \5547_nGdc3 );
nand \U$5503 ( \6216 , \6215 , \4811 );
and \U$5504 ( \6217 , \6214 , \6216 );
and \U$5505 ( \6218 , \4807 , \5547_nGdc3 );
and \U$5506 ( \6219 , \5520_nGe7a , \4937 );
nor \U$5507 ( \6220 , \6217 , \6218 , \6219 );
and \U$5508 ( \6221 , \6213 , \6220 );
and \U$5509 ( \6222 , \6205 , \6212 );
or \U$5510 ( \6223 , \6221 , \6222 );
nand \U$5511 ( \6224 , \4903_nG1319 , \5388 );
or \U$5512 ( \6225 , \5259 , \4800_nG140b );
nand \U$5513 ( \6226 , \6225 , \5478 );
and \U$5514 ( \6227 , \6224 , \6226 );
and \U$5515 ( \6228 , \5481 , \4800_nG140b );
and \U$5516 ( \6229 , \4903_nG1319 , \5391 );
nor \U$5517 ( \6230 , \6227 , \6228 , \6229 );
not \U$5518 ( \6231 , \6230 );
or \U$5519 ( \6232 , \5813 , \5262 );
or \U$5520 ( \6233 , \4683_nG1613 , \5491 );
or \U$5521 ( \6234 , \4762_nG1506 , \5490 );
nand \U$5522 ( \6235 , \6232 , \6233 , \6234 );
nand \U$5523 ( \6236 , \6231 , \6235 );
xor \U$5524 ( \6237 , \6223 , \6236 );
and \U$5525 ( \6238 , \5968_nGbd0 , \4566 );
and \U$5526 ( \6239 , \4559 , \6163_nGb55 );
nand \U$5527 ( \6240 , \5968_nGbd0 , \4557 );
or \U$5528 ( \6241 , \4527 , \6163_nGb55 );
nand \U$5529 ( \6242 , \6241 , \4562 );
and \U$5530 ( \6243 , \6240 , \6242 );
nor \U$5531 ( \6244 , \6238 , \6239 , \6243 );
nand \U$5532 ( \6245 , \5927_nGc6b , \4618 );
or \U$5533 ( \6246 , \4580 , \5588_nGcfd );
nand \U$5534 ( \6247 , \6246 , \4650 );
and \U$5535 ( \6248 , \6245 , \6247 );
and \U$5536 ( \6249 , \4653 , \5588_nGcfd );
and \U$5537 ( \6250 , \5927_nGc6b , \4621 );
nor \U$5538 ( \6251 , \6248 , \6249 , \6250 );
and \U$5539 ( \6252 , \6244 , \6251 );
not \U$5540 ( \6253 , \6252 );
and \U$5541 ( \6254 , \738 , RIb559888_522);
and \U$5542 ( \6255 , \724 , RIb559978_524);
and \U$5543 ( \6256 , RIb5599f0_525, \726 );
nor \U$5544 ( \6257 , \6255 , \6256 );
and \U$5545 ( \6258 , \710 , RIb559e28_534);
and \U$5546 ( \6259 , RIb559a68_526, \690 );
nor \U$5547 ( \6260 , \6258 , \6259 );
and \U$5548 ( \6261 , \716 , RIb559d38_532);
and \U$5549 ( \6262 , RIb559db0_533, \713 );
nor \U$5550 ( \6263 , \6261 , \6262 );
and \U$5551 ( \6264 , \695 , RIb559c48_530);
and \U$5552 ( \6265 , RIb559cc0_531, \719 );
nor \U$5553 ( \6266 , \6264 , \6265 );
nand \U$5554 ( \6267 , \6257 , \6260 , \6263 , \6266 );
nor \U$5555 ( \6268 , \6254 , \6267 );
and \U$5556 ( \6269 , \740 , RIb559900_523);
and \U$5557 ( \6270 , RIb559810_521, \734 );
nor \U$5558 ( \6271 , \6269 , \6270 );
and \U$5559 ( \6272 , \4505 , RIb559798_520);
and \U$5560 ( \6273 , RIb559bd0_529, \698 );
nor \U$5561 ( \6274 , \6272 , \6273 );
and \U$5562 ( \6275 , \703 , RIb559b58_528);
and \U$5563 ( \6276 , RIb559ae0_527, \705 );
nor \U$5564 ( \6277 , \6275 , \6276 );
nand \U$5565 ( \6278 , \6268 , \6271 , \6274 , \6277 );
_DC gadc ( \6279_nGadc , \6278 , \4513 );
nand \U$5566 ( \6280 , \6279_nGadc , \4485 );
not \U$5567 ( \6281 , \6280 );
and \U$5568 ( \6282 , \6253 , \6281 );
nor \U$5569 ( \6283 , \6244 , \6251 );
nor \U$5570 ( \6284 , \6282 , \6283 );
and \U$5571 ( \6285 , \6237 , \6284 );
and \U$5572 ( \6286 , \6223 , \6236 );
or \U$5573 ( \6287 , \6285 , \6286 );
and \U$5574 ( \6288 , \6198 , \6287 );
and \U$5575 ( \6289 , \6188 , \6197 );
nor \U$5576 ( \6290 , \6288 , \6289 );
and \U$5577 ( \6291 , \6186 , \6290 );
and \U$5578 ( \6292 , \6184 , \6185 );
or \U$5579 ( \6293 , \6291 , \6292 );
xor \U$5580 ( \6294 , \6056 , \6104 );
not \U$5581 ( \6295 , \5988 );
not \U$5582 ( \6296 , \5990 );
nand \U$5583 ( \6297 , \6296 , \5974 );
not \U$5584 ( \6298 , \6297 );
or \U$5585 ( \6299 , \6295 , \6298 );
or \U$5586 ( \6300 , \6297 , \5988 );
nand \U$5587 ( \6301 , \6299 , \6300 );
and \U$5588 ( \6302 , \6294 , \6301 );
xor \U$5589 ( \6303 , \6293 , \6302 );
xor \U$5590 ( \6304 , \6050 , \6105 );
xor \U$5591 ( \6305 , \6304 , \6113 );
and \U$5592 ( \6306 , \6303 , \6305 );
and \U$5593 ( \6307 , \6293 , \6302 );
or \U$5594 ( \6308 , \6306 , \6307 );
xor \U$5595 ( \6309 , \6131 , \6308 );
xor \U$5596 ( \6310 , \6293 , \6302 );
xor \U$5597 ( \6311 , \6310 , \6305 );
xor \U$5598 ( \6312 , \6294 , \6301 );
xor \U$5599 ( \6313 , \6184 , \6185 );
xor \U$5600 ( \6314 , \6313 , \6290 );
and \U$5601 ( \6315 , \6312 , \6314 );
nand \U$5602 ( \6316 , \4876_nG1212 , \5388 );
or \U$5603 ( \6317 , \5259 , \4903_nG1319 );
nand \U$5604 ( \6318 , \6317 , \5478 );
and \U$5605 ( \6319 , \6316 , \6318 );
and \U$5606 ( \6320 , \5481 , \4903_nG1319 );
and \U$5607 ( \6321 , \4876_nG1212 , \5391 );
nor \U$5608 ( \6322 , \6319 , \6320 , \6321 );
and \U$5609 ( \6323 , \5979 , \5810 );
not \U$5610 ( \6324 , \4800_nG140b );
and \U$5611 ( \6325 , \5489 , \6324 );
and \U$5612 ( \6326 , \4762_nG1506 , \5814 );
nor \U$5613 ( \6327 , \6323 , \6325 , \6326 );
xor \U$5614 ( \6328 , \6322 , \6327 );
nand \U$5615 ( \6329 , \5311_nG1029 , \5140 );
or \U$5616 ( \6330 , \5093 , \5065_nG112f );
nand \U$5617 ( \6331 , \6330 , \5248 );
and \U$5618 ( \6332 , \6329 , \6331 );
and \U$5619 ( \6333 , \5243 , \5065_nG112f );
and \U$5620 ( \6334 , \5311_nG1029 , \5143 );
nor \U$5621 ( \6335 , \6332 , \6333 , \6334 );
and \U$5622 ( \6336 , \6328 , \6335 );
and \U$5623 ( \6337 , \6322 , \6327 );
or \U$5624 ( \6338 , \6336 , \6337 );
not \U$5625 ( \6339 , \6338 );
nand \U$5626 ( \6340 , \5547_nGdc3 , \4805 );
or \U$5627 ( \6341 , \4696 , \5588_nGcfd );
nand \U$5628 ( \6342 , \6341 , \4811 );
and \U$5629 ( \6343 , \6340 , \6342 );
and \U$5630 ( \6344 , \4807 , \5588_nGcfd );
and \U$5631 ( \6345 , \5547_nGdc3 , \4937 );
nor \U$5632 ( \6346 , \6343 , \6344 , \6345 );
and \U$5633 ( \6347 , \5371_nGf4a , \5071 );
or \U$5634 ( \6348 , \4928 , \5371_nGf4a );
nand \U$5635 ( \6349 , \6348 , \5074 );
nand \U$5636 ( \6350 , \5520_nGe7a , \4925 );
and \U$5637 ( \6351 , \6349 , \6350 );
and \U$5638 ( \6352 , \5520_nGe7a , \4930 );
nor \U$5639 ( \6353 , \6347 , \6351 , \6352 );
xor \U$5640 ( \6354 , \6346 , \6353 );
nand \U$5641 ( \6355 , \5968_nGbd0 , \4618 );
or \U$5642 ( \6356 , \4580 , \5927_nGc6b );
nand \U$5643 ( \6357 , \6356 , \4650 );
and \U$5644 ( \6358 , \6355 , \6357 );
and \U$5645 ( \6359 , \4653 , \5927_nGc6b );
and \U$5646 ( \6360 , \5968_nGbd0 , \4621 );
nor \U$5647 ( \6361 , \6358 , \6359 , \6360 );
and \U$5648 ( \6362 , \6354 , \6361 );
and \U$5649 ( \6363 , \6346 , \6353 );
or \U$5650 ( \6364 , \6362 , \6363 );
not \U$5651 ( \6365 , \6364 );
nand \U$5652 ( \6366 , \6339 , \6365 );
xor \U$5653 ( \6367 , \6190 , \6192 );
xor \U$5654 ( \6368 , \6367 , \6194 );
and \U$5655 ( \6369 , \6366 , \6368 );
xor \U$5656 ( \6370 , \6205 , \6212 );
xor \U$5657 ( \6371 , \6370 , \6220 );
not \U$5658 ( \6372 , \6371 );
not \U$5659 ( \6373 , \6280 );
nor \U$5660 ( \6374 , \6252 , \6283 );
not \U$5661 ( \6375 , \6374 );
or \U$5662 ( \6376 , \6373 , \6375 );
or \U$5663 ( \6377 , \6374 , \6280 );
nand \U$5664 ( \6378 , \6376 , \6377 );
nand \U$5665 ( \6379 , \6372 , \6378 );
xor \U$5666 ( \6380 , \6190 , \6192 );
xor \U$5667 ( \6381 , \6380 , \6194 );
and \U$5668 ( \6382 , \6379 , \6381 );
and \U$5669 ( \6383 , \6366 , \6379 );
or \U$5670 ( \6384 , \6369 , \6382 , \6383 );
xnor \U$5671 ( \6385 , \6173 , \6182 );
not \U$5672 ( \6386 , \6385 );
not \U$5673 ( \6387 , \6132 );
and \U$5674 ( \6388 , \6386 , \6387 );
and \U$5675 ( \6389 , \6385 , \6132 );
nor \U$5676 ( \6390 , \6388 , \6389 );
xor \U$5677 ( \6391 , \6384 , \6390 );
xor \U$5678 ( \6392 , \6188 , \6197 );
xor \U$5679 ( \6393 , \6392 , \6287 );
and \U$5680 ( \6394 , \6391 , \6393 );
and \U$5681 ( \6395 , \6384 , \6390 );
or \U$5682 ( \6396 , \6394 , \6395 );
not \U$5683 ( \6397 , \6396 );
xor \U$5684 ( \6398 , \6184 , \6185 );
xor \U$5685 ( \6399 , \6398 , \6290 );
and \U$5686 ( \6400 , \6397 , \6399 );
and \U$5687 ( \6401 , \6312 , \6397 );
or \U$5688 ( \6402 , \6315 , \6400 , \6401 );
xor \U$5689 ( \6403 , \6311 , \6402 );
xor \U$5690 ( \6404 , \6184 , \6185 );
xor \U$5691 ( \6405 , \6404 , \6290 );
xor \U$5692 ( \6406 , \6312 , \6397 );
xor \U$5693 ( \6407 , \6405 , \6406 );
xor \U$5694 ( \6408 , \6384 , \6390 );
xor \U$5695 ( \6409 , \6408 , \6393 );
not \U$5696 ( \6410 , \6378 );
not \U$5697 ( \6411 , \6371 );
and \U$5698 ( \6412 , \6410 , \6411 );
and \U$5699 ( \6413 , \6378 , \6371 );
nor \U$5700 ( \6414 , \6412 , \6413 );
not \U$5701 ( \6415 , \6414 );
or \U$5702 ( \6416 , \6364 , \6339 );
or \U$5703 ( \6417 , \6338 , \6365 );
and \U$5704 ( \6418 , \738 , RIb55a878_556);
and \U$5705 ( \6419 , \724 , RIb55a968_558);
and \U$5706 ( \6420 , RIb55a9e0_559, \726 );
nor \U$5707 ( \6421 , \6419 , \6420 );
and \U$5708 ( \6422 , \716 , RIb55ad28_566);
and \U$5709 ( \6423 , RIb55ada0_567, \713 );
nor \U$5710 ( \6424 , \6422 , \6423 );
and \U$5711 ( \6425 , \710 , RIb55ae18_568);
and \U$5712 ( \6426 , RIb55abc0_563, \698 );
nor \U$5713 ( \6427 , \6425 , \6426 );
and \U$5714 ( \6428 , \695 , RIb55ac38_564);
and \U$5715 ( \6429 , RIb55acb0_565, \719 );
nor \U$5716 ( \6430 , \6428 , \6429 );
nand \U$5717 ( \6431 , \6421 , \6424 , \6427 , \6430 );
nor \U$5718 ( \6432 , \6418 , \6431 );
and \U$5719 ( \6433 , \690 , RIb55aa58_560);
and \U$5720 ( \6434 , RIb55aad0_561, \705 );
nor \U$5721 ( \6435 , \6433 , \6434 );
and \U$5722 ( \6436 , \740 , RIb55a8f0_557);
and \U$5723 ( \6437 , RIb55a800_555, \734 );
nor \U$5724 ( \6438 , \6436 , \6437 );
and \U$5725 ( \6439 , \4505 , RIb55a788_554);
and \U$5726 ( \6440 , RIb55ab48_562, \703 );
nor \U$5727 ( \6441 , \6439 , \6440 );
nand \U$5728 ( \6442 , \6432 , \6435 , \6438 , \6441 );
_DC ga88 ( \6443_nGa88 , \6442 , \4513 );
nand \U$5729 ( \6444 , \6443_nGa88 , \4485 );
and \U$5730 ( \6445 , \6163_nGb55 , \4566 );
and \U$5731 ( \6446 , \4559 , \6279_nGadc );
nand \U$5732 ( \6447 , \6163_nGb55 , \4557 );
or \U$5733 ( \6448 , \4527 , \6279_nGadc );
nand \U$5734 ( \6449 , \6448 , \4562 );
and \U$5735 ( \6450 , \6447 , \6449 );
nor \U$5736 ( \6451 , \6445 , \6446 , \6450 );
or \U$5737 ( \6452 , \6444 , \6451 );
nand \U$5738 ( \6453 , \6416 , \6417 , \6452 );
nand \U$5739 ( \6454 , \6415 , \6453 );
xor \U$5740 ( \6455 , \6223 , \6236 );
xor \U$5741 ( \6456 , \6455 , \6284 );
xor \U$5742 ( \6457 , \6454 , \6456 );
xor \U$5743 ( \6458 , \6346 , \6353 );
xor \U$5744 ( \6459 , \6458 , \6361 );
xor \U$5745 ( \6460 , \6322 , \6327 );
xor \U$5746 ( \6461 , \6460 , \6335 );
xor \U$5747 ( \6462 , \6459 , \6461 );
xnor \U$5748 ( \6463 , \6444 , \6451 );
and \U$5749 ( \6464 , \6462 , \6463 );
and \U$5750 ( \6465 , \6459 , \6461 );
or \U$5751 ( \6466 , \6464 , \6465 );
not \U$5752 ( \6467 , \6230 );
not \U$5753 ( \6468 , \6235 );
and \U$5754 ( \6469 , \6467 , \6468 );
and \U$5755 ( \6470 , \6230 , \6235 );
nor \U$5756 ( \6471 , \6469 , \6470 );
xor \U$5757 ( \6472 , \6466 , \6471 );
and \U$5758 ( \6473 , \5520_nGe7a , \5071 );
or \U$5759 ( \6474 , \4928 , \5520_nGe7a );
nand \U$5760 ( \6475 , \6474 , \5074 );
nand \U$5761 ( \6476 , \5547_nGdc3 , \4925 );
and \U$5762 ( \6477 , \6475 , \6476 );
and \U$5763 ( \6478 , \5547_nGdc3 , \4930 );
nor \U$5764 ( \6479 , \6473 , \6477 , \6478 );
and \U$5765 ( \6480 , \5371_nGf4a , \5143 );
or \U$5766 ( \6481 , \5093 , \5311_nG1029 );
nand \U$5767 ( \6482 , \6481 , \5248 );
nand \U$5768 ( \6483 , \5371_nGf4a , \5140 );
and \U$5769 ( \6484 , \6482 , \6483 );
and \U$5770 ( \6485 , \5311_nG1029 , \5243 );
nor \U$5771 ( \6486 , \6480 , \6484 , \6485 );
xor \U$5772 ( \6487 , \6479 , \6486 );
nand \U$5773 ( \6488 , \5588_nGcfd , \4805 );
or \U$5774 ( \6489 , \4696 , \5927_nGc6b );
nand \U$5775 ( \6490 , \6489 , \4811 );
and \U$5776 ( \6491 , \6488 , \6490 );
and \U$5777 ( \6492 , \4807 , \5927_nGc6b );
and \U$5778 ( \6493 , \5588_nGcfd , \4937 );
nor \U$5779 ( \6494 , \6491 , \6492 , \6493 );
and \U$5780 ( \6495 , \6487 , \6494 );
and \U$5781 ( \6496 , \6479 , \6486 );
or \U$5782 ( \6497 , \6495 , \6496 );
nand \U$5783 ( \6498 , \6163_nGb55 , \4618 );
or \U$5784 ( \6499 , \4580 , \5968_nGbd0 );
nand \U$5785 ( \6500 , \6499 , \4650 );
and \U$5786 ( \6501 , \6498 , \6500 );
and \U$5787 ( \6502 , \4653 , \5968_nGbd0 );
and \U$5788 ( \6503 , \6163_nGb55 , \4621 );
nor \U$5789 ( \6504 , \6501 , \6502 , \6503 );
and \U$5790 ( \6505 , \4505 , RIb55af80_571);
and \U$5791 ( \6506 , \695 , RIb55b430_581);
and \U$5792 ( \6507 , RIb55b4a8_582, \719 );
nor \U$5793 ( \6508 , \6506 , \6507 );
and \U$5794 ( \6509 , \724 , RIb55b160_575);
and \U$5795 ( \6510 , RIb55b1d8_576, \726 );
nor \U$5796 ( \6511 , \6509 , \6510 );
and \U$5797 ( \6512 , \710 , RIb55b610_585);
and \U$5798 ( \6513 , RIb55b250_577, \690 );
nor \U$5799 ( \6514 , \6512 , \6513 );
and \U$5800 ( \6515 , \716 , RIb55b520_583);
and \U$5801 ( \6516 , RIb55b598_584, \713 );
nor \U$5802 ( \6517 , \6515 , \6516 );
nand \U$5803 ( \6518 , \6508 , \6511 , \6514 , \6517 );
nor \U$5804 ( \6519 , \6505 , \6518 );
and \U$5805 ( \6520 , \703 , RIb55b340_579);
and \U$5806 ( \6521 , RIb55b3b8_580, \698 );
nor \U$5807 ( \6522 , \6520 , \6521 );
and \U$5808 ( \6523 , \740 , RIb55b0e8_574);
and \U$5809 ( \6524 , RIb55aff8_572, \734 );
nor \U$5810 ( \6525 , \6523 , \6524 );
and \U$5811 ( \6526 , \738 , RIb55b070_573);
and \U$5812 ( \6527 , RIb55b2c8_578, \705 );
nor \U$5813 ( \6528 , \6526 , \6527 );
nand \U$5814 ( \6529 , \6519 , \6522 , \6525 , \6528 );
_DC g97a ( \6530_nG97a , \6529 , \4513 );
nand \U$5815 ( \6531 , \6530_nG97a , \4485 );
xor \U$5816 ( \6532 , \6504 , \6531 );
and \U$5817 ( \6533 , \6443_nGa88 , \4559 );
or \U$5818 ( \6534 , \4527 , \6443_nGa88 );
nand \U$5819 ( \6535 , \6534 , \4562 );
nand \U$5820 ( \6536 , \6279_nGadc , \4557 );
and \U$5821 ( \6537 , \6535 , \6536 );
and \U$5822 ( \6538 , \6279_nGadc , \4566 );
nor \U$5823 ( \6539 , \6533 , \6537 , \6538 );
and \U$5824 ( \6540 , \6532 , \6539 );
and \U$5825 ( \6541 , \6504 , \6531 );
or \U$5826 ( \6542 , \6540 , \6541 );
nand \U$5827 ( \6543 , \6497 , \6542 );
or \U$5828 ( \6544 , \5813 , \6324 );
or \U$5829 ( \6545 , \4800_nG140b , \5491 );
or \U$5830 ( \6546 , \4903_nG1319 , \5490 );
nand \U$5831 ( \6547 , \6544 , \6545 , \6546 );
not \U$5832 ( \6548 , \5065_nG112f );
or \U$5833 ( \6549 , \5392 , \6548 );
not \U$5834 ( \6550 , \4876_nG1212 );
or \U$5835 ( \6551 , \6550 , \5981 );
or \U$5836 ( \6552 , \5389 , \6548 );
or \U$5837 ( \6553 , \5259 , \4876_nG1212 );
nand \U$5838 ( \6554 , \6553 , \5478 );
nand \U$5839 ( \6555 , \6552 , \6554 );
nand \U$5840 ( \6556 , \6549 , \6551 , \6555 );
and \U$5841 ( \6557 , \6547 , \6556 );
and \U$5842 ( \6558 , \6543 , \6557 );
nor \U$5843 ( \6559 , \6542 , \6497 );
nor \U$5844 ( \6560 , \6558 , \6559 );
and \U$5845 ( \6561 , \6472 , \6560 );
and \U$5846 ( \6562 , \6466 , \6471 );
or \U$5847 ( \6563 , \6561 , \6562 );
and \U$5848 ( \6564 , \6457 , \6563 );
and \U$5849 ( \6565 , \6454 , \6456 );
or \U$5850 ( \6566 , \6564 , \6565 );
nor \U$5851 ( \6567 , \6409 , \6566 );
xor \U$5852 ( \6568 , \6407 , \6567 );
and \U$5853 ( \6569 , \6409 , \6566 );
nor \U$5854 ( \6570 , \6569 , \6567 );
xor \U$5855 ( \6571 , \6454 , \6456 );
xor \U$5856 ( \6572 , \6571 , \6563 );
xor \U$5857 ( \6573 , \6190 , \6192 );
xor \U$5858 ( \6574 , \6573 , \6194 );
xor \U$5859 ( \6575 , \6366 , \6379 );
xor \U$5860 ( \6576 , \6574 , \6575 );
nor \U$5861 ( \6577 , \6572 , \6576 );
xor \U$5862 ( \6578 , \6570 , \6577 );
and \U$5863 ( \6579 , \6572 , \6576 );
nor \U$5864 ( \6580 , \6579 , \6577 );
nand \U$5865 ( \6581 , \5927_nGc6b , \4805 );
or \U$5866 ( \6582 , \4696 , \5968_nGbd0 );
nand \U$5867 ( \6583 , \6582 , \4811 );
and \U$5868 ( \6584 , \6581 , \6583 );
and \U$5869 ( \6585 , \4807 , \5968_nGbd0 );
and \U$5870 ( \6586 , \5927_nGc6b , \4937 );
nor \U$5871 ( \6587 , \6584 , \6585 , \6586 );
and \U$5872 ( \6588 , \5547_nGdc3 , \5071 );
or \U$5873 ( \6589 , \4928 , \5547_nGdc3 );
nand \U$5874 ( \6590 , \6589 , \5074 );
nand \U$5875 ( \6591 , \5588_nGcfd , \4925 );
and \U$5876 ( \6592 , \6590 , \6591 );
and \U$5877 ( \6593 , \5588_nGcfd , \4930 );
nor \U$5878 ( \6594 , \6588 , \6592 , \6593 );
xor \U$5879 ( \6595 , \6587 , \6594 );
nand \U$5880 ( \6596 , \6279_nGadc , \4618 );
or \U$5881 ( \6597 , \4580 , \6163_nGb55 );
nand \U$5882 ( \6598 , \6597 , \4650 );
and \U$5883 ( \6599 , \6596 , \6598 );
and \U$5884 ( \6600 , \4653 , \6163_nGb55 );
and \U$5885 ( \6601 , \6279_nGadc , \4621 );
nor \U$5886 ( \6602 , \6599 , \6600 , \6601 );
and \U$5887 ( \6603 , \6595 , \6602 );
and \U$5888 ( \6604 , \6587 , \6594 );
or \U$5889 ( \6605 , \6603 , \6604 );
nand \U$5890 ( \6606 , \5311_nG1029 , \5388 );
or \U$5891 ( \6607 , \5259 , \5065_nG112f );
nand \U$5892 ( \6608 , \6607 , \5478 );
and \U$5893 ( \6609 , \6606 , \6608 );
and \U$5894 ( \6610 , \5481 , \5065_nG112f );
and \U$5895 ( \6611 , \5311_nG1029 , \5391 );
nor \U$5896 ( \6612 , \6609 , \6610 , \6611 );
not \U$5897 ( \6613 , \4903_nG1319 );
and \U$5898 ( \6614 , \6613 , \5810 );
and \U$5899 ( \6615 , \5489 , \6550 );
and \U$5900 ( \6616 , \4903_nG1319 , \5814 );
nor \U$5901 ( \6617 , \6614 , \6615 , \6616 );
xor \U$5902 ( \6618 , \6612 , \6617 );
nand \U$5903 ( \6619 , \5520_nGe7a , \5140 );
or \U$5904 ( \6620 , \5093 , \5371_nGf4a );
nand \U$5905 ( \6621 , \6620 , \5248 );
and \U$5906 ( \6622 , \6619 , \6621 );
and \U$5907 ( \6623 , \5243 , \5371_nGf4a );
and \U$5908 ( \6624 , \5520_nGe7a , \5143 );
nor \U$5909 ( \6625 , \6622 , \6623 , \6624 );
and \U$5910 ( \6626 , \6618 , \6625 );
and \U$5911 ( \6627 , \6612 , \6617 );
or \U$5912 ( \6628 , \6626 , \6627 );
xor \U$5913 ( \6629 , \6605 , \6628 );
xor \U$5914 ( \6630 , \6504 , \6531 );
xor \U$5915 ( \6631 , \6630 , \6539 );
and \U$5916 ( \6632 , \6629 , \6631 );
and \U$5917 ( \6633 , \6605 , \6628 );
or \U$5918 ( \6634 , \6632 , \6633 );
xor \U$5919 ( \6635 , \6459 , \6461 );
xor \U$5920 ( \6636 , \6635 , \6463 );
nand \U$5921 ( \6637 , \6634 , \6636 );
xor \U$5922 ( \6638 , \6547 , \6556 );
not \U$5923 ( \6639 , \6638 );
xor \U$5924 ( \6640 , \6479 , \6486 );
xor \U$5925 ( \6641 , \6640 , \6494 );
nor \U$5926 ( \6642 , \6639 , \6641 );
and \U$5927 ( \6643 , \6637 , \6642 );
nor \U$5928 ( \6644 , \6636 , \6634 );
nor \U$5929 ( \6645 , \6643 , \6644 );
not \U$5930 ( \6646 , \6414 );
not \U$5931 ( \6647 , \6453 );
and \U$5932 ( \6648 , \6646 , \6647 );
and \U$5933 ( \6649 , \6414 , \6453 );
nor \U$5934 ( \6650 , \6648 , \6649 );
xor \U$5935 ( \6651 , \6645 , \6650 );
xor \U$5936 ( \6652 , \6466 , \6471 );
xor \U$5937 ( \6653 , \6652 , \6560 );
and \U$5938 ( \6654 , \6651 , \6653 );
and \U$5939 ( \6655 , \6645 , \6650 );
or \U$5940 ( \6656 , \6654 , \6655 );
not \U$5941 ( \6657 , \6656 );
xor \U$5942 ( \6658 , \6580 , \6657 );
xor \U$5943 ( \6659 , \6645 , \6650 );
xor \U$5944 ( \6660 , \6659 , \6653 );
not \U$5945 ( \6661 , \6660 );
not \U$5946 ( \6662 , \6642 );
not \U$5947 ( \6663 , \6644 );
nand \U$5948 ( \6664 , \6663 , \6637 );
not \U$5949 ( \6665 , \6664 );
or \U$5950 ( \6666 , \6662 , \6665 );
or \U$5951 ( \6667 , \6664 , \6642 );
nand \U$5952 ( \6668 , \6666 , \6667 );
not \U$5953 ( \6669 , \6557 );
not \U$5954 ( \6670 , \6559 );
nand \U$5955 ( \6671 , \6670 , \6543 );
not \U$5956 ( \6672 , \6671 );
or \U$5957 ( \6673 , \6669 , \6672 );
or \U$5958 ( \6674 , \6671 , \6557 );
nand \U$5959 ( \6675 , \6673 , \6674 );
nor \U$5960 ( \6676 , \6668 , \6675 );
nand \U$5961 ( \6677 , \5371_nGf4a , \5388 );
or \U$5962 ( \6678 , \5259 , \5311_nG1029 );
nand \U$5963 ( \6679 , \6678 , \5478 );
and \U$5964 ( \6680 , \6677 , \6679 );
and \U$5965 ( \6681 , \5481 , \5311_nG1029 );
and \U$5966 ( \6682 , \5371_nGf4a , \5391 );
nor \U$5967 ( \6683 , \6680 , \6681 , \6682 );
and \U$5968 ( \6684 , \6550 , \5810 );
and \U$5969 ( \6685 , \5489 , \6548 );
and \U$5970 ( \6686 , \4876_nG1212 , \5814 );
nor \U$5971 ( \6687 , \6684 , \6685 , \6686 );
xor \U$5972 ( \6688 , \6683 , \6687 );
and \U$5973 ( \6689 , \6688 , \4527 );
and \U$5974 ( \6690 , \6683 , \6687 );
or \U$5975 ( \6691 , \6689 , \6690 );
and \U$5976 ( \6692 , \5588_nGcfd , \5071 );
or \U$5977 ( \6693 , \4928 , \5588_nGcfd );
nand \U$5978 ( \6694 , \6693 , \5074 );
nand \U$5979 ( \6695 , \5927_nGc6b , \4925 );
and \U$5980 ( \6696 , \6694 , \6695 );
and \U$5981 ( \6697 , \5927_nGc6b , \4930 );
nor \U$5982 ( \6698 , \6692 , \6696 , \6697 );
and \U$5983 ( \6699 , \5547_nGdc3 , \5143 );
or \U$5984 ( \6700 , \5093 , \5520_nGe7a );
nand \U$5985 ( \6701 , \6700 , \5248 );
nand \U$5986 ( \6702 , \5547_nGdc3 , \5140 );
and \U$5987 ( \6703 , \6701 , \6702 );
and \U$5988 ( \6704 , \5520_nGe7a , \5243 );
nor \U$5989 ( \6705 , \6699 , \6703 , \6704 );
xor \U$5990 ( \6706 , \6698 , \6705 );
nand \U$5991 ( \6707 , \5968_nGbd0 , \4805 );
or \U$5992 ( \6708 , \4696 , \6163_nGb55 );
nand \U$5993 ( \6709 , \6708 , \4811 );
and \U$5994 ( \6710 , \6707 , \6709 );
and \U$5995 ( \6711 , \4807 , \6163_nGb55 );
and \U$5996 ( \6712 , \5968_nGbd0 , \4937 );
nor \U$5997 ( \6713 , \6710 , \6711 , \6712 );
and \U$5998 ( \6714 , \6706 , \6713 );
and \U$5999 ( \6715 , \6698 , \6705 );
or \U$6000 ( \6716 , \6714 , \6715 );
xor \U$6001 ( \6717 , \6691 , \6716 );
and \U$6002 ( \6718 , \6530_nG97a , \4559 );
or \U$6003 ( \6719 , \4527 , \6530_nG97a );
nand \U$6004 ( \6720 , \6719 , \4562 );
nand \U$6005 ( \6721 , \6443_nGa88 , \4557 );
and \U$6006 ( \6722 , \6720 , \6721 );
and \U$6007 ( \6723 , \6443_nGa88 , \4566 );
nor \U$6008 ( \6724 , \6718 , \6722 , \6723 );
and \U$6009 ( \6725 , \6717 , \6724 );
and \U$6010 ( \6726 , \6691 , \6716 );
or \U$6011 ( \6727 , \6725 , \6726 );
not \U$6012 ( \6728 , \6641 );
not \U$6013 ( \6729 , \6638 );
and \U$6014 ( \6730 , \6728 , \6729 );
and \U$6015 ( \6731 , \6641 , \6638 );
nor \U$6016 ( \6732 , \6730 , \6731 );
xor \U$6017 ( \6733 , \6727 , \6732 );
xor \U$6018 ( \6734 , \6605 , \6628 );
xor \U$6019 ( \6735 , \6734 , \6631 );
and \U$6020 ( \6736 , \6733 , \6735 );
and \U$6021 ( \6737 , \6727 , \6732 );
or \U$6022 ( \6738 , \6736 , \6737 );
or \U$6023 ( \6739 , \6676 , \6738 );
nand \U$6024 ( \6740 , \6675 , \6668 );
nand \U$6025 ( \6741 , \6739 , \6740 );
xor \U$6026 ( \6742 , \6661 , \6741 );
not \U$6027 ( \6743 , \6738 );
not \U$6028 ( \6744 , \6676 );
nand \U$6029 ( \6745 , \6744 , \6740 );
not \U$6030 ( \6746 , \6745 );
or \U$6031 ( \6747 , \6743 , \6746 );
or \U$6032 ( \6748 , \6745 , \6738 );
nand \U$6033 ( \6749 , \6747 , \6748 );
xor \U$6034 ( \6750 , \6691 , \6716 );
xor \U$6035 ( \6751 , \6750 , \6724 );
xor \U$6036 ( \6752 , \6612 , \6617 );
xor \U$6037 ( \6753 , \6752 , \6625 );
or \U$6038 ( \6754 , \6751 , \6753 );
nand \U$6039 ( \6755 , \6443_nGa88 , \4618 );
or \U$6040 ( \6756 , \4580 , \6279_nGadc );
nand \U$6041 ( \6757 , \6756 , \4650 );
and \U$6042 ( \6758 , \6755 , \6757 );
and \U$6043 ( \6759 , \4653 , \6279_nGadc );
and \U$6044 ( \6760 , \6443_nGa88 , \4621 );
nor \U$6045 ( \6761 , \6758 , \6759 , \6760 );
nand \U$6046 ( \6762 , \5520_nGe7a , \5388 );
or \U$6047 ( \6763 , \5259 , \5371_nGf4a );
nand \U$6048 ( \6764 , \6763 , \5478 );
and \U$6049 ( \6765 , \6762 , \6764 );
and \U$6050 ( \6766 , \5481 , \5371_nGf4a );
and \U$6051 ( \6767 , \5520_nGe7a , \5391 );
nor \U$6052 ( \6768 , \6765 , \6766 , \6767 );
and \U$6053 ( \6769 , \6548 , \5810 );
not \U$6054 ( \6770 , \5311_nG1029 );
and \U$6055 ( \6771 , \5489 , \6770 );
and \U$6056 ( \6772 , \5065_nG112f , \5814 );
nor \U$6057 ( \6773 , \6769 , \6771 , \6772 );
xor \U$6058 ( \6774 , \6768 , \6773 );
nand \U$6059 ( \6775 , \5588_nGcfd , \5140 );
or \U$6060 ( \6776 , \5093 , \5547_nGdc3 );
nand \U$6061 ( \6777 , \6776 , \5248 );
and \U$6062 ( \6778 , \6775 , \6777 );
and \U$6063 ( \6779 , \5243 , \5547_nGdc3 );
and \U$6064 ( \6780 , \5588_nGcfd , \5143 );
nor \U$6065 ( \6781 , \6778 , \6779 , \6780 );
and \U$6066 ( \6782 , \6774 , \6781 );
and \U$6067 ( \6783 , \6768 , \6773 );
or \U$6068 ( \6784 , \6782 , \6783 );
xor \U$6069 ( \6785 , \6761 , \6784 );
nand \U$6070 ( \6786 , \6163_nGb55 , \4805 );
or \U$6071 ( \6787 , \4696 , \6279_nGadc );
nand \U$6072 ( \6788 , \6787 , \4811 );
and \U$6073 ( \6789 , \6786 , \6788 );
and \U$6074 ( \6790 , \4807 , \6279_nGadc );
and \U$6075 ( \6791 , \6163_nGb55 , \4937 );
nor \U$6076 ( \6792 , \6789 , \6790 , \6791 );
and \U$6077 ( \6793 , \5927_nGc6b , \5071 );
or \U$6078 ( \6794 , \4928 , \5927_nGc6b );
nand \U$6079 ( \6795 , \6794 , \5074 );
nand \U$6080 ( \6796 , \5968_nGbd0 , \4925 );
and \U$6081 ( \6797 , \6795 , \6796 );
and \U$6082 ( \6798 , \5968_nGbd0 , \4930 );
nor \U$6083 ( \6799 , \6793 , \6797 , \6798 );
xor \U$6084 ( \6800 , \6792 , \6799 );
nand \U$6085 ( \6801 , \6530_nG97a , \4618 );
or \U$6086 ( \6802 , \4580 , \6443_nGa88 );
nand \U$6087 ( \6803 , \6802 , \4650 );
and \U$6088 ( \6804 , \6801 , \6803 );
and \U$6089 ( \6805 , \4653 , \6443_nGa88 );
and \U$6090 ( \6806 , \6530_nG97a , \4621 );
nor \U$6091 ( \6807 , \6804 , \6805 , \6806 );
and \U$6092 ( \6808 , \6800 , \6807 );
and \U$6093 ( \6809 , \6792 , \6799 );
or \U$6094 ( \6810 , \6808 , \6809 );
and \U$6095 ( \6811 , \6785 , \6810 );
and \U$6096 ( \6812 , \6761 , \6784 );
or \U$6097 ( \6813 , \6811 , \6812 );
xor \U$6098 ( \6814 , \6587 , \6594 );
xor \U$6099 ( \6815 , \6814 , \6602 );
xor \U$6100 ( \6816 , \6813 , \6815 );
xor \U$6101 ( \6817 , \6698 , \6705 );
xor \U$6102 ( \6818 , \6817 , \6713 );
xor \U$6103 ( \6819 , \6683 , \6687 );
xor \U$6104 ( \6820 , \6819 , \4527 );
and \U$6105 ( \6821 , \6818 , \6820 );
and \U$6106 ( \6822 , \4566 , \6530_nG97a );
nand \U$6107 ( \6823 , \6530_nG97a , \4557 );
and \U$6108 ( \6824 , \6823 , \4526 );
nor \U$6109 ( \6825 , \6822 , \6824 );
xor \U$6110 ( \6826 , \6683 , \6687 );
xor \U$6111 ( \6827 , \6826 , \4527 );
and \U$6112 ( \6828 , \6825 , \6827 );
and \U$6113 ( \6829 , \6818 , \6825 );
or \U$6114 ( \6830 , \6821 , \6828 , \6829 );
and \U$6115 ( \6831 , \6816 , \6830 );
and \U$6116 ( \6832 , \6813 , \6815 );
or \U$6117 ( \6833 , \6831 , \6832 );
xor \U$6118 ( \6834 , \6754 , \6833 );
xor \U$6119 ( \6835 , \6727 , \6732 );
xor \U$6120 ( \6836 , \6835 , \6735 );
and \U$6121 ( \6837 , \6834 , \6836 );
and \U$6122 ( \6838 , \6754 , \6833 );
or \U$6123 ( \6839 , \6837 , \6838 );
xor \U$6124 ( \6840 , \6749 , \6839 );
and \U$6125 ( \6841 , \5968_nGbd0 , \5071 );
or \U$6126 ( \6842 , \4928 , \5968_nGbd0 );
nand \U$6127 ( \6843 , \6842 , \5074 );
nand \U$6128 ( \6844 , \6163_nGb55 , \4925 );
and \U$6129 ( \6845 , \6843 , \6844 );
and \U$6130 ( \6846 , \6163_nGb55 , \4930 );
nor \U$6131 ( \6847 , \6841 , \6845 , \6846 );
and \U$6132 ( \6848 , \5927_nGc6b , \5143 );
or \U$6133 ( \6849 , \5093 , \5588_nGcfd );
nand \U$6134 ( \6850 , \6849 , \5248 );
nand \U$6135 ( \6851 , \5927_nGc6b , \5140 );
and \U$6136 ( \6852 , \6850 , \6851 );
and \U$6137 ( \6853 , \5588_nGcfd , \5243 );
nor \U$6138 ( \6854 , \6848 , \6852 , \6853 );
xor \U$6139 ( \6855 , \6847 , \6854 );
nand \U$6140 ( \6856 , \6279_nGadc , \4805 );
or \U$6141 ( \6857 , \4696 , \6443_nGa88 );
nand \U$6142 ( \6858 , \6857 , \4811 );
and \U$6143 ( \6859 , \6856 , \6858 );
and \U$6144 ( \6860 , \4807 , \6443_nGa88 );
and \U$6145 ( \6861 , \6279_nGadc , \4937 );
nor \U$6146 ( \6862 , \6859 , \6860 , \6861 );
and \U$6147 ( \6863 , \6855 , \6862 );
and \U$6148 ( \6864 , \6847 , \6854 );
or \U$6149 ( \6865 , \6863 , \6864 );
nand \U$6150 ( \6866 , \5547_nGdc3 , \5388 );
or \U$6151 ( \6867 , \5259 , \5520_nGe7a );
nand \U$6152 ( \6868 , \6867 , \5478 );
and \U$6153 ( \6869 , \6866 , \6868 );
and \U$6154 ( \6870 , \5481 , \5520_nGe7a );
and \U$6155 ( \6871 , \5547_nGdc3 , \5391 );
nor \U$6156 ( \6872 , \6869 , \6870 , \6871 );
and \U$6157 ( \6873 , \6770 , \5810 );
not \U$6158 ( \6874 , \5371_nGf4a );
and \U$6159 ( \6875 , \5489 , \6874 );
and \U$6160 ( \6876 , \5311_nG1029 , \5814 );
nor \U$6161 ( \6877 , \6873 , \6875 , \6876 );
xor \U$6162 ( \6878 , \6872 , \6877 );
and \U$6163 ( \6879 , \6878 , \4580 );
and \U$6164 ( \6880 , \6872 , \6877 );
or \U$6165 ( \6881 , \6879 , \6880 );
xor \U$6166 ( \6882 , \6865 , \6881 );
xor \U$6167 ( \6883 , \6792 , \6799 );
xor \U$6168 ( \6884 , \6883 , \6807 );
and \U$6169 ( \6885 , \6882 , \6884 );
and \U$6170 ( \6886 , \6865 , \6881 );
or \U$6171 ( \6887 , \6885 , \6886 );
xor \U$6172 ( \6888 , \6761 , \6784 );
xor \U$6173 ( \6889 , \6888 , \6810 );
xor \U$6174 ( \6890 , \6887 , \6889 );
xor \U$6175 ( \6891 , \6683 , \6687 );
xor \U$6176 ( \6892 , \6891 , \4527 );
xor \U$6177 ( \6893 , \6818 , \6825 );
xor \U$6178 ( \6894 , \6892 , \6893 );
and \U$6179 ( \6895 , \6890 , \6894 );
and \U$6180 ( \6896 , \6887 , \6889 );
or \U$6181 ( \6897 , \6895 , \6896 );
xor \U$6182 ( \6898 , \6813 , \6815 );
xor \U$6183 ( \6899 , \6898 , \6830 );
xor \U$6184 ( \6900 , \6897 , \6899 );
xnor \U$6185 ( \6901 , \6753 , \6751 );
xor \U$6186 ( \6902 , \6900 , \6901 );
not \U$6187 ( \6903 , \6902 );
xor \U$6188 ( \6904 , \6887 , \6889 );
xor \U$6189 ( \6905 , \6904 , \6894 );
nand \U$6190 ( \6906 , \5588_nGcfd , \5388 );
or \U$6191 ( \6907 , \5259 , \5547_nGdc3 );
nand \U$6192 ( \6908 , \6907 , \5478 );
and \U$6193 ( \6909 , \6906 , \6908 );
and \U$6194 ( \6910 , \5481 , \5547_nGdc3 );
and \U$6195 ( \6911 , \5588_nGcfd , \5391 );
nor \U$6196 ( \6912 , \6909 , \6910 , \6911 );
not \U$6197 ( \6913 , \6912 );
and \U$6198 ( \6914 , \6874 , \5810 );
not \U$6199 ( \6915 , \5520_nGe7a );
and \U$6200 ( \6916 , \5489 , \6915 );
and \U$6201 ( \6917 , \5371_nGf4a , \5814 );
nor \U$6202 ( \6918 , \6914 , \6916 , \6917 );
not \U$6203 ( \6919 , \6918 );
and \U$6204 ( \6920 , \6913 , \6919 );
and \U$6205 ( \6921 , \6912 , \6918 );
nand \U$6206 ( \6922 , \5968_nGbd0 , \5140 );
or \U$6207 ( \6923 , \5093 , \5927_nGc6b );
nand \U$6208 ( \6924 , \6923 , \5248 );
and \U$6209 ( \6925 , \6922 , \6924 );
and \U$6210 ( \6926 , \5243 , \5927_nGc6b );
and \U$6211 ( \6927 , \5968_nGbd0 , \5143 );
nor \U$6212 ( \6928 , \6925 , \6926 , \6927 );
nor \U$6213 ( \6929 , \6921 , \6928 );
nor \U$6214 ( \6930 , \6920 , \6929 );
xor \U$6215 ( \6931 , \6847 , \6854 );
xor \U$6216 ( \6932 , \6931 , \6862 );
and \U$6217 ( \6933 , \6930 , \6932 );
and \U$6218 ( \6934 , \6530_nG97a , \4653 );
not \U$6219 ( \6935 , \6530_nG97a );
and \U$6220 ( \6936 , \6935 , \4620 );
not \U$6221 ( \6937 , \4650 );
nor \U$6222 ( \6938 , \6934 , \6936 , \6937 );
xor \U$6223 ( \6939 , \6847 , \6854 );
xor \U$6224 ( \6940 , \6939 , \6862 );
and \U$6225 ( \6941 , \6938 , \6940 );
and \U$6226 ( \6942 , \6930 , \6938 );
or \U$6227 ( \6943 , \6933 , \6941 , \6942 );
xor \U$6228 ( \6944 , \6768 , \6773 );
xor \U$6229 ( \6945 , \6944 , \6781 );
xor \U$6230 ( \6946 , \6943 , \6945 );
xor \U$6231 ( \6947 , \6865 , \6881 );
xor \U$6232 ( \6948 , \6947 , \6884 );
and \U$6233 ( \6949 , \6946 , \6948 );
and \U$6234 ( \6950 , \6943 , \6945 );
or \U$6235 ( \6951 , \6949 , \6950 );
nor \U$6236 ( \6952 , \6905 , \6951 );
xor \U$6237 ( \6953 , \6903 , \6952 );
and \U$6238 ( \6954 , \6905 , \6951 );
nor \U$6239 ( \6955 , \6954 , \6952 );
xor \U$6240 ( \6956 , \6943 , \6945 );
xor \U$6241 ( \6957 , \6956 , \6948 );
nand \U$6242 ( \6958 , \5927_nGc6b , \5388 );
or \U$6243 ( \6959 , \5259 , \5588_nGcfd );
nand \U$6244 ( \6960 , \6959 , \5478 );
and \U$6245 ( \6961 , \6958 , \6960 );
and \U$6246 ( \6962 , \5481 , \5588_nGcfd );
and \U$6247 ( \6963 , \5927_nGc6b , \5391 );
nor \U$6248 ( \6964 , \6961 , \6962 , \6963 );
and \U$6249 ( \6965 , \6915 , \5810 );
not \U$6250 ( \6966 , \5547_nGdc3 );
and \U$6251 ( \6967 , \5489 , \6966 );
and \U$6252 ( \6968 , \5520_nGe7a , \5814 );
nor \U$6253 ( \6969 , \6965 , \6967 , \6968 );
xor \U$6254 ( \6970 , \6964 , \6969 );
and \U$6255 ( \6971 , \6970 , \4696 );
and \U$6256 ( \6972 , \6964 , \6969 );
or \U$6257 ( \6973 , \6971 , \6972 );
and \U$6258 ( \6974 , \6163_nGb55 , \5071 );
or \U$6259 ( \6975 , \4928 , \6163_nGb55 );
nand \U$6260 ( \6976 , \6975 , \5074 );
nand \U$6261 ( \6977 , \6279_nGadc , \4925 );
and \U$6262 ( \6978 , \6976 , \6977 );
and \U$6263 ( \6979 , \6279_nGadc , \4930 );
nor \U$6264 ( \6980 , \6974 , \6978 , \6979 );
xor \U$6265 ( \6981 , \6973 , \6980 );
and \U$6266 ( \6982 , \6279_nGadc , \5071 );
or \U$6267 ( \6983 , \4928 , \6279_nGadc );
nand \U$6268 ( \6984 , \6983 , \5074 );
nand \U$6269 ( \6985 , \6443_nGa88 , \4925 );
and \U$6270 ( \6986 , \6984 , \6985 );
and \U$6271 ( \6987 , \6443_nGa88 , \4930 );
nor \U$6272 ( \6988 , \6982 , \6986 , \6987 );
and \U$6273 ( \6989 , \6163_nGb55 , \5143 );
or \U$6274 ( \6990 , \5093 , \5968_nGbd0 );
nand \U$6275 ( \6991 , \6990 , \5248 );
nand \U$6276 ( \6992 , \6163_nGb55 , \5140 );
and \U$6277 ( \6993 , \6991 , \6992 );
and \U$6278 ( \6994 , \5968_nGbd0 , \5243 );
nor \U$6279 ( \6995 , \6989 , \6993 , \6994 );
xor \U$6280 ( \6996 , \6988 , \6995 );
and \U$6281 ( \6997 , \4937 , \6530_nG97a );
nand \U$6282 ( \6998 , \6530_nG97a , \4805 );
and \U$6283 ( \6999 , \6998 , \4809 );
nor \U$6284 ( \7000 , \6997 , \6999 );
and \U$6285 ( \7001 , \6996 , \7000 );
and \U$6286 ( \7002 , \6988 , \6995 );
or \U$6287 ( \7003 , \7001 , \7002 );
and \U$6288 ( \7004 , \6981 , \7003 );
and \U$6289 ( \7005 , \6973 , \6980 );
or \U$6290 ( \7006 , \7004 , \7005 );
xor \U$6291 ( \7007 , \6872 , \6877 );
xor \U$6292 ( \7008 , \7007 , \4580 );
nand \U$6293 ( \7009 , \7006 , \7008 );
not \U$6294 ( \7010 , \6912 );
xor \U$6295 ( \7011 , \6918 , \6928 );
not \U$6296 ( \7012 , \7011 );
or \U$6297 ( \7013 , \7010 , \7012 );
or \U$6298 ( \7014 , \7011 , \6912 );
nand \U$6299 ( \7015 , \7013 , \7014 );
not \U$6300 ( \7016 , \6443_nGa88 );
or \U$6301 ( \7017 , \4938 , \7016 );
or \U$6302 ( \7018 , \6935 , \4940 );
or \U$6303 ( \7019 , \4936 , \7016 );
or \U$6304 ( \7020 , \4696 , \6530_nG97a );
nand \U$6305 ( \7021 , \7020 , \4811 );
nand \U$6306 ( \7022 , \7019 , \7021 );
nand \U$6307 ( \7023 , \7017 , \7018 , \7022 );
and \U$6308 ( \7024 , \7015 , \7023 );
and \U$6309 ( \7025 , \7009 , \7024 );
nor \U$6310 ( \7026 , \7006 , \7008 );
nor \U$6311 ( \7027 , \7025 , \7026 );
nor \U$6312 ( \7028 , \6957 , \7027 );
xor \U$6313 ( \7029 , \6955 , \7028 );
not \U$6314 ( \7030 , \7024 );
not \U$6315 ( \7031 , \7026 );
nand \U$6316 ( \7032 , \7031 , \7009 );
not \U$6317 ( \7033 , \7032 );
or \U$6318 ( \7034 , \7030 , \7033 );
or \U$6319 ( \7035 , \7032 , \7024 );
nand \U$6320 ( \7036 , \7034 , \7035 );
xor \U$6321 ( \7037 , \6847 , \6854 );
xor \U$6322 ( \7038 , \7037 , \6862 );
xor \U$6323 ( \7039 , \6930 , \6938 );
xor \U$6324 ( \7040 , \7038 , \7039 );
not \U$6325 ( \7041 , \7040 );
xor \U$6326 ( \7042 , \7036 , \7041 );
xor \U$6327 ( \7043 , \6973 , \6980 );
xor \U$6328 ( \7044 , \7043 , \7003 );
nand \U$6329 ( \7045 , \5968_nGbd0 , \5388 );
or \U$6330 ( \7046 , \5259 , \5927_nGc6b );
nand \U$6331 ( \7047 , \7046 , \5478 );
and \U$6332 ( \7048 , \7045 , \7047 );
and \U$6333 ( \7049 , \5481 , \5927_nGc6b );
and \U$6334 ( \7050 , \5968_nGbd0 , \5391 );
nor \U$6335 ( \7051 , \7048 , \7049 , \7050 );
and \U$6336 ( \7052 , \6966 , \5810 );
not \U$6337 ( \7053 , \5588_nGcfd );
and \U$6338 ( \7054 , \5489 , \7053 );
and \U$6339 ( \7055 , \5547_nGdc3 , \5814 );
nor \U$6340 ( \7056 , \7052 , \7054 , \7055 );
xor \U$6341 ( \7057 , \7051 , \7056 );
nand \U$6342 ( \7058 , \6279_nGadc , \5140 );
or \U$6343 ( \7059 , \5093 , \6163_nGb55 );
nand \U$6344 ( \7060 , \7059 , \5248 );
and \U$6345 ( \7061 , \7058 , \7060 );
and \U$6346 ( \7062 , \5243 , \6163_nGb55 );
and \U$6347 ( \7063 , \6279_nGadc , \5143 );
nor \U$6348 ( \7064 , \7061 , \7062 , \7063 );
and \U$6349 ( \7065 , \7057 , \7064 );
and \U$6350 ( \7066 , \7051 , \7056 );
or \U$6351 ( \7067 , \7065 , \7066 );
xor \U$6352 ( \7068 , \6964 , \6969 );
xor \U$6353 ( \7069 , \7068 , \4696 );
and \U$6354 ( \7070 , \7067 , \7069 );
xor \U$6355 ( \7071 , \6988 , \6995 );
xor \U$6356 ( \7072 , \7071 , \7000 );
xor \U$6357 ( \7073 , \6964 , \6969 );
xor \U$6358 ( \7074 , \7073 , \4696 );
and \U$6359 ( \7075 , \7072 , \7074 );
and \U$6360 ( \7076 , \7067 , \7072 );
or \U$6361 ( \7077 , \7070 , \7075 , \7076 );
nor \U$6362 ( \7078 , \7044 , \7077 );
xor \U$6363 ( \7079 , \7015 , \7023 );
or \U$6364 ( \7080 , \7078 , \7079 );
nand \U$6365 ( \7081 , \7077 , \7044 );
nand \U$6366 ( \7082 , \7080 , \7081 );
not \U$6367 ( \7083 , \7082 );
xor \U$6368 ( \7084 , \7042 , \7083 );
not \U$6369 ( \7085 , \7081 );
nor \U$6370 ( \7086 , \7085 , \7078 );
not \U$6371 ( \7087 , \7086 );
not \U$6372 ( \7088 , \7079 );
and \U$6373 ( \7089 , \7087 , \7088 );
and \U$6374 ( \7090 , \7086 , \7079 );
nor \U$6375 ( \7091 , \7089 , \7090 );
xor \U$6376 ( \7092 , \6964 , \6969 );
xor \U$6377 ( \7093 , \7092 , \4696 );
xor \U$6378 ( \7094 , \7067 , \7072 );
xor \U$6379 ( \7095 , \7093 , \7094 );
nand \U$6380 ( \7096 , \6443_nGa88 , \5140 );
or \U$6381 ( \7097 , \5093 , \6279_nGadc );
nand \U$6382 ( \7098 , \7097 , \5248 );
and \U$6383 ( \7099 , \7096 , \7098 );
and \U$6384 ( \7100 , \5243 , \6279_nGadc );
and \U$6385 ( \7101 , \6443_nGa88 , \5143 );
nor \U$6386 ( \7102 , \7099 , \7100 , \7101 );
not \U$6387 ( \7103 , \7102 );
or \U$6388 ( \7104 , \5149 , \6935 );
or \U$6389 ( \7105 , \6530_nG97a , \4928 );
nand \U$6390 ( \7106 , \7104 , \7105 , \5074 );
nand \U$6391 ( \7107 , \7103 , \7106 );
nand \U$6392 ( \7108 , \6163_nGb55 , \5388 );
or \U$6393 ( \7109 , \5259 , \5968_nGbd0 );
nand \U$6394 ( \7110 , \7109 , \5478 );
and \U$6395 ( \7111 , \7108 , \7110 );
and \U$6396 ( \7112 , \5481 , \5968_nGbd0 );
and \U$6397 ( \7113 , \6163_nGb55 , \5391 );
nor \U$6398 ( \7114 , \7111 , \7112 , \7113 );
and \U$6399 ( \7115 , \7053 , \5810 );
not \U$6400 ( \7116 , \5927_nGc6b );
and \U$6401 ( \7117 , \5489 , \7116 );
and \U$6402 ( \7118 , \5588_nGcfd , \5814 );
nor \U$6403 ( \7119 , \7115 , \7117 , \7118 );
xor \U$6404 ( \7120 , \7114 , \7119 );
and \U$6405 ( \7121 , \7120 , \4928 );
and \U$6406 ( \7122 , \7114 , \7119 );
or \U$6407 ( \7123 , \7121 , \7122 );
xor \U$6408 ( \7124 , \7107 , \7123 );
and \U$6409 ( \7125 , \6443_nGa88 , \5071 );
or \U$6410 ( \7126 , \4928 , \6443_nGa88 );
nand \U$6411 ( \7127 , \7126 , \5074 );
nand \U$6412 ( \7128 , \6530_nG97a , \4925 );
and \U$6413 ( \7129 , \7127 , \7128 );
and \U$6414 ( \7130 , \6530_nG97a , \4930 );
nor \U$6415 ( \7131 , \7125 , \7129 , \7130 );
and \U$6416 ( \7132 , \7124 , \7131 );
and \U$6417 ( \7133 , \7107 , \7123 );
or \U$6418 ( \7134 , \7132 , \7133 );
nor \U$6419 ( \7135 , \7095 , \7134 );
xor \U$6420 ( \7136 , \7091 , \7135 );
not \U$6421 ( \7137 , \7102 );
not \U$6422 ( \7138 , \7106 );
or \U$6423 ( \7139 , \7137 , \7138 );
or \U$6424 ( \7140 , \7106 , \7102 );
nand \U$6425 ( \7141 , \7139 , \7140 );
not \U$6426 ( \7142 , \7141 );
xor \U$6427 ( \7143 , \7114 , \7119 );
xor \U$6428 ( \7144 , \7143 , \4928 );
nand \U$6429 ( \7145 , \6279_nGadc , \5388 );
or \U$6430 ( \7146 , \5259 , \6163_nGb55 );
nand \U$6431 ( \7147 , \7146 , \5478 );
and \U$6432 ( \7148 , \7145 , \7147 );
and \U$6433 ( \7149 , \5481 , \6163_nGb55 );
and \U$6434 ( \7150 , \6279_nGadc , \5391 );
nor \U$6435 ( \7151 , \7148 , \7149 , \7150 );
and \U$6436 ( \7152 , \7116 , \5810 );
not \U$6437 ( \7153 , \5968_nGbd0 );
and \U$6438 ( \7154 , \5489 , \7153 );
and \U$6439 ( \7155 , \5927_nGc6b , \5814 );
nor \U$6440 ( \7156 , \7152 , \7154 , \7155 );
xor \U$6441 ( \7157 , \7151 , \7156 );
nand \U$6442 ( \7158 , \6530_nG97a , \5140 );
or \U$6443 ( \7159 , \5093 , \6443_nGa88 );
nand \U$6444 ( \7160 , \7159 , \5248 );
and \U$6445 ( \7161 , \7158 , \7160 );
and \U$6446 ( \7162 , \5243 , \6443_nGa88 );
and \U$6447 ( \7163 , \6530_nG97a , \5143 );
nor \U$6448 ( \7164 , \7161 , \7162 , \7163 );
and \U$6449 ( \7165 , \7157 , \7164 );
and \U$6450 ( \7166 , \7151 , \7156 );
or \U$6451 ( \7167 , \7165 , \7166 );
nand \U$6452 ( \7168 , \7144 , \7167 );
not \U$6453 ( \7169 , \7168 );
nor \U$6454 ( \7170 , \7167 , \7144 );
nor \U$6455 ( \7171 , \7169 , \7170 );
not \U$6456 ( \7172 , \7171 );
and \U$6457 ( \7173 , \7142 , \7172 );
and \U$6458 ( \7174 , \7141 , \7171 );
nor \U$6459 ( \7175 , \7173 , \7174 );
xor \U$6460 ( \7176 , \7151 , \7156 );
xor \U$6461 ( \7177 , \7176 , \7164 );
and \U$6462 ( \7178 , \7153 , \5810 );
not \U$6463 ( \7179 , \6163_nGb55 );
and \U$6464 ( \7180 , \5489 , \7179 );
and \U$6465 ( \7181 , \5968_nGbd0 , \5814 );
nor \U$6466 ( \7182 , \7178 , \7180 , \7181 );
xor \U$6467 ( \7183 , \5093 , \7182 );
nand \U$6468 ( \7184 , \6443_nGa88 , \5388 );
or \U$6469 ( \7185 , \5259 , \6279_nGadc );
nand \U$6470 ( \7186 , \7185 , \5478 );
and \U$6471 ( \7187 , \7184 , \7186 );
and \U$6472 ( \7188 , \5481 , \6279_nGadc );
and \U$6473 ( \7189 , \6443_nGa88 , \5391 );
nor \U$6474 ( \7190 , \7187 , \7188 , \7189 );
and \U$6475 ( \7191 , \7183 , \7190 );
and \U$6476 ( \7192 , \5093 , \7182 );
or \U$6477 ( \7193 , \7191 , \7192 );
nor \U$6478 ( \7194 , \7177 , \7193 );
xor \U$6479 ( \7195 , \7175 , \7194 );
not \U$6480 ( \7196 , \6279_nGadc );
or \U$6481 ( \7197 , \5813 , \7196 );
or \U$6482 ( \7198 , \6279_nGadc , \5491 );
or \U$6483 ( \7199 , \6443_nGa88 , \5490 );
nand \U$6484 ( \7200 , \7197 , \7198 , \7199 );
xor \U$6485 ( \7201 , \7200 , \5390 );
and \U$6486 ( \7202 , \7016 , \5810 );
and \U$6487 ( \7203 , \5489 , \6935 );
and \U$6488 ( \7204 , \6443_nGa88 , \5814 );
nor \U$6489 ( \7205 , \7202 , \7203 , \7204 );
nand \U$6490 ( \7206 , \6530_nG97a , \5490 );
nand \U$6491 ( \7207 , \5254 , \7206 );
nor \U$6492 ( \7208 , \7205 , \7207 );
xor \U$6493 ( \7209 , \7201 , \7208 );
or \U$6494 ( \7210 , \5981 , \6935 );
or \U$6495 ( \7211 , \6530_nG97a , \5259 );
nand \U$6496 ( \7212 , \7210 , \7211 , \5478 );
and \U$6497 ( \7213 , \7209 , \7212 );
and \U$6498 ( \7214 , \7201 , \7208 );
or \U$6499 ( \7215 , \7213 , \7214 );
and \U$6500 ( \7216 , \7200 , \5390 );
xor \U$6501 ( \7217 , \7215 , \7216 );
nand \U$6502 ( \7218 , \6530_nG97a , \5388 );
or \U$6503 ( \7219 , \5259 , \6443_nGa88 );
nand \U$6504 ( \7220 , \7219 , \5478 );
and \U$6505 ( \7221 , \7218 , \7220 );
and \U$6506 ( \7222 , \5481 , \6443_nGa88 );
and \U$6507 ( \7223 , \6530_nG97a , \5391 );
nor \U$6508 ( \7224 , \7221 , \7222 , \7223 );
and \U$6509 ( \7225 , \7179 , \5810 );
and \U$6510 ( \7226 , \5489 , \7196 );
and \U$6511 ( \7227 , \6163_nGb55 , \5814 );
nor \U$6512 ( \7228 , \7225 , \7226 , \7227 );
and \U$6513 ( \7229 , \7224 , \7228 );
nor \U$6514 ( \7230 , \7224 , \7228 );
nor \U$6515 ( \7231 , \7229 , \7230 );
and \U$6516 ( \7232 , \7217 , \7231 );
and \U$6517 ( \7233 , \7215 , \7216 );
or \U$6518 ( \7234 , \7232 , \7233 );
xor \U$6519 ( \7235 , \7234 , \7230 );
and \U$6520 ( \7236 , \6530_nG97a , \5243 );
and \U$6521 ( \7237 , \6935 , \5142 );
not \U$6522 ( \7238 , \5248 );
nor \U$6523 ( \7239 , \7236 , \7237 , \7238 );
xor \U$6524 ( \7240 , \5093 , \7182 );
xor \U$6525 ( \7241 , \7240 , \7190 );
and \U$6526 ( \7242 , \7239 , \7241 );
nor \U$6527 ( \7243 , \7239 , \7241 );
nor \U$6528 ( \7244 , \7242 , \7243 );
and \U$6529 ( \7245 , \7235 , \7244 );
and \U$6530 ( \7246 , \7234 , \7230 );
or \U$6531 ( \7247 , \7245 , \7246 );
xor \U$6532 ( \7248 , \7247 , \7243 );
and \U$6533 ( \7249 , \7177 , \7193 );
nor \U$6534 ( \7250 , \7249 , \7194 );
and \U$6535 ( \7251 , \7248 , \7250 );
and \U$6536 ( \7252 , \7247 , \7243 );
or \U$6537 ( \7253 , \7251 , \7252 );
and \U$6538 ( \7254 , \7195 , \7253 );
and \U$6539 ( \7255 , \7175 , \7194 );
or \U$6540 ( \7256 , \7254 , \7255 );
or \U$6541 ( \7257 , \7141 , \7170 );
nand \U$6542 ( \7258 , \7257 , \7168 );
not \U$6543 ( \7259 , \7258 );
xor \U$6544 ( \7260 , \7256 , \7259 );
xor \U$6545 ( \7261 , \7107 , \7123 );
xor \U$6546 ( \7262 , \7261 , \7131 );
xor \U$6547 ( \7263 , \7051 , \7056 );
xor \U$6548 ( \7264 , \7263 , \7064 );
and \U$6549 ( \7265 , \7262 , \7264 );
nor \U$6550 ( \7266 , \7262 , \7264 );
nor \U$6551 ( \7267 , \7265 , \7266 );
and \U$6552 ( \7268 , \7260 , \7267 );
and \U$6553 ( \7269 , \7256 , \7259 );
or \U$6554 ( \7270 , \7268 , \7269 );
xor \U$6555 ( \7271 , \7270 , \7266 );
and \U$6556 ( \7272 , \7095 , \7134 );
nor \U$6557 ( \7273 , \7272 , \7135 );
and \U$6558 ( \7274 , \7271 , \7273 );
and \U$6559 ( \7275 , \7270 , \7266 );
or \U$6560 ( \7276 , \7274 , \7275 );
and \U$6561 ( \7277 , \7136 , \7276 );
and \U$6562 ( \7278 , \7091 , \7135 );
or \U$6563 ( \7279 , \7277 , \7278 );
and \U$6564 ( \7280 , \7084 , \7279 );
and \U$6565 ( \7281 , \7042 , \7083 );
or \U$6566 ( \7282 , \7280 , \7281 );
and \U$6567 ( \7283 , \7036 , \7041 );
xor \U$6568 ( \7284 , \7282 , \7283 );
and \U$6569 ( \7285 , \6957 , \7027 );
nor \U$6570 ( \7286 , \7285 , \7028 );
and \U$6571 ( \7287 , \7284 , \7286 );
and \U$6572 ( \7288 , \7282 , \7283 );
or \U$6573 ( \7289 , \7287 , \7288 );
and \U$6574 ( \7290 , \7029 , \7289 );
and \U$6575 ( \7291 , \6955 , \7028 );
or \U$6576 ( \7292 , \7290 , \7291 );
and \U$6577 ( \7293 , \6953 , \7292 );
and \U$6578 ( \7294 , \6903 , \6952 );
or \U$6579 ( \7295 , \7293 , \7294 );
xor \U$6580 ( \7296 , \6897 , \6899 );
and \U$6581 ( \7297 , \7296 , \6901 );
and \U$6582 ( \7298 , \6897 , \6899 );
or \U$6583 ( \7299 , \7297 , \7298 );
xor \U$6584 ( \7300 , \6754 , \6833 );
xor \U$6585 ( \7301 , \7300 , \6836 );
nand \U$6586 ( \7302 , \7299 , \7301 );
and \U$6587 ( \7303 , \7295 , \7302 );
nor \U$6588 ( \7304 , \7301 , \7299 );
nor \U$6589 ( \7305 , \7303 , \7304 );
and \U$6590 ( \7306 , \6840 , \7305 );
and \U$6591 ( \7307 , \6749 , \6839 );
or \U$6592 ( \7308 , \7306 , \7307 );
not \U$6593 ( \7309 , \7308 );
and \U$6594 ( \7310 , \6742 , \7309 );
and \U$6595 ( \7311 , \6661 , \6741 );
or \U$6596 ( \7312 , \7310 , \7311 );
and \U$6597 ( \7313 , \6658 , \7312 );
and \U$6598 ( \7314 , \6580 , \6657 );
or \U$6599 ( \7315 , \7313 , \7314 );
and \U$6600 ( \7316 , \6578 , \7315 );
and \U$6601 ( \7317 , \6570 , \6577 );
or \U$6602 ( \7318 , \7316 , \7317 );
and \U$6603 ( \7319 , \6568 , \7318 );
and \U$6604 ( \7320 , \6407 , \6567 );
or \U$6605 ( \7321 , \7319 , \7320 );
and \U$6606 ( \7322 , \6403 , \7321 );
and \U$6607 ( \7323 , \6311 , \6402 );
or \U$6608 ( \7324 , \7322 , \7323 );
and \U$6609 ( \7325 , \6309 , \7324 );
and \U$6610 ( \7326 , \6131 , \6308 );
or \U$6611 ( \7327 , \7325 , \7326 );
and \U$6612 ( \7328 , \6129 , \7327 );
and \U$6613 ( \7329 , \6045 , \6128 );
or \U$6614 ( \7330 , \7328 , \7329 );
not \U$6615 ( \7331 , \5863 );
not \U$6616 ( \7332 , \5772 );
or \U$6617 ( \7333 , \7331 , \7332 );
or \U$6618 ( \7334 , \5772 , \5863 );
nand \U$6619 ( \7335 , \7333 , \7334 );
not \U$6620 ( \7336 , \7335 );
not \U$6621 ( \7337 , \5764 );
and \U$6622 ( \7338 , \7336 , \7337 );
and \U$6623 ( \7339 , \7335 , \5764 );
nor \U$6624 ( \7340 , \7338 , \7339 );
not \U$6625 ( \7341 , \6034 );
not \U$6626 ( \7342 , \6041 );
and \U$6627 ( \7343 , \7341 , \7342 );
nor \U$6628 ( \7344 , \7343 , \6033 );
nand \U$6629 ( \7345 , \7340 , \7344 );
and \U$6630 ( \7346 , \7330 , \7345 );
nor \U$6631 ( \7347 , \7344 , \7340 );
nor \U$6632 ( \7348 , \7346 , \7347 );
nor \U$6633 ( \7349 , \5869 , \7348 );
nor \U$6634 ( \7350 , \5866 , \7349 );
not \U$6635 ( \7351 , \7350 );
and \U$6636 ( \7352 , \5755 , \7351 );
and \U$6637 ( \7353 , \5734 , \5754 );
or \U$6638 ( \7354 , \7352 , \7353 );
and \U$6639 ( \7355 , \5744 , \5750 );
nor \U$6640 ( \7356 , \7355 , \5746 );
not \U$6641 ( \7357 , \5442 );
not \U$6642 ( \7358 , \5340 );
nand \U$6643 ( \7359 , \7358 , \5444 );
not \U$6644 ( \7360 , \7359 );
or \U$6645 ( \7361 , \7357 , \7360 );
or \U$6646 ( \7362 , \7359 , \5442 );
nand \U$6647 ( \7363 , \7361 , \7362 );
nand \U$6648 ( \7364 , \7356 , \7363 );
and \U$6649 ( \7365 , \7354 , \7364 );
nor \U$6650 ( \7366 , \7363 , \7356 );
nor \U$6651 ( \7367 , \7365 , \7366 );
not \U$6652 ( \7368 , \7367 );
and \U$6653 ( \7369 , \5450 , \7368 );
and \U$6654 ( \7370 , \5445 , \5449 );
or \U$6655 ( \7371 , \7369 , \7370 );
and \U$6656 ( \7372 , \5336 , \7371 );
and \U$6657 ( \7373 , \5220 , \5335 );
or \U$6658 ( \7374 , \7372 , \7373 );
not \U$6659 ( \7375 , \5211 );
not \U$6660 ( \7376 , \5216 );
or \U$6661 ( \7377 , \7375 , \7376 );
nand \U$6662 ( \7378 , \7377 , \5212 );
xor \U$6663 ( \7379 , \5112 , \5114 );
xor \U$6664 ( \7380 , \7379 , \5117 );
nand \U$6665 ( \7381 , \7378 , \7380 );
and \U$6666 ( \7382 , \7374 , \7381 );
nor \U$6667 ( \7383 , \7380 , \7378 );
nor \U$6668 ( \7384 , \7382 , \7383 );
xor \U$6669 ( \7385 , \4841 , \4843 );
xor \U$6670 ( \7386 , \7385 , \5007 );
and \U$6671 ( \7387 , \7384 , \7386 );
and \U$6672 ( \7388 , \5120 , \7384 );
or \U$6673 ( \7389 , \5123 , \7387 , \7388 );
and \U$6674 ( \7390 , \5018 , \7389 );
and \U$6675 ( \7391 , \5010 , \5017 );
or \U$6676 ( \7392 , \7390 , \7391 );
not \U$6677 ( \7393 , \7392 );
and \U$6678 ( \7394 , \4836 , \7393 );
and \U$6679 ( \7395 , \4834 , \4835 );
or \U$6680 ( \7396 , \7394 , \7395 );
not \U$6681 ( \7397 , \7396 );
or \U$6682 ( \7398 , \4729 , \7397 );
or \U$6683 ( \7399 , \7396 , \4728 );
nand \U$6684 ( \7400 , \7398 , \7399 );
buf \U$6685 ( \7401 , \4098 );
buf \U$6686 ( \7402 , \750 );
_DC g476 ( \7403_nG476 , \7401 , \7402 );
not \U$6687 ( \7404 , \7403_nG476 );
buf \U$6688 ( \7405 , \745 );
buf \U$6689 ( \7406 , \750 );
_DC g473 ( \7407_nG473 , \7405 , \7406 );
and \U$6690 ( \7408 , \7404 , \7407_nG473 );
nor \U$6691 ( \7409 , \652 , RIb55b778_588);
and \U$6692 ( \7410 , \7409 , RIb54a798_8);
nand \U$6693 ( \7411 , RIb54a720_7, \7410 );
not \U$6694 ( \7412 , \7411 );
nand \U$6695 ( \7413 , \7412 , RIb54a6a8_6);
nor \U$6696 ( \7414 , \7413 , \902 );
nand \U$6697 ( \7415 , RIb54a5b8_4, \7414 );
nor \U$6698 ( \7416 , \7415 , \828 );
nand \U$6699 ( \7417 , RIb54a4c8_2, \7416 );
not \U$6700 ( \7418 , \7417 );
nand \U$6701 ( \7419 , \7418 , RIb54a450_1);
not \U$6702 ( \7420 , \7419 );
not \U$6703 ( \7421 , RIb5517a0_247);
and \U$6704 ( \7422 , \7420 , \7421 );
and \U$6705 ( \7423 , \7419 , RIb5517a0_247);
nor \U$6706 ( \7424 , \7422 , \7423 );
not \U$6707 ( \7425 , \7424 );
buf \U$6708 ( \7426 , \4098 );
buf \U$6709 ( \7427 , \750 );
_DC g2fa ( \7428_nG2fa , \7426 , \7427 );
not \U$6710 ( \7429 , \7428_nG2fa );
and \U$6711 ( \7430 , \7425 , \7429 );
and \U$6712 ( \7431 , \7428_nG2fa , \7424 );
buf \U$6713 ( \7432 , \4128 );
_DC g317 ( \7433_nG317 , \7432 , \7427 );
buf \U$6714 ( \7434 , \4157 );
_DC g334 ( \7435_nG334 , \7434 , \7427 );
not \U$6715 ( \7436 , \7435_nG334 );
or \U$6716 ( \7437 , \7416 , RIb54a4c8_2);
nand \U$6717 ( \7438 , \7437 , \7417 );
not \U$6718 ( \7439 , \7438 );
or \U$6719 ( \7440 , \7436 , \7439 );
buf \U$6720 ( \7441 , \4271 );
_DC g3a6 ( \7442_nG3a6 , \7441 , \7427 );
not \U$6721 ( \7443 , \7442_nG3a6 );
not \U$6722 ( \7444 , \938 );
not \U$6723 ( \7445 , \7411 );
or \U$6724 ( \7446 , \7444 , \7445 );
nand \U$6725 ( \7447 , \7446 , \7413 );
not \U$6726 ( \7448 , \7447 );
or \U$6727 ( \7449 , \7443 , \7448 );
or \U$6728 ( \7450 , \7447 , \7442_nG3a6 );
buf \U$6729 ( \7451 , \4300 );
_DC g3c3 ( \7452_nG3c3 , \7451 , \7427 );
xnor \U$6730 ( \7453 , RIb54a798_8, \7409 );
buf \U$6731 ( \7454 , \4329 );
_DC g3e0 ( \7455_nG3e0 , \7454 , \7427 );
and \U$6732 ( \7456 , \7453 , \7455_nG3e0 );
not \U$6733 ( \7457 , \7453 );
not \U$6734 ( \7458 , \7455_nG3e0 );
and \U$6735 ( \7459 , \7457 , \7458 );
buf \U$6736 ( \7460 , \4387 );
_DC g41a ( \7461_nG41a , \7460 , \7427 );
not \U$6737 ( \7462 , \7461_nG41a );
not \U$6738 ( \7463 , RIb55b778_588);
nand \U$6739 ( \7464 , RIb54a900_11, \7463 );
not \U$6740 ( \7465 , \7464 );
nor \U$6741 ( \7466 , \7463 , RIb54a900_11);
buf \U$6742 ( \7467 , \4416 );
_DC g437 ( \7468_nG437 , \7467 , \7427 );
or \U$6743 ( \7469 , \7465 , \7466 , \7468_nG437 );
buf \U$6744 ( \7470 , \4444 );
_DC g453 ( \7471_nG453 , \7470 , \7427 );
nand \U$6745 ( \7472 , \7469 , \7471_nG453 );
or \U$6746 ( \7473 , \7472 , RIb550378_204);
or \U$6747 ( \7474 , \7465 , \7466 );
nand \U$6748 ( \7475 , \7474 , \7468_nG437 );
nand \U$6749 ( \7476 , \7473 , \7475 );
not \U$6750 ( \7477 , \7476 );
or \U$6751 ( \7478 , \7462 , \7477 );
or \U$6752 ( \7479 , \7476 , \7461_nG41a );
or \U$6753 ( \7480 , RIb54a888_10, \7464 );
nand \U$6754 ( \7481 , RIb54a888_10, \7464 );
nand \U$6755 ( \7482 , \7479 , \7480 , \7481 );
nand \U$6756 ( \7483 , \7478 , \7482 );
buf \U$6757 ( \7484 , \4358 );
_DC g3fd ( \7485_nG3fd , \7484 , \7427 );
and \U$6758 ( \7486 , \7483 , \7485_nG3fd );
and \U$6759 ( \7487 , \651 , \7463 );
nor \U$6760 ( \7488 , \7487 , RIb54a810_9);
or \U$6761 ( \7489 , \7486 , \7409 , \7488 );
or \U$6762 ( \7490 , \7483 , \7485_nG3fd );
nand \U$6763 ( \7491 , \7489 , \7490 );
nor \U$6764 ( \7492 , \7459 , \7491 );
nor \U$6765 ( \7493 , \7456 , \7492 );
not \U$6766 ( \7494 , \7493 );
or \U$6767 ( \7495 , \7452_nG3c3 , \7494 );
not \U$6768 ( \7496 , \7452_nG3c3 );
or \U$6769 ( \7497 , \7493 , \7496 );
or \U$6770 ( \7498 , RIb54a720_7, \7410 );
nand \U$6771 ( \7499 , \7497 , \7498 , \7411 );
nand \U$6772 ( \7500 , \7450 , \7495 , \7499 );
nand \U$6773 ( \7501 , \7449 , \7500 );
buf \U$6774 ( \7502 , \4243 );
_DC g38a ( \7503_nG38a , \7502 , \7427 );
and \U$6775 ( \7504 , \7501 , \7503_nG38a );
and \U$6776 ( \7505 , \7413 , RIb54a630_5);
nor \U$6777 ( \7506 , \7501 , \7503_nG38a );
nor \U$6778 ( \7507 , \7413 , RIb54a630_5);
nor \U$6779 ( \7508 , \7505 , \7506 , \7507 );
nor \U$6780 ( \7509 , \7504 , \7508 );
or \U$6781 ( \7510 , \7414 , RIb54a5b8_4);
nand \U$6782 ( \7511 , \7510 , \7415 );
not \U$6783 ( \7512 , \7511 );
and \U$6784 ( \7513 , \7509 , \7512 );
not \U$6785 ( \7514 , \7509 );
not \U$6786 ( \7515 , \7512 );
and \U$6787 ( \7516 , \7514 , \7515 );
buf \U$6788 ( \7517 , \4214 );
_DC g36d ( \7518_nG36d , \7517 , \7427 );
nor \U$6789 ( \7519 , \7516 , \7518_nG36d );
nor \U$6790 ( \7520 , \7513 , \7519 );
buf \U$6791 ( \7521 , \4185 );
_DC g350 ( \7522_nG350 , \7521 , \7427 );
and \U$6792 ( \7523 , \7520 , \7522_nG350 );
not \U$6793 ( \7524 , \7415 );
not \U$6794 ( \7525 , RIb54a540_3);
and \U$6795 ( \7526 , \7524 , \7525 );
and \U$6796 ( \7527 , \7415 , RIb54a540_3);
nor \U$6797 ( \7528 , \7526 , \7527 );
or \U$6798 ( \7529 , \7523 , \7528 );
or \U$6799 ( \7530 , \7435_nG334 , \7438 );
or \U$6800 ( \7531 , \7522_nG350 , \7520 );
nand \U$6801 ( \7532 , \7529 , \7530 , \7531 );
nand \U$6802 ( \7533 , \7440 , \7532 );
and \U$6803 ( \7534 , \7433_nG317 , \7533 );
and \U$6804 ( \7535 , \7417 , RIb54a450_1);
nor \U$6805 ( \7536 , \7533 , \7433_nG317 );
nor \U$6806 ( \7537 , \7417 , RIb54a450_1);
nor \U$6807 ( \7538 , \7535 , \7536 , \7537 );
nor \U$6808 ( \7539 , \7431 , \7534 , \7538 );
nor \U$6809 ( \7540 , \7430 , \7539 );
buf \U$6810 ( \7541 , \4128 );
_DC g495 ( \7542_nG495 , \7541 , \7402 );
buf \U$6811 ( \7543 , \1137 );
_DC g5cd ( \7544_nG5cd , \7543 , \7406 );
not \U$6812 ( \7545 , \7544_nG5cd );
not \U$6813 ( \7546 , \7545 );
buf \U$6814 ( \7547 , \4416 );
_DC g5cf ( \7548_nG5cf , \7547 , \7402 );
not \U$6815 ( \7549 , \7548_nG5cf );
and \U$6816 ( \7550 , \7546 , \7549 );
buf \U$6817 ( \7551 , \1170 );
_DC g5ee ( \7552_nG5ee , \7551 , \7406 );
nor \U$6818 ( \7553 , \7550 , \7552_nG5ee );
buf \U$6819 ( \7554 , \4444 );
_DC g5f0 ( \7555_nG5f0 , \7554 , \7402 );
and \U$6820 ( \7556 , \7553 , \7555_nG5f0 );
and \U$6821 ( \7557 , \7548_nG5cf , \7545 );
nor \U$6822 ( \7558 , \7556 , \7557 );
buf \U$6823 ( \7559 , \4387 );
_DC g5b0 ( \7560_nG5b0 , \7559 , \7402 );
not \U$6824 ( \7561 , \7560_nG5b0 );
buf \U$6825 ( \7562 , \1106 );
_DC g5ae ( \7563_nG5ae , \7562 , \7406 );
and \U$6826 ( \7564 , \7561 , \7563_nG5ae );
or \U$6827 ( \7565 , \7558 , \7564 );
or \U$6828 ( \7566 , \7563_nG5ae , \7561 );
nand \U$6829 ( \7567 , \7565 , \7566 );
buf \U$6830 ( \7568 , \4358 );
_DC g591 ( \7569_nG591 , \7568 , \7402 );
and \U$6831 ( \7570 , \7567 , \7569_nG591 );
not \U$6832 ( \7571 , \7567 );
not \U$6833 ( \7572 , \7569_nG591 );
and \U$6834 ( \7573 , \7571 , \7572 );
buf \U$6835 ( \7574 , \1074 );
_DC g58f ( \7575_nG58f , \7574 , \7406 );
nor \U$6836 ( \7576 , \7573 , \7575_nG58f );
nor \U$6837 ( \7577 , \7570 , \7576 );
buf \U$6838 ( \7578 , \1042 );
_DC g570 ( \7579_nG570 , \7578 , \7406 );
or \U$6839 ( \7580 , \7577 , \7579_nG570 );
not \U$6840 ( \7581 , \7579_nG570 );
not \U$6841 ( \7582 , \7577 );
or \U$6842 ( \7583 , \7581 , \7582 );
buf \U$6843 ( \7584 , \4329 );
_DC g572 ( \7585_nG572 , \7584 , \7402 );
nand \U$6844 ( \7586 , \7583 , \7585_nG572 );
nand \U$6845 ( \7587 , \7580 , \7586 );
buf \U$6846 ( \7588 , \4300 );
_DC g553 ( \7589_nG553 , \7588 , \7402 );
and \U$6847 ( \7590 , \7587 , \7589_nG553 );
not \U$6848 ( \7591 , \7587 );
not \U$6849 ( \7592 , \7589_nG553 );
and \U$6850 ( \7593 , \7591 , \7592 );
buf \U$6851 ( \7594 , \1006 );
_DC g551 ( \7595_nG551 , \7594 , \7406 );
nor \U$6852 ( \7596 , \7593 , \7595_nG551 );
nor \U$6853 ( \7597 , \7590 , \7596 );
buf \U$6854 ( \7598 , \4271 );
_DC g534 ( \7599_nG534 , \7598 , \7402 );
not \U$6855 ( \7600 , \7599_nG534 );
buf \U$6856 ( \7601 , \970 );
_DC g532 ( \7602_nG532 , \7601 , \7406 );
and \U$6857 ( \7603 , \7600 , \7602_nG532 );
or \U$6858 ( \7604 , \7597 , \7603 );
or \U$6859 ( \7605 , \7602_nG532 , \7600 );
nand \U$6860 ( \7606 , \7604 , \7605 );
buf \U$6861 ( \7607 , \4243 );
_DC g513 ( \7608_nG513 , \7607 , \7402 );
and \U$6862 ( \7609 , \7606 , \7608_nG513 );
not \U$6863 ( \7610 , \7606 );
not \U$6864 ( \7611 , \7608_nG513 );
and \U$6865 ( \7612 , \7610 , \7611 );
buf \U$6866 ( \7613 , \932 );
_DC g511 ( \7614_nG511 , \7613 , \7406 );
nor \U$6867 ( \7615 , \7612 , \7614_nG511 );
nor \U$6868 ( \7616 , \7609 , \7615 );
buf \U$6869 ( \7617 , \4214 );
_DC g4f4 ( \7618_nG4f4 , \7617 , \7402 );
not \U$6870 ( \7619 , \7618_nG4f4 );
buf \U$6871 ( \7620 , \896 );
_DC g4f2 ( \7621_nG4f2 , \7620 , \7406 );
and \U$6872 ( \7622 , \7619 , \7621_nG4f2 );
or \U$6873 ( \7623 , \7616 , \7622 );
or \U$6874 ( \7624 , \7621_nG4f2 , \7619 );
nand \U$6875 ( \7625 , \7623 , \7624 );
buf \U$6876 ( \7626 , \4185 );
_DC g4d3 ( \7627_nG4d3 , \7626 , \7402 );
and \U$6877 ( \7628 , \7625 , \7627_nG4d3 );
not \U$6878 ( \7629 , \7625 );
not \U$6879 ( \7630 , \7627_nG4d3 );
and \U$6880 ( \7631 , \7629 , \7630 );
buf \U$6881 ( \7632 , \858 );
_DC g4d1 ( \7633_nG4d1 , \7632 , \7406 );
nor \U$6882 ( \7634 , \7631 , \7633_nG4d1 );
nor \U$6883 ( \7635 , \7628 , \7634 );
buf \U$6884 ( \7636 , \4157 );
_DC g4b4 ( \7637_nG4b4 , \7636 , \7402 );
not \U$6885 ( \7638 , \7637_nG4b4 );
buf \U$6886 ( \7639 , \822 );
_DC g4b2 ( \7640_nG4b2 , \7639 , \7406 );
and \U$6887 ( \7641 , \7638 , \7640_nG4b2 );
or \U$6888 ( \7642 , \7635 , \7641 );
or \U$6889 ( \7643 , \7640_nG4b2 , \7638 );
nand \U$6890 ( \7644 , \7642 , \7643 );
and \U$6891 ( \7645 , \7542_nG495 , \7644 );
not \U$6892 ( \7646 , \7407_nG473 );
and \U$6893 ( \7647 , \7403_nG476 , \7646 );
not \U$6894 ( \7648 , \7644 );
not \U$6895 ( \7649 , \7542_nG495 );
and \U$6896 ( \7650 , \7648 , \7649 );
buf \U$6897 ( \7651 , \786 );
_DC g493 ( \7652_nG493 , \7651 , \7406 );
nor \U$6898 ( \7653 , \7650 , \7652_nG493 );
nor \U$6899 ( \7654 , \7645 , \7647 , \7653 );
nor \U$6900 ( \7655 , \7408 , \7540 , \7654 );
not \U$6901 ( \7656 , \682 );
nand \U$6902 ( \7657 , \7656 , RIb54a9f0_13);
and \U$6903 ( \7658 , \7655 , \679 , \7657 );
_HMUX g2231_GF_PartitionCandidate ( \7659_nG2231 , \4070 , \7400 , \7658 );
buf \U$6904 ( \7660 , \7659_nG2231 );
xor \U$6905 ( \7661 , \1565 , \1566 );
xor \U$6906 ( \7662 , \7661 , \4063 );
xor \U$6907 ( \7663 , \4834 , \4835 );
xor \U$6908 ( \7664 , \7663 , \7393 );
_HMUX g21f6_GF_PartitionCandidate ( \7665_nG21f6 , \7662 , \7664 , \7658 );
buf \U$6909 ( \7666 , \7665_nG21f6 );
xor \U$6910 ( \7667 , \1569 , \1740 );
xor \U$6911 ( \7668 , \7667 , \4060 );
xor \U$6912 ( \7669 , \5010 , \5017 );
xor \U$6913 ( \7670 , \7669 , \7389 );
not \U$6914 ( \7671 , \7670 );
_HMUX g21c6_GF_PartitionCandidate ( \7672_nG21c6 , \7668 , \7671 , \7658 );
buf \U$6915 ( \7673 , \7672_nG21c6 );
xor \U$6916 ( \7674 , \1743 , \1849 );
xor \U$6917 ( \7675 , \7674 , \4057 );
xor \U$6918 ( \7676 , \4841 , \4843 );
xor \U$6919 ( \7677 , \7676 , \5007 );
xor \U$6920 ( \7678 , \5120 , \7384 );
xor \U$6921 ( \7679 , \7677 , \7678 );
not \U$6922 ( \7680 , \7679 );
_HMUX g2179_GF_PartitionCandidate ( \7681_nG2179 , \7675 , \7680 , \7658 );
buf \U$6923 ( \7682 , \7681_nG2179 );
xor \U$6924 ( \7683 , \1935 , \1937 );
xor \U$6925 ( \7684 , \7683 , \4054 );
not \U$6926 ( \7685 , \7383 );
nand \U$6927 ( \7686 , \7685 , \7381 );
not \U$6928 ( \7687 , \7686 );
not \U$6929 ( \7688 , \7374 );
or \U$6930 ( \7689 , \7687 , \7688 );
or \U$6931 ( \7690 , \7374 , \7686 );
nand \U$6932 ( \7691 , \7689 , \7690 );
_HMUX g2115_GF_PartitionCandidate ( \7692_nG2115 , \7684 , \7691 , \7658 );
buf \U$6933 ( \7693 , \7692_nG2115 );
xor \U$6934 ( \7694 , \1940 , \2048 );
xor \U$6935 ( \7695 , \7694 , \4051 );
xor \U$6936 ( \7696 , \5220 , \5335 );
xor \U$6937 ( \7697 , \7696 , \7371 );
_HMUX g209c_GF_PartitionCandidate ( \7698_nG209c , \7695 , \7697 , \7658 );
buf \U$6938 ( \7699 , \7698_nG209c );
xor \U$6939 ( \7700 , \2156 , \2160 );
xor \U$6940 ( \7701 , \7700 , \4048 );
xor \U$6941 ( \7702 , \5445 , \5449 );
xor \U$6942 ( \7703 , \7702 , \7368 );
_HMUX g2013_GF_PartitionCandidate ( \7704_nG2013 , \7701 , \7703 , \7658 );
buf \U$6943 ( \7705 , \7704_nG2013 );
xor \U$6944 ( \7706 , \2163 , \2301 );
xor \U$6945 ( \7707 , \7706 , \4045 );
not \U$6946 ( \7708 , \7366 );
nand \U$6947 ( \7709 , \7708 , \7364 );
not \U$6948 ( \7710 , \7709 );
not \U$6949 ( \7711 , \7354 );
or \U$6950 ( \7712 , \7710 , \7711 );
or \U$6951 ( \7713 , \7354 , \7709 );
nand \U$6952 ( \7714 , \7712 , \7713 );
_HMUX g1f8e_GF_PartitionCandidate ( \7715_nG1f8e , \7707 , \7714 , \7658 );
buf \U$6953 ( \7716 , \7715_nG1f8e );
not \U$6954 ( \7717 , \4043 );
nand \U$6955 ( \7718 , \7717 , \4041 );
not \U$6956 ( \7719 , \7718 );
not \U$6957 ( \7720 , \4029 );
or \U$6958 ( \7721 , \7719 , \7720 );
or \U$6959 ( \7722 , \4029 , \7718 );
nand \U$6960 ( \7723 , \7721 , \7722 );
xor \U$6961 ( \7724 , \5734 , \5754 );
xor \U$6962 ( \7725 , \7724 , \7351 );
_HMUX g1eef_GF_PartitionCandidate ( \7726_nG1eef , \7723 , \7725 , \7658 );
buf \U$6963 ( \7727 , \7726_nG1eef );
xor \U$6964 ( \7728 , \2470 , \2583 );
xor \U$6965 ( \7729 , \7728 , \4026 );
xor \U$6966 ( \7730 , \5865 , \5762 );
not \U$6967 ( \7731 , \7730 );
not \U$6968 ( \7732 , \7348 );
or \U$6969 ( \7733 , \7731 , \7732 );
or \U$6970 ( \7734 , \7348 , \7730 );
nand \U$6971 ( \7735 , \7733 , \7734 );
_HMUX g1e25_GF_PartitionCandidate ( \7736_nG1e25 , \7729 , \7735 , \7658 );
buf \U$6972 ( \7737 , \7736_nG1e25 );
xor \U$6973 ( \7738 , \2746 , \2748 );
xor \U$6974 ( \7739 , \7738 , \4023 );
not \U$6975 ( \7740 , \7347 );
nand \U$6976 ( \7741 , \7740 , \7345 );
not \U$6977 ( \7742 , \7741 );
not \U$6978 ( \7743 , \7330 );
or \U$6979 ( \7744 , \7742 , \7743 );
or \U$6980 ( \7745 , \7330 , \7741 );
nand \U$6981 ( \7746 , \7744 , \7745 );
_HMUX g1d58_GF_PartitionCandidate ( \7747_nG1d58 , \7739 , \7746 , \7658 );
buf \U$6982 ( \7748 , \7747_nG1d58 );
xor \U$6983 ( \7749 , \2820 , \2822 );
xor \U$6984 ( \7750 , \7749 , \4020 );
xor \U$6985 ( \7751 , \6045 , \6128 );
xor \U$6986 ( \7752 , \7751 , \7327 );
_HMUX g1c7b_GF_PartitionCandidate ( \7753_nG1c7b , \7750 , \7752 , \7658 );
buf \U$6987 ( \7754 , \7753_nG1c7b );
xor \U$6988 ( \7755 , \2825 , \2994 );
xor \U$6989 ( \7756 , \7755 , \4017 );
xor \U$6990 ( \7757 , \6131 , \6308 );
xor \U$6991 ( \7758 , \7757 , \7324 );
_HMUX g1baa_GF_PartitionCandidate ( \7759_nG1baa , \7756 , \7758 , \7658 );
buf \U$6992 ( \7760 , \7759_nG1baa );
xor \U$6993 ( \7761 , \2997 , \3077 );
xor \U$6994 ( \7762 , \7761 , \4014 );
xor \U$6995 ( \7763 , \6311 , \6402 );
xor \U$6996 ( \7764 , \7763 , \7321 );
_HMUX g1ad8_GF_PartitionCandidate ( \7765_nG1ad8 , \7762 , \7764 , \7658 );
buf \U$6997 ( \7766 , \7765_nG1ad8 );
xor \U$6998 ( \7767 , \3080 , \3249 );
xor \U$6999 ( \7768 , \7767 , \4011 );
xor \U$7000 ( \7769 , \6407 , \6567 );
xor \U$7001 ( \7770 , \7769 , \7318 );
_HMUX g19f9_GF_PartitionCandidate ( \7771_nG19f9 , \7768 , \7770 , \7658 );
buf \U$7002 ( \7772 , \7771_nG19f9 );
xor \U$7003 ( \7773 , \3252 , \3265 );
xor \U$7004 ( \7774 , \7773 , \4008 );
xor \U$7005 ( \7775 , \6570 , \6577 );
xor \U$7006 ( \7776 , \7775 , \7315 );
_HMUX g18ff_GF_PartitionCandidate ( \7777_nG18ff , \7774 , \7776 , \7658 );
buf \U$7007 ( \7778 , \7777_nG18ff );
xor \U$7008 ( \7779 , \3268 , \3350 );
xor \U$7009 ( \7780 , \7779 , \4005 );
xor \U$7010 ( \7781 , \6580 , \6657 );
xor \U$7011 ( \7782 , \7781 , \7312 );
_HMUX g17ec_GF_PartitionCandidate ( \7783_nG17ec , \7780 , \7782 , \7658 );
buf \U$7012 ( \7784 , \7783_nG17ec );
xor \U$7013 ( \7785 , \3353 , \3428 );
xor \U$7014 ( \7786 , \7785 , \4002 );
xor \U$7015 ( \7787 , \6661 , \6741 );
xor \U$7016 ( \7788 , \7787 , \7309 );
_HMUX g16f6_GF_PartitionCandidate ( \7789_nG16f6 , \7786 , \7788 , \7658 );
buf \U$7017 ( \7790 , \7789_nG16f6 );
xor \U$7018 ( \7791 , \3436 , \3526 );
xor \U$7019 ( \7792 , \7791 , \3998 );
not \U$7020 ( \7793 , \7792 );
xor \U$7021 ( \7794 , \6749 , \6839 );
xor \U$7022 ( \7795 , \7794 , \7305 );
not \U$7023 ( \7796 , \7795 );
_HMUX g15de_GF_PartitionCandidate ( \7797_nG15de , \7793 , \7796 , \7658 );
buf \U$7024 ( \7798 , \7797_nG15de );
not \U$7025 ( \7799 , \3997 );
nand \U$7026 ( \7800 , \7799 , \3995 );
not \U$7027 ( \7801 , \7800 );
not \U$7028 ( \7802 , \3988 );
or \U$7029 ( \7803 , \7801 , \7802 );
or \U$7030 ( \7804 , \3988 , \7800 );
nand \U$7031 ( \7805 , \7803 , \7804 );
not \U$7032 ( \7806 , \7304 );
nand \U$7033 ( \7807 , \7806 , \7302 );
not \U$7034 ( \7808 , \7807 );
not \U$7035 ( \7809 , \7295 );
or \U$7036 ( \7810 , \7808 , \7809 );
or \U$7037 ( \7811 , \7295 , \7807 );
nand \U$7038 ( \7812 , \7810 , \7811 );
_HMUX g14d2_GF_PartitionCandidate ( \7813_nG14d2 , \7805 , \7812 , \7658 );
buf \U$7039 ( \7814 , \7813_nG14d2 );
xor \U$7040 ( \7815 , \3590 , \3637 );
xor \U$7041 ( \7816 , \7815 , \3985 );
xor \U$7042 ( \7817 , \6903 , \6952 );
xor \U$7043 ( \7818 , \7817 , \7292 );
_HMUX g13d7_GF_PartitionCandidate ( \7819_nG13d7 , \7816 , \7818 , \7658 );
buf \U$7044 ( \7820 , \7819_nG13d7 );
xor \U$7045 ( \7821 , \3640 , \3709 );
xor \U$7046 ( \7822 , \7821 , \3982 );
xor \U$7047 ( \7823 , \6955 , \7028 );
xor \U$7048 ( \7824 , \7823 , \7289 );
_HMUX g12e5_GF_PartitionCandidate ( \7825_nG12e5 , \7822 , \7824 , \7658 );
buf \U$7049 ( \7826 , \7825_nG12e5 );
xor \U$7050 ( \7827 , \3974 , \3976 );
xor \U$7051 ( \7828 , \7827 , \3979 );
xor \U$7052 ( \7829 , \7282 , \7283 );
xor \U$7053 ( \7830 , \7829 , \7286 );
_HMUX g11da_GF_PartitionCandidate ( \7831_nG11da , \7828 , \7830 , \7658 );
buf \U$7054 ( \7832 , \7831_nG11da );
nor \U$7055 ( \7833 , \3972 , \3969 );
not \U$7056 ( \7834 , \7833 );
not \U$7057 ( \7835 , \3943 );
or \U$7058 ( \7836 , \7834 , \7835 );
or \U$7059 ( \7837 , \3943 , \7833 );
nand \U$7060 ( \7838 , \7836 , \7837 );
xor \U$7061 ( \7839 , \7042 , \7083 );
xor \U$7062 ( \7840 , \7839 , \7279 );
_HMUX g10fb_GF_PartitionCandidate ( \7841_nG10fb , \7838 , \7840 , \7658 );
buf \U$7063 ( \7842 , \7841_nG10fb );
not \U$7064 ( \7843 , \3939 );
nand \U$7065 ( \7844 , \7843 , \3942 );
not \U$7066 ( \7845 , \7844 );
not \U$7067 ( \7846 , \3920 );
or \U$7068 ( \7847 , \7845 , \7846 );
or \U$7069 ( \7848 , \3920 , \7844 );
nand \U$7070 ( \7849 , \7847 , \7848 );
xor \U$7071 ( \7850 , \7091 , \7135 );
xor \U$7072 ( \7851 , \7850 , \7276 );
_HMUX gfed_GF_PartitionCandidate ( \7852_nGfed , \7849 , \7851 , \7658 );
buf \U$7073 ( \7853 , \7852_nGfed );
xor \U$7074 ( \7854 , \3900 , \3901 );
xor \U$7075 ( \7855 , \7854 , \3917 );
xor \U$7076 ( \7856 , \7270 , \7266 );
xor \U$7077 ( \7857 , \7856 , \7273 );
_HMUX gf15_GF_PartitionCandidate ( \7858_nGf15 , \7855 , \7857 , \7658 );
buf \U$7078 ( \7859 , \7858_nGf15 );
xor \U$7079 ( \7860 , \3777 , \3814 );
xor \U$7080 ( \7861 , \7860 , \3897 );
xor \U$7081 ( \7862 , \7256 , \7259 );
xor \U$7082 ( \7863 , \7862 , \7267 );
_HMUX ge3d_GF_PartitionCandidate ( \7864_nGe3d , \7861 , \7863 , \7658 );
buf \U$7083 ( \7865 , \7864_nGe3d );
nand \U$7084 ( \7866 , RIb55bca0_599, RIb55bc28_598);
not \U$7085 ( \7867 , \7866 );
nand \U$7086 ( \7868 , \7867 , RIb55bbb0_597);
not \U$7087 ( \7869 , \7868 );
nand \U$7088 ( \7870 , \7869 , RIb55bb38_596);
not \U$7089 ( \7871 , \7870 );
nand \U$7090 ( \7872 , \7871 , RIb55bac0_595);
not \U$7091 ( \7873 , \7872 );
nand \U$7092 ( \7874 , \7873 , RIb55ba48_594);
not \U$7093 ( \7875 , \7874 );
nand \U$7094 ( \7876 , \7875 , RIb55b9d0_593);
not \U$7095 ( \7877 , \7876 );
nand \U$7096 ( \7878 , \7877 , RIb55b958_592);
not \U$7097 ( \7879 , \7878 );
nand \U$7098 ( \7880 , \7879 , RIb55b8e0_591);
not \U$7099 ( \7881 , \7880 );
nand \U$7100 ( \7882 , \7881 , RIb55b868_590);
not \U$7101 ( \7883 , \7882 );
nand \U$7102 ( \7884 , \7883 , RIb55b7f0_589);
not \U$7103 ( \7885 , \7884 );
not \U$7104 ( \7886 , RIb55c3a8_614);
and \U$7105 ( \7887 , \7885 , \7886 );
and \U$7106 ( \7888 , \7884 , RIb55c3a8_614);
nor \U$7107 ( \7889 , \7887 , \7888 );
not \U$7108 ( \7890 , RIb55be08_602);
nor \U$7109 ( \7891 , RIb55bfe8_606, RIb55c1c8_610);
not \U$7110 ( \7892 , \7891 );
or \U$7111 ( \7893 , RIb55c0d8_608, RIb55c150_609, RIb55c240_611, RIb55c2b8_612);
nor \U$7112 ( \7894 , \7892 , \7893 , RIb55c060_607, RIb55c330_613);
not \U$7113 ( \7895 , \7894 );
nor \U$7114 ( \7896 , \7895 , RIb55bef8_604);
nand \U$7115 ( \7897 , \7890 , \7896 );
and \U$7116 ( \7898 , RIb55bd18_600, RIb55bd90_601);
nand \U$7117 ( \7899 , RIb55be80_603, \7898 );
nor \U$7118 ( \7900 , \7897 , \7899 );
and \U$7119 ( \7901 , \7900 , RIb551a70_253);
not \U$7120 ( \7902 , RIb55be80_603);
nor \U$7121 ( \7903 , \7897 , \7902 );
not \U$7122 ( \7904 , RIb55bd18_600);
nor \U$7123 ( \7905 , \7904 , RIb55bd90_601);
and \U$7124 ( \7906 , \7903 , \7905 );
and \U$7125 ( \7907 , \7906 , RIb551b60_255);
nand \U$7126 ( \7908 , RIb55be08_602, \7896 );
nor \U$7127 ( \7909 , \7908 , RIb55be80_603);
and \U$7128 ( \7910 , \7909 , \7898 );
and \U$7129 ( \7911 , RIb551c50_257, \7910 );
nor \U$7130 ( \7912 , \7907 , \7911 );
nor \U$7131 ( \7913 , RIb55bd18_600, RIb55bd90_601);
and \U$7132 ( \7914 , \7903 , \7913 );
and \U$7133 ( \7915 , \7914 , RIb551bd8_256);
nor \U$7134 ( \7916 , \7908 , \7902 );
and \U$7135 ( \7917 , \7916 , \7905 );
and \U$7136 ( \7918 , RIb551980_251, \7917 );
nor \U$7137 ( \7919 , \7915 , \7918 );
and \U$7138 ( \7920 , \7904 , RIb55bd90_601);
and \U$7139 ( \7921 , \7916 , \7920 );
and \U$7140 ( \7922 , \7921 , RIb551908_250);
nor \U$7141 ( \7923 , \7908 , \7899 );
and \U$7142 ( \7924 , RIb551890_249, \7923 );
nor \U$7143 ( \7925 , \7922 , \7924 );
and \U$7144 ( \7926 , \7909 , \7920 );
and \U$7145 ( \7927 , \7926 , RIb551cc8_258);
not \U$7146 ( \7928 , \7913 );
nor \U$7147 ( \7929 , \7928 , RIb55be80_603, RIb55be08_602);
and \U$7148 ( \7930 , \7929 , \7894 , RIb55bef8_604);
nand \U$7149 ( \7931 , RIb551818_248, \7930 );
not \U$7150 ( \7932 , \7931 );
nor \U$7151 ( \7933 , \7927 , \7932 );
nand \U$7152 ( \7934 , \7912 , \7919 , \7925 , \7933 );
nor \U$7153 ( \7935 , \7897 , RIb55be80_603);
and \U$7154 ( \7936 , \7935 , \7905 );
and \U$7155 ( \7937 , \7936 , RIb551f20_263);
and \U$7156 ( \7938 , \7935 , \7920 );
and \U$7157 ( \7939 , RIb551ea8_262, \7938 );
nor \U$7158 ( \7940 , \7937 , \7939 );
not \U$7159 ( \7941 , \7940 );
nor \U$7160 ( \7942 , \7901 , \7934 , \7941 );
and \U$7161 ( \7943 , \7909 , \7913 );
and \U$7162 ( \7944 , \7943 , RIb551db8_260);
and \U$7163 ( \7945 , \7935 , \7898 );
and \U$7164 ( \7946 , RIb551e30_261, \7945 );
nor \U$7165 ( \7947 , \7944 , \7946 );
and \U$7166 ( \7948 , \7896 , \7929 );
and \U$7167 ( \7949 , \7948 , RIb551f98_264);
and \U$7168 ( \7950 , \7916 , \7913 );
and \U$7169 ( \7951 , RIb5519f8_252, \7950 );
nor \U$7170 ( \7952 , \7949 , \7951 );
and \U$7171 ( \7953 , \7903 , \7920 );
and \U$7172 ( \7954 , \7953 , RIb551ae8_254);
and \U$7173 ( \7955 , \7909 , \7905 );
and \U$7174 ( \7956 , RIb551d40_259, \7955 );
nor \U$7175 ( \7957 , \7954 , \7956 );
nand \U$7176 ( \7958 , \7942 , \7947 , \7952 , \7957 );
buf \U$7177 ( \7959 , \7958 );
not \U$7178 ( \7960 , \7929 );
nand \U$7179 ( \7961 , \7960 , RIb55bef8_604);
nand \U$7180 ( \7962 , \7961 , \7894 );
buf \U$7181 ( \7963 , \7962 );
_DC g2ace ( \7964_nG2ace , \7959 , \7963 );
xor \U$7182 ( \7965 , \7889 , \7964_nG2ace );
not \U$7183 ( \7966 , \7882 );
not \U$7184 ( \7967 , RIb55b7f0_589);
and \U$7185 ( \7968 , \7966 , \7967 );
and \U$7186 ( \7969 , \7882 , RIb55b7f0_589);
nor \U$7187 ( \7970 , \7968 , \7969 );
and \U$7188 ( \7971 , \7923 , RIb54ac48_18);
and \U$7189 ( \7972 , RIb54b1e8_30, \7945 );
and \U$7190 ( \7973 , \7938 , RIb54b260_31);
and \U$7191 ( \7974 , RIb54ae28_22, \7900 );
nor \U$7192 ( \7975 , \7972 , \7973 , \7974 );
and \U$7193 ( \7976 , \7953 , RIb54aea0_23);
and \U$7194 ( \7977 , RIb54adb0_21, \7950 );
nor \U$7195 ( \7978 , \7976 , \7977 );
and \U$7196 ( \7979 , \7948 , RIb54b350_33);
and \U$7197 ( \7980 , RIb54b2d8_32, \7936 );
nor \U$7198 ( \7981 , \7979 , \7980 );
and \U$7199 ( \7982 , \7943 , RIb54b170_29);
and \U$7200 ( \7983 , RIb54b0f8_28, \7955 );
nor \U$7201 ( \7984 , \7982 , \7983 );
nand \U$7202 ( \7985 , \7975 , \7978 , \7981 , \7984 );
nand \U$7203 ( \7986 , RIb54a978_12, \7930 );
not \U$7204 ( \7987 , \7986 );
nor \U$7205 ( \7988 , \7971 , \7985 , \7987 );
and \U$7206 ( \7989 , \7914 , RIb54af90_25);
and \U$7207 ( \7990 , RIb54af18_24, \7906 );
nor \U$7208 ( \7991 , \7989 , \7990 );
and \U$7209 ( \7992 , \7917 , RIb54ad38_20);
and \U$7210 ( \7993 , RIb54acc0_19, \7921 );
nor \U$7211 ( \7994 , \7992 , \7993 );
and \U$7212 ( \7995 , \7926 , RIb54b080_27);
and \U$7213 ( \7996 , RIb54b008_26, \7910 );
nor \U$7214 ( \7997 , \7995 , \7996 );
nand \U$7215 ( \7998 , \7988 , \7991 , \7994 , \7997 );
buf \U$7216 ( \7999 , \7998 );
_DC g28f2 ( \8000_nG28f2 , \7999 , \7963 );
xor \U$7217 ( \8001 , \7970 , \8000_nG28f2 );
not \U$7218 ( \8002 , \7880 );
not \U$7219 ( \8003 , RIb55b868_590);
and \U$7220 ( \8004 , \8002 , \8003 );
and \U$7221 ( \8005 , \7880 , RIb55b868_590);
nor \U$7222 ( \8006 , \8004 , \8005 );
and \U$7223 ( \8007 , \7900 , RIb54b620_39);
and \U$7224 ( \8008 , \7906 , RIb54b710_41);
and \U$7225 ( \8009 , RIb54b800_43, \7910 );
nor \U$7226 ( \8010 , \8008 , \8009 );
and \U$7227 ( \8011 , \7914 , RIb54b788_42);
and \U$7228 ( \8012 , RIb54b530_37, \7917 );
nor \U$7229 ( \8013 , \8011 , \8012 );
and \U$7230 ( \8014 , \7921 , RIb54b4b8_36);
and \U$7231 ( \8015 , RIb54b440_35, \7923 );
nor \U$7232 ( \8016 , \8014 , \8015 );
and \U$7233 ( \8017 , \7926 , RIb54b878_44);
nand \U$7234 ( \8018 , RIb54b3c8_34, \7930 );
not \U$7235 ( \8019 , \8018 );
nor \U$7236 ( \8020 , \8017 , \8019 );
nand \U$7237 ( \8021 , \8010 , \8013 , \8016 , \8020 );
and \U$7238 ( \8022 , \7936 , RIb54bad0_49);
and \U$7239 ( \8023 , RIb54ba58_48, \7938 );
nor \U$7240 ( \8024 , \8022 , \8023 );
not \U$7241 ( \8025 , \8024 );
nor \U$7242 ( \8026 , \8007 , \8021 , \8025 );
and \U$7243 ( \8027 , \7943 , RIb54b968_46);
and \U$7244 ( \8028 , RIb54b9e0_47, \7945 );
nor \U$7245 ( \8029 , \8027 , \8028 );
and \U$7246 ( \8030 , \7948 , RIb54bb48_50);
and \U$7247 ( \8031 , RIb54b5a8_38, \7950 );
nor \U$7248 ( \8032 , \8030 , \8031 );
and \U$7249 ( \8033 , \7953 , RIb54b698_40);
and \U$7250 ( \8034 , RIb54b8f0_45, \7955 );
nor \U$7251 ( \8035 , \8033 , \8034 );
nand \U$7252 ( \8036 , \8026 , \8029 , \8032 , \8035 );
buf \U$7253 ( \8037 , \8036 );
_DC g28f0 ( \8038_nG28f0 , \8037 , \7963 );
xor \U$7254 ( \8039 , \8006 , \8038_nG28f0 );
not \U$7255 ( \8040 , \7878 );
not \U$7256 ( \8041 , RIb55b8e0_591);
and \U$7257 ( \8042 , \8040 , \8041 );
and \U$7258 ( \8043 , \7878 , RIb55b8e0_591);
nor \U$7259 ( \8044 , \8042 , \8043 );
and \U$7260 ( \8045 , \7900 , RIb54be18_56);
and \U$7261 ( \8046 , \7906 , RIb54bf08_58);
and \U$7262 ( \8047 , RIb54bff8_60, \7910 );
nor \U$7263 ( \8048 , \8046 , \8047 );
and \U$7264 ( \8049 , \7914 , RIb54bf80_59);
and \U$7265 ( \8050 , RIb54bd28_54, \7917 );
nor \U$7266 ( \8051 , \8049 , \8050 );
and \U$7267 ( \8052 , \7921 , RIb54bcb0_53);
and \U$7268 ( \8053 , RIb54bc38_52, \7923 );
nor \U$7269 ( \8054 , \8052 , \8053 );
and \U$7270 ( \8055 , \7926 , RIb54c070_61);
nand \U$7271 ( \8056 , RIb54bbc0_51, \7930 );
not \U$7272 ( \8057 , \8056 );
nor \U$7273 ( \8058 , \8055 , \8057 );
nand \U$7274 ( \8059 , \8048 , \8051 , \8054 , \8058 );
and \U$7275 ( \8060 , \7936 , RIb54c2c8_66);
and \U$7276 ( \8061 , RIb54c250_65, \7938 );
nor \U$7277 ( \8062 , \8060 , \8061 );
not \U$7278 ( \8063 , \8062 );
nor \U$7279 ( \8064 , \8045 , \8059 , \8063 );
and \U$7280 ( \8065 , \7943 , RIb54c160_63);
and \U$7281 ( \8066 , RIb54c1d8_64, \7945 );
nor \U$7282 ( \8067 , \8065 , \8066 );
and \U$7283 ( \8068 , \7948 , RIb54c340_67);
and \U$7284 ( \8069 , RIb54bda0_55, \7950 );
nor \U$7285 ( \8070 , \8068 , \8069 );
and \U$7286 ( \8071 , \7953 , RIb54be90_57);
and \U$7287 ( \8072 , RIb54c0e8_62, \7955 );
nor \U$7288 ( \8073 , \8071 , \8072 );
nand \U$7289 ( \8074 , \8064 , \8067 , \8070 , \8073 );
buf \U$7290 ( \8075 , \8074 );
_DC g273d ( \8076_nG273d , \8075 , \7963 );
xor \U$7291 ( \8077 , \8044 , \8076_nG273d );
not \U$7292 ( \8078 , \7876 );
not \U$7293 ( \8079 , RIb55b958_592);
and \U$7294 ( \8080 , \8078 , \8079 );
and \U$7295 ( \8081 , \7876 , RIb55b958_592);
nor \U$7296 ( \8082 , \8080 , \8081 );
and \U$7297 ( \8083 , \7923 , RIb54c430_69);
and \U$7298 ( \8084 , RIb54c9d0_81, \7945 );
and \U$7299 ( \8085 , \7938 , RIb54ca48_82);
and \U$7300 ( \8086 , RIb54c610_73, \7900 );
nor \U$7301 ( \8087 , \8084 , \8085 , \8086 );
and \U$7302 ( \8088 , \7953 , RIb54c688_74);
and \U$7303 ( \8089 , RIb54c598_72, \7950 );
nor \U$7304 ( \8090 , \8088 , \8089 );
and \U$7305 ( \8091 , \7948 , RIb54cb38_84);
and \U$7306 ( \8092 , RIb54cac0_83, \7936 );
nor \U$7307 ( \8093 , \8091 , \8092 );
and \U$7308 ( \8094 , \7943 , RIb54c958_80);
and \U$7309 ( \8095 , RIb54c8e0_79, \7955 );
nor \U$7310 ( \8096 , \8094 , \8095 );
nand \U$7311 ( \8097 , \8087 , \8090 , \8093 , \8096 );
nand \U$7312 ( \8098 , RIb54c3b8_68, \7930 );
not \U$7313 ( \8099 , \8098 );
nor \U$7314 ( \8100 , \8083 , \8097 , \8099 );
and \U$7315 ( \8101 , \7914 , RIb54c778_76);
and \U$7316 ( \8102 , RIb54c700_75, \7906 );
nor \U$7317 ( \8103 , \8101 , \8102 );
and \U$7318 ( \8104 , \7917 , RIb54c520_71);
and \U$7319 ( \8105 , RIb54c4a8_70, \7921 );
nor \U$7320 ( \8106 , \8104 , \8105 );
and \U$7321 ( \8107 , \7926 , RIb54c868_78);
and \U$7322 ( \8108 , RIb54c7f0_77, \7910 );
nor \U$7323 ( \8109 , \8107 , \8108 );
nand \U$7324 ( \8110 , \8100 , \8103 , \8106 , \8109 );
buf \U$7325 ( \8111 , \8110 );
_DC g273b ( \8112_nG273b , \8111 , \7963 );
xor \U$7326 ( \8113 , \8082 , \8112_nG273b );
and \U$7327 ( \8114 , \7874 , RIb55b9d0_593);
not \U$7328 ( \8115 , \7874 );
not \U$7329 ( \8116 , RIb55b9d0_593);
and \U$7330 ( \8117 , \8115 , \8116 );
nor \U$7331 ( \8118 , \8114 , \8117 );
and \U$7332 ( \8119 , \7900 , RIb54ce08_90);
and \U$7333 ( \8120 , \7906 , RIb54cef8_92);
and \U$7334 ( \8121 , RIb54cfe8_94, \7910 );
nor \U$7335 ( \8122 , \8120 , \8121 );
and \U$7336 ( \8123 , \7914 , RIb54cf70_93);
and \U$7337 ( \8124 , RIb54cd18_88, \7917 );
nor \U$7338 ( \8125 , \8123 , \8124 );
and \U$7339 ( \8126 , \7921 , RIb54cca0_87);
and \U$7340 ( \8127 , RIb54cc28_86, \7923 );
nor \U$7341 ( \8128 , \8126 , \8127 );
and \U$7342 ( \8129 , \7926 , RIb54d060_95);
nand \U$7343 ( \8130 , RIb54cbb0_85, \7930 );
not \U$7344 ( \8131 , \8130 );
nor \U$7345 ( \8132 , \8129 , \8131 );
nand \U$7346 ( \8133 , \8122 , \8125 , \8128 , \8132 );
and \U$7347 ( \8134 , \7936 , RIb54d2b8_100);
and \U$7348 ( \8135 , RIb54d240_99, \7938 );
nor \U$7349 ( \8136 , \8134 , \8135 );
not \U$7350 ( \8137 , \8136 );
nor \U$7351 ( \8138 , \8119 , \8133 , \8137 );
and \U$7352 ( \8139 , \7943 , RIb54d150_97);
and \U$7353 ( \8140 , RIb54d1c8_98, \7945 );
nor \U$7354 ( \8141 , \8139 , \8140 );
and \U$7355 ( \8142 , \7948 , RIb54d330_101);
and \U$7356 ( \8143 , RIb54cd90_89, \7950 );
nor \U$7357 ( \8144 , \8142 , \8143 );
and \U$7358 ( \8145 , \7953 , RIb54ce80_91);
and \U$7359 ( \8146 , RIb54d0d8_96, \7955 );
nor \U$7360 ( \8147 , \8145 , \8146 );
nand \U$7361 ( \8148 , \8138 , \8141 , \8144 , \8147 );
buf \U$7362 ( \8149 , \8148 );
_DC g25c7 ( \8150_nG25c7 , \8149 , \7963 );
xor \U$7363 ( \8151 , \8118 , \8150_nG25c7 );
not \U$7364 ( \8152 , \7872 );
not \U$7365 ( \8153 , RIb55ba48_594);
and \U$7366 ( \8154 , \8152 , \8153 );
and \U$7367 ( \8155 , \7872 , RIb55ba48_594);
nor \U$7368 ( \8156 , \8154 , \8155 );
and \U$7369 ( \8157 , \7900 , RIb54d600_107);
and \U$7370 ( \8158 , \7906 , RIb54d6f0_109);
and \U$7371 ( \8159 , RIb54d7e0_111, \7910 );
nor \U$7372 ( \8160 , \8158 , \8159 );
and \U$7373 ( \8161 , \7914 , RIb54d768_110);
and \U$7374 ( \8162 , RIb54d510_105, \7917 );
nor \U$7375 ( \8163 , \8161 , \8162 );
and \U$7376 ( \8164 , \7921 , RIb54d498_104);
and \U$7377 ( \8165 , RIb54d420_103, \7923 );
nor \U$7378 ( \8166 , \8164 , \8165 );
and \U$7379 ( \8167 , \7926 , RIb54d858_112);
nand \U$7380 ( \8168 , RIb54d3a8_102, \7930 );
not \U$7381 ( \8169 , \8168 );
nor \U$7382 ( \8170 , \8167 , \8169 );
nand \U$7383 ( \8171 , \8160 , \8163 , \8166 , \8170 );
and \U$7384 ( \8172 , \7936 , RIb54dab0_117);
and \U$7385 ( \8173 , RIb54da38_116, \7938 );
nor \U$7386 ( \8174 , \8172 , \8173 );
not \U$7387 ( \8175 , \8174 );
nor \U$7388 ( \8176 , \8157 , \8171 , \8175 );
and \U$7389 ( \8177 , \7943 , RIb54d948_114);
and \U$7390 ( \8178 , RIb54d9c0_115, \7945 );
nor \U$7391 ( \8179 , \8177 , \8178 );
and \U$7392 ( \8180 , \7948 , RIb54db28_118);
and \U$7393 ( \8181 , RIb54d588_106, \7950 );
nor \U$7394 ( \8182 , \8180 , \8181 );
and \U$7395 ( \8183 , \7953 , RIb54d678_108);
and \U$7396 ( \8184 , RIb54d8d0_113, \7955 );
nor \U$7397 ( \8185 , \8183 , \8184 );
nand \U$7398 ( \8186 , \8176 , \8179 , \8182 , \8185 );
buf \U$7399 ( \8187 , \8186 );
_DC g25c5 ( \8188_nG25c5 , \8187 , \7963 );
xor \U$7400 ( \8189 , \8156 , \8188_nG25c5 );
not \U$7401 ( \8190 , \7870 );
not \U$7402 ( \8191 , RIb55bac0_595);
and \U$7403 ( \8192 , \8190 , \8191 );
and \U$7404 ( \8193 , \7870 , RIb55bac0_595);
nor \U$7405 ( \8194 , \8192 , \8193 );
and \U$7406 ( \8195 , \7900 , RIb54ddf8_124);
and \U$7407 ( \8196 , \7906 , RIb54dee8_126);
and \U$7408 ( \8197 , RIb54dfd8_128, \7910 );
nor \U$7409 ( \8198 , \8196 , \8197 );
and \U$7410 ( \8199 , \7914 , RIb54df60_127);
and \U$7411 ( \8200 , RIb54dd08_122, \7917 );
nor \U$7412 ( \8201 , \8199 , \8200 );
and \U$7413 ( \8202 , \7921 , RIb54dc90_121);
and \U$7414 ( \8203 , RIb54dc18_120, \7923 );
nor \U$7415 ( \8204 , \8202 , \8203 );
and \U$7416 ( \8205 , \7926 , RIb54e050_129);
nand \U$7417 ( \8206 , RIb54dba0_119, \7930 );
not \U$7418 ( \8207 , \8206 );
nor \U$7419 ( \8208 , \8205 , \8207 );
nand \U$7420 ( \8209 , \8198 , \8201 , \8204 , \8208 );
and \U$7421 ( \8210 , \7936 , RIb54e2a8_134);
and \U$7422 ( \8211 , RIb54e230_133, \7938 );
nor \U$7423 ( \8212 , \8210 , \8211 );
not \U$7424 ( \8213 , \8212 );
nor \U$7425 ( \8214 , \8195 , \8209 , \8213 );
and \U$7426 ( \8215 , \7943 , RIb54e140_131);
and \U$7427 ( \8216 , RIb54e1b8_132, \7945 );
nor \U$7428 ( \8217 , \8215 , \8216 );
and \U$7429 ( \8218 , \7948 , RIb54e320_135);
and \U$7430 ( \8219 , RIb54dd80_123, \7950 );
nor \U$7431 ( \8220 , \8218 , \8219 );
and \U$7432 ( \8221 , \7953 , RIb54de70_125);
and \U$7433 ( \8222 , RIb54e0c8_130, \7955 );
nor \U$7434 ( \8223 , \8221 , \8222 );
nand \U$7435 ( \8224 , \8214 , \8217 , \8220 , \8223 );
buf \U$7436 ( \8225 , \8224 );
_DC g2497 ( \8226_nG2497 , \8225 , \7963 );
xor \U$7437 ( \8227 , \8194 , \8226_nG2497 );
not \U$7438 ( \8228 , \7868 );
not \U$7439 ( \8229 , RIb55bb38_596);
and \U$7440 ( \8230 , \8228 , \8229 );
and \U$7441 ( \8231 , \7868 , RIb55bb38_596);
nor \U$7442 ( \8232 , \8230 , \8231 );
and \U$7443 ( \8233 , \7923 , RIb54e410_137);
and \U$7444 ( \8234 , RIb54e9b0_149, \7945 );
and \U$7445 ( \8235 , \7938 , RIb54ea28_150);
and \U$7446 ( \8236 , RIb54e5f0_141, \7900 );
nor \U$7447 ( \8237 , \8234 , \8235 , \8236 );
and \U$7448 ( \8238 , \7953 , RIb54e668_142);
and \U$7449 ( \8239 , RIb54e578_140, \7950 );
nor \U$7450 ( \8240 , \8238 , \8239 );
and \U$7451 ( \8241 , \7948 , RIb54eb18_152);
and \U$7452 ( \8242 , RIb54eaa0_151, \7936 );
nor \U$7453 ( \8243 , \8241 , \8242 );
and \U$7454 ( \8244 , \7943 , RIb54e938_148);
and \U$7455 ( \8245 , RIb54e8c0_147, \7955 );
nor \U$7456 ( \8246 , \8244 , \8245 );
nand \U$7457 ( \8247 , \8237 , \8240 , \8243 , \8246 );
nand \U$7458 ( \8248 , RIb54e398_136, \7930 );
not \U$7459 ( \8249 , \8248 );
nor \U$7460 ( \8250 , \8233 , \8247 , \8249 );
and \U$7461 ( \8251 , \7914 , RIb54e758_144);
and \U$7462 ( \8252 , RIb54e6e0_143, \7906 );
nor \U$7463 ( \8253 , \8251 , \8252 );
and \U$7464 ( \8254 , \7917 , RIb54e500_139);
and \U$7465 ( \8255 , RIb54e488_138, \7921 );
nor \U$7466 ( \8256 , \8254 , \8255 );
and \U$7467 ( \8257 , \7926 , RIb54e848_146);
and \U$7468 ( \8258 , RIb54e7d0_145, \7910 );
nor \U$7469 ( \8259 , \8257 , \8258 );
nand \U$7470 ( \8260 , \8250 , \8253 , \8256 , \8259 );
buf \U$7471 ( \8261 , \8260 );
_DC g2495 ( \8262_nG2495 , \8261 , \7963 );
xor \U$7472 ( \8263 , \8232 , \8262_nG2495 );
not \U$7473 ( \8264 , \7866 );
not \U$7474 ( \8265 , RIb55bbb0_597);
and \U$7475 ( \8266 , \8264 , \8265 );
and \U$7476 ( \8267 , \7866 , RIb55bbb0_597);
nor \U$7477 ( \8268 , \8266 , \8267 );
and \U$7478 ( \8269 , \7900 , RIb54ede8_158);
and \U$7479 ( \8270 , \7906 , RIb54eed8_160);
and \U$7480 ( \8271 , RIb54efc8_162, \7910 );
nor \U$7481 ( \8272 , \8270 , \8271 );
and \U$7482 ( \8273 , \7914 , RIb54ef50_161);
and \U$7483 ( \8274 , RIb54ecf8_156, \7917 );
nor \U$7484 ( \8275 , \8273 , \8274 );
and \U$7485 ( \8276 , \7921 , RIb54ec80_155);
and \U$7486 ( \8277 , RIb54ec08_154, \7923 );
nor \U$7487 ( \8278 , \8276 , \8277 );
and \U$7488 ( \8279 , \7926 , RIb54f040_163);
nand \U$7489 ( \8280 , RIb54eb90_153, \7930 );
not \U$7490 ( \8281 , \8280 );
nor \U$7491 ( \8282 , \8279 , \8281 );
nand \U$7492 ( \8283 , \8272 , \8275 , \8278 , \8282 );
and \U$7493 ( \8284 , \7936 , RIb54f298_168);
and \U$7494 ( \8285 , RIb54f220_167, \7938 );
nor \U$7495 ( \8286 , \8284 , \8285 );
not \U$7496 ( \8287 , \8286 );
nor \U$7497 ( \8288 , \8269 , \8283 , \8287 );
and \U$7498 ( \8289 , \7943 , RIb54f130_165);
and \U$7499 ( \8290 , RIb54f1a8_166, \7945 );
nor \U$7500 ( \8291 , \8289 , \8290 );
and \U$7501 ( \8292 , \7948 , RIb54f310_169);
and \U$7502 ( \8293 , RIb54ed70_157, \7950 );
nor \U$7503 ( \8294 , \8292 , \8293 );
and \U$7504 ( \8295 , \7953 , RIb54ee60_159);
and \U$7505 ( \8296 , RIb54f0b8_164, \7955 );
nor \U$7506 ( \8297 , \8295 , \8296 );
nand \U$7507 ( \8298 , \8288 , \8291 , \8294 , \8297 );
buf \U$7508 ( \8299 , \8298 );
_DC g23c0 ( \8300_nG23c0 , \8299 , \7963 );
xor \U$7509 ( \8301 , \8268 , \8300_nG23c0 );
xnor \U$7510 ( \8302 , RIb55bc28_598, RIb55bca0_599);
and \U$7511 ( \8303 , \7923 , RIb54f400_171);
and \U$7512 ( \8304 , RIb54f9a0_183, \7945 );
and \U$7513 ( \8305 , \7938 , RIb54fa18_184);
and \U$7514 ( \8306 , RIb54f5e0_175, \7900 );
nor \U$7515 ( \8307 , \8304 , \8305 , \8306 );
and \U$7516 ( \8308 , \7953 , RIb54f658_176);
and \U$7517 ( \8309 , RIb54f568_174, \7950 );
nor \U$7518 ( \8310 , \8308 , \8309 );
and \U$7519 ( \8311 , \7948 , RIb54fb08_186);
and \U$7520 ( \8312 , RIb54fa90_185, \7936 );
nor \U$7521 ( \8313 , \8311 , \8312 );
and \U$7522 ( \8314 , \7943 , RIb54f928_182);
and \U$7523 ( \8315 , RIb54f8b0_181, \7955 );
nor \U$7524 ( \8316 , \8314 , \8315 );
nand \U$7525 ( \8317 , \8307 , \8310 , \8313 , \8316 );
nand \U$7526 ( \8318 , RIb54f388_170, \7930 );
not \U$7527 ( \8319 , \8318 );
nor \U$7528 ( \8320 , \8303 , \8317 , \8319 );
and \U$7529 ( \8321 , \7914 , RIb54f748_178);
and \U$7530 ( \8322 , RIb54f6d0_177, \7906 );
nor \U$7531 ( \8323 , \8321 , \8322 );
and \U$7532 ( \8324 , \7917 , RIb54f4f0_173);
and \U$7533 ( \8325 , RIb54f478_172, \7921 );
nor \U$7534 ( \8326 , \8324 , \8325 );
and \U$7535 ( \8327 , \7926 , RIb54f838_180);
and \U$7536 ( \8328 , RIb54f7c0_179, \7910 );
nor \U$7537 ( \8329 , \8327 , \8328 );
nand \U$7538 ( \8330 , \8320 , \8323 , \8326 , \8329 );
buf \U$7539 ( \8331 , \8330 );
_DC g23c2 ( \8332_nG23c2 , \8331 , \7963 );
xor \U$7540 ( \8333 , \8302 , \8332_nG23c2 );
and \U$7541 ( \8334 , \7923 , RIb54fbf8_188);
and \U$7542 ( \8335 , RIb550198_200, \7945 );
and \U$7543 ( \8336 , \7938 , RIb550210_201);
and \U$7544 ( \8337 , RIb54fdd8_192, \7900 );
nor \U$7545 ( \8338 , \8335 , \8336 , \8337 );
and \U$7546 ( \8339 , \7953 , RIb54fe50_193);
and \U$7547 ( \8340 , RIb54fd60_191, \7950 );
nor \U$7548 ( \8341 , \8339 , \8340 );
and \U$7549 ( \8342 , \7948 , RIb550300_203);
and \U$7550 ( \8343 , RIb550288_202, \7936 );
nor \U$7551 ( \8344 , \8342 , \8343 );
and \U$7552 ( \8345 , \7943 , RIb550120_199);
and \U$7553 ( \8346 , RIb5500a8_198, \7955 );
nor \U$7554 ( \8347 , \8345 , \8346 );
nand \U$7555 ( \8348 , \8338 , \8341 , \8344 , \8347 );
nand \U$7556 ( \8349 , RIb54fb80_187, \7930 );
not \U$7557 ( \8350 , \8349 );
nor \U$7558 ( \8351 , \8334 , \8348 , \8350 );
and \U$7559 ( \8352 , \7914 , RIb54ff40_195);
and \U$7560 ( \8353 , RIb54fec8_194, \7906 );
nor \U$7561 ( \8354 , \8352 , \8353 );
and \U$7562 ( \8355 , \7917 , RIb54fce8_190);
and \U$7563 ( \8356 , RIb54fc70_189, \7921 );
nor \U$7564 ( \8357 , \8355 , \8356 );
and \U$7565 ( \8358 , \7926 , RIb550030_197);
and \U$7566 ( \8359 , RIb54ffb8_196, \7910 );
nor \U$7567 ( \8360 , \8358 , \8359 );
nand \U$7568 ( \8361 , \8351 , \8354 , \8357 , \8360 );
buf \U$7569 ( \8362 , \8361 );
_DC g2255 ( \8363_nG2255 , \8362 , \7963 );
xor \U$7570 ( \8364 , RIb55bca0_599, \8363_nG2255 );
and \U$7571 ( \8365 , \7923 , RIb550468_206);
and \U$7572 ( \8366 , RIb550a08_218, \7945 );
and \U$7573 ( \8367 , \7938 , RIb550a80_219);
and \U$7574 ( \8368 , RIb550648_210, \7900 );
nor \U$7575 ( \8369 , \8366 , \8367 , \8368 );
and \U$7576 ( \8370 , \7953 , RIb5506c0_211);
and \U$7577 ( \8371 , RIb5505d0_209, \7950 );
nor \U$7578 ( \8372 , \8370 , \8371 );
and \U$7579 ( \8373 , \7948 , RIb550b70_221);
and \U$7580 ( \8374 , RIb550af8_220, \7936 );
nor \U$7581 ( \8375 , \8373 , \8374 );
and \U$7582 ( \8376 , \7943 , RIb550990_217);
and \U$7583 ( \8377 , RIb550918_216, \7955 );
nor \U$7584 ( \8378 , \8376 , \8377 );
nand \U$7585 ( \8379 , \8369 , \8372 , \8375 , \8378 );
nand \U$7586 ( \8380 , RIb5503f0_205, \7930 );
not \U$7587 ( \8381 , \8380 );
nor \U$7588 ( \8382 , \8365 , \8379 , \8381 );
and \U$7589 ( \8383 , \7914 , RIb5507b0_213);
and \U$7590 ( \8384 , RIb550738_212, \7906 );
nor \U$7591 ( \8385 , \8383 , \8384 );
and \U$7592 ( \8386 , \7917 , RIb550558_208);
and \U$7593 ( \8387 , RIb5504e0_207, \7921 );
nor \U$7594 ( \8388 , \8386 , \8387 );
and \U$7595 ( \8389 , \7926 , RIb5508a0_215);
and \U$7596 ( \8390 , RIb550828_214, \7910 );
nor \U$7597 ( \8391 , \8389 , \8390 );
nand \U$7598 ( \8392 , \8382 , \8385 , \8388 , \8391 );
buf \U$7599 ( \8393 , \8392 );
_DC g2253 ( \8394_nG2253 , \8393 , \7963 );
not \U$7600 ( \8395 , RIb55bf70_605);
nand \U$7601 ( \8396 , \8394_nG2253 , \8395 );
not \U$7602 ( \8397 , \8396 );
and \U$7603 ( \8398 , \8364 , \8397 );
and \U$7604 ( \8399 , RIb55bca0_599, \8363_nG2255 );
or \U$7605 ( \8400 , \8398 , \8399 );
and \U$7606 ( \8401 , \8333 , \8400 );
and \U$7607 ( \8402 , \8302 , \8332_nG23c2 );
or \U$7608 ( \8403 , \8401 , \8402 );
and \U$7609 ( \8404 , \8301 , \8403 );
and \U$7610 ( \8405 , \8268 , \8300_nG23c0 );
or \U$7611 ( \8406 , \8404 , \8405 );
and \U$7612 ( \8407 , \8263 , \8406 );
and \U$7613 ( \8408 , \8232 , \8262_nG2495 );
or \U$7614 ( \8409 , \8407 , \8408 );
and \U$7615 ( \8410 , \8227 , \8409 );
and \U$7616 ( \8411 , \8194 , \8226_nG2497 );
or \U$7617 ( \8412 , \8410 , \8411 );
and \U$7618 ( \8413 , \8189 , \8412 );
and \U$7619 ( \8414 , \8156 , \8188_nG25c5 );
or \U$7620 ( \8415 , \8413 , \8414 );
and \U$7621 ( \8416 , \8151 , \8415 );
and \U$7622 ( \8417 , \8118 , \8150_nG25c7 );
or \U$7623 ( \8418 , \8416 , \8417 );
and \U$7624 ( \8419 , \8113 , \8418 );
and \U$7625 ( \8420 , \8082 , \8112_nG273b );
or \U$7626 ( \8421 , \8419 , \8420 );
and \U$7627 ( \8422 , \8077 , \8421 );
and \U$7628 ( \8423 , \8044 , \8076_nG273d );
or \U$7629 ( \8424 , \8422 , \8423 );
and \U$7630 ( \8425 , \8039 , \8424 );
and \U$7631 ( \8426 , \8006 , \8038_nG28f0 );
or \U$7632 ( \8427 , \8425 , \8426 );
and \U$7633 ( \8428 , \8001 , \8427 );
and \U$7634 ( \8429 , \7970 , \8000_nG28f2 );
or \U$7635 ( \8430 , \8428 , \8429 );
and \U$7636 ( \8431 , \7965 , \8430 );
and \U$7637 ( \8432 , \7889 , \7964_nG2ace );
or \U$7638 ( \8433 , \8431 , \8432 );
not \U$7639 ( \8434 , \7884 );
nand \U$7640 ( \8435 , \8434 , RIb55c3a8_614);
nor \U$7641 ( \8436 , \8433 , \8435 );
not \U$7642 ( \8437 , \8436 );
and \U$7643 ( \8438 , RIb551098_232, \7917 );
and \U$7644 ( \8439 , RIb5513e0_239, \7926 );
and \U$7645 ( \8440 , \7943 , RIb5514d0_241);
and \U$7646 ( \8441 , RIb551458_240, \7955 );
nor \U$7647 ( \8442 , \8440 , \8441 );
and \U$7648 ( \8443 , \7948 , RIb5516b0_245);
and \U$7649 ( \8444 , RIb551638_244, \7936 );
nor \U$7650 ( \8445 , \8443 , \8444 );
and \U$7651 ( \8446 , \7914 , RIb5512f0_237);
and \U$7652 ( \8447 , RIb551188_234, \7900 );
nor \U$7653 ( \8448 , \8446 , \8447 );
and \U$7654 ( \8449 , \7938 , RIb5515c0_243);
and \U$7655 ( \8450 , RIb551548_242, \7945 );
nor \U$7656 ( \8451 , \8449 , \8450 );
nand \U$7657 ( \8452 , \8442 , \8445 , \8448 , \8451 );
nor \U$7658 ( \8453 , \8438 , \8439 , \8452 );
and \U$7659 ( \8454 , \7910 , RIb551368_238);
and \U$7660 ( \8455 , RIb551020_231, \7921 );
nor \U$7661 ( \8456 , \8454 , \8455 );
and \U$7662 ( \8457 , \7953 , RIb551200_235);
and \U$7663 ( \8458 , RIb551110_233, \7950 );
nor \U$7664 ( \8459 , \8457 , \8458 );
not \U$7665 ( \8460 , \7923 );
not \U$7666 ( \8461 , \7930 );
nand \U$7667 ( \8462 , \8460 , \8461 );
and \U$7668 ( \8463 , \8462 , RIb550be8_222);
and \U$7669 ( \8464 , RIb551278_236, \7906 );
nor \U$7670 ( \8465 , \8463 , \8464 );
nand \U$7671 ( \8466 , \8453 , \8456 , \8459 , \8465 );
buf \U$7672 ( \8467 , \7962 );
_DC g310a ( \8468_nG310a , \8466 , \8467 );
not \U$7673 ( \8469 , \8468_nG310a );
nor \U$7674 ( \8470 , \8437 , \8469 );
xor \U$7675 ( \8471 , \7889 , \7964_nG2ace );
xor \U$7676 ( \8472 , \8471 , \8430 );
not \U$7677 ( \8473 , \8472 );
xor \U$7678 ( \8474 , \7970 , \8000_nG28f2 );
xor \U$7679 ( \8475 , \8474 , \8427 );
not \U$7680 ( \8476 , \8475 );
and \U$7681 ( \8477 , \8473 , \8476 );
and \U$7682 ( \8478 , \8433 , \8435 );
nor \U$7683 ( \8479 , \8478 , \8436 );
nor \U$7684 ( \8480 , \8477 , \8479 );
not \U$7685 ( \8481 , \8480 );
and \U$7686 ( \8482 , RIb552010_265, \8462 );
and \U$7687 ( \8483 , RIb552100_267, \7917 );
and \U$7688 ( \8484 , \7955 , RIb5524c0_275);
and \U$7689 ( \8485 , RIb552448_274, \7926 );
nor \U$7690 ( \8486 , \8484 , \8485 );
and \U$7691 ( \8487 , \7948 , RIb552718_280);
and \U$7692 ( \8488 , RIb5523d0_273, \7910 );
nor \U$7693 ( \8489 , \8487 , \8488 );
and \U$7694 ( \8490 , \7906 , RIb5522e0_271);
and \U$7695 ( \8491 , RIb5521f0_269, \7900 );
nor \U$7696 ( \8492 , \8490 , \8491 );
and \U$7697 ( \8493 , \7936 , RIb5526a0_279);
and \U$7698 ( \8494 , RIb552628_278, \7938 );
nor \U$7699 ( \8495 , \8493 , \8494 );
nand \U$7700 ( \8496 , \8486 , \8489 , \8492 , \8495 );
nor \U$7701 ( \8497 , \8482 , \8483 , \8496 );
and \U$7702 ( \8498 , \7945 , RIb5525b0_277);
and \U$7703 ( \8499 , RIb552178_268, \7950 );
nor \U$7704 ( \8500 , \8498 , \8499 );
and \U$7705 ( \8501 , \7953 , RIb552268_270);
and \U$7706 ( \8502 , RIb552088_266, \7921 );
nor \U$7707 ( \8503 , \8501 , \8502 );
and \U$7708 ( \8504 , \7914 , RIb552358_272);
and \U$7709 ( \8505 , RIb552538_276, \7943 );
nor \U$7710 ( \8506 , \8504 , \8505 );
nand \U$7711 ( \8507 , \8497 , \8500 , \8503 , \8506 );
_DC g3222 ( \8508_nG3222 , \8507 , \8467 );
or \U$7712 ( \8509 , \8481 , \8508_nG3222 );
not \U$7713 ( \8510 , \8508_nG3222 );
and \U$7714 ( \8511 , \8479 , \8472 );
nor \U$7715 ( \8512 , \8479 , \8472 );
xnor \U$7716 ( \8513 , \8475 , \8472 );
not \U$7717 ( \8514 , \8513 );
nor \U$7718 ( \8515 , \8511 , \8512 , \8514 );
nand \U$7719 ( \8516 , \8481 , \8515 );
or \U$7720 ( \8517 , \8510 , \8516 );
or \U$7721 ( \8518 , \8481 , \8515 );
nand \U$7722 ( \8519 , \8509 , \8517 , \8518 );
xnor \U$7723 ( \8520 , \8470 , \8519 );
nor \U$7724 ( \8521 , \8480 , \8513 );
not \U$7725 ( \8522 , \8521 );
or \U$7726 ( \8523 , \8522 , \8510 );
or \U$7727 ( \8524 , \8469 , \8516 );
or \U$7728 ( \8525 , \8513 , \8510 );
or \U$7729 ( \8526 , \8481 , \8468_nG310a );
nand \U$7730 ( \8527 , \8526 , \8518 );
nand \U$7731 ( \8528 , \8525 , \8527 );
nand \U$7732 ( \8529 , \8523 , \8524 , \8528 );
xor \U$7733 ( \8530 , \8006 , \8038_nG28f0 );
xor \U$7734 ( \8531 , \8530 , \8424 );
xor \U$7735 ( \8532 , \8044 , \8076_nG273d );
xor \U$7736 ( \8533 , \8532 , \8421 );
nor \U$7737 ( \8534 , \8531 , \8533 );
or \U$7738 ( \8535 , \8475 , \8534 );
and \U$7739 ( \8536 , \8529 , \8535 );
and \U$7740 ( \8537 , RIb5529e8_286, \7900 );
and \U$7741 ( \8538 , RIb552e98_296, \7936 );
and \U$7742 ( \8539 , \7943 , RIb552d30_293);
and \U$7743 ( \8540 , RIb552da8_294, \7945 );
nor \U$7744 ( \8541 , \8539 , \8540 );
and \U$7745 ( \8542 , \7953 , RIb552a60_287);
and \U$7746 ( \8543 , RIb552970_285, \7950 );
nor \U$7747 ( \8544 , \8542 , \8543 );
and \U$7748 ( \8545 , \7917 , RIb5528f8_284);
and \U$7749 ( \8546 , RIb552880_283, \7921 );
nor \U$7750 ( \8547 , \8545 , \8546 );
and \U$7751 ( \8548 , \8462 , RIb552808_282);
and \U$7752 ( \8549 , RIb552b50_289, \7914 );
nor \U$7753 ( \8550 , \8548 , \8549 );
nand \U$7754 ( \8551 , \8541 , \8544 , \8547 , \8550 );
nor \U$7755 ( \8552 , \8537 , \8538 , \8551 );
and \U$7756 ( \8553 , \7938 , RIb552e20_295);
and \U$7757 ( \8554 , RIb552bc8_290, \7910 );
nor \U$7758 ( \8555 , \8553 , \8554 );
and \U$7759 ( \8556 , \7948 , RIb552f10_297);
and \U$7760 ( \8557 , RIb552ad8_288, \7906 );
nor \U$7761 ( \8558 , \8556 , \8557 );
and \U$7762 ( \8559 , \7955 , RIb552cb8_292);
and \U$7763 ( \8560 , RIb552c40_291, \7926 );
nor \U$7764 ( \8561 , \8559 , \8560 );
nand \U$7765 ( \8562 , \8552 , \8555 , \8558 , \8561 );
_DC g3003 ( \8563_nG3003 , \8562 , \8467 );
not \U$7766 ( \8564 , \8563_nG3003 );
nor \U$7767 ( \8565 , \8437 , \8564 );
nor \U$7768 ( \8566 , \8536 , \8565 );
xor \U$7769 ( \8567 , \8520 , \8566 );
not \U$7770 ( \8568 , \8567 );
not \U$7771 ( \8569 , \8531 );
not \U$7772 ( \8570 , \8475 );
or \U$7773 ( \8571 , \8569 , \8570 );
or \U$7774 ( \8572 , \8475 , \8531 );
nand \U$7775 ( \8573 , \8571 , \8572 );
xor \U$7776 ( \8574 , \8533 , \8531 );
nor \U$7777 ( \8575 , \8573 , \8574 );
not \U$7778 ( \8576 , \8575 );
not \U$7779 ( \8577 , \8535 );
nor \U$7780 ( \8578 , \8576 , \8577 );
not \U$7781 ( \8579 , \8578 );
or \U$7782 ( \8580 , \8579 , \8510 );
or \U$7783 ( \8581 , \8576 , \8510 );
nand \U$7784 ( \8582 , \8581 , \8577 );
nand \U$7785 ( \8583 , \8580 , \8582 );
or \U$7786 ( \8584 , \8522 , \8469 );
or \U$7787 ( \8585 , \8564 , \8516 );
or \U$7788 ( \8586 , \8513 , \8469 );
or \U$7789 ( \8587 , \8481 , \8563_nG3003 );
nand \U$7790 ( \8588 , \8587 , \8518 );
nand \U$7791 ( \8589 , \8586 , \8588 );
nand \U$7792 ( \8590 , \8584 , \8585 , \8589 );
and \U$7793 ( \8591 , \8583 , \8590 );
not \U$7794 ( \8592 , \8591 );
and \U$7795 ( \8593 , \8529 , \8535 );
not \U$7796 ( \8594 , \8529 );
and \U$7797 ( \8595 , \8594 , \8577 );
nor \U$7798 ( \8596 , \8593 , \8595 );
xnor \U$7799 ( \8597 , \8596 , \8565 );
nor \U$7800 ( \8598 , \8592 , \8597 );
and \U$7801 ( \8599 , \8568 , \8598 );
or \U$7802 ( \8600 , \8599 , \8480 );
and \U$7803 ( \8601 , \8519 , \8470 );
and \U$7804 ( \8602 , \8480 , \8599 );
nor \U$7805 ( \8603 , \8601 , \8602 );
nand \U$7806 ( \8604 , \8600 , \8603 );
not \U$7807 ( \8605 , \8604 );
and \U$7808 ( \8606 , \8436 , \8508_nG3222 );
and \U$7809 ( \8607 , \8520 , \8566 );
nor \U$7810 ( \8608 , \8606 , \8607 );
not \U$7811 ( \8609 , \8608 );
and \U$7812 ( \8610 , \8605 , \8609 );
and \U$7813 ( \8611 , \8604 , \8608 );
nor \U$7814 ( \8612 , \8610 , \8611 );
not \U$7815 ( \8613 , \8612 );
xor \U$7816 ( \8614 , \8568 , \8598 );
not \U$7817 ( \8615 , \8614 );
not \U$7818 ( \8616 , \8597 );
not \U$7819 ( \8617 , \8591 );
and \U$7820 ( \8618 , \8616 , \8617 );
and \U$7821 ( \8619 , \8597 , \8591 );
nor \U$7822 ( \8620 , \8618 , \8619 );
not \U$7823 ( \8621 , \8620 );
and \U$7824 ( \8622 , \8468_nG310a , \8578 );
and \U$7825 ( \8623 , \8535 , \8574 );
and \U$7826 ( \8624 , \8623 , \8508_nG3222 );
nand \U$7827 ( \8625 , \8468_nG310a , \8575 );
or \U$7828 ( \8626 , \8535 , \8508_nG3222 );
or \U$7829 ( \8627 , \8535 , \8574 );
nand \U$7830 ( \8628 , \8626 , \8627 );
and \U$7831 ( \8629 , \8625 , \8628 );
nor \U$7832 ( \8630 , \8622 , \8624 , \8629 );
and \U$7833 ( \8631 , \8563_nG3003 , \8521 );
and \U$7834 ( \8632 , RIb5539d8_320, \7900 );
and \U$7835 ( \8633 , RIb553ca8_326, \7955 );
and \U$7836 ( \8634 , \7943 , RIb553d20_327);
and \U$7837 ( \8635 , RIb553d98_328, \7945 );
nor \U$7838 ( \8636 , \8634 , \8635 );
and \U$7839 ( \8637 , \7950 , RIb553960_319);
and \U$7840 ( \8638 , RIb553bb8_324, \7910 );
nor \U$7841 ( \8639 , \8637 , \8638 );
and \U$7842 ( \8640 , \7917 , RIb5538e8_318);
and \U$7843 ( \8641 , RIb553870_317, \7921 );
nor \U$7844 ( \8642 , \8640 , \8641 );
and \U$7845 ( \8643 , \8462 , RIb5537f8_316);
and \U$7846 ( \8644 , RIb553b40_323, \7914 );
nor \U$7847 ( \8645 , \8643 , \8644 );
nand \U$7848 ( \8646 , \8636 , \8639 , \8642 , \8645 );
nor \U$7849 ( \8647 , \8632 , \8633 , \8646 );
and \U$7850 ( \8648 , \7936 , RIb553e88_330);
and \U$7851 ( \8649 , RIb553c30_325, \7926 );
nor \U$7852 ( \8650 , \8648 , \8649 );
and \U$7853 ( \8651 , \7948 , RIb553f00_331);
and \U$7854 ( \8652 , RIb553e10_329, \7938 );
nor \U$7855 ( \8653 , \8651 , \8652 );
and \U$7856 ( \8654 , \7906 , RIb553ac8_322);
and \U$7857 ( \8655 , RIb553a50_321, \7953 );
nor \U$7858 ( \8656 , \8654 , \8655 );
nand \U$7859 ( \8657 , \8647 , \8650 , \8653 , \8656 );
_DC g2ee1 ( \8658_nG2ee1 , \8657 , \8467 );
or \U$7860 ( \8659 , \8481 , \8658_nG2ee1 );
nand \U$7861 ( \8660 , \8659 , \8518 );
nand \U$7862 ( \8661 , \8563_nG3003 , \8514 );
and \U$7863 ( \8662 , \8660 , \8661 );
not \U$7864 ( \8663 , \8516 );
and \U$7865 ( \8664 , \8658_nG2ee1 , \8663 );
nor \U$7866 ( \8665 , \8631 , \8662 , \8664 );
nand \U$7867 ( \8666 , \8630 , \8665 );
xor \U$7868 ( \8667 , \8082 , \8112_nG273b );
xor \U$7869 ( \8668 , \8667 , \8418 );
xor \U$7870 ( \8669 , \8118 , \8150_nG25c7 );
xor \U$7871 ( \8670 , \8669 , \8415 );
nor \U$7872 ( \8671 , \8668 , \8670 );
or \U$7873 ( \8672 , \8533 , \8671 );
and \U$7874 ( \8673 , \8666 , \8672 );
nor \U$7875 ( \8674 , \8665 , \8630 );
nor \U$7876 ( \8675 , \8673 , \8674 );
xor \U$7877 ( \8676 , \8583 , \8590 );
not \U$7878 ( \8677 , \8676 );
nand \U$7879 ( \8678 , \8658_nG2ee1 , \8436 );
not \U$7880 ( \8679 , \8678 );
and \U$7881 ( \8680 , \8677 , \8679 );
and \U$7882 ( \8681 , \8676 , \8678 );
nor \U$7883 ( \8682 , \8680 , \8681 );
nand \U$7884 ( \8683 , \8675 , \8682 );
nand \U$7885 ( \8684 , \8621 , \8683 );
nor \U$7886 ( \8685 , \8615 , \8684 );
not \U$7887 ( \8686 , \8685 );
and \U$7888 ( \8687 , \8613 , \8686 );
and \U$7889 ( \8688 , \8612 , \8685 );
nor \U$7890 ( \8689 , \8687 , \8688 );
not \U$7891 ( \8690 , \8689 );
not \U$7892 ( \8691 , \8620 );
not \U$7893 ( \8692 , \8683 );
and \U$7894 ( \8693 , \8691 , \8692 );
and \U$7895 ( \8694 , \8620 , \8683 );
nor \U$7896 ( \8695 , \8693 , \8694 );
not \U$7897 ( \8696 , \8672 );
not \U$7898 ( \8697 , \8674 );
nand \U$7899 ( \8698 , \8697 , \8666 );
not \U$7900 ( \8699 , \8698 );
or \U$7901 ( \8700 , \8696 , \8699 );
or \U$7902 ( \8701 , \8698 , \8672 );
nand \U$7903 ( \8702 , \8700 , \8701 );
not \U$7904 ( \8703 , \8702 );
and \U$7905 ( \8704 , RIb5531e0_303, \7900 );
and \U$7906 ( \8705 , RIb553690_313, \7936 );
and \U$7907 ( \8706 , \7943 , RIb553528_310);
and \U$7908 ( \8707 , RIb5535a0_311, \7945 );
nor \U$7909 ( \8708 , \8706 , \8707 );
and \U$7910 ( \8709 , \7953 , RIb553258_304);
and \U$7911 ( \8710 , RIb553168_302, \7950 );
nor \U$7912 ( \8711 , \8709 , \8710 );
and \U$7913 ( \8712 , \7917 , RIb5530f0_301);
and \U$7914 ( \8713 , RIb553078_300, \7921 );
nor \U$7915 ( \8714 , \8712 , \8713 );
and \U$7916 ( \8715 , \8462 , RIb553000_299);
and \U$7917 ( \8716 , RIb553348_306, \7914 );
nor \U$7918 ( \8717 , \8715 , \8716 );
nand \U$7919 ( \8718 , \8708 , \8711 , \8714 , \8717 );
nor \U$7920 ( \8719 , \8704 , \8705 , \8718 );
and \U$7921 ( \8720 , \7938 , RIb553618_312);
and \U$7922 ( \8721 , RIb5534b0_309, \7955 );
nor \U$7923 ( \8722 , \8720 , \8721 );
and \U$7924 ( \8723 , \7948 , RIb553708_314);
and \U$7925 ( \8724 , RIb553438_308, \7926 );
nor \U$7926 ( \8725 , \8723 , \8724 );
and \U$7927 ( \8726 , \7906 , RIb5532d0_305);
and \U$7928 ( \8727 , RIb5533c0_307, \7910 );
nor \U$7929 ( \8728 , \8726 , \8727 );
nand \U$7930 ( \8729 , \8719 , \8722 , \8725 , \8728 );
_DC g2df7 ( \8730_nG2df7 , \8729 , \8467 );
nand \U$7931 ( \8731 , \8730_nG2df7 , \8436 );
not \U$7932 ( \8732 , \8731 );
and \U$7933 ( \8733 , \8703 , \8732 );
and \U$7934 ( \8734 , \8702 , \8731 );
nor \U$7935 ( \8735 , \8733 , \8734 );
not \U$7936 ( \8736 , \8735 );
and \U$7937 ( \8737 , \8658_nG2ee1 , \8521 );
or \U$7938 ( \8738 , \8481 , \8730_nG2df7 );
nand \U$7939 ( \8739 , \8738 , \8518 );
nand \U$7940 ( \8740 , \8658_nG2ee1 , \8514 );
and \U$7941 ( \8741 , \8739 , \8740 );
and \U$7942 ( \8742 , \8730_nG2df7 , \8663 );
nor \U$7943 ( \8743 , \8737 , \8741 , \8742 );
and \U$7944 ( \8744 , RIb5541d0_337, \7900 );
and \U$7945 ( \8745 , RIb5544a0_343, \7955 );
and \U$7946 ( \8746 , \7943 , RIb554518_344);
and \U$7947 ( \8747 , RIb554590_345, \7945 );
nor \U$7948 ( \8748 , \8746 , \8747 );
and \U$7949 ( \8749 , \7914 , RIb554338_340);
and \U$7950 ( \8750 , RIb5540e0_335, \7917 );
nor \U$7951 ( \8751 , \8749 , \8750 );
and \U$7952 ( \8752 , \7953 , RIb554248_338);
and \U$7953 ( \8753 , RIb554158_336, \7950 );
nor \U$7954 ( \8754 , \8752 , \8753 );
and \U$7955 ( \8755 , \8462 , RIb553ff0_333);
and \U$7956 ( \8756 , RIb554068_334, \7921 );
nor \U$7957 ( \8757 , \8755 , \8756 );
nand \U$7958 ( \8758 , \8748 , \8751 , \8754 , \8757 );
nor \U$7959 ( \8759 , \8744 , \8745 , \8758 );
and \U$7960 ( \8760 , \7936 , RIb554680_347);
and \U$7961 ( \8761 , RIb554608_346, \7938 );
nor \U$7962 ( \8762 , \8760 , \8761 );
and \U$7963 ( \8763 , \7948 , RIb5546f8_348);
and \U$7964 ( \8764 , RIb5542c0_339, \7906 );
nor \U$7965 ( \8765 , \8763 , \8764 );
and \U$7966 ( \8766 , \7926 , RIb554428_342);
and \U$7967 ( \8767 , RIb5543b0_341, \7910 );
nor \U$7968 ( \8768 , \8766 , \8767 );
nand \U$7969 ( \8769 , \8759 , \8762 , \8765 , \8768 );
_DC g2cf7 ( \8770_nG2cf7 , \8769 , \8467 );
nand \U$7970 ( \8771 , \8770_nG2cf7 , \8436 );
or \U$7971 ( \8772 , \8743 , \8771 );
and \U$7972 ( \8773 , \8533 , \8668 );
nor \U$7973 ( \8774 , \8533 , \8668 );
xor \U$7974 ( \8775 , \8668 , \8670 );
nor \U$7975 ( \8776 , \8773 , \8774 , \8775 );
and \U$7976 ( \8777 , \8776 , \8672 );
and \U$7977 ( \8778 , \8508_nG3222 , \8777 );
not \U$7978 ( \8779 , \8672 );
and \U$7979 ( \8780 , \8510 , \8779 );
or \U$7980 ( \8781 , \8776 , \8672 );
not \U$7981 ( \8782 , \8781 );
nor \U$7982 ( \8783 , \8778 , \8780 , \8782 );
and \U$7983 ( \8784 , \8563_nG3003 , \8578 );
and \U$7984 ( \8785 , \8623 , \8468_nG310a );
nand \U$7985 ( \8786 , \8563_nG3003 , \8575 );
or \U$7986 ( \8787 , \8535 , \8468_nG310a );
nand \U$7987 ( \8788 , \8787 , \8627 );
and \U$7988 ( \8789 , \8786 , \8788 );
nor \U$7989 ( \8790 , \8784 , \8785 , \8789 );
or \U$7990 ( \8791 , \8783 , \8790 );
nand \U$7991 ( \8792 , \8772 , \8791 );
nand \U$7992 ( \8793 , \8736 , \8792 );
not \U$7993 ( \8794 , \8793 );
or \U$7994 ( \8795 , \8682 , \8675 );
nand \U$7995 ( \8796 , \8795 , \8683 );
nand \U$7996 ( \8797 , \8794 , \8796 );
nand \U$7997 ( \8798 , \8695 , \8797 );
not \U$7998 ( \8799 , \8798 );
nor \U$7999 ( \8800 , \8797 , \8695 );
nor \U$8000 ( \8801 , \8799 , \8800 );
not \U$8001 ( \8802 , \8801 );
not \U$8002 ( \8803 , \8676 );
nor \U$8003 ( \8804 , \8803 , \8678 );
not \U$8004 ( \8805 , \8804 );
and \U$8005 ( \8806 , \8802 , \8805 );
and \U$8006 ( \8807 , \8801 , \8804 );
nor \U$8007 ( \8808 , \8806 , \8807 );
not \U$8008 ( \8809 , \8702 );
nor \U$8009 ( \8810 , \8809 , \8731 );
not \U$8010 ( \8811 , \8796 );
not \U$8011 ( \8812 , \8793 );
or \U$8012 ( \8813 , \8811 , \8812 );
or \U$8013 ( \8814 , \8793 , \8796 );
nand \U$8014 ( \8815 , \8813 , \8814 );
nand \U$8015 ( \8816 , \8810 , \8815 );
xnor \U$8016 ( \8817 , \8783 , \8790 );
not \U$8017 ( \8818 , \8817 );
xor \U$8018 ( \8819 , \8771 , \8743 );
not \U$8019 ( \8820 , \8819 );
or \U$8020 ( \8821 , \8818 , \8820 );
or \U$8021 ( \8822 , \8819 , \8817 );
nand \U$8022 ( \8823 , \8821 , \8822 );
and \U$8023 ( \8824 , \8730_nG2df7 , \8521 );
or \U$8024 ( \8825 , \8481 , \8770_nG2cf7 );
nand \U$8025 ( \8826 , \8825 , \8518 );
nand \U$8026 ( \8827 , \8730_nG2df7 , \8514 );
and \U$8027 ( \8828 , \8826 , \8827 );
and \U$8028 ( \8829 , \8770_nG2cf7 , \8663 );
nor \U$8029 ( \8830 , \8824 , \8828 , \8829 );
and \U$8030 ( \8831 , RIb555058_368, \7921 );
and \U$8031 ( \8832 , RIb555328_374, \7914 );
and \U$8032 ( \8833 , \7955 , RIb555490_377);
and \U$8033 ( \8834 , RIb5553a0_375, \7910 );
nor \U$8034 ( \8835 , \8833 , \8834 );
and \U$8035 ( \8836 , \7938 , RIb5555f8_380);
and \U$8036 ( \8837 , RIb5551c0_371, \7900 );
nor \U$8037 ( \8838 , \8836 , \8837 );
and \U$8038 ( \8839 , \7948 , RIb5556e8_382);
and \U$8039 ( \8840 , RIb555670_381, \7936 );
nor \U$8040 ( \8841 , \8839 , \8840 );
and \U$8041 ( \8842 , \7906 , RIb5552b0_373);
and \U$8042 ( \8843 , RIb555418_376, \7926 );
nor \U$8043 ( \8844 , \8842 , \8843 );
nand \U$8044 ( \8845 , \8835 , \8838 , \8841 , \8844 );
nor \U$8045 ( \8846 , \8831 , \8832 , \8845 );
and \U$8046 ( \8847 , \7943 , RIb555508_378);
and \U$8047 ( \8848 , RIb555238_372, \7953 );
nor \U$8048 ( \8849 , \8847 , \8848 );
and \U$8049 ( \8850 , \7950 , RIb555148_370);
and \U$8050 ( \8851 , RIb5550d0_369, \7917 );
nor \U$8051 ( \8852 , \8850 , \8851 );
and \U$8052 ( \8853 , \8462 , RIb554fe0_367);
and \U$8053 ( \8854 , RIb555580_379, \7945 );
nor \U$8054 ( \8855 , \8853 , \8854 );
nand \U$8055 ( \8856 , \8846 , \8849 , \8852 , \8855 );
_DC g2bf3 ( \8857_nG2bf3 , \8856 , \8467 );
nand \U$8056 ( \8858 , \8857_nG2bf3 , \8436 );
or \U$8057 ( \8859 , \8830 , \8858 );
nand \U$8058 ( \8860 , \8508_nG3222 , \8775 );
or \U$8059 ( \8861 , \8672 , \8468_nG310a );
nand \U$8060 ( \8862 , \8861 , \8781 );
and \U$8061 ( \8863 , \8860 , \8862 );
and \U$8062 ( \8864 , \8777 , \8468_nG310a );
not \U$8063 ( \8865 , \8775 );
nor \U$8064 ( \8866 , \8779 , \8865 );
and \U$8065 ( \8867 , \8508_nG3222 , \8866 );
nor \U$8066 ( \8868 , \8863 , \8864 , \8867 );
not \U$8067 ( \8869 , \8868 );
xor \U$8068 ( \8870 , \8156 , \8188_nG25c5 );
xor \U$8069 ( \8871 , \8870 , \8412 );
xor \U$8070 ( \8872 , \8194 , \8226_nG2497 );
xor \U$8071 ( \8873 , \8872 , \8409 );
nor \U$8072 ( \8874 , \8871 , \8873 );
or \U$8073 ( \8875 , \8670 , \8874 );
not \U$8074 ( \8876 , \8875 );
not \U$8075 ( \8877 , \8876 );
and \U$8076 ( \8878 , \8869 , \8877 );
and \U$8077 ( \8879 , \8868 , \8876 );
and \U$8078 ( \8880 , \8658_nG2ee1 , \8578 );
and \U$8079 ( \8881 , \8623 , \8563_nG3003 );
nand \U$8080 ( \8882 , \8658_nG2ee1 , \8575 );
or \U$8081 ( \8883 , \8535 , \8563_nG3003 );
nand \U$8082 ( \8884 , \8883 , \8627 );
and \U$8083 ( \8885 , \8882 , \8884 );
nor \U$8084 ( \8886 , \8880 , \8881 , \8885 );
nor \U$8085 ( \8887 , \8879 , \8886 );
nor \U$8086 ( \8888 , \8878 , \8887 );
nand \U$8087 ( \8889 , \8859 , \8888 );
nor \U$8088 ( \8890 , \8823 , \8889 );
and \U$8089 ( \8891 , \8730_nG2df7 , \8578 );
and \U$8090 ( \8892 , \8623 , \8658_nG2ee1 );
nand \U$8091 ( \8893 , \8730_nG2df7 , \8575 );
or \U$8092 ( \8894 , \8535 , \8658_nG2ee1 );
nand \U$8093 ( \8895 , \8894 , \8627 );
and \U$8094 ( \8896 , \8893 , \8895 );
nor \U$8095 ( \8897 , \8891 , \8892 , \8896 );
and \U$8096 ( \8898 , RIb554860_351, \7921 );
and \U$8097 ( \8899 , RIb554c20_359, \7926 );
and \U$8098 ( \8900 , \7945 , RIb554d88_362);
and \U$8099 ( \8901 , RIb554ab8_356, \7906 );
nor \U$8100 ( \8902 , \8900 , \8901 );
and \U$8101 ( \8903 , \7955 , RIb554c98_360);
and \U$8102 ( \8904 , RIb5549c8_354, \7900 );
nor \U$8103 ( \8905 , \8903 , \8904 );
and \U$8104 ( \8906 , \7953 , RIb554a40_355);
and \U$8105 ( \8907 , RIb554950_353, \7950 );
nor \U$8106 ( \8908 , \8906 , \8907 );
and \U$8107 ( \8909 , \7948 , RIb554ef0_365);
and \U$8108 ( \8910 , RIb554d10_361, \7943 );
nor \U$8109 ( \8911 , \8909 , \8910 );
nand \U$8110 ( \8912 , \8902 , \8905 , \8908 , \8911 );
nor \U$8111 ( \8913 , \8898 , \8899 , \8912 );
and \U$8112 ( \8914 , \7914 , RIb554b30_357);
and \U$8113 ( \8915 , RIb554ba8_358, \7910 );
nor \U$8114 ( \8916 , \8914 , \8915 );
and \U$8115 ( \8917 , \7938 , RIb554e00_363);
and \U$8116 ( \8918 , RIb5548d8_352, \7917 );
nor \U$8117 ( \8919 , \8917 , \8918 );
and \U$8118 ( \8920 , \8462 , RIb5547e8_350);
and \U$8119 ( \8921 , RIb554e78_364, \7936 );
nor \U$8120 ( \8922 , \8920 , \8921 );
nand \U$8121 ( \8923 , \8913 , \8916 , \8919 , \8922 );
_DC g2ae9 ( \8924_nG2ae9 , \8923 , \8467 );
nand \U$8122 ( \8925 , \8924_nG2ae9 , \8436 );
xor \U$8123 ( \8926 , \8897 , \8925 );
and \U$8124 ( \8927 , \8770_nG2cf7 , \8521 );
or \U$8125 ( \8928 , \8481 , \8857_nG2bf3 );
nand \U$8126 ( \8929 , \8928 , \8518 );
nand \U$8127 ( \8930 , \8770_nG2cf7 , \8514 );
and \U$8128 ( \8931 , \8929 , \8930 );
and \U$8129 ( \8932 , \8857_nG2bf3 , \8663 );
nor \U$8130 ( \8933 , \8927 , \8931 , \8932 );
and \U$8131 ( \8934 , \8926 , \8933 );
and \U$8132 ( \8935 , \8897 , \8925 );
or \U$8133 ( \8936 , \8934 , \8935 );
not \U$8134 ( \8937 , \8936 );
not \U$8135 ( \8938 , \8871 );
not \U$8136 ( \8939 , \8670 );
or \U$8137 ( \8940 , \8938 , \8939 );
or \U$8138 ( \8941 , \8670 , \8871 );
nand \U$8139 ( \8942 , \8940 , \8941 );
xor \U$8140 ( \8943 , \8873 , \8871 );
nor \U$8141 ( \8944 , \8942 , \8943 );
nand \U$8142 ( \8945 , \8875 , \8944 );
or \U$8143 ( \8946 , \8945 , \8510 );
not \U$8144 ( \8947 , \8944 );
or \U$8145 ( \8948 , \8947 , \8510 );
nand \U$8146 ( \8949 , \8948 , \8876 );
nand \U$8147 ( \8950 , \8946 , \8949 );
not \U$8148 ( \8951 , \8866 );
or \U$8149 ( \8952 , \8951 , \8469 );
not \U$8150 ( \8953 , \8777 );
or \U$8151 ( \8954 , \8564 , \8953 );
or \U$8152 ( \8955 , \8865 , \8469 );
or \U$8153 ( \8956 , \8672 , \8563_nG3003 );
nand \U$8154 ( \8957 , \8956 , \8781 );
nand \U$8155 ( \8958 , \8955 , \8957 );
nand \U$8156 ( \8959 , \8952 , \8954 , \8958 );
and \U$8157 ( \8960 , \8950 , \8959 );
nand \U$8158 ( \8961 , \8937 , \8960 );
not \U$8159 ( \8962 , \8961 );
not \U$8160 ( \8963 , \8868 );
or \U$8161 ( \8964 , \8886 , \8875 );
nand \U$8162 ( \8965 , \8875 , \8886 );
nand \U$8163 ( \8966 , \8964 , \8965 );
not \U$8164 ( \8967 , \8966 );
or \U$8165 ( \8968 , \8963 , \8967 );
or \U$8166 ( \8969 , \8966 , \8868 );
nand \U$8167 ( \8970 , \8968 , \8969 );
xor \U$8168 ( \8971 , \8858 , \8830 );
and \U$8169 ( \8972 , \8970 , \8971 );
nand \U$8170 ( \8973 , \8962 , \8972 );
xor \U$8171 ( \8974 , \8890 , \8973 );
not \U$8172 ( \8975 , \8735 );
not \U$8173 ( \8976 , \8792 );
and \U$8174 ( \8977 , \8975 , \8976 );
and \U$8175 ( \8978 , \8735 , \8792 );
nor \U$8176 ( \8979 , \8977 , \8978 );
and \U$8177 ( \8980 , \8974 , \8979 );
and \U$8178 ( \8981 , \8890 , \8973 );
or \U$8179 ( \8982 , \8980 , \8981 );
and \U$8180 ( \8983 , \8816 , \8982 );
nor \U$8181 ( \8984 , \8815 , \8810 );
nor \U$8182 ( \8985 , \8983 , \8984 );
xor \U$8183 ( \8986 , \8808 , \8985 );
xor \U$8184 ( \8987 , \8897 , \8925 );
xor \U$8185 ( \8988 , \8987 , \8933 );
not \U$8186 ( \8989 , \8988 );
xor \U$8187 ( \8990 , \8950 , \8959 );
nand \U$8188 ( \8991 , \8989 , \8990 );
not \U$8189 ( \8992 , \8991 );
and \U$8190 ( \8993 , \8857_nG2bf3 , \8521 );
or \U$8191 ( \8994 , \8481 , \8924_nG2ae9 );
nand \U$8192 ( \8995 , \8994 , \8518 );
nand \U$8193 ( \8996 , \8857_nG2bf3 , \8514 );
and \U$8194 ( \8997 , \8995 , \8996 );
and \U$8195 ( \8998 , \8924_nG2ae9 , \8663 );
nor \U$8196 ( \8999 , \8993 , \8997 , \8998 );
and \U$8197 ( \9000 , \8770_nG2cf7 , \8578 );
and \U$8198 ( \9001 , \8623 , \8730_nG2df7 );
nand \U$8199 ( \9002 , \8770_nG2cf7 , \8575 );
or \U$8200 ( \9003 , \8535 , \8730_nG2df7 );
nand \U$8201 ( \9004 , \9003 , \8627 );
and \U$8202 ( \9005 , \9002 , \9004 );
nor \U$8203 ( \9006 , \9000 , \9001 , \9005 );
and \U$8204 ( \9007 , \8999 , \9006 );
not \U$8205 ( \9008 , \9007 );
and \U$8206 ( \9009 , RIb555fd0_401, \8462 );
and \U$8207 ( \9010 , RIb5560c0_403, \7917 );
and \U$8208 ( \9011 , \7955 , RIb556480_411);
and \U$8209 ( \9012 , RIb556408_410, \7926 );
nor \U$8210 ( \9013 , \9011 , \9012 );
and \U$8211 ( \9014 , \7938 , RIb5565e8_414);
and \U$8212 ( \9015 , RIb5561b0_405, \7900 );
nor \U$8213 ( \9016 , \9014 , \9015 );
and \U$8214 ( \9017 , \7948 , RIb5566d8_416);
and \U$8215 ( \9018 , RIb556660_415, \7936 );
nor \U$8216 ( \9019 , \9017 , \9018 );
and \U$8217 ( \9020 , \7906 , RIb5562a0_407);
and \U$8218 ( \9021 , RIb556390_409, \7910 );
nor \U$8219 ( \9022 , \9020 , \9021 );
nand \U$8220 ( \9023 , \9013 , \9016 , \9019 , \9022 );
nor \U$8221 ( \9024 , \9009 , \9010 , \9023 );
and \U$8222 ( \9025 , \7945 , RIb556570_413);
and \U$8223 ( \9026 , RIb556138_404, \7950 );
nor \U$8224 ( \9027 , \9025 , \9026 );
and \U$8225 ( \9028 , \7953 , RIb556228_406);
and \U$8226 ( \9029 , RIb556048_402, \7921 );
nor \U$8227 ( \9030 , \9028 , \9029 );
and \U$8228 ( \9031 , \7914 , RIb556318_408);
and \U$8229 ( \9032 , RIb5564f8_412, \7943 );
nor \U$8230 ( \9033 , \9031 , \9032 );
nand \U$8231 ( \9034 , \9024 , \9027 , \9030 , \9033 );
_DC g2a09 ( \9035_nG2a09 , \9034 , \8467 );
nand \U$8232 ( \9036 , \9035_nG2a09 , \8436 );
not \U$8233 ( \9037 , \9036 );
and \U$8234 ( \9038 , \9008 , \9037 );
nor \U$8235 ( \9039 , \8999 , \9006 );
nor \U$8236 ( \9040 , \9038 , \9039 );
or \U$8237 ( \9041 , \8945 , \8469 );
nand \U$8238 ( \9042 , \8943 , \8875 );
or \U$8239 ( \9043 , \8510 , \9042 );
or \U$8240 ( \9044 , \8947 , \8469 );
or \U$8241 ( \9045 , \8875 , \8508_nG3222 );
or \U$8242 ( \9046 , \8875 , \8943 );
nand \U$8243 ( \9047 , \9045 , \9046 );
nand \U$8244 ( \9048 , \9044 , \9047 );
nand \U$8245 ( \9049 , \9041 , \9043 , \9048 );
xor \U$8246 ( \9050 , \8268 , \8300_nG23c0 );
xor \U$8247 ( \9051 , \9050 , \8403 );
not \U$8248 ( \9052 , \9051 );
xor \U$8249 ( \9053 , \8232 , \8262_nG2495 );
xor \U$8250 ( \9054 , \9053 , \8406 );
not \U$8251 ( \9055 , \9054 );
and \U$8252 ( \9056 , \9052 , \9055 );
or \U$8253 ( \9057 , \8873 , \9056 );
and \U$8254 ( \9058 , \9049 , \9057 );
not \U$8255 ( \9059 , \9049 );
not \U$8256 ( \9060 , \9057 );
and \U$8257 ( \9061 , \9059 , \9060 );
nand \U$8258 ( \9062 , \8563_nG3003 , \8775 );
or \U$8259 ( \9063 , \8672 , \8658_nG2ee1 );
nand \U$8260 ( \9064 , \9063 , \8781 );
and \U$8261 ( \9065 , \9062 , \9064 );
and \U$8262 ( \9066 , \8777 , \8658_nG2ee1 );
and \U$8263 ( \9067 , \8563_nG3003 , \8866 );
nor \U$8264 ( \9068 , \9065 , \9066 , \9067 );
nor \U$8265 ( \9069 , \9061 , \9068 );
nor \U$8266 ( \9070 , \9058 , \9069 );
nor \U$8267 ( \9071 , \9040 , \9070 );
nand \U$8268 ( \9072 , \8992 , \9071 );
not \U$8269 ( \9073 , \8936 );
not \U$8270 ( \9074 , \8960 );
and \U$8271 ( \9075 , \9073 , \9074 );
and \U$8272 ( \9076 , \8936 , \8960 );
nor \U$8273 ( \9077 , \9075 , \9076 );
not \U$8274 ( \9078 , \9077 );
xor \U$8275 ( \9079 , \8970 , \8971 );
nand \U$8276 ( \9080 , \9078 , \9079 );
xor \U$8277 ( \9081 , \9072 , \9080 );
and \U$8278 ( \9082 , \8823 , \8889 );
nor \U$8279 ( \9083 , \9082 , \8890 );
and \U$8280 ( \9084 , \9081 , \9083 );
and \U$8281 ( \9085 , \9072 , \9080 );
or \U$8282 ( \9086 , \9084 , \9085 );
not \U$8283 ( \9087 , \8817 );
nand \U$8284 ( \9088 , \9087 , \8819 );
xor \U$8285 ( \9089 , \9086 , \9088 );
xor \U$8286 ( \9090 , \8890 , \8973 );
xor \U$8287 ( \9091 , \9090 , \8979 );
and \U$8288 ( \9092 , \9089 , \9091 );
and \U$8289 ( \9093 , \9086 , \9088 );
or \U$8290 ( \9094 , \9092 , \9093 );
not \U$8291 ( \9095 , \8982 );
not \U$8292 ( \9096 , \8984 );
nand \U$8293 ( \9097 , \9096 , \8816 );
not \U$8294 ( \9098 , \9097 );
or \U$8295 ( \9099 , \9095 , \9098 );
or \U$8296 ( \9100 , \9097 , \8982 );
nand \U$8297 ( \9101 , \9099 , \9100 );
xor \U$8298 ( \9102 , \9094 , \9101 );
not \U$8299 ( \9103 , \8972 );
not \U$8300 ( \9104 , \8961 );
or \U$8301 ( \9105 , \9103 , \9104 );
or \U$8302 ( \9106 , \8961 , \8972 );
nand \U$8303 ( \9107 , \9105 , \9106 );
not \U$8304 ( \9108 , \9079 );
not \U$8305 ( \9109 , \9077 );
or \U$8306 ( \9110 , \9108 , \9109 );
or \U$8307 ( \9111 , \9077 , \9079 );
nand \U$8308 ( \9112 , \9110 , \9111 );
not \U$8309 ( \9113 , \9054 );
not \U$8310 ( \9114 , \8873 );
or \U$8311 ( \9115 , \9113 , \9114 );
or \U$8312 ( \9116 , \8873 , \9054 );
nand \U$8313 ( \9117 , \9115 , \9116 );
xor \U$8314 ( \9118 , \9052 , \9055 );
nor \U$8315 ( \9119 , \9117 , \9118 );
not \U$8316 ( \9120 , \9119 );
not \U$8317 ( \9121 , \9057 );
nor \U$8318 ( \9122 , \9120 , \9121 );
not \U$8319 ( \9123 , \9122 );
or \U$8320 ( \9124 , \9123 , \8510 );
or \U$8321 ( \9125 , \9120 , \8510 );
nand \U$8322 ( \9126 , \9125 , \9121 );
nand \U$8323 ( \9127 , \9124 , \9126 );
or \U$8324 ( \9128 , \8945 , \8564 );
or \U$8325 ( \9129 , \8469 , \9042 );
or \U$8326 ( \9130 , \8947 , \8564 );
or \U$8327 ( \9131 , \8875 , \8468_nG310a );
nand \U$8328 ( \9132 , \9131 , \9046 );
nand \U$8329 ( \9133 , \9130 , \9132 );
nand \U$8330 ( \9134 , \9128 , \9129 , \9133 );
and \U$8331 ( \9135 , \9127 , \9134 );
and \U$8332 ( \9136 , \8857_nG2bf3 , \8578 );
and \U$8333 ( \9137 , \8623 , \8770_nG2cf7 );
nand \U$8334 ( \9138 , \8857_nG2bf3 , \8575 );
or \U$8335 ( \9139 , \8535 , \8770_nG2cf7 );
nand \U$8336 ( \9140 , \9139 , \8627 );
and \U$8337 ( \9141 , \9138 , \9140 );
nor \U$8338 ( \9142 , \9136 , \9137 , \9141 );
nand \U$8339 ( \9143 , \8658_nG2ee1 , \8775 );
or \U$8340 ( \9144 , \8672 , \8730_nG2df7 );
nand \U$8341 ( \9145 , \9144 , \8781 );
and \U$8342 ( \9146 , \9143 , \9145 );
and \U$8343 ( \9147 , \8777 , \8730_nG2df7 );
and \U$8344 ( \9148 , \8658_nG2ee1 , \8866 );
nor \U$8345 ( \9149 , \9146 , \9147 , \9148 );
xor \U$8346 ( \9150 , \9142 , \9149 );
and \U$8347 ( \9151 , \8924_nG2ae9 , \8521 );
or \U$8348 ( \9152 , \8481 , \9035_nG2a09 );
nand \U$8349 ( \9153 , \9152 , \8518 );
nand \U$8350 ( \9154 , \8924_nG2ae9 , \8514 );
and \U$8351 ( \9155 , \9153 , \9154 );
and \U$8352 ( \9156 , \9035_nG2a09 , \8663 );
nor \U$8353 ( \9157 , \9151 , \9155 , \9156 );
and \U$8354 ( \9158 , \9150 , \9157 );
and \U$8355 ( \9159 , \9142 , \9149 );
or \U$8356 ( \9160 , \9158 , \9159 );
not \U$8357 ( \9161 , \9160 );
and \U$8358 ( \9162 , \9135 , \9161 );
and \U$8359 ( \9163 , \9049 , \9057 );
not \U$8360 ( \9164 , \9049 );
and \U$8361 ( \9165 , \9164 , \9121 );
nor \U$8362 ( \9166 , \9163 , \9165 );
not \U$8363 ( \9167 , \9166 );
not \U$8364 ( \9168 , \9068 );
or \U$8365 ( \9169 , \9167 , \9168 );
or \U$8366 ( \9170 , \9068 , \9166 );
nand \U$8367 ( \9171 , \9169 , \9170 );
not \U$8368 ( \9172 , \9036 );
nor \U$8369 ( \9173 , \9007 , \9039 );
not \U$8370 ( \9174 , \9173 );
or \U$8371 ( \9175 , \9172 , \9174 );
or \U$8372 ( \9176 , \9173 , \9036 );
nand \U$8373 ( \9177 , \9175 , \9176 );
and \U$8374 ( \9178 , \9171 , \9177 );
and \U$8375 ( \9179 , \9162 , \9178 );
xor \U$8376 ( \9180 , \9112 , \9179 );
xnor \U$8377 ( \9181 , \9070 , \9040 );
not \U$8378 ( \9182 , \8988 );
not \U$8379 ( \9183 , \8990 );
and \U$8380 ( \9184 , \9182 , \9183 );
and \U$8381 ( \9185 , \8988 , \8990 );
nor \U$8382 ( \9186 , \9184 , \9185 );
nand \U$8383 ( \9187 , \9181 , \9186 );
and \U$8384 ( \9188 , \9180 , \9187 );
and \U$8385 ( \9189 , \9112 , \9179 );
or \U$8386 ( \9190 , \9188 , \9189 );
nand \U$8387 ( \9191 , \9107 , \9190 );
or \U$8388 ( \9192 , \9190 , \9107 );
nand \U$8389 ( \9193 , \9191 , \9192 );
not \U$8390 ( \9194 , \9193 );
xor \U$8391 ( \9195 , \9072 , \9080 );
xor \U$8392 ( \9196 , \9195 , \9083 );
not \U$8393 ( \9197 , \9196 );
and \U$8394 ( \9198 , \9194 , \9197 );
and \U$8395 ( \9199 , \9193 , \9196 );
nor \U$8396 ( \9200 , \9198 , \9199 );
not \U$8397 ( \9201 , \9071 );
not \U$8398 ( \9202 , \8991 );
or \U$8399 ( \9203 , \9201 , \9202 );
or \U$8400 ( \9204 , \8991 , \9071 );
nand \U$8401 ( \9205 , \9203 , \9204 );
xor \U$8402 ( \9206 , \9112 , \9179 );
xor \U$8403 ( \9207 , \9206 , \9187 );
and \U$8404 ( \9208 , \9205 , \9207 );
xor \U$8405 ( \9209 , \9135 , \9161 );
xor \U$8406 ( \9210 , \9171 , \9177 );
and \U$8407 ( \9211 , \9209 , \9210 );
xor \U$8408 ( \9212 , \9127 , \9134 );
xor \U$8409 ( \9213 , \9142 , \9149 );
xor \U$8410 ( \9214 , \9213 , \9157 );
not \U$8411 ( \9215 , \9214 );
and \U$8412 ( \9216 , \9212 , \9215 );
or \U$8413 ( \9217 , \9123 , \8469 );
and \U$8414 ( \9218 , \9057 , \9118 );
not \U$8415 ( \9219 , \9218 );
or \U$8416 ( \9220 , \8510 , \9219 );
or \U$8417 ( \9221 , \9120 , \8469 );
or \U$8418 ( \9222 , \9057 , \8508_nG3222 );
or \U$8419 ( \9223 , \9057 , \9118 );
nand \U$8420 ( \9224 , \9222 , \9223 );
nand \U$8421 ( \9225 , \9221 , \9224 );
nand \U$8422 ( \9226 , \9217 , \9220 , \9225 );
xor \U$8423 ( \9227 , RIb55bca0_599, \8363_nG2255 );
xor \U$8424 ( \9228 , \9227 , \8397 );
not \U$8425 ( \9229 , \9228 );
xor \U$8426 ( \9230 , \8302 , \8332_nG23c2 );
xor \U$8427 ( \9231 , \9230 , \8400 );
not \U$8428 ( \9232 , \9231 );
and \U$8429 ( \9233 , \9229 , \9232 );
or \U$8430 ( \9234 , \9051 , \9233 );
xor \U$8431 ( \9235 , \9226 , \9234 );
not \U$8432 ( \9236 , \8658_nG2ee1 );
or \U$8433 ( \9237 , \8945 , \9236 );
or \U$8434 ( \9238 , \8564 , \9042 );
or \U$8435 ( \9239 , \8947 , \9236 );
or \U$8436 ( \9240 , \8875 , \8563_nG3003 );
nand \U$8437 ( \9241 , \9240 , \9046 );
nand \U$8438 ( \9242 , \9239 , \9241 );
nand \U$8439 ( \9243 , \9237 , \9238 , \9242 );
and \U$8440 ( \9244 , \9235 , \9243 );
and \U$8441 ( \9245 , \9226 , \9234 );
or \U$8442 ( \9246 , \9244 , \9245 );
and \U$8443 ( \9247 , \8924_nG2ae9 , \8578 );
and \U$8444 ( \9248 , \8623 , \8857_nG2bf3 );
nand \U$8445 ( \9249 , \8924_nG2ae9 , \8575 );
or \U$8446 ( \9250 , \8535 , \8857_nG2bf3 );
nand \U$8447 ( \9251 , \9250 , \8627 );
and \U$8448 ( \9252 , \9249 , \9251 );
nor \U$8449 ( \9253 , \9247 , \9248 , \9252 );
nand \U$8450 ( \9254 , \8730_nG2df7 , \8775 );
or \U$8451 ( \9255 , \8672 , \8770_nG2cf7 );
nand \U$8452 ( \9256 , \9255 , \8781 );
and \U$8453 ( \9257 , \9254 , \9256 );
and \U$8454 ( \9258 , \8777 , \8770_nG2cf7 );
and \U$8455 ( \9259 , \8730_nG2df7 , \8866 );
nor \U$8456 ( \9260 , \9257 , \9258 , \9259 );
xor \U$8457 ( \9261 , \9253 , \9260 );
and \U$8458 ( \9262 , \9035_nG2a09 , \8521 );
and \U$8459 ( \9263 , RIb5559b8_388, \7900 );
and \U$8460 ( \9264 , RIb555e68_398, \7936 );
and \U$8461 ( \9265 , \7943 , RIb555d00_395);
and \U$8462 ( \9266 , RIb555d78_396, \7945 );
nor \U$8463 ( \9267 , \9265 , \9266 );
and \U$8464 ( \9268 , \7953 , RIb555a30_389);
and \U$8465 ( \9269 , RIb555940_387, \7950 );
nor \U$8466 ( \9270 , \9268 , \9269 );
and \U$8467 ( \9271 , \7917 , RIb5558c8_386);
and \U$8468 ( \9272 , RIb555850_385, \7921 );
nor \U$8469 ( \9273 , \9271 , \9272 );
and \U$8470 ( \9274 , \8462 , RIb5557d8_384);
and \U$8471 ( \9275 , RIb555b20_391, \7914 );
nor \U$8472 ( \9276 , \9274 , \9275 );
nand \U$8473 ( \9277 , \9267 , \9270 , \9273 , \9276 );
nor \U$8474 ( \9278 , \9263 , \9264 , \9277 );
and \U$8475 ( \9279 , \7938 , RIb555df0_397);
and \U$8476 ( \9280 , RIb555c88_394, \7955 );
nor \U$8477 ( \9281 , \9279 , \9280 );
and \U$8478 ( \9282 , \7948 , RIb555ee0_399);
and \U$8479 ( \9283 , RIb555c10_393, \7926 );
nor \U$8480 ( \9284 , \9282 , \9283 );
and \U$8481 ( \9285 , \7906 , RIb555aa8_390);
and \U$8482 ( \9286 , RIb555b98_392, \7910 );
nor \U$8483 ( \9287 , \9285 , \9286 );
nand \U$8484 ( \9288 , \9278 , \9281 , \9284 , \9287 );
_DC g290d ( \9289_nG290d , \9288 , \8467 );
or \U$8485 ( \9290 , \8481 , \9289_nG290d );
nand \U$8486 ( \9291 , \9290 , \8518 );
nand \U$8487 ( \9292 , \9035_nG2a09 , \8514 );
and \U$8488 ( \9293 , \9291 , \9292 );
and \U$8489 ( \9294 , \9289_nG290d , \8663 );
nor \U$8490 ( \9295 , \9262 , \9293 , \9294 );
and \U$8491 ( \9296 , \9261 , \9295 );
and \U$8492 ( \9297 , \9253 , \9260 );
or \U$8493 ( \9298 , \9296 , \9297 );
not \U$8494 ( \9299 , \9298 );
and \U$8495 ( \9300 , \9246 , \9299 );
and \U$8496 ( \9301 , \9216 , \9300 );
xor \U$8497 ( \9302 , \9211 , \9301 );
or \U$8498 ( \9303 , \9186 , \9181 );
nand \U$8499 ( \9304 , \9303 , \9187 );
and \U$8500 ( \9305 , \9302 , \9304 );
and \U$8501 ( \9306 , \9211 , \9301 );
or \U$8502 ( \9307 , \9305 , \9306 );
xor \U$8503 ( \9308 , \9112 , \9179 );
xor \U$8504 ( \9309 , \9308 , \9187 );
and \U$8505 ( \9310 , \9307 , \9309 );
and \U$8506 ( \9311 , \9205 , \9307 );
or \U$8507 ( \9312 , \9208 , \9310 , \9311 );
xor \U$8508 ( \9313 , \9200 , \9312 );
xor \U$8509 ( \9314 , \9212 , \9215 );
nand \U$8510 ( \9315 , \9289_nG290d , \8436 );
and \U$8511 ( \9316 , \9314 , \9315 );
xor \U$8512 ( \9317 , \9246 , \9299 );
nor \U$8513 ( \9318 , \9316 , \9317 );
and \U$8514 ( \9319 , RIb5571a0_439, \7900 );
and \U$8515 ( \9320 , RIb557470_445, \7955 );
and \U$8516 ( \9321 , \7943 , RIb5574e8_446);
and \U$8517 ( \9322 , RIb557560_447, \7945 );
nor \U$8518 ( \9323 , \9321 , \9322 );
and \U$8519 ( \9324 , \7953 , RIb557218_440);
and \U$8520 ( \9325 , RIb557128_438, \7950 );
nor \U$8521 ( \9326 , \9324 , \9325 );
and \U$8522 ( \9327 , \7917 , RIb5570b0_437);
and \U$8523 ( \9328 , RIb557038_436, \7921 );
nor \U$8524 ( \9329 , \9327 , \9328 );
and \U$8525 ( \9330 , \8462 , RIb556fc0_435);
and \U$8526 ( \9331 , RIb557308_442, \7914 );
nor \U$8527 ( \9332 , \9330 , \9331 );
nand \U$8528 ( \9333 , \9323 , \9326 , \9329 , \9332 );
nor \U$8529 ( \9334 , \9319 , \9320 , \9333 );
and \U$8530 ( \9335 , \7936 , RIb557650_449);
and \U$8531 ( \9336 , RIb5575d8_448, \7938 );
nor \U$8532 ( \9337 , \9335 , \9336 );
and \U$8533 ( \9338 , \7948 , RIb5576c8_450);
and \U$8534 ( \9339 , RIb557290_441, \7906 );
nor \U$8535 ( \9340 , \9338 , \9339 );
and \U$8536 ( \9341 , \7926 , RIb5573f8_444);
and \U$8537 ( \9342 , RIb557380_443, \7910 );
nor \U$8538 ( \9343 , \9341 , \9342 );
nand \U$8539 ( \9344 , \9334 , \9337 , \9340 , \9343 );
_DC g282e ( \9345_nG282e , \9344 , \8467 );
nand \U$8540 ( \9346 , \9345_nG282e , \8436 );
not \U$8541 ( \9347 , \9346 );
xor \U$8542 ( \9348 , \9226 , \9234 );
xor \U$8543 ( \9349 , \9348 , \9243 );
xor \U$8544 ( \9350 , \9253 , \9260 );
xor \U$8545 ( \9351 , \9350 , \9295 );
not \U$8546 ( \9352 , \9351 );
and \U$8547 ( \9353 , \9349 , \9352 );
nor \U$8548 ( \9354 , \9347 , \9353 );
not \U$8549 ( \9355 , \9354 );
or \U$8550 ( \9356 , \9051 , \9231 );
nand \U$8551 ( \9357 , \9231 , \9051 );
nand \U$8552 ( \9358 , \9356 , \9357 );
xor \U$8553 ( \9359 , \9229 , \9232 );
nor \U$8554 ( \9360 , \9358 , \9359 );
not \U$8555 ( \9361 , \9360 );
not \U$8556 ( \9362 , \9234 );
nor \U$8557 ( \9363 , \9361 , \9362 );
not \U$8558 ( \9364 , \9363 );
or \U$8559 ( \9365 , \9364 , \8510 );
or \U$8560 ( \9366 , \9361 , \8510 );
nand \U$8561 ( \9367 , \9366 , \9362 );
nand \U$8562 ( \9368 , \9365 , \9367 );
not \U$8563 ( \9369 , \9368 );
nand \U$8564 ( \9370 , \8563_nG3003 , \9119 );
or \U$8565 ( \9371 , \9057 , \8468_nG310a );
nand \U$8566 ( \9372 , \9371 , \9223 );
and \U$8567 ( \9373 , \9370 , \9372 );
and \U$8568 ( \9374 , \9218 , \8468_nG310a );
and \U$8569 ( \9375 , \8563_nG3003 , \9122 );
nor \U$8570 ( \9376 , \9373 , \9374 , \9375 );
nor \U$8571 ( \9377 , \9369 , \9376 );
not \U$8572 ( \9378 , \9377 );
nand \U$8573 ( \9379 , \8770_nG2cf7 , \8775 );
or \U$8574 ( \9380 , \8672 , \8857_nG2bf3 );
nand \U$8575 ( \9381 , \9380 , \8781 );
and \U$8576 ( \9382 , \9379 , \9381 );
and \U$8577 ( \9383 , \8777 , \8857_nG2bf3 );
and \U$8578 ( \9384 , \8770_nG2cf7 , \8866 );
nor \U$8579 ( \9385 , \9382 , \9383 , \9384 );
nand \U$8580 ( \9386 , \8730_nG2df7 , \8944 );
or \U$8581 ( \9387 , \8875 , \8658_nG2ee1 );
nand \U$8582 ( \9388 , \9387 , \9046 );
and \U$8583 ( \9389 , \9386 , \9388 );
not \U$8584 ( \9390 , \9042 );
and \U$8585 ( \9391 , \9390 , \8658_nG2ee1 );
not \U$8586 ( \9392 , \8945 );
and \U$8587 ( \9393 , \8730_nG2df7 , \9392 );
nor \U$8588 ( \9394 , \9389 , \9391 , \9393 );
xor \U$8589 ( \9395 , \9385 , \9394 );
and \U$8590 ( \9396 , \9035_nG2a09 , \8578 );
and \U$8591 ( \9397 , \8623 , \8924_nG2ae9 );
nand \U$8592 ( \9398 , \9035_nG2a09 , \8575 );
or \U$8593 ( \9399 , \8535 , \8924_nG2ae9 );
nand \U$8594 ( \9400 , \9399 , \8627 );
and \U$8595 ( \9401 , \9398 , \9400 );
nor \U$8596 ( \9402 , \9396 , \9397 , \9401 );
and \U$8597 ( \9403 , \9395 , \9402 );
and \U$8598 ( \9404 , \9385 , \9394 );
or \U$8599 ( \9405 , \9403 , \9404 );
nor \U$8600 ( \9406 , \9378 , \9405 );
nand \U$8601 ( \9407 , \9355 , \9406 );
or \U$8602 ( \9408 , \9318 , \9407 );
not \U$8603 ( \9409 , \9407 );
not \U$8604 ( \9410 , \9318 );
or \U$8605 ( \9411 , \9409 , \9410 );
xor \U$8606 ( \9412 , \9209 , \9210 );
nand \U$8607 ( \9413 , \9411 , \9412 );
nand \U$8608 ( \9414 , \9408 , \9413 );
xor \U$8609 ( \9415 , \9162 , \9178 );
xor \U$8610 ( \9416 , \9414 , \9415 );
xor \U$8611 ( \9417 , \9211 , \9301 );
xor \U$8612 ( \9418 , \9417 , \9304 );
and \U$8613 ( \9419 , \9416 , \9418 );
and \U$8614 ( \9420 , \9414 , \9415 );
or \U$8615 ( \9421 , \9419 , \9420 );
xor \U$8616 ( \9422 , \9112 , \9179 );
xor \U$8617 ( \9423 , \9422 , \9187 );
xor \U$8618 ( \9424 , \9205 , \9307 );
xor \U$8619 ( \9425 , \9423 , \9424 );
xor \U$8620 ( \9426 , \9421 , \9425 );
xor \U$8621 ( \9427 , \9414 , \9415 );
xor \U$8622 ( \9428 , \9427 , \9418 );
xnor \U$8623 ( \9429 , \9407 , \9318 );
not \U$8624 ( \9430 , \9429 );
not \U$8625 ( \9431 , \9412 );
and \U$8626 ( \9432 , \9430 , \9431 );
and \U$8627 ( \9433 , \9429 , \9412 );
nor \U$8628 ( \9434 , \9432 , \9433 );
not \U$8629 ( \9435 , \9314 );
not \U$8630 ( \9436 , \9317 );
nand \U$8631 ( \9437 , \9436 , \9315 );
not \U$8632 ( \9438 , \9437 );
and \U$8633 ( \9439 , \9435 , \9438 );
and \U$8634 ( \9440 , \9314 , \9437 );
nor \U$8635 ( \9441 , \9439 , \9440 );
not \U$8636 ( \9442 , \9376 );
not \U$8637 ( \9443 , \9368 );
and \U$8638 ( \9444 , \9442 , \9443 );
and \U$8639 ( \9445 , \9376 , \9368 );
nor \U$8640 ( \9446 , \9444 , \9445 );
xor \U$8641 ( \9447 , \9385 , \9394 );
xor \U$8642 ( \9448 , \9447 , \9402 );
and \U$8643 ( \9449 , \9446 , \9448 );
and \U$8644 ( \9450 , RIb556840_419, \7921 );
and \U$8645 ( \9451 , RIb556d68_430, \7945 );
and \U$8646 ( \9452 , \7906 , RIb556a98_424);
and \U$8647 ( \9453 , RIb556b88_426, \7910 );
nor \U$8648 ( \9454 , \9452 , \9453 );
and \U$8649 ( \9455 , \7948 , RIb556ed0_433);
and \U$8650 ( \9456 , RIb556c78_428, \7955 );
nor \U$8651 ( \9457 , \9455 , \9456 );
and \U$8652 ( \9458 , \7926 , RIb556c00_427);
and \U$8653 ( \9459 , RIb5569a8_422, \7900 );
nor \U$8654 ( \9460 , \9458 , \9459 );
and \U$8655 ( \9461 , \7936 , RIb556e58_432);
and \U$8656 ( \9462 , RIb556de0_431, \7938 );
nor \U$8657 ( \9463 , \9461 , \9462 );
nand \U$8658 ( \9464 , \9454 , \9457 , \9460 , \9463 );
nor \U$8659 ( \9465 , \9450 , \9451 , \9464 );
and \U$8660 ( \9466 , \7914 , RIb556b10_425);
and \U$8661 ( \9467 , RIb556cf0_429, \7943 );
nor \U$8662 ( \9468 , \9466 , \9467 );
and \U$8663 ( \9469 , \7950 , RIb556930_421);
and \U$8664 ( \9470 , RIb5568b8_420, \7917 );
nor \U$8665 ( \9471 , \9469 , \9470 );
and \U$8666 ( \9472 , \8462 , RIb5567c8_418);
and \U$8667 ( \9473 , RIb556a20_423, \7953 );
nor \U$8668 ( \9474 , \9472 , \9473 );
nand \U$8669 ( \9475 , \9465 , \9468 , \9471 , \9474 );
_DC g2758 ( \9476_nG2758 , \9475 , \8467 );
nand \U$8670 ( \9477 , \9476_nG2758 , \8436 );
and \U$8671 ( \9478 , \9289_nG290d , \8521 );
or \U$8672 ( \9479 , \8481 , \9345_nG282e );
nand \U$8673 ( \9480 , \9479 , \8518 );
nand \U$8674 ( \9481 , \9289_nG290d , \8514 );
and \U$8675 ( \9482 , \9480 , \9481 );
and \U$8676 ( \9483 , \9345_nG282e , \8663 );
nor \U$8677 ( \9484 , \9478 , \9482 , \9483 );
xnor \U$8678 ( \9485 , \9477 , \9484 );
xor \U$8679 ( \9486 , \9385 , \9394 );
xor \U$8680 ( \9487 , \9486 , \9402 );
and \U$8681 ( \9488 , \9485 , \9487 );
and \U$8682 ( \9489 , \9446 , \9485 );
or \U$8683 ( \9490 , \9449 , \9488 , \9489 );
not \U$8684 ( \9491 , \9490 );
nand \U$8685 ( \9492 , \8857_nG2bf3 , \8775 );
or \U$8686 ( \9493 , \8672 , \8924_nG2ae9 );
nand \U$8687 ( \9494 , \9493 , \8781 );
and \U$8688 ( \9495 , \9492 , \9494 );
and \U$8689 ( \9496 , \8777 , \8924_nG2ae9 );
and \U$8690 ( \9497 , \8857_nG2bf3 , \8866 );
nor \U$8691 ( \9498 , \9495 , \9496 , \9497 );
nand \U$8692 ( \9499 , \8770_nG2cf7 , \8944 );
or \U$8693 ( \9500 , \8875 , \8730_nG2df7 );
nand \U$8694 ( \9501 , \9500 , \9046 );
and \U$8695 ( \9502 , \9499 , \9501 );
and \U$8696 ( \9503 , \9390 , \8730_nG2df7 );
and \U$8697 ( \9504 , \8770_nG2cf7 , \9392 );
nor \U$8698 ( \9505 , \9502 , \9503 , \9504 );
xor \U$8699 ( \9506 , \9498 , \9505 );
and \U$8700 ( \9507 , \9289_nG290d , \8578 );
and \U$8701 ( \9508 , \8623 , \9035_nG2a09 );
nand \U$8702 ( \9509 , \9289_nG290d , \8575 );
or \U$8703 ( \9510 , \8535 , \9035_nG2a09 );
nand \U$8704 ( \9511 , \9510 , \8627 );
and \U$8705 ( \9512 , \9509 , \9511 );
nor \U$8706 ( \9513 , \9507 , \9508 , \9512 );
and \U$8707 ( \9514 , \9506 , \9513 );
and \U$8708 ( \9515 , \9498 , \9505 );
or \U$8709 ( \9516 , \9514 , \9515 );
nand \U$8710 ( \9517 , \8468_nG310a , \9360 );
or \U$8711 ( \9518 , \9234 , \8508_nG3222 );
or \U$8712 ( \9519 , \9234 , \9359 );
nand \U$8713 ( \9520 , \9518 , \9519 );
and \U$8714 ( \9521 , \9517 , \9520 );
and \U$8715 ( \9522 , \9234 , \9359 );
and \U$8716 ( \9523 , \9522 , \8508_nG3222 );
and \U$8717 ( \9524 , \8468_nG310a , \9363 );
nor \U$8718 ( \9525 , \9521 , \9523 , \9524 );
nand \U$8719 ( \9526 , \8658_nG2ee1 , \9119 );
or \U$8720 ( \9527 , \9057 , \8563_nG3003 );
nand \U$8721 ( \9528 , \9527 , \9223 );
and \U$8722 ( \9529 , \9526 , \9528 );
and \U$8723 ( \9530 , \9218 , \8563_nG3003 );
and \U$8724 ( \9531 , \8658_nG2ee1 , \9122 );
nor \U$8725 ( \9532 , \9529 , \9530 , \9531 );
nand \U$8726 ( \9533 , \9525 , \9532 );
and \U$8727 ( \9534 , \9533 , \9228 );
nor \U$8728 ( \9535 , \9532 , \9525 );
nor \U$8729 ( \9536 , \9534 , \9535 );
nor \U$8730 ( \9537 , \9516 , \9536 );
nand \U$8731 ( \9538 , \9491 , \9537 );
xor \U$8732 ( \9539 , \9441 , \9538 );
xor \U$8733 ( \9540 , \9349 , \9352 );
not \U$8734 ( \9541 , \9540 );
not \U$8735 ( \9542 , \9346 );
and \U$8736 ( \9543 , \9541 , \9542 );
and \U$8737 ( \9544 , \9540 , \9346 );
nor \U$8738 ( \9545 , \9543 , \9544 );
not \U$8739 ( \9546 , \9545 );
or \U$8740 ( \9547 , \9405 , \9377 );
or \U$8741 ( \9548 , \9477 , \9484 );
nand \U$8742 ( \9549 , \9377 , \9405 );
nand \U$8743 ( \9550 , \9547 , \9548 , \9549 );
nand \U$8744 ( \9551 , \9546 , \9550 );
and \U$8745 ( \9552 , \9539 , \9551 );
and \U$8746 ( \9553 , \9441 , \9538 );
or \U$8747 ( \9554 , \9552 , \9553 );
nor \U$8748 ( \9555 , \9434 , \9554 );
not \U$8749 ( \9556 , \9555 );
not \U$8750 ( \9557 , \9315 );
nor \U$8751 ( \9558 , \9557 , \9300 );
not \U$8752 ( \9559 , \9558 );
not \U$8753 ( \9560 , \9216 );
or \U$8754 ( \9561 , \9559 , \9560 );
or \U$8755 ( \9562 , \9216 , \9558 );
nand \U$8756 ( \9563 , \9561 , \9562 );
not \U$8757 ( \9564 , \9563 );
and \U$8758 ( \9565 , \9556 , \9564 );
and \U$8759 ( \9566 , \9434 , \9554 );
nor \U$8760 ( \9567 , \9565 , \9566 );
xor \U$8761 ( \9568 , \9428 , \9567 );
xor \U$8762 ( \9569 , \9441 , \9538 );
xor \U$8763 ( \9570 , \9569 , \9551 );
not \U$8764 ( \9571 , \9550 );
not \U$8765 ( \9572 , \9545 );
or \U$8766 ( \9573 , \9571 , \9572 );
or \U$8767 ( \9574 , \9545 , \9550 );
nand \U$8768 ( \9575 , \9573 , \9574 );
not \U$8769 ( \9576 , \9537 );
not \U$8770 ( \9577 , \9490 );
or \U$8771 ( \9578 , \9576 , \9577 );
or \U$8772 ( \9579 , \9490 , \9537 );
nand \U$8773 ( \9580 , \9578 , \9579 );
and \U$8774 ( \9581 , \9575 , \9580 );
not \U$8775 ( \9582 , \9575 );
not \U$8776 ( \9583 , \9580 );
and \U$8777 ( \9584 , \9582 , \9583 );
nand \U$8778 ( \9585 , \8857_nG2bf3 , \8944 );
or \U$8779 ( \9586 , \8875 , \8770_nG2cf7 );
nand \U$8780 ( \9587 , \9586 , \9046 );
and \U$8781 ( \9588 , \9585 , \9587 );
and \U$8782 ( \9589 , \9390 , \8770_nG2cf7 );
and \U$8783 ( \9590 , \8857_nG2bf3 , \9392 );
nor \U$8784 ( \9591 , \9588 , \9589 , \9590 );
nand \U$8785 ( \9592 , \8730_nG2df7 , \9119 );
or \U$8786 ( \9593 , \9057 , \8658_nG2ee1 );
nand \U$8787 ( \9594 , \9593 , \9223 );
and \U$8788 ( \9595 , \9592 , \9594 );
and \U$8789 ( \9596 , \9218 , \8658_nG2ee1 );
and \U$8790 ( \9597 , \8730_nG2df7 , \9122 );
nor \U$8791 ( \9598 , \9595 , \9596 , \9597 );
xor \U$8792 ( \9599 , \9591 , \9598 );
nand \U$8793 ( \9600 , \8924_nG2ae9 , \8775 );
or \U$8794 ( \9601 , \8672 , \9035_nG2a09 );
nand \U$8795 ( \9602 , \9601 , \8781 );
and \U$8796 ( \9603 , \9600 , \9602 );
and \U$8797 ( \9604 , \8777 , \9035_nG2a09 );
and \U$8798 ( \9605 , \8924_nG2ae9 , \8866 );
nor \U$8799 ( \9606 , \9603 , \9604 , \9605 );
and \U$8800 ( \9607 , \9599 , \9606 );
and \U$8801 ( \9608 , \9591 , \9598 );
or \U$8802 ( \9609 , \9607 , \9608 );
and \U$8803 ( \9610 , \9476_nG2758 , \8521 );
and \U$8804 ( \9611 , RIb557fb0_469, \8462 );
and \U$8805 ( \9612 , RIb5580a0_471, \7917 );
and \U$8806 ( \9613 , \7955 , RIb558460_479);
and \U$8807 ( \9614 , RIb5583e8_478, \7926 );
nor \U$8808 ( \9615 , \9613 , \9614 );
and \U$8809 ( \9616 , \7948 , RIb5586b8_484);
and \U$8810 ( \9617 , RIb558370_477, \7910 );
nor \U$8811 ( \9618 , \9616 , \9617 );
and \U$8812 ( \9619 , \7906 , RIb558280_475);
and \U$8813 ( \9620 , RIb558190_473, \7900 );
nor \U$8814 ( \9621 , \9619 , \9620 );
and \U$8815 ( \9622 , \7936 , RIb558640_483);
and \U$8816 ( \9623 , RIb5585c8_482, \7938 );
nor \U$8817 ( \9624 , \9622 , \9623 );
nand \U$8818 ( \9625 , \9615 , \9618 , \9621 , \9624 );
nor \U$8819 ( \9626 , \9611 , \9612 , \9625 );
and \U$8820 ( \9627 , \7945 , RIb558550_481);
and \U$8821 ( \9628 , RIb558118_472, \7950 );
nor \U$8822 ( \9629 , \9627 , \9628 );
and \U$8823 ( \9630 , \7953 , RIb558208_474);
and \U$8824 ( \9631 , RIb558028_470, \7921 );
nor \U$8825 ( \9632 , \9630 , \9631 );
and \U$8826 ( \9633 , \7914 , RIb5582f8_476);
and \U$8827 ( \9634 , RIb5584d8_480, \7943 );
nor \U$8828 ( \9635 , \9633 , \9634 );
nand \U$8829 ( \9636 , \9626 , \9629 , \9632 , \9635 );
_DC g26ac ( \9637_nG26ac , \9636 , \8467 );
or \U$8830 ( \9638 , \8481 , \9637_nG26ac );
nand \U$8831 ( \9639 , \9638 , \8518 );
nand \U$8832 ( \9640 , \9476_nG2758 , \8514 );
and \U$8833 ( \9641 , \9639 , \9640 );
and \U$8834 ( \9642 , \9637_nG26ac , \8663 );
nor \U$8835 ( \9643 , \9610 , \9641 , \9642 );
and \U$8836 ( \9644 , \9345_nG282e , \8578 );
and \U$8837 ( \9645 , \8623 , \9289_nG290d );
nand \U$8838 ( \9646 , \9345_nG282e , \8575 );
or \U$8839 ( \9647 , \8535 , \9289_nG290d );
nand \U$8840 ( \9648 , \9647 , \8627 );
and \U$8841 ( \9649 , \9646 , \9648 );
nor \U$8842 ( \9650 , \9644 , \9645 , \9649 );
and \U$8843 ( \9651 , \9643 , \9650 );
not \U$8844 ( \9652 , \9651 );
and \U$8845 ( \9653 , RIb557830_453, \7921 );
and \U$8846 ( \9654 , RIb557d58_464, \7945 );
and \U$8847 ( \9655 , \7955 , RIb557c68_462);
and \U$8848 ( \9656 , RIb557bf0_461, \7926 );
nor \U$8849 ( \9657 , \9655 , \9656 );
and \U$8850 ( \9658 , \7938 , RIb557dd0_465);
and \U$8851 ( \9659 , RIb557998_456, \7900 );
nor \U$8852 ( \9660 , \9658 , \9659 );
and \U$8853 ( \9661 , \7948 , RIb557ec0_467);
and \U$8854 ( \9662 , RIb557e48_466, \7936 );
nor \U$8855 ( \9663 , \9661 , \9662 );
and \U$8856 ( \9664 , \7906 , RIb557a88_458);
and \U$8857 ( \9665 , RIb557b78_460, \7910 );
nor \U$8858 ( \9666 , \9664 , \9665 );
nand \U$8859 ( \9667 , \9657 , \9660 , \9663 , \9666 );
nor \U$8860 ( \9668 , \9653 , \9654 , \9667 );
and \U$8861 ( \9669 , \7914 , RIb557b00_459);
and \U$8862 ( \9670 , RIb557ce0_463, \7943 );
nor \U$8863 ( \9671 , \9669 , \9670 );
and \U$8864 ( \9672 , \7950 , RIb557920_455);
and \U$8865 ( \9673 , RIb5578a8_454, \7917 );
nor \U$8866 ( \9674 , \9672 , \9673 );
and \U$8867 ( \9675 , \8462 , RIb5577b8_452);
and \U$8868 ( \9676 , RIb557a10_457, \7953 );
nor \U$8869 ( \9677 , \9675 , \9676 );
nand \U$8870 ( \9678 , \9668 , \9671 , \9674 , \9677 );
_DC g25e2 ( \9679_nG25e2 , \9678 , \8467 );
nand \U$8871 ( \9680 , \9679_nG25e2 , \8436 );
not \U$8872 ( \9681 , \9680 );
and \U$8873 ( \9682 , \9652 , \9681 );
nor \U$8874 ( \9683 , \9643 , \9650 );
nor \U$8875 ( \9684 , \9682 , \9683 );
nand \U$8876 ( \9685 , \9609 , \9684 );
or \U$8877 ( \9686 , \9228 , \8508_nG3222 );
or \U$8878 ( \9687 , \8395 , \8394_nG2253 );
nand \U$8879 ( \9688 , \9687 , \8396 );
nor \U$8880 ( \9689 , \9228 , \9688 );
not \U$8881 ( \9690 , \9689 );
nand \U$8882 ( \9691 , \9229 , \9690 );
nand \U$8883 ( \9692 , \9686 , \9691 );
or \U$8884 ( \9693 , \9364 , \8564 );
not \U$8885 ( \9694 , \9522 );
or \U$8886 ( \9695 , \8469 , \9694 );
or \U$8887 ( \9696 , \9361 , \8564 );
or \U$8888 ( \9697 , \9234 , \8468_nG310a );
nand \U$8889 ( \9698 , \9697 , \9519 );
nand \U$8890 ( \9699 , \9696 , \9698 );
nand \U$8891 ( \9700 , \9693 , \9695 , \9699 );
and \U$8892 ( \9701 , \9692 , \9700 );
and \U$8893 ( \9702 , \9685 , \9701 );
nor \U$8894 ( \9703 , \9684 , \9609 );
nor \U$8895 ( \9704 , \9702 , \9703 );
nand \U$8896 ( \9705 , \9637_nG26ac , \8436 );
and \U$8897 ( \9706 , \9345_nG282e , \8521 );
or \U$8898 ( \9707 , \8481 , \9476_nG2758 );
nand \U$8899 ( \9708 , \9707 , \8518 );
nand \U$8900 ( \9709 , \9345_nG282e , \8514 );
and \U$8901 ( \9710 , \9708 , \9709 );
and \U$8902 ( \9711 , \9476_nG2758 , \8663 );
nor \U$8903 ( \9712 , \9706 , \9710 , \9711 );
xnor \U$8904 ( \9713 , \9705 , \9712 );
xor \U$8905 ( \9714 , \9704 , \9713 );
xor \U$8906 ( \9715 , \9385 , \9394 );
xor \U$8907 ( \9716 , \9715 , \9402 );
xor \U$8908 ( \9717 , \9446 , \9485 );
xor \U$8909 ( \9718 , \9716 , \9717 );
and \U$8910 ( \9719 , \9714 , \9718 );
and \U$8911 ( \9720 , \9704 , \9713 );
or \U$8912 ( \9721 , \9719 , \9720 );
nor \U$8913 ( \9722 , \9584 , \9721 );
nor \U$8914 ( \9723 , \9581 , \9722 );
nand \U$8915 ( \9724 , \9570 , \9723 );
not \U$8916 ( \9725 , \9724 );
nor \U$8917 ( \9726 , \9723 , \9570 );
nor \U$8918 ( \9727 , \9725 , \9726 );
not \U$8919 ( \9728 , \9727 );
not \U$8920 ( \9729 , \9406 );
not \U$8921 ( \9730 , \9354 );
or \U$8922 ( \9731 , \9729 , \9730 );
or \U$8923 ( \9732 , \9354 , \9406 );
nand \U$8924 ( \9733 , \9731 , \9732 );
not \U$8925 ( \9734 , \9733 );
and \U$8926 ( \9735 , \9728 , \9734 );
and \U$8927 ( \9736 , \9727 , \9733 );
nor \U$8928 ( \9737 , \9735 , \9736 );
or \U$8929 ( \9738 , \9712 , \9705 );
not \U$8930 ( \9739 , \9536 );
or \U$8931 ( \9740 , \9739 , \9516 );
not \U$8932 ( \9741 , \9516 );
or \U$8933 ( \9742 , \9536 , \9741 );
nand \U$8934 ( \9743 , \9738 , \9740 , \9742 );
xor \U$8935 ( \9744 , \9704 , \9713 );
xor \U$8936 ( \9745 , \9744 , \9718 );
not \U$8937 ( \9746 , \9745 );
and \U$8938 ( \9747 , \9743 , \9746 );
not \U$8939 ( \9748 , \9228 );
not \U$8940 ( \9749 , \9535 );
nand \U$8941 ( \9750 , \9749 , \9533 );
not \U$8942 ( \9751 , \9750 );
or \U$8943 ( \9752 , \9748 , \9751 );
or \U$8944 ( \9753 , \9750 , \9228 );
nand \U$8945 ( \9754 , \9752 , \9753 );
xor \U$8946 ( \9755 , \9713 , \9754 );
not \U$8947 ( \9756 , \9701 );
not \U$8948 ( \9757 , \9703 );
nand \U$8949 ( \9758 , \9757 , \9685 );
not \U$8950 ( \9759 , \9758 );
or \U$8951 ( \9760 , \9756 , \9759 );
or \U$8952 ( \9761 , \9758 , \9701 );
nand \U$8953 ( \9762 , \9760 , \9761 );
and \U$8954 ( \9763 , \9755 , \9762 );
and \U$8955 ( \9764 , \9713 , \9754 );
or \U$8956 ( \9765 , \9763 , \9764 );
not \U$8957 ( \9766 , \9765 );
xor \U$8958 ( \9767 , \9591 , \9598 );
xor \U$8959 ( \9768 , \9767 , \9606 );
not \U$8960 ( \9769 , \9768 );
not \U$8961 ( \9770 , \9680 );
nor \U$8962 ( \9771 , \9651 , \9683 );
not \U$8963 ( \9772 , \9771 );
or \U$8964 ( \9773 , \9770 , \9772 );
or \U$8965 ( \9774 , \9771 , \9680 );
nand \U$8966 ( \9775 , \9773 , \9774 );
and \U$8967 ( \9776 , \9769 , \9775 );
nand \U$8968 ( \9777 , \9035_nG2a09 , \8775 );
or \U$8969 ( \9778 , \8672 , \9289_nG290d );
nand \U$8970 ( \9779 , \9778 , \8781 );
and \U$8971 ( \9780 , \9777 , \9779 );
and \U$8972 ( \9781 , \8777 , \9289_nG290d );
and \U$8973 ( \9782 , \9035_nG2a09 , \8866 );
nor \U$8974 ( \9783 , \9780 , \9781 , \9782 );
nand \U$8975 ( \9784 , \8924_nG2ae9 , \8944 );
or \U$8976 ( \9785 , \8875 , \8857_nG2bf3 );
nand \U$8977 ( \9786 , \9785 , \9046 );
and \U$8978 ( \9787 , \9784 , \9786 );
and \U$8979 ( \9788 , \9390 , \8857_nG2bf3 );
and \U$8980 ( \9789 , \8924_nG2ae9 , \9392 );
nor \U$8981 ( \9790 , \9787 , \9788 , \9789 );
xor \U$8982 ( \9791 , \9783 , \9790 );
and \U$8983 ( \9792 , \9476_nG2758 , \8578 );
and \U$8984 ( \9793 , \8623 , \9345_nG282e );
nand \U$8985 ( \9794 , \9476_nG2758 , \8575 );
or \U$8986 ( \9795 , \8535 , \9345_nG282e );
nand \U$8987 ( \9796 , \9795 , \8627 );
and \U$8988 ( \9797 , \9794 , \9796 );
nor \U$8989 ( \9798 , \9792 , \9793 , \9797 );
and \U$8990 ( \9799 , \9791 , \9798 );
and \U$8991 ( \9800 , \9783 , \9790 );
or \U$8992 ( \9801 , \9799 , \9800 );
nand \U$8993 ( \9802 , \8658_nG2ee1 , \9360 );
or \U$8994 ( \9803 , \9234 , \8563_nG3003 );
nand \U$8995 ( \9804 , \9803 , \9519 );
and \U$8996 ( \9805 , \9802 , \9804 );
and \U$8997 ( \9806 , \9522 , \8563_nG3003 );
and \U$8998 ( \9807 , \8658_nG2ee1 , \9363 );
nor \U$8999 ( \9808 , \9805 , \9806 , \9807 );
not \U$9000 ( \9809 , \9808 );
not \U$9001 ( \9810 , \9691 );
and \U$9002 ( \9811 , \8510 , \9810 );
and \U$9003 ( \9812 , \9689 , \8469 );
nand \U$9004 ( \9813 , \9688 , \9228 );
not \U$9005 ( \9814 , \9813 );
and \U$9006 ( \9815 , \8508_nG3222 , \9814 );
nor \U$9007 ( \9816 , \9811 , \9812 , \9815 );
not \U$9008 ( \9817 , \9816 );
and \U$9009 ( \9818 , \9809 , \9817 );
and \U$9010 ( \9819 , \9808 , \9816 );
nand \U$9011 ( \9820 , \8770_nG2cf7 , \9119 );
or \U$9012 ( \9821 , \9057 , \8730_nG2df7 );
nand \U$9013 ( \9822 , \9821 , \9223 );
and \U$9014 ( \9823 , \9820 , \9822 );
and \U$9015 ( \9824 , \9218 , \8730_nG2df7 );
and \U$9016 ( \9825 , \8770_nG2cf7 , \9122 );
nor \U$9017 ( \9826 , \9823 , \9824 , \9825 );
nor \U$9018 ( \9827 , \9819 , \9826 );
nor \U$9019 ( \9828 , \9818 , \9827 );
nor \U$9020 ( \9829 , \9801 , \9828 );
not \U$9021 ( \9830 , \9829 );
xor \U$9022 ( \9831 , \9498 , \9505 );
xor \U$9023 ( \9832 , \9831 , \9513 );
nand \U$9024 ( \9833 , \9830 , \9832 );
and \U$9025 ( \9834 , \9776 , \9833 );
not \U$9026 ( \9835 , \9832 );
and \U$9027 ( \9836 , \9835 , \9829 );
nor \U$9028 ( \9837 , \9834 , \9836 );
nand \U$9029 ( \9838 , \9766 , \9837 );
xor \U$9030 ( \9839 , \9747 , \9838 );
not \U$9031 ( \9840 , \9721 );
xor \U$9032 ( \9841 , \9580 , \9575 );
not \U$9033 ( \9842 , \9841 );
or \U$9034 ( \9843 , \9840 , \9842 );
or \U$9035 ( \9844 , \9841 , \9721 );
nand \U$9036 ( \9845 , \9843 , \9844 );
and \U$9037 ( \9846 , \9839 , \9845 );
and \U$9038 ( \9847 , \9747 , \9838 );
or \U$9039 ( \9848 , \9846 , \9847 );
xor \U$9040 ( \9849 , \9737 , \9848 );
xor \U$9041 ( \9850 , \9743 , \9746 );
not \U$9042 ( \9851 , \9765 );
not \U$9043 ( \9852 , \9837 );
and \U$9044 ( \9853 , \9851 , \9852 );
and \U$9045 ( \9854 , \9765 , \9837 );
nor \U$9046 ( \9855 , \9853 , \9854 );
xor \U$9047 ( \9856 , \9850 , \9855 );
xor \U$9048 ( \9857 , \9783 , \9790 );
xor \U$9049 ( \9858 , \9857 , \9798 );
not \U$9050 ( \9859 , \9858 );
and \U$9051 ( \9860 , RIb559450_513, \7955 );
and \U$9052 ( \9861 , RIb5595b8_516, \7938 );
and \U$9053 ( \9862 , \7926 , RIb5593d8_512);
and \U$9054 ( \9863 , RIb559360_511, \7910 );
nor \U$9055 ( \9864 , \9862 , \9863 );
and \U$9056 ( \9865 , \8462 , RIb558fa0_503);
and \U$9057 ( \9866 , RIb559018_504, \7921 );
nor \U$9058 ( \9867 , \9865 , \9866 );
and \U$9059 ( \9868 , \7950 , RIb559108_506);
and \U$9060 ( \9869 , RIb559090_505, \7917 );
nor \U$9061 ( \9870 , \9868 , \9869 );
and \U$9062 ( \9871 , \7906 , RIb559270_509);
and \U$9063 ( \9872 , RIb5591f8_508, \7953 );
nor \U$9064 ( \9873 , \9871 , \9872 );
nand \U$9065 ( \9874 , \9864 , \9867 , \9870 , \9873 );
nor \U$9066 ( \9875 , \9860 , \9861 , \9874 );
and \U$9067 ( \9876 , \7914 , RIb5592e8_510);
and \U$9068 ( \9877 , RIb559540_515, \7945 );
nor \U$9069 ( \9878 , \9876 , \9877 );
and \U$9070 ( \9879 , \7948 , RIb5596a8_518);
and \U$9071 ( \9880 , RIb559180_507, \7900 );
nor \U$9072 ( \9881 , \9879 , \9880 );
and \U$9073 ( \9882 , \7936 , RIb559630_517);
and \U$9074 ( \9883 , RIb5594c8_514, \7943 );
nor \U$9075 ( \9884 , \9882 , \9883 );
nand \U$9076 ( \9885 , \9875 , \9878 , \9881 , \9884 );
_DC g2554 ( \9886_nG2554 , \9885 , \8467 );
nand \U$9077 ( \9887 , \9886_nG2554 , \8436 );
and \U$9078 ( \9888 , \9637_nG26ac , \8521 );
or \U$9079 ( \9889 , \8481 , \9679_nG25e2 );
nand \U$9080 ( \9890 , \9889 , \8518 );
nand \U$9081 ( \9891 , \9637_nG26ac , \8514 );
and \U$9082 ( \9892 , \9890 , \9891 );
and \U$9083 ( \9893 , \9679_nG25e2 , \8663 );
nor \U$9084 ( \9894 , \9888 , \9892 , \9893 );
xor \U$9085 ( \9895 , \9887 , \9894 );
and \U$9086 ( \9896 , \9859 , \9895 );
xor \U$9087 ( \9897 , \9692 , \9700 );
xor \U$9088 ( \9898 , \9896 , \9897 );
nand \U$9089 ( \9899 , \9035_nG2a09 , \8944 );
or \U$9090 ( \9900 , \8875 , \8924_nG2ae9 );
nand \U$9091 ( \9901 , \9900 , \9046 );
and \U$9092 ( \9902 , \9899 , \9901 );
and \U$9093 ( \9903 , \9390 , \8924_nG2ae9 );
and \U$9094 ( \9904 , \9035_nG2a09 , \9392 );
nor \U$9095 ( \9905 , \9902 , \9903 , \9904 );
nand \U$9096 ( \9906 , \8857_nG2bf3 , \9119 );
or \U$9097 ( \9907 , \9057 , \8770_nG2cf7 );
nand \U$9098 ( \9908 , \9907 , \9223 );
and \U$9099 ( \9909 , \9906 , \9908 );
and \U$9100 ( \9910 , \9218 , \8770_nG2cf7 );
and \U$9101 ( \9911 , \8857_nG2bf3 , \9122 );
nor \U$9102 ( \9912 , \9909 , \9910 , \9911 );
xor \U$9103 ( \9913 , \9905 , \9912 );
nand \U$9104 ( \9914 , \9289_nG290d , \8775 );
or \U$9105 ( \9915 , \8672 , \9345_nG282e );
nand \U$9106 ( \9916 , \9915 , \8781 );
and \U$9107 ( \9917 , \9914 , \9916 );
and \U$9108 ( \9918 , \8777 , \9345_nG282e );
and \U$9109 ( \9919 , \9289_nG290d , \8866 );
nor \U$9110 ( \9920 , \9917 , \9918 , \9919 );
and \U$9111 ( \9921 , \9913 , \9920 );
and \U$9112 ( \9922 , \9905 , \9912 );
or \U$9113 ( \9923 , \9921 , \9922 );
not \U$9114 ( \9924 , \9923 );
or \U$9115 ( \9925 , \9813 , \8469 );
or \U$9116 ( \9926 , \8468_nG310a , \9691 );
or \U$9117 ( \9927 , \8563_nG3003 , \9690 );
nand \U$9118 ( \9928 , \9925 , \9926 , \9927 );
not \U$9119 ( \9929 , \8730_nG2df7 );
or \U$9120 ( \9930 , \9364 , \9929 );
or \U$9121 ( \9931 , \9236 , \9694 );
or \U$9122 ( \9932 , \9361 , \9929 );
or \U$9123 ( \9933 , \9234 , \8658_nG2ee1 );
nand \U$9124 ( \9934 , \9933 , \9519 );
nand \U$9125 ( \9935 , \9932 , \9934 );
nand \U$9126 ( \9936 , \9930 , \9931 , \9935 );
and \U$9127 ( \9937 , \9928 , \9936 );
xor \U$9128 ( \9938 , \9924 , \9937 );
not \U$9129 ( \9939 , \9637_nG26ac );
or \U$9130 ( \9940 , \8579 , \9939 );
and \U$9131 ( \9941 , \8623 , \9476_nG2758 );
nand \U$9132 ( \9942 , \9637_nG26ac , \8575 );
or \U$9133 ( \9943 , \8535 , \9476_nG2758 );
nand \U$9134 ( \9944 , \9943 , \8627 );
and \U$9135 ( \9945 , \9942 , \9944 );
nor \U$9136 ( \9946 , \9941 , \9945 );
nand \U$9137 ( \9947 , \9940 , \9946 );
and \U$9138 ( \9948 , RIb558988_490, \7900 );
and \U$9139 ( \9949 , RIb558c58_496, \7955 );
and \U$9140 ( \9950 , \7943 , RIb558cd0_497);
and \U$9141 ( \9951 , RIb558d48_498, \7945 );
nor \U$9142 ( \9952 , \9950 , \9951 );
and \U$9143 ( \9953 , \7953 , RIb558a00_491);
and \U$9144 ( \9954 , RIb558910_489, \7950 );
nor \U$9145 ( \9955 , \9953 , \9954 );
and \U$9146 ( \9956 , \7917 , RIb558898_488);
and \U$9147 ( \9957 , RIb558820_487, \7921 );
nor \U$9148 ( \9958 , \9956 , \9957 );
and \U$9149 ( \9959 , \8462 , RIb5587a8_486);
and \U$9150 ( \9960 , RIb558af0_493, \7914 );
nor \U$9151 ( \9961 , \9959 , \9960 );
nand \U$9152 ( \9962 , \9952 , \9955 , \9958 , \9961 );
nor \U$9153 ( \9963 , \9948 , \9949 , \9962 );
and \U$9154 ( \9964 , \7936 , RIb558e38_500);
and \U$9155 ( \9965 , RIb558dc0_499, \7938 );
nor \U$9156 ( \9966 , \9964 , \9965 );
and \U$9157 ( \9967 , \7948 , RIb558eb0_501);
and \U$9158 ( \9968 , RIb558a78_492, \7906 );
nor \U$9159 ( \9969 , \9967 , \9968 );
and \U$9160 ( \9970 , \7926 , RIb558be0_495);
and \U$9161 ( \9971 , RIb558b68_494, \7910 );
nor \U$9162 ( \9972 , \9970 , \9971 );
nand \U$9163 ( \9973 , \9963 , \9966 , \9969 , \9972 );
_DC g24b2 ( \9974_nG24b2 , \9973 , \8467 );
not \U$9164 ( \9975 , \9974_nG24b2 );
nor \U$9165 ( \9976 , \8437 , \9975 );
xor \U$9166 ( \9977 , \9947 , \9976 );
not \U$9167 ( \9978 , \9679_nG25e2 );
or \U$9168 ( \9979 , \8522 , \9978 );
not \U$9169 ( \9980 , \9886_nG2554 );
or \U$9170 ( \9981 , \9980 , \8516 );
or \U$9171 ( \9982 , \8513 , \9978 );
or \U$9172 ( \9983 , \8481 , \9886_nG2554 );
nand \U$9173 ( \9984 , \9983 , \8518 );
nand \U$9174 ( \9985 , \9982 , \9984 );
nand \U$9175 ( \9986 , \9979 , \9981 , \9985 );
and \U$9176 ( \9987 , \9977 , \9986 );
and \U$9177 ( \9988 , \9947 , \9976 );
or \U$9178 ( \9989 , \9987 , \9988 );
and \U$9179 ( \9990 , \9938 , \9989 );
and \U$9180 ( \9991 , \9924 , \9937 );
or \U$9181 ( \9992 , \9990 , \9991 );
and \U$9182 ( \9993 , \9898 , \9992 );
and \U$9183 ( \9994 , \9896 , \9897 );
or \U$9184 ( \9995 , \9993 , \9994 );
or \U$9185 ( \9996 , \9894 , \9887 );
not \U$9186 ( \9997 , \9828 );
or \U$9187 ( \9998 , \9997 , \9801 );
not \U$9188 ( \9999 , \9801 );
or \U$9189 ( \10000 , \9828 , \9999 );
nand \U$9190 ( \10001 , \9996 , \9998 , \10000 );
xor \U$9191 ( \10002 , \9769 , \9775 );
and \U$9192 ( \10003 , \10001 , \10002 );
xor \U$9193 ( \10004 , \9995 , \10003 );
xor \U$9194 ( \10005 , \9713 , \9754 );
xor \U$9195 ( \10006 , \10005 , \9762 );
and \U$9196 ( \10007 , \10004 , \10006 );
and \U$9197 ( \10008 , \9995 , \10003 );
or \U$9198 ( \10009 , \10007 , \10008 );
and \U$9199 ( \10010 , \9856 , \10009 );
and \U$9200 ( \10011 , \9850 , \9855 );
or \U$9201 ( \10012 , \10010 , \10011 );
xor \U$9202 ( \10013 , \9747 , \9838 );
xor \U$9203 ( \10014 , \10013 , \9845 );
xor \U$9204 ( \10015 , \10012 , \10014 );
xor \U$9205 ( \10016 , \10001 , \10002 );
not \U$9206 ( \10017 , \9808 );
xor \U$9207 ( \10018 , \9816 , \9826 );
not \U$9208 ( \10019 , \10018 );
or \U$9209 ( \10020 , \10017 , \10019 );
or \U$9210 ( \10021 , \10018 , \9808 );
nand \U$9211 ( \10022 , \10020 , \10021 );
nand \U$9212 ( \10023 , \9345_nG282e , \8775 );
or \U$9213 ( \10024 , \8672 , \9476_nG2758 );
nand \U$9214 ( \10025 , \10024 , \8781 );
and \U$9215 ( \10026 , \10023 , \10025 );
and \U$9216 ( \10027 , \8777 , \9476_nG2758 );
and \U$9217 ( \10028 , \9345_nG282e , \8866 );
nor \U$9218 ( \10029 , \10026 , \10027 , \10028 );
nand \U$9219 ( \10030 , \9289_nG290d , \8944 );
or \U$9220 ( \10031 , \8875 , \9035_nG2a09 );
nand \U$9221 ( \10032 , \10031 , \9046 );
and \U$9222 ( \10033 , \10030 , \10032 );
and \U$9223 ( \10034 , \9390 , \9035_nG2a09 );
and \U$9224 ( \10035 , \9289_nG290d , \9392 );
nor \U$9225 ( \10036 , \10033 , \10034 , \10035 );
xor \U$9226 ( \10037 , \10029 , \10036 );
and \U$9227 ( \10038 , \9679_nG25e2 , \8578 );
and \U$9228 ( \10039 , \8623 , \9637_nG26ac );
nand \U$9229 ( \10040 , \9679_nG25e2 , \8575 );
or \U$9230 ( \10041 , \8535 , \9637_nG26ac );
nand \U$9231 ( \10042 , \10041 , \8627 );
and \U$9232 ( \10043 , \10040 , \10042 );
nor \U$9233 ( \10044 , \10038 , \10039 , \10043 );
and \U$9234 ( \10045 , \10037 , \10044 );
and \U$9235 ( \10046 , \10029 , \10036 );
or \U$9236 ( \10047 , \10045 , \10046 );
nand \U$9237 ( \10048 , \8770_nG2cf7 , \9360 );
or \U$9238 ( \10049 , \9234 , \8730_nG2df7 );
nand \U$9239 ( \10050 , \10049 , \9519 );
and \U$9240 ( \10051 , \10048 , \10050 );
and \U$9241 ( \10052 , \9522 , \8730_nG2df7 );
and \U$9242 ( \10053 , \8770_nG2cf7 , \9363 );
nor \U$9243 ( \10054 , \10051 , \10052 , \10053 );
and \U$9244 ( \10055 , \8564 , \9810 );
and \U$9245 ( \10056 , \9689 , \9236 );
and \U$9246 ( \10057 , \8563_nG3003 , \9814 );
nor \U$9247 ( \10058 , \10055 , \10056 , \10057 );
xor \U$9248 ( \10059 , \10054 , \10058 );
nand \U$9249 ( \10060 , \8924_nG2ae9 , \9119 );
or \U$9250 ( \10061 , \9057 , \8857_nG2bf3 );
nand \U$9251 ( \10062 , \10061 , \9223 );
and \U$9252 ( \10063 , \10060 , \10062 );
and \U$9253 ( \10064 , \9218 , \8857_nG2bf3 );
and \U$9254 ( \10065 , \8924_nG2ae9 , \9122 );
nor \U$9255 ( \10066 , \10063 , \10064 , \10065 );
and \U$9256 ( \10067 , \10059 , \10066 );
and \U$9257 ( \10068 , \10054 , \10058 );
or \U$9258 ( \10069 , \10067 , \10068 );
nor \U$9259 ( \10070 , \10047 , \10069 );
and \U$9260 ( \10071 , \10022 , \10070 );
xor \U$9261 ( \10072 , \10016 , \10071 );
xor \U$9262 ( \10073 , \9896 , \9897 );
xor \U$9263 ( \10074 , \10073 , \9992 );
and \U$9264 ( \10075 , \10072 , \10074 );
and \U$9265 ( \10076 , \10016 , \10071 );
or \U$9266 ( \10077 , \10075 , \10076 );
not \U$9267 ( \10078 , \9832 );
xor \U$9268 ( \10079 , \9829 , \9776 );
not \U$9269 ( \10080 , \10079 );
or \U$9270 ( \10081 , \10078 , \10080 );
or \U$9271 ( \10082 , \10079 , \9832 );
nand \U$9272 ( \10083 , \10081 , \10082 );
xor \U$9273 ( \10084 , \10077 , \10083 );
xor \U$9274 ( \10085 , \9995 , \10003 );
xor \U$9275 ( \10086 , \10085 , \10006 );
and \U$9276 ( \10087 , \10084 , \10086 );
and \U$9277 ( \10088 , \10077 , \10083 );
or \U$9278 ( \10089 , \10087 , \10088 );
xor \U$9279 ( \10090 , \9850 , \9855 );
xor \U$9280 ( \10091 , \10090 , \10009 );
xor \U$9281 ( \10092 , \10089 , \10091 );
xor \U$9282 ( \10093 , \10077 , \10083 );
xor \U$9283 ( \10094 , \10093 , \10086 );
and \U$9284 ( \10095 , \9886_nG2554 , \8521 );
or \U$9285 ( \10096 , \8481 , \9974_nG24b2 );
nand \U$9286 ( \10097 , \10096 , \8518 );
nand \U$9287 ( \10098 , \9886_nG2554 , \8514 );
and \U$9288 ( \10099 , \10097 , \10098 );
and \U$9289 ( \10100 , \9974_nG24b2 , \8663 );
nor \U$9290 ( \10101 , \10095 , \10099 , \10100 );
and \U$9291 ( \10102 , RIb55a008_538, \7921 );
and \U$9292 ( \10103 , RIb55a1e8_542, \7953 );
and \U$9293 ( \10104 , \7955 , RIb55a440_547);
and \U$9294 ( \10105 , RIb55a3c8_546, \7926 );
nor \U$9295 ( \10106 , \10104 , \10105 );
and \U$9296 ( \10107 , \7938 , RIb55a5a8_550);
and \U$9297 ( \10108 , RIb55a170_541, \7900 );
nor \U$9298 ( \10109 , \10107 , \10108 );
and \U$9299 ( \10110 , \7948 , RIb55a698_552);
and \U$9300 ( \10111 , RIb55a620_551, \7936 );
nor \U$9301 ( \10112 , \10110 , \10111 );
and \U$9302 ( \10113 , \7906 , RIb55a260_543);
and \U$9303 ( \10114 , RIb55a350_545, \7910 );
nor \U$9304 ( \10115 , \10113 , \10114 );
nand \U$9305 ( \10116 , \10106 , \10109 , \10112 , \10115 );
nor \U$9306 ( \10117 , \10102 , \10103 , \10116 );
and \U$9307 ( \10118 , \7943 , RIb55a4b8_548);
and \U$9308 ( \10119 , RIb55a080_539, \7917 );
nor \U$9309 ( \10120 , \10118 , \10119 );
and \U$9310 ( \10121 , \7914 , RIb55a2d8_544);
and \U$9311 ( \10122 , RIb55a0f8_540, \7950 );
nor \U$9312 ( \10123 , \10121 , \10122 );
and \U$9313 ( \10124 , \8462 , RIb559f90_537);
and \U$9314 ( \10125 , RIb55a530_549, \7945 );
nor \U$9315 ( \10126 , \10124 , \10125 );
nand \U$9316 ( \10127 , \10117 , \10120 , \10123 , \10126 );
_DC g2440 ( \10128_nG2440 , \10127 , \8467 );
nand \U$9317 ( \10129 , \10128_nG2440 , \8436 );
or \U$9318 ( \10130 , \10101 , \10129 );
not \U$9319 ( \10131 , \10069 );
or \U$9320 ( \10132 , \10131 , \10047 );
not \U$9321 ( \10133 , \10047 );
or \U$9322 ( \10134 , \10069 , \10133 );
nand \U$9323 ( \10135 , \10130 , \10132 , \10134 );
xor \U$9324 ( \10136 , \9928 , \9936 );
xor \U$9325 ( \10137 , \10135 , \10136 );
xor \U$9326 ( \10138 , \9947 , \9976 );
xor \U$9327 ( \10139 , \10138 , \9986 );
and \U$9328 ( \10140 , \10137 , \10139 );
and \U$9329 ( \10141 , \10135 , \10136 );
or \U$9330 ( \10142 , \10140 , \10141 );
xor \U$9331 ( \10143 , \9859 , \9895 );
xor \U$9332 ( \10144 , \10142 , \10143 );
xor \U$9333 ( \10145 , \10029 , \10036 );
xor \U$9334 ( \10146 , \10145 , \10044 );
xor \U$9335 ( \10147 , \10054 , \10058 );
xor \U$9336 ( \10148 , \10147 , \10066 );
xor \U$9337 ( \10149 , \10146 , \10148 );
xnor \U$9338 ( \10150 , \10129 , \10101 );
and \U$9339 ( \10151 , \10149 , \10150 );
and \U$9340 ( \10152 , \10146 , \10148 );
or \U$9341 ( \10153 , \10151 , \10152 );
xor \U$9342 ( \10154 , \9905 , \9912 );
xor \U$9343 ( \10155 , \10154 , \9920 );
xor \U$9344 ( \10156 , \10153 , \10155 );
nand \U$9345 ( \10157 , \9345_nG282e , \8944 );
or \U$9346 ( \10158 , \8875 , \9289_nG290d );
nand \U$9347 ( \10159 , \10158 , \9046 );
and \U$9348 ( \10160 , \10157 , \10159 );
and \U$9349 ( \10161 , \9390 , \9289_nG290d );
and \U$9350 ( \10162 , \9345_nG282e , \9392 );
nor \U$9351 ( \10163 , \10160 , \10161 , \10162 );
nand \U$9352 ( \10164 , \9035_nG2a09 , \9119 );
or \U$9353 ( \10165 , \9057 , \8924_nG2ae9 );
nand \U$9354 ( \10166 , \10165 , \9223 );
and \U$9355 ( \10167 , \10164 , \10166 );
and \U$9356 ( \10168 , \9218 , \8924_nG2ae9 );
and \U$9357 ( \10169 , \9035_nG2a09 , \9122 );
nor \U$9358 ( \10170 , \10167 , \10168 , \10169 );
xor \U$9359 ( \10171 , \10163 , \10170 );
nand \U$9360 ( \10172 , \9476_nG2758 , \8775 );
or \U$9361 ( \10173 , \8672 , \9637_nG26ac );
nand \U$9362 ( \10174 , \10173 , \8781 );
and \U$9363 ( \10175 , \10172 , \10174 );
and \U$9364 ( \10176 , \8777 , \9637_nG26ac );
and \U$9365 ( \10177 , \9476_nG2758 , \8866 );
nor \U$9366 ( \10178 , \10175 , \10176 , \10177 );
and \U$9367 ( \10179 , \10171 , \10178 );
and \U$9368 ( \10180 , \10163 , \10170 );
or \U$9369 ( \10181 , \10179 , \10180 );
nand \U$9370 ( \10182 , \8857_nG2bf3 , \9360 );
or \U$9371 ( \10183 , \9234 , \8770_nG2cf7 );
nand \U$9372 ( \10184 , \10183 , \9519 );
and \U$9373 ( \10185 , \10182 , \10184 );
and \U$9374 ( \10186 , \9522 , \8770_nG2cf7 );
and \U$9375 ( \10187 , \8857_nG2bf3 , \9363 );
nor \U$9376 ( \10188 , \10185 , \10186 , \10187 );
not \U$9377 ( \10189 , \10188 );
or \U$9378 ( \10190 , \9813 , \9236 );
or \U$9379 ( \10191 , \8658_nG2ee1 , \9691 );
or \U$9380 ( \10192 , \8730_nG2df7 , \9690 );
nand \U$9381 ( \10193 , \10190 , \10191 , \10192 );
nand \U$9382 ( \10194 , \10189 , \10193 );
xor \U$9383 ( \10195 , \10181 , \10194 );
and \U$9384 ( \10196 , \9974_nG24b2 , \8521 );
or \U$9385 ( \10197 , \8481 , \10128_nG2440 );
nand \U$9386 ( \10198 , \10197 , \8518 );
nand \U$9387 ( \10199 , \9974_nG24b2 , \8514 );
and \U$9388 ( \10200 , \10198 , \10199 );
and \U$9389 ( \10201 , \10128_nG2440 , \8663 );
nor \U$9390 ( \10202 , \10196 , \10200 , \10201 );
and \U$9391 ( \10203 , \9886_nG2554 , \8578 );
and \U$9392 ( \10204 , \8623 , \9679_nG25e2 );
nand \U$9393 ( \10205 , \9886_nG2554 , \8575 );
or \U$9394 ( \10206 , \8535 , \9679_nG25e2 );
nand \U$9395 ( \10207 , \10206 , \8627 );
and \U$9396 ( \10208 , \10205 , \10207 );
nor \U$9397 ( \10209 , \10203 , \10204 , \10208 );
and \U$9398 ( \10210 , \10202 , \10209 );
not \U$9399 ( \10211 , \10210 );
and \U$9400 ( \10212 , RIb559978_524, \7900 );
and \U$9401 ( \10213 , RIb559c48_530, \7955 );
and \U$9402 ( \10214 , \7943 , RIb559cc0_531);
and \U$9403 ( \10215 , RIb559d38_532, \7945 );
nor \U$9404 ( \10216 , \10214 , \10215 );
and \U$9405 ( \10217 , \7950 , RIb559900_523);
and \U$9406 ( \10218 , RIb559b58_528, \7910 );
nor \U$9407 ( \10219 , \10217 , \10218 );
and \U$9408 ( \10220 , \7917 , RIb559888_522);
and \U$9409 ( \10221 , RIb559810_521, \7921 );
nor \U$9410 ( \10222 , \10220 , \10221 );
and \U$9411 ( \10223 , \8462 , RIb559798_520);
and \U$9412 ( \10224 , RIb559ae0_527, \7914 );
nor \U$9413 ( \10225 , \10223 , \10224 );
nand \U$9414 ( \10226 , \10216 , \10219 , \10222 , \10225 );
nor \U$9415 ( \10227 , \10212 , \10213 , \10226 );
and \U$9416 ( \10228 , \7906 , RIb559a68_526);
and \U$9417 ( \10229 , RIb559bd0_529, \7926 );
nor \U$9418 ( \10230 , \10228 , \10229 );
and \U$9419 ( \10231 , \7948 , RIb559ea0_535);
and \U$9420 ( \10232 , RIb5599f0_525, \7953 );
nor \U$9421 ( \10233 , \10231 , \10232 );
and \U$9422 ( \10234 , \7936 , RIb559e28_534);
and \U$9423 ( \10235 , RIb559db0_533, \7938 );
nor \U$9424 ( \10236 , \10234 , \10235 );
nand \U$9425 ( \10237 , \10227 , \10230 , \10233 , \10236 );
_DC g23be ( \10238_nG23be , \10237 , \8467 );
nand \U$9426 ( \10239 , \10238_nG23be , \8436 );
not \U$9427 ( \10240 , \10239 );
and \U$9428 ( \10241 , \10211 , \10240 );
nor \U$9429 ( \10242 , \10202 , \10209 );
nor \U$9430 ( \10243 , \10241 , \10242 );
and \U$9431 ( \10244 , \10195 , \10243 );
and \U$9432 ( \10245 , \10181 , \10194 );
or \U$9433 ( \10246 , \10244 , \10245 );
and \U$9434 ( \10247 , \10156 , \10246 );
and \U$9435 ( \10248 , \10153 , \10155 );
or \U$9436 ( \10249 , \10247 , \10248 );
not \U$9437 ( \10250 , \10249 );
and \U$9438 ( \10251 , \10144 , \10250 );
and \U$9439 ( \10252 , \10142 , \10143 );
or \U$9440 ( \10253 , \10251 , \10252 );
xor \U$9441 ( \10254 , \10022 , \10070 );
xor \U$9442 ( \10255 , \9924 , \9937 );
xor \U$9443 ( \10256 , \10255 , \9989 );
and \U$9444 ( \10257 , \10254 , \10256 );
xor \U$9445 ( \10258 , \10253 , \10257 );
xor \U$9446 ( \10259 , \10016 , \10071 );
xor \U$9447 ( \10260 , \10259 , \10074 );
and \U$9448 ( \10261 , \10258 , \10260 );
and \U$9449 ( \10262 , \10253 , \10257 );
or \U$9450 ( \10263 , \10261 , \10262 );
xor \U$9451 ( \10264 , \10094 , \10263 );
xor \U$9452 ( \10265 , \10253 , \10257 );
xor \U$9453 ( \10266 , \10265 , \10260 );
xor \U$9454 ( \10267 , \10254 , \10256 );
xor \U$9455 ( \10268 , \10142 , \10143 );
xor \U$9456 ( \10269 , \10268 , \10250 );
and \U$9457 ( \10270 , \10267 , \10269 );
xor \U$9458 ( \10271 , \10163 , \10170 );
xor \U$9459 ( \10272 , \10271 , \10178 );
not \U$9460 ( \10273 , \10272 );
not \U$9461 ( \10274 , \10239 );
nor \U$9462 ( \10275 , \10210 , \10242 );
not \U$9463 ( \10276 , \10275 );
or \U$9464 ( \10277 , \10274 , \10276 );
or \U$9465 ( \10278 , \10275 , \10239 );
nand \U$9466 ( \10279 , \10277 , \10278 );
nand \U$9467 ( \10280 , \10273 , \10279 );
nand \U$9468 ( \10281 , \8924_nG2ae9 , \9360 );
or \U$9469 ( \10282 , \9234 , \8857_nG2bf3 );
nand \U$9470 ( \10283 , \10282 , \9519 );
and \U$9471 ( \10284 , \10281 , \10283 );
and \U$9472 ( \10285 , \9522 , \8857_nG2bf3 );
and \U$9473 ( \10286 , \8924_nG2ae9 , \9363 );
nor \U$9474 ( \10287 , \10284 , \10285 , \10286 );
and \U$9475 ( \10288 , \9929 , \9810 );
not \U$9476 ( \10289 , \8770_nG2cf7 );
and \U$9477 ( \10290 , \9689 , \10289 );
and \U$9478 ( \10291 , \8730_nG2df7 , \9814 );
nor \U$9479 ( \10292 , \10288 , \10290 , \10291 );
xor \U$9480 ( \10293 , \10287 , \10292 );
nand \U$9481 ( \10294 , \9289_nG290d , \9119 );
or \U$9482 ( \10295 , \9057 , \9035_nG2a09 );
nand \U$9483 ( \10296 , \10295 , \9223 );
and \U$9484 ( \10297 , \10294 , \10296 );
and \U$9485 ( \10298 , \9218 , \9035_nG2a09 );
and \U$9486 ( \10299 , \9289_nG290d , \9122 );
nor \U$9487 ( \10300 , \10297 , \10298 , \10299 );
and \U$9488 ( \10301 , \10293 , \10300 );
and \U$9489 ( \10302 , \10287 , \10292 );
or \U$9490 ( \10303 , \10301 , \10302 );
not \U$9491 ( \10304 , \10303 );
nand \U$9492 ( \10305 , \9637_nG26ac , \8775 );
or \U$9493 ( \10306 , \8672 , \9679_nG25e2 );
nand \U$9494 ( \10307 , \10306 , \8781 );
and \U$9495 ( \10308 , \10305 , \10307 );
and \U$9496 ( \10309 , \8777 , \9679_nG25e2 );
and \U$9497 ( \10310 , \9637_nG26ac , \8866 );
nor \U$9498 ( \10311 , \10308 , \10309 , \10310 );
nand \U$9499 ( \10312 , \9476_nG2758 , \8944 );
or \U$9500 ( \10313 , \8875 , \9345_nG282e );
nand \U$9501 ( \10314 , \10313 , \9046 );
and \U$9502 ( \10315 , \10312 , \10314 );
and \U$9503 ( \10316 , \9390 , \9345_nG282e );
and \U$9504 ( \10317 , \9476_nG2758 , \9392 );
nor \U$9505 ( \10318 , \10315 , \10316 , \10317 );
xor \U$9506 ( \10319 , \10311 , \10318 );
and \U$9507 ( \10320 , \9974_nG24b2 , \8578 );
and \U$9508 ( \10321 , \8623 , \9886_nG2554 );
nand \U$9509 ( \10322 , \9974_nG24b2 , \8575 );
or \U$9510 ( \10323 , \8535 , \9886_nG2554 );
nand \U$9511 ( \10324 , \10323 , \8627 );
and \U$9512 ( \10325 , \10322 , \10324 );
nor \U$9513 ( \10326 , \10320 , \10321 , \10325 );
and \U$9514 ( \10327 , \10319 , \10326 );
and \U$9515 ( \10328 , \10311 , \10318 );
or \U$9516 ( \10329 , \10327 , \10328 );
not \U$9517 ( \10330 , \10329 );
nand \U$9518 ( \10331 , \10304 , \10330 );
xor \U$9519 ( \10332 , \10280 , \10331 );
xor \U$9520 ( \10333 , \10146 , \10148 );
xor \U$9521 ( \10334 , \10333 , \10150 );
and \U$9522 ( \10335 , \10332 , \10334 );
and \U$9523 ( \10336 , \10280 , \10331 );
or \U$9524 ( \10337 , \10335 , \10336 );
not \U$9525 ( \10338 , \10337 );
xor \U$9526 ( \10339 , \10135 , \10136 );
xor \U$9527 ( \10340 , \10339 , \10139 );
nor \U$9528 ( \10341 , \10338 , \10340 );
xor \U$9529 ( \10342 , \10153 , \10155 );
xor \U$9530 ( \10343 , \10342 , \10246 );
or \U$9531 ( \10344 , \10341 , \10343 );
not \U$9532 ( \10345 , \10337 );
nand \U$9533 ( \10346 , \10345 , \10340 );
nand \U$9534 ( \10347 , \10344 , \10346 );
xor \U$9535 ( \10348 , \10142 , \10143 );
xor \U$9536 ( \10349 , \10348 , \10250 );
and \U$9537 ( \10350 , \10347 , \10349 );
and \U$9538 ( \10351 , \10267 , \10347 );
or \U$9539 ( \10352 , \10270 , \10350 , \10351 );
xor \U$9540 ( \10353 , \10266 , \10352 );
xor \U$9541 ( \10354 , \10142 , \10143 );
xor \U$9542 ( \10355 , \10354 , \10250 );
xor \U$9543 ( \10356 , \10267 , \10347 );
xor \U$9544 ( \10357 , \10355 , \10356 );
not \U$9545 ( \10358 , \10340 );
not \U$9546 ( \10359 , \10343 );
or \U$9547 ( \10360 , \10358 , \10359 );
or \U$9548 ( \10361 , \10343 , \10340 );
nand \U$9549 ( \10362 , \10360 , \10361 );
not \U$9550 ( \10363 , \10362 );
not \U$9551 ( \10364 , \10337 );
and \U$9552 ( \10365 , \10363 , \10364 );
and \U$9553 ( \10366 , \10362 , \10337 );
nor \U$9554 ( \10367 , \10365 , \10366 );
not \U$9555 ( \10368 , \10279 );
not \U$9556 ( \10369 , \10272 );
and \U$9557 ( \10370 , \10368 , \10369 );
and \U$9558 ( \10371 , \10279 , \10272 );
nor \U$9559 ( \10372 , \10370 , \10371 );
not \U$9560 ( \10373 , \10372 );
and \U$9561 ( \10374 , \10128_nG2440 , \8521 );
or \U$9562 ( \10375 , \8481 , \10238_nG23be );
nand \U$9563 ( \10376 , \10375 , \8518 );
nand \U$9564 ( \10377 , \10128_nG2440 , \8514 );
and \U$9565 ( \10378 , \10376 , \10377 );
and \U$9566 ( \10379 , \10238_nG23be , \8663 );
nor \U$9567 ( \10380 , \10374 , \10378 , \10379 );
and \U$9568 ( \10381 , RIb55aad0_561, \7914 );
and \U$9569 ( \10382 , RIb55aa58_560, \7906 );
and \U$9570 ( \10383 , \7953 , RIb55a9e0_559);
and \U$9571 ( \10384 , RIb55a8f0_557, \7950 );
nor \U$9572 ( \10385 , \10383 , \10384 );
and \U$9573 ( \10386 , \7948 , RIb55ae90_569);
and \U$9574 ( \10387 , RIb55ae18_568, \7936 );
nor \U$9575 ( \10388 , \10386 , \10387 );
and \U$9576 ( \10389 , \7917 , RIb55a878_556);
and \U$9577 ( \10390 , RIb55a800_555, \7921 );
nor \U$9578 ( \10391 , \10389 , \10390 );
and \U$9579 ( \10392 , \7938 , RIb55ada0_567);
and \U$9580 ( \10393 , RIb55a968_558, \7900 );
nor \U$9581 ( \10394 , \10392 , \10393 );
nand \U$9582 ( \10395 , \10385 , \10388 , \10391 , \10394 );
nor \U$9583 ( \10396 , \10381 , \10382 , \10395 );
and \U$9584 ( \10397 , \7926 , RIb55abc0_563);
and \U$9585 ( \10398 , RIb55ab48_562, \7910 );
nor \U$9586 ( \10399 , \10397 , \10398 );
and \U$9587 ( \10400 , \8462 , RIb55a788_554);
and \U$9588 ( \10401 , RIb55ad28_566, \7945 );
nor \U$9589 ( \10402 , \10400 , \10401 );
and \U$9590 ( \10403 , \7943 , RIb55acb0_565);
and \U$9591 ( \10404 , RIb55ac38_564, \7955 );
nor \U$9592 ( \10405 , \10403 , \10404 );
nand \U$9593 ( \10406 , \10396 , \10399 , \10402 , \10405 );
_DC g236e ( \10407_nG236e , \10406 , \8467 );
nand \U$9594 ( \10408 , \10407_nG236e , \8436 );
or \U$9595 ( \10409 , \10380 , \10408 );
or \U$9596 ( \10410 , \10304 , \10329 );
or \U$9597 ( \10411 , \10303 , \10330 );
nand \U$9598 ( \10412 , \10409 , \10410 , \10411 );
nand \U$9599 ( \10413 , \10373 , \10412 );
xor \U$9600 ( \10414 , \10181 , \10194 );
xor \U$9601 ( \10415 , \10414 , \10243 );
xor \U$9602 ( \10416 , \10413 , \10415 );
xor \U$9603 ( \10417 , \10311 , \10318 );
xor \U$9604 ( \10418 , \10417 , \10326 );
xor \U$9605 ( \10419 , \10287 , \10292 );
xor \U$9606 ( \10420 , \10419 , \10300 );
xor \U$9607 ( \10421 , \10418 , \10420 );
xnor \U$9608 ( \10422 , \10408 , \10380 );
and \U$9609 ( \10423 , \10421 , \10422 );
and \U$9610 ( \10424 , \10418 , \10420 );
or \U$9611 ( \10425 , \10423 , \10424 );
not \U$9612 ( \10426 , \10188 );
not \U$9613 ( \10427 , \10193 );
and \U$9614 ( \10428 , \10426 , \10427 );
and \U$9615 ( \10429 , \10188 , \10193 );
nor \U$9616 ( \10430 , \10428 , \10429 );
xor \U$9617 ( \10431 , \10425 , \10430 );
nand \U$9618 ( \10432 , \9637_nG26ac , \8944 );
or \U$9619 ( \10433 , \8875 , \9476_nG2758 );
nand \U$9620 ( \10434 , \10433 , \9046 );
and \U$9621 ( \10435 , \10432 , \10434 );
and \U$9622 ( \10436 , \9390 , \9476_nG2758 );
and \U$9623 ( \10437 , \9637_nG26ac , \9392 );
nor \U$9624 ( \10438 , \10435 , \10436 , \10437 );
nand \U$9625 ( \10439 , \9345_nG282e , \9119 );
or \U$9626 ( \10440 , \9057 , \9289_nG290d );
nand \U$9627 ( \10441 , \10440 , \9223 );
and \U$9628 ( \10442 , \10439 , \10441 );
and \U$9629 ( \10443 , \9218 , \9289_nG290d );
and \U$9630 ( \10444 , \9345_nG282e , \9122 );
nor \U$9631 ( \10445 , \10442 , \10443 , \10444 );
xor \U$9632 ( \10446 , \10438 , \10445 );
nand \U$9633 ( \10447 , \9679_nG25e2 , \8775 );
or \U$9634 ( \10448 , \8672 , \9886_nG2554 );
nand \U$9635 ( \10449 , \10448 , \8781 );
and \U$9636 ( \10450 , \10447 , \10449 );
and \U$9637 ( \10451 , \8777 , \9886_nG2554 );
and \U$9638 ( \10452 , \9679_nG25e2 , \8866 );
nor \U$9639 ( \10453 , \10450 , \10451 , \10452 );
and \U$9640 ( \10454 , \10446 , \10453 );
and \U$9641 ( \10455 , \10438 , \10445 );
or \U$9642 ( \10456 , \10454 , \10455 );
nand \U$9643 ( \10457 , \9035_nG2a09 , \9360 );
or \U$9644 ( \10458 , \9234 , \8924_nG2ae9 );
nand \U$9645 ( \10459 , \10458 , \9519 );
and \U$9646 ( \10460 , \10457 , \10459 );
and \U$9647 ( \10461 , \9522 , \8924_nG2ae9 );
and \U$9648 ( \10462 , \9035_nG2a09 , \9363 );
nor \U$9649 ( \10463 , \10460 , \10461 , \10462 );
not \U$9650 ( \10464 , \10463 );
or \U$9651 ( \10465 , \9813 , \10289 );
or \U$9652 ( \10466 , \8770_nG2cf7 , \9691 );
or \U$9653 ( \10467 , \8857_nG2bf3 , \9690 );
nand \U$9654 ( \10468 , \10465 , \10466 , \10467 );
nand \U$9655 ( \10469 , \10464 , \10468 );
xor \U$9656 ( \10470 , \10456 , \10469 );
and \U$9657 ( \10471 , \10128_nG2440 , \8578 );
and \U$9658 ( \10472 , \8623 , \9974_nG24b2 );
nand \U$9659 ( \10473 , \10128_nG2440 , \8575 );
or \U$9660 ( \10474 , \8535 , \9974_nG24b2 );
nand \U$9661 ( \10475 , \10474 , \8627 );
and \U$9662 ( \10476 , \10473 , \10475 );
nor \U$9663 ( \10477 , \10471 , \10472 , \10476 );
and \U$9664 ( \10478 , RIb55aff8_572, \7921 );
and \U$9665 ( \10479 , RIb55b2c8_578, \7914 );
and \U$9666 ( \10480 , \7955 , RIb55b430_581);
and \U$9667 ( \10481 , RIb55b3b8_580, \7926 );
nor \U$9668 ( \10482 , \10480 , \10481 );
and \U$9669 ( \10483 , \7938 , RIb55b598_584);
and \U$9670 ( \10484 , RIb55b160_575, \7900 );
nor \U$9671 ( \10485 , \10483 , \10484 );
and \U$9672 ( \10486 , \7948 , RIb55b688_586);
and \U$9673 ( \10487 , RIb55b610_585, \7936 );
nor \U$9674 ( \10488 , \10486 , \10487 );
and \U$9675 ( \10489 , \7906 , RIb55b250_577);
and \U$9676 ( \10490 , RIb55b340_579, \7910 );
nor \U$9677 ( \10491 , \10489 , \10490 );
nand \U$9678 ( \10492 , \10482 , \10485 , \10488 , \10491 );
nor \U$9679 ( \10493 , \10478 , \10479 , \10492 );
and \U$9680 ( \10494 , \7943 , RIb55b4a8_582);
and \U$9681 ( \10495 , RIb55b1d8_576, \7953 );
nor \U$9682 ( \10496 , \10494 , \10495 );
and \U$9683 ( \10497 , \7950 , RIb55b0e8_574);
and \U$9684 ( \10498 , RIb55b070_573, \7917 );
nor \U$9685 ( \10499 , \10497 , \10498 );
and \U$9686 ( \10500 , \8462 , RIb55af80_571);
and \U$9687 ( \10501 , RIb55b520_583, \7945 );
nor \U$9688 ( \10502 , \10500 , \10501 );
nand \U$9689 ( \10503 , \10493 , \10496 , \10499 , \10502 );
_DC g2250 ( \10504_nG2250 , \10503 , \8467 );
nand \U$9690 ( \10505 , \10504_nG2250 , \8436 );
xor \U$9691 ( \10506 , \10477 , \10505 );
and \U$9692 ( \10507 , \10238_nG23be , \8521 );
or \U$9693 ( \10508 , \8481 , \10407_nG236e );
nand \U$9694 ( \10509 , \10508 , \8518 );
nand \U$9695 ( \10510 , \10238_nG23be , \8514 );
and \U$9696 ( \10511 , \10509 , \10510 );
and \U$9697 ( \10512 , \10407_nG236e , \8663 );
nor \U$9698 ( \10513 , \10507 , \10511 , \10512 );
and \U$9699 ( \10514 , \10506 , \10513 );
and \U$9700 ( \10515 , \10477 , \10505 );
or \U$9701 ( \10516 , \10514 , \10515 );
and \U$9702 ( \10517 , \10470 , \10516 );
and \U$9703 ( \10518 , \10456 , \10469 );
or \U$9704 ( \10519 , \10517 , \10518 );
and \U$9705 ( \10520 , \10431 , \10519 );
and \U$9706 ( \10521 , \10425 , \10430 );
or \U$9707 ( \10522 , \10520 , \10521 );
and \U$9708 ( \10523 , \10416 , \10522 );
and \U$9709 ( \10524 , \10413 , \10415 );
or \U$9710 ( \10525 , \10523 , \10524 );
nor \U$9711 ( \10526 , \10367 , \10525 );
xor \U$9712 ( \10527 , \10357 , \10526 );
and \U$9713 ( \10528 , \10367 , \10525 );
nor \U$9714 ( \10529 , \10528 , \10526 );
xor \U$9715 ( \10530 , \10413 , \10415 );
xor \U$9716 ( \10531 , \10530 , \10522 );
xor \U$9717 ( \10532 , \10280 , \10331 );
xor \U$9718 ( \10533 , \10532 , \10334 );
nor \U$9719 ( \10534 , \10531 , \10533 );
xor \U$9720 ( \10535 , \10529 , \10534 );
and \U$9721 ( \10536 , \10531 , \10533 );
nor \U$9722 ( \10537 , \10536 , \10534 );
nand \U$9723 ( \10538 , \9886_nG2554 , \8775 );
or \U$9724 ( \10539 , \8672 , \9974_nG24b2 );
nand \U$9725 ( \10540 , \10539 , \8781 );
and \U$9726 ( \10541 , \10538 , \10540 );
and \U$9727 ( \10542 , \8777 , \9974_nG24b2 );
and \U$9728 ( \10543 , \9886_nG2554 , \8866 );
nor \U$9729 ( \10544 , \10541 , \10542 , \10543 );
nand \U$9730 ( \10545 , \9679_nG25e2 , \8944 );
or \U$9731 ( \10546 , \8875 , \9637_nG26ac );
nand \U$9732 ( \10547 , \10546 , \9046 );
and \U$9733 ( \10548 , \10545 , \10547 );
and \U$9734 ( \10549 , \9390 , \9637_nG26ac );
and \U$9735 ( \10550 , \9679_nG25e2 , \9392 );
nor \U$9736 ( \10551 , \10548 , \10549 , \10550 );
xor \U$9737 ( \10552 , \10544 , \10551 );
and \U$9738 ( \10553 , \10238_nG23be , \8578 );
and \U$9739 ( \10554 , \8623 , \10128_nG2440 );
nand \U$9740 ( \10555 , \10238_nG23be , \8575 );
or \U$9741 ( \10556 , \8535 , \10128_nG2440 );
nand \U$9742 ( \10557 , \10556 , \8627 );
and \U$9743 ( \10558 , \10555 , \10557 );
nor \U$9744 ( \10559 , \10553 , \10554 , \10558 );
and \U$9745 ( \10560 , \10552 , \10559 );
and \U$9746 ( \10561 , \10544 , \10551 );
or \U$9747 ( \10562 , \10560 , \10561 );
nand \U$9748 ( \10563 , \9289_nG290d , \9360 );
or \U$9749 ( \10564 , \9234 , \9035_nG2a09 );
nand \U$9750 ( \10565 , \10564 , \9519 );
and \U$9751 ( \10566 , \10563 , \10565 );
and \U$9752 ( \10567 , \9522 , \9035_nG2a09 );
and \U$9753 ( \10568 , \9289_nG290d , \9363 );
nor \U$9754 ( \10569 , \10566 , \10567 , \10568 );
not \U$9755 ( \10570 , \8857_nG2bf3 );
and \U$9756 ( \10571 , \10570 , \9810 );
not \U$9757 ( \10572 , \8924_nG2ae9 );
and \U$9758 ( \10573 , \9689 , \10572 );
and \U$9759 ( \10574 , \8857_nG2bf3 , \9814 );
nor \U$9760 ( \10575 , \10571 , \10573 , \10574 );
xor \U$9761 ( \10576 , \10569 , \10575 );
nand \U$9762 ( \10577 , \9476_nG2758 , \9119 );
or \U$9763 ( \10578 , \9057 , \9345_nG282e );
nand \U$9764 ( \10579 , \10578 , \9223 );
and \U$9765 ( \10580 , \10577 , \10579 );
and \U$9766 ( \10581 , \9218 , \9345_nG282e );
and \U$9767 ( \10582 , \9476_nG2758 , \9122 );
nor \U$9768 ( \10583 , \10580 , \10581 , \10582 );
and \U$9769 ( \10584 , \10576 , \10583 );
and \U$9770 ( \10585 , \10569 , \10575 );
or \U$9771 ( \10586 , \10584 , \10585 );
xor \U$9772 ( \10587 , \10562 , \10586 );
xor \U$9773 ( \10588 , \10477 , \10505 );
xor \U$9774 ( \10589 , \10588 , \10513 );
and \U$9775 ( \10590 , \10587 , \10589 );
and \U$9776 ( \10591 , \10562 , \10586 );
or \U$9777 ( \10592 , \10590 , \10591 );
xor \U$9778 ( \10593 , \10438 , \10445 );
xor \U$9779 ( \10594 , \10593 , \10453 );
not \U$9780 ( \10595 , \10594 );
not \U$9781 ( \10596 , \10468 );
not \U$9782 ( \10597 , \10463 );
or \U$9783 ( \10598 , \10596 , \10597 );
or \U$9784 ( \10599 , \10463 , \10468 );
nand \U$9785 ( \10600 , \10598 , \10599 );
nand \U$9786 ( \10601 , \10595 , \10600 );
xor \U$9787 ( \10602 , \10592 , \10601 );
xor \U$9788 ( \10603 , \10418 , \10420 );
xor \U$9789 ( \10604 , \10603 , \10422 );
and \U$9790 ( \10605 , \10602 , \10604 );
and \U$9791 ( \10606 , \10592 , \10601 );
or \U$9792 ( \10607 , \10605 , \10606 );
not \U$9793 ( \10608 , \10372 );
not \U$9794 ( \10609 , \10412 );
and \U$9795 ( \10610 , \10608 , \10609 );
and \U$9796 ( \10611 , \10372 , \10412 );
nor \U$9797 ( \10612 , \10610 , \10611 );
xor \U$9798 ( \10613 , \10607 , \10612 );
xor \U$9799 ( \10614 , \10425 , \10430 );
xor \U$9800 ( \10615 , \10614 , \10519 );
and \U$9801 ( \10616 , \10613 , \10615 );
and \U$9802 ( \10617 , \10607 , \10612 );
or \U$9803 ( \10618 , \10616 , \10617 );
not \U$9804 ( \10619 , \10618 );
xor \U$9805 ( \10620 , \10537 , \10619 );
nand \U$9806 ( \10621 , \9345_nG282e , \9360 );
or \U$9807 ( \10622 , \9234 , \9289_nG290d );
nand \U$9808 ( \10623 , \10622 , \9519 );
and \U$9809 ( \10624 , \10621 , \10623 );
and \U$9810 ( \10625 , \9522 , \9289_nG290d );
and \U$9811 ( \10626 , \9345_nG282e , \9363 );
nor \U$9812 ( \10627 , \10624 , \10625 , \10626 );
and \U$9813 ( \10628 , \10572 , \9810 );
not \U$9814 ( \10629 , \9035_nG2a09 );
and \U$9815 ( \10630 , \9689 , \10629 );
and \U$9816 ( \10631 , \8924_nG2ae9 , \9814 );
nor \U$9817 ( \10632 , \10628 , \10630 , \10631 );
xor \U$9818 ( \10633 , \10627 , \10632 );
and \U$9819 ( \10634 , \10633 , \8481 );
and \U$9820 ( \10635 , \10627 , \10632 );
or \U$9821 ( \10636 , \10634 , \10635 );
nand \U$9822 ( \10637 , \9886_nG2554 , \8944 );
or \U$9823 ( \10638 , \8875 , \9679_nG25e2 );
nand \U$9824 ( \10639 , \10638 , \9046 );
and \U$9825 ( \10640 , \10637 , \10639 );
and \U$9826 ( \10641 , \9390 , \9679_nG25e2 );
and \U$9827 ( \10642 , \9886_nG2554 , \9392 );
nor \U$9828 ( \10643 , \10640 , \10641 , \10642 );
nand \U$9829 ( \10644 , \9637_nG26ac , \9119 );
or \U$9830 ( \10645 , \9057 , \9476_nG2758 );
nand \U$9831 ( \10646 , \10645 , \9223 );
and \U$9832 ( \10647 , \10644 , \10646 );
and \U$9833 ( \10648 , \9218 , \9476_nG2758 );
and \U$9834 ( \10649 , \9637_nG26ac , \9122 );
nor \U$9835 ( \10650 , \10647 , \10648 , \10649 );
xor \U$9836 ( \10651 , \10643 , \10650 );
nand \U$9837 ( \10652 , \9974_nG24b2 , \8775 );
or \U$9838 ( \10653 , \8672 , \10128_nG2440 );
nand \U$9839 ( \10654 , \10653 , \8781 );
and \U$9840 ( \10655 , \10652 , \10654 );
and \U$9841 ( \10656 , \8777 , \10128_nG2440 );
and \U$9842 ( \10657 , \9974_nG24b2 , \8866 );
nor \U$9843 ( \10658 , \10655 , \10656 , \10657 );
and \U$9844 ( \10659 , \10651 , \10658 );
and \U$9845 ( \10660 , \10643 , \10650 );
or \U$9846 ( \10661 , \10659 , \10660 );
xor \U$9847 ( \10662 , \10636 , \10661 );
and \U$9848 ( \10663 , \10407_nG236e , \8521 );
or \U$9849 ( \10664 , \8481 , \10504_nG2250 );
nand \U$9850 ( \10665 , \10664 , \8518 );
nand \U$9851 ( \10666 , \10407_nG236e , \8514 );
and \U$9852 ( \10667 , \10665 , \10666 );
and \U$9853 ( \10668 , \10504_nG2250 , \8663 );
nor \U$9854 ( \10669 , \10663 , \10667 , \10668 );
and \U$9855 ( \10670 , \10662 , \10669 );
and \U$9856 ( \10671 , \10636 , \10661 );
or \U$9857 ( \10672 , \10670 , \10671 );
not \U$9858 ( \10673 , \10594 );
not \U$9859 ( \10674 , \10600 );
and \U$9860 ( \10675 , \10673 , \10674 );
and \U$9861 ( \10676 , \10594 , \10600 );
nor \U$9862 ( \10677 , \10675 , \10676 );
xor \U$9863 ( \10678 , \10672 , \10677 );
xor \U$9864 ( \10679 , \10562 , \10586 );
xor \U$9865 ( \10680 , \10679 , \10589 );
and \U$9866 ( \10681 , \10678 , \10680 );
and \U$9867 ( \10682 , \10672 , \10677 );
or \U$9868 ( \10683 , \10681 , \10682 );
xor \U$9869 ( \10684 , \10456 , \10469 );
xor \U$9870 ( \10685 , \10684 , \10516 );
xor \U$9871 ( \10686 , \10683 , \10685 );
xor \U$9872 ( \10687 , \10592 , \10601 );
xor \U$9873 ( \10688 , \10687 , \10604 );
and \U$9874 ( \10689 , \10686 , \10688 );
and \U$9875 ( \10690 , \10683 , \10685 );
or \U$9876 ( \10691 , \10689 , \10690 );
xor \U$9877 ( \10692 , \10607 , \10612 );
xor \U$9878 ( \10693 , \10692 , \10615 );
and \U$9879 ( \10694 , \10691 , \10693 );
xor \U$9880 ( \10695 , \10636 , \10661 );
xor \U$9881 ( \10696 , \10695 , \10669 );
xor \U$9882 ( \10697 , \10569 , \10575 );
xor \U$9883 ( \10698 , \10697 , \10583 );
or \U$9884 ( \10699 , \10696 , \10698 );
and \U$9885 ( \10700 , \10407_nG236e , \8578 );
and \U$9886 ( \10701 , \8623 , \10238_nG23be );
nand \U$9887 ( \10702 , \10407_nG236e , \8575 );
or \U$9888 ( \10703 , \8535 , \10238_nG23be );
nand \U$9889 ( \10704 , \10703 , \8627 );
and \U$9890 ( \10705 , \10702 , \10704 );
nor \U$9891 ( \10706 , \10700 , \10701 , \10705 );
nand \U$9892 ( \10707 , \9476_nG2758 , \9360 );
or \U$9893 ( \10708 , \9234 , \9345_nG282e );
nand \U$9894 ( \10709 , \10708 , \9519 );
and \U$9895 ( \10710 , \10707 , \10709 );
and \U$9896 ( \10711 , \9522 , \9345_nG282e );
and \U$9897 ( \10712 , \9476_nG2758 , \9363 );
nor \U$9898 ( \10713 , \10710 , \10711 , \10712 );
and \U$9899 ( \10714 , \10629 , \9810 );
not \U$9900 ( \10715 , \9289_nG290d );
and \U$9901 ( \10716 , \9689 , \10715 );
and \U$9902 ( \10717 , \9035_nG2a09 , \9814 );
nor \U$9903 ( \10718 , \10714 , \10716 , \10717 );
xor \U$9904 ( \10719 , \10713 , \10718 );
nand \U$9905 ( \10720 , \9679_nG25e2 , \9119 );
or \U$9906 ( \10721 , \9057 , \9637_nG26ac );
nand \U$9907 ( \10722 , \10721 , \9223 );
and \U$9908 ( \10723 , \10720 , \10722 );
and \U$9909 ( \10724 , \9218 , \9637_nG26ac );
and \U$9910 ( \10725 , \9679_nG25e2 , \9122 );
nor \U$9911 ( \10726 , \10723 , \10724 , \10725 );
and \U$9912 ( \10727 , \10719 , \10726 );
and \U$9913 ( \10728 , \10713 , \10718 );
or \U$9914 ( \10729 , \10727 , \10728 );
xor \U$9915 ( \10730 , \10706 , \10729 );
nand \U$9916 ( \10731 , \10128_nG2440 , \8775 );
or \U$9917 ( \10732 , \8672 , \10238_nG23be );
nand \U$9918 ( \10733 , \10732 , \8781 );
and \U$9919 ( \10734 , \10731 , \10733 );
and \U$9920 ( \10735 , \8777 , \10238_nG23be );
and \U$9921 ( \10736 , \10128_nG2440 , \8866 );
nor \U$9922 ( \10737 , \10734 , \10735 , \10736 );
nand \U$9923 ( \10738 , \9974_nG24b2 , \8944 );
or \U$9924 ( \10739 , \8875 , \9886_nG2554 );
nand \U$9925 ( \10740 , \10739 , \9046 );
and \U$9926 ( \10741 , \10738 , \10740 );
and \U$9927 ( \10742 , \9390 , \9886_nG2554 );
and \U$9928 ( \10743 , \9974_nG24b2 , \9392 );
nor \U$9929 ( \10744 , \10741 , \10742 , \10743 );
xor \U$9930 ( \10745 , \10737 , \10744 );
and \U$9931 ( \10746 , \10504_nG2250 , \8578 );
and \U$9932 ( \10747 , \8623 , \10407_nG236e );
nand \U$9933 ( \10748 , \10504_nG2250 , \8575 );
or \U$9934 ( \10749 , \8535 , \10407_nG236e );
nand \U$9935 ( \10750 , \10749 , \8627 );
and \U$9936 ( \10751 , \10748 , \10750 );
nor \U$9937 ( \10752 , \10746 , \10747 , \10751 );
and \U$9938 ( \10753 , \10745 , \10752 );
and \U$9939 ( \10754 , \10737 , \10744 );
or \U$9940 ( \10755 , \10753 , \10754 );
and \U$9941 ( \10756 , \10730 , \10755 );
and \U$9942 ( \10757 , \10706 , \10729 );
or \U$9943 ( \10758 , \10756 , \10757 );
xor \U$9944 ( \10759 , \10544 , \10551 );
xor \U$9945 ( \10760 , \10759 , \10559 );
xor \U$9946 ( \10761 , \10758 , \10760 );
xor \U$9947 ( \10762 , \10643 , \10650 );
xor \U$9948 ( \10763 , \10762 , \10658 );
xor \U$9949 ( \10764 , \10627 , \10632 );
xor \U$9950 ( \10765 , \10764 , \8481 );
and \U$9951 ( \10766 , \10763 , \10765 );
nand \U$9952 ( \10767 , \10504_nG2250 , \8514 );
and \U$9953 ( \10768 , \8480 , \10767 );
and \U$9954 ( \10769 , \10504_nG2250 , \8521 );
nor \U$9955 ( \10770 , \10768 , \10769 );
xor \U$9956 ( \10771 , \10627 , \10632 );
xor \U$9957 ( \10772 , \10771 , \8481 );
and \U$9958 ( \10773 , \10770 , \10772 );
and \U$9959 ( \10774 , \10763 , \10770 );
or \U$9960 ( \10775 , \10766 , \10773 , \10774 );
and \U$9961 ( \10776 , \10761 , \10775 );
and \U$9962 ( \10777 , \10758 , \10760 );
or \U$9963 ( \10778 , \10776 , \10777 );
xor \U$9964 ( \10779 , \10699 , \10778 );
xor \U$9965 ( \10780 , \10672 , \10677 );
xor \U$9966 ( \10781 , \10780 , \10680 );
and \U$9967 ( \10782 , \10779 , \10781 );
and \U$9968 ( \10783 , \10699 , \10778 );
or \U$9969 ( \10784 , \10782 , \10783 );
xor \U$9970 ( \10785 , \10683 , \10685 );
xor \U$9971 ( \10786 , \10785 , \10688 );
and \U$9972 ( \10787 , \10784 , \10786 );
nand \U$9973 ( \10788 , \10128_nG2440 , \8944 );
or \U$9974 ( \10789 , \8875 , \9974_nG24b2 );
nand \U$9975 ( \10790 , \10789 , \9046 );
and \U$9976 ( \10791 , \10788 , \10790 );
and \U$9977 ( \10792 , \9390 , \9974_nG24b2 );
and \U$9978 ( \10793 , \10128_nG2440 , \9392 );
nor \U$9979 ( \10794 , \10791 , \10792 , \10793 );
nand \U$9980 ( \10795 , \9886_nG2554 , \9119 );
or \U$9981 ( \10796 , \9057 , \9679_nG25e2 );
nand \U$9982 ( \10797 , \10796 , \9223 );
and \U$9983 ( \10798 , \10795 , \10797 );
and \U$9984 ( \10799 , \9218 , \9679_nG25e2 );
and \U$9985 ( \10800 , \9886_nG2554 , \9122 );
nor \U$9986 ( \10801 , \10798 , \10799 , \10800 );
xor \U$9987 ( \10802 , \10794 , \10801 );
nand \U$9988 ( \10803 , \10238_nG23be , \8775 );
or \U$9989 ( \10804 , \8672 , \10407_nG236e );
nand \U$9990 ( \10805 , \10804 , \8781 );
and \U$9991 ( \10806 , \10803 , \10805 );
and \U$9992 ( \10807 , \8777 , \10407_nG236e );
and \U$9993 ( \10808 , \10238_nG23be , \8866 );
nor \U$9994 ( \10809 , \10806 , \10807 , \10808 );
and \U$9995 ( \10810 , \10802 , \10809 );
and \U$9996 ( \10811 , \10794 , \10801 );
or \U$9997 ( \10812 , \10810 , \10811 );
nand \U$9998 ( \10813 , \9637_nG26ac , \9360 );
or \U$9999 ( \10814 , \9234 , \9476_nG2758 );
nand \U$10000 ( \10815 , \10814 , \9519 );
and \U$10001 ( \10816 , \10813 , \10815 );
and \U$10002 ( \10817 , \9522 , \9476_nG2758 );
and \U$10003 ( \10818 , \9637_nG26ac , \9363 );
nor \U$10004 ( \10819 , \10816 , \10817 , \10818 );
and \U$10005 ( \10820 , \10715 , \9810 );
not \U$10006 ( \10821 , \9345_nG282e );
and \U$10007 ( \10822 , \9689 , \10821 );
and \U$10008 ( \10823 , \9289_nG290d , \9814 );
nor \U$10009 ( \10824 , \10820 , \10822 , \10823 );
xor \U$10010 ( \10825 , \10819 , \10824 );
and \U$10011 ( \10826 , \10825 , \8535 );
and \U$10012 ( \10827 , \10819 , \10824 );
or \U$10013 ( \10828 , \10826 , \10827 );
xor \U$10014 ( \10829 , \10812 , \10828 );
xor \U$10015 ( \10830 , \10737 , \10744 );
xor \U$10016 ( \10831 , \10830 , \10752 );
and \U$10017 ( \10832 , \10829 , \10831 );
and \U$10018 ( \10833 , \10812 , \10828 );
or \U$10019 ( \10834 , \10832 , \10833 );
xor \U$10020 ( \10835 , \10706 , \10729 );
xor \U$10021 ( \10836 , \10835 , \10755 );
xor \U$10022 ( \10837 , \10834 , \10836 );
xor \U$10023 ( \10838 , \10627 , \10632 );
xor \U$10024 ( \10839 , \10838 , \8481 );
xor \U$10025 ( \10840 , \10763 , \10770 );
xor \U$10026 ( \10841 , \10839 , \10840 );
and \U$10027 ( \10842 , \10837 , \10841 );
and \U$10028 ( \10843 , \10834 , \10836 );
or \U$10029 ( \10844 , \10842 , \10843 );
xor \U$10030 ( \10845 , \10758 , \10760 );
xor \U$10031 ( \10846 , \10845 , \10775 );
xor \U$10032 ( \10847 , \10844 , \10846 );
xnor \U$10033 ( \10848 , \10698 , \10696 );
xor \U$10034 ( \10849 , \10847 , \10848 );
not \U$10035 ( \10850 , \10849 );
xor \U$10036 ( \10851 , \10834 , \10836 );
xor \U$10037 ( \10852 , \10851 , \10841 );
or \U$10038 ( \10853 , \9123 , \9975 );
or \U$10039 ( \10854 , \9980 , \9219 );
or \U$10040 ( \10855 , \9120 , \9975 );
or \U$10041 ( \10856 , \9057 , \9886_nG2554 );
nand \U$10042 ( \10857 , \10856 , \9223 );
nand \U$10043 ( \10858 , \10855 , \10857 );
nand \U$10044 ( \10859 , \10853 , \10854 , \10858 );
and \U$10045 ( \10860 , \10821 , \9810 );
not \U$10046 ( \10861 , \9476_nG2758 );
and \U$10047 ( \10862 , \9689 , \10861 );
and \U$10048 ( \10863 , \9345_nG282e , \9814 );
nor \U$10049 ( \10864 , \10860 , \10862 , \10863 );
nand \U$10050 ( \10865 , \9679_nG25e2 , \9360 );
or \U$10051 ( \10866 , \9234 , \9637_nG26ac );
nand \U$10052 ( \10867 , \10866 , \9519 );
and \U$10053 ( \10868 , \10865 , \10867 );
and \U$10054 ( \10869 , \9522 , \9637_nG26ac );
and \U$10055 ( \10870 , \9679_nG25e2 , \9363 );
nor \U$10056 ( \10871 , \10868 , \10869 , \10870 );
nand \U$10057 ( \10872 , \10864 , \10871 );
and \U$10058 ( \10873 , \10859 , \10872 );
nor \U$10059 ( \10874 , \10871 , \10864 );
nor \U$10060 ( \10875 , \10873 , \10874 );
xor \U$10061 ( \10876 , \10794 , \10801 );
xor \U$10062 ( \10877 , \10876 , \10809 );
and \U$10063 ( \10878 , \10875 , \10877 );
and \U$10064 ( \10879 , \10504_nG2250 , \8623 );
not \U$10065 ( \10880 , \10504_nG2250 );
and \U$10066 ( \10881 , \10880 , \8577 );
not \U$10067 ( \10882 , \8627 );
nor \U$10068 ( \10883 , \10879 , \10881 , \10882 );
xor \U$10069 ( \10884 , \10794 , \10801 );
xor \U$10070 ( \10885 , \10884 , \10809 );
and \U$10071 ( \10886 , \10883 , \10885 );
and \U$10072 ( \10887 , \10875 , \10883 );
or \U$10073 ( \10888 , \10878 , \10886 , \10887 );
xor \U$10074 ( \10889 , \10713 , \10718 );
xor \U$10075 ( \10890 , \10889 , \10726 );
xor \U$10076 ( \10891 , \10888 , \10890 );
xor \U$10077 ( \10892 , \10812 , \10828 );
xor \U$10078 ( \10893 , \10892 , \10831 );
and \U$10079 ( \10894 , \10891 , \10893 );
and \U$10080 ( \10895 , \10888 , \10890 );
or \U$10081 ( \10896 , \10894 , \10895 );
nor \U$10082 ( \10897 , \10852 , \10896 );
xor \U$10083 ( \10898 , \10850 , \10897 );
and \U$10084 ( \10899 , \10852 , \10896 );
nor \U$10085 ( \10900 , \10899 , \10897 );
xor \U$10086 ( \10901 , \10888 , \10890 );
xor \U$10087 ( \10902 , \10901 , \10893 );
xor \U$10088 ( \10903 , \10819 , \10824 );
xor \U$10089 ( \10904 , \10903 , \8535 );
nand \U$10090 ( \10905 , \9886_nG2554 , \9360 );
or \U$10091 ( \10906 , \9234 , \9679_nG25e2 );
nand \U$10092 ( \10907 , \10906 , \9519 );
and \U$10093 ( \10908 , \10905 , \10907 );
and \U$10094 ( \10909 , \9522 , \9679_nG25e2 );
and \U$10095 ( \10910 , \9886_nG2554 , \9363 );
nor \U$10096 ( \10911 , \10908 , \10909 , \10910 );
and \U$10097 ( \10912 , \10861 , \9810 );
and \U$10098 ( \10913 , \9689 , \9939 );
and \U$10099 ( \10914 , \9476_nG2758 , \9814 );
nor \U$10100 ( \10915 , \10912 , \10913 , \10914 );
xor \U$10101 ( \10916 , \10911 , \10915 );
and \U$10102 ( \10917 , \10916 , \8672 );
and \U$10103 ( \10918 , \10911 , \10915 );
or \U$10104 ( \10919 , \10917 , \10918 );
nand \U$10105 ( \10920 , \10238_nG23be , \8944 );
or \U$10106 ( \10921 , \8875 , \10128_nG2440 );
nand \U$10107 ( \10922 , \10921 , \9046 );
and \U$10108 ( \10923 , \10920 , \10922 );
and \U$10109 ( \10924 , \9390 , \10128_nG2440 );
and \U$10110 ( \10925 , \10238_nG23be , \9392 );
nor \U$10111 ( \10926 , \10923 , \10924 , \10925 );
xor \U$10112 ( \10927 , \10919 , \10926 );
nand \U$10113 ( \10928 , \10407_nG236e , \8944 );
or \U$10114 ( \10929 , \8875 , \10238_nG23be );
nand \U$10115 ( \10930 , \10929 , \9046 );
and \U$10116 ( \10931 , \10928 , \10930 );
and \U$10117 ( \10932 , \9390 , \10238_nG23be );
and \U$10118 ( \10933 , \10407_nG236e , \9392 );
nor \U$10119 ( \10934 , \10931 , \10932 , \10933 );
nand \U$10120 ( \10935 , \10128_nG2440 , \9119 );
or \U$10121 ( \10936 , \9057 , \9974_nG24b2 );
nand \U$10122 ( \10937 , \10936 , \9223 );
and \U$10123 ( \10938 , \10935 , \10937 );
and \U$10124 ( \10939 , \9218 , \9974_nG24b2 );
and \U$10125 ( \10940 , \10128_nG2440 , \9122 );
nor \U$10126 ( \10941 , \10938 , \10939 , \10940 );
xor \U$10127 ( \10942 , \10934 , \10941 );
and \U$10128 ( \10943 , \8866 , \10504_nG2250 );
nand \U$10129 ( \10944 , \10504_nG2250 , \8775 );
and \U$10130 ( \10945 , \10944 , \8779 );
nor \U$10131 ( \10946 , \10943 , \10945 );
and \U$10132 ( \10947 , \10942 , \10946 );
and \U$10133 ( \10948 , \10934 , \10941 );
or \U$10134 ( \10949 , \10947 , \10948 );
and \U$10135 ( \10950 , \10927 , \10949 );
and \U$10136 ( \10951 , \10919 , \10926 );
or \U$10137 ( \10952 , \10950 , \10951 );
nand \U$10138 ( \10953 , \10904 , \10952 );
not \U$10139 ( \10954 , \10874 );
nand \U$10140 ( \10955 , \10954 , \10872 );
not \U$10141 ( \10956 , \10955 );
not \U$10142 ( \10957 , \10859 );
or \U$10143 ( \10958 , \10956 , \10957 );
or \U$10144 ( \10959 , \10859 , \10955 );
nand \U$10145 ( \10960 , \10958 , \10959 );
not \U$10146 ( \10961 , \10407_nG236e );
or \U$10147 ( \10962 , \8951 , \10961 );
or \U$10148 ( \10963 , \10880 , \8953 );
or \U$10149 ( \10964 , \8865 , \10961 );
or \U$10150 ( \10965 , \8672 , \10504_nG2250 );
nand \U$10151 ( \10966 , \10965 , \8781 );
nand \U$10152 ( \10967 , \10964 , \10966 );
nand \U$10153 ( \10968 , \10962 , \10963 , \10967 );
and \U$10154 ( \10969 , \10960 , \10968 );
and \U$10155 ( \10970 , \10953 , \10969 );
nor \U$10156 ( \10971 , \10952 , \10904 );
nor \U$10157 ( \10972 , \10970 , \10971 );
nor \U$10158 ( \10973 , \10902 , \10972 );
xor \U$10159 ( \10974 , \10900 , \10973 );
not \U$10160 ( \10975 , \10969 );
not \U$10161 ( \10976 , \10971 );
nand \U$10162 ( \10977 , \10976 , \10953 );
not \U$10163 ( \10978 , \10977 );
or \U$10164 ( \10979 , \10975 , \10978 );
or \U$10165 ( \10980 , \10977 , \10969 );
nand \U$10166 ( \10981 , \10979 , \10980 );
xor \U$10167 ( \10982 , \10794 , \10801 );
xor \U$10168 ( \10983 , \10982 , \10809 );
xor \U$10169 ( \10984 , \10875 , \10883 );
xor \U$10170 ( \10985 , \10983 , \10984 );
not \U$10171 ( \10986 , \10985 );
xor \U$10172 ( \10987 , \10981 , \10986 );
xor \U$10173 ( \10988 , \10919 , \10926 );
xor \U$10174 ( \10989 , \10988 , \10949 );
nand \U$10175 ( \10990 , \9974_nG24b2 , \9360 );
or \U$10176 ( \10991 , \9234 , \9886_nG2554 );
nand \U$10177 ( \10992 , \10991 , \9519 );
and \U$10178 ( \10993 , \10990 , \10992 );
and \U$10179 ( \10994 , \9522 , \9886_nG2554 );
and \U$10180 ( \10995 , \9974_nG24b2 , \9363 );
nor \U$10181 ( \10996 , \10993 , \10994 , \10995 );
and \U$10182 ( \10997 , \9939 , \9810 );
and \U$10183 ( \10998 , \9689 , \9978 );
and \U$10184 ( \10999 , \9637_nG26ac , \9814 );
nor \U$10185 ( \11000 , \10997 , \10998 , \10999 );
xor \U$10186 ( \11001 , \10996 , \11000 );
nand \U$10187 ( \11002 , \10238_nG23be , \9119 );
or \U$10188 ( \11003 , \9057 , \10128_nG2440 );
nand \U$10189 ( \11004 , \11003 , \9223 );
and \U$10190 ( \11005 , \11002 , \11004 );
and \U$10191 ( \11006 , \9218 , \10128_nG2440 );
and \U$10192 ( \11007 , \10238_nG23be , \9122 );
nor \U$10193 ( \11008 , \11005 , \11006 , \11007 );
and \U$10194 ( \11009 , \11001 , \11008 );
and \U$10195 ( \11010 , \10996 , \11000 );
or \U$10196 ( \11011 , \11009 , \11010 );
xor \U$10197 ( \11012 , \10911 , \10915 );
xor \U$10198 ( \11013 , \11012 , \8672 );
and \U$10199 ( \11014 , \11011 , \11013 );
xor \U$10200 ( \11015 , \10934 , \10941 );
xor \U$10201 ( \11016 , \11015 , \10946 );
xor \U$10202 ( \11017 , \10911 , \10915 );
xor \U$10203 ( \11018 , \11017 , \8672 );
and \U$10204 ( \11019 , \11016 , \11018 );
and \U$10205 ( \11020 , \11011 , \11016 );
or \U$10206 ( \11021 , \11014 , \11019 , \11020 );
nor \U$10207 ( \11022 , \10989 , \11021 );
xor \U$10208 ( \11023 , \10960 , \10968 );
or \U$10209 ( \11024 , \11022 , \11023 );
nand \U$10210 ( \11025 , \11021 , \10989 );
nand \U$10211 ( \11026 , \11024 , \11025 );
not \U$10212 ( \11027 , \11026 );
xor \U$10213 ( \11028 , \10987 , \11027 );
not \U$10214 ( \11029 , \11025 );
nor \U$10215 ( \11030 , \11029 , \11022 );
not \U$10216 ( \11031 , \11030 );
not \U$10217 ( \11032 , \11023 );
and \U$10218 ( \11033 , \11031 , \11032 );
and \U$10219 ( \11034 , \11030 , \11023 );
nor \U$10220 ( \11035 , \11033 , \11034 );
xor \U$10221 ( \11036 , \10911 , \10915 );
xor \U$10222 ( \11037 , \11036 , \8672 );
xor \U$10223 ( \11038 , \11011 , \11016 );
xor \U$10224 ( \11039 , \11037 , \11038 );
nand \U$10225 ( \11040 , \10504_nG2250 , \8944 );
or \U$10226 ( \11041 , \8875 , \10407_nG236e );
nand \U$10227 ( \11042 , \11041 , \9046 );
and \U$10228 ( \11043 , \11040 , \11042 );
and \U$10229 ( \11044 , \9390 , \10407_nG236e );
and \U$10230 ( \11045 , \10504_nG2250 , \9392 );
nor \U$10231 ( \11046 , \11043 , \11044 , \11045 );
nand \U$10232 ( \11047 , \10128_nG2440 , \9360 );
or \U$10233 ( \11048 , \9234 , \9974_nG24b2 );
nand \U$10234 ( \11049 , \11048 , \9519 );
and \U$10235 ( \11050 , \11047 , \11049 );
and \U$10236 ( \11051 , \9522 , \9974_nG24b2 );
and \U$10237 ( \11052 , \10128_nG2440 , \9363 );
nor \U$10238 ( \11053 , \11050 , \11051 , \11052 );
and \U$10239 ( \11054 , \9978 , \9810 );
and \U$10240 ( \11055 , \9689 , \9980 );
and \U$10241 ( \11056 , \9679_nG25e2 , \9814 );
nor \U$10242 ( \11057 , \11054 , \11055 , \11056 );
xor \U$10243 ( \11058 , \11053 , \11057 );
and \U$10244 ( \11059 , \11058 , \8875 );
and \U$10245 ( \11060 , \11053 , \11057 );
or \U$10246 ( \11061 , \11059 , \11060 );
xor \U$10247 ( \11062 , \11046 , \11061 );
nand \U$10248 ( \11063 , \10407_nG236e , \9119 );
or \U$10249 ( \11064 , \9057 , \10238_nG23be );
nand \U$10250 ( \11065 , \11064 , \9223 );
and \U$10251 ( \11066 , \11063 , \11065 );
and \U$10252 ( \11067 , \9218 , \10238_nG23be );
and \U$10253 ( \11068 , \10407_nG236e , \9122 );
nor \U$10254 ( \11069 , \11066 , \11067 , \11068 );
not \U$10255 ( \11070 , \11069 );
or \U$10256 ( \11071 , \9042 , \10880 );
or \U$10257 ( \11072 , \10504_nG2250 , \8875 );
nand \U$10258 ( \11073 , \11071 , \11072 , \9046 );
nand \U$10259 ( \11074 , \11070 , \11073 );
and \U$10260 ( \11075 , \11062 , \11074 );
and \U$10261 ( \11076 , \11046 , \11061 );
or \U$10262 ( \11077 , \11075 , \11076 );
nor \U$10263 ( \11078 , \11039 , \11077 );
xor \U$10264 ( \11079 , \11035 , \11078 );
xor \U$10265 ( \11080 , \11046 , \11061 );
xor \U$10266 ( \11081 , \11080 , \11074 );
xor \U$10267 ( \11082 , \10996 , \11000 );
xor \U$10268 ( \11083 , \11082 , \11008 );
and \U$10269 ( \11084 , \11081 , \11083 );
nor \U$10270 ( \11085 , \11081 , \11083 );
nor \U$10271 ( \11086 , \11084 , \11085 );
not \U$10272 ( \11087 , \11069 );
not \U$10273 ( \11088 , \11073 );
or \U$10274 ( \11089 , \11087 , \11088 );
or \U$10275 ( \11090 , \11073 , \11069 );
nand \U$10276 ( \11091 , \11089 , \11090 );
xor \U$10277 ( \11092 , \11053 , \11057 );
xor \U$10278 ( \11093 , \11092 , \8875 );
nand \U$10279 ( \11094 , \10238_nG23be , \9360 );
or \U$10280 ( \11095 , \9234 , \10128_nG2440 );
nand \U$10281 ( \11096 , \11095 , \9519 );
and \U$10282 ( \11097 , \11094 , \11096 );
and \U$10283 ( \11098 , \9522 , \10128_nG2440 );
and \U$10284 ( \11099 , \10238_nG23be , \9363 );
nor \U$10285 ( \11100 , \11097 , \11098 , \11099 );
and \U$10286 ( \11101 , \9980 , \9810 );
and \U$10287 ( \11102 , \9689 , \9975 );
and \U$10288 ( \11103 , \9886_nG2554 , \9814 );
nor \U$10289 ( \11104 , \11101 , \11102 , \11103 );
xor \U$10290 ( \11105 , \11100 , \11104 );
nand \U$10291 ( \11106 , \10504_nG2250 , \9119 );
or \U$10292 ( \11107 , \9057 , \10407_nG236e );
nand \U$10293 ( \11108 , \11107 , \9223 );
and \U$10294 ( \11109 , \11106 , \11108 );
and \U$10295 ( \11110 , \9218 , \10407_nG236e );
and \U$10296 ( \11111 , \10504_nG2250 , \9122 );
nor \U$10297 ( \11112 , \11109 , \11110 , \11111 );
and \U$10298 ( \11113 , \11105 , \11112 );
and \U$10299 ( \11114 , \11100 , \11104 );
or \U$10300 ( \11115 , \11113 , \11114 );
nand \U$10301 ( \11116 , \11093 , \11115 );
and \U$10302 ( \11117 , \11091 , \11116 );
nor \U$10303 ( \11118 , \11115 , \11093 );
nor \U$10304 ( \11119 , \11117 , \11118 );
not \U$10305 ( \11120 , \11119 );
xor \U$10306 ( \11121 , \11086 , \11120 );
not \U$10307 ( \11122 , \11091 );
not \U$10308 ( \11123 , \11116 );
nor \U$10309 ( \11124 , \11123 , \11118 );
not \U$10310 ( \11125 , \11124 );
and \U$10311 ( \11126 , \11122 , \11125 );
and \U$10312 ( \11127 , \11091 , \11124 );
nor \U$10313 ( \11128 , \11126 , \11127 );
xor \U$10314 ( \11129 , \11100 , \11104 );
xor \U$10315 ( \11130 , \11129 , \11112 );
and \U$10316 ( \11131 , \9975 , \9810 );
not \U$10317 ( \11132 , \10128_nG2440 );
and \U$10318 ( \11133 , \9689 , \11132 );
and \U$10319 ( \11134 , \9974_nG24b2 , \9814 );
nor \U$10320 ( \11135 , \11131 , \11133 , \11134 );
xor \U$10321 ( \11136 , \9057 , \11135 );
nand \U$10322 ( \11137 , \10407_nG236e , \9360 );
or \U$10323 ( \11138 , \9234 , \10238_nG23be );
nand \U$10324 ( \11139 , \11138 , \9519 );
and \U$10325 ( \11140 , \11137 , \11139 );
and \U$10326 ( \11141 , \9522 , \10238_nG23be );
and \U$10327 ( \11142 , \10407_nG236e , \9363 );
nor \U$10328 ( \11143 , \11140 , \11141 , \11142 );
and \U$10329 ( \11144 , \11136 , \11143 );
and \U$10330 ( \11145 , \9057 , \11135 );
or \U$10331 ( \11146 , \11144 , \11145 );
nor \U$10332 ( \11147 , \11130 , \11146 );
xor \U$10333 ( \11148 , \11128 , \11147 );
not \U$10334 ( \11149 , \10238_nG23be );
or \U$10335 ( \11150 , \9813 , \11149 );
or \U$10336 ( \11151 , \10238_nG23be , \9691 );
or \U$10337 ( \11152 , \10407_nG236e , \9690 );
nand \U$10338 ( \11153 , \11150 , \11151 , \11152 );
xor \U$10339 ( \11154 , \11153 , \9362 );
and \U$10340 ( \11155 , \10961 , \9810 );
and \U$10341 ( \11156 , \9689 , \10880 );
and \U$10342 ( \11157 , \10407_nG236e , \9814 );
nor \U$10343 ( \11158 , \11155 , \11156 , \11157 );
nand \U$10344 ( \11159 , \10504_nG2250 , \9690 );
nand \U$10345 ( \11160 , \9229 , \11159 );
nor \U$10346 ( \11161 , \11158 , \11160 );
xor \U$10347 ( \11162 , \11154 , \11161 );
or \U$10348 ( \11163 , \9694 , \10880 );
or \U$10349 ( \11164 , \10504_nG2250 , \9234 );
nand \U$10350 ( \11165 , \11163 , \11164 , \9519 );
and \U$10351 ( \11166 , \11162 , \11165 );
and \U$10352 ( \11167 , \11154 , \11161 );
or \U$10353 ( \11168 , \11166 , \11167 );
and \U$10354 ( \11169 , \11153 , \9362 );
xor \U$10355 ( \11170 , \11168 , \11169 );
nand \U$10356 ( \11171 , \10504_nG2250 , \9360 );
or \U$10357 ( \11172 , \9234 , \10407_nG236e );
nand \U$10358 ( \11173 , \11172 , \9519 );
and \U$10359 ( \11174 , \11171 , \11173 );
and \U$10360 ( \11175 , \9522 , \10407_nG236e );
and \U$10361 ( \11176 , \10504_nG2250 , \9363 );
nor \U$10362 ( \11177 , \11174 , \11175 , \11176 );
and \U$10363 ( \11178 , \11132 , \9810 );
and \U$10364 ( \11179 , \9689 , \11149 );
and \U$10365 ( \11180 , \10128_nG2440 , \9814 );
nor \U$10366 ( \11181 , \11178 , \11179 , \11180 );
and \U$10367 ( \11182 , \11177 , \11181 );
nor \U$10368 ( \11183 , \11177 , \11181 );
nor \U$10369 ( \11184 , \11182 , \11183 );
and \U$10370 ( \11185 , \11170 , \11184 );
and \U$10371 ( \11186 , \11168 , \11169 );
or \U$10372 ( \11187 , \11185 , \11186 );
xor \U$10373 ( \11188 , \11187 , \11183 );
and \U$10374 ( \11189 , \10504_nG2250 , \9218 );
and \U$10375 ( \11190 , \10880 , \9121 );
not \U$10376 ( \11191 , \9223 );
nor \U$10377 ( \11192 , \11189 , \11190 , \11191 );
xor \U$10378 ( \11193 , \9057 , \11135 );
xor \U$10379 ( \11194 , \11193 , \11143 );
and \U$10380 ( \11195 , \11192 , \11194 );
nor \U$10381 ( \11196 , \11192 , \11194 );
nor \U$10382 ( \11197 , \11195 , \11196 );
and \U$10383 ( \11198 , \11188 , \11197 );
and \U$10384 ( \11199 , \11187 , \11183 );
or \U$10385 ( \11200 , \11198 , \11199 );
xor \U$10386 ( \11201 , \11200 , \11196 );
and \U$10387 ( \11202 , \11130 , \11146 );
nor \U$10388 ( \11203 , \11202 , \11147 );
and \U$10389 ( \11204 , \11201 , \11203 );
and \U$10390 ( \11205 , \11200 , \11196 );
or \U$10391 ( \11206 , \11204 , \11205 );
and \U$10392 ( \11207 , \11148 , \11206 );
and \U$10393 ( \11208 , \11128 , \11147 );
or \U$10394 ( \11209 , \11207 , \11208 );
and \U$10395 ( \11210 , \11121 , \11209 );
and \U$10396 ( \11211 , \11086 , \11120 );
or \U$10397 ( \11212 , \11210 , \11211 );
xor \U$10398 ( \11213 , \11212 , \11085 );
and \U$10399 ( \11214 , \11039 , \11077 );
nor \U$10400 ( \11215 , \11214 , \11078 );
and \U$10401 ( \11216 , \11213 , \11215 );
and \U$10402 ( \11217 , \11212 , \11085 );
or \U$10403 ( \11218 , \11216 , \11217 );
and \U$10404 ( \11219 , \11079 , \11218 );
and \U$10405 ( \11220 , \11035 , \11078 );
or \U$10406 ( \11221 , \11219 , \11220 );
and \U$10407 ( \11222 , \11028 , \11221 );
and \U$10408 ( \11223 , \10987 , \11027 );
or \U$10409 ( \11224 , \11222 , \11223 );
and \U$10410 ( \11225 , \10981 , \10986 );
xor \U$10411 ( \11226 , \11224 , \11225 );
and \U$10412 ( \11227 , \10902 , \10972 );
nor \U$10413 ( \11228 , \11227 , \10973 );
and \U$10414 ( \11229 , \11226 , \11228 );
and \U$10415 ( \11230 , \11224 , \11225 );
or \U$10416 ( \11231 , \11229 , \11230 );
and \U$10417 ( \11232 , \10974 , \11231 );
and \U$10418 ( \11233 , \10900 , \10973 );
or \U$10419 ( \11234 , \11232 , \11233 );
and \U$10420 ( \11235 , \10898 , \11234 );
and \U$10421 ( \11236 , \10850 , \10897 );
or \U$10422 ( \11237 , \11235 , \11236 );
xor \U$10423 ( \11238 , \10844 , \10846 );
and \U$10424 ( \11239 , \11238 , \10848 );
and \U$10425 ( \11240 , \10844 , \10846 );
or \U$10426 ( \11241 , \11239 , \11240 );
xor \U$10427 ( \11242 , \10699 , \10778 );
xor \U$10428 ( \11243 , \11242 , \10781 );
nand \U$10429 ( \11244 , \11241 , \11243 );
and \U$10430 ( \11245 , \11237 , \11244 );
nor \U$10431 ( \11246 , \11243 , \11241 );
nor \U$10432 ( \11247 , \11245 , \11246 );
xor \U$10433 ( \11248 , \10683 , \10685 );
xor \U$10434 ( \11249 , \11248 , \10688 );
and \U$10435 ( \11250 , \11247 , \11249 );
and \U$10436 ( \11251 , \10784 , \11247 );
or \U$10437 ( \11252 , \10787 , \11250 , \11251 );
xor \U$10438 ( \11253 , \10607 , \10612 );
xor \U$10439 ( \11254 , \11253 , \10615 );
and \U$10440 ( \11255 , \11252 , \11254 );
and \U$10441 ( \11256 , \10691 , \11252 );
or \U$10442 ( \11257 , \10694 , \11255 , \11256 );
not \U$10443 ( \11258 , \11257 );
and \U$10444 ( \11259 , \10620 , \11258 );
and \U$10445 ( \11260 , \10537 , \10619 );
or \U$10446 ( \11261 , \11259 , \11260 );
and \U$10447 ( \11262 , \10535 , \11261 );
and \U$10448 ( \11263 , \10529 , \10534 );
or \U$10449 ( \11264 , \11262 , \11263 );
and \U$10450 ( \11265 , \10527 , \11264 );
and \U$10451 ( \11266 , \10357 , \10526 );
or \U$10452 ( \11267 , \11265 , \11266 );
and \U$10453 ( \11268 , \10353 , \11267 );
and \U$10454 ( \11269 , \10266 , \10352 );
or \U$10455 ( \11270 , \11268 , \11269 );
and \U$10456 ( \11271 , \10264 , \11270 );
and \U$10457 ( \11272 , \10094 , \10263 );
or \U$10458 ( \11273 , \11271 , \11272 );
and \U$10459 ( \11274 , \10092 , \11273 );
and \U$10460 ( \11275 , \10089 , \10091 );
or \U$10461 ( \11276 , \11274 , \11275 );
and \U$10462 ( \11277 , \10015 , \11276 );
and \U$10463 ( \11278 , \10012 , \10014 );
or \U$10464 ( \11279 , \11277 , \11278 );
and \U$10465 ( \11280 , \9849 , \11279 );
and \U$10466 ( \11281 , \9737 , \9848 );
or \U$10467 ( \11282 , \11280 , \11281 );
and \U$10468 ( \11283 , \9724 , \9733 );
nor \U$10469 ( \11284 , \11283 , \9726 );
not \U$10470 ( \11285 , \9563 );
nor \U$10471 ( \11286 , \9555 , \9566 );
not \U$10472 ( \11287 , \11286 );
or \U$10473 ( \11288 , \11285 , \11287 );
or \U$10474 ( \11289 , \11286 , \9563 );
nand \U$10475 ( \11290 , \11288 , \11289 );
nand \U$10476 ( \11291 , \11284 , \11290 );
and \U$10477 ( \11292 , \11282 , \11291 );
nor \U$10478 ( \11293 , \11290 , \11284 );
nor \U$10479 ( \11294 , \11292 , \11293 );
not \U$10480 ( \11295 , \11294 );
and \U$10481 ( \11296 , \9568 , \11295 );
and \U$10482 ( \11297 , \9428 , \9567 );
or \U$10483 ( \11298 , \11296 , \11297 );
and \U$10484 ( \11299 , \9426 , \11298 );
and \U$10485 ( \11300 , \9421 , \9425 );
or \U$10486 ( \11301 , \11299 , \11300 );
and \U$10487 ( \11302 , \9313 , \11301 );
and \U$10488 ( \11303 , \9200 , \9312 );
or \U$10489 ( \11304 , \11302 , \11303 );
not \U$10490 ( \11305 , \9191 );
not \U$10491 ( \11306 , \9196 );
or \U$10492 ( \11307 , \11305 , \11306 );
nand \U$10493 ( \11308 , \11307 , \9192 );
xor \U$10494 ( \11309 , \9086 , \9088 );
xor \U$10495 ( \11310 , \11309 , \9091 );
nand \U$10496 ( \11311 , \11308 , \11310 );
and \U$10497 ( \11312 , \11304 , \11311 );
nor \U$10498 ( \11313 , \11310 , \11308 );
nor \U$10499 ( \11314 , \11312 , \11313 );
and \U$10500 ( \11315 , \9102 , \11314 );
and \U$10501 ( \11316 , \9094 , \9101 );
or \U$10502 ( \11317 , \11315 , \11316 );
not \U$10503 ( \11318 , \11317 );
and \U$10504 ( \11319 , \8986 , \11318 );
and \U$10505 ( \11320 , \8808 , \8985 );
or \U$10506 ( \11321 , \11319 , \11320 );
not \U$10507 ( \11322 , \8614 );
not \U$10508 ( \11323 , \8684 );
and \U$10509 ( \11324 , \11322 , \11323 );
and \U$10510 ( \11325 , \8684 , \8614 );
nor \U$10511 ( \11326 , \11324 , \11325 );
and \U$10512 ( \11327 , \8798 , \8804 );
nor \U$10513 ( \11328 , \11327 , \8800 );
nand \U$10514 ( \11329 , \11326 , \11328 );
and \U$10515 ( \11330 , \11321 , \11329 );
nor \U$10516 ( \11331 , \11328 , \11326 );
nor \U$10517 ( \11332 , \11330 , \11331 );
not \U$10518 ( \11333 , \11332 );
or \U$10519 ( \11334 , \8690 , \11333 );
or \U$10520 ( \11335 , \11332 , \8689 );
nand \U$10521 ( \11336 , \11334 , \11335 );
and \U$10522 ( \11337 , \7896 , \7899 );
not \U$10523 ( \11338 , \7897 );
nor \U$10524 ( \11339 , \11337 , \11338 );
xnor \U$10525 ( \11340 , RIb55bd18_600, \11339 );
and \U$10526 ( \11341 , \11340 , \7916 , RIb55bd90_601);
and \U$10527 ( \11342 , \11341 , RIb551890_249);
and \U$10528 ( \11343 , \7943 , RIb551d40_259);
and \U$10529 ( \11344 , RIb551cc8_258, \7955 );
nor \U$10530 ( \11345 , \11343 , \11344 );
and \U$10531 ( \11346 , \7914 , RIb551b60_255);
and \U$10532 ( \11347 , RIb551ae8_254, \7906 );
nor \U$10533 ( \11348 , \11346 , \11347 );
and \U$10534 ( \11349 , \7953 , RIb551a70_253);
and \U$10535 ( \11350 , RIb5519f8_252, \7900 );
nor \U$10536 ( \11351 , \11349 , \11350 );
and \U$10537 ( \11352 , \7926 , RIb551c50_257);
and \U$10538 ( \11353 , RIb551bd8_256, \7910 );
nor \U$10539 ( \11354 , \11352 , \11353 );
nand \U$10540 ( \11355 , \11345 , \11348 , \11351 , \11354 );
and \U$10541 ( \11356 , \7950 , RIb551980_251);
and \U$10542 ( \11357 , RIb551908_250, \7917 );
nor \U$10543 ( \11358 , \11356 , \11357 );
not \U$10544 ( \11359 , \11358 );
nor \U$10545 ( \11360 , \11342 , \11355 , \11359 );
and \U$10546 ( \11361 , \7948 , RIb551f20_263);
and \U$10547 ( \11362 , RIb551ea8_262, \7936 );
nor \U$10548 ( \11363 , \11361 , \11362 );
and \U$10549 ( \11364 , \7938 , RIb551e30_261);
and \U$10550 ( \11365 , RIb551db8_260, \7945 );
nor \U$10551 ( \11366 , \11364 , \11365 );
nand \U$10552 ( \11367 , \11360 , \11363 , \7931 , \11366 );
buf \U$10553 ( \11368 , \11367 );
buf \U$10554 ( \11369 , \7962 );
_DC g2aeb ( \11370_nG2aeb , \11368 , \11369 );
xor \U$10555 ( \11371 , \7889 , \11370_nG2aeb );
and \U$10556 ( \11372 , \11341 , RIb54ac48_18);
and \U$10557 ( \11373 , \7943 , RIb54b0f8_28);
and \U$10558 ( \11374 , RIb54b080_27, \7955 );
nor \U$10559 ( \11375 , \11373 , \11374 );
and \U$10560 ( \11376 , \7914 , RIb54af18_24);
and \U$10561 ( \11377 , RIb54aea0_23, \7906 );
nor \U$10562 ( \11378 , \11376 , \11377 );
and \U$10563 ( \11379 , \7953 , RIb54ae28_22);
and \U$10564 ( \11380 , RIb54adb0_21, \7900 );
nor \U$10565 ( \11381 , \11379 , \11380 );
and \U$10566 ( \11382 , \7926 , RIb54b008_26);
and \U$10567 ( \11383 , RIb54af90_25, \7910 );
nor \U$10568 ( \11384 , \11382 , \11383 );
nand \U$10569 ( \11385 , \11375 , \11378 , \11381 , \11384 );
and \U$10570 ( \11386 , \7950 , RIb54ad38_20);
and \U$10571 ( \11387 , RIb54acc0_19, \7917 );
nor \U$10572 ( \11388 , \11386 , \11387 );
not \U$10573 ( \11389 , \11388 );
nor \U$10574 ( \11390 , \11372 , \11385 , \11389 );
and \U$10575 ( \11391 , \7948 , RIb54b2d8_32);
and \U$10576 ( \11392 , RIb54b260_31, \7936 );
nor \U$10577 ( \11393 , \11391 , \11392 );
and \U$10578 ( \11394 , \7938 , RIb54b1e8_30);
and \U$10579 ( \11395 , RIb54b170_29, \7945 );
nor \U$10580 ( \11396 , \11394 , \11395 );
nand \U$10581 ( \11397 , \11390 , \11393 , \7986 , \11396 );
buf \U$10582 ( \11398 , \11397 );
_DC g2911 ( \11399_nG2911 , \11398 , \11369 );
xor \U$10583 ( \11400 , \7970 , \11399_nG2911 );
and \U$10584 ( \11401 , \11341 , RIb54b440_35);
and \U$10585 ( \11402 , \7943 , RIb54b8f0_45);
and \U$10586 ( \11403 , RIb54b878_44, \7955 );
nor \U$10587 ( \11404 , \11402 , \11403 );
and \U$10588 ( \11405 , \7914 , RIb54b710_41);
and \U$10589 ( \11406 , RIb54b698_40, \7906 );
nor \U$10590 ( \11407 , \11405 , \11406 );
and \U$10591 ( \11408 , \7953 , RIb54b620_39);
and \U$10592 ( \11409 , RIb54b5a8_38, \7900 );
nor \U$10593 ( \11410 , \11408 , \11409 );
and \U$10594 ( \11411 , \7926 , RIb54b800_43);
and \U$10595 ( \11412 , RIb54b788_42, \7910 );
nor \U$10596 ( \11413 , \11411 , \11412 );
nand \U$10597 ( \11414 , \11404 , \11407 , \11410 , \11413 );
and \U$10598 ( \11415 , \7950 , RIb54b530_37);
and \U$10599 ( \11416 , RIb54b4b8_36, \7917 );
nor \U$10600 ( \11417 , \11415 , \11416 );
not \U$10601 ( \11418 , \11417 );
nor \U$10602 ( \11419 , \11401 , \11414 , \11418 );
and \U$10603 ( \11420 , \7948 , RIb54bad0_49);
and \U$10604 ( \11421 , RIb54ba58_48, \7936 );
nor \U$10605 ( \11422 , \11420 , \11421 );
and \U$10606 ( \11423 , \7938 , RIb54b9e0_47);
and \U$10607 ( \11424 , RIb54b968_46, \7945 );
nor \U$10608 ( \11425 , \11423 , \11424 );
nand \U$10609 ( \11426 , \11419 , \11422 , \8018 , \11425 );
buf \U$10610 ( \11427 , \11426 );
_DC g290f ( \11428_nG290f , \11427 , \11369 );
xor \U$10611 ( \11429 , \8006 , \11428_nG290f );
and \U$10612 ( \11430 , \11341 , RIb54bc38_52);
and \U$10613 ( \11431 , \7943 , RIb54c0e8_62);
and \U$10614 ( \11432 , RIb54c070_61, \7955 );
nor \U$10615 ( \11433 , \11431 , \11432 );
and \U$10616 ( \11434 , \7914 , RIb54bf08_58);
and \U$10617 ( \11435 , RIb54be90_57, \7906 );
nor \U$10618 ( \11436 , \11434 , \11435 );
and \U$10619 ( \11437 , \7953 , RIb54be18_56);
and \U$10620 ( \11438 , RIb54bda0_55, \7900 );
nor \U$10621 ( \11439 , \11437 , \11438 );
and \U$10622 ( \11440 , \7926 , RIb54bff8_60);
and \U$10623 ( \11441 , RIb54bf80_59, \7910 );
nor \U$10624 ( \11442 , \11440 , \11441 );
nand \U$10625 ( \11443 , \11433 , \11436 , \11439 , \11442 );
and \U$10626 ( \11444 , \7950 , RIb54bd28_54);
and \U$10627 ( \11445 , RIb54bcb0_53, \7917 );
nor \U$10628 ( \11446 , \11444 , \11445 );
not \U$10629 ( \11447 , \11446 );
nor \U$10630 ( \11448 , \11430 , \11443 , \11447 );
and \U$10631 ( \11449 , \7948 , RIb54c2c8_66);
and \U$10632 ( \11450 , RIb54c250_65, \7936 );
nor \U$10633 ( \11451 , \11449 , \11450 );
and \U$10634 ( \11452 , \7938 , RIb54c1d8_64);
and \U$10635 ( \11453 , RIb54c160_63, \7945 );
nor \U$10636 ( \11454 , \11452 , \11453 );
nand \U$10637 ( \11455 , \11448 , \11451 , \8056 , \11454 );
buf \U$10638 ( \11456 , \11455 );
_DC g275c ( \11457_nG275c , \11456 , \11369 );
xor \U$10639 ( \11458 , \8044 , \11457_nG275c );
and \U$10640 ( \11459 , \11341 , RIb54c430_69);
and \U$10641 ( \11460 , \7943 , RIb54c8e0_79);
and \U$10642 ( \11461 , RIb54c868_78, \7955 );
nor \U$10643 ( \11462 , \11460 , \11461 );
and \U$10644 ( \11463 , \7914 , RIb54c700_75);
and \U$10645 ( \11464 , RIb54c688_74, \7906 );
nor \U$10646 ( \11465 , \11463 , \11464 );
and \U$10647 ( \11466 , \7953 , RIb54c610_73);
and \U$10648 ( \11467 , RIb54c598_72, \7900 );
nor \U$10649 ( \11468 , \11466 , \11467 );
and \U$10650 ( \11469 , \7926 , RIb54c7f0_77);
and \U$10651 ( \11470 , RIb54c778_76, \7910 );
nor \U$10652 ( \11471 , \11469 , \11470 );
nand \U$10653 ( \11472 , \11462 , \11465 , \11468 , \11471 );
and \U$10654 ( \11473 , \7950 , RIb54c520_71);
and \U$10655 ( \11474 , RIb54c4a8_70, \7917 );
nor \U$10656 ( \11475 , \11473 , \11474 );
not \U$10657 ( \11476 , \11475 );
nor \U$10658 ( \11477 , \11459 , \11472 , \11476 );
and \U$10659 ( \11478 , \7948 , RIb54cac0_83);
and \U$10660 ( \11479 , RIb54ca48_82, \7936 );
nor \U$10661 ( \11480 , \11478 , \11479 );
and \U$10662 ( \11481 , \7938 , RIb54c9d0_81);
and \U$10663 ( \11482 , RIb54c958_80, \7945 );
nor \U$10664 ( \11483 , \11481 , \11482 );
nand \U$10665 ( \11484 , \11477 , \11480 , \8098 , \11483 );
buf \U$10666 ( \11485 , \11484 );
_DC g275a ( \11486_nG275a , \11485 , \11369 );
xor \U$10667 ( \11487 , \8082 , \11486_nG275a );
and \U$10668 ( \11488 , \11341 , RIb54cc28_86);
and \U$10669 ( \11489 , \7943 , RIb54d0d8_96);
and \U$10670 ( \11490 , RIb54d060_95, \7955 );
nor \U$10671 ( \11491 , \11489 , \11490 );
and \U$10672 ( \11492 , \7914 , RIb54cef8_92);
and \U$10673 ( \11493 , RIb54ce80_91, \7906 );
nor \U$10674 ( \11494 , \11492 , \11493 );
and \U$10675 ( \11495 , \7953 , RIb54ce08_90);
and \U$10676 ( \11496 , RIb54cd90_89, \7900 );
nor \U$10677 ( \11497 , \11495 , \11496 );
and \U$10678 ( \11498 , \7926 , RIb54cfe8_94);
and \U$10679 ( \11499 , RIb54cf70_93, \7910 );
nor \U$10680 ( \11500 , \11498 , \11499 );
nand \U$10681 ( \11501 , \11491 , \11494 , \11497 , \11500 );
and \U$10682 ( \11502 , \7950 , RIb54cd18_88);
and \U$10683 ( \11503 , RIb54cca0_87, \7917 );
nor \U$10684 ( \11504 , \11502 , \11503 );
not \U$10685 ( \11505 , \11504 );
nor \U$10686 ( \11506 , \11488 , \11501 , \11505 );
and \U$10687 ( \11507 , \7948 , RIb54d2b8_100);
and \U$10688 ( \11508 , RIb54d240_99, \7936 );
nor \U$10689 ( \11509 , \11507 , \11508 );
and \U$10690 ( \11510 , \7938 , RIb54d1c8_98);
and \U$10691 ( \11511 , RIb54d150_97, \7945 );
nor \U$10692 ( \11512 , \11510 , \11511 );
nand \U$10693 ( \11513 , \11506 , \11509 , \8130 , \11512 );
buf \U$10694 ( \11514 , \11513 );
_DC g25e6 ( \11515_nG25e6 , \11514 , \11369 );
xor \U$10695 ( \11516 , \8118 , \11515_nG25e6 );
and \U$10696 ( \11517 , \11341 , RIb54d420_103);
and \U$10697 ( \11518 , \7943 , RIb54d8d0_113);
and \U$10698 ( \11519 , RIb54d858_112, \7955 );
nor \U$10699 ( \11520 , \11518 , \11519 );
and \U$10700 ( \11521 , \7914 , RIb54d6f0_109);
and \U$10701 ( \11522 , RIb54d678_108, \7906 );
nor \U$10702 ( \11523 , \11521 , \11522 );
and \U$10703 ( \11524 , \7953 , RIb54d600_107);
and \U$10704 ( \11525 , RIb54d588_106, \7900 );
nor \U$10705 ( \11526 , \11524 , \11525 );
and \U$10706 ( \11527 , \7926 , RIb54d7e0_111);
and \U$10707 ( \11528 , RIb54d768_110, \7910 );
nor \U$10708 ( \11529 , \11527 , \11528 );
nand \U$10709 ( \11530 , \11520 , \11523 , \11526 , \11529 );
and \U$10710 ( \11531 , \7950 , RIb54d510_105);
and \U$10711 ( \11532 , RIb54d498_104, \7917 );
nor \U$10712 ( \11533 , \11531 , \11532 );
not \U$10713 ( \11534 , \11533 );
nor \U$10714 ( \11535 , \11517 , \11530 , \11534 );
and \U$10715 ( \11536 , \7948 , RIb54dab0_117);
and \U$10716 ( \11537 , RIb54da38_116, \7936 );
nor \U$10717 ( \11538 , \11536 , \11537 );
and \U$10718 ( \11539 , \7938 , RIb54d9c0_115);
and \U$10719 ( \11540 , RIb54d948_114, \7945 );
nor \U$10720 ( \11541 , \11539 , \11540 );
nand \U$10721 ( \11542 , \11535 , \11538 , \8168 , \11541 );
buf \U$10722 ( \11543 , \11542 );
_DC g25e4 ( \11544_nG25e4 , \11543 , \11369 );
xor \U$10723 ( \11545 , \8156 , \11544_nG25e4 );
and \U$10724 ( \11546 , \11341 , RIb54dc18_120);
and \U$10725 ( \11547 , \7914 , RIb54dee8_126);
and \U$10726 ( \11548 , RIb54de70_125, \7906 );
nor \U$10727 ( \11549 , \11547 , \11548 );
and \U$10728 ( \11550 , \7936 , RIb54e230_133);
and \U$10729 ( \11551 , RIb54e1b8_132, \7938 );
nor \U$10730 ( \11552 , \11550 , \11551 );
and \U$10731 ( \11553 , \7953 , RIb54ddf8_124);
and \U$10732 ( \11554 , RIb54dd80_123, \7900 );
nor \U$10733 ( \11555 , \11553 , \11554 );
and \U$10734 ( \11556 , \7943 , RIb54e0c8_130);
and \U$10735 ( \11557 , RIb54e140_131, \7945 );
nor \U$10736 ( \11558 , \11556 , \11557 );
nand \U$10737 ( \11559 , \11549 , \11552 , \11555 , \11558 );
and \U$10738 ( \11560 , \7950 , RIb54dd08_122);
and \U$10739 ( \11561 , RIb54dc90_121, \7917 );
nor \U$10740 ( \11562 , \11560 , \11561 );
not \U$10741 ( \11563 , \11562 );
nor \U$10742 ( \11564 , \11546 , \11559 , \11563 );
and \U$10743 ( \11565 , \7948 , RIb54e2a8_134);
and \U$10744 ( \11566 , RIb54e050_129, \7955 );
nor \U$10745 ( \11567 , \11565 , \11566 );
and \U$10746 ( \11568 , \7926 , RIb54dfd8_128);
and \U$10747 ( \11569 , RIb54df60_127, \7910 );
nor \U$10748 ( \11570 , \11568 , \11569 );
nand \U$10749 ( \11571 , \11564 , \11567 , \8206 , \11570 );
buf \U$10750 ( \11572 , \11571 );
_DC g24b6 ( \11573_nG24b6 , \11572 , \11369 );
xor \U$10751 ( \11574 , \8194 , \11573_nG24b6 );
and \U$10752 ( \11575 , \11341 , RIb54e410_137);
and \U$10753 ( \11576 , \7943 , RIb54e8c0_147);
and \U$10754 ( \11577 , RIb54e848_146, \7955 );
nor \U$10755 ( \11578 , \11576 , \11577 );
and \U$10756 ( \11579 , \7914 , RIb54e6e0_143);
and \U$10757 ( \11580 , RIb54e668_142, \7906 );
nor \U$10758 ( \11581 , \11579 , \11580 );
and \U$10759 ( \11582 , \7953 , RIb54e5f0_141);
and \U$10760 ( \11583 , RIb54e578_140, \7900 );
nor \U$10761 ( \11584 , \11582 , \11583 );
and \U$10762 ( \11585 , \7926 , RIb54e7d0_145);
and \U$10763 ( \11586 , RIb54e758_144, \7910 );
nor \U$10764 ( \11587 , \11585 , \11586 );
nand \U$10765 ( \11588 , \11578 , \11581 , \11584 , \11587 );
and \U$10766 ( \11589 , \7950 , RIb54e500_139);
and \U$10767 ( \11590 , RIb54e488_138, \7917 );
nor \U$10768 ( \11591 , \11589 , \11590 );
not \U$10769 ( \11592 , \11591 );
nor \U$10770 ( \11593 , \11575 , \11588 , \11592 );
and \U$10771 ( \11594 , \7948 , RIb54eaa0_151);
and \U$10772 ( \11595 , RIb54ea28_150, \7936 );
nor \U$10773 ( \11596 , \11594 , \11595 );
and \U$10774 ( \11597 , \7938 , RIb54e9b0_149);
and \U$10775 ( \11598 , RIb54e938_148, \7945 );
nor \U$10776 ( \11599 , \11597 , \11598 );
nand \U$10777 ( \11600 , \11593 , \11596 , \8248 , \11599 );
buf \U$10778 ( \11601 , \11600 );
_DC g24b4 ( \11602_nG24b4 , \11601 , \11369 );
xor \U$10779 ( \11603 , \8232 , \11602_nG24b4 );
and \U$10780 ( \11604 , \11341 , RIb54ec08_154);
and \U$10781 ( \11605 , \7943 , RIb54f0b8_164);
and \U$10782 ( \11606 , RIb54f040_163, \7955 );
nor \U$10783 ( \11607 , \11605 , \11606 );
and \U$10784 ( \11608 , \7914 , RIb54eed8_160);
and \U$10785 ( \11609 , RIb54ee60_159, \7906 );
nor \U$10786 ( \11610 , \11608 , \11609 );
and \U$10787 ( \11611 , \7953 , RIb54ede8_158);
and \U$10788 ( \11612 , RIb54ed70_157, \7900 );
nor \U$10789 ( \11613 , \11611 , \11612 );
and \U$10790 ( \11614 , \7926 , RIb54efc8_162);
and \U$10791 ( \11615 , RIb54ef50_161, \7910 );
nor \U$10792 ( \11616 , \11614 , \11615 );
nand \U$10793 ( \11617 , \11607 , \11610 , \11613 , \11616 );
and \U$10794 ( \11618 , \7950 , RIb54ecf8_156);
and \U$10795 ( \11619 , RIb54ec80_155, \7917 );
nor \U$10796 ( \11620 , \11618 , \11619 );
not \U$10797 ( \11621 , \11620 );
nor \U$10798 ( \11622 , \11604 , \11617 , \11621 );
and \U$10799 ( \11623 , \7948 , RIb54f298_168);
and \U$10800 ( \11624 , RIb54f220_167, \7936 );
nor \U$10801 ( \11625 , \11623 , \11624 );
and \U$10802 ( \11626 , \7938 , RIb54f1a8_166);
and \U$10803 ( \11627 , RIb54f130_165, \7945 );
nor \U$10804 ( \11628 , \11626 , \11627 );
nand \U$10805 ( \11629 , \11622 , \11625 , \8280 , \11628 );
buf \U$10806 ( \11630 , \11629 );
_DC g23de ( \11631_nG23de , \11630 , \11369 );
xor \U$10807 ( \11632 , \8268 , \11631_nG23de );
and \U$10808 ( \11633 , \11341 , RIb54f400_171);
and \U$10809 ( \11634 , \7943 , RIb54f8b0_181);
and \U$10810 ( \11635 , RIb54f838_180, \7955 );
nor \U$10811 ( \11636 , \11634 , \11635 );
and \U$10812 ( \11637 , \7914 , RIb54f6d0_177);
and \U$10813 ( \11638 , RIb54f658_176, \7906 );
nor \U$10814 ( \11639 , \11637 , \11638 );
and \U$10815 ( \11640 , \7953 , RIb54f5e0_175);
and \U$10816 ( \11641 , RIb54f568_174, \7900 );
nor \U$10817 ( \11642 , \11640 , \11641 );
and \U$10818 ( \11643 , \7926 , RIb54f7c0_179);
and \U$10819 ( \11644 , RIb54f748_178, \7910 );
nor \U$10820 ( \11645 , \11643 , \11644 );
nand \U$10821 ( \11646 , \11636 , \11639 , \11642 , \11645 );
and \U$10822 ( \11647 , \7950 , RIb54f4f0_173);
and \U$10823 ( \11648 , RIb54f478_172, \7917 );
nor \U$10824 ( \11649 , \11647 , \11648 );
not \U$10825 ( \11650 , \11649 );
nor \U$10826 ( \11651 , \11633 , \11646 , \11650 );
and \U$10827 ( \11652 , \7948 , RIb54fa90_185);
and \U$10828 ( \11653 , RIb54fa18_184, \7936 );
nor \U$10829 ( \11654 , \11652 , \11653 );
and \U$10830 ( \11655 , \7938 , RIb54f9a0_183);
and \U$10831 ( \11656 , RIb54f928_182, \7945 );
nor \U$10832 ( \11657 , \11655 , \11656 );
nand \U$10833 ( \11658 , \11651 , \11654 , \8318 , \11657 );
buf \U$10834 ( \11659 , \11658 );
_DC g23e0 ( \11660_nG23e0 , \11659 , \11369 );
xor \U$10835 ( \11661 , \8302 , \11660_nG23e0 );
and \U$10836 ( \11662 , \11341 , RIb54fbf8_188);
and \U$10837 ( \11663 , \7943 , RIb5500a8_198);
and \U$10838 ( \11664 , RIb550030_197, \7955 );
nor \U$10839 ( \11665 , \11663 , \11664 );
and \U$10840 ( \11666 , \7914 , RIb54fec8_194);
and \U$10841 ( \11667 , RIb54fe50_193, \7906 );
nor \U$10842 ( \11668 , \11666 , \11667 );
and \U$10843 ( \11669 , \7953 , RIb54fdd8_192);
and \U$10844 ( \11670 , RIb54fd60_191, \7900 );
nor \U$10845 ( \11671 , \11669 , \11670 );
and \U$10846 ( \11672 , \7926 , RIb54ffb8_196);
and \U$10847 ( \11673 , RIb54ff40_195, \7910 );
nor \U$10848 ( \11674 , \11672 , \11673 );
nand \U$10849 ( \11675 , \11665 , \11668 , \11671 , \11674 );
and \U$10850 ( \11676 , \7950 , RIb54fce8_190);
and \U$10851 ( \11677 , RIb54fc70_189, \7917 );
nor \U$10852 ( \11678 , \11676 , \11677 );
not \U$10853 ( \11679 , \11678 );
nor \U$10854 ( \11680 , \11662 , \11675 , \11679 );
and \U$10855 ( \11681 , \7948 , RIb550288_202);
and \U$10856 ( \11682 , RIb550210_201, \7936 );
nor \U$10857 ( \11683 , \11681 , \11682 );
and \U$10858 ( \11684 , \7938 , RIb550198_200);
and \U$10859 ( \11685 , RIb550120_199, \7945 );
nor \U$10860 ( \11686 , \11684 , \11685 );
nand \U$10861 ( \11687 , \11680 , \11683 , \8349 , \11686 );
buf \U$10862 ( \11688 , \11687 );
_DC g2277 ( \11689_nG2277 , \11688 , \11369 );
xor \U$10863 ( \11690 , RIb55bca0_599, \11689_nG2277 );
and \U$10864 ( \11691 , \11341 , RIb550468_206);
and \U$10865 ( \11692 , \7943 , RIb550918_216);
and \U$10866 ( \11693 , RIb5508a0_215, \7955 );
nor \U$10867 ( \11694 , \11692 , \11693 );
and \U$10868 ( \11695 , \7914 , RIb550738_212);
and \U$10869 ( \11696 , RIb5506c0_211, \7906 );
nor \U$10870 ( \11697 , \11695 , \11696 );
and \U$10871 ( \11698 , \7953 , RIb550648_210);
and \U$10872 ( \11699 , RIb5505d0_209, \7900 );
nor \U$10873 ( \11700 , \11698 , \11699 );
and \U$10874 ( \11701 , \7926 , RIb550828_214);
and \U$10875 ( \11702 , RIb5507b0_213, \7910 );
nor \U$10876 ( \11703 , \11701 , \11702 );
nand \U$10877 ( \11704 , \11694 , \11697 , \11700 , \11703 );
and \U$10878 ( \11705 , \7950 , RIb550558_208);
and \U$10879 ( \11706 , RIb5504e0_207, \7917 );
nor \U$10880 ( \11707 , \11705 , \11706 );
not \U$10881 ( \11708 , \11707 );
nor \U$10882 ( \11709 , \11691 , \11704 , \11708 );
and \U$10883 ( \11710 , \7948 , RIb550af8_220);
and \U$10884 ( \11711 , RIb550a80_219, \7936 );
nor \U$10885 ( \11712 , \11710 , \11711 );
and \U$10886 ( \11713 , \7938 , RIb550a08_218);
and \U$10887 ( \11714 , RIb550990_217, \7945 );
nor \U$10888 ( \11715 , \11713 , \11714 );
nand \U$10889 ( \11716 , \11709 , \11712 , \8380 , \11715 );
buf \U$10890 ( \11717 , \11716 );
_DC g2275 ( \11718_nG2275 , \11717 , \11369 );
nand \U$10891 ( \11719 , \11718_nG2275 , \8395 );
not \U$10892 ( \11720 , \11719 );
and \U$10893 ( \11721 , \11690 , \11720 );
and \U$10894 ( \11722 , RIb55bca0_599, \11689_nG2277 );
or \U$10895 ( \11723 , \11721 , \11722 );
and \U$10896 ( \11724 , \11661 , \11723 );
and \U$10897 ( \11725 , \8302 , \11660_nG23e0 );
or \U$10898 ( \11726 , \11724 , \11725 );
and \U$10899 ( \11727 , \11632 , \11726 );
and \U$10900 ( \11728 , \8268 , \11631_nG23de );
or \U$10901 ( \11729 , \11727 , \11728 );
and \U$10902 ( \11730 , \11603 , \11729 );
and \U$10903 ( \11731 , \8232 , \11602_nG24b4 );
or \U$10904 ( \11732 , \11730 , \11731 );
and \U$10905 ( \11733 , \11574 , \11732 );
and \U$10906 ( \11734 , \8194 , \11573_nG24b6 );
or \U$10907 ( \11735 , \11733 , \11734 );
and \U$10908 ( \11736 , \11545 , \11735 );
and \U$10909 ( \11737 , \8156 , \11544_nG25e4 );
or \U$10910 ( \11738 , \11736 , \11737 );
and \U$10911 ( \11739 , \11516 , \11738 );
and \U$10912 ( \11740 , \8118 , \11515_nG25e6 );
or \U$10913 ( \11741 , \11739 , \11740 );
and \U$10914 ( \11742 , \11487 , \11741 );
and \U$10915 ( \11743 , \8082 , \11486_nG275a );
or \U$10916 ( \11744 , \11742 , \11743 );
and \U$10917 ( \11745 , \11458 , \11744 );
and \U$10918 ( \11746 , \8044 , \11457_nG275c );
or \U$10919 ( \11747 , \11745 , \11746 );
and \U$10920 ( \11748 , \11429 , \11747 );
and \U$10921 ( \11749 , \8006 , \11428_nG290f );
or \U$10922 ( \11750 , \11748 , \11749 );
and \U$10923 ( \11751 , \11400 , \11750 );
and \U$10924 ( \11752 , \7970 , \11399_nG2911 );
or \U$10925 ( \11753 , \11751 , \11752 );
and \U$10926 ( \11754 , \11371 , \11753 );
and \U$10927 ( \11755 , \7889 , \11370_nG2aeb );
or \U$10928 ( \11756 , \11754 , \11755 );
nor \U$10929 ( \11757 , \11756 , \8435 );
not \U$10930 ( \11758 , \11757 );
not \U$10931 ( \11759 , \11341 );
nand \U$10932 ( \11760 , \11759 , \8461 );
and \U$10933 ( \11761 , \11760 , RIb550be8_222);
and \U$10934 ( \11762 , RIb5514d0_241, \7945 );
nor \U$10935 ( \11763 , \11761 , \11762 );
and \U$10936 ( \11764 , \7936 , RIb5515c0_243);
and \U$10937 ( \11765 , RIb5513e0_239, \7955 );
nor \U$10938 ( \11766 , \11764 , \11765 );
and \U$10939 ( \11767 , \7950 , RIb551098_232);
and \U$10940 ( \11768 , RIb551110_233, \7900 );
nor \U$10941 ( \11769 , \11767 , \11768 );
and \U$10942 ( \11770 , \7917 , RIb551020_231);
and \U$10943 ( \11771 , \7938 , RIb551548_242);
and \U$10944 ( \11772 , RIb551458_240, \7943 );
nor \U$10945 ( \11773 , \11771 , \11772 );
and \U$10946 ( \11774 , \7906 , RIb551200_235);
and \U$10947 ( \11775 , RIb551188_234, \7953 );
nor \U$10948 ( \11776 , \11774 , \11775 );
and \U$10949 ( \11777 , \7948 , RIb551638_244);
and \U$10950 ( \11778 , RIb551368_238, \7926 );
nor \U$10951 ( \11779 , \11777 , \11778 );
and \U$10952 ( \11780 , \7914 , RIb551278_236);
and \U$10953 ( \11781 , RIb5512f0_237, \7910 );
nor \U$10954 ( \11782 , \11780 , \11781 );
nand \U$10955 ( \11783 , \11773 , \11776 , \11779 , \11782 );
nor \U$10956 ( \11784 , \11770 , \11783 );
nand \U$10957 ( \11785 , \11763 , \11766 , \11769 , \11784 );
buf \U$10958 ( \11786 , \7962 );
_DC g3124 ( \11787_nG3124 , \11785 , \11786 );
not \U$10959 ( \11788 , \11787_nG3124 );
nor \U$10960 ( \11789 , \11758 , \11788 );
xor \U$10961 ( \11790 , \7889 , \11370_nG2aeb );
xor \U$10962 ( \11791 , \11790 , \11753 );
not \U$10963 ( \11792 , \11791 );
xor \U$10964 ( \11793 , \7970 , \11399_nG2911 );
xor \U$10965 ( \11794 , \11793 , \11750 );
not \U$10966 ( \11795 , \11794 );
and \U$10967 ( \11796 , \11792 , \11795 );
and \U$10968 ( \11797 , \11756 , \8435 );
nor \U$10969 ( \11798 , \11797 , \11757 );
nor \U$10970 ( \11799 , \11796 , \11798 );
not \U$10971 ( \11800 , \11799 );
and \U$10972 ( \11801 , \11798 , \11791 );
nor \U$10973 ( \11802 , \11798 , \11791 );
xnor \U$10974 ( \11803 , \11794 , \11791 );
not \U$10975 ( \11804 , \11803 );
nor \U$10976 ( \11805 , \11801 , \11802 , \11804 );
nand \U$10977 ( \11806 , \11800 , \11805 );
and \U$10978 ( \11807 , \11760 , RIb552010_265);
and \U$10979 ( \11808 , RIb552628_278, \7936 );
nor \U$10980 ( \11809 , \11807 , \11808 );
and \U$10981 ( \11810 , \7938 , RIb5525b0_277);
and \U$10982 ( \11811 , RIb552448_274, \7955 );
nor \U$10983 ( \11812 , \11810 , \11811 );
and \U$10984 ( \11813 , \7950 , RIb552100_267);
and \U$10985 ( \11814 , RIb552178_268, \7900 );
nor \U$10986 ( \11815 , \11813 , \11814 );
and \U$10987 ( \11816 , \7917 , RIb552088_266);
and \U$10988 ( \11817 , \7906 , RIb552268_270);
and \U$10989 ( \11818 , RIb5521f0_269, \7953 );
nor \U$10990 ( \11819 , \11817 , \11818 );
and \U$10991 ( \11820 , \7914 , RIb5522e0_271);
and \U$10992 ( \11821 , RIb552358_272, \7910 );
nor \U$10993 ( \11822 , \11820 , \11821 );
and \U$10994 ( \11823 , \7948 , RIb5526a0_279);
and \U$10995 ( \11824 , RIb5523d0_273, \7926 );
nor \U$10996 ( \11825 , \11823 , \11824 );
and \U$10997 ( \11826 , \7943 , RIb5524c0_275);
and \U$10998 ( \11827 , RIb552538_276, \7945 );
nor \U$10999 ( \11828 , \11826 , \11827 );
nand \U$11000 ( \11829 , \11819 , \11822 , \11825 , \11828 );
nor \U$11001 ( \11830 , \11816 , \11829 );
nand \U$11002 ( \11831 , \11809 , \11812 , \11815 , \11830 );
_DC g323c ( \11832_nG323c , \11831 , \11786 );
not \U$11003 ( \11833 , \11832_nG323c );
or \U$11004 ( \11834 , \11806 , \11833 );
or \U$11005 ( \11835 , \11832_nG323c , \11800 );
or \U$11006 ( \11836 , \11805 , \11800 );
nand \U$11007 ( \11837 , \11834 , \11835 , \11836 );
xnor \U$11008 ( \11838 , \11789 , \11837 );
nand \U$11009 ( \11839 , \11804 , \11800 );
or \U$11010 ( \11840 , \11839 , \11833 );
or \U$11011 ( \11841 , \11788 , \11806 );
or \U$11012 ( \11842 , \11803 , \11833 );
or \U$11013 ( \11843 , \11800 , \11787_nG3124 );
nand \U$11014 ( \11844 , \11843 , \11836 );
nand \U$11015 ( \11845 , \11842 , \11844 );
nand \U$11016 ( \11846 , \11840 , \11841 , \11845 );
xor \U$11017 ( \11847 , \8006 , \11428_nG290f );
xor \U$11018 ( \11848 , \11847 , \11747 );
xor \U$11019 ( \11849 , \8044 , \11457_nG275c );
xor \U$11020 ( \11850 , \11849 , \11744 );
nor \U$11021 ( \11851 , \11848 , \11850 );
or \U$11022 ( \11852 , \11794 , \11851 );
and \U$11023 ( \11853 , \11846 , \11852 );
and \U$11024 ( \11854 , \11760 , RIb552808_282);
and \U$11025 ( \11855 , RIb552e20_295, \7936 );
nor \U$11026 ( \11856 , \11854 , \11855 );
and \U$11027 ( \11857 , \7938 , RIb552da8_294);
and \U$11028 ( \11858 , RIb552c40_291, \7955 );
nor \U$11029 ( \11859 , \11857 , \11858 );
and \U$11030 ( \11860 , \7950 , RIb5528f8_284);
and \U$11031 ( \11861 , RIb552970_285, \7900 );
nor \U$11032 ( \11862 , \11860 , \11861 );
and \U$11033 ( \11863 , \7917 , RIb552880_283);
and \U$11034 ( \11864 , \7906 , RIb552a60_287);
and \U$11035 ( \11865 , RIb5529e8_286, \7953 );
nor \U$11036 ( \11866 , \11864 , \11865 );
and \U$11037 ( \11867 , \7914 , RIb552ad8_288);
and \U$11038 ( \11868 , RIb552b50_289, \7910 );
nor \U$11039 ( \11869 , \11867 , \11868 );
and \U$11040 ( \11870 , \7948 , RIb552e98_296);
and \U$11041 ( \11871 , RIb552bc8_290, \7926 );
nor \U$11042 ( \11872 , \11870 , \11871 );
and \U$11043 ( \11873 , \7943 , RIb552cb8_292);
and \U$11044 ( \11874 , RIb552d30_293, \7945 );
nor \U$11045 ( \11875 , \11873 , \11874 );
nand \U$11046 ( \11876 , \11866 , \11869 , \11872 , \11875 );
nor \U$11047 ( \11877 , \11863 , \11876 );
nand \U$11048 ( \11878 , \11856 , \11859 , \11862 , \11877 );
_DC g301d ( \11879_nG301d , \11878 , \11786 );
nand \U$11049 ( \11880 , \11879_nG301d , \11757 );
not \U$11050 ( \11881 , \11880 );
nor \U$11051 ( \11882 , \11853 , \11881 );
xor \U$11052 ( \11883 , \11838 , \11882 );
not \U$11053 ( \11884 , \11883 );
not \U$11054 ( \11885 , \11848 );
not \U$11055 ( \11886 , \11794 );
or \U$11056 ( \11887 , \11885 , \11886 );
or \U$11057 ( \11888 , \11794 , \11848 );
nand \U$11058 ( \11889 , \11887 , \11888 );
xor \U$11059 ( \11890 , \11850 , \11848 );
nor \U$11060 ( \11891 , \11889 , \11890 );
not \U$11061 ( \11892 , \11891 );
not \U$11062 ( \11893 , \11852 );
nor \U$11063 ( \11894 , \11892 , \11893 );
not \U$11064 ( \11895 , \11894 );
or \U$11065 ( \11896 , \11895 , \11833 );
or \U$11066 ( \11897 , \11892 , \11833 );
nand \U$11067 ( \11898 , \11897 , \11893 );
nand \U$11068 ( \11899 , \11896 , \11898 );
or \U$11069 ( \11900 , \11839 , \11788 );
not \U$11070 ( \11901 , \11879_nG301d );
or \U$11071 ( \11902 , \11901 , \11806 );
or \U$11072 ( \11903 , \11803 , \11788 );
or \U$11073 ( \11904 , \11800 , \11879_nG301d );
nand \U$11074 ( \11905 , \11904 , \11836 );
nand \U$11075 ( \11906 , \11903 , \11905 );
nand \U$11076 ( \11907 , \11900 , \11902 , \11906 );
and \U$11077 ( \11908 , \11899 , \11907 );
not \U$11078 ( \11909 , \11880 );
and \U$11079 ( \11910 , \11846 , \11852 );
not \U$11080 ( \11911 , \11846 );
and \U$11081 ( \11912 , \11911 , \11893 );
nor \U$11082 ( \11913 , \11910 , \11912 );
not \U$11083 ( \11914 , \11913 );
or \U$11084 ( \11915 , \11909 , \11914 );
or \U$11085 ( \11916 , \11913 , \11880 );
nand \U$11086 ( \11917 , \11915 , \11916 );
and \U$11087 ( \11918 , \11908 , \11917 );
and \U$11088 ( \11919 , \11884 , \11918 );
or \U$11089 ( \11920 , \11919 , \11799 );
and \U$11090 ( \11921 , \11919 , \11799 );
and \U$11091 ( \11922 , \11789 , \11837 );
nor \U$11092 ( \11923 , \11921 , \11922 );
nand \U$11093 ( \11924 , \11920 , \11923 );
not \U$11094 ( \11925 , \11924 );
and \U$11095 ( \11926 , \11757 , \11832_nG323c );
and \U$11096 ( \11927 , \11838 , \11882 );
nor \U$11097 ( \11928 , \11926 , \11927 );
not \U$11098 ( \11929 , \11928 );
and \U$11099 ( \11930 , \11925 , \11929 );
and \U$11100 ( \11931 , \11924 , \11928 );
nor \U$11101 ( \11932 , \11930 , \11931 );
not \U$11102 ( \11933 , \11932 );
xor \U$11103 ( \11934 , \11884 , \11918 );
and \U$11104 ( \11935 , \11787_nG3124 , \11894 );
and \U$11105 ( \11936 , \11852 , \11890 );
and \U$11106 ( \11937 , \11936 , \11832_nG323c );
nand \U$11107 ( \11938 , \11787_nG3124 , \11891 );
or \U$11108 ( \11939 , \11852 , \11832_nG323c );
or \U$11109 ( \11940 , \11852 , \11890 );
nand \U$11110 ( \11941 , \11939 , \11940 );
and \U$11111 ( \11942 , \11938 , \11941 );
nor \U$11112 ( \11943 , \11935 , \11937 , \11942 );
not \U$11113 ( \11944 , \11839 );
and \U$11114 ( \11945 , \11879_nG301d , \11944 );
not \U$11115 ( \11946 , \11806 );
and \U$11116 ( \11947 , \11760 , RIb5537f8_316);
and \U$11117 ( \11948 , RIb553e10_329, \7936 );
nor \U$11118 ( \11949 , \11947 , \11948 );
and \U$11119 ( \11950 , \7938 , RIb553d98_328);
and \U$11120 ( \11951 , RIb553c30_325, \7955 );
nor \U$11121 ( \11952 , \11950 , \11951 );
and \U$11122 ( \11953 , \7950 , RIb5538e8_318);
and \U$11123 ( \11954 , RIb553960_319, \7900 );
nor \U$11124 ( \11955 , \11953 , \11954 );
and \U$11125 ( \11956 , \7917 , RIb553870_317);
and \U$11126 ( \11957 , \7943 , RIb553ca8_326);
and \U$11127 ( \11958 , RIb553bb8_324, \7926 );
nor \U$11128 ( \11959 , \11957 , \11958 );
and \U$11129 ( \11960 , \7914 , RIb553ac8_322);
and \U$11130 ( \11961 , RIb553b40_323, \7910 );
nor \U$11131 ( \11962 , \11960 , \11961 );
and \U$11132 ( \11963 , \7948 , RIb553e88_330);
and \U$11133 ( \11964 , RIb553d20_327, \7945 );
nor \U$11134 ( \11965 , \11963 , \11964 );
and \U$11135 ( \11966 , \7906 , RIb553a50_321);
and \U$11136 ( \11967 , RIb5539d8_320, \7953 );
nor \U$11137 ( \11968 , \11966 , \11967 );
nand \U$11138 ( \11969 , \11959 , \11962 , \11965 , \11968 );
nor \U$11139 ( \11970 , \11956 , \11969 );
nand \U$11140 ( \11971 , \11949 , \11952 , \11955 , \11970 );
_DC g2efb ( \11972_nG2efb , \11971 , \11786 );
and \U$11141 ( \11973 , \11946 , \11972_nG2efb );
nand \U$11142 ( \11974 , \11879_nG301d , \11804 );
or \U$11143 ( \11975 , \11800 , \11972_nG2efb );
nand \U$11144 ( \11976 , \11975 , \11836 );
and \U$11145 ( \11977 , \11974 , \11976 );
nor \U$11146 ( \11978 , \11945 , \11973 , \11977 );
nand \U$11147 ( \11979 , \11943 , \11978 );
xor \U$11148 ( \11980 , \8082 , \11486_nG275a );
xor \U$11149 ( \11981 , \11980 , \11741 );
xor \U$11150 ( \11982 , \8118 , \11515_nG25e6 );
xor \U$11151 ( \11983 , \11982 , \11738 );
nor \U$11152 ( \11984 , \11981 , \11983 );
or \U$11153 ( \11985 , \11850 , \11984 );
and \U$11154 ( \11986 , \11979 , \11985 );
nor \U$11155 ( \11987 , \11978 , \11943 );
nor \U$11156 ( \11988 , \11986 , \11987 );
xor \U$11157 ( \11989 , \11899 , \11907 );
not \U$11158 ( \11990 , \11989 );
nand \U$11159 ( \11991 , \11972_nG2efb , \11757 );
not \U$11160 ( \11992 , \11991 );
and \U$11161 ( \11993 , \11990 , \11992 );
and \U$11162 ( \11994 , \11989 , \11991 );
nor \U$11163 ( \11995 , \11993 , \11994 );
nand \U$11164 ( \11996 , \11988 , \11995 );
xor \U$11165 ( \11997 , \11908 , \11917 );
and \U$11166 ( \11998 , \11996 , \11997 );
and \U$11167 ( \11999 , \11934 , \11998 );
not \U$11168 ( \12000 , \11999 );
and \U$11169 ( \12001 , \11933 , \12000 );
and \U$11170 ( \12002 , \11932 , \11999 );
nor \U$11171 ( \12003 , \12001 , \12002 );
not \U$11172 ( \12004 , \12003 );
not \U$11173 ( \12005 , \11985 );
not \U$11174 ( \12006 , \11987 );
nand \U$11175 ( \12007 , \12006 , \11979 );
not \U$11176 ( \12008 , \12007 );
or \U$11177 ( \12009 , \12005 , \12008 );
or \U$11178 ( \12010 , \12007 , \11985 );
nand \U$11179 ( \12011 , \12009 , \12010 );
not \U$11180 ( \12012 , \12011 );
and \U$11181 ( \12013 , \11760 , RIb553000_299);
and \U$11182 ( \12014 , RIb553618_312, \7936 );
nor \U$11183 ( \12015 , \12013 , \12014 );
and \U$11184 ( \12016 , \7938 , RIb5535a0_311);
and \U$11185 ( \12017 , RIb553438_308, \7955 );
nor \U$11186 ( \12018 , \12016 , \12017 );
and \U$11187 ( \12019 , \7950 , RIb5530f0_301);
and \U$11188 ( \12020 , RIb553168_302, \7900 );
nor \U$11189 ( \12021 , \12019 , \12020 );
and \U$11190 ( \12022 , \7917 , RIb553078_300);
and \U$11191 ( \12023 , \7906 , RIb553258_304);
and \U$11192 ( \12024 , RIb5531e0_303, \7953 );
nor \U$11193 ( \12025 , \12023 , \12024 );
and \U$11194 ( \12026 , \7943 , RIb5534b0_309);
and \U$11195 ( \12027 , RIb553528_310, \7945 );
nor \U$11196 ( \12028 , \12026 , \12027 );
and \U$11197 ( \12029 , \7948 , RIb553690_313);
and \U$11198 ( \12030 , RIb5533c0_307, \7926 );
nor \U$11199 ( \12031 , \12029 , \12030 );
and \U$11200 ( \12032 , \7914 , RIb5532d0_305);
and \U$11201 ( \12033 , RIb553348_306, \7910 );
nor \U$11202 ( \12034 , \12032 , \12033 );
nand \U$11203 ( \12035 , \12025 , \12028 , \12031 , \12034 );
nor \U$11204 ( \12036 , \12022 , \12035 );
nand \U$11205 ( \12037 , \12015 , \12018 , \12021 , \12036 );
_DC g2e11 ( \12038_nG2e11 , \12037 , \11786 );
nand \U$11206 ( \12039 , \12038_nG2e11 , \11757 );
not \U$11207 ( \12040 , \12039 );
and \U$11208 ( \12041 , \12012 , \12040 );
and \U$11209 ( \12042 , \12011 , \12039 );
nor \U$11210 ( \12043 , \12041 , \12042 );
not \U$11211 ( \12044 , \12043 );
and \U$11212 ( \12045 , \11879_nG301d , \11894 );
and \U$11213 ( \12046 , \11936 , \11787_nG3124 );
nand \U$11214 ( \12047 , \11879_nG301d , \11891 );
or \U$11215 ( \12048 , \11852 , \11787_nG3124 );
nand \U$11216 ( \12049 , \12048 , \11940 );
and \U$11217 ( \12050 , \12047 , \12049 );
nor \U$11218 ( \12051 , \12045 , \12046 , \12050 );
and \U$11219 ( \12052 , \11850 , \11981 );
nor \U$11220 ( \12053 , \11850 , \11981 );
xor \U$11221 ( \12054 , \11981 , \11983 );
nor \U$11222 ( \12055 , \12052 , \12053 , \12054 );
and \U$11223 ( \12056 , \12055 , \11985 );
and \U$11224 ( \12057 , \11832_nG323c , \12056 );
not \U$11225 ( \12058 , \11985 );
and \U$11226 ( \12059 , \11833 , \12058 );
or \U$11227 ( \12060 , \12055 , \11985 );
not \U$11228 ( \12061 , \12060 );
nor \U$11229 ( \12062 , \12057 , \12059 , \12061 );
or \U$11230 ( \12063 , \12051 , \12062 );
and \U$11231 ( \12064 , \11760 , RIb553ff0_333);
and \U$11232 ( \12065 , RIb554608_346, \7936 );
nor \U$11233 ( \12066 , \12064 , \12065 );
and \U$11234 ( \12067 , \7938 , RIb554590_345);
and \U$11235 ( \12068 , RIb554428_342, \7955 );
nor \U$11236 ( \12069 , \12067 , \12068 );
and \U$11237 ( \12070 , \7950 , RIb5540e0_335);
and \U$11238 ( \12071 , RIb554158_336, \7900 );
nor \U$11239 ( \12072 , \12070 , \12071 );
and \U$11240 ( \12073 , \7917 , RIb554068_334);
and \U$11241 ( \12074 , \7906 , RIb554248_338);
and \U$11242 ( \12075 , RIb5541d0_337, \7953 );
nor \U$11243 ( \12076 , \12074 , \12075 );
and \U$11244 ( \12077 , \7914 , RIb5542c0_339);
and \U$11245 ( \12078 , RIb554338_340, \7910 );
nor \U$11246 ( \12079 , \12077 , \12078 );
and \U$11247 ( \12080 , \7948 , RIb554680_347);
and \U$11248 ( \12081 , RIb5543b0_341, \7926 );
nor \U$11249 ( \12082 , \12080 , \12081 );
and \U$11250 ( \12083 , \7943 , RIb5544a0_343);
and \U$11251 ( \12084 , RIb554518_344, \7945 );
nor \U$11252 ( \12085 , \12083 , \12084 );
nand \U$11253 ( \12086 , \12076 , \12079 , \12082 , \12085 );
nor \U$11254 ( \12087 , \12073 , \12086 );
nand \U$11255 ( \12088 , \12066 , \12069 , \12072 , \12087 );
_DC g2d11 ( \12089_nG2d11 , \12088 , \11786 );
nand \U$11256 ( \12090 , \12089_nG2d11 , \11757 );
and \U$11257 ( \12091 , \11972_nG2efb , \11944 );
and \U$11258 ( \12092 , \11946 , \12038_nG2e11 );
nand \U$11259 ( \12093 , \11972_nG2efb , \11804 );
or \U$11260 ( \12094 , \11800 , \12038_nG2e11 );
nand \U$11261 ( \12095 , \12094 , \11836 );
and \U$11262 ( \12096 , \12093 , \12095 );
nor \U$11263 ( \12097 , \12091 , \12092 , \12096 );
or \U$11264 ( \12098 , \12090 , \12097 );
nand \U$11265 ( \12099 , \12063 , \12098 );
nand \U$11266 ( \12100 , \12044 , \12099 );
not \U$11267 ( \12101 , \12100 );
or \U$11268 ( \12102 , \11995 , \11988 );
nand \U$11269 ( \12103 , \12102 , \11996 );
nand \U$11270 ( \12104 , \12101 , \12103 );
xor \U$11271 ( \12105 , \11996 , \11997 );
not \U$11272 ( \12106 , \11989 );
nor \U$11273 ( \12107 , \12106 , \11991 );
nor \U$11274 ( \12108 , \12105 , \12107 );
or \U$11275 ( \12109 , \12104 , \12108 );
nand \U$11276 ( \12110 , \12107 , \12105 );
nand \U$11277 ( \12111 , \12109 , \12110 );
xor \U$11278 ( \12112 , \11934 , \11998 );
and \U$11279 ( \12113 , \12111 , \12112 );
not \U$11280 ( \12114 , \12111 );
not \U$11281 ( \12115 , \12112 );
and \U$11282 ( \12116 , \12114 , \12115 );
and \U$11283 ( \12117 , \11760 , RIb554fe0_367);
and \U$11284 ( \12118 , RIb555418_376, \7955 );
nor \U$11285 ( \12119 , \12117 , \12118 );
and \U$11286 ( \12120 , \7926 , RIb5553a0_375);
and \U$11287 ( \12121 , RIb555328_374, \7910 );
nor \U$11288 ( \12122 , \12120 , \12121 );
and \U$11289 ( \12123 , \7906 , RIb555238_372);
and \U$11290 ( \12124 , RIb5551c0_371, \7953 );
nor \U$11291 ( \12125 , \12123 , \12124 );
and \U$11292 ( \12126 , \7914 , RIb5552b0_373);
and \U$11293 ( \12127 , \7943 , RIb555490_377);
and \U$11294 ( \12128 , RIb555508_378, \7945 );
nor \U$11295 ( \12129 , \12127 , \12128 );
and \U$11296 ( \12130 , \7950 , RIb5550d0_369);
and \U$11297 ( \12131 , RIb555058_368, \7917 );
nor \U$11298 ( \12132 , \12130 , \12131 );
and \U$11299 ( \12133 , \7948 , RIb555670_381);
and \U$11300 ( \12134 , RIb555148_370, \7900 );
nor \U$11301 ( \12135 , \12133 , \12134 );
and \U$11302 ( \12136 , \7936 , RIb5555f8_380);
and \U$11303 ( \12137 , RIb555580_379, \7938 );
nor \U$11304 ( \12138 , \12136 , \12137 );
nand \U$11305 ( \12139 , \12129 , \12132 , \12135 , \12138 );
nor \U$11306 ( \12140 , \12126 , \12139 );
nand \U$11307 ( \12141 , \12119 , \12122 , \12125 , \12140 );
_DC g2c0d ( \12142_nG2c0d , \12141 , \11786 );
and \U$11308 ( \12143 , \12142_nG2c0d , \11944 );
and \U$11309 ( \12144 , \11760 , RIb5547e8_350);
and \U$11310 ( \12145 , RIb554e00_363, \7936 );
nor \U$11311 ( \12146 , \12144 , \12145 );
and \U$11312 ( \12147 , \7938 , RIb554d88_362);
and \U$11313 ( \12148 , RIb554c20_359, \7955 );
nor \U$11314 ( \12149 , \12147 , \12148 );
and \U$11315 ( \12150 , \7950 , RIb5548d8_352);
and \U$11316 ( \12151 , RIb554950_353, \7900 );
nor \U$11317 ( \12152 , \12150 , \12151 );
and \U$11318 ( \12153 , \7917 , RIb554860_351);
and \U$11319 ( \12154 , \7914 , RIb554ab8_356);
and \U$11320 ( \12155 , RIb554b30_357, \7910 );
nor \U$11321 ( \12156 , \12154 , \12155 );
and \U$11322 ( \12157 , \7906 , RIb554a40_355);
and \U$11323 ( \12158 , RIb5549c8_354, \7953 );
nor \U$11324 ( \12159 , \12157 , \12158 );
and \U$11325 ( \12160 , \7948 , RIb554e78_364);
and \U$11326 ( \12161 , RIb554ba8_358, \7926 );
nor \U$11327 ( \12162 , \12160 , \12161 );
and \U$11328 ( \12163 , \7943 , RIb554c98_360);
and \U$11329 ( \12164 , RIb554d10_361, \7945 );
nor \U$11330 ( \12165 , \12163 , \12164 );
nand \U$11331 ( \12166 , \12156 , \12159 , \12162 , \12165 );
nor \U$11332 ( \12167 , \12153 , \12166 );
nand \U$11333 ( \12168 , \12146 , \12149 , \12152 , \12167 );
_DC g2b05 ( \12169_nG2b05 , \12168 , \11786 );
and \U$11334 ( \12170 , \11946 , \12169_nG2b05 );
nand \U$11335 ( \12171 , \12142_nG2c0d , \11804 );
or \U$11336 ( \12172 , \11800 , \12169_nG2b05 );
nand \U$11337 ( \12173 , \12172 , \11836 );
and \U$11338 ( \12174 , \12171 , \12173 );
nor \U$11339 ( \12175 , \12143 , \12170 , \12174 );
and \U$11340 ( \12176 , \12089_nG2d11 , \11894 );
and \U$11341 ( \12177 , \11936 , \12038_nG2e11 );
nand \U$11342 ( \12178 , \12089_nG2d11 , \11891 );
or \U$11343 ( \12179 , \11852 , \12038_nG2e11 );
nand \U$11344 ( \12180 , \12179 , \11940 );
and \U$11345 ( \12181 , \12178 , \12180 );
nor \U$11346 ( \12182 , \12176 , \12177 , \12181 );
and \U$11347 ( \12183 , \12175 , \12182 );
not \U$11348 ( \12184 , \12183 );
and \U$11349 ( \12185 , \11760 , RIb555fd0_401);
and \U$11350 ( \12186 , RIb5565e8_414, \7936 );
nor \U$11351 ( \12187 , \12185 , \12186 );
and \U$11352 ( \12188 , \7938 , RIb556570_413);
and \U$11353 ( \12189 , RIb556408_410, \7955 );
nor \U$11354 ( \12190 , \12188 , \12189 );
and \U$11355 ( \12191 , \7950 , RIb5560c0_403);
and \U$11356 ( \12192 , RIb556138_404, \7900 );
nor \U$11357 ( \12193 , \12191 , \12192 );
and \U$11358 ( \12194 , \7917 , RIb556048_402);
and \U$11359 ( \12195 , \7906 , RIb556228_406);
and \U$11360 ( \12196 , RIb5561b0_405, \7953 );
nor \U$11361 ( \12197 , \12195 , \12196 );
and \U$11362 ( \12198 , \7943 , RIb556480_411);
and \U$11363 ( \12199 , RIb5564f8_412, \7945 );
nor \U$11364 ( \12200 , \12198 , \12199 );
and \U$11365 ( \12201 , \7948 , RIb556660_415);
and \U$11366 ( \12202 , RIb556390_409, \7926 );
nor \U$11367 ( \12203 , \12201 , \12202 );
and \U$11368 ( \12204 , \7914 , RIb5562a0_407);
and \U$11369 ( \12205 , RIb556318_408, \7910 );
nor \U$11370 ( \12206 , \12204 , \12205 );
nand \U$11371 ( \12207 , \12197 , \12200 , \12203 , \12206 );
nor \U$11372 ( \12208 , \12194 , \12207 );
nand \U$11373 ( \12209 , \12187 , \12190 , \12193 , \12208 );
_DC g2a23 ( \12210_nG2a23 , \12209 , \11786 );
nand \U$11374 ( \12211 , \12210_nG2a23 , \11757 );
not \U$11375 ( \12212 , \12211 );
and \U$11376 ( \12213 , \12184 , \12212 );
nor \U$11377 ( \12214 , \12175 , \12182 );
nor \U$11378 ( \12215 , \12213 , \12214 );
xor \U$11379 ( \12216 , \8156 , \11544_nG25e4 );
xor \U$11380 ( \12217 , \12216 , \11735 );
not \U$11381 ( \12218 , \12217 );
not \U$11382 ( \12219 , \11983 );
or \U$11383 ( \12220 , \12218 , \12219 );
or \U$11384 ( \12221 , \11983 , \12217 );
nand \U$11385 ( \12222 , \12220 , \12221 );
xor \U$11386 ( \12223 , \8194 , \11573_nG24b6 );
xor \U$11387 ( \12224 , \12223 , \11732 );
xor \U$11388 ( \12225 , \12224 , \12217 );
nor \U$11389 ( \12226 , \12222 , \12225 );
nand \U$11390 ( \12227 , \11787_nG3124 , \12226 );
nor \U$11391 ( \12228 , \12217 , \12224 );
or \U$11392 ( \12229 , \11983 , \12228 );
or \U$11393 ( \12230 , \12229 , \11832_nG323c );
or \U$11394 ( \12231 , \12229 , \12225 );
nand \U$11395 ( \12232 , \12230 , \12231 );
and \U$11396 ( \12233 , \12227 , \12232 );
and \U$11397 ( \12234 , \12229 , \12225 );
and \U$11398 ( \12235 , \12234 , \11832_nG323c );
not \U$11399 ( \12236 , \12226 );
not \U$11400 ( \12237 , \12229 );
nor \U$11401 ( \12238 , \12236 , \12237 );
and \U$11402 ( \12239 , \11787_nG3124 , \12238 );
nor \U$11403 ( \12240 , \12233 , \12235 , \12239 );
nand \U$11404 ( \12241 , \11879_nG301d , \12054 );
or \U$11405 ( \12242 , \11985 , \11972_nG2efb );
nand \U$11406 ( \12243 , \12242 , \12060 );
and \U$11407 ( \12244 , \12241 , \12243 );
and \U$11408 ( \12245 , \12056 , \11972_nG2efb );
not \U$11409 ( \12246 , \12054 );
nor \U$11410 ( \12247 , \12058 , \12246 );
and \U$11411 ( \12248 , \11879_nG301d , \12247 );
nor \U$11412 ( \12249 , \12244 , \12245 , \12248 );
nand \U$11413 ( \12250 , \12240 , \12249 );
xor \U$11414 ( \12251 , \8268 , \11631_nG23de );
xor \U$11415 ( \12252 , \12251 , \11726 );
not \U$11416 ( \12253 , \12252 );
xor \U$11417 ( \12254 , \8232 , \11602_nG24b4 );
xor \U$11418 ( \12255 , \12254 , \11729 );
not \U$11419 ( \12256 , \12255 );
and \U$11420 ( \12257 , \12253 , \12256 );
or \U$11421 ( \12258 , \12257 , \12224 );
and \U$11422 ( \12259 , \12250 , \12258 );
nor \U$11423 ( \12260 , \12249 , \12240 );
nor \U$11424 ( \12261 , \12259 , \12260 );
nor \U$11425 ( \12262 , \12215 , \12261 );
not \U$11426 ( \12263 , \12238 );
or \U$11427 ( \12264 , \12263 , \11833 );
or \U$11428 ( \12265 , \12236 , \11833 );
nand \U$11429 ( \12266 , \12265 , \12237 );
nand \U$11430 ( \12267 , \12264 , \12266 );
not \U$11431 ( \12268 , \12247 );
or \U$11432 ( \12269 , \12268 , \11788 );
not \U$11433 ( \12270 , \12056 );
or \U$11434 ( \12271 , \11901 , \12270 );
or \U$11435 ( \12272 , \12246 , \11788 );
or \U$11436 ( \12273 , \11985 , \11879_nG301d );
nand \U$11437 ( \12274 , \12273 , \12060 );
nand \U$11438 ( \12275 , \12272 , \12274 );
nand \U$11439 ( \12276 , \12269 , \12271 , \12275 );
xor \U$11440 ( \12277 , \12267 , \12276 );
not \U$11441 ( \12278 , \12277 );
and \U$11442 ( \12279 , \12089_nG2d11 , \11944 );
and \U$11443 ( \12280 , \11946 , \12142_nG2c0d );
nand \U$11444 ( \12281 , \12089_nG2d11 , \11804 );
or \U$11445 ( \12282 , \11800 , \12142_nG2c0d );
nand \U$11446 ( \12283 , \12282 , \11836 );
and \U$11447 ( \12284 , \12281 , \12283 );
nor \U$11448 ( \12285 , \12279 , \12280 , \12284 );
and \U$11449 ( \12286 , \12038_nG2e11 , \11894 );
and \U$11450 ( \12287 , \11936 , \11972_nG2efb );
nand \U$11451 ( \12288 , \12038_nG2e11 , \11891 );
or \U$11452 ( \12289 , \11852 , \11972_nG2efb );
nand \U$11453 ( \12290 , \12289 , \11940 );
and \U$11454 ( \12291 , \12288 , \12290 );
nor \U$11455 ( \12292 , \12286 , \12287 , \12291 );
or \U$11456 ( \12293 , \12285 , \12292 );
not \U$11457 ( \12294 , \12293 );
and \U$11458 ( \12295 , \12285 , \12292 );
nor \U$11459 ( \12296 , \12294 , \12295 );
not \U$11460 ( \12297 , \12296 );
nand \U$11461 ( \12298 , \12169_nG2b05 , \11757 );
not \U$11462 ( \12299 , \12298 );
and \U$11463 ( \12300 , \12297 , \12299 );
and \U$11464 ( \12301 , \12296 , \12298 );
nor \U$11465 ( \12302 , \12300 , \12301 );
nor \U$11466 ( \12303 , \12278 , \12302 );
and \U$11467 ( \12304 , \12262 , \12303 );
not \U$11468 ( \12305 , \12229 );
and \U$11469 ( \12306 , \11972_nG2efb , \11894 );
and \U$11470 ( \12307 , \11936 , \11879_nG301d );
nand \U$11471 ( \12308 , \11972_nG2efb , \11891 );
or \U$11472 ( \12309 , \11852 , \11879_nG301d );
nand \U$11473 ( \12310 , \12309 , \11940 );
and \U$11474 ( \12311 , \12308 , \12310 );
nor \U$11475 ( \12312 , \12306 , \12307 , \12311 );
nand \U$11476 ( \12313 , \11832_nG323c , \12054 );
or \U$11477 ( \12314 , \11985 , \11787_nG3124 );
nand \U$11478 ( \12315 , \12314 , \12060 );
and \U$11479 ( \12316 , \12313 , \12315 );
and \U$11480 ( \12317 , \12056 , \11787_nG3124 );
and \U$11481 ( \12318 , \11832_nG323c , \12247 );
nor \U$11482 ( \12319 , \12316 , \12317 , \12318 );
nor \U$11483 ( \12320 , \12312 , \12319 );
not \U$11484 ( \12321 , \12320 );
nand \U$11485 ( \12322 , \12319 , \12312 );
nand \U$11486 ( \12323 , \12321 , \12322 );
not \U$11487 ( \12324 , \12323 );
or \U$11488 ( \12325 , \12305 , \12324 );
or \U$11489 ( \12326 , \12323 , \12229 );
nand \U$11490 ( \12327 , \12325 , \12326 );
not \U$11491 ( \12328 , \12142_nG2c0d );
nor \U$11492 ( \12329 , \11758 , \12328 );
not \U$11493 ( \12330 , \12038_nG2e11 );
or \U$11494 ( \12331 , \11839 , \12330 );
not \U$11495 ( \12332 , \12089_nG2d11 );
or \U$11496 ( \12333 , \12332 , \11806 );
or \U$11497 ( \12334 , \11803 , \12330 );
or \U$11498 ( \12335 , \11800 , \12089_nG2d11 );
nand \U$11499 ( \12336 , \12335 , \11836 );
nand \U$11500 ( \12337 , \12334 , \12336 );
nand \U$11501 ( \12338 , \12331 , \12333 , \12337 );
xor \U$11502 ( \12339 , \12329 , \12338 );
xor \U$11503 ( \12340 , \12327 , \12339 );
and \U$11504 ( \12341 , \12267 , \12276 );
or \U$11505 ( \12342 , \12295 , \12298 );
nand \U$11506 ( \12343 , \12342 , \12293 );
xor \U$11507 ( \12344 , \12341 , \12343 );
and \U$11508 ( \12345 , \12340 , \12344 );
xor \U$11509 ( \12346 , \12304 , \12345 );
xnor \U$11510 ( \12347 , \12090 , \12097 );
not \U$11511 ( \12348 , \12347 );
xor \U$11512 ( \12349 , \12062 , \12051 );
not \U$11513 ( \12350 , \12349 );
and \U$11514 ( \12351 , \12348 , \12350 );
and \U$11515 ( \12352 , \12347 , \12349 );
nor \U$11516 ( \12353 , \12351 , \12352 );
and \U$11517 ( \12354 , \12322 , \12229 );
and \U$11518 ( \12355 , \12329 , \12338 );
nor \U$11519 ( \12356 , \12354 , \12355 , \12320 );
or \U$11520 ( \12357 , \12353 , \12356 );
nand \U$11521 ( \12358 , \12356 , \12353 );
nand \U$11522 ( \12359 , \12357 , \12358 );
and \U$11523 ( \12360 , \12346 , \12359 );
and \U$11524 ( \12361 , \12304 , \12345 );
or \U$11525 ( \12362 , \12360 , \12361 );
not \U$11526 ( \12363 , \12349 );
nor \U$11527 ( \12364 , \12363 , \12347 );
xor \U$11528 ( \12365 , \12362 , \12364 );
and \U$11529 ( \12366 , \12327 , \12339 );
and \U$11530 ( \12367 , \12341 , \12343 );
and \U$11531 ( \12368 , \12366 , \12367 );
xor \U$11532 ( \12369 , \12368 , \12358 );
not \U$11533 ( \12370 , \12099 );
not \U$11534 ( \12371 , \12043 );
or \U$11535 ( \12372 , \12370 , \12371 );
or \U$11536 ( \12373 , \12043 , \12099 );
nand \U$11537 ( \12374 , \12372 , \12373 );
xor \U$11538 ( \12375 , \12369 , \12374 );
and \U$11539 ( \12376 , \12365 , \12375 );
and \U$11540 ( \12377 , \12362 , \12364 );
or \U$11541 ( \12378 , \12376 , \12377 );
not \U$11542 ( \12379 , \12039 );
nand \U$11543 ( \12380 , \12379 , \12011 );
not \U$11544 ( \12381 , \12100 );
not \U$11545 ( \12382 , \12103 );
and \U$11546 ( \12383 , \12381 , \12382 );
and \U$11547 ( \12384 , \12100 , \12103 );
nor \U$11548 ( \12385 , \12383 , \12384 );
nand \U$11549 ( \12386 , \12380 , \12385 );
not \U$11550 ( \12387 , \12386 );
nor \U$11551 ( \12388 , \12385 , \12380 );
nor \U$11552 ( \12389 , \12387 , \12388 );
not \U$11553 ( \12390 , \12389 );
xor \U$11554 ( \12391 , \12368 , \12358 );
and \U$11555 ( \12392 , \12391 , \12374 );
and \U$11556 ( \12393 , \12368 , \12358 );
or \U$11557 ( \12394 , \12392 , \12393 );
not \U$11558 ( \12395 , \12394 );
and \U$11559 ( \12396 , \12390 , \12395 );
and \U$11560 ( \12397 , \12389 , \12394 );
nor \U$11561 ( \12398 , \12396 , \12397 );
xor \U$11562 ( \12399 , \12378 , \12398 );
xor \U$11563 ( \12400 , \12362 , \12364 );
xor \U$11564 ( \12401 , \12400 , \12375 );
xor \U$11565 ( \12402 , \12340 , \12344 );
not \U$11566 ( \12403 , \12255 );
not \U$11567 ( \12404 , \12224 );
or \U$11568 ( \12405 , \12403 , \12404 );
or \U$11569 ( \12406 , \12224 , \12255 );
nand \U$11570 ( \12407 , \12405 , \12406 );
xor \U$11571 ( \12408 , \12253 , \12256 );
nor \U$11572 ( \12409 , \12407 , \12408 );
not \U$11573 ( \12410 , \12409 );
not \U$11574 ( \12411 , \12258 );
nor \U$11575 ( \12412 , \12410 , \12411 );
not \U$11576 ( \12413 , \12412 );
or \U$11577 ( \12414 , \12413 , \11833 );
or \U$11578 ( \12415 , \12410 , \11833 );
nand \U$11579 ( \12416 , \12415 , \12411 );
nand \U$11580 ( \12417 , \12414 , \12416 );
or \U$11581 ( \12418 , \12263 , \11901 );
not \U$11582 ( \12419 , \12234 );
or \U$11583 ( \12420 , \11788 , \12419 );
or \U$11584 ( \12421 , \12236 , \11901 );
or \U$11585 ( \12422 , \12229 , \11787_nG3124 );
nand \U$11586 ( \12423 , \12422 , \12231 );
nand \U$11587 ( \12424 , \12421 , \12423 );
nand \U$11588 ( \12425 , \12418 , \12420 , \12424 );
and \U$11589 ( \12426 , \12417 , \12425 );
and \U$11590 ( \12427 , \12142_nG2c0d , \11894 );
and \U$11591 ( \12428 , \11936 , \12089_nG2d11 );
nand \U$11592 ( \12429 , \12142_nG2c0d , \11891 );
or \U$11593 ( \12430 , \11852 , \12089_nG2d11 );
nand \U$11594 ( \12431 , \12430 , \11940 );
and \U$11595 ( \12432 , \12429 , \12431 );
nor \U$11596 ( \12433 , \12427 , \12428 , \12432 );
nand \U$11597 ( \12434 , \11972_nG2efb , \12054 );
or \U$11598 ( \12435 , \11985 , \12038_nG2e11 );
nand \U$11599 ( \12436 , \12435 , \12060 );
and \U$11600 ( \12437 , \12434 , \12436 );
and \U$11601 ( \12438 , \12056 , \12038_nG2e11 );
and \U$11602 ( \12439 , \11972_nG2efb , \12247 );
nor \U$11603 ( \12440 , \12437 , \12438 , \12439 );
xor \U$11604 ( \12441 , \12433 , \12440 );
and \U$11605 ( \12442 , \12169_nG2b05 , \11944 );
and \U$11606 ( \12443 , \11946 , \12210_nG2a23 );
nand \U$11607 ( \12444 , \12169_nG2b05 , \11804 );
or \U$11608 ( \12445 , \11800 , \12210_nG2a23 );
nand \U$11609 ( \12446 , \12445 , \11836 );
and \U$11610 ( \12447 , \12444 , \12446 );
nor \U$11611 ( \12448 , \12442 , \12443 , \12447 );
and \U$11612 ( \12449 , \12441 , \12448 );
and \U$11613 ( \12450 , \12433 , \12440 );
or \U$11614 ( \12451 , \12449 , \12450 );
not \U$11615 ( \12452 , \12451 );
and \U$11616 ( \12453 , \12426 , \12452 );
not \U$11617 ( \12454 , \12258 );
not \U$11618 ( \12455 , \12260 );
nand \U$11619 ( \12456 , \12455 , \12250 );
not \U$11620 ( \12457 , \12456 );
or \U$11621 ( \12458 , \12454 , \12457 );
or \U$11622 ( \12459 , \12456 , \12258 );
nand \U$11623 ( \12460 , \12458 , \12459 );
not \U$11624 ( \12461 , \12211 );
nor \U$11625 ( \12462 , \12183 , \12214 );
not \U$11626 ( \12463 , \12462 );
or \U$11627 ( \12464 , \12461 , \12463 );
or \U$11628 ( \12465 , \12462 , \12211 );
nand \U$11629 ( \12466 , \12464 , \12465 );
and \U$11630 ( \12467 , \12460 , \12466 );
and \U$11631 ( \12468 , \12453 , \12467 );
xor \U$11632 ( \12469 , \12402 , \12468 );
xnor \U$11633 ( \12470 , \12261 , \12215 );
not \U$11634 ( \12471 , \12302 );
not \U$11635 ( \12472 , \12277 );
and \U$11636 ( \12473 , \12471 , \12472 );
and \U$11637 ( \12474 , \12302 , \12277 );
nor \U$11638 ( \12475 , \12473 , \12474 );
nand \U$11639 ( \12476 , \12470 , \12475 );
and \U$11640 ( \12477 , \12469 , \12476 );
and \U$11641 ( \12478 , \12402 , \12468 );
or \U$11642 ( \12479 , \12477 , \12478 );
xor \U$11643 ( \12480 , \12366 , \12367 );
xor \U$11644 ( \12481 , \12479 , \12480 );
xor \U$11645 ( \12482 , \12304 , \12345 );
xor \U$11646 ( \12483 , \12482 , \12359 );
and \U$11647 ( \12484 , \12481 , \12483 );
and \U$11648 ( \12485 , \12479 , \12480 );
or \U$11649 ( \12486 , \12484 , \12485 );
xor \U$11650 ( \12487 , \12401 , \12486 );
xor \U$11651 ( \12488 , \12479 , \12480 );
xor \U$11652 ( \12489 , \12488 , \12483 );
xor \U$11653 ( \12490 , \12262 , \12303 );
xor \U$11654 ( \12491 , \12402 , \12468 );
xor \U$11655 ( \12492 , \12491 , \12476 );
and \U$11656 ( \12493 , \12490 , \12492 );
xor \U$11657 ( \12494 , \12426 , \12452 );
xor \U$11658 ( \12495 , \12460 , \12466 );
and \U$11659 ( \12496 , \12494 , \12495 );
xor \U$11660 ( \12497 , \12417 , \12425 );
xor \U$11661 ( \12498 , \12433 , \12440 );
xor \U$11662 ( \12499 , \12498 , \12448 );
not \U$11663 ( \12500 , \12499 );
and \U$11664 ( \12501 , \12497 , \12500 );
and \U$11665 ( \12502 , \12169_nG2b05 , \11894 );
and \U$11666 ( \12503 , \11936 , \12142_nG2c0d );
nand \U$11667 ( \12504 , \12169_nG2b05 , \11891 );
or \U$11668 ( \12505 , \11852 , \12142_nG2c0d );
nand \U$11669 ( \12506 , \12505 , \11940 );
and \U$11670 ( \12507 , \12504 , \12506 );
nor \U$11671 ( \12508 , \12502 , \12503 , \12507 );
nand \U$11672 ( \12509 , \12038_nG2e11 , \12054 );
or \U$11673 ( \12510 , \11985 , \12089_nG2d11 );
nand \U$11674 ( \12511 , \12510 , \12060 );
and \U$11675 ( \12512 , \12509 , \12511 );
and \U$11676 ( \12513 , \12056 , \12089_nG2d11 );
and \U$11677 ( \12514 , \12038_nG2e11 , \12247 );
nor \U$11678 ( \12515 , \12512 , \12513 , \12514 );
xor \U$11679 ( \12516 , \12508 , \12515 );
and \U$11680 ( \12517 , \12210_nG2a23 , \11944 );
and \U$11681 ( \12518 , \11760 , RIb5557d8_384);
and \U$11682 ( \12519 , RIb555df0_397, \7936 );
nor \U$11683 ( \12520 , \12518 , \12519 );
and \U$11684 ( \12521 , \7938 , RIb555d78_396);
and \U$11685 ( \12522 , RIb555c10_393, \7955 );
nor \U$11686 ( \12523 , \12521 , \12522 );
and \U$11687 ( \12524 , \7950 , RIb5558c8_386);
and \U$11688 ( \12525 , RIb555940_387, \7900 );
nor \U$11689 ( \12526 , \12524 , \12525 );
and \U$11690 ( \12527 , \7917 , RIb555850_385);
and \U$11691 ( \12528 , \7906 , RIb555a30_389);
and \U$11692 ( \12529 , RIb5559b8_388, \7953 );
nor \U$11693 ( \12530 , \12528 , \12529 );
and \U$11694 ( \12531 , \7943 , RIb555c88_394);
and \U$11695 ( \12532 , RIb555d00_395, \7945 );
nor \U$11696 ( \12533 , \12531 , \12532 );
and \U$11697 ( \12534 , \7948 , RIb555e68_398);
and \U$11698 ( \12535 , RIb555b98_392, \7926 );
nor \U$11699 ( \12536 , \12534 , \12535 );
and \U$11700 ( \12537 , \7914 , RIb555aa8_390);
and \U$11701 ( \12538 , RIb555b20_391, \7910 );
nor \U$11702 ( \12539 , \12537 , \12538 );
nand \U$11703 ( \12540 , \12530 , \12533 , \12536 , \12539 );
nor \U$11704 ( \12541 , \12527 , \12540 );
nand \U$11705 ( \12542 , \12520 , \12523 , \12526 , \12541 );
_DC g292b ( \12543_nG292b , \12542 , \11786 );
and \U$11706 ( \12544 , \11946 , \12543_nG292b );
nand \U$11707 ( \12545 , \12210_nG2a23 , \11804 );
or \U$11708 ( \12546 , \11800 , \12543_nG292b );
nand \U$11709 ( \12547 , \12546 , \11836 );
and \U$11710 ( \12548 , \12545 , \12547 );
nor \U$11711 ( \12549 , \12517 , \12544 , \12548 );
and \U$11712 ( \12550 , \12516 , \12549 );
and \U$11713 ( \12551 , \12508 , \12515 );
or \U$11714 ( \12552 , \12550 , \12551 );
and \U$11715 ( \12553 , \12258 , \12408 );
and \U$11716 ( \12554 , \11832_nG323c , \12553 );
or \U$11717 ( \12555 , \12258 , \11832_nG323c );
or \U$11718 ( \12556 , \12258 , \12408 );
nand \U$11719 ( \12557 , \12555 , \12556 );
nand \U$11720 ( \12558 , \11787_nG3124 , \12409 );
and \U$11721 ( \12559 , \12557 , \12558 );
and \U$11722 ( \12560 , \11787_nG3124 , \12412 );
nor \U$11723 ( \12561 , \12554 , \12559 , \12560 );
xor \U$11724 ( \12562 , RIb55bca0_599, \11689_nG2277 );
xor \U$11725 ( \12563 , \12562 , \11720 );
not \U$11726 ( \12564 , \12563 );
xor \U$11727 ( \12565 , \8302 , \11660_nG23e0 );
xor \U$11728 ( \12566 , \12565 , \11723 );
not \U$11729 ( \12567 , \12566 );
and \U$11730 ( \12568 , \12564 , \12567 );
or \U$11731 ( \12569 , \12252 , \12568 );
not \U$11732 ( \12570 , \12569 );
xor \U$11733 ( \12571 , \12561 , \12570 );
nand \U$11734 ( \12572 , \11972_nG2efb , \12226 );
or \U$11735 ( \12573 , \12229 , \11879_nG301d );
nand \U$11736 ( \12574 , \12573 , \12231 );
and \U$11737 ( \12575 , \12572 , \12574 );
and \U$11738 ( \12576 , \12234 , \11879_nG301d );
and \U$11739 ( \12577 , \11972_nG2efb , \12238 );
nor \U$11740 ( \12578 , \12575 , \12576 , \12577 );
and \U$11741 ( \12579 , \12571 , \12578 );
and \U$11742 ( \12580 , \12561 , \12570 );
or \U$11743 ( \12581 , \12579 , \12580 );
nor \U$11744 ( \12582 , \12552 , \12581 );
and \U$11745 ( \12583 , \12501 , \12582 );
xor \U$11746 ( \12584 , \12496 , \12583 );
or \U$11747 ( \12585 , \12475 , \12470 );
nand \U$11748 ( \12586 , \12585 , \12476 );
and \U$11749 ( \12587 , \12584 , \12586 );
and \U$11750 ( \12588 , \12496 , \12583 );
or \U$11751 ( \12589 , \12587 , \12588 );
xor \U$11752 ( \12590 , \12402 , \12468 );
xor \U$11753 ( \12591 , \12590 , \12476 );
and \U$11754 ( \12592 , \12589 , \12591 );
and \U$11755 ( \12593 , \12490 , \12589 );
or \U$11756 ( \12594 , \12493 , \12592 , \12593 );
xor \U$11757 ( \12595 , \12489 , \12594 );
nand \U$11758 ( \12596 , \12543_nG292b , \11757 );
not \U$11759 ( \12597 , \12596 );
xor \U$11760 ( \12598 , \12497 , \12500 );
not \U$11761 ( \12599 , \12598 );
or \U$11762 ( \12600 , \12597 , \12599 );
xnor \U$11763 ( \12601 , \12581 , \12552 );
nand \U$11764 ( \12602 , \12600 , \12601 );
or \U$11765 ( \12603 , \12252 , \12566 );
nand \U$11766 ( \12604 , \12566 , \12252 );
nand \U$11767 ( \12605 , \12603 , \12604 );
xor \U$11768 ( \12606 , \12564 , \12567 );
nor \U$11769 ( \12607 , \12605 , \12606 );
not \U$11770 ( \12608 , \12607 );
nor \U$11771 ( \12609 , \12608 , \12570 );
not \U$11772 ( \12610 , \12609 );
or \U$11773 ( \12611 , \12610 , \11833 );
or \U$11774 ( \12612 , \12608 , \11833 );
nand \U$11775 ( \12613 , \12612 , \12570 );
nand \U$11776 ( \12614 , \12611 , \12613 );
not \U$11777 ( \12615 , \12614 );
and \U$11778 ( \12616 , \11787_nG3124 , \12553 );
or \U$11779 ( \12617 , \12258 , \11787_nG3124 );
nand \U$11780 ( \12618 , \12617 , \12556 );
nand \U$11781 ( \12619 , \11879_nG301d , \12409 );
and \U$11782 ( \12620 , \12618 , \12619 );
and \U$11783 ( \12621 , \11879_nG301d , \12412 );
nor \U$11784 ( \12622 , \12616 , \12620 , \12621 );
nor \U$11785 ( \12623 , \12615 , \12622 );
not \U$11786 ( \12624 , \12623 );
nand \U$11787 ( \12625 , \12089_nG2d11 , \12054 );
or \U$11788 ( \12626 , \11985 , \12142_nG2c0d );
nand \U$11789 ( \12627 , \12626 , \12060 );
and \U$11790 ( \12628 , \12625 , \12627 );
and \U$11791 ( \12629 , \12056 , \12142_nG2c0d );
and \U$11792 ( \12630 , \12089_nG2d11 , \12247 );
nor \U$11793 ( \12631 , \12628 , \12629 , \12630 );
nand \U$11794 ( \12632 , \12038_nG2e11 , \12226 );
or \U$11795 ( \12633 , \12229 , \11972_nG2efb );
nand \U$11796 ( \12634 , \12633 , \12231 );
and \U$11797 ( \12635 , \12632 , \12634 );
and \U$11798 ( \12636 , \12234 , \11972_nG2efb );
and \U$11799 ( \12637 , \12038_nG2e11 , \12238 );
nor \U$11800 ( \12638 , \12635 , \12636 , \12637 );
xor \U$11801 ( \12639 , \12631 , \12638 );
and \U$11802 ( \12640 , \12210_nG2a23 , \11894 );
and \U$11803 ( \12641 , \11936 , \12169_nG2b05 );
nand \U$11804 ( \12642 , \12210_nG2a23 , \11891 );
or \U$11805 ( \12643 , \11852 , \12169_nG2b05 );
nand \U$11806 ( \12644 , \12643 , \11940 );
and \U$11807 ( \12645 , \12642 , \12644 );
nor \U$11808 ( \12646 , \12640 , \12641 , \12645 );
and \U$11809 ( \12647 , \12639 , \12646 );
and \U$11810 ( \12648 , \12631 , \12638 );
or \U$11811 ( \12649 , \12647 , \12648 );
nor \U$11812 ( \12650 , \12624 , \12649 );
xor \U$11813 ( \12651 , \12508 , \12515 );
xor \U$11814 ( \12652 , \12651 , \12549 );
xor \U$11815 ( \12653 , \12561 , \12570 );
xor \U$11816 ( \12654 , \12653 , \12578 );
nor \U$11817 ( \12655 , \12652 , \12654 );
not \U$11818 ( \12656 , \12655 );
and \U$11819 ( \12657 , \11760 , RIb556fc0_435);
and \U$11820 ( \12658 , RIb5575d8_448, \7936 );
nor \U$11821 ( \12659 , \12657 , \12658 );
and \U$11822 ( \12660 , \7938 , RIb557560_447);
and \U$11823 ( \12661 , RIb5573f8_444, \7955 );
nor \U$11824 ( \12662 , \12660 , \12661 );
and \U$11825 ( \12663 , \7950 , RIb5570b0_437);
and \U$11826 ( \12664 , RIb557128_438, \7900 );
nor \U$11827 ( \12665 , \12663 , \12664 );
and \U$11828 ( \12666 , \7917 , RIb557038_436);
and \U$11829 ( \12667 , \7943 , RIb557470_445);
and \U$11830 ( \12668 , RIb557380_443, \7926 );
nor \U$11831 ( \12669 , \12667 , \12668 );
and \U$11832 ( \12670 , \7914 , RIb557290_441);
and \U$11833 ( \12671 , RIb557308_442, \7910 );
nor \U$11834 ( \12672 , \12670 , \12671 );
and \U$11835 ( \12673 , \7948 , RIb557650_449);
and \U$11836 ( \12674 , RIb5574e8_446, \7945 );
nor \U$11837 ( \12675 , \12673 , \12674 );
and \U$11838 ( \12676 , \7906 , RIb557218_440);
and \U$11839 ( \12677 , RIb5571a0_439, \7953 );
nor \U$11840 ( \12678 , \12676 , \12677 );
nand \U$11841 ( \12679 , \12669 , \12672 , \12675 , \12678 );
nor \U$11842 ( \12680 , \12666 , \12679 );
nand \U$11843 ( \12681 , \12659 , \12662 , \12665 , \12680 );
_DC g2848 ( \12682_nG2848 , \12681 , \11786 );
nand \U$11844 ( \12683 , \12682_nG2848 , \11757 );
nand \U$11845 ( \12684 , \12656 , \12683 );
and \U$11846 ( \12685 , \12650 , \12684 );
xor \U$11847 ( \12686 , \12602 , \12685 );
xor \U$11848 ( \12687 , \12494 , \12495 );
and \U$11849 ( \12688 , \12686 , \12687 );
and \U$11850 ( \12689 , \12602 , \12685 );
or \U$11851 ( \12690 , \12688 , \12689 );
xor \U$11852 ( \12691 , \12453 , \12467 );
xor \U$11853 ( \12692 , \12690 , \12691 );
xor \U$11854 ( \12693 , \12496 , \12583 );
xor \U$11855 ( \12694 , \12693 , \12586 );
and \U$11856 ( \12695 , \12692 , \12694 );
and \U$11857 ( \12696 , \12690 , \12691 );
or \U$11858 ( \12697 , \12695 , \12696 );
xor \U$11859 ( \12698 , \12402 , \12468 );
xor \U$11860 ( \12699 , \12698 , \12476 );
xor \U$11861 ( \12700 , \12490 , \12589 );
xor \U$11862 ( \12701 , \12699 , \12700 );
xor \U$11863 ( \12702 , \12697 , \12701 );
xor \U$11864 ( \12703 , \12690 , \12691 );
xor \U$11865 ( \12704 , \12703 , \12694 );
not \U$11866 ( \12705 , \12596 );
nor \U$11867 ( \12706 , \12705 , \12582 );
not \U$11868 ( \12707 , \12706 );
not \U$11869 ( \12708 , \12501 );
or \U$11870 ( \12709 , \12707 , \12708 );
or \U$11871 ( \12710 , \12501 , \12706 );
nand \U$11872 ( \12711 , \12709 , \12710 );
xor \U$11873 ( \12712 , \12602 , \12685 );
xor \U$11874 ( \12713 , \12712 , \12687 );
and \U$11875 ( \12714 , \12711 , \12713 );
or \U$11876 ( \12715 , \12649 , \12623 );
and \U$11877 ( \12716 , \11760 , RIb5567c8_418);
and \U$11878 ( \12717 , RIb556de0_431, \7936 );
nor \U$11879 ( \12718 , \12716 , \12717 );
and \U$11880 ( \12719 , \7938 , RIb556d68_430);
and \U$11881 ( \12720 , RIb556c00_427, \7955 );
nor \U$11882 ( \12721 , \12719 , \12720 );
and \U$11883 ( \12722 , \7950 , RIb5568b8_420);
and \U$11884 ( \12723 , RIb556930_421, \7900 );
nor \U$11885 ( \12724 , \12722 , \12723 );
and \U$11886 ( \12725 , \7917 , RIb556840_419);
and \U$11887 ( \12726 , \7943 , RIb556c78_428);
and \U$11888 ( \12727 , RIb556b88_426, \7926 );
nor \U$11889 ( \12728 , \12726 , \12727 );
and \U$11890 ( \12729 , \7914 , RIb556a98_424);
and \U$11891 ( \12730 , RIb556b10_425, \7910 );
nor \U$11892 ( \12731 , \12729 , \12730 );
and \U$11893 ( \12732 , \7948 , RIb556e58_432);
and \U$11894 ( \12733 , RIb556cf0_429, \7945 );
nor \U$11895 ( \12734 , \12732 , \12733 );
and \U$11896 ( \12735 , \7906 , RIb556a20_423);
and \U$11897 ( \12736 , RIb5569a8_422, \7953 );
nor \U$11898 ( \12737 , \12735 , \12736 );
nand \U$11899 ( \12738 , \12728 , \12731 , \12734 , \12737 );
nor \U$11900 ( \12739 , \12725 , \12738 );
nand \U$11901 ( \12740 , \12718 , \12721 , \12724 , \12739 );
_DC g2776 ( \12741_nG2776 , \12740 , \11786 );
nand \U$11902 ( \12742 , \12741_nG2776 , \11757 );
and \U$11903 ( \12743 , \12543_nG292b , \11944 );
and \U$11904 ( \12744 , \11946 , \12682_nG2848 );
nand \U$11905 ( \12745 , \12543_nG292b , \11804 );
or \U$11906 ( \12746 , \11800 , \12682_nG2848 );
nand \U$11907 ( \12747 , \12746 , \11836 );
and \U$11908 ( \12748 , \12745 , \12747 );
nor \U$11909 ( \12749 , \12743 , \12744 , \12748 );
or \U$11910 ( \12750 , \12742 , \12749 );
nand \U$11911 ( \12751 , \12623 , \12649 );
nand \U$11912 ( \12752 , \12715 , \12750 , \12751 );
not \U$11913 ( \12753 , \12752 );
and \U$11914 ( \12754 , \12652 , \12654 );
nor \U$11915 ( \12755 , \12754 , \12655 );
not \U$11916 ( \12756 , \12755 );
not \U$11917 ( \12757 , \12683 );
and \U$11918 ( \12758 , \12756 , \12757 );
and \U$11919 ( \12759 , \12755 , \12683 );
nor \U$11920 ( \12760 , \12758 , \12759 );
nor \U$11921 ( \12761 , \12753 , \12760 );
not \U$11922 ( \12762 , \12543_nG292b );
or \U$11923 ( \12763 , \11895 , \12762 );
and \U$11924 ( \12764 , \11936 , \12210_nG2a23 );
nand \U$11925 ( \12765 , \12543_nG292b , \11891 );
or \U$11926 ( \12766 , \11852 , \12210_nG2a23 );
nand \U$11927 ( \12767 , \12766 , \11940 );
and \U$11928 ( \12768 , \12765 , \12767 );
nor \U$11929 ( \12769 , \12764 , \12768 );
nand \U$11930 ( \12770 , \12763 , \12769 );
nand \U$11931 ( \12771 , \12089_nG2d11 , \12226 );
or \U$11932 ( \12772 , \12229 , \12038_nG2e11 );
nand \U$11933 ( \12773 , \12772 , \12231 );
and \U$11934 ( \12774 , \12771 , \12773 );
and \U$11935 ( \12775 , \12234 , \12038_nG2e11 );
and \U$11936 ( \12776 , \12089_nG2d11 , \12238 );
nor \U$11937 ( \12777 , \12774 , \12775 , \12776 );
nand \U$11938 ( \12778 , \12142_nG2c0d , \12054 );
or \U$11939 ( \12779 , \11985 , \12169_nG2b05 );
nand \U$11940 ( \12780 , \12779 , \12060 );
and \U$11941 ( \12781 , \12778 , \12780 );
and \U$11942 ( \12782 , \12056 , \12169_nG2b05 );
and \U$11943 ( \12783 , \12142_nG2c0d , \12247 );
nor \U$11944 ( \12784 , \12781 , \12782 , \12783 );
nand \U$11945 ( \12785 , \12777 , \12784 );
and \U$11946 ( \12786 , \12770 , \12785 );
nor \U$11947 ( \12787 , \12784 , \12777 );
nor \U$11948 ( \12788 , \12786 , \12787 );
nand \U$11949 ( \12789 , \11787_nG3124 , \12607 );
or \U$11950 ( \12790 , \12569 , \11832_nG323c );
or \U$11951 ( \12791 , \12569 , \12606 );
nand \U$11952 ( \12792 , \12790 , \12791 );
and \U$11953 ( \12793 , \12789 , \12792 );
and \U$11954 ( \12794 , \12569 , \12606 );
and \U$11955 ( \12795 , \12794 , \11832_nG323c );
and \U$11956 ( \12796 , \11787_nG3124 , \12609 );
nor \U$11957 ( \12797 , \12793 , \12795 , \12796 );
xor \U$11958 ( \12798 , \12797 , \12564 );
and \U$11959 ( \12799 , \11879_nG301d , \12553 );
or \U$11960 ( \12800 , \12258 , \11879_nG301d );
nand \U$11961 ( \12801 , \12800 , \12556 );
nand \U$11962 ( \12802 , \11972_nG2efb , \12409 );
and \U$11963 ( \12803 , \12801 , \12802 );
and \U$11964 ( \12804 , \11972_nG2efb , \12412 );
nor \U$11965 ( \12805 , \12799 , \12803 , \12804 );
and \U$11966 ( \12806 , \12798 , \12805 );
and \U$11967 ( \12807 , \12797 , \12564 );
or \U$11968 ( \12808 , \12806 , \12807 );
nor \U$11969 ( \12809 , \12788 , \12808 );
not \U$11970 ( \12810 , \12809 );
not \U$11971 ( \12811 , \12622 );
not \U$11972 ( \12812 , \12614 );
and \U$11973 ( \12813 , \12811 , \12812 );
and \U$11974 ( \12814 , \12622 , \12614 );
nor \U$11975 ( \12815 , \12813 , \12814 );
xor \U$11976 ( \12816 , \12631 , \12638 );
xor \U$11977 ( \12817 , \12816 , \12646 );
and \U$11978 ( \12818 , \12815 , \12817 );
xnor \U$11979 ( \12819 , \12742 , \12749 );
xor \U$11980 ( \12820 , \12631 , \12638 );
xor \U$11981 ( \12821 , \12820 , \12646 );
and \U$11982 ( \12822 , \12819 , \12821 );
and \U$11983 ( \12823 , \12815 , \12819 );
or \U$11984 ( \12824 , \12818 , \12822 , \12823 );
nor \U$11985 ( \12825 , \12810 , \12824 );
xor \U$11986 ( \12826 , \12761 , \12825 );
not \U$11987 ( \12827 , \12596 );
xor \U$11988 ( \12828 , \12601 , \12598 );
not \U$11989 ( \12829 , \12828 );
or \U$11990 ( \12830 , \12827 , \12829 );
or \U$11991 ( \12831 , \12828 , \12596 );
nand \U$11992 ( \12832 , \12830 , \12831 );
and \U$11993 ( \12833 , \12826 , \12832 );
and \U$11994 ( \12834 , \12761 , \12825 );
or \U$11995 ( \12835 , \12833 , \12834 );
xor \U$11996 ( \12836 , \12602 , \12685 );
xor \U$11997 ( \12837 , \12836 , \12687 );
and \U$11998 ( \12838 , \12835 , \12837 );
and \U$11999 ( \12839 , \12711 , \12835 );
or \U$12000 ( \12840 , \12714 , \12838 , \12839 );
xor \U$12001 ( \12841 , \12704 , \12840 );
xor \U$12002 ( \12842 , \12602 , \12685 );
xor \U$12003 ( \12843 , \12842 , \12687 );
xor \U$12004 ( \12844 , \12711 , \12835 );
xor \U$12005 ( \12845 , \12843 , \12844 );
xor \U$12006 ( \12846 , \12761 , \12825 );
xor \U$12007 ( \12847 , \12846 , \12832 );
xor \U$12008 ( \12848 , \12650 , \12684 );
nor \U$12009 ( \12849 , \12847 , \12848 );
nand \U$12010 ( \12850 , \12142_nG2c0d , \12226 );
or \U$12011 ( \12851 , \12229 , \12089_nG2d11 );
nand \U$12012 ( \12852 , \12851 , \12231 );
and \U$12013 ( \12853 , \12850 , \12852 );
and \U$12014 ( \12854 , \12234 , \12089_nG2d11 );
and \U$12015 ( \12855 , \12142_nG2c0d , \12238 );
nor \U$12016 ( \12856 , \12853 , \12854 , \12855 );
and \U$12017 ( \12857 , \11972_nG2efb , \12553 );
or \U$12018 ( \12858 , \12258 , \11972_nG2efb );
nand \U$12019 ( \12859 , \12858 , \12556 );
nand \U$12020 ( \12860 , \12038_nG2e11 , \12409 );
and \U$12021 ( \12861 , \12859 , \12860 );
and \U$12022 ( \12862 , \12038_nG2e11 , \12412 );
nor \U$12023 ( \12863 , \12857 , \12861 , \12862 );
xor \U$12024 ( \12864 , \12856 , \12863 );
nand \U$12025 ( \12865 , \12169_nG2b05 , \12054 );
or \U$12026 ( \12866 , \11985 , \12210_nG2a23 );
nand \U$12027 ( \12867 , \12866 , \12060 );
and \U$12028 ( \12868 , \12865 , \12867 );
and \U$12029 ( \12869 , \12056 , \12210_nG2a23 );
and \U$12030 ( \12870 , \12169_nG2b05 , \12247 );
nor \U$12031 ( \12871 , \12868 , \12869 , \12870 );
and \U$12032 ( \12872 , \12864 , \12871 );
and \U$12033 ( \12873 , \12856 , \12863 );
or \U$12034 ( \12874 , \12872 , \12873 );
nand \U$12035 ( \12875 , \11879_nG301d , \12607 );
or \U$12036 ( \12876 , \12569 , \11787_nG3124 );
nand \U$12037 ( \12877 , \12876 , \12791 );
and \U$12038 ( \12878 , \12875 , \12877 );
and \U$12039 ( \12879 , \12794 , \11787_nG3124 );
and \U$12040 ( \12880 , \11879_nG301d , \12609 );
nor \U$12041 ( \12881 , \12878 , \12879 , \12880 );
not \U$12042 ( \12882 , \12881 );
or \U$12043 ( \12883 , \12563 , \11832_nG323c );
or \U$12044 ( \12884 , \8395 , \11718_nG2275 );
nand \U$12045 ( \12885 , \12884 , \11719 );
nor \U$12046 ( \12886 , \12563 , \12885 );
not \U$12047 ( \12887 , \12886 );
nand \U$12048 ( \12888 , \12564 , \12887 );
nand \U$12049 ( \12889 , \12883 , \12888 );
nand \U$12050 ( \12890 , \12882 , \12889 );
xor \U$12051 ( \12891 , \12874 , \12890 );
and \U$12052 ( \12892 , \12741_nG2776 , \11944 );
and \U$12053 ( \12893 , \11760 , RIb557fb0_469);
and \U$12054 ( \12894 , RIb5585c8_482, \7936 );
nor \U$12055 ( \12895 , \12893 , \12894 );
and \U$12056 ( \12896 , \7938 , RIb558550_481);
and \U$12057 ( \12897 , RIb5583e8_478, \7955 );
nor \U$12058 ( \12898 , \12896 , \12897 );
and \U$12059 ( \12899 , \7950 , RIb5580a0_471);
and \U$12060 ( \12900 , RIb558118_472, \7900 );
nor \U$12061 ( \12901 , \12899 , \12900 );
and \U$12062 ( \12902 , \7917 , RIb558028_470);
and \U$12063 ( \12903 , \7943 , RIb558460_479);
and \U$12064 ( \12904 , RIb558370_477, \7926 );
nor \U$12065 ( \12905 , \12903 , \12904 );
and \U$12066 ( \12906 , \7914 , RIb558280_475);
and \U$12067 ( \12907 , RIb5582f8_476, \7910 );
nor \U$12068 ( \12908 , \12906 , \12907 );
and \U$12069 ( \12909 , \7948 , RIb558640_483);
and \U$12070 ( \12910 , RIb5584d8_480, \7945 );
nor \U$12071 ( \12911 , \12909 , \12910 );
and \U$12072 ( \12912 , \7906 , RIb558208_474);
and \U$12073 ( \12913 , RIb558190_473, \7953 );
nor \U$12074 ( \12914 , \12912 , \12913 );
nand \U$12075 ( \12915 , \12905 , \12908 , \12911 , \12914 );
nor \U$12076 ( \12916 , \12902 , \12915 );
nand \U$12077 ( \12917 , \12895 , \12898 , \12901 , \12916 );
_DC g26c6 ( \12918_nG26c6 , \12917 , \11786 );
and \U$12078 ( \12919 , \11946 , \12918_nG26c6 );
nand \U$12079 ( \12920 , \12741_nG2776 , \11804 );
or \U$12080 ( \12921 , \11800 , \12918_nG26c6 );
nand \U$12081 ( \12922 , \12921 , \11836 );
and \U$12082 ( \12923 , \12920 , \12922 );
nor \U$12083 ( \12924 , \12892 , \12919 , \12923 );
and \U$12084 ( \12925 , \12682_nG2848 , \11894 );
and \U$12085 ( \12926 , \11936 , \12543_nG292b );
nand \U$12086 ( \12927 , \12682_nG2848 , \11891 );
or \U$12087 ( \12928 , \11852 , \12543_nG292b );
nand \U$12088 ( \12929 , \12928 , \11940 );
and \U$12089 ( \12930 , \12927 , \12929 );
nor \U$12090 ( \12931 , \12925 , \12926 , \12930 );
and \U$12091 ( \12932 , \12924 , \12931 );
not \U$12092 ( \12933 , \12932 );
and \U$12093 ( \12934 , \11760 , RIb5577b8_452);
and \U$12094 ( \12935 , RIb557dd0_465, \7936 );
nor \U$12095 ( \12936 , \12934 , \12935 );
and \U$12096 ( \12937 , \7938 , RIb557d58_464);
and \U$12097 ( \12938 , RIb557bf0_461, \7955 );
nor \U$12098 ( \12939 , \12937 , \12938 );
and \U$12099 ( \12940 , \7950 , RIb5578a8_454);
and \U$12100 ( \12941 , RIb557920_455, \7900 );
nor \U$12101 ( \12942 , \12940 , \12941 );
and \U$12102 ( \12943 , \7917 , RIb557830_453);
and \U$12103 ( \12944 , \7906 , RIb557a10_457);
and \U$12104 ( \12945 , RIb557998_456, \7953 );
nor \U$12105 ( \12946 , \12944 , \12945 );
and \U$12106 ( \12947 , \7914 , RIb557a88_458);
and \U$12107 ( \12948 , RIb557b00_459, \7910 );
nor \U$12108 ( \12949 , \12947 , \12948 );
and \U$12109 ( \12950 , \7948 , RIb557e48_466);
and \U$12110 ( \12951 , RIb557b78_460, \7926 );
nor \U$12111 ( \12952 , \12950 , \12951 );
and \U$12112 ( \12953 , \7943 , RIb557c68_462);
and \U$12113 ( \12954 , RIb557ce0_463, \7945 );
nor \U$12114 ( \12955 , \12953 , \12954 );
nand \U$12115 ( \12956 , \12946 , \12949 , \12952 , \12955 );
nor \U$12116 ( \12957 , \12943 , \12956 );
nand \U$12117 ( \12958 , \12936 , \12939 , \12942 , \12957 );
_DC g2600 ( \12959_nG2600 , \12958 , \11786 );
nand \U$12118 ( \12960 , \12959_nG2600 , \11757 );
not \U$12119 ( \12961 , \12960 );
and \U$12120 ( \12962 , \12933 , \12961 );
nor \U$12121 ( \12963 , \12924 , \12931 );
nor \U$12122 ( \12964 , \12962 , \12963 );
and \U$12123 ( \12965 , \12891 , \12964 );
and \U$12124 ( \12966 , \12874 , \12890 );
or \U$12125 ( \12967 , \12965 , \12966 );
nand \U$12126 ( \12968 , \12918_nG26c6 , \11757 );
and \U$12127 ( \12969 , \12682_nG2848 , \11944 );
and \U$12128 ( \12970 , \11946 , \12741_nG2776 );
nand \U$12129 ( \12971 , \12682_nG2848 , \11804 );
or \U$12130 ( \12972 , \11800 , \12741_nG2776 );
nand \U$12131 ( \12973 , \12972 , \11836 );
and \U$12132 ( \12974 , \12971 , \12973 );
nor \U$12133 ( \12975 , \12969 , \12970 , \12974 );
xnor \U$12134 ( \12976 , \12968 , \12975 );
xor \U$12135 ( \12977 , \12967 , \12976 );
xor \U$12136 ( \12978 , \12631 , \12638 );
xor \U$12137 ( \12979 , \12978 , \12646 );
xor \U$12138 ( \12980 , \12815 , \12819 );
xor \U$12139 ( \12981 , \12979 , \12980 );
and \U$12140 ( \12982 , \12977 , \12981 );
and \U$12141 ( \12983 , \12967 , \12976 );
or \U$12142 ( \12984 , \12982 , \12983 );
not \U$12143 ( \12985 , \12824 );
not \U$12144 ( \12986 , \12809 );
and \U$12145 ( \12987 , \12985 , \12986 );
and \U$12146 ( \12988 , \12824 , \12809 );
nor \U$12147 ( \12989 , \12987 , \12988 );
xor \U$12148 ( \12990 , \12984 , \12989 );
not \U$12149 ( \12991 , \12760 );
not \U$12150 ( \12992 , \12752 );
and \U$12151 ( \12993 , \12991 , \12992 );
and \U$12152 ( \12994 , \12760 , \12752 );
nor \U$12153 ( \12995 , \12993 , \12994 );
and \U$12154 ( \12996 , \12990 , \12995 );
and \U$12155 ( \12997 , \12984 , \12989 );
or \U$12156 ( \12998 , \12996 , \12997 );
or \U$12157 ( \12999 , \12849 , \12998 );
nand \U$12158 ( \13000 , \12848 , \12847 );
nand \U$12159 ( \13001 , \12999 , \13000 );
xor \U$12160 ( \13002 , \12845 , \13001 );
not \U$12161 ( \13003 , \12998 );
not \U$12162 ( \13004 , \12849 );
nand \U$12163 ( \13005 , \13004 , \13000 );
not \U$12164 ( \13006 , \13005 );
or \U$12165 ( \13007 , \13003 , \13006 );
or \U$12166 ( \13008 , \13005 , \12998 );
nand \U$12167 ( \13009 , \13007 , \13008 );
xor \U$12168 ( \13010 , \12967 , \12976 );
xor \U$12169 ( \13011 , \13010 , \12981 );
not \U$12170 ( \13012 , \13011 );
not \U$12171 ( \13013 , \12808 );
or \U$12172 ( \13014 , \12788 , \13013 );
or \U$12173 ( \13015 , \12968 , \12975 );
not \U$12174 ( \13016 , \12788 );
or \U$12175 ( \13017 , \12808 , \13016 );
nand \U$12176 ( \13018 , \13014 , \13015 , \13017 );
nand \U$12177 ( \13019 , \13012 , \13018 );
not \U$12178 ( \13020 , \12976 );
xor \U$12179 ( \13021 , \12797 , \12564 );
xor \U$12180 ( \13022 , \13021 , \12805 );
xor \U$12181 ( \13023 , \13020 , \13022 );
xor \U$12182 ( \13024 , \12874 , \12890 );
xor \U$12183 ( \13025 , \13024 , \12964 );
and \U$12184 ( \13026 , \13023 , \13025 );
and \U$12185 ( \13027 , \13020 , \13022 );
or \U$12186 ( \13028 , \13026 , \13027 );
not \U$12187 ( \13029 , \13028 );
nand \U$12188 ( \13030 , \12210_nG2a23 , \12054 );
or \U$12189 ( \13031 , \11985 , \12543_nG292b );
nand \U$12190 ( \13032 , \13031 , \12060 );
and \U$12191 ( \13033 , \13030 , \13032 );
and \U$12192 ( \13034 , \12056 , \12543_nG292b );
and \U$12193 ( \13035 , \12210_nG2a23 , \12247 );
nor \U$12194 ( \13036 , \13033 , \13034 , \13035 );
nand \U$12195 ( \13037 , \12169_nG2b05 , \12226 );
or \U$12196 ( \13038 , \12229 , \12142_nG2c0d );
nand \U$12197 ( \13039 , \13038 , \12231 );
and \U$12198 ( \13040 , \13037 , \13039 );
and \U$12199 ( \13041 , \12234 , \12142_nG2c0d );
and \U$12200 ( \13042 , \12169_nG2b05 , \12238 );
nor \U$12201 ( \13043 , \13040 , \13041 , \13042 );
xor \U$12202 ( \13044 , \13036 , \13043 );
and \U$12203 ( \13045 , \12741_nG2776 , \11894 );
and \U$12204 ( \13046 , \11936 , \12682_nG2848 );
nand \U$12205 ( \13047 , \12741_nG2776 , \11891 );
or \U$12206 ( \13048 , \11852 , \12682_nG2848 );
nand \U$12207 ( \13049 , \13048 , \11940 );
and \U$12208 ( \13050 , \13047 , \13049 );
nor \U$12209 ( \13051 , \13045 , \13046 , \13050 );
and \U$12210 ( \13052 , \13044 , \13051 );
and \U$12211 ( \13053 , \13036 , \13043 );
or \U$12212 ( \13054 , \13052 , \13053 );
nand \U$12213 ( \13055 , \11972_nG2efb , \12607 );
or \U$12214 ( \13056 , \12569 , \11879_nG301d );
nand \U$12215 ( \13057 , \13056 , \12791 );
and \U$12216 ( \13058 , \13055 , \13057 );
and \U$12217 ( \13059 , \12794 , \11879_nG301d );
and \U$12218 ( \13060 , \11972_nG2efb , \12609 );
nor \U$12219 ( \13061 , \13058 , \13059 , \13060 );
not \U$12220 ( \13062 , \13061 );
not \U$12221 ( \13063 , \12888 );
and \U$12222 ( \13064 , \11833 , \13063 );
and \U$12223 ( \13065 , \12886 , \11788 );
nand \U$12224 ( \13066 , \12885 , \12563 );
not \U$12225 ( \13067 , \13066 );
and \U$12226 ( \13068 , \11832_nG323c , \13067 );
nor \U$12227 ( \13069 , \13064 , \13065 , \13068 );
not \U$12228 ( \13070 , \13069 );
and \U$12229 ( \13071 , \13062 , \13070 );
and \U$12230 ( \13072 , \13061 , \13069 );
and \U$12231 ( \13073 , \12038_nG2e11 , \12553 );
or \U$12232 ( \13074 , \12258 , \12038_nG2e11 );
nand \U$12233 ( \13075 , \13074 , \12556 );
nand \U$12234 ( \13076 , \12089_nG2d11 , \12409 );
and \U$12235 ( \13077 , \13075 , \13076 );
and \U$12236 ( \13078 , \12089_nG2d11 , \12412 );
nor \U$12237 ( \13079 , \13073 , \13077 , \13078 );
nor \U$12238 ( \13080 , \13072 , \13079 );
nor \U$12239 ( \13081 , \13071 , \13080 );
nor \U$12240 ( \13082 , \13054 , \13081 );
not \U$12241 ( \13083 , \12787 );
nand \U$12242 ( \13084 , \13083 , \12785 );
not \U$12243 ( \13085 , \13084 );
not \U$12244 ( \13086 , \12770 );
or \U$12245 ( \13087 , \13085 , \13086 );
or \U$12246 ( \13088 , \12770 , \13084 );
nand \U$12247 ( \13089 , \13087 , \13088 );
xor \U$12248 ( \13090 , \13082 , \13089 );
not \U$12249 ( \13091 , \12960 );
nor \U$12250 ( \13092 , \12932 , \12963 );
not \U$12251 ( \13093 , \13092 );
or \U$12252 ( \13094 , \13091 , \13093 );
or \U$12253 ( \13095 , \13092 , \12960 );
nand \U$12254 ( \13096 , \13094 , \13095 );
not \U$12255 ( \13097 , \13096 );
xor \U$12256 ( \13098 , \12856 , \12863 );
xor \U$12257 ( \13099 , \13098 , \12871 );
nor \U$12258 ( \13100 , \13097 , \13099 );
and \U$12259 ( \13101 , \13090 , \13100 );
and \U$12260 ( \13102 , \13082 , \13089 );
or \U$12261 ( \13103 , \13101 , \13102 );
nor \U$12262 ( \13104 , \13029 , \13103 );
xor \U$12263 ( \13105 , \13019 , \13104 );
xor \U$12264 ( \13106 , \12984 , \12989 );
xor \U$12265 ( \13107 , \13106 , \12995 );
and \U$12266 ( \13108 , \13105 , \13107 );
and \U$12267 ( \13109 , \13019 , \13104 );
or \U$12268 ( \13110 , \13108 , \13109 );
xor \U$12269 ( \13111 , \13009 , \13110 );
not \U$12270 ( \13112 , \13081 );
or \U$12271 ( \13113 , \13054 , \13112 );
and \U$12272 ( \13114 , \11760 , RIb558fa0_503);
and \U$12273 ( \13115 , RIb5595b8_516, \7936 );
nor \U$12274 ( \13116 , \13114 , \13115 );
and \U$12275 ( \13117 , \7938 , RIb559540_515);
and \U$12276 ( \13118 , RIb5593d8_512, \7955 );
nor \U$12277 ( \13119 , \13117 , \13118 );
and \U$12278 ( \13120 , \7950 , RIb559090_505);
and \U$12279 ( \13121 , RIb559108_506, \7900 );
nor \U$12280 ( \13122 , \13120 , \13121 );
and \U$12281 ( \13123 , \7917 , RIb559018_504);
and \U$12282 ( \13124 , \7906 , RIb5591f8_508);
and \U$12283 ( \13125 , RIb559180_507, \7953 );
nor \U$12284 ( \13126 , \13124 , \13125 );
and \U$12285 ( \13127 , \7943 , RIb559450_513);
and \U$12286 ( \13128 , RIb5594c8_514, \7945 );
nor \U$12287 ( \13129 , \13127 , \13128 );
and \U$12288 ( \13130 , \7948 , RIb559630_517);
and \U$12289 ( \13131 , RIb559360_511, \7926 );
nor \U$12290 ( \13132 , \13130 , \13131 );
and \U$12291 ( \13133 , \7914 , RIb559270_509);
and \U$12292 ( \13134 , RIb5592e8_510, \7910 );
nor \U$12293 ( \13135 , \13133 , \13134 );
nand \U$12294 ( \13136 , \13126 , \13129 , \13132 , \13135 );
nor \U$12295 ( \13137 , \13123 , \13136 );
nand \U$12296 ( \13138 , \13116 , \13119 , \13122 , \13137 );
_DC g256e ( \13139_nG256e , \13138 , \11786 );
nand \U$12297 ( \13140 , \13139_nG256e , \11757 );
and \U$12298 ( \13141 , \12918_nG26c6 , \11944 );
and \U$12299 ( \13142 , \11946 , \12959_nG2600 );
nand \U$12300 ( \13143 , \12918_nG26c6 , \11804 );
or \U$12301 ( \13144 , \11800 , \12959_nG2600 );
nand \U$12302 ( \13145 , \13144 , \11836 );
and \U$12303 ( \13146 , \13143 , \13145 );
nor \U$12304 ( \13147 , \13141 , \13142 , \13146 );
or \U$12305 ( \13148 , \13140 , \13147 );
not \U$12306 ( \13149 , \13054 );
or \U$12307 ( \13150 , \13081 , \13149 );
nand \U$12308 ( \13151 , \13113 , \13148 , \13150 );
not \U$12309 ( \13152 , \13151 );
not \U$12310 ( \13153 , \13096 );
not \U$12311 ( \13154 , \13099 );
and \U$12312 ( \13155 , \13153 , \13154 );
and \U$12313 ( \13156 , \13096 , \13099 );
nor \U$12314 ( \13157 , \13155 , \13156 );
not \U$12315 ( \13158 , \13157 );
or \U$12316 ( \13159 , \13152 , \13158 );
or \U$12317 ( \13160 , \13157 , \13151 );
nand \U$12318 ( \13161 , \13159 , \13160 );
not \U$12319 ( \13162 , \13061 );
xor \U$12320 ( \13163 , \13069 , \13079 );
not \U$12321 ( \13164 , \13163 );
or \U$12322 ( \13165 , \13162 , \13164 );
or \U$12323 ( \13166 , \13163 , \13061 );
nand \U$12324 ( \13167 , \13165 , \13166 );
nand \U$12325 ( \13168 , \12682_nG2848 , \12054 );
or \U$12326 ( \13169 , \11985 , \12741_nG2776 );
nand \U$12327 ( \13170 , \13169 , \12060 );
and \U$12328 ( \13171 , \13168 , \13170 );
and \U$12329 ( \13172 , \12056 , \12741_nG2776 );
and \U$12330 ( \13173 , \12682_nG2848 , \12247 );
nor \U$12331 ( \13174 , \13171 , \13172 , \13173 );
nand \U$12332 ( \13175 , \12543_nG292b , \12226 );
or \U$12333 ( \13176 , \12229 , \12210_nG2a23 );
nand \U$12334 ( \13177 , \13176 , \12231 );
and \U$12335 ( \13178 , \13175 , \13177 );
and \U$12336 ( \13179 , \12234 , \12210_nG2a23 );
and \U$12337 ( \13180 , \12543_nG292b , \12238 );
nor \U$12338 ( \13181 , \13178 , \13179 , \13180 );
xor \U$12339 ( \13182 , \13174 , \13181 );
and \U$12340 ( \13183 , \12959_nG2600 , \11894 );
and \U$12341 ( \13184 , \11936 , \12918_nG26c6 );
nand \U$12342 ( \13185 , \12959_nG2600 , \11891 );
or \U$12343 ( \13186 , \11852 , \12918_nG26c6 );
nand \U$12344 ( \13187 , \13186 , \11940 );
and \U$12345 ( \13188 , \13185 , \13187 );
nor \U$12346 ( \13189 , \13183 , \13184 , \13188 );
and \U$12347 ( \13190 , \13182 , \13189 );
and \U$12348 ( \13191 , \13174 , \13181 );
or \U$12349 ( \13192 , \13190 , \13191 );
nand \U$12350 ( \13193 , \12089_nG2d11 , \12607 );
or \U$12351 ( \13194 , \12569 , \12038_nG2e11 );
nand \U$12352 ( \13195 , \13194 , \12791 );
and \U$12353 ( \13196 , \13193 , \13195 );
and \U$12354 ( \13197 , \12794 , \12038_nG2e11 );
and \U$12355 ( \13198 , \12089_nG2d11 , \12609 );
nor \U$12356 ( \13199 , \13196 , \13197 , \13198 );
and \U$12357 ( \13200 , \11901 , \13063 );
not \U$12358 ( \13201 , \11972_nG2efb );
and \U$12359 ( \13202 , \12886 , \13201 );
and \U$12360 ( \13203 , \11879_nG301d , \13067 );
nor \U$12361 ( \13204 , \13200 , \13202 , \13203 );
xor \U$12362 ( \13205 , \13199 , \13204 );
and \U$12363 ( \13206 , \12142_nG2c0d , \12553 );
or \U$12364 ( \13207 , \12258 , \12142_nG2c0d );
nand \U$12365 ( \13208 , \13207 , \12556 );
nand \U$12366 ( \13209 , \12169_nG2b05 , \12409 );
and \U$12367 ( \13210 , \13208 , \13209 );
and \U$12368 ( \13211 , \12169_nG2b05 , \12412 );
nor \U$12369 ( \13212 , \13206 , \13210 , \13211 );
and \U$12370 ( \13213 , \13205 , \13212 );
and \U$12371 ( \13214 , \13199 , \13204 );
or \U$12372 ( \13215 , \13213 , \13214 );
nor \U$12373 ( \13216 , \13192 , \13215 );
and \U$12374 ( \13217 , \13167 , \13216 );
xor \U$12375 ( \13218 , \13161 , \13217 );
xor \U$12376 ( \13219 , \13036 , \13043 );
xor \U$12377 ( \13220 , \13219 , \13051 );
not \U$12378 ( \13221 , \13220 );
xor \U$12379 ( \13222 , \13140 , \13147 );
and \U$12380 ( \13223 , \13221 , \13222 );
not \U$12381 ( \13224 , \13223 );
nand \U$12382 ( \13225 , \12210_nG2a23 , \12226 );
or \U$12383 ( \13226 , \12229 , \12169_nG2b05 );
nand \U$12384 ( \13227 , \13226 , \12231 );
and \U$12385 ( \13228 , \13225 , \13227 );
and \U$12386 ( \13229 , \12234 , \12169_nG2b05 );
and \U$12387 ( \13230 , \12210_nG2a23 , \12238 );
nor \U$12388 ( \13231 , \13228 , \13229 , \13230 );
and \U$12389 ( \13232 , \12089_nG2d11 , \12553 );
or \U$12390 ( \13233 , \12258 , \12089_nG2d11 );
nand \U$12391 ( \13234 , \13233 , \12556 );
nand \U$12392 ( \13235 , \12142_nG2c0d , \12409 );
and \U$12393 ( \13236 , \13234 , \13235 );
and \U$12394 ( \13237 , \12142_nG2c0d , \12412 );
nor \U$12395 ( \13238 , \13232 , \13236 , \13237 );
xor \U$12396 ( \13239 , \13231 , \13238 );
nand \U$12397 ( \13240 , \12543_nG292b , \12054 );
or \U$12398 ( \13241 , \11985 , \12682_nG2848 );
nand \U$12399 ( \13242 , \13241 , \12060 );
and \U$12400 ( \13243 , \13240 , \13242 );
and \U$12401 ( \13244 , \12056 , \12682_nG2848 );
and \U$12402 ( \13245 , \12543_nG292b , \12247 );
nor \U$12403 ( \13246 , \13243 , \13244 , \13245 );
and \U$12404 ( \13247 , \13239 , \13246 );
and \U$12405 ( \13248 , \13231 , \13238 );
or \U$12406 ( \13249 , \13247 , \13248 );
and \U$12407 ( \13250 , \12959_nG2600 , \11944 );
and \U$12408 ( \13251 , \11946 , \13139_nG256e );
nand \U$12409 ( \13252 , \12959_nG2600 , \11804 );
or \U$12410 ( \13253 , \11800 , \13139_nG256e );
nand \U$12411 ( \13254 , \13253 , \11836 );
and \U$12412 ( \13255 , \13252 , \13254 );
nor \U$12413 ( \13256 , \13250 , \13251 , \13255 );
and \U$12414 ( \13257 , \12918_nG26c6 , \11894 );
and \U$12415 ( \13258 , \11936 , \12741_nG2776 );
nand \U$12416 ( \13259 , \12918_nG26c6 , \11891 );
or \U$12417 ( \13260 , \11852 , \12741_nG2776 );
nand \U$12418 ( \13261 , \13260 , \11940 );
and \U$12419 ( \13262 , \13259 , \13261 );
nor \U$12420 ( \13263 , \13257 , \13258 , \13262 );
and \U$12421 ( \13264 , \13256 , \13263 );
not \U$12422 ( \13265 , \13264 );
and \U$12423 ( \13266 , \11760 , RIb5587a8_486);
and \U$12424 ( \13267 , RIb558dc0_499, \7936 );
nor \U$12425 ( \13268 , \13266 , \13267 );
and \U$12426 ( \13269 , \7938 , RIb558d48_498);
and \U$12427 ( \13270 , RIb558be0_495, \7955 );
nor \U$12428 ( \13271 , \13269 , \13270 );
and \U$12429 ( \13272 , \7950 , RIb558898_488);
and \U$12430 ( \13273 , RIb558910_489, \7900 );
nor \U$12431 ( \13274 , \13272 , \13273 );
and \U$12432 ( \13275 , \7917 , RIb558820_487);
and \U$12433 ( \13276 , \7943 , RIb558c58_496);
and \U$12434 ( \13277 , RIb558b68_494, \7926 );
nor \U$12435 ( \13278 , \13276 , \13277 );
and \U$12436 ( \13279 , \7914 , RIb558a78_492);
and \U$12437 ( \13280 , RIb558af0_493, \7910 );
nor \U$12438 ( \13281 , \13279 , \13280 );
and \U$12439 ( \13282 , \7948 , RIb558e38_500);
and \U$12440 ( \13283 , RIb558cd0_497, \7945 );
nor \U$12441 ( \13284 , \13282 , \13283 );
and \U$12442 ( \13285 , \7906 , RIb558a00_491);
and \U$12443 ( \13286 , RIb558988_490, \7953 );
nor \U$12444 ( \13287 , \13285 , \13286 );
nand \U$12445 ( \13288 , \13278 , \13281 , \13284 , \13287 );
nor \U$12446 ( \13289 , \13275 , \13288 );
nand \U$12447 ( \13290 , \13268 , \13271 , \13274 , \13289 );
_DC g24d0 ( \13291_nG24d0 , \13290 , \11786 );
nand \U$12448 ( \13292 , \13291_nG24d0 , \11757 );
not \U$12449 ( \13293 , \13292 );
and \U$12450 ( \13294 , \13265 , \13293 );
nor \U$12451 ( \13295 , \13256 , \13263 );
nor \U$12452 ( \13296 , \13294 , \13295 );
nand \U$12453 ( \13297 , \13249 , \13296 );
or \U$12454 ( \13298 , \13066 , \11788 );
or \U$12455 ( \13299 , \11787_nG3124 , \12888 );
or \U$12456 ( \13300 , \11879_nG301d , \12887 );
nand \U$12457 ( \13301 , \13298 , \13299 , \13300 );
or \U$12458 ( \13302 , \12610 , \12330 );
or \U$12459 ( \13303 , \12569 , \11972_nG2efb );
nand \U$12460 ( \13304 , \13303 , \12791 );
nand \U$12461 ( \13305 , \12038_nG2e11 , \12607 );
and \U$12462 ( \13306 , \13304 , \13305 );
and \U$12463 ( \13307 , \11972_nG2efb , \12794 );
nor \U$12464 ( \13308 , \13306 , \13307 );
nand \U$12465 ( \13309 , \13302 , \13308 );
and \U$12466 ( \13310 , \13301 , \13309 );
and \U$12467 ( \13311 , \13297 , \13310 );
nor \U$12468 ( \13312 , \13296 , \13249 );
nor \U$12469 ( \13313 , \13311 , \13312 );
not \U$12470 ( \13314 , \12881 );
not \U$12471 ( \13315 , \12889 );
and \U$12472 ( \13316 , \13314 , \13315 );
and \U$12473 ( \13317 , \12881 , \12889 );
nor \U$12474 ( \13318 , \13316 , \13317 );
nor \U$12475 ( \13319 , \13313 , \13318 );
not \U$12476 ( \13320 , \13319 );
nand \U$12477 ( \13321 , \13318 , \13313 );
nand \U$12478 ( \13322 , \13320 , \13321 );
not \U$12479 ( \13323 , \13322 );
or \U$12480 ( \13324 , \13224 , \13323 );
or \U$12481 ( \13325 , \13322 , \13223 );
nand \U$12482 ( \13326 , \13324 , \13325 );
and \U$12483 ( \13327 , \13218 , \13326 );
and \U$12484 ( \13328 , \13161 , \13217 );
or \U$12485 ( \13329 , \13327 , \13328 );
xor \U$12486 ( \13330 , \13082 , \13089 );
xor \U$12487 ( \13331 , \13330 , \13100 );
xor \U$12488 ( \13332 , \13329 , \13331 );
not \U$12489 ( \13333 , \13157 );
nand \U$12490 ( \13334 , \13333 , \13151 );
not \U$12491 ( \13335 , \13334 );
and \U$12492 ( \13336 , \13321 , \13223 );
nor \U$12493 ( \13337 , \13336 , \13319 );
xor \U$12494 ( \13338 , \13020 , \13022 );
xor \U$12495 ( \13339 , \13338 , \13025 );
nor \U$12496 ( \13340 , \13337 , \13339 );
and \U$12497 ( \13341 , \13337 , \13339 );
nor \U$12498 ( \13342 , \13340 , \13341 );
not \U$12499 ( \13343 , \13342 );
or \U$12500 ( \13344 , \13335 , \13343 );
or \U$12501 ( \13345 , \13342 , \13334 );
nand \U$12502 ( \13346 , \13344 , \13345 );
and \U$12503 ( \13347 , \13332 , \13346 );
and \U$12504 ( \13348 , \13329 , \13331 );
or \U$12505 ( \13349 , \13347 , \13348 );
not \U$12506 ( \13350 , \13341 );
not \U$12507 ( \13351 , \13334 );
and \U$12508 ( \13352 , \13350 , \13351 );
nor \U$12509 ( \13353 , \13352 , \13340 );
not \U$12510 ( \13354 , \13011 );
not \U$12511 ( \13355 , \13018 );
and \U$12512 ( \13356 , \13354 , \13355 );
and \U$12513 ( \13357 , \13011 , \13018 );
nor \U$12514 ( \13358 , \13356 , \13357 );
nand \U$12515 ( \13359 , \13353 , \13358 );
not \U$12516 ( \13360 , \13359 );
nor \U$12517 ( \13361 , \13358 , \13353 );
nor \U$12518 ( \13362 , \13360 , \13361 );
not \U$12519 ( \13363 , \13362 );
not \U$12520 ( \13364 , \13028 );
not \U$12521 ( \13365 , \13103 );
and \U$12522 ( \13366 , \13364 , \13365 );
and \U$12523 ( \13367 , \13028 , \13103 );
nor \U$12524 ( \13368 , \13366 , \13367 );
not \U$12525 ( \13369 , \13368 );
and \U$12526 ( \13370 , \13363 , \13369 );
and \U$12527 ( \13371 , \13362 , \13368 );
nor \U$12528 ( \13372 , \13370 , \13371 );
xor \U$12529 ( \13373 , \13349 , \13372 );
xor \U$12530 ( \13374 , \13329 , \13331 );
xor \U$12531 ( \13375 , \13374 , \13346 );
not \U$12532 ( \13376 , \13215 );
or \U$12533 ( \13377 , \13192 , \13376 );
and \U$12534 ( \13378 , \11760 , RIb559f90_537);
and \U$12535 ( \13379 , RIb55a5a8_550, \7936 );
nor \U$12536 ( \13380 , \13378 , \13379 );
and \U$12537 ( \13381 , \7938 , RIb55a530_549);
and \U$12538 ( \13382 , RIb55a3c8_546, \7955 );
nor \U$12539 ( \13383 , \13381 , \13382 );
and \U$12540 ( \13384 , \7950 , RIb55a080_539);
and \U$12541 ( \13385 , RIb55a0f8_540, \7900 );
nor \U$12542 ( \13386 , \13384 , \13385 );
and \U$12543 ( \13387 , \7917 , RIb55a008_538);
and \U$12544 ( \13388 , \7943 , RIb55a440_547);
and \U$12545 ( \13389 , RIb55a350_545, \7926 );
nor \U$12546 ( \13390 , \13388 , \13389 );
and \U$12547 ( \13391 , \7914 , RIb55a260_543);
and \U$12548 ( \13392 , RIb55a2d8_544, \7910 );
nor \U$12549 ( \13393 , \13391 , \13392 );
and \U$12550 ( \13394 , \7948 , RIb55a620_551);
and \U$12551 ( \13395 , RIb55a4b8_548, \7945 );
nor \U$12552 ( \13396 , \13394 , \13395 );
and \U$12553 ( \13397 , \7906 , RIb55a1e8_542);
and \U$12554 ( \13398 , RIb55a170_541, \7953 );
nor \U$12555 ( \13399 , \13397 , \13398 );
nand \U$12556 ( \13400 , \13390 , \13393 , \13396 , \13399 );
nor \U$12557 ( \13401 , \13387 , \13400 );
nand \U$12558 ( \13402 , \13380 , \13383 , \13386 , \13401 );
_DC g245a ( \13403_nG245a , \13402 , \11786 );
nand \U$12559 ( \13404 , \13403_nG245a , \11757 );
and \U$12560 ( \13405 , \13139_nG256e , \11944 );
and \U$12561 ( \13406 , \11946 , \13291_nG24d0 );
nand \U$12562 ( \13407 , \13139_nG256e , \11804 );
or \U$12563 ( \13408 , \11800 , \13291_nG24d0 );
nand \U$12564 ( \13409 , \13408 , \11836 );
and \U$12565 ( \13410 , \13407 , \13409 );
nor \U$12566 ( \13411 , \13405 , \13406 , \13410 );
or \U$12567 ( \13412 , \13404 , \13411 );
not \U$12568 ( \13413 , \13192 );
or \U$12569 ( \13414 , \13215 , \13413 );
nand \U$12570 ( \13415 , \13377 , \13412 , \13414 );
xor \U$12571 ( \13416 , \13301 , \13309 );
xor \U$12572 ( \13417 , \13415 , \13416 );
not \U$12573 ( \13418 , \13292 );
nor \U$12574 ( \13419 , \13264 , \13295 );
not \U$12575 ( \13420 , \13419 );
or \U$12576 ( \13421 , \13418 , \13420 );
or \U$12577 ( \13422 , \13419 , \13292 );
nand \U$12578 ( \13423 , \13421 , \13422 );
and \U$12579 ( \13424 , \13417 , \13423 );
and \U$12580 ( \13425 , \13415 , \13416 );
or \U$12581 ( \13426 , \13424 , \13425 );
xor \U$12582 ( \13427 , \13221 , \13222 );
xor \U$12583 ( \13428 , \13426 , \13427 );
xnor \U$12584 ( \13429 , \13404 , \13411 );
xor \U$12585 ( \13430 , \13174 , \13181 );
xor \U$12586 ( \13431 , \13430 , \13189 );
and \U$12587 ( \13432 , \13429 , \13431 );
not \U$12588 ( \13433 , \13432 );
xor \U$12589 ( \13434 , \13199 , \13204 );
xor \U$12590 ( \13435 , \13434 , \13212 );
not \U$12591 ( \13436 , \13435 );
and \U$12592 ( \13437 , \13433 , \13436 );
nor \U$12593 ( \13438 , \13429 , \13431 );
nor \U$12594 ( \13439 , \13437 , \13438 );
xor \U$12595 ( \13440 , \13231 , \13238 );
xor \U$12596 ( \13441 , \13440 , \13246 );
xor \U$12597 ( \13442 , \13439 , \13441 );
nand \U$12598 ( \13443 , \12682_nG2848 , \12226 );
or \U$12599 ( \13444 , \12229 , \12543_nG292b );
nand \U$12600 ( \13445 , \13444 , \12231 );
and \U$12601 ( \13446 , \13443 , \13445 );
and \U$12602 ( \13447 , \12234 , \12543_nG292b );
and \U$12603 ( \13448 , \12682_nG2848 , \12238 );
nor \U$12604 ( \13449 , \13446 , \13447 , \13448 );
and \U$12605 ( \13450 , \12169_nG2b05 , \12553 );
or \U$12606 ( \13451 , \12258 , \12169_nG2b05 );
nand \U$12607 ( \13452 , \13451 , \12556 );
nand \U$12608 ( \13453 , \12210_nG2a23 , \12409 );
and \U$12609 ( \13454 , \13452 , \13453 );
and \U$12610 ( \13455 , \12210_nG2a23 , \12412 );
nor \U$12611 ( \13456 , \13450 , \13454 , \13455 );
xor \U$12612 ( \13457 , \13449 , \13456 );
nand \U$12613 ( \13458 , \12741_nG2776 , \12054 );
or \U$12614 ( \13459 , \11985 , \12918_nG26c6 );
nand \U$12615 ( \13460 , \13459 , \12060 );
and \U$12616 ( \13461 , \13458 , \13460 );
and \U$12617 ( \13462 , \12056 , \12918_nG26c6 );
and \U$12618 ( \13463 , \12741_nG2776 , \12247 );
nor \U$12619 ( \13464 , \13461 , \13462 , \13463 );
and \U$12620 ( \13465 , \13457 , \13464 );
and \U$12621 ( \13466 , \13449 , \13456 );
or \U$12622 ( \13467 , \13465 , \13466 );
nand \U$12623 ( \13468 , \12142_nG2c0d , \12607 );
or \U$12624 ( \13469 , \12569 , \12089_nG2d11 );
nand \U$12625 ( \13470 , \13469 , \12791 );
and \U$12626 ( \13471 , \13468 , \13470 );
and \U$12627 ( \13472 , \12794 , \12089_nG2d11 );
and \U$12628 ( \13473 , \12142_nG2c0d , \12609 );
nor \U$12629 ( \13474 , \13471 , \13472 , \13473 );
not \U$12630 ( \13475 , \13474 );
or \U$12631 ( \13476 , \13066 , \13201 );
or \U$12632 ( \13477 , \11972_nG2efb , \12888 );
or \U$12633 ( \13478 , \12038_nG2e11 , \12887 );
nand \U$12634 ( \13479 , \13476 , \13477 , \13478 );
nand \U$12635 ( \13480 , \13475 , \13479 );
xor \U$12636 ( \13481 , \13467 , \13480 );
and \U$12637 ( \13482 , \13291_nG24d0 , \11944 );
and \U$12638 ( \13483 , \11946 , \13403_nG245a );
nand \U$12639 ( \13484 , \13291_nG24d0 , \11804 );
or \U$12640 ( \13485 , \11800 , \13403_nG245a );
nand \U$12641 ( \13486 , \13485 , \11836 );
and \U$12642 ( \13487 , \13484 , \13486 );
nor \U$12643 ( \13488 , \13482 , \13483 , \13487 );
and \U$12644 ( \13489 , \13139_nG256e , \11894 );
and \U$12645 ( \13490 , \11936 , \12959_nG2600 );
nand \U$12646 ( \13491 , \13139_nG256e , \11891 );
or \U$12647 ( \13492 , \11852 , \12959_nG2600 );
nand \U$12648 ( \13493 , \13492 , \11940 );
and \U$12649 ( \13494 , \13491 , \13493 );
nor \U$12650 ( \13495 , \13489 , \13490 , \13494 );
and \U$12651 ( \13496 , \13488 , \13495 );
not \U$12652 ( \13497 , \13496 );
and \U$12653 ( \13498 , \11760 , RIb559798_520);
and \U$12654 ( \13499 , RIb559db0_533, \7936 );
nor \U$12655 ( \13500 , \13498 , \13499 );
and \U$12656 ( \13501 , \7938 , RIb559d38_532);
and \U$12657 ( \13502 , RIb559bd0_529, \7955 );
nor \U$12658 ( \13503 , \13501 , \13502 );
and \U$12659 ( \13504 , \7950 , RIb559888_522);
and \U$12660 ( \13505 , RIb559900_523, \7900 );
nor \U$12661 ( \13506 , \13504 , \13505 );
and \U$12662 ( \13507 , \7917 , RIb559810_521);
and \U$12663 ( \13508 , \7906 , RIb5599f0_525);
and \U$12664 ( \13509 , RIb559978_524, \7953 );
nor \U$12665 ( \13510 , \13508 , \13509 );
and \U$12666 ( \13511 , \7943 , RIb559c48_530);
and \U$12667 ( \13512 , RIb559cc0_531, \7945 );
nor \U$12668 ( \13513 , \13511 , \13512 );
and \U$12669 ( \13514 , \7948 , RIb559e28_534);
and \U$12670 ( \13515 , RIb559b58_528, \7926 );
nor \U$12671 ( \13516 , \13514 , \13515 );
and \U$12672 ( \13517 , \7914 , RIb559a68_526);
and \U$12673 ( \13518 , RIb559ae0_527, \7910 );
nor \U$12674 ( \13519 , \13517 , \13518 );
nand \U$12675 ( \13520 , \13510 , \13513 , \13516 , \13519 );
nor \U$12676 ( \13521 , \13507 , \13520 );
nand \U$12677 ( \13522 , \13500 , \13503 , \13506 , \13521 );
_DC g23dc ( \13523_nG23dc , \13522 , \11786 );
nand \U$12678 ( \13524 , \13523_nG23dc , \11757 );
not \U$12679 ( \13525 , \13524 );
and \U$12680 ( \13526 , \13497 , \13525 );
nor \U$12681 ( \13527 , \13488 , \13495 );
nor \U$12682 ( \13528 , \13526 , \13527 );
and \U$12683 ( \13529 , \13481 , \13528 );
and \U$12684 ( \13530 , \13467 , \13480 );
or \U$12685 ( \13531 , \13529 , \13530 );
and \U$12686 ( \13532 , \13442 , \13531 );
and \U$12687 ( \13533 , \13439 , \13441 );
or \U$12688 ( \13534 , \13532 , \13533 );
not \U$12689 ( \13535 , \13534 );
and \U$12690 ( \13536 , \13428 , \13535 );
and \U$12691 ( \13537 , \13426 , \13427 );
or \U$12692 ( \13538 , \13536 , \13537 );
xor \U$12693 ( \13539 , \13167 , \13216 );
not \U$12694 ( \13540 , \13310 );
not \U$12695 ( \13541 , \13312 );
nand \U$12696 ( \13542 , \13541 , \13297 );
not \U$12697 ( \13543 , \13542 );
or \U$12698 ( \13544 , \13540 , \13543 );
or \U$12699 ( \13545 , \13542 , \13310 );
nand \U$12700 ( \13546 , \13544 , \13545 );
and \U$12701 ( \13547 , \13539 , \13546 );
xor \U$12702 ( \13548 , \13538 , \13547 );
xor \U$12703 ( \13549 , \13161 , \13217 );
xor \U$12704 ( \13550 , \13549 , \13326 );
and \U$12705 ( \13551 , \13548 , \13550 );
and \U$12706 ( \13552 , \13538 , \13547 );
or \U$12707 ( \13553 , \13551 , \13552 );
xor \U$12708 ( \13554 , \13375 , \13553 );
xor \U$12709 ( \13555 , \13415 , \13416 );
xor \U$12710 ( \13556 , \13555 , \13423 );
not \U$12711 ( \13557 , \13556 );
not \U$12712 ( \13558 , \13524 );
nor \U$12713 ( \13559 , \13496 , \13527 );
not \U$12714 ( \13560 , \13559 );
or \U$12715 ( \13561 , \13558 , \13560 );
or \U$12716 ( \13562 , \13559 , \13524 );
nand \U$12717 ( \13563 , \13561 , \13562 );
not \U$12718 ( \13564 , \13563 );
xor \U$12719 ( \13565 , \13449 , \13456 );
xor \U$12720 ( \13566 , \13565 , \13464 );
nor \U$12721 ( \13567 , \13564 , \13566 );
nand \U$12722 ( \13568 , \12918_nG26c6 , \12054 );
or \U$12723 ( \13569 , \11985 , \12959_nG2600 );
nand \U$12724 ( \13570 , \13569 , \12060 );
and \U$12725 ( \13571 , \13568 , \13570 );
and \U$12726 ( \13572 , \12056 , \12959_nG2600 );
and \U$12727 ( \13573 , \12918_nG26c6 , \12247 );
nor \U$12728 ( \13574 , \13571 , \13572 , \13573 );
nand \U$12729 ( \13575 , \12741_nG2776 , \12226 );
or \U$12730 ( \13576 , \12229 , \12682_nG2848 );
nand \U$12731 ( \13577 , \13576 , \12231 );
and \U$12732 ( \13578 , \13575 , \13577 );
and \U$12733 ( \13579 , \12234 , \12682_nG2848 );
and \U$12734 ( \13580 , \12741_nG2776 , \12238 );
nor \U$12735 ( \13581 , \13578 , \13579 , \13580 );
xor \U$12736 ( \13582 , \13574 , \13581 );
and \U$12737 ( \13583 , \13291_nG24d0 , \11894 );
and \U$12738 ( \13584 , \11936 , \13139_nG256e );
nand \U$12739 ( \13585 , \13291_nG24d0 , \11891 );
or \U$12740 ( \13586 , \11852 , \13139_nG256e );
nand \U$12741 ( \13587 , \13586 , \11940 );
and \U$12742 ( \13588 , \13585 , \13587 );
nor \U$12743 ( \13589 , \13583 , \13584 , \13588 );
and \U$12744 ( \13590 , \13582 , \13589 );
and \U$12745 ( \13591 , \13574 , \13581 );
or \U$12746 ( \13592 , \13590 , \13591 );
nand \U$12747 ( \13593 , \12169_nG2b05 , \12607 );
or \U$12748 ( \13594 , \12569 , \12142_nG2c0d );
nand \U$12749 ( \13595 , \13594 , \12791 );
and \U$12750 ( \13596 , \13593 , \13595 );
and \U$12751 ( \13597 , \12794 , \12142_nG2c0d );
and \U$12752 ( \13598 , \12169_nG2b05 , \12609 );
nor \U$12753 ( \13599 , \13596 , \13597 , \13598 );
and \U$12754 ( \13600 , \12330 , \13063 );
and \U$12755 ( \13601 , \12886 , \12332 );
and \U$12756 ( \13602 , \12038_nG2e11 , \13067 );
nor \U$12757 ( \13603 , \13600 , \13601 , \13602 );
xor \U$12758 ( \13604 , \13599 , \13603 );
and \U$12759 ( \13605 , \12210_nG2a23 , \12553 );
or \U$12760 ( \13606 , \12258 , \12210_nG2a23 );
nand \U$12761 ( \13607 , \13606 , \12556 );
nand \U$12762 ( \13608 , \12543_nG292b , \12409 );
and \U$12763 ( \13609 , \13607 , \13608 );
and \U$12764 ( \13610 , \12543_nG292b , \12412 );
nor \U$12765 ( \13611 , \13605 , \13609 , \13610 );
and \U$12766 ( \13612 , \13604 , \13611 );
and \U$12767 ( \13613 , \13599 , \13603 );
or \U$12768 ( \13614 , \13612 , \13613 );
nor \U$12769 ( \13615 , \13592 , \13614 );
xor \U$12770 ( \13616 , \13567 , \13615 );
not \U$12771 ( \13617 , \13435 );
nor \U$12772 ( \13618 , \13432 , \13438 );
not \U$12773 ( \13619 , \13618 );
or \U$12774 ( \13620 , \13617 , \13619 );
or \U$12775 ( \13621 , \13618 , \13435 );
nand \U$12776 ( \13622 , \13620 , \13621 );
and \U$12777 ( \13623 , \13616 , \13622 );
and \U$12778 ( \13624 , \13567 , \13615 );
or \U$12779 ( \13625 , \13623 , \13624 );
not \U$12780 ( \13626 , \13625 );
or \U$12781 ( \13627 , \13557 , \13626 );
xor \U$12782 ( \13628 , \13439 , \13441 );
xor \U$12783 ( \13629 , \13628 , \13531 );
nor \U$12784 ( \13630 , \13625 , \13556 );
or \U$12785 ( \13631 , \13629 , \13630 );
nand \U$12786 ( \13632 , \13627 , \13631 );
xor \U$12787 ( \13633 , \13539 , \13546 );
xor \U$12788 ( \13634 , \13632 , \13633 );
xor \U$12789 ( \13635 , \13426 , \13427 );
xor \U$12790 ( \13636 , \13635 , \13535 );
and \U$12791 ( \13637 , \13634 , \13636 );
and \U$12792 ( \13638 , \13632 , \13633 );
or \U$12793 ( \13639 , \13637 , \13638 );
xor \U$12794 ( \13640 , \13538 , \13547 );
xor \U$12795 ( \13641 , \13640 , \13550 );
xor \U$12796 ( \13642 , \13639 , \13641 );
xor \U$12797 ( \13643 , \13632 , \13633 );
xor \U$12798 ( \13644 , \13643 , \13636 );
not \U$12799 ( \13645 , \13629 );
not \U$12800 ( \13646 , \13625 );
and \U$12801 ( \13647 , \13645 , \13646 );
and \U$12802 ( \13648 , \13629 , \13625 );
nor \U$12803 ( \13649 , \13647 , \13648 );
not \U$12804 ( \13650 , \13649 );
not \U$12805 ( \13651 , \13556 );
and \U$12806 ( \13652 , \13650 , \13651 );
and \U$12807 ( \13653 , \13649 , \13556 );
nor \U$12808 ( \13654 , \13652 , \13653 );
xor \U$12809 ( \13655 , \13574 , \13581 );
xor \U$12810 ( \13656 , \13655 , \13589 );
xor \U$12811 ( \13657 , \13599 , \13603 );
xor \U$12812 ( \13658 , \13657 , \13611 );
xor \U$12813 ( \13659 , \13656 , \13658 );
and \U$12814 ( \13660 , \11760 , RIb55a788_554);
and \U$12815 ( \13661 , RIb55acb0_565, \7945 );
nor \U$12816 ( \13662 , \13660 , \13661 );
and \U$12817 ( \13663 , \7943 , RIb55ac38_564);
and \U$12818 ( \13664 , RIb55abc0_563, \7955 );
nor \U$12819 ( \13665 , \13663 , \13664 );
and \U$12820 ( \13666 , \7950 , RIb55a878_556);
and \U$12821 ( \13667 , RIb55a8f0_557, \7900 );
nor \U$12822 ( \13668 , \13666 , \13667 );
and \U$12823 ( \13669 , \7917 , RIb55a800_555);
and \U$12824 ( \13670 , \7906 , RIb55a9e0_559);
and \U$12825 ( \13671 , RIb55a968_558, \7953 );
nor \U$12826 ( \13672 , \13670 , \13671 );
and \U$12827 ( \13673 , \7938 , RIb55ad28_566);
and \U$12828 ( \13674 , RIb55ab48_562, \7926 );
nor \U$12829 ( \13675 , \13673 , \13674 );
and \U$12830 ( \13676 , \7948 , RIb55ae18_568);
and \U$12831 ( \13677 , RIb55ada0_567, \7936 );
nor \U$12832 ( \13678 , \13676 , \13677 );
and \U$12833 ( \13679 , \7914 , RIb55aa58_560);
and \U$12834 ( \13680 , RIb55aad0_561, \7910 );
nor \U$12835 ( \13681 , \13679 , \13680 );
nand \U$12836 ( \13682 , \13672 , \13675 , \13678 , \13681 );
nor \U$12837 ( \13683 , \13669 , \13682 );
nand \U$12838 ( \13684 , \13662 , \13665 , \13668 , \13683 );
_DC g2388 ( \13685_nG2388 , \13684 , \11786 );
nand \U$12839 ( \13686 , \13685_nG2388 , \11757 );
and \U$12840 ( \13687 , \13403_nG245a , \11944 );
and \U$12841 ( \13688 , \11946 , \13523_nG23dc );
nand \U$12842 ( \13689 , \13403_nG245a , \11804 );
or \U$12843 ( \13690 , \11800 , \13523_nG23dc );
nand \U$12844 ( \13691 , \13690 , \11836 );
and \U$12845 ( \13692 , \13689 , \13691 );
nor \U$12846 ( \13693 , \13687 , \13688 , \13692 );
xnor \U$12847 ( \13694 , \13686 , \13693 );
and \U$12848 ( \13695 , \13659 , \13694 );
and \U$12849 ( \13696 , \13656 , \13658 );
or \U$12850 ( \13697 , \13695 , \13696 );
not \U$12851 ( \13698 , \13474 );
not \U$12852 ( \13699 , \13479 );
and \U$12853 ( \13700 , \13698 , \13699 );
and \U$12854 ( \13701 , \13474 , \13479 );
nor \U$12855 ( \13702 , \13700 , \13701 );
xor \U$12856 ( \13703 , \13697 , \13702 );
nand \U$12857 ( \13704 , \12918_nG26c6 , \12226 );
or \U$12858 ( \13705 , \12229 , \12741_nG2776 );
nand \U$12859 ( \13706 , \13705 , \12231 );
and \U$12860 ( \13707 , \13704 , \13706 );
and \U$12861 ( \13708 , \12234 , \12741_nG2776 );
and \U$12862 ( \13709 , \12918_nG26c6 , \12238 );
nor \U$12863 ( \13710 , \13707 , \13708 , \13709 );
and \U$12864 ( \13711 , \12543_nG292b , \12553 );
or \U$12865 ( \13712 , \12258 , \12543_nG292b );
nand \U$12866 ( \13713 , \13712 , \12556 );
nand \U$12867 ( \13714 , \12682_nG2848 , \12409 );
and \U$12868 ( \13715 , \13713 , \13714 );
and \U$12869 ( \13716 , \12682_nG2848 , \12412 );
nor \U$12870 ( \13717 , \13711 , \13715 , \13716 );
xor \U$12871 ( \13718 , \13710 , \13717 );
nand \U$12872 ( \13719 , \12959_nG2600 , \12054 );
or \U$12873 ( \13720 , \11985 , \13139_nG256e );
nand \U$12874 ( \13721 , \13720 , \12060 );
and \U$12875 ( \13722 , \13719 , \13721 );
and \U$12876 ( \13723 , \12056 , \13139_nG256e );
and \U$12877 ( \13724 , \12959_nG2600 , \12247 );
nor \U$12878 ( \13725 , \13722 , \13723 , \13724 );
and \U$12879 ( \13726 , \13718 , \13725 );
and \U$12880 ( \13727 , \13710 , \13717 );
or \U$12881 ( \13728 , \13726 , \13727 );
nand \U$12882 ( \13729 , \12210_nG2a23 , \12607 );
or \U$12883 ( \13730 , \12569 , \12169_nG2b05 );
nand \U$12884 ( \13731 , \13730 , \12791 );
and \U$12885 ( \13732 , \13729 , \13731 );
and \U$12886 ( \13733 , \12794 , \12169_nG2b05 );
and \U$12887 ( \13734 , \12210_nG2a23 , \12609 );
nor \U$12888 ( \13735 , \13732 , \13733 , \13734 );
not \U$12889 ( \13736 , \13735 );
or \U$12890 ( \13737 , \13066 , \12332 );
or \U$12891 ( \13738 , \12089_nG2d11 , \12888 );
or \U$12892 ( \13739 , \12142_nG2c0d , \12887 );
nand \U$12893 ( \13740 , \13737 , \13738 , \13739 );
nand \U$12894 ( \13741 , \13736 , \13740 );
xor \U$12895 ( \13742 , \13728 , \13741 );
and \U$12896 ( \13743 , \13403_nG245a , \11894 );
and \U$12897 ( \13744 , \11936 , \13291_nG24d0 );
nand \U$12898 ( \13745 , \13403_nG245a , \11891 );
or \U$12899 ( \13746 , \11852 , \13291_nG24d0 );
nand \U$12900 ( \13747 , \13746 , \11940 );
and \U$12901 ( \13748 , \13745 , \13747 );
nor \U$12902 ( \13749 , \13743 , \13744 , \13748 );
and \U$12903 ( \13750 , \11760 , RIb55af80_571);
and \U$12904 ( \13751 , RIb55b598_584, \7936 );
nor \U$12905 ( \13752 , \13750 , \13751 );
and \U$12906 ( \13753 , \7938 , RIb55b520_583);
and \U$12907 ( \13754 , RIb55b3b8_580, \7955 );
nor \U$12908 ( \13755 , \13753 , \13754 );
and \U$12909 ( \13756 , \7950 , RIb55b070_573);
and \U$12910 ( \13757 , RIb55b0e8_574, \7900 );
nor \U$12911 ( \13758 , \13756 , \13757 );
and \U$12912 ( \13759 , \7917 , RIb55aff8_572);
and \U$12913 ( \13760 , \7906 , RIb55b1d8_576);
and \U$12914 ( \13761 , RIb55b160_575, \7953 );
nor \U$12915 ( \13762 , \13760 , \13761 );
and \U$12916 ( \13763 , \7914 , RIb55b250_577);
and \U$12917 ( \13764 , RIb55b2c8_578, \7910 );
nor \U$12918 ( \13765 , \13763 , \13764 );
and \U$12919 ( \13766 , \7948 , RIb55b610_585);
and \U$12920 ( \13767 , RIb55b340_579, \7926 );
nor \U$12921 ( \13768 , \13766 , \13767 );
and \U$12922 ( \13769 , \7943 , RIb55b430_581);
and \U$12923 ( \13770 , RIb55b4a8_582, \7945 );
nor \U$12924 ( \13771 , \13769 , \13770 );
nand \U$12925 ( \13772 , \13762 , \13765 , \13768 , \13771 );
nor \U$12926 ( \13773 , \13759 , \13772 );
nand \U$12927 ( \13774 , \13752 , \13755 , \13758 , \13773 );
_DC g2272 ( \13775_nG2272 , \13774 , \11786 );
nand \U$12928 ( \13776 , \13775_nG2272 , \11757 );
xor \U$12929 ( \13777 , \13749 , \13776 );
and \U$12930 ( \13778 , \13523_nG23dc , \11944 );
and \U$12931 ( \13779 , \11946 , \13685_nG2388 );
nand \U$12932 ( \13780 , \13523_nG23dc , \11804 );
or \U$12933 ( \13781 , \11800 , \13685_nG2388 );
nand \U$12934 ( \13782 , \13781 , \11836 );
and \U$12935 ( \13783 , \13780 , \13782 );
nor \U$12936 ( \13784 , \13778 , \13779 , \13783 );
and \U$12937 ( \13785 , \13777 , \13784 );
and \U$12938 ( \13786 , \13749 , \13776 );
or \U$12939 ( \13787 , \13785 , \13786 );
and \U$12940 ( \13788 , \13742 , \13787 );
and \U$12941 ( \13789 , \13728 , \13741 );
or \U$12942 ( \13790 , \13788 , \13789 );
and \U$12943 ( \13791 , \13703 , \13790 );
and \U$12944 ( \13792 , \13697 , \13702 );
or \U$12945 ( \13793 , \13791 , \13792 );
xor \U$12946 ( \13794 , \13467 , \13480 );
xor \U$12947 ( \13795 , \13794 , \13528 );
and \U$12948 ( \13796 , \13793 , \13795 );
not \U$12949 ( \13797 , \13796 );
not \U$12950 ( \13798 , \13563 );
not \U$12951 ( \13799 , \13566 );
and \U$12952 ( \13800 , \13798 , \13799 );
and \U$12953 ( \13801 , \13563 , \13566 );
nor \U$12954 ( \13802 , \13800 , \13801 );
not \U$12955 ( \13803 , \13802 );
not \U$12956 ( \13804 , \13614 );
or \U$12957 ( \13805 , \13592 , \13804 );
or \U$12958 ( \13806 , \13686 , \13693 );
not \U$12959 ( \13807 , \13592 );
or \U$12960 ( \13808 , \13614 , \13807 );
nand \U$12961 ( \13809 , \13805 , \13806 , \13808 );
nand \U$12962 ( \13810 , \13803 , \13809 );
not \U$12963 ( \13811 , \13810 );
and \U$12964 ( \13812 , \13797 , \13811 );
nor \U$12965 ( \13813 , \13793 , \13795 );
nor \U$12966 ( \13814 , \13812 , \13813 );
nor \U$12967 ( \13815 , \13654 , \13814 );
xor \U$12968 ( \13816 , \13644 , \13815 );
and \U$12969 ( \13817 , \13654 , \13814 );
nor \U$12970 ( \13818 , \13817 , \13815 );
xor \U$12971 ( \13819 , \13567 , \13615 );
xor \U$12972 ( \13820 , \13819 , \13622 );
not \U$12973 ( \13821 , \13810 );
nor \U$12974 ( \13822 , \13813 , \13796 );
not \U$12975 ( \13823 , \13822 );
or \U$12976 ( \13824 , \13821 , \13823 );
or \U$12977 ( \13825 , \13822 , \13810 );
nand \U$12978 ( \13826 , \13824 , \13825 );
nand \U$12979 ( \13827 , \13820 , \13826 );
not \U$12980 ( \13828 , \13827 );
xor \U$12981 ( \13829 , \13818 , \13828 );
or \U$12982 ( \13830 , \13826 , \13820 );
nand \U$12983 ( \13831 , \13830 , \13827 );
nand \U$12984 ( \13832 , \13139_nG256e , \12054 );
or \U$12985 ( \13833 , \11985 , \13291_nG24d0 );
nand \U$12986 ( \13834 , \13833 , \12060 );
and \U$12987 ( \13835 , \13832 , \13834 );
and \U$12988 ( \13836 , \12056 , \13291_nG24d0 );
and \U$12989 ( \13837 , \13139_nG256e , \12247 );
nor \U$12990 ( \13838 , \13835 , \13836 , \13837 );
nand \U$12991 ( \13839 , \12959_nG2600 , \12226 );
or \U$12992 ( \13840 , \12229 , \12918_nG26c6 );
nand \U$12993 ( \13841 , \13840 , \12231 );
and \U$12994 ( \13842 , \13839 , \13841 );
and \U$12995 ( \13843 , \12234 , \12918_nG26c6 );
and \U$12996 ( \13844 , \12959_nG2600 , \12238 );
nor \U$12997 ( \13845 , \13842 , \13843 , \13844 );
xor \U$12998 ( \13846 , \13838 , \13845 );
and \U$12999 ( \13847 , \13523_nG23dc , \11894 );
and \U$13000 ( \13848 , \11936 , \13403_nG245a );
nand \U$13001 ( \13849 , \13523_nG23dc , \11891 );
or \U$13002 ( \13850 , \11852 , \13403_nG245a );
nand \U$13003 ( \13851 , \13850 , \11940 );
and \U$13004 ( \13852 , \13849 , \13851 );
nor \U$13005 ( \13853 , \13847 , \13848 , \13852 );
and \U$13006 ( \13854 , \13846 , \13853 );
and \U$13007 ( \13855 , \13838 , \13845 );
or \U$13008 ( \13856 , \13854 , \13855 );
nand \U$13009 ( \13857 , \12543_nG292b , \12607 );
or \U$13010 ( \13858 , \12569 , \12210_nG2a23 );
nand \U$13011 ( \13859 , \13858 , \12791 );
and \U$13012 ( \13860 , \13857 , \13859 );
and \U$13013 ( \13861 , \12794 , \12210_nG2a23 );
and \U$13014 ( \13862 , \12543_nG292b , \12609 );
nor \U$13015 ( \13863 , \13860 , \13861 , \13862 );
and \U$13016 ( \13864 , \12328 , \13063 );
not \U$13017 ( \13865 , \12169_nG2b05 );
and \U$13018 ( \13866 , \12886 , \13865 );
and \U$13019 ( \13867 , \12142_nG2c0d , \13067 );
nor \U$13020 ( \13868 , \13864 , \13866 , \13867 );
xor \U$13021 ( \13869 , \13863 , \13868 );
and \U$13022 ( \13870 , \12682_nG2848 , \12553 );
or \U$13023 ( \13871 , \12258 , \12682_nG2848 );
nand \U$13024 ( \13872 , \13871 , \12556 );
nand \U$13025 ( \13873 , \12741_nG2776 , \12409 );
and \U$13026 ( \13874 , \13872 , \13873 );
and \U$13027 ( \13875 , \12741_nG2776 , \12412 );
nor \U$13028 ( \13876 , \13870 , \13874 , \13875 );
and \U$13029 ( \13877 , \13869 , \13876 );
and \U$13030 ( \13878 , \13863 , \13868 );
or \U$13031 ( \13879 , \13877 , \13878 );
xor \U$13032 ( \13880 , \13856 , \13879 );
xor \U$13033 ( \13881 , \13749 , \13776 );
xor \U$13034 ( \13882 , \13881 , \13784 );
and \U$13035 ( \13883 , \13880 , \13882 );
and \U$13036 ( \13884 , \13856 , \13879 );
or \U$13037 ( \13885 , \13883 , \13884 );
xor \U$13038 ( \13886 , \13710 , \13717 );
xor \U$13039 ( \13887 , \13886 , \13725 );
not \U$13040 ( \13888 , \13887 );
not \U$13041 ( \13889 , \13740 );
not \U$13042 ( \13890 , \13735 );
or \U$13043 ( \13891 , \13889 , \13890 );
or \U$13044 ( \13892 , \13735 , \13740 );
nand \U$13045 ( \13893 , \13891 , \13892 );
nand \U$13046 ( \13894 , \13888 , \13893 );
xor \U$13047 ( \13895 , \13885 , \13894 );
xor \U$13048 ( \13896 , \13656 , \13658 );
xor \U$13049 ( \13897 , \13896 , \13694 );
and \U$13050 ( \13898 , \13895 , \13897 );
and \U$13051 ( \13899 , \13885 , \13894 );
or \U$13052 ( \13900 , \13898 , \13899 );
not \U$13053 ( \13901 , \13802 );
not \U$13054 ( \13902 , \13809 );
and \U$13055 ( \13903 , \13901 , \13902 );
and \U$13056 ( \13904 , \13802 , \13809 );
nor \U$13057 ( \13905 , \13903 , \13904 );
xor \U$13058 ( \13906 , \13900 , \13905 );
xor \U$13059 ( \13907 , \13697 , \13702 );
xor \U$13060 ( \13908 , \13907 , \13790 );
and \U$13061 ( \13909 , \13906 , \13908 );
and \U$13062 ( \13910 , \13900 , \13905 );
or \U$13063 ( \13911 , \13909 , \13910 );
xor \U$13064 ( \13912 , \13831 , \13911 );
not \U$13065 ( \13913 , \13685_nG2388 );
or \U$13066 ( \13914 , \11839 , \13913 );
not \U$13067 ( \13915 , \13775_nG2272 );
or \U$13068 ( \13916 , \13915 , \11806 );
or \U$13069 ( \13917 , \11803 , \13913 );
or \U$13070 ( \13918 , \11800 , \13775_nG2272 );
nand \U$13071 ( \13919 , \13918 , \11836 );
nand \U$13072 ( \13920 , \13917 , \13919 );
nand \U$13073 ( \13921 , \13914 , \13916 , \13920 );
nand \U$13074 ( \13922 , \13139_nG256e , \12226 );
or \U$13075 ( \13923 , \12229 , \12959_nG2600 );
nand \U$13076 ( \13924 , \13923 , \12231 );
and \U$13077 ( \13925 , \13922 , \13924 );
and \U$13078 ( \13926 , \12234 , \12959_nG2600 );
and \U$13079 ( \13927 , \13139_nG256e , \12238 );
nor \U$13080 ( \13928 , \13925 , \13926 , \13927 );
and \U$13081 ( \13929 , \12741_nG2776 , \12553 );
or \U$13082 ( \13930 , \12258 , \12741_nG2776 );
nand \U$13083 ( \13931 , \13930 , \12556 );
nand \U$13084 ( \13932 , \12918_nG26c6 , \12409 );
and \U$13085 ( \13933 , \13931 , \13932 );
and \U$13086 ( \13934 , \12918_nG26c6 , \12412 );
nor \U$13087 ( \13935 , \13929 , \13933 , \13934 );
xor \U$13088 ( \13936 , \13928 , \13935 );
nand \U$13089 ( \13937 , \13291_nG24d0 , \12054 );
or \U$13090 ( \13938 , \11985 , \13403_nG245a );
nand \U$13091 ( \13939 , \13938 , \12060 );
and \U$13092 ( \13940 , \13937 , \13939 );
and \U$13093 ( \13941 , \12056 , \13403_nG245a );
and \U$13094 ( \13942 , \13291_nG24d0 , \12247 );
nor \U$13095 ( \13943 , \13940 , \13941 , \13942 );
and \U$13096 ( \13944 , \13936 , \13943 );
and \U$13097 ( \13945 , \13928 , \13935 );
or \U$13098 ( \13946 , \13944 , \13945 );
nand \U$13099 ( \13947 , \12682_nG2848 , \12607 );
or \U$13100 ( \13948 , \12569 , \12543_nG292b );
nand \U$13101 ( \13949 , \13948 , \12791 );
and \U$13102 ( \13950 , \13947 , \13949 );
and \U$13103 ( \13951 , \12794 , \12543_nG292b );
and \U$13104 ( \13952 , \12682_nG2848 , \12609 );
nor \U$13105 ( \13953 , \13950 , \13951 , \13952 );
and \U$13106 ( \13954 , \13865 , \13063 );
not \U$13107 ( \13955 , \12210_nG2a23 );
and \U$13108 ( \13956 , \12886 , \13955 );
and \U$13109 ( \13957 , \12169_nG2b05 , \13067 );
nor \U$13110 ( \13958 , \13954 , \13956 , \13957 );
xor \U$13111 ( \13959 , \13953 , \13958 );
and \U$13112 ( \13960 , \13959 , \11800 );
and \U$13113 ( \13961 , \13953 , \13958 );
or \U$13114 ( \13962 , \13960 , \13961 );
nand \U$13115 ( \13963 , \13946 , \13962 );
and \U$13116 ( \13964 , \13921 , \13963 );
nor \U$13117 ( \13965 , \13962 , \13946 );
nor \U$13118 ( \13966 , \13964 , \13965 );
not \U$13119 ( \13967 , \13887 );
not \U$13120 ( \13968 , \13893 );
and \U$13121 ( \13969 , \13967 , \13968 );
and \U$13122 ( \13970 , \13887 , \13893 );
nor \U$13123 ( \13971 , \13969 , \13970 );
xor \U$13124 ( \13972 , \13966 , \13971 );
xor \U$13125 ( \13973 , \13856 , \13879 );
xor \U$13126 ( \13974 , \13973 , \13882 );
and \U$13127 ( \13975 , \13972 , \13974 );
and \U$13128 ( \13976 , \13966 , \13971 );
or \U$13129 ( \13977 , \13975 , \13976 );
xor \U$13130 ( \13978 , \13728 , \13741 );
xor \U$13131 ( \13979 , \13978 , \13787 );
xor \U$13132 ( \13980 , \13977 , \13979 );
xor \U$13133 ( \13981 , \13885 , \13894 );
xor \U$13134 ( \13982 , \13981 , \13897 );
and \U$13135 ( \13983 , \13980 , \13982 );
and \U$13136 ( \13984 , \13977 , \13979 );
or \U$13137 ( \13985 , \13983 , \13984 );
xor \U$13138 ( \13986 , \13900 , \13905 );
xor \U$13139 ( \13987 , \13986 , \13908 );
and \U$13140 ( \13988 , \13985 , \13987 );
xor \U$13141 ( \13989 , \13863 , \13868 );
xor \U$13142 ( \13990 , \13989 , \13876 );
not \U$13143 ( \13991 , \13990 );
not \U$13144 ( \13992 , \13965 );
nand \U$13145 ( \13993 , \13992 , \13963 );
not \U$13146 ( \13994 , \13993 );
not \U$13147 ( \13995 , \13921 );
or \U$13148 ( \13996 , \13994 , \13995 );
or \U$13149 ( \13997 , \13921 , \13993 );
nand \U$13150 ( \13998 , \13996 , \13997 );
nand \U$13151 ( \13999 , \13991 , \13998 );
and \U$13152 ( \14000 , \13685_nG2388 , \11894 );
and \U$13153 ( \14001 , \11936 , \13523_nG23dc );
nand \U$13154 ( \14002 , \13685_nG2388 , \11891 );
or \U$13155 ( \14003 , \11852 , \13523_nG23dc );
nand \U$13156 ( \14004 , \14003 , \11940 );
and \U$13157 ( \14005 , \14002 , \14004 );
nor \U$13158 ( \14006 , \14000 , \14001 , \14005 );
nand \U$13159 ( \14007 , \12741_nG2776 , \12607 );
or \U$13160 ( \14008 , \12569 , \12682_nG2848 );
nand \U$13161 ( \14009 , \14008 , \12791 );
and \U$13162 ( \14010 , \14007 , \14009 );
and \U$13163 ( \14011 , \12794 , \12682_nG2848 );
and \U$13164 ( \14012 , \12741_nG2776 , \12609 );
nor \U$13165 ( \14013 , \14010 , \14011 , \14012 );
and \U$13166 ( \14014 , \13955 , \13063 );
and \U$13167 ( \14015 , \12886 , \12762 );
and \U$13168 ( \14016 , \12210_nG2a23 , \13067 );
nor \U$13169 ( \14017 , \14014 , \14015 , \14016 );
xor \U$13170 ( \14018 , \14013 , \14017 );
and \U$13171 ( \14019 , \12918_nG26c6 , \12553 );
or \U$13172 ( \14020 , \12258 , \12918_nG26c6 );
nand \U$13173 ( \14021 , \14020 , \12556 );
nand \U$13174 ( \14022 , \12959_nG2600 , \12409 );
and \U$13175 ( \14023 , \14021 , \14022 );
and \U$13176 ( \14024 , \12959_nG2600 , \12412 );
nor \U$13177 ( \14025 , \14019 , \14023 , \14024 );
and \U$13178 ( \14026 , \14018 , \14025 );
and \U$13179 ( \14027 , \14013 , \14017 );
or \U$13180 ( \14028 , \14026 , \14027 );
xor \U$13181 ( \14029 , \14006 , \14028 );
nand \U$13182 ( \14030 , \13403_nG245a , \12054 );
or \U$13183 ( \14031 , \11985 , \13523_nG23dc );
nand \U$13184 ( \14032 , \14031 , \12060 );
and \U$13185 ( \14033 , \14030 , \14032 );
and \U$13186 ( \14034 , \12056 , \13523_nG23dc );
and \U$13187 ( \14035 , \13403_nG245a , \12247 );
nor \U$13188 ( \14036 , \14033 , \14034 , \14035 );
nand \U$13189 ( \14037 , \13291_nG24d0 , \12226 );
or \U$13190 ( \14038 , \12229 , \13139_nG256e );
nand \U$13191 ( \14039 , \14038 , \12231 );
and \U$13192 ( \14040 , \14037 , \14039 );
and \U$13193 ( \14041 , \12234 , \13139_nG256e );
and \U$13194 ( \14042 , \13291_nG24d0 , \12238 );
nor \U$13195 ( \14043 , \14040 , \14041 , \14042 );
xor \U$13196 ( \14044 , \14036 , \14043 );
and \U$13197 ( \14045 , \13775_nG2272 , \11894 );
and \U$13198 ( \14046 , \11936 , \13685_nG2388 );
nand \U$13199 ( \14047 , \13775_nG2272 , \11891 );
or \U$13200 ( \14048 , \11852 , \13685_nG2388 );
nand \U$13201 ( \14049 , \14048 , \11940 );
and \U$13202 ( \14050 , \14047 , \14049 );
nor \U$13203 ( \14051 , \14045 , \14046 , \14050 );
and \U$13204 ( \14052 , \14044 , \14051 );
and \U$13205 ( \14053 , \14036 , \14043 );
or \U$13206 ( \14054 , \14052 , \14053 );
and \U$13207 ( \14055 , \14029 , \14054 );
and \U$13208 ( \14056 , \14006 , \14028 );
or \U$13209 ( \14057 , \14055 , \14056 );
xor \U$13210 ( \14058 , \13838 , \13845 );
xor \U$13211 ( \14059 , \14058 , \13853 );
xor \U$13212 ( \14060 , \14057 , \14059 );
xor \U$13213 ( \14061 , \13928 , \13935 );
xor \U$13214 ( \14062 , \14061 , \13943 );
xor \U$13215 ( \14063 , \13953 , \13958 );
xor \U$13216 ( \14064 , \14063 , \11800 );
and \U$13217 ( \14065 , \14062 , \14064 );
and \U$13218 ( \14066 , \11944 , \13775_nG2272 );
nand \U$13219 ( \14067 , \13775_nG2272 , \11804 );
and \U$13220 ( \14068 , \14067 , \11799 );
nor \U$13221 ( \14069 , \14066 , \14068 );
xor \U$13222 ( \14070 , \13953 , \13958 );
xor \U$13223 ( \14071 , \14070 , \11800 );
and \U$13224 ( \14072 , \14069 , \14071 );
and \U$13225 ( \14073 , \14062 , \14069 );
or \U$13226 ( \14074 , \14065 , \14072 , \14073 );
and \U$13227 ( \14075 , \14060 , \14074 );
and \U$13228 ( \14076 , \14057 , \14059 );
or \U$13229 ( \14077 , \14075 , \14076 );
xor \U$13230 ( \14078 , \13999 , \14077 );
xor \U$13231 ( \14079 , \13966 , \13971 );
xor \U$13232 ( \14080 , \14079 , \13974 );
and \U$13233 ( \14081 , \14078 , \14080 );
and \U$13234 ( \14082 , \13999 , \14077 );
or \U$13235 ( \14083 , \14081 , \14082 );
xor \U$13236 ( \14084 , \13977 , \13979 );
xor \U$13237 ( \14085 , \14084 , \13982 );
and \U$13238 ( \14086 , \14083 , \14085 );
xor \U$13239 ( \14087 , \14057 , \14059 );
xor \U$13240 ( \14088 , \14087 , \14074 );
nand \U$13241 ( \14089 , \13403_nG245a , \12226 );
or \U$13242 ( \14090 , \12229 , \13291_nG24d0 );
nand \U$13243 ( \14091 , \14090 , \12231 );
and \U$13244 ( \14092 , \14089 , \14091 );
and \U$13245 ( \14093 , \12234 , \13291_nG24d0 );
and \U$13246 ( \14094 , \13403_nG245a , \12238 );
nor \U$13247 ( \14095 , \14092 , \14093 , \14094 );
and \U$13248 ( \14096 , \12959_nG2600 , \12553 );
or \U$13249 ( \14097 , \12258 , \12959_nG2600 );
nand \U$13250 ( \14098 , \14097 , \12556 );
nand \U$13251 ( \14099 , \13139_nG256e , \12409 );
and \U$13252 ( \14100 , \14098 , \14099 );
and \U$13253 ( \14101 , \13139_nG256e , \12412 );
nor \U$13254 ( \14102 , \14096 , \14100 , \14101 );
xor \U$13255 ( \14103 , \14095 , \14102 );
nand \U$13256 ( \14104 , \13523_nG23dc , \12054 );
or \U$13257 ( \14105 , \11985 , \13685_nG2388 );
nand \U$13258 ( \14106 , \14105 , \12060 );
and \U$13259 ( \14107 , \14104 , \14106 );
and \U$13260 ( \14108 , \12056 , \13685_nG2388 );
and \U$13261 ( \14109 , \13523_nG23dc , \12247 );
nor \U$13262 ( \14110 , \14107 , \14108 , \14109 );
and \U$13263 ( \14111 , \14103 , \14110 );
and \U$13264 ( \14112 , \14095 , \14102 );
or \U$13265 ( \14113 , \14111 , \14112 );
nand \U$13266 ( \14114 , \12918_nG26c6 , \12607 );
or \U$13267 ( \14115 , \12569 , \12741_nG2776 );
nand \U$13268 ( \14116 , \14115 , \12791 );
and \U$13269 ( \14117 , \14114 , \14116 );
and \U$13270 ( \14118 , \12794 , \12741_nG2776 );
and \U$13271 ( \14119 , \12918_nG26c6 , \12609 );
nor \U$13272 ( \14120 , \14117 , \14118 , \14119 );
and \U$13273 ( \14121 , \12762 , \13063 );
not \U$13274 ( \14122 , \12682_nG2848 );
and \U$13275 ( \14123 , \12886 , \14122 );
and \U$13276 ( \14124 , \12543_nG292b , \13067 );
nor \U$13277 ( \14125 , \14121 , \14123 , \14124 );
xor \U$13278 ( \14126 , \14120 , \14125 );
and \U$13279 ( \14127 , \14126 , \11852 );
and \U$13280 ( \14128 , \14120 , \14125 );
or \U$13281 ( \14129 , \14127 , \14128 );
xor \U$13282 ( \14130 , \14113 , \14129 );
xor \U$13283 ( \14131 , \14036 , \14043 );
xor \U$13284 ( \14132 , \14131 , \14051 );
and \U$13285 ( \14133 , \14130 , \14132 );
and \U$13286 ( \14134 , \14113 , \14129 );
or \U$13287 ( \14135 , \14133 , \14134 );
xor \U$13288 ( \14136 , \14006 , \14028 );
xor \U$13289 ( \14137 , \14136 , \14054 );
xor \U$13290 ( \14138 , \14135 , \14137 );
xor \U$13291 ( \14139 , \13953 , \13958 );
xor \U$13292 ( \14140 , \14139 , \11800 );
xor \U$13293 ( \14141 , \14062 , \14069 );
xor \U$13294 ( \14142 , \14140 , \14141 );
and \U$13295 ( \14143 , \14138 , \14142 );
and \U$13296 ( \14144 , \14135 , \14137 );
or \U$13297 ( \14145 , \14143 , \14144 );
nand \U$13298 ( \14146 , \14088 , \14145 );
not \U$13299 ( \14147 , \14146 );
nor \U$13300 ( \14148 , \14145 , \14088 );
nor \U$13301 ( \14149 , \14147 , \14148 );
not \U$13302 ( \14150 , \14149 );
not \U$13303 ( \14151 , \13990 );
not \U$13304 ( \14152 , \13998 );
or \U$13305 ( \14153 , \14151 , \14152 );
or \U$13306 ( \14154 , \13998 , \13990 );
nand \U$13307 ( \14155 , \14153 , \14154 );
not \U$13308 ( \14156 , \14155 );
and \U$13309 ( \14157 , \14150 , \14156 );
and \U$13310 ( \14158 , \14149 , \14155 );
nor \U$13311 ( \14159 , \14157 , \14158 );
xor \U$13312 ( \14160 , \14135 , \14137 );
xor \U$13313 ( \14161 , \14160 , \14142 );
nand \U$13314 ( \14162 , \12959_nG2600 , \12607 );
or \U$13315 ( \14163 , \12569 , \12918_nG26c6 );
nand \U$13316 ( \14164 , \14163 , \12791 );
and \U$13317 ( \14165 , \14162 , \14164 );
and \U$13318 ( \14166 , \12794 , \12918_nG26c6 );
and \U$13319 ( \14167 , \12959_nG2600 , \12609 );
nor \U$13320 ( \14168 , \14165 , \14166 , \14167 );
not \U$13321 ( \14169 , \14168 );
and \U$13322 ( \14170 , \14122 , \13063 );
not \U$13323 ( \14171 , \12741_nG2776 );
and \U$13324 ( \14172 , \12886 , \14171 );
and \U$13325 ( \14173 , \12682_nG2848 , \13067 );
nor \U$13326 ( \14174 , \14170 , \14172 , \14173 );
not \U$13327 ( \14175 , \14174 );
and \U$13328 ( \14176 , \14169 , \14175 );
and \U$13329 ( \14177 , \14168 , \14174 );
and \U$13330 ( \14178 , \13139_nG256e , \12553 );
or \U$13331 ( \14179 , \12258 , \13139_nG256e );
nand \U$13332 ( \14180 , \14179 , \12556 );
nand \U$13333 ( \14181 , \13291_nG24d0 , \12409 );
and \U$13334 ( \14182 , \14180 , \14181 );
and \U$13335 ( \14183 , \13291_nG24d0 , \12412 );
nor \U$13336 ( \14184 , \14178 , \14182 , \14183 );
nor \U$13337 ( \14185 , \14177 , \14184 );
nor \U$13338 ( \14186 , \14176 , \14185 );
xor \U$13339 ( \14187 , \14095 , \14102 );
xor \U$13340 ( \14188 , \14187 , \14110 );
and \U$13341 ( \14189 , \14186 , \14188 );
and \U$13342 ( \14190 , \13775_nG2272 , \11936 );
and \U$13343 ( \14191 , \13915 , \11893 );
not \U$13344 ( \14192 , \11940 );
nor \U$13345 ( \14193 , \14190 , \14191 , \14192 );
xor \U$13346 ( \14194 , \14095 , \14102 );
xor \U$13347 ( \14195 , \14194 , \14110 );
and \U$13348 ( \14196 , \14193 , \14195 );
and \U$13349 ( \14197 , \14186 , \14193 );
or \U$13350 ( \14198 , \14189 , \14196 , \14197 );
xor \U$13351 ( \14199 , \14013 , \14017 );
xor \U$13352 ( \14200 , \14199 , \14025 );
xor \U$13353 ( \14201 , \14198 , \14200 );
xor \U$13354 ( \14202 , \14113 , \14129 );
xor \U$13355 ( \14203 , \14202 , \14132 );
and \U$13356 ( \14204 , \14201 , \14203 );
and \U$13357 ( \14205 , \14198 , \14200 );
or \U$13358 ( \14206 , \14204 , \14205 );
nor \U$13359 ( \14207 , \14161 , \14206 );
xor \U$13360 ( \14208 , \14159 , \14207 );
and \U$13361 ( \14209 , \14161 , \14206 );
nor \U$13362 ( \14210 , \14209 , \14207 );
xor \U$13363 ( \14211 , \14198 , \14200 );
xor \U$13364 ( \14212 , \14211 , \14203 );
xor \U$13365 ( \14213 , \14120 , \14125 );
xor \U$13366 ( \14214 , \14213 , \11852 );
nand \U$13367 ( \14215 , \13139_nG256e , \12607 );
or \U$13368 ( \14216 , \12569 , \12959_nG2600 );
nand \U$13369 ( \14217 , \14216 , \12791 );
and \U$13370 ( \14218 , \14215 , \14217 );
and \U$13371 ( \14219 , \12794 , \12959_nG2600 );
and \U$13372 ( \14220 , \13139_nG256e , \12609 );
nor \U$13373 ( \14221 , \14218 , \14219 , \14220 );
and \U$13374 ( \14222 , \14171 , \13063 );
not \U$13375 ( \14223 , \12918_nG26c6 );
and \U$13376 ( \14224 , \12886 , \14223 );
and \U$13377 ( \14225 , \12741_nG2776 , \13067 );
nor \U$13378 ( \14226 , \14222 , \14224 , \14225 );
xor \U$13379 ( \14227 , \14221 , \14226 );
and \U$13380 ( \14228 , \14227 , \11985 );
and \U$13381 ( \14229 , \14221 , \14226 );
or \U$13382 ( \14230 , \14228 , \14229 );
nand \U$13383 ( \14231 , \13523_nG23dc , \12226 );
or \U$13384 ( \14232 , \12229 , \13403_nG245a );
nand \U$13385 ( \14233 , \14232 , \12231 );
and \U$13386 ( \14234 , \14231 , \14233 );
and \U$13387 ( \14235 , \12234 , \13403_nG245a );
and \U$13388 ( \14236 , \13523_nG23dc , \12238 );
nor \U$13389 ( \14237 , \14234 , \14235 , \14236 );
xor \U$13390 ( \14238 , \14230 , \14237 );
nand \U$13391 ( \14239 , \13685_nG2388 , \12226 );
or \U$13392 ( \14240 , \12229 , \13523_nG23dc );
nand \U$13393 ( \14241 , \14240 , \12231 );
and \U$13394 ( \14242 , \14239 , \14241 );
and \U$13395 ( \14243 , \12234 , \13523_nG23dc );
and \U$13396 ( \14244 , \13685_nG2388 , \12238 );
nor \U$13397 ( \14245 , \14242 , \14243 , \14244 );
and \U$13398 ( \14246 , \13291_nG24d0 , \12553 );
or \U$13399 ( \14247 , \12258 , \13291_nG24d0 );
nand \U$13400 ( \14248 , \14247 , \12556 );
nand \U$13401 ( \14249 , \13403_nG245a , \12409 );
and \U$13402 ( \14250 , \14248 , \14249 );
and \U$13403 ( \14251 , \13403_nG245a , \12412 );
nor \U$13404 ( \14252 , \14246 , \14250 , \14251 );
xor \U$13405 ( \14253 , \14245 , \14252 );
and \U$13406 ( \14254 , \12247 , \13775_nG2272 );
nand \U$13407 ( \14255 , \13775_nG2272 , \12054 );
and \U$13408 ( \14256 , \14255 , \12058 );
nor \U$13409 ( \14257 , \14254 , \14256 );
and \U$13410 ( \14258 , \14253 , \14257 );
and \U$13411 ( \14259 , \14245 , \14252 );
or \U$13412 ( \14260 , \14258 , \14259 );
and \U$13413 ( \14261 , \14238 , \14260 );
and \U$13414 ( \14262 , \14230 , \14237 );
or \U$13415 ( \14263 , \14261 , \14262 );
nand \U$13416 ( \14264 , \14214 , \14263 );
not \U$13417 ( \14265 , \14168 );
xor \U$13418 ( \14266 , \14174 , \14184 );
not \U$13419 ( \14267 , \14266 );
or \U$13420 ( \14268 , \14265 , \14267 );
or \U$13421 ( \14269 , \14266 , \14168 );
nand \U$13422 ( \14270 , \14268 , \14269 );
or \U$13423 ( \14271 , \12268 , \13913 );
or \U$13424 ( \14272 , \13915 , \12270 );
or \U$13425 ( \14273 , \12246 , \13913 );
or \U$13426 ( \14274 , \11985 , \13775_nG2272 );
nand \U$13427 ( \14275 , \14274 , \12060 );
nand \U$13428 ( \14276 , \14273 , \14275 );
nand \U$13429 ( \14277 , \14271 , \14272 , \14276 );
and \U$13430 ( \14278 , \14270 , \14277 );
and \U$13431 ( \14279 , \14264 , \14278 );
nor \U$13432 ( \14280 , \14263 , \14214 );
nor \U$13433 ( \14281 , \14279 , \14280 );
nor \U$13434 ( \14282 , \14212 , \14281 );
xor \U$13435 ( \14283 , \14210 , \14282 );
not \U$13436 ( \14284 , \14278 );
not \U$13437 ( \14285 , \14280 );
nand \U$13438 ( \14286 , \14285 , \14264 );
not \U$13439 ( \14287 , \14286 );
or \U$13440 ( \14288 , \14284 , \14287 );
or \U$13441 ( \14289 , \14286 , \14278 );
nand \U$13442 ( \14290 , \14288 , \14289 );
xor \U$13443 ( \14291 , \14095 , \14102 );
xor \U$13444 ( \14292 , \14291 , \14110 );
xor \U$13445 ( \14293 , \14186 , \14193 );
xor \U$13446 ( \14294 , \14292 , \14293 );
not \U$13447 ( \14295 , \14294 );
xor \U$13448 ( \14296 , \14290 , \14295 );
xor \U$13449 ( \14297 , \14230 , \14237 );
xor \U$13450 ( \14298 , \14297 , \14260 );
nand \U$13451 ( \14299 , \13291_nG24d0 , \12607 );
or \U$13452 ( \14300 , \12569 , \13139_nG256e );
nand \U$13453 ( \14301 , \14300 , \12791 );
and \U$13454 ( \14302 , \14299 , \14301 );
and \U$13455 ( \14303 , \12794 , \13139_nG256e );
and \U$13456 ( \14304 , \13291_nG24d0 , \12609 );
nor \U$13457 ( \14305 , \14302 , \14303 , \14304 );
and \U$13458 ( \14306 , \14223 , \13063 );
not \U$13459 ( \14307 , \12959_nG2600 );
and \U$13460 ( \14308 , \12886 , \14307 );
and \U$13461 ( \14309 , \12918_nG26c6 , \13067 );
nor \U$13462 ( \14310 , \14306 , \14308 , \14309 );
xor \U$13463 ( \14311 , \14305 , \14310 );
and \U$13464 ( \14312 , \13403_nG245a , \12553 );
or \U$13465 ( \14313 , \12258 , \13403_nG245a );
nand \U$13466 ( \14314 , \14313 , \12556 );
nand \U$13467 ( \14315 , \13523_nG23dc , \12409 );
and \U$13468 ( \14316 , \14314 , \14315 );
and \U$13469 ( \14317 , \13523_nG23dc , \12412 );
nor \U$13470 ( \14318 , \14312 , \14316 , \14317 );
and \U$13471 ( \14319 , \14311 , \14318 );
and \U$13472 ( \14320 , \14305 , \14310 );
or \U$13473 ( \14321 , \14319 , \14320 );
xor \U$13474 ( \14322 , \14221 , \14226 );
xor \U$13475 ( \14323 , \14322 , \11985 );
and \U$13476 ( \14324 , \14321 , \14323 );
xor \U$13477 ( \14325 , \14245 , \14252 );
xor \U$13478 ( \14326 , \14325 , \14257 );
xor \U$13479 ( \14327 , \14221 , \14226 );
xor \U$13480 ( \14328 , \14327 , \11985 );
and \U$13481 ( \14329 , \14326 , \14328 );
and \U$13482 ( \14330 , \14321 , \14326 );
or \U$13483 ( \14331 , \14324 , \14329 , \14330 );
nand \U$13484 ( \14332 , \14298 , \14331 );
xor \U$13485 ( \14333 , \14270 , \14277 );
and \U$13486 ( \14334 , \14332 , \14333 );
nor \U$13487 ( \14335 , \14331 , \14298 );
nor \U$13488 ( \14336 , \14334 , \14335 );
not \U$13489 ( \14337 , \14336 );
xor \U$13490 ( \14338 , \14296 , \14337 );
not \U$13491 ( \14339 , \14332 );
nor \U$13492 ( \14340 , \14339 , \14335 );
not \U$13493 ( \14341 , \14340 );
not \U$13494 ( \14342 , \14333 );
and \U$13495 ( \14343 , \14341 , \14342 );
and \U$13496 ( \14344 , \14340 , \14333 );
nor \U$13497 ( \14345 , \14343 , \14344 );
xor \U$13498 ( \14346 , \14221 , \14226 );
xor \U$13499 ( \14347 , \14346 , \11985 );
xor \U$13500 ( \14348 , \14321 , \14326 );
xor \U$13501 ( \14349 , \14347 , \14348 );
nand \U$13502 ( \14350 , \13775_nG2272 , \12226 );
or \U$13503 ( \14351 , \12229 , \13685_nG2388 );
nand \U$13504 ( \14352 , \14351 , \12231 );
and \U$13505 ( \14353 , \14350 , \14352 );
and \U$13506 ( \14354 , \12234 , \13685_nG2388 );
and \U$13507 ( \14355 , \13775_nG2272 , \12238 );
nor \U$13508 ( \14356 , \14353 , \14354 , \14355 );
not \U$13509 ( \14357 , \13403_nG245a );
or \U$13510 ( \14358 , \12610 , \14357 );
or \U$13511 ( \14359 , \12569 , \13291_nG24d0 );
nand \U$13512 ( \14360 , \14359 , \12791 );
nand \U$13513 ( \14361 , \13403_nG245a , \12607 );
and \U$13514 ( \14362 , \14360 , \14361 );
and \U$13515 ( \14363 , \13291_nG24d0 , \12794 );
nor \U$13516 ( \14364 , \14362 , \14363 );
nand \U$13517 ( \14365 , \14358 , \14364 );
or \U$13518 ( \14366 , \13066 , \14307 );
or \U$13519 ( \14367 , \12959_nG2600 , \12888 );
or \U$13520 ( \14368 , \13139_nG256e , \12887 );
nand \U$13521 ( \14369 , \14366 , \14367 , \14368 );
or \U$13522 ( \14370 , \14365 , \14369 );
and \U$13523 ( \14371 , \12237 , \14370 );
and \U$13524 ( \14372 , \14369 , \14365 );
nor \U$13525 ( \14373 , \14371 , \14372 );
xor \U$13526 ( \14374 , \14356 , \14373 );
and \U$13527 ( \14375 , \13523_nG23dc , \12553 );
or \U$13528 ( \14376 , \12258 , \13523_nG23dc );
nand \U$13529 ( \14377 , \14376 , \12556 );
nand \U$13530 ( \14378 , \13685_nG2388 , \12409 );
and \U$13531 ( \14379 , \14377 , \14378 );
and \U$13532 ( \14380 , \13685_nG2388 , \12412 );
nor \U$13533 ( \14381 , \14375 , \14379 , \14380 );
not \U$13534 ( \14382 , \14381 );
or \U$13535 ( \14383 , \12419 , \13915 );
or \U$13536 ( \14384 , \13775_nG2272 , \12229 );
nand \U$13537 ( \14385 , \14383 , \14384 , \12231 );
nand \U$13538 ( \14386 , \14382 , \14385 );
and \U$13539 ( \14387 , \14374 , \14386 );
and \U$13540 ( \14388 , \14356 , \14373 );
or \U$13541 ( \14389 , \14387 , \14388 );
nor \U$13542 ( \14390 , \14349 , \14389 );
xor \U$13543 ( \14391 , \14345 , \14390 );
xor \U$13544 ( \14392 , \14356 , \14373 );
xor \U$13545 ( \14393 , \14392 , \14386 );
xor \U$13546 ( \14394 , \14305 , \14310 );
xor \U$13547 ( \14395 , \14394 , \14318 );
and \U$13548 ( \14396 , \14393 , \14395 );
nor \U$13549 ( \14397 , \14393 , \14395 );
nor \U$13550 ( \14398 , \14396 , \14397 );
nand \U$13551 ( \14399 , \13523_nG23dc , \12607 );
or \U$13552 ( \14400 , \12569 , \13403_nG245a );
nand \U$13553 ( \14401 , \14400 , \12791 );
and \U$13554 ( \14402 , \14399 , \14401 );
and \U$13555 ( \14403 , \12794 , \13403_nG245a );
and \U$13556 ( \14404 , \13523_nG23dc , \12609 );
nor \U$13557 ( \14405 , \14402 , \14403 , \14404 );
not \U$13558 ( \14406 , \13139_nG256e );
and \U$13559 ( \14407 , \14406 , \13063 );
not \U$13560 ( \14408 , \13291_nG24d0 );
and \U$13561 ( \14409 , \12886 , \14408 );
and \U$13562 ( \14410 , \13139_nG256e , \13067 );
nor \U$13563 ( \14411 , \14407 , \14409 , \14410 );
xor \U$13564 ( \14412 , \14405 , \14411 );
and \U$13565 ( \14413 , \13685_nG2388 , \12553 );
or \U$13566 ( \14414 , \12258 , \13685_nG2388 );
nand \U$13567 ( \14415 , \14414 , \12556 );
nand \U$13568 ( \14416 , \13775_nG2272 , \12409 );
and \U$13569 ( \14417 , \14415 , \14416 );
and \U$13570 ( \14418 , \13775_nG2272 , \12412 );
nor \U$13571 ( \14419 , \14413 , \14417 , \14418 );
and \U$13572 ( \14420 , \14412 , \14419 );
and \U$13573 ( \14421 , \14405 , \14411 );
or \U$13574 ( \14422 , \14420 , \14421 );
not \U$13575 ( \14423 , \14422 );
xnor \U$13576 ( \14424 , \14369 , \14365 );
and \U$13577 ( \14425 , \14424 , \12229 );
not \U$13578 ( \14426 , \14424 );
and \U$13579 ( \14427 , \14426 , \12237 );
nor \U$13580 ( \14428 , \14425 , \14427 );
xor \U$13581 ( \14429 , \14423 , \14428 );
not \U$13582 ( \14430 , \14381 );
not \U$13583 ( \14431 , \14385 );
or \U$13584 ( \14432 , \14430 , \14431 );
or \U$13585 ( \14433 , \14385 , \14381 );
nand \U$13586 ( \14434 , \14432 , \14433 );
and \U$13587 ( \14435 , \14429 , \14434 );
and \U$13588 ( \14436 , \14423 , \14428 );
or \U$13589 ( \14437 , \14435 , \14436 );
xor \U$13590 ( \14438 , \14398 , \14437 );
not \U$13591 ( \14439 , \13523_nG23dc );
or \U$13592 ( \14440 , \13066 , \14439 );
or \U$13593 ( \14441 , \13523_nG23dc , \12888 );
or \U$13594 ( \14442 , \13685_nG2388 , \12887 );
nand \U$13595 ( \14443 , \14440 , \14441 , \14442 );
xor \U$13596 ( \14444 , \14443 , \12570 );
and \U$13597 ( \14445 , \13913 , \13063 );
and \U$13598 ( \14446 , \12886 , \13915 );
and \U$13599 ( \14447 , \13685_nG2388 , \13067 );
nor \U$13600 ( \14448 , \14445 , \14446 , \14447 );
nand \U$13601 ( \14449 , \13775_nG2272 , \12887 );
nand \U$13602 ( \14450 , \12564 , \14449 );
nor \U$13603 ( \14451 , \14448 , \14450 );
xor \U$13604 ( \14452 , \14444 , \14451 );
not \U$13605 ( \14453 , \12794 );
or \U$13606 ( \14454 , \14453 , \13915 );
or \U$13607 ( \14455 , \13775_nG2272 , \12569 );
nand \U$13608 ( \14456 , \14454 , \14455 , \12791 );
and \U$13609 ( \14457 , \14452 , \14456 );
and \U$13610 ( \14458 , \14444 , \14451 );
or \U$13611 ( \14459 , \14457 , \14458 );
and \U$13612 ( \14460 , \14443 , \12570 );
xor \U$13613 ( \14461 , \14459 , \14460 );
nand \U$13614 ( \14462 , \13775_nG2272 , \12607 );
or \U$13615 ( \14463 , \12569 , \13685_nG2388 );
nand \U$13616 ( \14464 , \14463 , \12791 );
and \U$13617 ( \14465 , \14462 , \14464 );
and \U$13618 ( \14466 , \12794 , \13685_nG2388 );
and \U$13619 ( \14467 , \13775_nG2272 , \12609 );
nor \U$13620 ( \14468 , \14465 , \14466 , \14467 );
and \U$13621 ( \14469 , \14357 , \13063 );
and \U$13622 ( \14470 , \12886 , \14439 );
and \U$13623 ( \14471 , \13403_nG245a , \13067 );
nor \U$13624 ( \14472 , \14469 , \14470 , \14471 );
and \U$13625 ( \14473 , \14468 , \14472 );
nor \U$13626 ( \14474 , \14468 , \14472 );
nor \U$13627 ( \14475 , \14473 , \14474 );
and \U$13628 ( \14476 , \14461 , \14475 );
and \U$13629 ( \14477 , \14459 , \14460 );
or \U$13630 ( \14478 , \14476 , \14477 );
xor \U$13631 ( \14479 , \14478 , \14474 );
and \U$13632 ( \14480 , \14408 , \13063 );
and \U$13633 ( \14481 , \12886 , \14357 );
and \U$13634 ( \14482 , \13291_nG24d0 , \13067 );
nor \U$13635 ( \14483 , \14480 , \14481 , \14482 );
xor \U$13636 ( \14484 , \12258 , \14483 );
nand \U$13637 ( \14485 , \13685_nG2388 , \12607 );
or \U$13638 ( \14486 , \12569 , \13523_nG23dc );
nand \U$13639 ( \14487 , \14486 , \12791 );
and \U$13640 ( \14488 , \14485 , \14487 );
and \U$13641 ( \14489 , \12794 , \13523_nG23dc );
and \U$13642 ( \14490 , \13685_nG2388 , \12609 );
nor \U$13643 ( \14491 , \14488 , \14489 , \14490 );
xor \U$13644 ( \14492 , \14484 , \14491 );
and \U$13645 ( \14493 , \13775_nG2272 , \12553 );
and \U$13646 ( \14494 , \13915 , \12411 );
not \U$13647 ( \14495 , \12556 );
nor \U$13648 ( \14496 , \14493 , \14494 , \14495 );
and \U$13649 ( \14497 , \14492 , \14496 );
nor \U$13650 ( \14498 , \14492 , \14496 );
nor \U$13651 ( \14499 , \14497 , \14498 );
and \U$13652 ( \14500 , \14479 , \14499 );
and \U$13653 ( \14501 , \14478 , \14474 );
or \U$13654 ( \14502 , \14500 , \14501 );
xor \U$13655 ( \14503 , \14502 , \14498 );
xor \U$13656 ( \14504 , \14405 , \14411 );
xor \U$13657 ( \14505 , \14504 , \14419 );
xor \U$13658 ( \14506 , \12258 , \14483 );
and \U$13659 ( \14507 , \14506 , \14491 );
and \U$13660 ( \14508 , \12258 , \14483 );
or \U$13661 ( \14509 , \14507 , \14508 );
and \U$13662 ( \14510 , \14505 , \14509 );
nor \U$13663 ( \14511 , \14505 , \14509 );
nor \U$13664 ( \14512 , \14510 , \14511 );
and \U$13665 ( \14513 , \14503 , \14512 );
and \U$13666 ( \14514 , \14502 , \14498 );
or \U$13667 ( \14515 , \14513 , \14514 );
xor \U$13668 ( \14516 , \14515 , \14511 );
xor \U$13669 ( \14517 , \14423 , \14428 );
xor \U$13670 ( \14518 , \14517 , \14434 );
and \U$13671 ( \14519 , \14516 , \14518 );
and \U$13672 ( \14520 , \14515 , \14511 );
or \U$13673 ( \14521 , \14519 , \14520 );
and \U$13674 ( \14522 , \14438 , \14521 );
and \U$13675 ( \14523 , \14398 , \14437 );
or \U$13676 ( \14524 , \14522 , \14523 );
xor \U$13677 ( \14525 , \14524 , \14397 );
and \U$13678 ( \14526 , \14349 , \14389 );
nor \U$13679 ( \14527 , \14526 , \14390 );
and \U$13680 ( \14528 , \14525 , \14527 );
and \U$13681 ( \14529 , \14524 , \14397 );
or \U$13682 ( \14530 , \14528 , \14529 );
and \U$13683 ( \14531 , \14391 , \14530 );
and \U$13684 ( \14532 , \14345 , \14390 );
or \U$13685 ( \14533 , \14531 , \14532 );
and \U$13686 ( \14534 , \14338 , \14533 );
and \U$13687 ( \14535 , \14296 , \14337 );
or \U$13688 ( \14536 , \14534 , \14535 );
and \U$13689 ( \14537 , \14290 , \14295 );
xor \U$13690 ( \14538 , \14536 , \14537 );
and \U$13691 ( \14539 , \14212 , \14281 );
nor \U$13692 ( \14540 , \14539 , \14282 );
and \U$13693 ( \14541 , \14538 , \14540 );
and \U$13694 ( \14542 , \14536 , \14537 );
or \U$13695 ( \14543 , \14541 , \14542 );
and \U$13696 ( \14544 , \14283 , \14543 );
and \U$13697 ( \14545 , \14210 , \14282 );
or \U$13698 ( \14546 , \14544 , \14545 );
and \U$13699 ( \14547 , \14208 , \14546 );
and \U$13700 ( \14548 , \14159 , \14207 );
or \U$13701 ( \14549 , \14547 , \14548 );
or \U$13702 ( \14550 , \14148 , \14155 );
nand \U$13703 ( \14551 , \14550 , \14146 );
xor \U$13704 ( \14552 , \13999 , \14077 );
xor \U$13705 ( \14553 , \14552 , \14080 );
nand \U$13706 ( \14554 , \14551 , \14553 );
and \U$13707 ( \14555 , \14549 , \14554 );
nor \U$13708 ( \14556 , \14553 , \14551 );
nor \U$13709 ( \14557 , \14555 , \14556 );
xor \U$13710 ( \14558 , \13977 , \13979 );
xor \U$13711 ( \14559 , \14558 , \13982 );
and \U$13712 ( \14560 , \14557 , \14559 );
and \U$13713 ( \14561 , \14083 , \14557 );
or \U$13714 ( \14562 , \14086 , \14560 , \14561 );
xor \U$13715 ( \14563 , \13900 , \13905 );
xor \U$13716 ( \14564 , \14563 , \13908 );
and \U$13717 ( \14565 , \14562 , \14564 );
and \U$13718 ( \14566 , \13985 , \14562 );
or \U$13719 ( \14567 , \13988 , \14565 , \14566 );
and \U$13720 ( \14568 , \13912 , \14567 );
and \U$13721 ( \14569 , \13831 , \13911 );
or \U$13722 ( \14570 , \14568 , \14569 );
not \U$13723 ( \14571 , \14570 );
and \U$13724 ( \14572 , \13829 , \14571 );
and \U$13725 ( \14573 , \13818 , \13828 );
or \U$13726 ( \14574 , \14572 , \14573 );
and \U$13727 ( \14575 , \13816 , \14574 );
and \U$13728 ( \14576 , \13644 , \13815 );
or \U$13729 ( \14577 , \14575 , \14576 );
and \U$13730 ( \14578 , \13642 , \14577 );
and \U$13731 ( \14579 , \13639 , \13641 );
or \U$13732 ( \14580 , \14578 , \14579 );
and \U$13733 ( \14581 , \13554 , \14580 );
and \U$13734 ( \14582 , \13375 , \13553 );
or \U$13735 ( \14583 , \14581 , \14582 );
and \U$13736 ( \14584 , \13373 , \14583 );
and \U$13737 ( \14585 , \13349 , \13372 );
or \U$13738 ( \14586 , \14584 , \14585 );
and \U$13739 ( \14587 , \13359 , \13368 );
nor \U$13740 ( \14588 , \14587 , \13361 );
xor \U$13741 ( \14589 , \13019 , \13104 );
xor \U$13742 ( \14590 , \14589 , \13107 );
nand \U$13743 ( \14591 , \14588 , \14590 );
and \U$13744 ( \14592 , \14586 , \14591 );
nor \U$13745 ( \14593 , \14590 , \14588 );
nor \U$13746 ( \14594 , \14592 , \14593 );
and \U$13747 ( \14595 , \13111 , \14594 );
and \U$13748 ( \14596 , \13009 , \13110 );
or \U$13749 ( \14597 , \14595 , \14596 );
not \U$13750 ( \14598 , \14597 );
and \U$13751 ( \14599 , \13002 , \14598 );
and \U$13752 ( \14600 , \12845 , \13001 );
or \U$13753 ( \14601 , \14599 , \14600 );
and \U$13754 ( \14602 , \12841 , \14601 );
and \U$13755 ( \14603 , \12704 , \12840 );
or \U$13756 ( \14604 , \14602 , \14603 );
and \U$13757 ( \14605 , \12702 , \14604 );
and \U$13758 ( \14606 , \12697 , \12701 );
or \U$13759 ( \14607 , \14605 , \14606 );
and \U$13760 ( \14608 , \12595 , \14607 );
and \U$13761 ( \14609 , \12489 , \12594 );
or \U$13762 ( \14610 , \14608 , \14609 );
and \U$13763 ( \14611 , \12487 , \14610 );
and \U$13764 ( \14612 , \12401 , \12486 );
or \U$13765 ( \14613 , \14611 , \14612 );
and \U$13766 ( \14614 , \12399 , \14613 );
and \U$13767 ( \14615 , \12378 , \12398 );
or \U$13768 ( \14616 , \14614 , \14615 );
not \U$13769 ( \14617 , \12104 );
not \U$13770 ( \14618 , \12108 );
nand \U$13771 ( \14619 , \14618 , \12110 );
not \U$13772 ( \14620 , \14619 );
or \U$13773 ( \14621 , \14617 , \14620 );
or \U$13774 ( \14622 , \14619 , \12104 );
nand \U$13775 ( \14623 , \14621 , \14622 );
or \U$13776 ( \14624 , \12388 , \12394 );
nand \U$13777 ( \14625 , \14624 , \12386 );
nand \U$13778 ( \14626 , \14623 , \14625 );
and \U$13779 ( \14627 , \14616 , \14626 );
nor \U$13780 ( \14628 , \14625 , \14623 );
nor \U$13781 ( \14629 , \14627 , \14628 );
nor \U$13782 ( \14630 , \12116 , \14629 );
nor \U$13783 ( \14631 , \12113 , \14630 );
not \U$13784 ( \14632 , \14631 );
or \U$13785 ( \14633 , \12004 , \14632 );
or \U$13786 ( \14634 , \14631 , \12003 );
nand \U$13787 ( \14635 , \14633 , \14634 );
buf \U$13788 ( \14636 , \11367 );
buf \U$13789 ( \14637 , \7962 );
_DC g7bc ( \14638_nG7bc , \14636 , \14637 );
not \U$13790 ( \14639 , \14638_nG7bc );
buf \U$13791 ( \14640 , \7958 );
buf \U$13792 ( \14641 , \7962 );
_DC g7b9 ( \14642_nG7b9 , \14640 , \14641 );
and \U$13793 ( \14643 , \14639 , \14642_nG7b9 );
buf \U$13794 ( \14644 , \8361 );
_DC g91b ( \14645_nG91b , \14644 , \14641 );
not \U$13795 ( \14646 , \14645_nG91b );
not \U$13796 ( \14647 , \14646 );
buf \U$13797 ( \14648 , \11687 );
_DC g91d ( \14649_nG91d , \14648 , \14637 );
not \U$13798 ( \14650 , \14649_nG91d );
and \U$13799 ( \14651 , \14647 , \14650 );
buf \U$13800 ( \14652 , \8392 );
_DC g93a ( \14653_nG93a , \14652 , \14641 );
nor \U$13801 ( \14654 , \14651 , \14653_nG93a );
buf \U$13802 ( \14655 , \11716 );
_DC g93c ( \14656_nG93c , \14655 , \14637 );
and \U$13803 ( \14657 , \14654 , \14656_nG93c );
and \U$13804 ( \14658 , \14649_nG91d , \14646 );
nor \U$13805 ( \14659 , \14657 , \14658 );
buf \U$13806 ( \14660 , \11658 );
_DC g8fe ( \14661_nG8fe , \14660 , \14637 );
not \U$13807 ( \14662 , \14661_nG8fe );
and \U$13808 ( \14663 , \14659 , \14662 );
buf \U$13809 ( \14664 , \8330 );
_DC g8fc ( \14665_nG8fc , \14664 , \14641 );
or \U$13810 ( \14666 , \14663 , \14665_nG8fc );
or \U$13811 ( \14667 , \14662 , \14659 );
nand \U$13812 ( \14668 , \14666 , \14667 );
buf \U$13813 ( \14669 , \11629 );
_DC g8df ( \14670_nG8df , \14669 , \14637 );
not \U$13814 ( \14671 , \14670_nG8df );
buf \U$13815 ( \14672 , \8298 );
_DC g8dd ( \14673_nG8dd , \14672 , \14641 );
nand \U$13816 ( \14674 , \14671 , \14673_nG8dd );
and \U$13817 ( \14675 , \14668 , \14674 );
not \U$13818 ( \14676 , \14673_nG8dd );
and \U$13819 ( \14677 , \14670_nG8df , \14676 );
nor \U$13820 ( \14678 , \14675 , \14677 );
buf \U$13821 ( \14679 , \8260 );
_DC g8bc ( \14680_nG8bc , \14679 , \14641 );
or \U$13822 ( \14681 , \14678 , \14680_nG8bc );
not \U$13823 ( \14682 , \14680_nG8bc );
not \U$13824 ( \14683 , \14678 );
or \U$13825 ( \14684 , \14682 , \14683 );
buf \U$13826 ( \14685 , \11600 );
_DC g8be ( \14686_nG8be , \14685 , \14637 );
nand \U$13827 ( \14687 , \14684 , \14686_nG8be );
nand \U$13828 ( \14688 , \14681 , \14687 );
buf \U$13829 ( \14689 , \11571 );
_DC g89f ( \14690_nG89f , \14689 , \14637 );
and \U$13830 ( \14691 , \14688 , \14690_nG89f );
not \U$13831 ( \14692 , \14688 );
not \U$13832 ( \14693 , \14690_nG89f );
and \U$13833 ( \14694 , \14692 , \14693 );
buf \U$13834 ( \14695 , \8224 );
_DC g89d ( \14696_nG89d , \14695 , \14641 );
nor \U$13835 ( \14697 , \14694 , \14696_nG89d );
nor \U$13836 ( \14698 , \14691 , \14697 );
buf \U$13837 ( \14699 , \8186 );
_DC g87c ( \14700_nG87c , \14699 , \14641 );
or \U$13838 ( \14701 , \14698 , \14700_nG87c );
not \U$13839 ( \14702 , \14700_nG87c );
not \U$13840 ( \14703 , \14698 );
or \U$13841 ( \14704 , \14702 , \14703 );
buf \U$13842 ( \14705 , \11542 );
_DC g87e ( \14706_nG87e , \14705 , \14637 );
nand \U$13843 ( \14707 , \14704 , \14706_nG87e );
nand \U$13844 ( \14708 , \14701 , \14707 );
buf \U$13845 ( \14709 , \11513 );
_DC g85d ( \14710_nG85d , \14709 , \14637 );
and \U$13846 ( \14711 , \14708 , \14710_nG85d );
not \U$13847 ( \14712 , \14708 );
not \U$13848 ( \14713 , \14710_nG85d );
and \U$13849 ( \14714 , \14712 , \14713 );
buf \U$13850 ( \14715 , \8148 );
_DC g85b ( \14716_nG85b , \14715 , \14641 );
nor \U$13851 ( \14717 , \14714 , \14716_nG85b );
nor \U$13852 ( \14718 , \14711 , \14717 );
buf \U$13853 ( \14719 , \11484 );
_DC g83c ( \14720_nG83c , \14719 , \14637 );
not \U$13854 ( \14721 , \14720_nG83c );
buf \U$13855 ( \14722 , \8110 );
_DC g83a ( \14723_nG83a , \14722 , \14641 );
and \U$13856 ( \14724 , \14721 , \14723_nG83a );
or \U$13857 ( \14725 , \14718 , \14724 );
or \U$13858 ( \14726 , \14723_nG83a , \14721 );
nand \U$13859 ( \14727 , \14725 , \14726 );
buf \U$13860 ( \14728 , \11455 );
_DC g81d ( \14729_nG81d , \14728 , \14637 );
and \U$13861 ( \14730 , \14727 , \14729_nG81d );
not \U$13862 ( \14731 , \14727 );
not \U$13863 ( \14732 , \14729_nG81d );
and \U$13864 ( \14733 , \14731 , \14732 );
buf \U$13865 ( \14734 , \8074 );
_DC g81b ( \14735_nG81b , \14734 , \14641 );
nor \U$13866 ( \14736 , \14733 , \14735_nG81b );
nor \U$13867 ( \14737 , \14730 , \14736 );
buf \U$13868 ( \14738 , \8036 );
_DC g7fa ( \14739_nG7fa , \14738 , \14641 );
or \U$13869 ( \14740 , \14737 , \14739_nG7fa );
not \U$13870 ( \14741 , \14739_nG7fa );
not \U$13871 ( \14742 , \14737 );
or \U$13872 ( \14743 , \14741 , \14742 );
buf \U$13873 ( \14744 , \11426 );
_DC g7fc ( \14745_nG7fc , \14744 , \14637 );
nand \U$13874 ( \14746 , \14743 , \14745_nG7fc );
nand \U$13875 ( \14747 , \14740 , \14746 );
buf \U$13876 ( \14748 , \11397 );
_DC g7db ( \14749_nG7db , \14748 , \14637 );
and \U$13877 ( \14750 , \14747 , \14749_nG7db );
not \U$13878 ( \14751 , \14747 );
not \U$13879 ( \14752 , \14749_nG7db );
and \U$13880 ( \14753 , \14751 , \14752 );
buf \U$13881 ( \14754 , \7998 );
_DC g7d9 ( \14755_nG7d9 , \14754 , \14641 );
nor \U$13882 ( \14756 , \14753 , \14755_nG7d9 );
nor \U$13883 ( \14757 , \14750 , \14756 );
nor \U$13884 ( \14758 , \14643 , \14757 );
nor \U$13885 ( \14759 , \14639 , \14642_nG7b9 );
or \U$13886 ( \14760 , \14758 , \14759 );
not \U$13887 ( \14761 , RIb55b8e0_591);
nor \U$13888 ( \14762 , \7870 , RIb55b778_588);
nand \U$13889 ( \14763 , RIb55bac0_595, \14762 );
not \U$13890 ( \14764 , \14763 );
nand \U$13891 ( \14765 , \14764 , RIb55ba48_594);
nor \U$13892 ( \14766 , \14765 , \8116 );
nand \U$13893 ( \14767 , RIb55b958_592, \14766 );
nor \U$13894 ( \14768 , \14761 , \14767 );
nand \U$13895 ( \14769 , RIb55b868_590, \14768 );
not \U$13896 ( \14770 , \14769 );
nand \U$13897 ( \14771 , RIb55b7f0_589, \14770 );
not \U$13898 ( \14772 , \14771 );
not \U$13899 ( \14773 , RIb55c3a8_614);
and \U$13900 ( \14774 , \14772 , \14773 );
and \U$13901 ( \14775 , \14771 , RIb55c3a8_614);
nor \U$13902 ( \14776 , \14774 , \14775 );
buf \U$13903 ( \14777 , \11367 );
buf \U$13904 ( \14778 , \7962 );
_DC g63b ( \14779_nG63b , \14777 , \14778 );
nor \U$13905 ( \14780 , \14776 , \14779_nG63b );
and \U$13906 ( \14781 , \14776 , \14779_nG63b );
or \U$13907 ( \14782 , \14770 , RIb55b7f0_589);
nand \U$13908 ( \14783 , \14782 , \14771 );
not \U$13909 ( \14784 , \14783 );
buf \U$13910 ( \14785 , \11397 );
_DC g658 ( \14786_nG658 , \14785 , \14778 );
not \U$13911 ( \14787 , \14786_nG658 );
and \U$13912 ( \14788 , \14784 , \14787 );
and \U$13913 ( \14789 , \14786_nG658 , \14783 );
or \U$13914 ( \14790 , \14768 , RIb55b868_590);
nand \U$13915 ( \14791 , \14790 , \14769 );
buf \U$13916 ( \14792 , \11455 );
_DC g692 ( \14793_nG692 , \14792 , \14778 );
not \U$13917 ( \14794 , \14793_nG692 );
not \U$13918 ( \14795 , \14767 );
not \U$13919 ( \14796 , RIb55b8e0_591);
and \U$13920 ( \14797 , \14795 , \14796 );
and \U$13921 ( \14798 , \14767 , RIb55b8e0_591);
nor \U$13922 ( \14799 , \14797 , \14798 );
not \U$13923 ( \14800 , \14799 );
or \U$13924 ( \14801 , \14794 , \14800 );
buf \U$13925 ( \14802 , \11513 );
_DC g6cc ( \14803_nG6cc , \14802 , \14778 );
buf \U$13926 ( \14804 , \11542 );
_DC g6e9 ( \14805_nG6e9 , \14804 , \14778 );
not \U$13927 ( \14806 , \14805_nG6e9 );
not \U$13928 ( \14807 , \14763 );
not \U$13929 ( \14808 , RIb55ba48_594);
and \U$13930 ( \14809 , \14807 , \14808 );
and \U$13931 ( \14810 , \14763 , RIb55ba48_594);
nor \U$13932 ( \14811 , \14809 , \14810 );
not \U$13933 ( \14812 , \14811 );
or \U$13934 ( \14813 , \14806 , \14812 );
or \U$13935 ( \14814 , \14762 , RIb55bac0_595);
nand \U$13936 ( \14815 , \14814 , \14763 );
buf \U$13937 ( \14816 , \11600 );
_DC g723 ( \14817_nG723 , \14816 , \14778 );
not \U$13938 ( \14818 , \14817_nG723 );
not \U$13939 ( \14819 , \7868 );
not \U$13940 ( \14820 , RIb55b778_588);
and \U$13941 ( \14821 , \14819 , \14820 );
nor \U$13942 ( \14822 , \14821 , RIb55bb38_596);
or \U$13943 ( \14823 , \14762 , \14822 );
not \U$13944 ( \14824 , \14823 );
or \U$13945 ( \14825 , \14818 , \14824 );
or \U$13946 ( \14826 , \14823 , \14817_nG723 );
buf \U$13947 ( \14827 , \11629 );
_DC g740 ( \14828_nG740 , \14827 , \14778 );
not \U$13948 ( \14829 , \7866 );
nand \U$13949 ( \14830 , \14829 , \7463 );
not \U$13950 ( \14831 , \14830 );
not \U$13951 ( \14832 , RIb55bbb0_597);
and \U$13952 ( \14833 , \14831 , \14832 );
and \U$13953 ( \14834 , \14830 , RIb55bbb0_597);
nor \U$13954 ( \14835 , \14833 , \14834 );
or \U$13955 ( \14836 , \14828_nG740 , \14835 );
and \U$13956 ( \14837 , \14835 , \14828_nG740 );
buf \U$13957 ( \14838 , \11658 );
_DC g75d ( \14839_nG75d , \14838 , \14778 );
nand \U$13958 ( \14840 , RIb55bca0_599, \7463 );
not \U$13959 ( \14841 , \14840 );
not \U$13960 ( \14842 , RIb55bc28_598);
and \U$13961 ( \14843 , \14841 , \14842 );
and \U$13962 ( \14844 , \14840 , RIb55bc28_598);
nor \U$13963 ( \14845 , \14843 , \14844 );
and \U$13964 ( \14846 , \14839_nG75d , \14845 );
nor \U$13965 ( \14847 , \14837 , \14846 );
or \U$13966 ( \14848 , \14845 , \14839_nG75d );
buf \U$13967 ( \14849 , \11687 );
_DC g77a ( \14850_nG77a , \14849 , \14778 );
or \U$13968 ( \14851 , \7463 , RIb55bca0_599);
nand \U$13969 ( \14852 , \14851 , \14840 );
or \U$13970 ( \14853 , \14850_nG77a , \14852 );
and \U$13971 ( \14854 , \14852 , \14850_nG77a );
buf \U$13972 ( \14855 , \11716 );
_DC g797 ( \14856_nG797 , \14855 , \14778 );
and \U$13973 ( \14857 , \14856_nG797 , \8395 );
nor \U$13974 ( \14858 , \14854 , \14857 );
not \U$13975 ( \14859 , \14858 );
nand \U$13976 ( \14860 , \14848 , \14853 , \14859 );
nand \U$13977 ( \14861 , \14847 , \14860 );
nand \U$13978 ( \14862 , \14826 , \14836 , \14861 );
nand \U$13979 ( \14863 , \14825 , \14862 );
buf \U$13980 ( \14864 , \11571 );
_DC g706 ( \14865_nG706 , \14864 , \14778 );
or \U$13981 ( \14866 , \14863 , \14865_nG706 );
and \U$13982 ( \14867 , \14815 , \14866 );
and \U$13983 ( \14868 , \14865_nG706 , \14863 );
nor \U$13984 ( \14869 , \14867 , \14868 );
nor \U$13985 ( \14870 , \14811 , \14805_nG6e9 );
or \U$13986 ( \14871 , \14869 , \14870 );
nand \U$13987 ( \14872 , \14813 , \14871 );
and \U$13988 ( \14873 , \14803_nG6cc , \14872 );
buf \U$13989 ( \14874 , \11484 );
_DC g6af ( \14875_nG6af , \14874 , \14778 );
or \U$13990 ( \14876 , \14766 , RIb55b958_592);
nand \U$13991 ( \14877 , \14876 , \14767 );
and \U$13992 ( \14878 , \14875_nG6af , \14877 );
and \U$13993 ( \14879 , \14765 , RIb55b9d0_593);
or \U$13994 ( \14880 , \14872 , \14803_nG6cc );
or \U$13995 ( \14881 , RIb55b9d0_593, \14765 );
nand \U$13996 ( \14882 , \14880 , \14881 );
nor \U$13997 ( \14883 , \14879 , \14882 );
nor \U$13998 ( \14884 , \14873 , \14878 , \14883 );
or \U$13999 ( \14885 , \14799 , \14793_nG692 );
or \U$14000 ( \14886 , \14875_nG6af , \14877 );
nand \U$14001 ( \14887 , \14885 , \14886 );
or \U$14002 ( \14888 , \14884 , \14887 );
nand \U$14003 ( \14889 , \14801 , \14888 );
or \U$14004 ( \14890 , \14791 , \14889 );
buf \U$14005 ( \14891 , \11426 );
_DC g675 ( \14892_nG675 , \14891 , \14778 );
and \U$14006 ( \14893 , \14890 , \14892_nG675 );
and \U$14007 ( \14894 , \14889 , \14791 );
nor \U$14008 ( \14895 , \14789 , \14893 , \14894 );
nor \U$14009 ( \14896 , \14788 , \14895 );
nor \U$14010 ( \14897 , \14781 , \14896 );
or \U$14011 ( \14898 , \14780 , \14897 );
nand \U$14012 ( \14899 , \14760 , \14898 );
nor \U$14013 ( \14900 , \14899 , \11339 );
_HMUX g3b42_GF_PartitionCandidate ( \14901_nG3b42 , \11336 , \14635 , \14900 );
buf \U$14014 ( \14902 , \14901_nG3b42 );
not \U$14015 ( \14903 , \11331 );
nand \U$14016 ( \14904 , \14903 , \11329 );
not \U$14017 ( \14905 , \14904 );
not \U$14018 ( \14906 , \11321 );
or \U$14019 ( \14907 , \14905 , \14906 );
or \U$14020 ( \14908 , \11321 , \14904 );
nand \U$14021 ( \14909 , \14907 , \14908 );
not \U$14022 ( \14910 , \12111 );
not \U$14023 ( \14911 , \14629 );
not \U$14024 ( \14912 , \12112 );
and \U$14025 ( \14913 , \14911 , \14912 );
and \U$14026 ( \14914 , \14629 , \12112 );
nor \U$14027 ( \14915 , \14913 , \14914 );
not \U$14028 ( \14916 , \14915 );
or \U$14029 ( \14917 , \14910 , \14916 );
or \U$14030 ( \14918 , \14915 , \12111 );
nand \U$14031 ( \14919 , \14917 , \14918 );
_HMUX g3b06_GF_PartitionCandidate ( \14920_nG3b06 , \14909 , \14919 , \14900 );
buf \U$14032 ( \14921 , \14920_nG3b06 );
xor \U$14033 ( \14922 , \8808 , \8985 );
xor \U$14034 ( \14923 , \14922 , \11318 );
not \U$14035 ( \14924 , \14628 );
nand \U$14036 ( \14925 , \14924 , \14626 );
not \U$14037 ( \14926 , \14925 );
not \U$14038 ( \14927 , \14616 );
or \U$14039 ( \14928 , \14926 , \14927 );
or \U$14040 ( \14929 , \14616 , \14925 );
nand \U$14041 ( \14930 , \14928 , \14929 );
_HMUX g3ac7_GF_PartitionCandidate ( \14931_nG3ac7 , \14923 , \14930 , \14900 );
buf \U$14042 ( \14932 , \14931_nG3ac7 );
xor \U$14043 ( \14933 , \9094 , \9101 );
xor \U$14044 ( \14934 , \14933 , \11314 );
not \U$14045 ( \14935 , \14934 );
xor \U$14046 ( \14936 , \12378 , \12398 );
xor \U$14047 ( \14937 , \14936 , \14613 );
_HMUX g3a68_GF_PartitionCandidate ( \14938_nG3a68 , \14935 , \14937 , \14900 );
buf \U$14048 ( \14939 , \14938_nG3a68 );
not \U$14049 ( \14940 , \11313 );
nand \U$14050 ( \14941 , \14940 , \11311 );
not \U$14051 ( \14942 , \14941 );
not \U$14052 ( \14943 , \11304 );
or \U$14053 ( \14944 , \14942 , \14943 );
or \U$14054 ( \14945 , \11304 , \14941 );
nand \U$14055 ( \14946 , \14944 , \14945 );
xor \U$14056 ( \14947 , \12401 , \12486 );
xor \U$14057 ( \14948 , \14947 , \14610 );
_HMUX g39fa_GF_PartitionCandidate ( \14949_nG39fa , \14946 , \14948 , \14900 );
buf \U$14058 ( \14950 , \14949_nG39fa );
xor \U$14059 ( \14951 , \9200 , \9312 );
xor \U$14060 ( \14952 , \14951 , \11301 );
xor \U$14061 ( \14953 , \12489 , \12594 );
xor \U$14062 ( \14954 , \14953 , \14607 );
_HMUX g397d_GF_PartitionCandidate ( \14955_nG397d , \14952 , \14954 , \14900 );
buf \U$14063 ( \14956 , \14955_nG397d );
xor \U$14064 ( \14957 , \9421 , \9425 );
xor \U$14065 ( \14958 , \14957 , \11298 );
xor \U$14066 ( \14959 , \12697 , \12701 );
xor \U$14067 ( \14960 , \14959 , \14604 );
_HMUX g38f4_GF_PartitionCandidate ( \14961_nG38f4 , \14958 , \14960 , \14900 );
buf \U$14068 ( \14962 , \14961_nG38f4 );
xor \U$14069 ( \14963 , \9428 , \9567 );
xor \U$14070 ( \14964 , \14963 , \11295 );
xor \U$14071 ( \14965 , \12704 , \12840 );
xor \U$14072 ( \14966 , \14965 , \14601 );
_HMUX g386b_GF_PartitionCandidate ( \14967_nG386b , \14964 , \14966 , \14900 );
buf \U$14073 ( \14968 , \14967_nG386b );
not \U$14074 ( \14969 , \11293 );
nand \U$14075 ( \14970 , \14969 , \11291 );
not \U$14076 ( \14971 , \14970 );
not \U$14077 ( \14972 , \11282 );
or \U$14078 ( \14973 , \14971 , \14972 );
or \U$14079 ( \14974 , \11282 , \14970 );
nand \U$14080 ( \14975 , \14973 , \14974 );
xor \U$14081 ( \14976 , \12845 , \13001 );
xor \U$14082 ( \14977 , \14976 , \14598 );
_HMUX g37d3_GF_PartitionCandidate ( \14978_nG37d3 , \14975 , \14977 , \14900 );
buf \U$14083 ( \14979 , \14978_nG37d3 );
xor \U$14084 ( \14980 , \9737 , \9848 );
xor \U$14085 ( \14981 , \14980 , \11279 );
xor \U$14086 ( \14982 , \13009 , \13110 );
xor \U$14087 ( \14983 , \14982 , \14594 );
not \U$14088 ( \14984 , \14983 );
_HMUX g3717_GF_PartitionCandidate ( \14985_nG3717 , \14981 , \14984 , \14900 );
buf \U$14089 ( \14986 , \14985_nG3717 );
xor \U$14090 ( \14987 , \10012 , \10014 );
xor \U$14091 ( \14988 , \14987 , \11276 );
not \U$14092 ( \14989 , \14593 );
nand \U$14093 ( \14990 , \14989 , \14591 );
not \U$14094 ( \14991 , \14990 );
not \U$14095 ( \14992 , \14586 );
or \U$14096 ( \14993 , \14991 , \14992 );
or \U$14097 ( \14994 , \14586 , \14990 );
nand \U$14098 ( \14995 , \14993 , \14994 );
_HMUX g365e_GF_PartitionCandidate ( \14996_nG365e , \14988 , \14995 , \14900 );
buf \U$14099 ( \14997 , \14996_nG365e );
xor \U$14100 ( \14998 , \10089 , \10091 );
xor \U$14101 ( \14999 , \14998 , \11273 );
xor \U$14102 ( \15000 , \13349 , \13372 );
xor \U$14103 ( \15001 , \15000 , \14583 );
_HMUX g358f_GF_PartitionCandidate ( \15002_nG358f , \14999 , \15001 , \14900 );
buf \U$14104 ( \15003 , \15002_nG358f );
xor \U$14105 ( \15004 , \10094 , \10263 );
xor \U$14106 ( \15005 , \15004 , \11270 );
xor \U$14107 ( \15006 , \13375 , \13553 );
xor \U$14108 ( \15007 , \15006 , \14580 );
_HMUX g34be_GF_PartitionCandidate ( \15008_nG34be , \15005 , \15007 , \14900 );
buf \U$14109 ( \15009 , \15008_nG34be );
xor \U$14110 ( \15010 , \10266 , \10352 );
xor \U$14111 ( \15011 , \15010 , \11267 );
xor \U$14112 ( \15012 , \13639 , \13641 );
xor \U$14113 ( \15013 , \15012 , \14577 );
_HMUX g33ea_GF_PartitionCandidate ( \15014_nG33ea , \15011 , \15013 , \14900 );
buf \U$14114 ( \15015 , \15014_nG33ea );
xor \U$14115 ( \15016 , \10357 , \10526 );
xor \U$14116 ( \15017 , \15016 , \11264 );
xor \U$14117 ( \15018 , \13644 , \13815 );
xor \U$14118 ( \15019 , \15018 , \14574 );
_HMUX g3309_GF_PartitionCandidate ( \15020_nG3309 , \15017 , \15019 , \14900 );
buf \U$14119 ( \15021 , \15020_nG3309 );
xor \U$14120 ( \15022 , \10529 , \10534 );
xor \U$14121 ( \15023 , \15022 , \11261 );
xor \U$14122 ( \15024 , \13818 , \13828 );
xor \U$14123 ( \15025 , \15024 , \14571 );
_HMUX g3207_GF_PartitionCandidate ( \15026_nG3207 , \15023 , \15025 , \14900 );
buf \U$14124 ( \15027 , \15026_nG3207 );
xor \U$14125 ( \15028 , \10537 , \10619 );
xor \U$14126 ( \15029 , \15028 , \11258 );
xor \U$14127 ( \15030 , \13831 , \13911 );
xor \U$14128 ( \15031 , \15030 , \14567 );
not \U$14129 ( \15032 , \15031 );
_HMUX g30ef_GF_PartitionCandidate ( \15033_nG30ef , \15029 , \15032 , \14900 );
buf \U$14130 ( \15034 , \15033_nG30ef );
xor \U$14131 ( \15035 , \10607 , \10612 );
xor \U$14132 ( \15036 , \15035 , \10615 );
xor \U$14133 ( \15037 , \10691 , \11252 );
xor \U$14134 ( \15038 , \15036 , \15037 );
not \U$14135 ( \15039 , \15038 );
xor \U$14136 ( \15040 , \13900 , \13905 );
xor \U$14137 ( \15041 , \15040 , \13908 );
xor \U$14138 ( \15042 , \13985 , \14562 );
xor \U$14139 ( \15043 , \15041 , \15042 );
not \U$14140 ( \15044 , \15043 );
_HMUX g2fe8_GF_PartitionCandidate ( \15045_nG2fe8 , \15039 , \15044 , \14900 );
buf \U$14141 ( \15046 , \15045_nG2fe8 );
xor \U$14142 ( \15047 , \10683 , \10685 );
xor \U$14143 ( \15048 , \15047 , \10688 );
xor \U$14144 ( \15049 , \10784 , \11247 );
xor \U$14145 ( \15050 , \15048 , \15049 );
not \U$14146 ( \15051 , \15050 );
xor \U$14147 ( \15052 , \13977 , \13979 );
xor \U$14148 ( \15053 , \15052 , \13982 );
xor \U$14149 ( \15054 , \14083 , \14557 );
xor \U$14150 ( \15055 , \15053 , \15054 );
not \U$14151 ( \15056 , \15055 );
_HMUX g2ec6_GF_PartitionCandidate ( \15057_nG2ec6 , \15051 , \15056 , \14900 );
buf \U$14152 ( \15058 , \15057_nG2ec6 );
not \U$14153 ( \15059 , \11246 );
nand \U$14154 ( \15060 , \15059 , \11244 );
not \U$14155 ( \15061 , \15060 );
not \U$14156 ( \15062 , \11237 );
or \U$14157 ( \15063 , \15061 , \15062 );
or \U$14158 ( \15064 , \11237 , \15060 );
nand \U$14159 ( \15065 , \15063 , \15064 );
not \U$14160 ( \15066 , \14556 );
nand \U$14161 ( \15067 , \15066 , \14554 );
not \U$14162 ( \15068 , \15067 );
not \U$14163 ( \15069 , \14549 );
or \U$14164 ( \15070 , \15068 , \15069 );
or \U$14165 ( \15071 , \14549 , \15067 );
nand \U$14166 ( \15072 , \15070 , \15071 );
_HMUX g2ddc_GF_PartitionCandidate ( \15073_nG2ddc , \15065 , \15072 , \14900 );
buf \U$14167 ( \15074 , \15073_nG2ddc );
xor \U$14168 ( \15075 , \10850 , \10897 );
xor \U$14169 ( \15076 , \15075 , \11234 );
xor \U$14170 ( \15077 , \14159 , \14207 );
xor \U$14171 ( \15078 , \15077 , \14546 );
_HMUX g2cdc_GF_PartitionCandidate ( \15079_nG2cdc , \15076 , \15078 , \14900 );
buf \U$14172 ( \15080 , \15079_nG2cdc );
xor \U$14173 ( \15081 , \10900 , \10973 );
xor \U$14174 ( \15082 , \15081 , \11231 );
xor \U$14175 ( \15083 , \14210 , \14282 );
xor \U$14176 ( \15084 , \15083 , \14543 );
_HMUX g2bd8_GF_PartitionCandidate ( \15085_nG2bd8 , \15082 , \15084 , \14900 );
buf \U$14177 ( \15086 , \15085_nG2bd8 );
xor \U$14178 ( \15087 , \11224 , \11225 );
xor \U$14179 ( \15088 , \15087 , \11228 );
xor \U$14180 ( \15089 , \14536 , \14537 );
xor \U$14181 ( \15090 , \15089 , \14540 );
_HMUX g2acc_GF_PartitionCandidate ( \15091_nG2acc , \15088 , \15090 , \14900 );
buf \U$14182 ( \15092 , \15091_nG2acc );
xor \U$14183 ( \15093 , \10987 , \11027 );
xor \U$14184 ( \15094 , \15093 , \11221 );
xor \U$14185 ( \15095 , \14296 , \14337 );
xor \U$14186 ( \15096 , \15095 , \14533 );
_HMUX g29ee_GF_PartitionCandidate ( \15097_nG29ee , \15094 , \15096 , \14900 );
buf \U$14187 ( \15098 , \15097_nG29ee );
xor \U$14188 ( \15099 , \11035 , \11078 );
xor \U$14189 ( \15100 , \15099 , \11218 );
xor \U$14190 ( \15101 , \14345 , \14390 );
xor \U$14191 ( \15102 , \15101 , \14530 );
_HMUX g28ee_GF_PartitionCandidate ( \15103_nG28ee , \15100 , \15102 , \14900 );
buf \U$14192 ( \15104 , \15103_nG28ee );
xor \U$14193 ( \15105 , \11212 , \11085 );
xor \U$14194 ( \15106 , \15105 , \11215 );
xor \U$14195 ( \15107 , \14524 , \14397 );
xor \U$14196 ( \15108 , \15107 , \14527 );
_HMUX g2813_GF_PartitionCandidate ( \15109_nG2813 , \15106 , \15108 , \14900 );
buf \U$14197 ( \15110 , \15109_nG2813 );
xor \U$14198 ( \15111 , \11086 , \11120 );
xor \U$14199 ( \15112 , \15111 , \11209 );
xor \U$14200 ( \15113 , \14398 , \14437 );
xor \U$14201 ( \15114 , \15113 , \14521 );
_HMUX g2739_GF_PartitionCandidate ( \15115_nG2739 , \15112 , \15114 , \14900 );
buf \U$14202 ( \15116 , \15115_nG2739 );
endmodule

