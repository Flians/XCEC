//
// Conformal-LEC Version 20.10-d214 (03-Sep-2020)
//
module top(RI9148f90_243,RI91589e0_777,RI9158968_776,RI91588f0_775,RI9158878_774,RI9158800_773,RI9158788_772,RI9158710_771,RI9158698_770,
        RI9158620_769,RI9148810_227,RI9148090_211,RI9147910_195,RI9147190_179,RI9146a10_163,RI9146290_147,RI9145b10_131,RI9145390_115,RI9144c10_99,
        RI9144490_83,RI9143d10_67,RI9143590_51,RI90f3658_35,RI90f99b8_19,RI9138b68_3,RI91506a0_497,RI9158e18_786,RI9158da0_785,RI9158d28_784,
        RI9158cb0_783,RI9158c38_782,RI9158bc0_781,RI9158b48_780,RI9158ad0_779,RI9158a58_778,RI914ff20_481,RI914f7a0_465,RI914f020_449,RI914e8a0_433,
        RI914e120_417,RI914d9a0_401,RI914d220_385,RI914caa0_369,RI914c320_353,RI914bba0_337,RI914b420_321,RI914aca0_305,RI914a520_289,RI9149da0_273,
        RI9149620_257,RI9148f18_242,RI9148798_226,RI9148018_210,RI9147898_194,RI9147118_178,RI9146998_162,RI9146218_146,RI9145a98_130,RI9145318_114,
        RI9144b98_98,RI9144418_82,RI9143c98_66,RI9143518_50,RI90f36d0_34,RI912e758_18,RI9138be0_2,RI9150718_498,RI914ff98_482,RI914f818_466,
        RI914f098_450,RI914e918_434,RI914e198_418,RI914da18_402,RI914d298_386,RI914cb18_370,RI914c398_354,RI914bc18_338,RI914b498_322,RI914ad18_306,
        RI914a598_290,RI9149e18_274,RI9149698_258,RI9148ea0_241,RI9148720_225,RI9147fa0_209,RI9147820_193,RI91470a0_177,RI9146920_161,RI91461a0_145,
        RI9145a20_129,RI91452a0_113,RI9144b20_97,RI91443a0_81,RI9143c20_65,RI91434a0_49,RI90f3748_33,RI912e7d0_17,RI9138c58_1,RI9149008_244,
        RI9148888_228,RI9148108_212,RI9147988_196,RI9147208_180,RI9146a88_164,RI9146308_148,RI9145b88_132,RI9145408_116,RI9144c88_100,RI9144508_84,
        RI9143d88_68,RI9143608_52,RI90f35e0_36,RI90f9940_20,RI9138af0_4,RI9150790_499,RI9150010_483,RI914f890_467,RI914f110_451,RI914e990_435,
        RI914e210_419,RI914da90_403,RI914d310_387,RI914cb90_371,RI914c410_355,RI914bc90_339,RI914b510_323,RI914ad90_307,RI914a610_291,RI9149e90_275,
        RI9149710_259,RI91490f8_246,RI9148978_230,RI91481f8_214,RI9147a78_198,RI91472f8_182,RI9146b78_166,RI91463f8_150,RI9145c78_134,RI91454f8_118,
        RI9144d78_102,RI91445f8_86,RI9143e78_70,RI91436f8_54,RI90f34f0_38,RI90f9850_22,RI9138a00_6,RI9149080_245,RI9148900_229,RI9148180_213,
        RI9147a00_197,RI9147280_181,RI9146b00_165,RI9146380_149,RI9145c00_133,RI9145480_117,RI9144d00_101,RI9144580_85,RI9143e00_69,RI9143680_53,
        RI90f3568_37,RI90f98c8_21,RI9138a78_5,RI9150808_500,RI9150088_484,RI914f908_468,RI914f188_452,RI914ea08_436,RI914e288_420,RI914db08_404,
        RI914d388_388,RI914cc08_372,RI914c488_356,RI914bd08_340,RI914b588_324,RI914ae08_308,RI914a688_292,RI9149f08_276,RI9149788_260,RI9149170_247,
        RI91489f0_231,RI9148270_215,RI9147af0_199,RI9147370_183,RI9146bf0_167,RI9146470_151,RI9145cf0_135,RI9145570_119,RI9144df0_103,RI9144670_87,
        RI9143ef0_71,RI9143770_55,RI90f3478_39,RI90f97d8_23,RI9138988_7,RI9150880_501,RI9150100_485,RI914f980_469,RI914f200_453,RI914ea80_437,
        RI914e300_421,RI914db80_405,RI914d400_389,RI914cc80_373,RI914c500_357,RI914bd80_341,RI914b600_325,RI914ae80_309,RI914a700_293,RI9149f80_277,
        RI9149800_261,RI91508f8_502,RI9150178_486,RI914f9f8_470,RI914f278_454,RI914eaf8_438,RI914e378_422,RI914dbf8_406,RI914d478_390,RI914ccf8_374,
        RI914c578_358,RI914bdf8_342,RI914b678_326,RI914aef8_310,RI914a778_294,RI9149ff8_278,RI9149878_262,RI9150970_503,RI91501f0_487,RI914fa70_471,
        RI914f2f0_455,RI914eb70_439,RI914e3f0_423,RI914dc70_407,RI914d4f0_391,RI914cd70_375,RI914c5f0_359,RI914be70_343,RI914b6f0_327,RI914af70_311,
        RI914a7f0_295,RI914a070_279,RI91498f0_263,RI9149260_249,RI9148ae0_233,RI9148360_217,RI9147be0_201,RI9147460_185,RI9146ce0_169,RI9146560_153,
        RI9145de0_137,RI9145660_121,RI9144ee0_105,RI9144760_89,RI9143fe0_73,RI9143860_57,RI90f3388_41,RI90f96e8_25,RI9138898_9,RI91491e8_248,
        RI9148a68_232,RI91482e8_216,RI9147b68_200,RI91473e8_184,RI9146c68_168,RI91464e8_152,RI9145d68_136,RI91455e8_120,RI9144e68_104,RI91446e8_88,
        RI9143f68_72,RI91437e8_56,RI90f3400_40,RI90f9760_24,RI9138910_8,RI91509e8_504,RI9150268_488,RI914fae8_472,RI914f368_456,RI914ebe8_440,
        RI914e468_424,RI914dce8_408,RI914d568_392,RI914cde8_376,RI914c668_360,RI914bee8_344,RI914b768_328,RI914afe8_312,RI914a868_296,RI914a0e8_280,
        RI9149968_264,RI91492d8_250,RI9148b58_234,RI91483d8_218,RI9147c58_202,RI91474d8_186,RI9146d58_170,RI91465d8_154,RI9145e58_138,RI91456d8_122,
        RI9144f58_106,RI91447d8_90,RI9144058_74,RI91438d8_58,RI90f3310_42,RI90f9670_26,RI912eb18_10,RI9150a60_505,RI91502e0_489,RI914fb60_473,
        RI914f3e0_457,RI914ec60_441,RI914e4e0_425,RI914dd60_409,RI914d5e0_393,RI914ce60_377,RI914c6e0_361,RI914bf60_345,RI914b7e0_329,RI914b060_313,
        RI914a8e0_297,RI914a160_281,RI91499e0_265,RI91493c8_252,RI9148c48_236,RI91484c8_220,RI9147d48_204,RI91475c8_188,RI9146e48_172,RI91466c8_156,
        RI9145f48_140,RI91457c8_124,RI9145048_108,RI91448c8_92,RI9144148_76,RI91439c8_60,RI9143248_44,RI90f39a0_28,RI912ea28_12,RI9149350_251,
        RI9148bd0_235,RI9148450_219,RI9147cd0_203,RI9147550_187,RI9146dd0_171,RI9146650_155,RI9145ed0_139,RI9145750_123,RI9144fd0_107,RI9144850_91,
        RI91440d0_75,RI9143950_59,RI90f3298_43,RI90f95f8_27,RI912eaa0_11,RI9150ad8_506,RI9150358_490,RI914fbd8_474,RI914f458_458,RI914ecd8_442,
        RI914e558_426,RI914ddd8_410,RI914d658_394,RI914ced8_378,RI914c758_362,RI914bfd8_346,RI914b858_330,RI914b0d8_314,RI914a958_298,RI914a1d8_282,
        RI9149a58_266,RI9149440_253,RI9148cc0_237,RI9148540_221,RI9147dc0_205,RI9147640_189,RI9146ec0_173,RI9146740_157,RI9145fc0_141,RI9145840_125,
        RI91450c0_109,RI9144940_93,RI91441c0_77,RI9143a40_61,RI91432c0_45,RI90f3928_29,RI912e9b0_13,RI9150b50_507,RI91503d0_491,RI914fc50_475,
        RI914f4d0_459,RI914ed50_443,RI914e5d0_427,RI914de50_411,RI914d6d0_395,RI914cf50_379,RI914c7d0_363,RI914c050_347,RI914b8d0_331,RI914b150_315,
        RI914a9d0_299,RI914a250_283,RI9149ad0_267,RI9150bc8_508,RI9150448_492,RI914fcc8_476,RI914f548_460,RI914edc8_444,RI914e648_428,RI914dec8_412,
        RI914d748_396,RI914cfc8_380,RI914c848_364,RI914c0c8_348,RI914b948_332,RI914b1c8_316,RI914aa48_300,RI914a2c8_284,RI9149b48_268,RI9149530_255,
        RI9148db0_239,RI9148630_223,RI9147eb0_207,RI9147730_191,RI9146fb0_175,RI9146830_159,RI91460b0_143,RI9145930_127,RI91451b0_111,RI9144a30_95,
        RI91442b0_79,RI9143b30_63,RI91433b0_47,RI90f3838_31,RI912e8c0_15,RI91494b8_254,RI9148d38_238,RI91485b8_222,RI9147e38_206,RI91476b8_190,
        RI9146f38_174,RI91467b8_158,RI9146038_142,RI91458b8_126,RI9145138_110,RI91449b8_94,RI9144238_78,RI9143ab8_62,RI9143338_46,RI90f38b0_30,
        RI912e938_14,RI9150c40_509,RI91504c0_493,RI914fd40_477,RI914f5c0_461,RI914ee40_445,RI914e6c0_429,RI914df40_413,RI914d7c0_397,RI914d040_381,
        RI914c8c0_365,RI914c140_349,RI914b9c0_333,RI914b240_317,RI914aac0_301,RI914a340_285,RI9149bc0_269,RI91495a8_256,RI9148e28_240,RI91486a8_224,
        RI9147f28_208,RI91477a8_192,RI9147028_176,RI91468a8_160,RI9146128_144,RI91459a8_128,RI9145228_112,RI9144aa8_96,RI9144328_80,RI9143ba8_64,
        RI9143428_48,RI90f37c0_32,RI912e848_16,RI9150cb8_510,RI9150538_494,RI914fdb8_478,RI914f638_462,RI914eeb8_446,RI914e738_430,RI914dfb8_414,
        RI914d838_398,RI914d0b8_382,RI914c938_366,RI914c1b8_350,RI914ba38_334,RI914b2b8_318,RI914ab38_302,RI914a3b8_286,RI9149c38_270,RI9150d30_511,
        RI91505b0_495,RI914fe30_479,RI914f6b0_463,RI914ef30_447,RI914e7b0_431,RI914e030_415,RI914d8b0_399,RI914d130_383,RI914c9b0_367,RI914c230_351,
        RI914bab0_335,RI914b330_319,RI914abb0_303,RI914a430_287,RI9149cb0_271,RI9150da8_512,RI9150628_496,RI914fea8_480,RI914f728_464,RI914efa8_448,
        RI914e828_432,RI914e0a8_416,RI914d928_400,RI914d1a8_384,RI914ca28_368,RI914c2a8_352,RI914bb28_336,RI914b3a8_320,RI914ac28_304,RI914a4a8_288,
        RI9149d28_272,RI9157ea0_753,RI9157720_737,RI9156fa0_721,RI9156820_705,RI91560a0_689,RI9155920_673,RI91551a0_657,RI9154a20_641,RI91542a0_625,
        RI9153b20_609,RI91533a0_593,RI9152c20_577,RI91524a0_561,RI9151d20_545,RI91515a0_529,RI9150e20_513,RI9157f18_754,RI9157798_738,RI9157018_722,
        RI9156898_706,RI9156118_690,RI9155998_674,RI9155218_658,RI9154a98_642,RI9154318_626,RI9153b98_610,RI9153418_594,RI9152c98_578,RI9152518_562,
        RI9151d98_546,RI9151618_530,RI9150e98_514,RI9157f90_755,RI9157810_739,RI9157090_723,RI9156910_707,RI9156190_691,RI9155a10_675,RI9155290_659,
        RI9154b10_643,RI9154390_627,RI9153c10_611,RI9153490_595,RI9152d10_579,RI9152590_563,RI9151e10_547,RI9151690_531,RI9150f10_515,RI9158008_756,
        RI9157888_740,RI9157108_724,RI9156988_708,RI9156208_692,RI9155a88_676,RI9155308_660,RI9154b88_644,RI9154408_628,RI9153c88_612,RI9153508_596,
        RI9152d88_580,RI9152608_564,RI9151e88_548,RI9151708_532,RI9150f88_516,RI9158080_757,RI9157900_741,RI9157180_725,RI9156a00_709,RI9156280_693,
        RI9155b00_677,RI9155380_661,RI9154c00_645,RI9154480_629,RI9153d00_613,RI9153580_597,RI9152e00_581,RI9152680_565,RI9151f00_549,RI9151780_533,
        RI9151000_517,RI91580f8_758,RI9157978_742,RI91571f8_726,RI9156a78_710,RI91562f8_694,RI9155b78_678,RI91553f8_662,RI9154c78_646,RI91544f8_630,
        RI9153d78_614,RI91535f8_598,RI9152e78_582,RI91526f8_566,RI9151f78_550,RI91517f8_534,RI9151078_518,RI9158170_759,RI91579f0_743,RI9157270_727,
        RI9156af0_711,RI9156370_695,RI9155bf0_679,RI9155470_663,RI9154cf0_647,RI9154570_631,RI9153df0_615,RI9153670_599,RI9152ef0_583,RI9152770_567,
        RI9151ff0_551,RI9151870_535,RI91510f0_519,RI91581e8_760,RI9157a68_744,RI91572e8_728,RI9156b68_712,RI91563e8_696,RI9155c68_680,RI91554e8_664,
        RI9154d68_648,RI91545e8_632,RI9153e68_616,RI91536e8_600,RI9152f68_584,RI91527e8_568,RI9152068_552,RI91518e8_536,RI9151168_520,RI9158260_761,
        RI9157ae0_745,RI9157360_729,RI9156be0_713,RI9156460_697,RI9155ce0_681,RI9155560_665,RI9154de0_649,RI9154660_633,RI9153ee0_617,RI9153760_601,
        RI9152fe0_585,RI9152860_569,RI91520e0_553,RI9151960_537,RI91511e0_521,RI91582d8_762,RI9157b58_746,RI91573d8_730,RI9156c58_714,RI91564d8_698,
        RI9155d58_682,RI91555d8_666,RI9154e58_650,RI91546d8_634,RI9153f58_618,RI91537d8_602,RI9153058_586,RI91528d8_570,RI9152158_554,RI91519d8_538,
        RI9151258_522,RI9158350_763,RI9157bd0_747,RI9157450_731,RI9156cd0_715,RI9156550_699,RI9155dd0_683,RI9155650_667,RI9154ed0_651,RI9154750_635,
        RI9153fd0_619,RI9153850_603,RI91530d0_587,RI9152950_571,RI91521d0_555,RI9151a50_539,RI91512d0_523,RI91583c8_764,RI9157c48_748,RI91574c8_732,
        RI9156d48_716,RI91565c8_700,RI9155e48_684,RI91556c8_668,RI9154f48_652,RI91547c8_636,RI9154048_620,RI91538c8_604,RI9153148_588,RI91529c8_572,
        RI9152248_556,RI9151ac8_540,RI9151348_524,RI9158440_765,RI9157cc0_749,RI9157540_733,RI9156dc0_717,RI9156640_701,RI9155ec0_685,RI9155740_669,
        RI9154fc0_653,RI9154840_637,RI91540c0_621,RI9153940_605,RI91531c0_589,RI9152a40_573,RI91522c0_557,RI9151b40_541,RI91513c0_525,RI91584b8_766,
        RI9157d38_750,RI91575b8_734,RI9156e38_718,RI91566b8_702,RI9155f38_686,RI91557b8_670,RI9155038_654,RI91548b8_638,RI9154138_622,RI91539b8_606,
        RI9153238_590,RI9152ab8_574,RI9152338_558,RI9151bb8_542,RI9151438_526,RI9158530_767,RI9157db0_751,RI9157630_735,RI9156eb0_719,RI9156730_703,
        RI9155fb0_687,RI9155830_671,RI91550b0_655,RI9154930_639,RI91541b0_623,RI9153a30_607,RI91532b0_591,RI9152b30_575,RI91523b0_559,RI9151c30_543,
        RI91514b0_527,RI91585a8_768,RI9157e28_752,RI91576a8_736,RI9156f28_720,RI91567a8_704,RI9156028_688,RI91558a8_672,RI9155128_656,RI91549a8_640,
        RI9154228_624,RI9153aa8_608,RI9153328_592,RI9152ba8_576,RI9152428_560,RI9151ca8_544,RI9151528_528,R_313_9fdbc38,R_314_9fdbce0,R_315_9fdbd88,
        R_316_9fdbe30,R_317_9fdbed8,R_318_9fdbf80,R_319_9fdc028,R_31a_9fdc0d0,R_31b_9fdc178,R_31c_9fdc220,R_31d_9fdc2c8,R_31e_9fdc370,R_31f_9fdc418,
        R_320_9fdc4c0,R_321_9fdc568,R_322_9fdc610,R_323_9fdc6b8,R_324_9fdc760,R_325_9fdc808,R_326_9fdc8b0,R_327_9fdc958,R_328_9fdca00,R_329_9fdcaa8,
        R_32a_9fdcb50,R_32b_9fdcbf8,R_32c_9fdcca0,R_32d_9fdcd48);
input RI9148f90_243,RI91589e0_777,RI9158968_776,RI91588f0_775,RI9158878_774,RI9158800_773,RI9158788_772,RI9158710_771,RI9158698_770,
        RI9158620_769,RI9148810_227,RI9148090_211,RI9147910_195,RI9147190_179,RI9146a10_163,RI9146290_147,RI9145b10_131,RI9145390_115,RI9144c10_99,
        RI9144490_83,RI9143d10_67,RI9143590_51,RI90f3658_35,RI90f99b8_19,RI9138b68_3,RI91506a0_497,RI9158e18_786,RI9158da0_785,RI9158d28_784,
        RI9158cb0_783,RI9158c38_782,RI9158bc0_781,RI9158b48_780,RI9158ad0_779,RI9158a58_778,RI914ff20_481,RI914f7a0_465,RI914f020_449,RI914e8a0_433,
        RI914e120_417,RI914d9a0_401,RI914d220_385,RI914caa0_369,RI914c320_353,RI914bba0_337,RI914b420_321,RI914aca0_305,RI914a520_289,RI9149da0_273,
        RI9149620_257,RI9148f18_242,RI9148798_226,RI9148018_210,RI9147898_194,RI9147118_178,RI9146998_162,RI9146218_146,RI9145a98_130,RI9145318_114,
        RI9144b98_98,RI9144418_82,RI9143c98_66,RI9143518_50,RI90f36d0_34,RI912e758_18,RI9138be0_2,RI9150718_498,RI914ff98_482,RI914f818_466,
        RI914f098_450,RI914e918_434,RI914e198_418,RI914da18_402,RI914d298_386,RI914cb18_370,RI914c398_354,RI914bc18_338,RI914b498_322,RI914ad18_306,
        RI914a598_290,RI9149e18_274,RI9149698_258,RI9148ea0_241,RI9148720_225,RI9147fa0_209,RI9147820_193,RI91470a0_177,RI9146920_161,RI91461a0_145,
        RI9145a20_129,RI91452a0_113,RI9144b20_97,RI91443a0_81,RI9143c20_65,RI91434a0_49,RI90f3748_33,RI912e7d0_17,RI9138c58_1,RI9149008_244,
        RI9148888_228,RI9148108_212,RI9147988_196,RI9147208_180,RI9146a88_164,RI9146308_148,RI9145b88_132,RI9145408_116,RI9144c88_100,RI9144508_84,
        RI9143d88_68,RI9143608_52,RI90f35e0_36,RI90f9940_20,RI9138af0_4,RI9150790_499,RI9150010_483,RI914f890_467,RI914f110_451,RI914e990_435,
        RI914e210_419,RI914da90_403,RI914d310_387,RI914cb90_371,RI914c410_355,RI914bc90_339,RI914b510_323,RI914ad90_307,RI914a610_291,RI9149e90_275,
        RI9149710_259,RI91490f8_246,RI9148978_230,RI91481f8_214,RI9147a78_198,RI91472f8_182,RI9146b78_166,RI91463f8_150,RI9145c78_134,RI91454f8_118,
        RI9144d78_102,RI91445f8_86,RI9143e78_70,RI91436f8_54,RI90f34f0_38,RI90f9850_22,RI9138a00_6,RI9149080_245,RI9148900_229,RI9148180_213,
        RI9147a00_197,RI9147280_181,RI9146b00_165,RI9146380_149,RI9145c00_133,RI9145480_117,RI9144d00_101,RI9144580_85,RI9143e00_69,RI9143680_53,
        RI90f3568_37,RI90f98c8_21,RI9138a78_5,RI9150808_500,RI9150088_484,RI914f908_468,RI914f188_452,RI914ea08_436,RI914e288_420,RI914db08_404,
        RI914d388_388,RI914cc08_372,RI914c488_356,RI914bd08_340,RI914b588_324,RI914ae08_308,RI914a688_292,RI9149f08_276,RI9149788_260,RI9149170_247,
        RI91489f0_231,RI9148270_215,RI9147af0_199,RI9147370_183,RI9146bf0_167,RI9146470_151,RI9145cf0_135,RI9145570_119,RI9144df0_103,RI9144670_87,
        RI9143ef0_71,RI9143770_55,RI90f3478_39,RI90f97d8_23,RI9138988_7,RI9150880_501,RI9150100_485,RI914f980_469,RI914f200_453,RI914ea80_437,
        RI914e300_421,RI914db80_405,RI914d400_389,RI914cc80_373,RI914c500_357,RI914bd80_341,RI914b600_325,RI914ae80_309,RI914a700_293,RI9149f80_277,
        RI9149800_261,RI91508f8_502,RI9150178_486,RI914f9f8_470,RI914f278_454,RI914eaf8_438,RI914e378_422,RI914dbf8_406,RI914d478_390,RI914ccf8_374,
        RI914c578_358,RI914bdf8_342,RI914b678_326,RI914aef8_310,RI914a778_294,RI9149ff8_278,RI9149878_262,RI9150970_503,RI91501f0_487,RI914fa70_471,
        RI914f2f0_455,RI914eb70_439,RI914e3f0_423,RI914dc70_407,RI914d4f0_391,RI914cd70_375,RI914c5f0_359,RI914be70_343,RI914b6f0_327,RI914af70_311,
        RI914a7f0_295,RI914a070_279,RI91498f0_263,RI9149260_249,RI9148ae0_233,RI9148360_217,RI9147be0_201,RI9147460_185,RI9146ce0_169,RI9146560_153,
        RI9145de0_137,RI9145660_121,RI9144ee0_105,RI9144760_89,RI9143fe0_73,RI9143860_57,RI90f3388_41,RI90f96e8_25,RI9138898_9,RI91491e8_248,
        RI9148a68_232,RI91482e8_216,RI9147b68_200,RI91473e8_184,RI9146c68_168,RI91464e8_152,RI9145d68_136,RI91455e8_120,RI9144e68_104,RI91446e8_88,
        RI9143f68_72,RI91437e8_56,RI90f3400_40,RI90f9760_24,RI9138910_8,RI91509e8_504,RI9150268_488,RI914fae8_472,RI914f368_456,RI914ebe8_440,
        RI914e468_424,RI914dce8_408,RI914d568_392,RI914cde8_376,RI914c668_360,RI914bee8_344,RI914b768_328,RI914afe8_312,RI914a868_296,RI914a0e8_280,
        RI9149968_264,RI91492d8_250,RI9148b58_234,RI91483d8_218,RI9147c58_202,RI91474d8_186,RI9146d58_170,RI91465d8_154,RI9145e58_138,RI91456d8_122,
        RI9144f58_106,RI91447d8_90,RI9144058_74,RI91438d8_58,RI90f3310_42,RI90f9670_26,RI912eb18_10,RI9150a60_505,RI91502e0_489,RI914fb60_473,
        RI914f3e0_457,RI914ec60_441,RI914e4e0_425,RI914dd60_409,RI914d5e0_393,RI914ce60_377,RI914c6e0_361,RI914bf60_345,RI914b7e0_329,RI914b060_313,
        RI914a8e0_297,RI914a160_281,RI91499e0_265,RI91493c8_252,RI9148c48_236,RI91484c8_220,RI9147d48_204,RI91475c8_188,RI9146e48_172,RI91466c8_156,
        RI9145f48_140,RI91457c8_124,RI9145048_108,RI91448c8_92,RI9144148_76,RI91439c8_60,RI9143248_44,RI90f39a0_28,RI912ea28_12,RI9149350_251,
        RI9148bd0_235,RI9148450_219,RI9147cd0_203,RI9147550_187,RI9146dd0_171,RI9146650_155,RI9145ed0_139,RI9145750_123,RI9144fd0_107,RI9144850_91,
        RI91440d0_75,RI9143950_59,RI90f3298_43,RI90f95f8_27,RI912eaa0_11,RI9150ad8_506,RI9150358_490,RI914fbd8_474,RI914f458_458,RI914ecd8_442,
        RI914e558_426,RI914ddd8_410,RI914d658_394,RI914ced8_378,RI914c758_362,RI914bfd8_346,RI914b858_330,RI914b0d8_314,RI914a958_298,RI914a1d8_282,
        RI9149a58_266,RI9149440_253,RI9148cc0_237,RI9148540_221,RI9147dc0_205,RI9147640_189,RI9146ec0_173,RI9146740_157,RI9145fc0_141,RI9145840_125,
        RI91450c0_109,RI9144940_93,RI91441c0_77,RI9143a40_61,RI91432c0_45,RI90f3928_29,RI912e9b0_13,RI9150b50_507,RI91503d0_491,RI914fc50_475,
        RI914f4d0_459,RI914ed50_443,RI914e5d0_427,RI914de50_411,RI914d6d0_395,RI914cf50_379,RI914c7d0_363,RI914c050_347,RI914b8d0_331,RI914b150_315,
        RI914a9d0_299,RI914a250_283,RI9149ad0_267,RI9150bc8_508,RI9150448_492,RI914fcc8_476,RI914f548_460,RI914edc8_444,RI914e648_428,RI914dec8_412,
        RI914d748_396,RI914cfc8_380,RI914c848_364,RI914c0c8_348,RI914b948_332,RI914b1c8_316,RI914aa48_300,RI914a2c8_284,RI9149b48_268,RI9149530_255,
        RI9148db0_239,RI9148630_223,RI9147eb0_207,RI9147730_191,RI9146fb0_175,RI9146830_159,RI91460b0_143,RI9145930_127,RI91451b0_111,RI9144a30_95,
        RI91442b0_79,RI9143b30_63,RI91433b0_47,RI90f3838_31,RI912e8c0_15,RI91494b8_254,RI9148d38_238,RI91485b8_222,RI9147e38_206,RI91476b8_190,
        RI9146f38_174,RI91467b8_158,RI9146038_142,RI91458b8_126,RI9145138_110,RI91449b8_94,RI9144238_78,RI9143ab8_62,RI9143338_46,RI90f38b0_30,
        RI912e938_14,RI9150c40_509,RI91504c0_493,RI914fd40_477,RI914f5c0_461,RI914ee40_445,RI914e6c0_429,RI914df40_413,RI914d7c0_397,RI914d040_381,
        RI914c8c0_365,RI914c140_349,RI914b9c0_333,RI914b240_317,RI914aac0_301,RI914a340_285,RI9149bc0_269,RI91495a8_256,RI9148e28_240,RI91486a8_224,
        RI9147f28_208,RI91477a8_192,RI9147028_176,RI91468a8_160,RI9146128_144,RI91459a8_128,RI9145228_112,RI9144aa8_96,RI9144328_80,RI9143ba8_64,
        RI9143428_48,RI90f37c0_32,RI912e848_16,RI9150cb8_510,RI9150538_494,RI914fdb8_478,RI914f638_462,RI914eeb8_446,RI914e738_430,RI914dfb8_414,
        RI914d838_398,RI914d0b8_382,RI914c938_366,RI914c1b8_350,RI914ba38_334,RI914b2b8_318,RI914ab38_302,RI914a3b8_286,RI9149c38_270,RI9150d30_511,
        RI91505b0_495,RI914fe30_479,RI914f6b0_463,RI914ef30_447,RI914e7b0_431,RI914e030_415,RI914d8b0_399,RI914d130_383,RI914c9b0_367,RI914c230_351,
        RI914bab0_335,RI914b330_319,RI914abb0_303,RI914a430_287,RI9149cb0_271,RI9150da8_512,RI9150628_496,RI914fea8_480,RI914f728_464,RI914efa8_448,
        RI914e828_432,RI914e0a8_416,RI914d928_400,RI914d1a8_384,RI914ca28_368,RI914c2a8_352,RI914bb28_336,RI914b3a8_320,RI914ac28_304,RI914a4a8_288,
        RI9149d28_272,RI9157ea0_753,RI9157720_737,RI9156fa0_721,RI9156820_705,RI91560a0_689,RI9155920_673,RI91551a0_657,RI9154a20_641,RI91542a0_625,
        RI9153b20_609,RI91533a0_593,RI9152c20_577,RI91524a0_561,RI9151d20_545,RI91515a0_529,RI9150e20_513,RI9157f18_754,RI9157798_738,RI9157018_722,
        RI9156898_706,RI9156118_690,RI9155998_674,RI9155218_658,RI9154a98_642,RI9154318_626,RI9153b98_610,RI9153418_594,RI9152c98_578,RI9152518_562,
        RI9151d98_546,RI9151618_530,RI9150e98_514,RI9157f90_755,RI9157810_739,RI9157090_723,RI9156910_707,RI9156190_691,RI9155a10_675,RI9155290_659,
        RI9154b10_643,RI9154390_627,RI9153c10_611,RI9153490_595,RI9152d10_579,RI9152590_563,RI9151e10_547,RI9151690_531,RI9150f10_515,RI9158008_756,
        RI9157888_740,RI9157108_724,RI9156988_708,RI9156208_692,RI9155a88_676,RI9155308_660,RI9154b88_644,RI9154408_628,RI9153c88_612,RI9153508_596,
        RI9152d88_580,RI9152608_564,RI9151e88_548,RI9151708_532,RI9150f88_516,RI9158080_757,RI9157900_741,RI9157180_725,RI9156a00_709,RI9156280_693,
        RI9155b00_677,RI9155380_661,RI9154c00_645,RI9154480_629,RI9153d00_613,RI9153580_597,RI9152e00_581,RI9152680_565,RI9151f00_549,RI9151780_533,
        RI9151000_517,RI91580f8_758,RI9157978_742,RI91571f8_726,RI9156a78_710,RI91562f8_694,RI9155b78_678,RI91553f8_662,RI9154c78_646,RI91544f8_630,
        RI9153d78_614,RI91535f8_598,RI9152e78_582,RI91526f8_566,RI9151f78_550,RI91517f8_534,RI9151078_518,RI9158170_759,RI91579f0_743,RI9157270_727,
        RI9156af0_711,RI9156370_695,RI9155bf0_679,RI9155470_663,RI9154cf0_647,RI9154570_631,RI9153df0_615,RI9153670_599,RI9152ef0_583,RI9152770_567,
        RI9151ff0_551,RI9151870_535,RI91510f0_519,RI91581e8_760,RI9157a68_744,RI91572e8_728,RI9156b68_712,RI91563e8_696,RI9155c68_680,RI91554e8_664,
        RI9154d68_648,RI91545e8_632,RI9153e68_616,RI91536e8_600,RI9152f68_584,RI91527e8_568,RI9152068_552,RI91518e8_536,RI9151168_520,RI9158260_761,
        RI9157ae0_745,RI9157360_729,RI9156be0_713,RI9156460_697,RI9155ce0_681,RI9155560_665,RI9154de0_649,RI9154660_633,RI9153ee0_617,RI9153760_601,
        RI9152fe0_585,RI9152860_569,RI91520e0_553,RI9151960_537,RI91511e0_521,RI91582d8_762,RI9157b58_746,RI91573d8_730,RI9156c58_714,RI91564d8_698,
        RI9155d58_682,RI91555d8_666,RI9154e58_650,RI91546d8_634,RI9153f58_618,RI91537d8_602,RI9153058_586,RI91528d8_570,RI9152158_554,RI91519d8_538,
        RI9151258_522,RI9158350_763,RI9157bd0_747,RI9157450_731,RI9156cd0_715,RI9156550_699,RI9155dd0_683,RI9155650_667,RI9154ed0_651,RI9154750_635,
        RI9153fd0_619,RI9153850_603,RI91530d0_587,RI9152950_571,RI91521d0_555,RI9151a50_539,RI91512d0_523,RI91583c8_764,RI9157c48_748,RI91574c8_732,
        RI9156d48_716,RI91565c8_700,RI9155e48_684,RI91556c8_668,RI9154f48_652,RI91547c8_636,RI9154048_620,RI91538c8_604,RI9153148_588,RI91529c8_572,
        RI9152248_556,RI9151ac8_540,RI9151348_524,RI9158440_765,RI9157cc0_749,RI9157540_733,RI9156dc0_717,RI9156640_701,RI9155ec0_685,RI9155740_669,
        RI9154fc0_653,RI9154840_637,RI91540c0_621,RI9153940_605,RI91531c0_589,RI9152a40_573,RI91522c0_557,RI9151b40_541,RI91513c0_525,RI91584b8_766,
        RI9157d38_750,RI91575b8_734,RI9156e38_718,RI91566b8_702,RI9155f38_686,RI91557b8_670,RI9155038_654,RI91548b8_638,RI9154138_622,RI91539b8_606,
        RI9153238_590,RI9152ab8_574,RI9152338_558,RI9151bb8_542,RI9151438_526,RI9158530_767,RI9157db0_751,RI9157630_735,RI9156eb0_719,RI9156730_703,
        RI9155fb0_687,RI9155830_671,RI91550b0_655,RI9154930_639,RI91541b0_623,RI9153a30_607,RI91532b0_591,RI9152b30_575,RI91523b0_559,RI9151c30_543,
        RI91514b0_527,RI91585a8_768,RI9157e28_752,RI91576a8_736,RI9156f28_720,RI91567a8_704,RI9156028_688,RI91558a8_672,RI9155128_656,RI91549a8_640,
        RI9154228_624,RI9153aa8_608,RI9153328_592,RI9152ba8_576,RI9152428_560,RI9151ca8_544,RI9151528_528;
output R_313_9fdbc38,R_314_9fdbce0,R_315_9fdbd88,R_316_9fdbe30,R_317_9fdbed8,R_318_9fdbf80,R_319_9fdc028,R_31a_9fdc0d0,R_31b_9fdc178,
        R_31c_9fdc220,R_31d_9fdc2c8,R_31e_9fdc370,R_31f_9fdc418,R_320_9fdc4c0,R_321_9fdc568,R_322_9fdc610,R_323_9fdc6b8,R_324_9fdc760,R_325_9fdc808,
        R_326_9fdc8b0,R_327_9fdc958,R_328_9fdca00,R_329_9fdcaa8,R_32a_9fdcb50,R_32b_9fdcbf8,R_32c_9fdcca0,R_32d_9fdcd48;

wire \814 , \815_ZERO , \816_ONE , \817 , \818 , \819 , \820 , \821 , \822 ,
         \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 ,
         \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 ,
         \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 ,
         \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861_nG395 , \862 ,
         \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 ,
         \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 ,
         \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 ,
         \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 ,
         \903 , \904 , \905 , \906 , \907 , \908 , \909_nG3c5 , \910 , \911 , \912 ,
         \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 ,
         \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932_nG3dc ,
         \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 ,
         \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952_nG3f0 ,
         \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 ,
         \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 ,
         \973 , \974_nG406 , \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 ,
         \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 ,
         \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 ,
         \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010_nG42b , \1011 , \1012 ,
         \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 ,
         \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 ,
         \1033 , \1034 , \1035_nG444 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 ,
         \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 ,
         \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059_nG45c , \1060 , \1061 , \1062 ,
         \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 ,
         \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082_nG473 ,
         \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 ,
         \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 ,
         \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111_nG490 , \1112 ,
         \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 ,
         \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 ,
         \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
         \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 ,
         \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 ,
         \1163_nG4c4 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 ,
         \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 ,
         \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 ,
         \1193 , \1194 , \1195_nG4e4 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 ,
         \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 ,
         \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 ,
         \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 ,
         \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 ,
         \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 ,
         \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259_nG524 , \1260 , \1261 , \1262 ,
         \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 ,
         \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 ,
         \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 ,
         \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 ,
         \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 ,
         \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 ,
         \1323 , \1324_nG565 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 ,
         \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 ,
         \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352_nG581 ,
         \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 ,
         \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 ,
         \1373 , \1374 , \1375_nG598 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 ,
         \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 ,
         \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 ,
         \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 ,
         \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 ,
         \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 ,
         \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 ,
         \1443 , \1444_nG5dd , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 ,
         \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 ,
         \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469_nG5f6 , \1470 , \1471 , \1472 ,
         \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 ,
         \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 ,
         \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 ,
         \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 ,
         \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 ,
         \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 ,
         \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 ,
         \1543 , \1544 , \1545 , \1546 , \1547 , \1548_nG645 , \1549 , \1550 , \1551 , \1552 ,
         \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 ,
         \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 ,
         \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 ,
         \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 ,
         \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 ,
         \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 ,
         \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 ,
         \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631_nG698 , \1632 ,
         \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 ,
         \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 ,
         \1653 , \1654_nG6af , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 ,
         \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 ,
         \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 ,
         \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 ,
         \1693 , \1694 , \1695_nG6d8 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 ,
         \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 ,
         \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 ,
         \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 ,
         \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 ,
         \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 ,
         \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 ,
         \1763 , \1764 , \1765 , \1766 , \1767_nG720 , \1768 , \1769 , \1770 , \1771 , \1772 ,
         \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 ,
         \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 ,
         \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 ,
         \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 ,
         \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822_nG757 ,
         \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 ,
         \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 ,
         \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 ,
         \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 ,
         \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 ,
         \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 ,
         \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 ,
         \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 ,
         \1903 , \1904 , \1905 , \1906_nG7ab , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 ,
         \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 ,
         \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 ,
         \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 ,
         \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 ,
         \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 ,
         \1963 , \1964_nG7e5 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 ,
         \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 ,
         \1983 , \1984 , \1985 , \1986 , \1987_nG7fc , \1988 , \1989 , \1990 , \1991 , \1992 ,
         \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 ,
         \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 ,
         \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 ,
         \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 ,
         \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 ,
         \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 ,
         \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 ,
         \2063 , \2064 , \2065_nG84a , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 ,
         \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 ,
         \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 ,
         \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 ,
         \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 ,
         \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 ,
         \2123 , \2124 , \2125 , \2126_nG887 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 ,
         \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 ,
         \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 ,
         \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 ,
         \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 ,
         \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 ,
         \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 ,
         \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 ,
         \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210_nG8db , \2211 , \2212 ,
         \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 ,
         \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 ,
         \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 ,
         \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 ,
         \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 ,
         \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 ,
         \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 ,
         \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 ,
         \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 ,
         \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 ,
         \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 ,
         \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 ,
         \2333 , \2334_nG957 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 ,
         \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 ,
         \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 ,
         \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 ,
         \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 ,
         \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 ,
         \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 ,
         \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 ,
         \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 ,
         \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 ,
         \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 ,
         \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 ,
         \2453 , \2454 , \2455 , \2456 , \2457 , \2458_nG9d3 , \2459 , \2460 , \2461 , \2462 ,
         \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 ,
         \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 ,
         \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 ,
         \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 ,
         \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 ,
         \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 ,
         \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 ,
         \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 ,
         \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 ,
         \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 ,
         \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 ,
         \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 ,
         \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 ,
         \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 ,
         \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 ,
         \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 ,
         \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 ,
         \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 ,
         \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 ,
         \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 ,
         \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 ,
         \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 ,
         \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 ,
         \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 ,
         \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 ,
         \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 ,
         \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 ,
         \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 ,
         \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 ,
         \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 ,
         \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 ,
         \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 ,
         \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 ,
         \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 ,
         \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 ,
         \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 ,
         \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 ,
         \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 ,
         \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 ,
         \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 ,
         \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 ,
         \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 ,
         \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 ,
         \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 ,
         \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 ,
         \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 ,
         \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 ,
         \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 ,
         \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 ,
         \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 ,
         \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 ,
         \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 ,
         \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 ,
         \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 ,
         \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 ,
         \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 ,
         \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 ,
         \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 ,
         \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 ,
         \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 ,
         \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 ,
         \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 ,
         \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 ,
         \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 ,
         \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 ,
         \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 ,
         \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 ,
         \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 ,
         \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 ,
         \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 ,
         \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 ,
         \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 ,
         \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191_nGcb0 , \3192 ,
         \3193 , \3194_nGcb3 , \3195 , \3196 , \3197_nGcb6 , \3198 , \3199 , \3200_nGcb9 , \3201 , \3202 ,
         \3203_nGcbc , \3204 , \3205 , \3206_nGcbf , \3207 , \3208 , \3209_nGcc2 , \3210 , \3211 , \3212_nGcc5 ,
         \3213 , \3214 , \3215_nGcc8 , \3216 , \3217 , \3218_nGccb , \3219 , \3220 , \3221_nGcce , \3222 ,
         \3223 , \3224_nGcd1 , \3225 , \3226 , \3227_nGcd4 , \3228 , \3229 , \3230_nGcd7 , \3231 , \3232 ,
         \3233_nGcda , \3234 , \3235 , \3236_nGcdd , \3237 , \3238 , \3239_nGce0 , \3240 , \3241 , \3242 ,
         \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 ,
         \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 ,
         \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 ,
         \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281_nGd37 , \3282 ,
         \3283 , \3284 , \3285_nGce3 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 ,
         \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 ,
         \3303 , \3304_nGd4a , \3305 , \3306 , \3307 , \3308_nGce6 , \3309 , \3310 , \3311 , \3312 ,
         \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 ,
         \3323 , \3324 , \3325 , \3326 , \3327_nGd5d , \3328 , \3329 , \3330 , \3331_nGce9 , \3332 ,
         \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 ,
         \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350_nGd70 , \3351 , \3352 ,
         \3353 , \3354_nGcec , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 ,
         \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 ,
         \3373_nGd83 , \3374 , \3375 , \3376 , \3377_nGcef , \3378 , \3379 , \3380 , \3381 , \3382 ,
         \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 ,
         \3393 , \3394 , \3395 , \3396_nGd96 , \3397 , \3398 , \3399 , \3400_nGcf2 , \3401 , \3402 ,
         \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 ,
         \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419_nGda9 , \3420 , \3421 , \3422 ,
         \3423_nGcf5 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 ,
         \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442_nGdbc ,
         \3443 , \3444 , \3445 , \3446_nGcf8 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 ,
         \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 ,
         \3463 , \3464 , \3465_nGdcf , \3466 , \3467 , \3468 , \3469_nGcfb , \3470 , \3471 , \3472 ,
         \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 ,
         \3483 , \3484 , \3485 , \3486 , \3487 , \3488_nGde2 , \3489 , \3490 , \3491 , \3492_nGcfe ,
         \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 ,
         \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511_nGdf5 , \3512 ,
         \3513 , \3514 , \3515_nGd01 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 ,
         \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 ,
         \3533 , \3534_nGe08 , \3535 , \3536 , \3537 , \3538_nGd04 , \3539 , \3540 , \3541 , \3542 ,
         \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 ,
         \3553 , \3554 , \3555 , \3556 , \3557_nGe1b , \3558 , \3559 , \3560 , \3561_nGd07 , \3562 ,
         \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 ,
         \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580_nGe2e , \3581 , \3582 ,
         \3583 , \3584_nGd0a , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 ,
         \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 ,
         \3603_nGe41 , \3604 , \3605 , \3606 , \3607_nGd0d , \3608 , \3609 , \3610 , \3611 , \3612 ,
         \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 ,
         \3623 , \3624 , \3625 , \3626_nGe54 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 ,
         \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 ,
         \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 ,
         \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 ,
         \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 ,
         \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 ,
         \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 ,
         \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 ,
         \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 ,
         \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 ,
         \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 ,
         \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 ,
         \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 ,
         \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 ,
         \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 ,
         \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 ;
buf \U$labajz466 ( R_313_9fdbc38, \3691 );
buf \U$labajz467 ( R_314_9fdbce0, \3694 );
buf \U$labajz468 ( R_315_9fdbd88, \3697 );
buf \U$labajz469 ( R_316_9fdbe30, \3700 );
buf \U$labajz470 ( R_317_9fdbed8, \3703 );
buf \U$labajz471 ( R_318_9fdbf80, \3706 );
buf \U$labajz472 ( R_319_9fdc028, \3709 );
buf \U$labajz473 ( R_31a_9fdc0d0, \3712 );
buf \U$labajz474 ( R_31b_9fdc178, \3715 );
buf \U$labajz475 ( R_31c_9fdc220, \3718 );
buf \U$labajz476 ( R_31d_9fdc2c8, \3721 );
buf \U$labajz477 ( R_31e_9fdc370, \3724 );
buf \U$labajz478 ( R_31f_9fdc418, \3727 );
buf \U$labajz479 ( R_320_9fdc4c0, \3730 );
buf \U$labajz480 ( R_321_9fdc568, \3733 );
buf \U$labajz481 ( R_322_9fdc610, \3736 );
buf \U$labajz482 ( R_323_9fdc6b8, \3740 );
buf \U$labajz483 ( R_324_9fdc760, \3744 );
buf \U$labajz484 ( R_325_9fdc808, \3748 );
buf \U$labajz485 ( R_326_9fdc8b0, \3752 );
buf \U$labajz486 ( R_327_9fdc958, \3756 );
buf \U$labajz487 ( R_328_9fdca00, \3760 );
buf \U$labajz488 ( R_329_9fdcaa8, \3764 );
buf \U$labajz489 ( R_32a_9fdcb50, \3768 );
buf \U$labajz490 ( R_32b_9fdcbf8, \3772 );
buf \U$labajz491 ( R_32c_9fdcca0, \3776 );
buf \U$labajz492 ( R_32d_9fdcd48, \3780 );
not \U$1 ( \817 , RI91589e0_777);
not \U$2 ( \818 , RI9158968_776);
not \U$3 ( \819 , RI91588f0_775);
not \U$4 ( \820 , RI9158878_774);
nor \U$5 ( \821 , \817 , \818 , \819 , \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$6 ( \822 , RI9148f90_243, \821 );
nor \U$7 ( \823 , RI91589e0_777, \818 , \819 , \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$8 ( \824 , RI9148810_227, \823 );
nor \U$9 ( \825 , \817 , RI9158968_776, \819 , \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$10 ( \826 , RI9148090_211, \825 );
nor \U$11 ( \827 , RI91589e0_777, RI9158968_776, \819 , \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$12 ( \828 , RI9147910_195, \827 );
nor \U$13 ( \829 , \817 , \818 , RI91588f0_775, \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$14 ( \830 , RI9147190_179, \829 );
nor \U$15 ( \831 , RI91589e0_777, \818 , RI91588f0_775, \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$16 ( \832 , RI9146a10_163, \831 );
nor \U$17 ( \833 , \817 , RI9158968_776, RI91588f0_775, \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$18 ( \834 , RI9146290_147, \833 );
nor \U$19 ( \835 , RI91589e0_777, RI9158968_776, RI91588f0_775, \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$20 ( \836 , RI9145b10_131, \835 );
nor \U$21 ( \837 , \817 , \818 , \819 , RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$22 ( \838 , RI9145390_115, \837 );
nor \U$23 ( \839 , RI91589e0_777, \818 , \819 , RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$24 ( \840 , RI9144c10_99, \839 );
nor \U$25 ( \841 , \817 , RI9158968_776, \819 , RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$26 ( \842 , RI9144490_83, \841 );
nor \U$27 ( \843 , RI91589e0_777, RI9158968_776, \819 , RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$28 ( \844 , RI9143d10_67, \843 );
nor \U$29 ( \845 , \817 , \818 , RI91588f0_775, RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$30 ( \846 , RI9143590_51, \845 );
nor \U$31 ( \847 , RI91589e0_777, \818 , RI91588f0_775, RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$32 ( \848 , RI90f3658_35, \847 );
nor \U$33 ( \849 , \817 , RI9158968_776, RI91588f0_775, RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$34 ( \850 , RI90f99b8_19, \849 );
nor \U$35 ( \851 , RI91589e0_777, RI9158968_776, RI91588f0_775, RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$36 ( \852 , RI9138b68_3, \851 );
or \U$37 ( \853 , \822 , \824 , \826 , \828 , \830 , \832 , \834 , \836 , \838 , \840 , \842 , \844 , \846 , \848 , \850 , \852 );
buf \U$38 ( \854 , RI9158800_773);
buf \U$39 ( \855 , RI9158788_772);
buf \U$40 ( \856 , RI9158710_771);
buf \U$41 ( \857 , RI9158698_770);
buf \U$42 ( \858 , RI9158620_769);
or \U$43 ( \859 , \854 , \855 , \856 , \857 , \858 );
buf \U$44 ( \860 , \859 );
_DC g395 ( \861_nG395 , \853 , \860 );
buf \U$45 ( \862 , \861_nG395 );
buf \U$46 ( \863 , \862 );
not \U$47 ( \864 , \863 );
not \U$48 ( \865 , RI9158e18_786);
not \U$49 ( \866 , RI9158da0_785);
not \U$50 ( \867 , RI9158d28_784);
not \U$51 ( \868 , RI9158cb0_783);
nor \U$52 ( \869 , \865 , \866 , \867 , \868 , RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$53 ( \870 , RI91506a0_497, \869 );
nor \U$54 ( \871 , RI9158e18_786, \866 , \867 , \868 , RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$55 ( \872 , RI914ff20_481, \871 );
nor \U$56 ( \873 , \865 , RI9158da0_785, \867 , \868 , RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$57 ( \874 , RI914f7a0_465, \873 );
nor \U$58 ( \875 , RI9158e18_786, RI9158da0_785, \867 , \868 , RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$59 ( \876 , RI914f020_449, \875 );
nor \U$60 ( \877 , \865 , \866 , RI9158d28_784, \868 , RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$61 ( \878 , RI914e8a0_433, \877 );
nor \U$62 ( \879 , RI9158e18_786, \866 , RI9158d28_784, \868 , RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$63 ( \880 , RI914e120_417, \879 );
nor \U$64 ( \881 , \865 , RI9158da0_785, RI9158d28_784, \868 , RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$65 ( \882 , RI914d9a0_401, \881 );
nor \U$66 ( \883 , RI9158e18_786, RI9158da0_785, RI9158d28_784, \868 , RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$67 ( \884 , RI914d220_385, \883 );
nor \U$68 ( \885 , \865 , \866 , \867 , RI9158cb0_783, RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$69 ( \886 , RI914caa0_369, \885 );
nor \U$70 ( \887 , RI9158e18_786, \866 , \867 , RI9158cb0_783, RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$71 ( \888 , RI914c320_353, \887 );
nor \U$72 ( \889 , \865 , RI9158da0_785, \867 , RI9158cb0_783, RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$73 ( \890 , RI914bba0_337, \889 );
nor \U$74 ( \891 , RI9158e18_786, RI9158da0_785, \867 , RI9158cb0_783, RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$75 ( \892 , RI914b420_321, \891 );
nor \U$76 ( \893 , \865 , \866 , RI9158d28_784, RI9158cb0_783, RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$77 ( \894 , RI914aca0_305, \893 );
nor \U$78 ( \895 , RI9158e18_786, \866 , RI9158d28_784, RI9158cb0_783, RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$79 ( \896 , RI914a520_289, \895 );
nor \U$80 ( \897 , \865 , RI9158da0_785, RI9158d28_784, RI9158cb0_783, RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$81 ( \898 , RI9149da0_273, \897 );
nor \U$82 ( \899 , RI9158e18_786, RI9158da0_785, RI9158d28_784, RI9158cb0_783, RI9158c38_782, RI9158bc0_781, RI9158b48_780, RI9158ad0_779, RI9158a58_778);
and \U$83 ( \900 , RI9149620_257, \899 );
or \U$84 ( \901 , \870 , \872 , \874 , \876 , \878 , \880 , \882 , \884 , \886 , \888 , \890 , \892 , \894 , \896 , \898 , \900 );
buf \U$85 ( \902 , RI9158c38_782);
buf \U$86 ( \903 , RI9158bc0_781);
buf \U$87 ( \904 , RI9158b48_780);
buf \U$88 ( \905 , RI9158ad0_779);
buf \U$89 ( \906 , RI9158a58_778);
or \U$90 ( \907 , \902 , \903 , \904 , \905 , \906 );
buf \U$91 ( \908 , \907 );
_DC g3c5 ( \909_nG3c5 , \901 , \908 );
buf \U$92 ( \910 , \909_nG3c5 );
buf \U$93 ( \911 , \910 );
not \U$94 ( \912 , \911 );
and \U$95 ( \913 , \912 , \863 );
nor \U$96 ( \914 , \864 , \913 );
and \U$97 ( \915 , RI9148f18_242, \821 );
and \U$98 ( \916 , RI9148798_226, \823 );
and \U$99 ( \917 , RI9148018_210, \825 );
and \U$100 ( \918 , RI9147898_194, \827 );
and \U$101 ( \919 , RI9147118_178, \829 );
and \U$102 ( \920 , RI9146998_162, \831 );
and \U$103 ( \921 , RI9146218_146, \833 );
and \U$104 ( \922 , RI9145a98_130, \835 );
and \U$105 ( \923 , RI9145318_114, \837 );
and \U$106 ( \924 , RI9144b98_98, \839 );
and \U$107 ( \925 , RI9144418_82, \841 );
and \U$108 ( \926 , RI9143c98_66, \843 );
and \U$109 ( \927 , RI9143518_50, \845 );
and \U$110 ( \928 , RI90f36d0_34, \847 );
and \U$111 ( \929 , RI912e758_18, \849 );
and \U$112 ( \930 , RI9138be0_2, \851 );
or \U$113 ( \931 , \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 );
_DC g3dc ( \932_nG3dc , \931 , \860 );
buf \U$114 ( \933 , \932_nG3dc );
buf \U$115 ( \934 , \933 );
and \U$116 ( \935 , RI9150718_498, \869 );
and \U$117 ( \936 , RI914ff98_482, \871 );
and \U$118 ( \937 , RI914f818_466, \873 );
and \U$119 ( \938 , RI914f098_450, \875 );
and \U$120 ( \939 , RI914e918_434, \877 );
and \U$121 ( \940 , RI914e198_418, \879 );
and \U$122 ( \941 , RI914da18_402, \881 );
and \U$123 ( \942 , RI914d298_386, \883 );
and \U$124 ( \943 , RI914cb18_370, \885 );
and \U$125 ( \944 , RI914c398_354, \887 );
and \U$126 ( \945 , RI914bc18_338, \889 );
and \U$127 ( \946 , RI914b498_322, \891 );
and \U$128 ( \947 , RI914ad18_306, \893 );
and \U$129 ( \948 , RI914a598_290, \895 );
and \U$130 ( \949 , RI9149e18_274, \897 );
and \U$131 ( \950 , RI9149698_258, \899 );
or \U$132 ( \951 , \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 );
_DC g3f0 ( \952_nG3f0 , \951 , \908 );
buf \U$133 ( \953 , \952_nG3f0 );
buf \U$134 ( \954 , \953 );
and \U$135 ( \955 , \934 , \954 );
and \U$136 ( \956 , \914 , \955 );
and \U$137 ( \957 , RI9148ea0_241, \821 );
and \U$138 ( \958 , RI9148720_225, \823 );
and \U$139 ( \959 , RI9147fa0_209, \825 );
and \U$140 ( \960 , RI9147820_193, \827 );
and \U$141 ( \961 , RI91470a0_177, \829 );
and \U$142 ( \962 , RI9146920_161, \831 );
and \U$143 ( \963 , RI91461a0_145, \833 );
and \U$144 ( \964 , RI9145a20_129, \835 );
and \U$145 ( \965 , RI91452a0_113, \837 );
and \U$146 ( \966 , RI9144b20_97, \839 );
and \U$147 ( \967 , RI91443a0_81, \841 );
and \U$148 ( \968 , RI9143c20_65, \843 );
and \U$149 ( \969 , RI91434a0_49, \845 );
and \U$150 ( \970 , RI90f3748_33, \847 );
and \U$151 ( \971 , RI912e7d0_17, \849 );
and \U$152 ( \972 , RI9138c58_1, \851 );
or \U$153 ( \973 , \957 , \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 );
_DC g406 ( \974_nG406 , \973 , \860 );
buf \U$154 ( \975 , \974_nG406 );
buf \U$155 ( \976 , \975 );
not \U$156 ( \977 , \976 );
and \U$157 ( \978 , \977 , \954 );
not \U$158 ( \979 , \954 );
nor \U$159 ( \980 , \978 , \979 );
and \U$160 ( \981 , \956 , \980 );
not \U$161 ( \982 , \934 );
and \U$162 ( \983 , \912 , \934 );
nor \U$163 ( \984 , \982 , \983 );
xor \U$164 ( \985 , \956 , \980 );
and \U$165 ( \986 , \984 , \985 );
and \U$167 ( \987 , \976 , \911 );
and \U$168 ( \988 , \986 , \987 );
and \U$169 ( \989 , \981 , \987 );
or \U$170 ( \990 , 1'b0 , \988 , \989 );
xor \U$171 ( \991 , \981 , \986 );
xor \U$172 ( \992 , \991 , \987 );
and \U$173 ( \993 , RI9149008_244, \821 );
and \U$174 ( \994 , RI9148888_228, \823 );
and \U$175 ( \995 , RI9148108_212, \825 );
and \U$176 ( \996 , RI9147988_196, \827 );
and \U$177 ( \997 , RI9147208_180, \829 );
and \U$178 ( \998 , RI9146a88_164, \831 );
and \U$179 ( \999 , RI9146308_148, \833 );
and \U$180 ( \1000 , RI9145b88_132, \835 );
and \U$181 ( \1001 , RI9145408_116, \837 );
and \U$182 ( \1002 , RI9144c88_100, \839 );
and \U$183 ( \1003 , RI9144508_84, \841 );
and \U$184 ( \1004 , RI9143d88_68, \843 );
and \U$185 ( \1005 , RI9143608_52, \845 );
and \U$186 ( \1006 , RI90f35e0_36, \847 );
and \U$187 ( \1007 , RI90f9940_20, \849 );
and \U$188 ( \1008 , RI9138af0_4, \851 );
or \U$189 ( \1009 , \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 );
_DC g42b ( \1010_nG42b , \1009 , \860 );
buf \U$190 ( \1011 , \1010_nG42b );
buf \U$191 ( \1012 , \1011 );
not \U$192 ( \1013 , \1012 );
and \U$193 ( \1014 , \912 , \1012 );
nor \U$194 ( \1015 , \1013 , \1014 );
and \U$195 ( \1016 , \863 , \954 );
and \U$196 ( \1017 , \1015 , \1016 );
and \U$197 ( \1018 , RI9150790_499, \869 );
and \U$198 ( \1019 , RI9150010_483, \871 );
and \U$199 ( \1020 , RI914f890_467, \873 );
and \U$200 ( \1021 , RI914f110_451, \875 );
and \U$201 ( \1022 , RI914e990_435, \877 );
and \U$202 ( \1023 , RI914e210_419, \879 );
and \U$203 ( \1024 , RI914da90_403, \881 );
and \U$204 ( \1025 , RI914d310_387, \883 );
and \U$205 ( \1026 , RI914cb90_371, \885 );
and \U$206 ( \1027 , RI914c410_355, \887 );
and \U$207 ( \1028 , RI914bc90_339, \889 );
and \U$208 ( \1029 , RI914b510_323, \891 );
and \U$209 ( \1030 , RI914ad90_307, \893 );
and \U$210 ( \1031 , RI914a610_291, \895 );
and \U$211 ( \1032 , RI9149e90_275, \897 );
and \U$212 ( \1033 , RI9149710_259, \899 );
or \U$213 ( \1034 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 );
_DC g444 ( \1035_nG444 , \1034 , \908 );
buf \U$214 ( \1036 , \1035_nG444 );
buf \U$215 ( \1037 , \1036 );
and \U$216 ( \1038 , \934 , \1037 );
and \U$217 ( \1039 , \1016 , \1038 );
and \U$218 ( \1040 , \1015 , \1038 );
or \U$219 ( \1041 , \1017 , \1039 , \1040 );
and \U$220 ( \1042 , RI91490f8_246, \821 );
and \U$221 ( \1043 , RI9148978_230, \823 );
and \U$222 ( \1044 , RI91481f8_214, \825 );
and \U$223 ( \1045 , RI9147a78_198, \827 );
and \U$224 ( \1046 , RI91472f8_182, \829 );
and \U$225 ( \1047 , RI9146b78_166, \831 );
and \U$226 ( \1048 , RI91463f8_150, \833 );
and \U$227 ( \1049 , RI9145c78_134, \835 );
and \U$228 ( \1050 , RI91454f8_118, \837 );
and \U$229 ( \1051 , RI9144d78_102, \839 );
and \U$230 ( \1052 , RI91445f8_86, \841 );
and \U$231 ( \1053 , RI9143e78_70, \843 );
and \U$232 ( \1054 , RI91436f8_54, \845 );
and \U$233 ( \1055 , RI90f34f0_38, \847 );
and \U$234 ( \1056 , RI90f9850_22, \849 );
and \U$235 ( \1057 , RI9138a00_6, \851 );
or \U$236 ( \1058 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 );
_DC g45c ( \1059_nG45c , \1058 , \860 );
buf \U$237 ( \1060 , \1059_nG45c );
buf \U$238 ( \1061 , \1060 );
not \U$239 ( \1062 , \1061 );
and \U$240 ( \1063 , \912 , \1061 );
nor \U$241 ( \1064 , \1062 , \1063 );
and \U$242 ( \1065 , RI9149080_245, \821 );
and \U$243 ( \1066 , RI9148900_229, \823 );
and \U$244 ( \1067 , RI9148180_213, \825 );
and \U$245 ( \1068 , RI9147a00_197, \827 );
and \U$246 ( \1069 , RI9147280_181, \829 );
and \U$247 ( \1070 , RI9146b00_165, \831 );
and \U$248 ( \1071 , RI9146380_149, \833 );
and \U$249 ( \1072 , RI9145c00_133, \835 );
and \U$250 ( \1073 , RI9145480_117, \837 );
and \U$251 ( \1074 , RI9144d00_101, \839 );
and \U$252 ( \1075 , RI9144580_85, \841 );
and \U$253 ( \1076 , RI9143e00_69, \843 );
and \U$254 ( \1077 , RI9143680_53, \845 );
and \U$255 ( \1078 , RI90f3568_37, \847 );
and \U$256 ( \1079 , RI90f98c8_21, \849 );
and \U$257 ( \1080 , RI9138a78_5, \851 );
or \U$258 ( \1081 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 );
_DC g473 ( \1082_nG473 , \1081 , \860 );
buf \U$259 ( \1083 , \1082_nG473 );
buf \U$260 ( \1084 , \1083 );
and \U$261 ( \1085 , \1084 , \954 );
and \U$262 ( \1086 , \1064 , \1085 );
not \U$263 ( \1087 , \1084 );
and \U$264 ( \1088 , \912 , \1084 );
nor \U$265 ( \1089 , \1087 , \1088 );
and \U$266 ( \1090 , \1086 , \1089 );
and \U$267 ( \1091 , \1012 , \954 );
and \U$268 ( \1092 , \863 , \1037 );
xor \U$269 ( \1093 , \1091 , \1092 );
and \U$270 ( \1094 , RI9150808_500, \869 );
and \U$271 ( \1095 , RI9150088_484, \871 );
and \U$272 ( \1096 , RI914f908_468, \873 );
and \U$273 ( \1097 , RI914f188_452, \875 );
and \U$274 ( \1098 , RI914ea08_436, \877 );
and \U$275 ( \1099 , RI914e288_420, \879 );
and \U$276 ( \1100 , RI914db08_404, \881 );
and \U$277 ( \1101 , RI914d388_388, \883 );
and \U$278 ( \1102 , RI914cc08_372, \885 );
and \U$279 ( \1103 , RI914c488_356, \887 );
and \U$280 ( \1104 , RI914bd08_340, \889 );
and \U$281 ( \1105 , RI914b588_324, \891 );
and \U$282 ( \1106 , RI914ae08_308, \893 );
and \U$283 ( \1107 , RI914a688_292, \895 );
and \U$284 ( \1108 , RI9149f08_276, \897 );
and \U$285 ( \1109 , RI9149788_260, \899 );
or \U$286 ( \1110 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 );
_DC g490 ( \1111_nG490 , \1110 , \908 );
buf \U$287 ( \1112 , \1111_nG490 );
buf \U$288 ( \1113 , \1112 );
and \U$289 ( \1114 , \934 , \1113 );
xor \U$290 ( \1115 , \1093 , \1114 );
and \U$291 ( \1116 , \1089 , \1115 );
and \U$292 ( \1117 , \1086 , \1115 );
or \U$293 ( \1118 , \1090 , \1116 , \1117 );
xor \U$294 ( \1119 , \1015 , \1016 );
xor \U$295 ( \1120 , \1119 , \1038 );
and \U$296 ( \1121 , \1118 , \1120 );
and \U$297 ( \1122 , \1041 , \1121 );
and \U$298 ( \1123 , \977 , \1037 );
not \U$299 ( \1124 , \1037 );
nor \U$300 ( \1125 , \1123 , \1124 );
and \U$301 ( \1126 , \1121 , \1125 );
and \U$302 ( \1127 , \1041 , \1125 );
or \U$303 ( \1128 , \1122 , \1126 , \1127 );
xor \U$304 ( \1129 , \1041 , \1121 );
xor \U$305 ( \1130 , \1129 , \1125 );
xor \U$306 ( \1131 , \914 , \955 );
and \U$307 ( \1132 , \1130 , \1131 );
and \U$308 ( \1133 , \1128 , \1132 );
xor \U$309 ( \1134 , \984 , \985 );
and \U$310 ( \1135 , \1132 , \1134 );
and \U$311 ( \1136 , \1128 , \1134 );
or \U$312 ( \1137 , \1133 , \1135 , \1136 );
and \U$313 ( \1138 , \992 , \1137 );
xor \U$314 ( \1139 , \992 , \1137 );
xor \U$315 ( \1140 , \1128 , \1132 );
xor \U$316 ( \1141 , \1140 , \1134 );
and \U$317 ( \1142 , \1091 , \1092 );
and \U$318 ( \1143 , \1092 , \1114 );
and \U$319 ( \1144 , \1091 , \1114 );
or \U$320 ( \1145 , \1142 , \1143 , \1144 );
and \U$321 ( \1146 , RI9149170_247, \821 );
and \U$322 ( \1147 , RI91489f0_231, \823 );
and \U$323 ( \1148 , RI9148270_215, \825 );
and \U$324 ( \1149 , RI9147af0_199, \827 );
and \U$325 ( \1150 , RI9147370_183, \829 );
and \U$326 ( \1151 , RI9146bf0_167, \831 );
and \U$327 ( \1152 , RI9146470_151, \833 );
and \U$328 ( \1153 , RI9145cf0_135, \835 );
and \U$329 ( \1154 , RI9145570_119, \837 );
and \U$330 ( \1155 , RI9144df0_103, \839 );
and \U$331 ( \1156 , RI9144670_87, \841 );
and \U$332 ( \1157 , RI9143ef0_71, \843 );
and \U$333 ( \1158 , RI9143770_55, \845 );
and \U$334 ( \1159 , RI90f3478_39, \847 );
and \U$335 ( \1160 , RI90f97d8_23, \849 );
and \U$336 ( \1161 , RI9138988_7, \851 );
or \U$337 ( \1162 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 );
_DC g4c4 ( \1163_nG4c4 , \1162 , \860 );
buf \U$338 ( \1164 , \1163_nG4c4 );
buf \U$339 ( \1165 , \1164 );
not \U$340 ( \1166 , \1165 );
and \U$341 ( \1167 , \912 , \1165 );
nor \U$342 ( \1168 , \1166 , \1167 );
and \U$343 ( \1169 , \1061 , \954 );
and \U$344 ( \1170 , \1168 , \1169 );
and \U$345 ( \1171 , \1084 , \1037 );
and \U$346 ( \1172 , \1169 , \1171 );
and \U$347 ( \1173 , \1168 , \1171 );
or \U$348 ( \1174 , \1170 , \1172 , \1173 );
and \U$349 ( \1175 , \1012 , \1037 );
and \U$350 ( \1176 , \863 , \1113 );
xor \U$351 ( \1177 , \1175 , \1176 );
and \U$352 ( \1178 , RI9150880_501, \869 );
and \U$353 ( \1179 , RI9150100_485, \871 );
and \U$354 ( \1180 , RI914f980_469, \873 );
and \U$355 ( \1181 , RI914f200_453, \875 );
and \U$356 ( \1182 , RI914ea80_437, \877 );
and \U$357 ( \1183 , RI914e300_421, \879 );
and \U$358 ( \1184 , RI914db80_405, \881 );
and \U$359 ( \1185 , RI914d400_389, \883 );
and \U$360 ( \1186 , RI914cc80_373, \885 );
and \U$361 ( \1187 , RI914c500_357, \887 );
and \U$362 ( \1188 , RI914bd80_341, \889 );
and \U$363 ( \1189 , RI914b600_325, \891 );
and \U$364 ( \1190 , RI914ae80_309, \893 );
and \U$365 ( \1191 , RI914a700_293, \895 );
and \U$366 ( \1192 , RI9149f80_277, \897 );
and \U$367 ( \1193 , RI9149800_261, \899 );
or \U$368 ( \1194 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 );
_DC g4e4 ( \1195_nG4e4 , \1194 , \908 );
buf \U$369 ( \1196 , \1195_nG4e4 );
buf \U$370 ( \1197 , \1196 );
and \U$371 ( \1198 , \934 , \1197 );
xor \U$372 ( \1199 , \1177 , \1198 );
and \U$373 ( \1200 , \1174 , \1199 );
xor \U$374 ( \1201 , \1064 , \1085 );
and \U$375 ( \1202 , \1199 , \1201 );
and \U$376 ( \1203 , \1174 , \1201 );
or \U$377 ( \1204 , \1200 , \1202 , \1203 );
xor \U$378 ( \1205 , \1086 , \1089 );
xor \U$379 ( \1206 , \1205 , \1115 );
and \U$380 ( \1207 , \1204 , \1206 );
and \U$381 ( \1208 , \1145 , \1207 );
and \U$382 ( \1209 , \977 , \1113 );
not \U$383 ( \1210 , \1113 );
nor \U$384 ( \1211 , \1209 , \1210 );
and \U$385 ( \1212 , \1207 , \1211 );
and \U$386 ( \1213 , \1145 , \1211 );
or \U$387 ( \1214 , \1208 , \1212 , \1213 );
xor \U$388 ( \1215 , \1145 , \1207 );
xor \U$389 ( \1216 , \1215 , \1211 );
xor \U$390 ( \1217 , \1118 , \1120 );
and \U$391 ( \1218 , \1216 , \1217 );
and \U$392 ( \1219 , \1214 , \1218 );
xor \U$393 ( \1220 , \1130 , \1131 );
and \U$394 ( \1221 , \1218 , \1220 );
and \U$395 ( \1222 , \1214 , \1220 );
or \U$396 ( \1223 , \1219 , \1221 , \1222 );
and \U$397 ( \1224 , \1141 , \1223 );
xor \U$398 ( \1225 , \1141 , \1223 );
xor \U$399 ( \1226 , \1214 , \1218 );
xor \U$400 ( \1227 , \1226 , \1220 );
and \U$401 ( \1228 , \1175 , \1176 );
and \U$402 ( \1229 , \1176 , \1198 );
and \U$403 ( \1230 , \1175 , \1198 );
or \U$404 ( \1231 , \1228 , \1229 , \1230 );
and \U$405 ( \1232 , \1165 , \954 );
and \U$406 ( \1233 , \1061 , \1037 );
and \U$407 ( \1234 , \1232 , \1233 );
and \U$408 ( \1235 , \1084 , \1113 );
and \U$409 ( \1236 , \1233 , \1235 );
and \U$410 ( \1237 , \1232 , \1235 );
or \U$411 ( \1238 , \1234 , \1236 , \1237 );
and \U$412 ( \1239 , \1012 , \1113 );
and \U$413 ( \1240 , \863 , \1197 );
xor \U$414 ( \1241 , \1239 , \1240 );
and \U$415 ( \1242 , RI91508f8_502, \869 );
and \U$416 ( \1243 , RI9150178_486, \871 );
and \U$417 ( \1244 , RI914f9f8_470, \873 );
and \U$418 ( \1245 , RI914f278_454, \875 );
and \U$419 ( \1246 , RI914eaf8_438, \877 );
and \U$420 ( \1247 , RI914e378_422, \879 );
and \U$421 ( \1248 , RI914dbf8_406, \881 );
and \U$422 ( \1249 , RI914d478_390, \883 );
and \U$423 ( \1250 , RI914ccf8_374, \885 );
and \U$424 ( \1251 , RI914c578_358, \887 );
and \U$425 ( \1252 , RI914bdf8_342, \889 );
and \U$426 ( \1253 , RI914b678_326, \891 );
and \U$427 ( \1254 , RI914aef8_310, \893 );
and \U$428 ( \1255 , RI914a778_294, \895 );
and \U$429 ( \1256 , RI9149ff8_278, \897 );
and \U$430 ( \1257 , RI9149878_262, \899 );
or \U$431 ( \1258 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 );
_DC g524 ( \1259_nG524 , \1258 , \908 );
buf \U$432 ( \1260 , \1259_nG524 );
buf \U$433 ( \1261 , \1260 );
and \U$434 ( \1262 , \934 , \1261 );
xor \U$435 ( \1263 , \1241 , \1262 );
and \U$436 ( \1264 , \1238 , \1263 );
xor \U$437 ( \1265 , \1168 , \1169 );
xor \U$438 ( \1266 , \1265 , \1171 );
and \U$439 ( \1267 , \1263 , \1266 );
and \U$440 ( \1268 , \1238 , \1266 );
or \U$441 ( \1269 , \1264 , \1267 , \1268 );
xor \U$442 ( \1270 , \1174 , \1199 );
xor \U$443 ( \1271 , \1270 , \1201 );
and \U$444 ( \1272 , \1269 , \1271 );
and \U$445 ( \1273 , \1231 , \1272 );
and \U$446 ( \1274 , \977 , \1197 );
not \U$447 ( \1275 , \1197 );
nor \U$448 ( \1276 , \1274 , \1275 );
and \U$449 ( \1277 , \1272 , \1276 );
and \U$450 ( \1278 , \1231 , \1276 );
or \U$451 ( \1279 , \1273 , \1277 , \1278 );
xor \U$452 ( \1280 , \1231 , \1272 );
xor \U$453 ( \1281 , \1280 , \1276 );
xor \U$454 ( \1282 , \1204 , \1206 );
and \U$455 ( \1283 , \1281 , \1282 );
and \U$456 ( \1284 , \1279 , \1283 );
xor \U$457 ( \1285 , \1216 , \1217 );
and \U$458 ( \1286 , \1283 , \1285 );
and \U$459 ( \1287 , \1279 , \1285 );
or \U$460 ( \1288 , \1284 , \1286 , \1287 );
and \U$461 ( \1289 , \1227 , \1288 );
xor \U$462 ( \1290 , \1227 , \1288 );
xor \U$463 ( \1291 , \1279 , \1283 );
xor \U$464 ( \1292 , \1291 , \1285 );
and \U$465 ( \1293 , \1239 , \1240 );
and \U$466 ( \1294 , \1240 , \1262 );
and \U$467 ( \1295 , \1239 , \1262 );
or \U$468 ( \1296 , \1293 , \1294 , \1295 );
and \U$469 ( \1297 , \1165 , \1037 );
and \U$470 ( \1298 , \1061 , \1113 );
and \U$471 ( \1299 , \1297 , \1298 );
and \U$472 ( \1300 , \1084 , \1197 );
and \U$473 ( \1301 , \1298 , \1300 );
and \U$474 ( \1302 , \1297 , \1300 );
or \U$475 ( \1303 , \1299 , \1301 , \1302 );
and \U$476 ( \1304 , \1012 , \1197 );
and \U$477 ( \1305 , \863 , \1261 );
xor \U$478 ( \1306 , \1304 , \1305 );
and \U$479 ( \1307 , RI9150970_503, \869 );
and \U$480 ( \1308 , RI91501f0_487, \871 );
and \U$481 ( \1309 , RI914fa70_471, \873 );
and \U$482 ( \1310 , RI914f2f0_455, \875 );
and \U$483 ( \1311 , RI914eb70_439, \877 );
and \U$484 ( \1312 , RI914e3f0_423, \879 );
and \U$485 ( \1313 , RI914dc70_407, \881 );
and \U$486 ( \1314 , RI914d4f0_391, \883 );
and \U$487 ( \1315 , RI914cd70_375, \885 );
and \U$488 ( \1316 , RI914c5f0_359, \887 );
and \U$489 ( \1317 , RI914be70_343, \889 );
and \U$490 ( \1318 , RI914b6f0_327, \891 );
and \U$491 ( \1319 , RI914af70_311, \893 );
and \U$492 ( \1320 , RI914a7f0_295, \895 );
and \U$493 ( \1321 , RI914a070_279, \897 );
and \U$494 ( \1322 , RI91498f0_263, \899 );
or \U$495 ( \1323 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 );
_DC g565 ( \1324_nG565 , \1323 , \908 );
buf \U$496 ( \1325 , \1324_nG565 );
buf \U$497 ( \1326 , \1325 );
and \U$498 ( \1327 , \934 , \1326 );
xor \U$499 ( \1328 , \1306 , \1327 );
and \U$500 ( \1329 , \1303 , \1328 );
xor \U$501 ( \1330 , \1232 , \1233 );
xor \U$502 ( \1331 , \1330 , \1235 );
and \U$503 ( \1332 , \1328 , \1331 );
and \U$504 ( \1333 , \1303 , \1331 );
or \U$505 ( \1334 , \1329 , \1332 , \1333 );
and \U$506 ( \1335 , RI9149260_249, \821 );
and \U$507 ( \1336 , RI9148ae0_233, \823 );
and \U$508 ( \1337 , RI9148360_217, \825 );
and \U$509 ( \1338 , RI9147be0_201, \827 );
and \U$510 ( \1339 , RI9147460_185, \829 );
and \U$511 ( \1340 , RI9146ce0_169, \831 );
and \U$512 ( \1341 , RI9146560_153, \833 );
and \U$513 ( \1342 , RI9145de0_137, \835 );
and \U$514 ( \1343 , RI9145660_121, \837 );
and \U$515 ( \1344 , RI9144ee0_105, \839 );
and \U$516 ( \1345 , RI9144760_89, \841 );
and \U$517 ( \1346 , RI9143fe0_73, \843 );
and \U$518 ( \1347 , RI9143860_57, \845 );
and \U$519 ( \1348 , RI90f3388_41, \847 );
and \U$520 ( \1349 , RI90f96e8_25, \849 );
and \U$521 ( \1350 , RI9138898_9, \851 );
or \U$522 ( \1351 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 );
_DC g581 ( \1352_nG581 , \1351 , \860 );
buf \U$523 ( \1353 , \1352_nG581 );
buf \U$524 ( \1354 , \1353 );
not \U$525 ( \1355 , \1354 );
and \U$526 ( \1356 , \912 , \1354 );
nor \U$527 ( \1357 , \1355 , \1356 );
and \U$528 ( \1358 , RI91491e8_248, \821 );
and \U$529 ( \1359 , RI9148a68_232, \823 );
and \U$530 ( \1360 , RI91482e8_216, \825 );
and \U$531 ( \1361 , RI9147b68_200, \827 );
and \U$532 ( \1362 , RI91473e8_184, \829 );
and \U$533 ( \1363 , RI9146c68_168, \831 );
and \U$534 ( \1364 , RI91464e8_152, \833 );
and \U$535 ( \1365 , RI9145d68_136, \835 );
and \U$536 ( \1366 , RI91455e8_120, \837 );
and \U$537 ( \1367 , RI9144e68_104, \839 );
and \U$538 ( \1368 , RI91446e8_88, \841 );
and \U$539 ( \1369 , RI9143f68_72, \843 );
and \U$540 ( \1370 , RI91437e8_56, \845 );
and \U$541 ( \1371 , RI90f3400_40, \847 );
and \U$542 ( \1372 , RI90f9760_24, \849 );
and \U$543 ( \1373 , RI9138910_8, \851 );
or \U$544 ( \1374 , \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 );
_DC g598 ( \1375_nG598 , \1374 , \860 );
buf \U$545 ( \1376 , \1375_nG598 );
buf \U$546 ( \1377 , \1376 );
and \U$547 ( \1378 , \1377 , \954 );
and \U$548 ( \1379 , \1357 , \1378 );
not \U$549 ( \1380 , \1377 );
and \U$550 ( \1381 , \912 , \1377 );
nor \U$551 ( \1382 , \1380 , \1381 );
and \U$552 ( \1383 , \1379 , \1382 );
and \U$553 ( \1384 , \1334 , \1383 );
xor \U$554 ( \1385 , \1238 , \1263 );
xor \U$555 ( \1386 , \1385 , \1266 );
and \U$556 ( \1387 , \1383 , \1386 );
and \U$557 ( \1388 , \1334 , \1386 );
or \U$558 ( \1389 , \1384 , \1387 , \1388 );
and \U$559 ( \1390 , \1296 , \1389 );
and \U$560 ( \1391 , \977 , \1261 );
not \U$561 ( \1392 , \1261 );
nor \U$562 ( \1393 , \1391 , \1392 );
and \U$563 ( \1394 , \1389 , \1393 );
and \U$564 ( \1395 , \1296 , \1393 );
or \U$565 ( \1396 , \1390 , \1394 , \1395 );
xor \U$566 ( \1397 , \1296 , \1389 );
xor \U$567 ( \1398 , \1397 , \1393 );
xor \U$568 ( \1399 , \1269 , \1271 );
and \U$569 ( \1400 , \1398 , \1399 );
and \U$570 ( \1401 , \1396 , \1400 );
xor \U$571 ( \1402 , \1281 , \1282 );
and \U$572 ( \1403 , \1400 , \1402 );
and \U$573 ( \1404 , \1396 , \1402 );
or \U$574 ( \1405 , \1401 , \1403 , \1404 );
and \U$575 ( \1406 , \1292 , \1405 );
xor \U$576 ( \1407 , \1292 , \1405 );
xor \U$577 ( \1408 , \1396 , \1400 );
xor \U$578 ( \1409 , \1408 , \1402 );
and \U$579 ( \1410 , \1304 , \1305 );
and \U$580 ( \1411 , \1305 , \1327 );
and \U$581 ( \1412 , \1304 , \1327 );
or \U$582 ( \1413 , \1410 , \1411 , \1412 );
and \U$583 ( \1414 , \1165 , \1113 );
and \U$584 ( \1415 , \1061 , \1197 );
and \U$585 ( \1416 , \1414 , \1415 );
and \U$586 ( \1417 , \1084 , \1261 );
and \U$587 ( \1418 , \1415 , \1417 );
and \U$588 ( \1419 , \1414 , \1417 );
or \U$589 ( \1420 , \1416 , \1418 , \1419 );
xor \U$590 ( \1421 , \1297 , \1298 );
xor \U$591 ( \1422 , \1421 , \1300 );
and \U$592 ( \1423 , \1420 , \1422 );
and \U$593 ( \1424 , \1012 , \1261 );
and \U$594 ( \1425 , \863 , \1326 );
xor \U$595 ( \1426 , \1424 , \1425 );
and \U$596 ( \1427 , RI91509e8_504, \869 );
and \U$597 ( \1428 , RI9150268_488, \871 );
and \U$598 ( \1429 , RI914fae8_472, \873 );
and \U$599 ( \1430 , RI914f368_456, \875 );
and \U$600 ( \1431 , RI914ebe8_440, \877 );
and \U$601 ( \1432 , RI914e468_424, \879 );
and \U$602 ( \1433 , RI914dce8_408, \881 );
and \U$603 ( \1434 , RI914d568_392, \883 );
and \U$604 ( \1435 , RI914cde8_376, \885 );
and \U$605 ( \1436 , RI914c668_360, \887 );
and \U$606 ( \1437 , RI914bee8_344, \889 );
and \U$607 ( \1438 , RI914b768_328, \891 );
and \U$608 ( \1439 , RI914afe8_312, \893 );
and \U$609 ( \1440 , RI914a868_296, \895 );
and \U$610 ( \1441 , RI914a0e8_280, \897 );
and \U$611 ( \1442 , RI9149968_264, \899 );
or \U$612 ( \1443 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 );
_DC g5dd ( \1444_nG5dd , \1443 , \908 );
buf \U$613 ( \1445 , \1444_nG5dd );
buf \U$614 ( \1446 , \1445 );
and \U$615 ( \1447 , \934 , \1446 );
xor \U$616 ( \1448 , \1426 , \1447 );
and \U$617 ( \1449 , \1422 , \1448 );
and \U$618 ( \1450 , \1420 , \1448 );
or \U$619 ( \1451 , \1423 , \1449 , \1450 );
and \U$620 ( \1452 , RI91492d8_250, \821 );
and \U$621 ( \1453 , RI9148b58_234, \823 );
and \U$622 ( \1454 , RI91483d8_218, \825 );
and \U$623 ( \1455 , RI9147c58_202, \827 );
and \U$624 ( \1456 , RI91474d8_186, \829 );
and \U$625 ( \1457 , RI9146d58_170, \831 );
and \U$626 ( \1458 , RI91465d8_154, \833 );
and \U$627 ( \1459 , RI9145e58_138, \835 );
and \U$628 ( \1460 , RI91456d8_122, \837 );
and \U$629 ( \1461 , RI9144f58_106, \839 );
and \U$630 ( \1462 , RI91447d8_90, \841 );
and \U$631 ( \1463 , RI9144058_74, \843 );
and \U$632 ( \1464 , RI91438d8_58, \845 );
and \U$633 ( \1465 , RI90f3310_42, \847 );
and \U$634 ( \1466 , RI90f9670_26, \849 );
and \U$635 ( \1467 , RI912eb18_10, \851 );
or \U$636 ( \1468 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 );
_DC g5f6 ( \1469_nG5f6 , \1468 , \860 );
buf \U$637 ( \1470 , \1469_nG5f6 );
buf \U$638 ( \1471 , \1470 );
not \U$639 ( \1472 , \1471 );
and \U$640 ( \1473 , \912 , \1471 );
nor \U$641 ( \1474 , \1472 , \1473 );
and \U$642 ( \1475 , \1354 , \954 );
and \U$643 ( \1476 , \1474 , \1475 );
and \U$644 ( \1477 , \1377 , \1037 );
and \U$645 ( \1478 , \1475 , \1477 );
and \U$646 ( \1479 , \1474 , \1477 );
or \U$647 ( \1480 , \1476 , \1478 , \1479 );
xor \U$648 ( \1481 , \1357 , \1378 );
and \U$649 ( \1482 , \1480 , \1481 );
and \U$650 ( \1483 , \1451 , \1482 );
xor \U$651 ( \1484 , \1303 , \1328 );
xor \U$652 ( \1485 , \1484 , \1331 );
and \U$653 ( \1486 , \1482 , \1485 );
and \U$654 ( \1487 , \1451 , \1485 );
or \U$655 ( \1488 , \1483 , \1486 , \1487 );
and \U$656 ( \1489 , \1413 , \1488 );
and \U$657 ( \1490 , \977 , \1326 );
not \U$658 ( \1491 , \1326 );
nor \U$659 ( \1492 , \1490 , \1491 );
and \U$660 ( \1493 , \1488 , \1492 );
and \U$661 ( \1494 , \1413 , \1492 );
or \U$662 ( \1495 , \1489 , \1493 , \1494 );
xor \U$663 ( \1496 , \1451 , \1482 );
xor \U$664 ( \1497 , \1496 , \1485 );
xor \U$665 ( \1498 , \1379 , \1382 );
and \U$666 ( \1499 , \1497 , \1498 );
xor \U$667 ( \1500 , \1413 , \1488 );
xor \U$668 ( \1501 , \1500 , \1492 );
and \U$669 ( \1502 , \1499 , \1501 );
xor \U$670 ( \1503 , \1334 , \1383 );
xor \U$671 ( \1504 , \1503 , \1386 );
and \U$672 ( \1505 , \1501 , \1504 );
and \U$673 ( \1506 , \1499 , \1504 );
or \U$674 ( \1507 , \1502 , \1505 , \1506 );
and \U$675 ( \1508 , \1495 , \1507 );
xor \U$676 ( \1509 , \1398 , \1399 );
and \U$677 ( \1510 , \1507 , \1509 );
and \U$678 ( \1511 , \1495 , \1509 );
or \U$679 ( \1512 , \1508 , \1510 , \1511 );
and \U$680 ( \1513 , \1409 , \1512 );
xor \U$681 ( \1514 , \1409 , \1512 );
xor \U$682 ( \1515 , \1495 , \1507 );
xor \U$683 ( \1516 , \1515 , \1509 );
and \U$684 ( \1517 , \1424 , \1425 );
and \U$685 ( \1518 , \1425 , \1447 );
and \U$686 ( \1519 , \1424 , \1447 );
or \U$687 ( \1520 , \1517 , \1518 , \1519 );
and \U$688 ( \1521 , \1165 , \1197 );
and \U$689 ( \1522 , \1061 , \1261 );
and \U$690 ( \1523 , \1521 , \1522 );
and \U$691 ( \1524 , \1084 , \1326 );
and \U$692 ( \1525 , \1522 , \1524 );
and \U$693 ( \1526 , \1521 , \1524 );
or \U$694 ( \1527 , \1523 , \1525 , \1526 );
and \U$695 ( \1528 , \1012 , \1326 );
and \U$696 ( \1529 , \863 , \1446 );
xor \U$697 ( \1530 , \1528 , \1529 );
and \U$698 ( \1531 , RI9150a60_505, \869 );
and \U$699 ( \1532 , RI91502e0_489, \871 );
and \U$700 ( \1533 , RI914fb60_473, \873 );
and \U$701 ( \1534 , RI914f3e0_457, \875 );
and \U$702 ( \1535 , RI914ec60_441, \877 );
and \U$703 ( \1536 , RI914e4e0_425, \879 );
and \U$704 ( \1537 , RI914dd60_409, \881 );
and \U$705 ( \1538 , RI914d5e0_393, \883 );
and \U$706 ( \1539 , RI914ce60_377, \885 );
and \U$707 ( \1540 , RI914c6e0_361, \887 );
and \U$708 ( \1541 , RI914bf60_345, \889 );
and \U$709 ( \1542 , RI914b7e0_329, \891 );
and \U$710 ( \1543 , RI914b060_313, \893 );
and \U$711 ( \1544 , RI914a8e0_297, \895 );
and \U$712 ( \1545 , RI914a160_281, \897 );
and \U$713 ( \1546 , RI91499e0_265, \899 );
or \U$714 ( \1547 , \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 , \1546 );
_DC g645 ( \1548_nG645 , \1547 , \908 );
buf \U$715 ( \1549 , \1548_nG645 );
buf \U$716 ( \1550 , \1549 );
and \U$717 ( \1551 , \934 , \1550 );
xor \U$718 ( \1552 , \1530 , \1551 );
and \U$719 ( \1553 , \1527 , \1552 );
xor \U$720 ( \1554 , \1414 , \1415 );
xor \U$721 ( \1555 , \1554 , \1417 );
and \U$722 ( \1556 , \1552 , \1555 );
and \U$723 ( \1557 , \1527 , \1555 );
or \U$724 ( \1558 , \1553 , \1556 , \1557 );
and \U$725 ( \1559 , \1471 , \954 );
and \U$726 ( \1560 , \1354 , \1037 );
and \U$727 ( \1561 , \1559 , \1560 );
and \U$728 ( \1562 , \1377 , \1113 );
and \U$729 ( \1563 , \1560 , \1562 );
and \U$730 ( \1564 , \1559 , \1562 );
or \U$731 ( \1565 , \1561 , \1563 , \1564 );
xor \U$732 ( \1566 , \1474 , \1475 );
xor \U$733 ( \1567 , \1566 , \1477 );
and \U$734 ( \1568 , \1565 , \1567 );
and \U$735 ( \1569 , \1558 , \1568 );
xor \U$736 ( \1570 , \1420 , \1422 );
xor \U$737 ( \1571 , \1570 , \1448 );
and \U$738 ( \1572 , \1568 , \1571 );
and \U$739 ( \1573 , \1558 , \1571 );
or \U$740 ( \1574 , \1569 , \1572 , \1573 );
and \U$741 ( \1575 , \1520 , \1574 );
and \U$742 ( \1576 , \977 , \1446 );
not \U$743 ( \1577 , \1446 );
nor \U$744 ( \1578 , \1576 , \1577 );
and \U$745 ( \1579 , \1574 , \1578 );
and \U$746 ( \1580 , \1520 , \1578 );
or \U$747 ( \1581 , \1575 , \1579 , \1580 );
xor \U$748 ( \1582 , \1558 , \1568 );
xor \U$749 ( \1583 , \1582 , \1571 );
xor \U$750 ( \1584 , \1480 , \1481 );
and \U$751 ( \1585 , \1583 , \1584 );
xor \U$752 ( \1586 , \1520 , \1574 );
xor \U$753 ( \1587 , \1586 , \1578 );
and \U$754 ( \1588 , \1585 , \1587 );
xor \U$755 ( \1589 , \1497 , \1498 );
and \U$756 ( \1590 , \1587 , \1589 );
and \U$757 ( \1591 , \1585 , \1589 );
or \U$758 ( \1592 , \1588 , \1590 , \1591 );
and \U$759 ( \1593 , \1581 , \1592 );
xor \U$760 ( \1594 , \1499 , \1501 );
xor \U$761 ( \1595 , \1594 , \1504 );
and \U$762 ( \1596 , \1592 , \1595 );
and \U$763 ( \1597 , \1581 , \1595 );
or \U$764 ( \1598 , \1593 , \1596 , \1597 );
and \U$765 ( \1599 , \1516 , \1598 );
xor \U$766 ( \1600 , \1516 , \1598 );
xor \U$767 ( \1601 , \1581 , \1592 );
xor \U$768 ( \1602 , \1601 , \1595 );
and \U$769 ( \1603 , \1528 , \1529 );
and \U$770 ( \1604 , \1529 , \1551 );
and \U$771 ( \1605 , \1528 , \1551 );
or \U$772 ( \1606 , \1603 , \1604 , \1605 );
and \U$773 ( \1607 , \1471 , \1037 );
and \U$774 ( \1608 , \1354 , \1113 );
and \U$775 ( \1609 , \1607 , \1608 );
and \U$776 ( \1610 , \1377 , \1197 );
and \U$777 ( \1611 , \1608 , \1610 );
and \U$778 ( \1612 , \1607 , \1610 );
or \U$779 ( \1613 , \1609 , \1611 , \1612 );
and \U$780 ( \1614 , RI91493c8_252, \821 );
and \U$781 ( \1615 , RI9148c48_236, \823 );
and \U$782 ( \1616 , RI91484c8_220, \825 );
and \U$783 ( \1617 , RI9147d48_204, \827 );
and \U$784 ( \1618 , RI91475c8_188, \829 );
and \U$785 ( \1619 , RI9146e48_172, \831 );
and \U$786 ( \1620 , RI91466c8_156, \833 );
and \U$787 ( \1621 , RI9145f48_140, \835 );
and \U$788 ( \1622 , RI91457c8_124, \837 );
and \U$789 ( \1623 , RI9145048_108, \839 );
and \U$790 ( \1624 , RI91448c8_92, \841 );
and \U$791 ( \1625 , RI9144148_76, \843 );
and \U$792 ( \1626 , RI91439c8_60, \845 );
and \U$793 ( \1627 , RI9143248_44, \847 );
and \U$794 ( \1628 , RI90f39a0_28, \849 );
and \U$795 ( \1629 , RI912ea28_12, \851 );
or \U$796 ( \1630 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 );
_DC g698 ( \1631_nG698 , \1630 , \860 );
buf \U$797 ( \1632 , \1631_nG698 );
buf \U$798 ( \1633 , \1632 );
not \U$799 ( \1634 , \1633 );
and \U$800 ( \1635 , \912 , \1633 );
nor \U$801 ( \1636 , \1634 , \1635 );
and \U$802 ( \1637 , RI9149350_251, \821 );
and \U$803 ( \1638 , RI9148bd0_235, \823 );
and \U$804 ( \1639 , RI9148450_219, \825 );
and \U$805 ( \1640 , RI9147cd0_203, \827 );
and \U$806 ( \1641 , RI9147550_187, \829 );
and \U$807 ( \1642 , RI9146dd0_171, \831 );
and \U$808 ( \1643 , RI9146650_155, \833 );
and \U$809 ( \1644 , RI9145ed0_139, \835 );
and \U$810 ( \1645 , RI9145750_123, \837 );
and \U$811 ( \1646 , RI9144fd0_107, \839 );
and \U$812 ( \1647 , RI9144850_91, \841 );
and \U$813 ( \1648 , RI91440d0_75, \843 );
and \U$814 ( \1649 , RI9143950_59, \845 );
and \U$815 ( \1650 , RI90f3298_43, \847 );
and \U$816 ( \1651 , RI90f95f8_27, \849 );
and \U$817 ( \1652 , RI912eaa0_11, \851 );
or \U$818 ( \1653 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 );
_DC g6af ( \1654_nG6af , \1653 , \860 );
buf \U$819 ( \1655 , \1654_nG6af );
buf \U$820 ( \1656 , \1655 );
and \U$821 ( \1657 , \1656 , \954 );
and \U$822 ( \1658 , \1636 , \1657 );
and \U$823 ( \1659 , \1613 , \1658 );
xor \U$824 ( \1660 , \1559 , \1560 );
xor \U$825 ( \1661 , \1660 , \1562 );
and \U$826 ( \1662 , \1658 , \1661 );
and \U$827 ( \1663 , \1613 , \1661 );
or \U$828 ( \1664 , \1659 , \1662 , \1663 );
and \U$829 ( \1665 , \1165 , \1261 );
and \U$830 ( \1666 , \1061 , \1326 );
and \U$831 ( \1667 , \1665 , \1666 );
and \U$832 ( \1668 , \1084 , \1446 );
and \U$833 ( \1669 , \1666 , \1668 );
and \U$834 ( \1670 , \1665 , \1668 );
or \U$835 ( \1671 , \1667 , \1669 , \1670 );
xor \U$836 ( \1672 , \1521 , \1522 );
xor \U$837 ( \1673 , \1672 , \1524 );
and \U$838 ( \1674 , \1671 , \1673 );
and \U$839 ( \1675 , \1012 , \1446 );
and \U$840 ( \1676 , \863 , \1550 );
xor \U$841 ( \1677 , \1675 , \1676 );
and \U$842 ( \1678 , RI9150ad8_506, \869 );
and \U$843 ( \1679 , RI9150358_490, \871 );
and \U$844 ( \1680 , RI914fbd8_474, \873 );
and \U$845 ( \1681 , RI914f458_458, \875 );
and \U$846 ( \1682 , RI914ecd8_442, \877 );
and \U$847 ( \1683 , RI914e558_426, \879 );
and \U$848 ( \1684 , RI914ddd8_410, \881 );
and \U$849 ( \1685 , RI914d658_394, \883 );
and \U$850 ( \1686 , RI914ced8_378, \885 );
and \U$851 ( \1687 , RI914c758_362, \887 );
and \U$852 ( \1688 , RI914bfd8_346, \889 );
and \U$853 ( \1689 , RI914b858_330, \891 );
and \U$854 ( \1690 , RI914b0d8_314, \893 );
and \U$855 ( \1691 , RI914a958_298, \895 );
and \U$856 ( \1692 , RI914a1d8_282, \897 );
and \U$857 ( \1693 , RI9149a58_266, \899 );
or \U$858 ( \1694 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 );
_DC g6d8 ( \1695_nG6d8 , \1694 , \908 );
buf \U$859 ( \1696 , \1695_nG6d8 );
buf \U$860 ( \1697 , \1696 );
and \U$861 ( \1698 , \934 , \1697 );
xor \U$862 ( \1699 , \1677 , \1698 );
and \U$863 ( \1700 , \1673 , \1699 );
and \U$864 ( \1701 , \1671 , \1699 );
or \U$865 ( \1702 , \1674 , \1700 , \1701 );
and \U$866 ( \1703 , \1664 , \1702 );
xor \U$867 ( \1704 , \1527 , \1552 );
xor \U$868 ( \1705 , \1704 , \1555 );
and \U$869 ( \1706 , \1702 , \1705 );
and \U$870 ( \1707 , \1664 , \1705 );
or \U$871 ( \1708 , \1703 , \1706 , \1707 );
and \U$872 ( \1709 , \1606 , \1708 );
and \U$873 ( \1710 , \977 , \1550 );
not \U$874 ( \1711 , \1550 );
nor \U$875 ( \1712 , \1710 , \1711 );
and \U$876 ( \1713 , \1708 , \1712 );
and \U$877 ( \1714 , \1606 , \1712 );
or \U$878 ( \1715 , \1709 , \1713 , \1714 );
not \U$879 ( \1716 , \1656 );
and \U$880 ( \1717 , \912 , \1656 );
nor \U$881 ( \1718 , \1716 , \1717 );
xor \U$882 ( \1719 , \1613 , \1658 );
xor \U$883 ( \1720 , \1719 , \1661 );
and \U$884 ( \1721 , \1718 , \1720 );
xor \U$885 ( \1722 , \1664 , \1702 );
xor \U$886 ( \1723 , \1722 , \1705 );
and \U$887 ( \1724 , \1721 , \1723 );
xor \U$888 ( \1725 , \1565 , \1567 );
and \U$889 ( \1726 , \1723 , \1725 );
and \U$890 ( \1727 , \1721 , \1725 );
or \U$891 ( \1728 , \1724 , \1726 , \1727 );
xor \U$892 ( \1729 , \1606 , \1708 );
xor \U$893 ( \1730 , \1729 , \1712 );
and \U$894 ( \1731 , \1728 , \1730 );
xor \U$895 ( \1732 , \1583 , \1584 );
and \U$896 ( \1733 , \1730 , \1732 );
and \U$897 ( \1734 , \1728 , \1732 );
or \U$898 ( \1735 , \1731 , \1733 , \1734 );
and \U$899 ( \1736 , \1715 , \1735 );
xor \U$900 ( \1737 , \1585 , \1587 );
xor \U$901 ( \1738 , \1737 , \1589 );
and \U$902 ( \1739 , \1735 , \1738 );
and \U$903 ( \1740 , \1715 , \1738 );
or \U$904 ( \1741 , \1736 , \1739 , \1740 );
and \U$905 ( \1742 , \1602 , \1741 );
xor \U$906 ( \1743 , \1602 , \1741 );
xor \U$907 ( \1744 , \1715 , \1735 );
xor \U$908 ( \1745 , \1744 , \1738 );
and \U$909 ( \1746 , \1675 , \1676 );
and \U$910 ( \1747 , \1676 , \1698 );
and \U$911 ( \1748 , \1675 , \1698 );
or \U$912 ( \1749 , \1746 , \1747 , \1748 );
and \U$913 ( \1750 , RI9149440_253, \821 );
and \U$914 ( \1751 , RI9148cc0_237, \823 );
and \U$915 ( \1752 , RI9148540_221, \825 );
and \U$916 ( \1753 , RI9147dc0_205, \827 );
and \U$917 ( \1754 , RI9147640_189, \829 );
and \U$918 ( \1755 , RI9146ec0_173, \831 );
and \U$919 ( \1756 , RI9146740_157, \833 );
and \U$920 ( \1757 , RI9145fc0_141, \835 );
and \U$921 ( \1758 , RI9145840_125, \837 );
and \U$922 ( \1759 , RI91450c0_109, \839 );
and \U$923 ( \1760 , RI9144940_93, \841 );
and \U$924 ( \1761 , RI91441c0_77, \843 );
and \U$925 ( \1762 , RI9143a40_61, \845 );
and \U$926 ( \1763 , RI91432c0_45, \847 );
and \U$927 ( \1764 , RI90f3928_29, \849 );
and \U$928 ( \1765 , RI912e9b0_13, \851 );
or \U$929 ( \1766 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 , \1765 );
_DC g720 ( \1767_nG720 , \1766 , \860 );
buf \U$930 ( \1768 , \1767_nG720 );
buf \U$931 ( \1769 , \1768 );
not \U$932 ( \1770 , \1769 );
and \U$933 ( \1771 , \912 , \1769 );
nor \U$934 ( \1772 , \1770 , \1771 );
and \U$935 ( \1773 , \1633 , \954 );
and \U$936 ( \1774 , \1772 , \1773 );
and \U$937 ( \1775 , \1656 , \1037 );
and \U$938 ( \1776 , \1773 , \1775 );
and \U$939 ( \1777 , \1772 , \1775 );
or \U$940 ( \1778 , \1774 , \1776 , \1777 );
and \U$941 ( \1779 , \1471 , \1113 );
and \U$942 ( \1780 , \1354 , \1197 );
and \U$943 ( \1781 , \1779 , \1780 );
and \U$944 ( \1782 , \1377 , \1261 );
and \U$945 ( \1783 , \1780 , \1782 );
and \U$946 ( \1784 , \1779 , \1782 );
or \U$947 ( \1785 , \1781 , \1783 , \1784 );
and \U$948 ( \1786 , \1778 , \1785 );
xor \U$949 ( \1787 , \1607 , \1608 );
xor \U$950 ( \1788 , \1787 , \1610 );
and \U$951 ( \1789 , \1785 , \1788 );
and \U$952 ( \1790 , \1778 , \1788 );
or \U$953 ( \1791 , \1786 , \1789 , \1790 );
and \U$954 ( \1792 , \1165 , \1326 );
and \U$955 ( \1793 , \1061 , \1446 );
and \U$956 ( \1794 , \1792 , \1793 );
and \U$957 ( \1795 , \1084 , \1550 );
and \U$958 ( \1796 , \1793 , \1795 );
and \U$959 ( \1797 , \1792 , \1795 );
or \U$960 ( \1798 , \1794 , \1796 , \1797 );
xor \U$961 ( \1799 , \1665 , \1666 );
xor \U$962 ( \1800 , \1799 , \1668 );
and \U$963 ( \1801 , \1798 , \1800 );
and \U$964 ( \1802 , \1012 , \1550 );
and \U$965 ( \1803 , \863 , \1697 );
xor \U$966 ( \1804 , \1802 , \1803 );
and \U$967 ( \1805 , RI9150b50_507, \869 );
and \U$968 ( \1806 , RI91503d0_491, \871 );
and \U$969 ( \1807 , RI914fc50_475, \873 );
and \U$970 ( \1808 , RI914f4d0_459, \875 );
and \U$971 ( \1809 , RI914ed50_443, \877 );
and \U$972 ( \1810 , RI914e5d0_427, \879 );
and \U$973 ( \1811 , RI914de50_411, \881 );
and \U$974 ( \1812 , RI914d6d0_395, \883 );
and \U$975 ( \1813 , RI914cf50_379, \885 );
and \U$976 ( \1814 , RI914c7d0_363, \887 );
and \U$977 ( \1815 , RI914c050_347, \889 );
and \U$978 ( \1816 , RI914b8d0_331, \891 );
and \U$979 ( \1817 , RI914b150_315, \893 );
and \U$980 ( \1818 , RI914a9d0_299, \895 );
and \U$981 ( \1819 , RI914a250_283, \897 );
and \U$982 ( \1820 , RI9149ad0_267, \899 );
or \U$983 ( \1821 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 );
_DC g757 ( \1822_nG757 , \1821 , \908 );
buf \U$984 ( \1823 , \1822_nG757 );
buf \U$985 ( \1824 , \1823 );
and \U$986 ( \1825 , \934 , \1824 );
xor \U$987 ( \1826 , \1804 , \1825 );
and \U$988 ( \1827 , \1800 , \1826 );
and \U$989 ( \1828 , \1798 , \1826 );
or \U$990 ( \1829 , \1801 , \1827 , \1828 );
and \U$991 ( \1830 , \1791 , \1829 );
xor \U$992 ( \1831 , \1671 , \1673 );
xor \U$993 ( \1832 , \1831 , \1699 );
and \U$994 ( \1833 , \1829 , \1832 );
and \U$995 ( \1834 , \1791 , \1832 );
or \U$996 ( \1835 , \1830 , \1833 , \1834 );
and \U$997 ( \1836 , \1749 , \1835 );
and \U$998 ( \1837 , \977 , \1697 );
not \U$999 ( \1838 , \1697 );
nor \U$1000 ( \1839 , \1837 , \1838 );
and \U$1001 ( \1840 , \1835 , \1839 );
and \U$1002 ( \1841 , \1749 , \1839 );
or \U$1003 ( \1842 , \1836 , \1840 , \1841 );
xor \U$1004 ( \1843 , \1778 , \1785 );
xor \U$1005 ( \1844 , \1843 , \1788 );
xor \U$1006 ( \1845 , \1636 , \1657 );
and \U$1007 ( \1846 , \1844 , \1845 );
xor \U$1008 ( \1847 , \1791 , \1829 );
xor \U$1009 ( \1848 , \1847 , \1832 );
and \U$1010 ( \1849 , \1846 , \1848 );
xor \U$1011 ( \1850 , \1718 , \1720 );
and \U$1012 ( \1851 , \1848 , \1850 );
and \U$1013 ( \1852 , \1846 , \1850 );
or \U$1014 ( \1853 , \1849 , \1851 , \1852 );
xor \U$1015 ( \1854 , \1749 , \1835 );
xor \U$1016 ( \1855 , \1854 , \1839 );
and \U$1017 ( \1856 , \1853 , \1855 );
xor \U$1018 ( \1857 , \1721 , \1723 );
xor \U$1019 ( \1858 , \1857 , \1725 );
and \U$1020 ( \1859 , \1855 , \1858 );
and \U$1021 ( \1860 , \1853 , \1858 );
or \U$1022 ( \1861 , \1856 , \1859 , \1860 );
and \U$1023 ( \1862 , \1842 , \1861 );
xor \U$1024 ( \1863 , \1728 , \1730 );
xor \U$1025 ( \1864 , \1863 , \1732 );
and \U$1026 ( \1865 , \1861 , \1864 );
and \U$1027 ( \1866 , \1842 , \1864 );
or \U$1028 ( \1867 , \1862 , \1865 , \1866 );
and \U$1029 ( \1868 , \1745 , \1867 );
xor \U$1030 ( \1869 , \1745 , \1867 );
xor \U$1031 ( \1870 , \1842 , \1861 );
xor \U$1032 ( \1871 , \1870 , \1864 );
and \U$1033 ( \1872 , \1802 , \1803 );
and \U$1034 ( \1873 , \1803 , \1825 );
and \U$1035 ( \1874 , \1802 , \1825 );
or \U$1036 ( \1875 , \1872 , \1873 , \1874 );
and \U$1037 ( \1876 , \1165 , \1446 );
and \U$1038 ( \1877 , \1061 , \1550 );
and \U$1039 ( \1878 , \1876 , \1877 );
and \U$1040 ( \1879 , \1084 , \1697 );
and \U$1041 ( \1880 , \1877 , \1879 );
and \U$1042 ( \1881 , \1876 , \1879 );
or \U$1043 ( \1882 , \1878 , \1880 , \1881 );
xor \U$1044 ( \1883 , \1792 , \1793 );
xor \U$1045 ( \1884 , \1883 , \1795 );
and \U$1046 ( \1885 , \1882 , \1884 );
and \U$1047 ( \1886 , \1012 , \1697 );
and \U$1048 ( \1887 , \863 , \1824 );
xor \U$1049 ( \1888 , \1886 , \1887 );
and \U$1050 ( \1889 , RI9150bc8_508, \869 );
and \U$1051 ( \1890 , RI9150448_492, \871 );
and \U$1052 ( \1891 , RI914fcc8_476, \873 );
and \U$1053 ( \1892 , RI914f548_460, \875 );
and \U$1054 ( \1893 , RI914edc8_444, \877 );
and \U$1055 ( \1894 , RI914e648_428, \879 );
and \U$1056 ( \1895 , RI914dec8_412, \881 );
and \U$1057 ( \1896 , RI914d748_396, \883 );
and \U$1058 ( \1897 , RI914cfc8_380, \885 );
and \U$1059 ( \1898 , RI914c848_364, \887 );
and \U$1060 ( \1899 , RI914c0c8_348, \889 );
and \U$1061 ( \1900 , RI914b948_332, \891 );
and \U$1062 ( \1901 , RI914b1c8_316, \893 );
and \U$1063 ( \1902 , RI914aa48_300, \895 );
and \U$1064 ( \1903 , RI914a2c8_284, \897 );
and \U$1065 ( \1904 , RI9149b48_268, \899 );
or \U$1066 ( \1905 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 );
_DC g7ab ( \1906_nG7ab , \1905 , \908 );
buf \U$1067 ( \1907 , \1906_nG7ab );
buf \U$1068 ( \1908 , \1907 );
and \U$1069 ( \1909 , \934 , \1908 );
xor \U$1070 ( \1910 , \1888 , \1909 );
and \U$1071 ( \1911 , \1884 , \1910 );
and \U$1072 ( \1912 , \1882 , \1910 );
or \U$1073 ( \1913 , \1885 , \1911 , \1912 );
and \U$1074 ( \1914 , \1471 , \1197 );
and \U$1075 ( \1915 , \1354 , \1261 );
and \U$1076 ( \1916 , \1914 , \1915 );
and \U$1077 ( \1917 , \1377 , \1326 );
and \U$1078 ( \1918 , \1915 , \1917 );
and \U$1079 ( \1919 , \1914 , \1917 );
or \U$1080 ( \1920 , \1916 , \1918 , \1919 );
and \U$1081 ( \1921 , \1769 , \954 );
and \U$1082 ( \1922 , \1633 , \1037 );
and \U$1083 ( \1923 , \1921 , \1922 );
and \U$1084 ( \1924 , \1656 , \1113 );
and \U$1085 ( \1925 , \1922 , \1924 );
and \U$1086 ( \1926 , \1921 , \1924 );
or \U$1087 ( \1927 , \1923 , \1925 , \1926 );
and \U$1088 ( \1928 , \1920 , \1927 );
xor \U$1089 ( \1929 , \1779 , \1780 );
xor \U$1090 ( \1930 , \1929 , \1782 );
and \U$1091 ( \1931 , \1927 , \1930 );
and \U$1092 ( \1932 , \1920 , \1930 );
or \U$1093 ( \1933 , \1928 , \1931 , \1932 );
and \U$1094 ( \1934 , \1913 , \1933 );
xor \U$1095 ( \1935 , \1798 , \1800 );
xor \U$1096 ( \1936 , \1935 , \1826 );
and \U$1097 ( \1937 , \1933 , \1936 );
and \U$1098 ( \1938 , \1913 , \1936 );
or \U$1099 ( \1939 , \1934 , \1937 , \1938 );
and \U$1100 ( \1940 , \1875 , \1939 );
and \U$1101 ( \1941 , \977 , \1824 );
not \U$1102 ( \1942 , \1824 );
nor \U$1103 ( \1943 , \1941 , \1942 );
and \U$1104 ( \1944 , \1939 , \1943 );
and \U$1105 ( \1945 , \1875 , \1943 );
or \U$1106 ( \1946 , \1940 , \1944 , \1945 );
and \U$1107 ( \1947 , RI9149530_255, \821 );
and \U$1108 ( \1948 , RI9148db0_239, \823 );
and \U$1109 ( \1949 , RI9148630_223, \825 );
and \U$1110 ( \1950 , RI9147eb0_207, \827 );
and \U$1111 ( \1951 , RI9147730_191, \829 );
and \U$1112 ( \1952 , RI9146fb0_175, \831 );
and \U$1113 ( \1953 , RI9146830_159, \833 );
and \U$1114 ( \1954 , RI91460b0_143, \835 );
and \U$1115 ( \1955 , RI9145930_127, \837 );
and \U$1116 ( \1956 , RI91451b0_111, \839 );
and \U$1117 ( \1957 , RI9144a30_95, \841 );
and \U$1118 ( \1958 , RI91442b0_79, \843 );
and \U$1119 ( \1959 , RI9143b30_63, \845 );
and \U$1120 ( \1960 , RI91433b0_47, \847 );
and \U$1121 ( \1961 , RI90f3838_31, \849 );
and \U$1122 ( \1962 , RI912e8c0_15, \851 );
or \U$1123 ( \1963 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 );
_DC g7e5 ( \1964_nG7e5 , \1963 , \860 );
buf \U$1124 ( \1965 , \1964_nG7e5 );
buf \U$1125 ( \1966 , \1965 );
not \U$1126 ( \1967 , \1966 );
and \U$1127 ( \1968 , \912 , \1966 );
nor \U$1128 ( \1969 , \1967 , \1968 );
and \U$1129 ( \1970 , RI91494b8_254, \821 );
and \U$1130 ( \1971 , RI9148d38_238, \823 );
and \U$1131 ( \1972 , RI91485b8_222, \825 );
and \U$1132 ( \1973 , RI9147e38_206, \827 );
and \U$1133 ( \1974 , RI91476b8_190, \829 );
and \U$1134 ( \1975 , RI9146f38_174, \831 );
and \U$1135 ( \1976 , RI91467b8_158, \833 );
and \U$1136 ( \1977 , RI9146038_142, \835 );
and \U$1137 ( \1978 , RI91458b8_126, \837 );
and \U$1138 ( \1979 , RI9145138_110, \839 );
and \U$1139 ( \1980 , RI91449b8_94, \841 );
and \U$1140 ( \1981 , RI9144238_78, \843 );
and \U$1141 ( \1982 , RI9143ab8_62, \845 );
and \U$1142 ( \1983 , RI9143338_46, \847 );
and \U$1143 ( \1984 , RI90f38b0_30, \849 );
and \U$1144 ( \1985 , RI912e938_14, \851 );
or \U$1145 ( \1986 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 );
_DC g7fc ( \1987_nG7fc , \1986 , \860 );
buf \U$1146 ( \1988 , \1987_nG7fc );
buf \U$1147 ( \1989 , \1988 );
and \U$1148 ( \1990 , \1989 , \954 );
and \U$1149 ( \1991 , \1969 , \1990 );
not \U$1150 ( \1992 , \1989 );
and \U$1151 ( \1993 , \912 , \1989 );
nor \U$1152 ( \1994 , \1992 , \1993 );
and \U$1153 ( \1995 , \1991 , \1994 );
xor \U$1154 ( \1996 , \1921 , \1922 );
xor \U$1155 ( \1997 , \1996 , \1924 );
and \U$1156 ( \1998 , \1994 , \1997 );
and \U$1157 ( \1999 , \1991 , \1997 );
or \U$1158 ( \2000 , \1995 , \1998 , \1999 );
xor \U$1159 ( \2001 , \1772 , \1773 );
xor \U$1160 ( \2002 , \2001 , \1775 );
and \U$1161 ( \2003 , \2000 , \2002 );
xor \U$1162 ( \2004 , \1920 , \1927 );
xor \U$1163 ( \2005 , \2004 , \1930 );
and \U$1164 ( \2006 , \2002 , \2005 );
and \U$1165 ( \2007 , \2000 , \2005 );
or \U$1166 ( \2008 , \2003 , \2006 , \2007 );
xor \U$1167 ( \2009 , \1913 , \1933 );
xor \U$1168 ( \2010 , \2009 , \1936 );
and \U$1169 ( \2011 , \2008 , \2010 );
xor \U$1170 ( \2012 , \1844 , \1845 );
and \U$1171 ( \2013 , \2010 , \2012 );
and \U$1172 ( \2014 , \2008 , \2012 );
or \U$1173 ( \2015 , \2011 , \2013 , \2014 );
xor \U$1174 ( \2016 , \1875 , \1939 );
xor \U$1175 ( \2017 , \2016 , \1943 );
and \U$1176 ( \2018 , \2015 , \2017 );
xor \U$1177 ( \2019 , \1846 , \1848 );
xor \U$1178 ( \2020 , \2019 , \1850 );
and \U$1179 ( \2021 , \2017 , \2020 );
and \U$1180 ( \2022 , \2015 , \2020 );
or \U$1181 ( \2023 , \2018 , \2021 , \2022 );
and \U$1182 ( \2024 , \1946 , \2023 );
xor \U$1183 ( \2025 , \1853 , \1855 );
xor \U$1184 ( \2026 , \2025 , \1858 );
and \U$1185 ( \2027 , \2023 , \2026 );
and \U$1186 ( \2028 , \1946 , \2026 );
or \U$1187 ( \2029 , \2024 , \2027 , \2028 );
and \U$1188 ( \2030 , \1871 , \2029 );
xor \U$1189 ( \2031 , \1871 , \2029 );
xor \U$1190 ( \2032 , \1946 , \2023 );
xor \U$1191 ( \2033 , \2032 , \2026 );
and \U$1192 ( \2034 , \1886 , \1887 );
and \U$1193 ( \2035 , \1887 , \1909 );
and \U$1194 ( \2036 , \1886 , \1909 );
or \U$1195 ( \2037 , \2034 , \2035 , \2036 );
and \U$1196 ( \2038 , \1165 , \1550 );
and \U$1197 ( \2039 , \1061 , \1697 );
and \U$1198 ( \2040 , \2038 , \2039 );
and \U$1199 ( \2041 , \1084 , \1824 );
and \U$1200 ( \2042 , \2039 , \2041 );
and \U$1201 ( \2043 , \2038 , \2041 );
or \U$1202 ( \2044 , \2040 , \2042 , \2043 );
and \U$1203 ( \2045 , \1012 , \1824 );
and \U$1204 ( \2046 , \863 , \1908 );
xor \U$1205 ( \2047 , \2045 , \2046 );
and \U$1206 ( \2048 , RI9150c40_509, \869 );
and \U$1207 ( \2049 , RI91504c0_493, \871 );
and \U$1208 ( \2050 , RI914fd40_477, \873 );
and \U$1209 ( \2051 , RI914f5c0_461, \875 );
and \U$1210 ( \2052 , RI914ee40_445, \877 );
and \U$1211 ( \2053 , RI914e6c0_429, \879 );
and \U$1212 ( \2054 , RI914df40_413, \881 );
and \U$1213 ( \2055 , RI914d7c0_397, \883 );
and \U$1214 ( \2056 , RI914d040_381, \885 );
and \U$1215 ( \2057 , RI914c8c0_365, \887 );
and \U$1216 ( \2058 , RI914c140_349, \889 );
and \U$1217 ( \2059 , RI914b9c0_333, \891 );
and \U$1218 ( \2060 , RI914b240_317, \893 );
and \U$1219 ( \2061 , RI914aac0_301, \895 );
and \U$1220 ( \2062 , RI914a340_285, \897 );
and \U$1221 ( \2063 , RI9149bc0_269, \899 );
or \U$1222 ( \2064 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 );
_DC g84a ( \2065_nG84a , \2064 , \908 );
buf \U$1223 ( \2066 , \2065_nG84a );
buf \U$1224 ( \2067 , \2066 );
and \U$1225 ( \2068 , \934 , \2067 );
xor \U$1226 ( \2069 , \2047 , \2068 );
and \U$1227 ( \2070 , \2044 , \2069 );
xor \U$1228 ( \2071 , \1876 , \1877 );
xor \U$1229 ( \2072 , \2071 , \1879 );
and \U$1230 ( \2073 , \2069 , \2072 );
and \U$1231 ( \2074 , \2044 , \2072 );
or \U$1232 ( \2075 , \2070 , \2073 , \2074 );
and \U$1233 ( \2076 , \1471 , \1261 );
and \U$1234 ( \2077 , \1354 , \1326 );
and \U$1235 ( \2078 , \2076 , \2077 );
and \U$1236 ( \2079 , \1377 , \1446 );
and \U$1237 ( \2080 , \2077 , \2079 );
and \U$1238 ( \2081 , \2076 , \2079 );
or \U$1239 ( \2082 , \2078 , \2080 , \2081 );
and \U$1240 ( \2083 , \1769 , \1037 );
and \U$1241 ( \2084 , \1633 , \1113 );
and \U$1242 ( \2085 , \2083 , \2084 );
and \U$1243 ( \2086 , \1656 , \1197 );
and \U$1244 ( \2087 , \2084 , \2086 );
and \U$1245 ( \2088 , \2083 , \2086 );
or \U$1246 ( \2089 , \2085 , \2087 , \2088 );
and \U$1247 ( \2090 , \2082 , \2089 );
xor \U$1248 ( \2091 , \1914 , \1915 );
xor \U$1249 ( \2092 , \2091 , \1917 );
and \U$1250 ( \2093 , \2089 , \2092 );
and \U$1251 ( \2094 , \2082 , \2092 );
or \U$1252 ( \2095 , \2090 , \2093 , \2094 );
and \U$1253 ( \2096 , \2075 , \2095 );
xor \U$1254 ( \2097 , \1882 , \1884 );
xor \U$1255 ( \2098 , \2097 , \1910 );
and \U$1256 ( \2099 , \2095 , \2098 );
and \U$1257 ( \2100 , \2075 , \2098 );
or \U$1258 ( \2101 , \2096 , \2099 , \2100 );
and \U$1259 ( \2102 , \2037 , \2101 );
and \U$1260 ( \2103 , \977 , \1908 );
not \U$1261 ( \2104 , \1908 );
nor \U$1262 ( \2105 , \2103 , \2104 );
and \U$1263 ( \2106 , \2101 , \2105 );
and \U$1264 ( \2107 , \2037 , \2105 );
or \U$1265 ( \2108 , \2102 , \2106 , \2107 );
and \U$1266 ( \2109 , RI91495a8_256, \821 );
and \U$1267 ( \2110 , RI9148e28_240, \823 );
and \U$1268 ( \2111 , RI91486a8_224, \825 );
and \U$1269 ( \2112 , RI9147f28_208, \827 );
and \U$1270 ( \2113 , RI91477a8_192, \829 );
and \U$1271 ( \2114 , RI9147028_176, \831 );
and \U$1272 ( \2115 , RI91468a8_160, \833 );
and \U$1273 ( \2116 , RI9146128_144, \835 );
and \U$1274 ( \2117 , RI91459a8_128, \837 );
and \U$1275 ( \2118 , RI9145228_112, \839 );
and \U$1276 ( \2119 , RI9144aa8_96, \841 );
and \U$1277 ( \2120 , RI9144328_80, \843 );
and \U$1278 ( \2121 , RI9143ba8_64, \845 );
and \U$1279 ( \2122 , RI9143428_48, \847 );
and \U$1280 ( \2123 , RI90f37c0_32, \849 );
and \U$1281 ( \2124 , RI912e848_16, \851 );
or \U$1282 ( \2125 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 );
_DC g887 ( \2126_nG887 , \2125 , \860 );
buf \U$1283 ( \2127 , \2126_nG887 );
buf \U$1284 ( \2128 , \2127 );
not \U$1285 ( \2129 , \2128 );
and \U$1286 ( \2130 , \912 , \2128 );
nor \U$1287 ( \2131 , \2129 , \2130 );
and \U$1288 ( \2132 , \1966 , \954 );
and \U$1289 ( \2133 , \2131 , \2132 );
and \U$1290 ( \2134 , \1989 , \1037 );
and \U$1291 ( \2135 , \2132 , \2134 );
and \U$1292 ( \2136 , \2131 , \2134 );
or \U$1293 ( \2137 , \2133 , \2135 , \2136 );
xor \U$1294 ( \2138 , \2083 , \2084 );
xor \U$1295 ( \2139 , \2138 , \2086 );
and \U$1296 ( \2140 , \2137 , \2139 );
xor \U$1297 ( \2141 , \1969 , \1990 );
and \U$1298 ( \2142 , \2139 , \2141 );
and \U$1299 ( \2143 , \2137 , \2141 );
or \U$1300 ( \2144 , \2140 , \2142 , \2143 );
xor \U$1301 ( \2145 , \2082 , \2089 );
xor \U$1302 ( \2146 , \2145 , \2092 );
and \U$1303 ( \2147 , \2144 , \2146 );
xor \U$1304 ( \2148 , \1991 , \1994 );
xor \U$1305 ( \2149 , \2148 , \1997 );
and \U$1306 ( \2150 , \2146 , \2149 );
and \U$1307 ( \2151 , \2144 , \2149 );
or \U$1308 ( \2152 , \2147 , \2150 , \2151 );
xor \U$1309 ( \2153 , \2075 , \2095 );
xor \U$1310 ( \2154 , \2153 , \2098 );
and \U$1311 ( \2155 , \2152 , \2154 );
xor \U$1312 ( \2156 , \2000 , \2002 );
xor \U$1313 ( \2157 , \2156 , \2005 );
and \U$1314 ( \2158 , \2154 , \2157 );
and \U$1315 ( \2159 , \2152 , \2157 );
or \U$1316 ( \2160 , \2155 , \2158 , \2159 );
xor \U$1317 ( \2161 , \2037 , \2101 );
xor \U$1318 ( \2162 , \2161 , \2105 );
and \U$1319 ( \2163 , \2160 , \2162 );
xor \U$1320 ( \2164 , \2008 , \2010 );
xor \U$1321 ( \2165 , \2164 , \2012 );
and \U$1322 ( \2166 , \2162 , \2165 );
and \U$1323 ( \2167 , \2160 , \2165 );
or \U$1324 ( \2168 , \2163 , \2166 , \2167 );
and \U$1325 ( \2169 , \2108 , \2168 );
xor \U$1326 ( \2170 , \2015 , \2017 );
xor \U$1327 ( \2171 , \2170 , \2020 );
and \U$1328 ( \2172 , \2168 , \2171 );
and \U$1329 ( \2173 , \2108 , \2171 );
or \U$1330 ( \2174 , \2169 , \2172 , \2173 );
and \U$1331 ( \2175 , \2033 , \2174 );
xor \U$1332 ( \2176 , \2033 , \2174 );
xor \U$1333 ( \2177 , \2108 , \2168 );
xor \U$1334 ( \2178 , \2177 , \2171 );
and \U$1335 ( \2179 , \2045 , \2046 );
and \U$1336 ( \2180 , \2046 , \2068 );
and \U$1337 ( \2181 , \2045 , \2068 );
or \U$1338 ( \2182 , \2179 , \2180 , \2181 );
and \U$1339 ( \2183 , \1165 , \1697 );
and \U$1340 ( \2184 , \1061 , \1824 );
and \U$1341 ( \2185 , \2183 , \2184 );
and \U$1342 ( \2186 , \1084 , \1908 );
and \U$1343 ( \2187 , \2184 , \2186 );
and \U$1344 ( \2188 , \2183 , \2186 );
or \U$1345 ( \2189 , \2185 , \2187 , \2188 );
and \U$1346 ( \2190 , \1012 , \1908 );
and \U$1347 ( \2191 , \863 , \2067 );
xor \U$1348 ( \2192 , \2190 , \2191 );
and \U$1349 ( \2193 , RI9150cb8_510, \869 );
and \U$1350 ( \2194 , RI9150538_494, \871 );
and \U$1351 ( \2195 , RI914fdb8_478, \873 );
and \U$1352 ( \2196 , RI914f638_462, \875 );
and \U$1353 ( \2197 , RI914eeb8_446, \877 );
and \U$1354 ( \2198 , RI914e738_430, \879 );
and \U$1355 ( \2199 , RI914dfb8_414, \881 );
and \U$1356 ( \2200 , RI914d838_398, \883 );
and \U$1357 ( \2201 , RI914d0b8_382, \885 );
and \U$1358 ( \2202 , RI914c938_366, \887 );
and \U$1359 ( \2203 , RI914c1b8_350, \889 );
and \U$1360 ( \2204 , RI914ba38_334, \891 );
and \U$1361 ( \2205 , RI914b2b8_318, \893 );
and \U$1362 ( \2206 , RI914ab38_302, \895 );
and \U$1363 ( \2207 , RI914a3b8_286, \897 );
and \U$1364 ( \2208 , RI9149c38_270, \899 );
or \U$1365 ( \2209 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 );
_DC g8db ( \2210_nG8db , \2209 , \908 );
buf \U$1366 ( \2211 , \2210_nG8db );
buf \U$1367 ( \2212 , \2211 );
and \U$1368 ( \2213 , \934 , \2212 );
xor \U$1369 ( \2214 , \2192 , \2213 );
and \U$1370 ( \2215 , \2189 , \2214 );
xor \U$1371 ( \2216 , \2038 , \2039 );
xor \U$1372 ( \2217 , \2216 , \2041 );
and \U$1373 ( \2218 , \2214 , \2217 );
and \U$1374 ( \2219 , \2189 , \2217 );
or \U$1375 ( \2220 , \2215 , \2218 , \2219 );
and \U$1376 ( \2221 , \1471 , \1326 );
and \U$1377 ( \2222 , \1354 , \1446 );
and \U$1378 ( \2223 , \2221 , \2222 );
and \U$1379 ( \2224 , \1377 , \1550 );
and \U$1380 ( \2225 , \2222 , \2224 );
and \U$1381 ( \2226 , \2221 , \2224 );
or \U$1382 ( \2227 , \2223 , \2225 , \2226 );
and \U$1383 ( \2228 , \1769 , \1113 );
and \U$1384 ( \2229 , \1633 , \1197 );
and \U$1385 ( \2230 , \2228 , \2229 );
and \U$1386 ( \2231 , \1656 , \1261 );
and \U$1387 ( \2232 , \2229 , \2231 );
and \U$1388 ( \2233 , \2228 , \2231 );
or \U$1389 ( \2234 , \2230 , \2232 , \2233 );
and \U$1390 ( \2235 , \2227 , \2234 );
xor \U$1391 ( \2236 , \2076 , \2077 );
xor \U$1392 ( \2237 , \2236 , \2079 );
and \U$1393 ( \2238 , \2234 , \2237 );
and \U$1394 ( \2239 , \2227 , \2237 );
or \U$1395 ( \2240 , \2235 , \2238 , \2239 );
and \U$1396 ( \2241 , \2220 , \2240 );
xor \U$1397 ( \2242 , \2044 , \2069 );
xor \U$1398 ( \2243 , \2242 , \2072 );
and \U$1399 ( \2244 , \2240 , \2243 );
and \U$1400 ( \2245 , \2220 , \2243 );
or \U$1401 ( \2246 , \2241 , \2244 , \2245 );
and \U$1402 ( \2247 , \2182 , \2246 );
and \U$1403 ( \2248 , \977 , \2067 );
not \U$1404 ( \2249 , \2067 );
nor \U$1405 ( \2250 , \2248 , \2249 );
and \U$1406 ( \2251 , \2246 , \2250 );
and \U$1407 ( \2252 , \2182 , \2250 );
or \U$1408 ( \2253 , \2247 , \2251 , \2252 );
and \U$1409 ( \2254 , \2128 , \954 );
and \U$1410 ( \2255 , \1966 , \1037 );
and \U$1411 ( \2256 , \2254 , \2255 );
and \U$1412 ( \2257 , \1989 , \1113 );
and \U$1413 ( \2258 , \2255 , \2257 );
and \U$1414 ( \2259 , \2254 , \2257 );
or \U$1415 ( \2260 , \2256 , \2258 , \2259 );
xor \U$1416 ( \2261 , \2228 , \2229 );
xor \U$1417 ( \2262 , \2261 , \2231 );
and \U$1418 ( \2263 , \2260 , \2262 );
xor \U$1419 ( \2264 , \2131 , \2132 );
xor \U$1420 ( \2265 , \2264 , \2134 );
and \U$1421 ( \2266 , \2262 , \2265 );
and \U$1422 ( \2267 , \2260 , \2265 );
or \U$1423 ( \2268 , \2263 , \2266 , \2267 );
xor \U$1424 ( \2269 , \2227 , \2234 );
xor \U$1425 ( \2270 , \2269 , \2237 );
and \U$1426 ( \2271 , \2268 , \2270 );
xor \U$1427 ( \2272 , \2137 , \2139 );
xor \U$1428 ( \2273 , \2272 , \2141 );
and \U$1429 ( \2274 , \2270 , \2273 );
and \U$1430 ( \2275 , \2268 , \2273 );
or \U$1431 ( \2276 , \2271 , \2274 , \2275 );
xor \U$1432 ( \2277 , \2220 , \2240 );
xor \U$1433 ( \2278 , \2277 , \2243 );
and \U$1434 ( \2279 , \2276 , \2278 );
xor \U$1435 ( \2280 , \2144 , \2146 );
xor \U$1436 ( \2281 , \2280 , \2149 );
and \U$1437 ( \2282 , \2278 , \2281 );
and \U$1438 ( \2283 , \2276 , \2281 );
or \U$1439 ( \2284 , \2279 , \2282 , \2283 );
xor \U$1440 ( \2285 , \2182 , \2246 );
xor \U$1441 ( \2286 , \2285 , \2250 );
and \U$1442 ( \2287 , \2284 , \2286 );
xor \U$1443 ( \2288 , \2152 , \2154 );
xor \U$1444 ( \2289 , \2288 , \2157 );
and \U$1445 ( \2290 , \2286 , \2289 );
and \U$1446 ( \2291 , \2284 , \2289 );
or \U$1447 ( \2292 , \2287 , \2290 , \2291 );
and \U$1448 ( \2293 , \2253 , \2292 );
xor \U$1449 ( \2294 , \2160 , \2162 );
xor \U$1450 ( \2295 , \2294 , \2165 );
and \U$1451 ( \2296 , \2292 , \2295 );
and \U$1452 ( \2297 , \2253 , \2295 );
or \U$1453 ( \2298 , \2293 , \2296 , \2297 );
and \U$1454 ( \2299 , \2178 , \2298 );
xor \U$1455 ( \2300 , \2178 , \2298 );
xor \U$1456 ( \2301 , \2253 , \2292 );
xor \U$1457 ( \2302 , \2301 , \2295 );
and \U$1458 ( \2303 , \2190 , \2191 );
and \U$1459 ( \2304 , \2191 , \2213 );
and \U$1460 ( \2305 , \2190 , \2213 );
or \U$1461 ( \2306 , \2303 , \2304 , \2305 );
and \U$1462 ( \2307 , \1165 , \1824 );
and \U$1463 ( \2308 , \1061 , \1908 );
and \U$1464 ( \2309 , \2307 , \2308 );
and \U$1465 ( \2310 , \1084 , \2067 );
and \U$1466 ( \2311 , \2308 , \2310 );
and \U$1467 ( \2312 , \2307 , \2310 );
or \U$1468 ( \2313 , \2309 , \2311 , \2312 );
and \U$1469 ( \2314 , \1012 , \2067 );
and \U$1470 ( \2315 , \863 , \2212 );
xor \U$1471 ( \2316 , \2314 , \2315 );
and \U$1472 ( \2317 , RI9150d30_511, \869 );
and \U$1473 ( \2318 , RI91505b0_495, \871 );
and \U$1474 ( \2319 , RI914fe30_479, \873 );
and \U$1475 ( \2320 , RI914f6b0_463, \875 );
and \U$1476 ( \2321 , RI914ef30_447, \877 );
and \U$1477 ( \2322 , RI914e7b0_431, \879 );
and \U$1478 ( \2323 , RI914e030_415, \881 );
and \U$1479 ( \2324 , RI914d8b0_399, \883 );
and \U$1480 ( \2325 , RI914d130_383, \885 );
and \U$1481 ( \2326 , RI914c9b0_367, \887 );
and \U$1482 ( \2327 , RI914c230_351, \889 );
and \U$1483 ( \2328 , RI914bab0_335, \891 );
and \U$1484 ( \2329 , RI914b330_319, \893 );
and \U$1485 ( \2330 , RI914abb0_303, \895 );
and \U$1486 ( \2331 , RI914a430_287, \897 );
and \U$1487 ( \2332 , RI9149cb0_271, \899 );
or \U$1488 ( \2333 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 );
_DC g957 ( \2334_nG957 , \2333 , \908 );
buf \U$1489 ( \2335 , \2334_nG957 );
buf \U$1490 ( \2336 , \2335 );
and \U$1491 ( \2337 , \934 , \2336 );
xor \U$1492 ( \2338 , \2316 , \2337 );
and \U$1493 ( \2339 , \2313 , \2338 );
xor \U$1494 ( \2340 , \2183 , \2184 );
xor \U$1495 ( \2341 , \2340 , \2186 );
and \U$1496 ( \2342 , \2338 , \2341 );
and \U$1497 ( \2343 , \2313 , \2341 );
or \U$1498 ( \2344 , \2339 , \2342 , \2343 );
and \U$1499 ( \2345 , \1471 , \1446 );
and \U$1500 ( \2346 , \1354 , \1550 );
and \U$1501 ( \2347 , \2345 , \2346 );
and \U$1502 ( \2348 , \1377 , \1697 );
and \U$1503 ( \2349 , \2346 , \2348 );
and \U$1504 ( \2350 , \2345 , \2348 );
or \U$1505 ( \2351 , \2347 , \2349 , \2350 );
and \U$1506 ( \2352 , \1769 , \1197 );
and \U$1507 ( \2353 , \1633 , \1261 );
and \U$1508 ( \2354 , \2352 , \2353 );
and \U$1509 ( \2355 , \1656 , \1326 );
and \U$1510 ( \2356 , \2353 , \2355 );
and \U$1511 ( \2357 , \2352 , \2355 );
or \U$1512 ( \2358 , \2354 , \2356 , \2357 );
and \U$1513 ( \2359 , \2351 , \2358 );
xor \U$1514 ( \2360 , \2221 , \2222 );
xor \U$1515 ( \2361 , \2360 , \2224 );
and \U$1516 ( \2362 , \2358 , \2361 );
and \U$1517 ( \2363 , \2351 , \2361 );
or \U$1518 ( \2364 , \2359 , \2362 , \2363 );
and \U$1519 ( \2365 , \2344 , \2364 );
xor \U$1520 ( \2366 , \2189 , \2214 );
xor \U$1521 ( \2367 , \2366 , \2217 );
and \U$1522 ( \2368 , \2364 , \2367 );
and \U$1523 ( \2369 , \2344 , \2367 );
or \U$1524 ( \2370 , \2365 , \2368 , \2369 );
and \U$1525 ( \2371 , \2306 , \2370 );
and \U$1526 ( \2372 , \977 , \2212 );
not \U$1527 ( \2373 , \2212 );
nor \U$1528 ( \2374 , \2372 , \2373 );
and \U$1529 ( \2375 , \2370 , \2374 );
and \U$1530 ( \2376 , \2306 , \2374 );
or \U$1531 ( \2377 , \2371 , \2375 , \2376 );
and \U$1532 ( \2378 , \2128 , \1037 );
and \U$1533 ( \2379 , \1966 , \1113 );
and \U$1534 ( \2380 , \2378 , \2379 );
and \U$1535 ( \2381 , \1989 , \1197 );
and \U$1536 ( \2382 , \2379 , \2381 );
and \U$1537 ( \2383 , \2378 , \2381 );
or \U$1538 ( \2384 , \2380 , \2382 , \2383 );
xor \U$1539 ( \2385 , \2352 , \2353 );
xor \U$1540 ( \2386 , \2385 , \2355 );
and \U$1541 ( \2387 , \2384 , \2386 );
xor \U$1542 ( \2388 , \2254 , \2255 );
xor \U$1543 ( \2389 , \2388 , \2257 );
and \U$1544 ( \2390 , \2386 , \2389 );
and \U$1545 ( \2391 , \2384 , \2389 );
or \U$1546 ( \2392 , \2387 , \2390 , \2391 );
xor \U$1547 ( \2393 , \2351 , \2358 );
xor \U$1548 ( \2394 , \2393 , \2361 );
and \U$1549 ( \2395 , \2392 , \2394 );
xor \U$1550 ( \2396 , \2260 , \2262 );
xor \U$1551 ( \2397 , \2396 , \2265 );
and \U$1552 ( \2398 , \2394 , \2397 );
and \U$1553 ( \2399 , \2392 , \2397 );
or \U$1554 ( \2400 , \2395 , \2398 , \2399 );
xor \U$1555 ( \2401 , \2344 , \2364 );
xor \U$1556 ( \2402 , \2401 , \2367 );
and \U$1557 ( \2403 , \2400 , \2402 );
xor \U$1558 ( \2404 , \2268 , \2270 );
xor \U$1559 ( \2405 , \2404 , \2273 );
and \U$1560 ( \2406 , \2402 , \2405 );
and \U$1561 ( \2407 , \2400 , \2405 );
or \U$1562 ( \2408 , \2403 , \2406 , \2407 );
xor \U$1563 ( \2409 , \2306 , \2370 );
xor \U$1564 ( \2410 , \2409 , \2374 );
and \U$1565 ( \2411 , \2408 , \2410 );
xor \U$1566 ( \2412 , \2276 , \2278 );
xor \U$1567 ( \2413 , \2412 , \2281 );
and \U$1568 ( \2414 , \2410 , \2413 );
and \U$1569 ( \2415 , \2408 , \2413 );
or \U$1570 ( \2416 , \2411 , \2414 , \2415 );
and \U$1571 ( \2417 , \2377 , \2416 );
xor \U$1572 ( \2418 , \2284 , \2286 );
xor \U$1573 ( \2419 , \2418 , \2289 );
and \U$1574 ( \2420 , \2416 , \2419 );
and \U$1575 ( \2421 , \2377 , \2419 );
or \U$1576 ( \2422 , \2417 , \2420 , \2421 );
and \U$1577 ( \2423 , \2302 , \2422 );
xor \U$1578 ( \2424 , \2302 , \2422 );
xor \U$1579 ( \2425 , \2377 , \2416 );
xor \U$1580 ( \2426 , \2425 , \2419 );
and \U$1581 ( \2427 , \2314 , \2315 );
and \U$1582 ( \2428 , \2315 , \2337 );
and \U$1583 ( \2429 , \2314 , \2337 );
or \U$1584 ( \2430 , \2427 , \2428 , \2429 );
and \U$1585 ( \2431 , \1165 , \1908 );
and \U$1586 ( \2432 , \1061 , \2067 );
and \U$1587 ( \2433 , \2431 , \2432 );
and \U$1588 ( \2434 , \1084 , \2212 );
and \U$1589 ( \2435 , \2432 , \2434 );
and \U$1590 ( \2436 , \2431 , \2434 );
or \U$1591 ( \2437 , \2433 , \2435 , \2436 );
and \U$1592 ( \2438 , \1012 , \2212 );
and \U$1593 ( \2439 , \863 , \2336 );
xor \U$1594 ( \2440 , \2438 , \2439 );
and \U$1595 ( \2441 , RI9150da8_512, \869 );
and \U$1596 ( \2442 , RI9150628_496, \871 );
and \U$1597 ( \2443 , RI914fea8_480, \873 );
and \U$1598 ( \2444 , RI914f728_464, \875 );
and \U$1599 ( \2445 , RI914efa8_448, \877 );
and \U$1600 ( \2446 , RI914e828_432, \879 );
and \U$1601 ( \2447 , RI914e0a8_416, \881 );
and \U$1602 ( \2448 , RI914d928_400, \883 );
and \U$1603 ( \2449 , RI914d1a8_384, \885 );
and \U$1604 ( \2450 , RI914ca28_368, \887 );
and \U$1605 ( \2451 , RI914c2a8_352, \889 );
and \U$1606 ( \2452 , RI914bb28_336, \891 );
and \U$1607 ( \2453 , RI914b3a8_320, \893 );
and \U$1608 ( \2454 , RI914ac28_304, \895 );
and \U$1609 ( \2455 , RI914a4a8_288, \897 );
and \U$1610 ( \2456 , RI9149d28_272, \899 );
or \U$1611 ( \2457 , \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 );
_DC g9d3 ( \2458_nG9d3 , \2457 , \908 );
buf \U$1612 ( \2459 , \2458_nG9d3 );
buf \U$1613 ( \2460 , \2459 );
and \U$1614 ( \2461 , \934 , \2460 );
xor \U$1615 ( \2462 , \2440 , \2461 );
and \U$1616 ( \2463 , \2437 , \2462 );
xor \U$1617 ( \2464 , \2307 , \2308 );
xor \U$1618 ( \2465 , \2464 , \2310 );
and \U$1619 ( \2466 , \2462 , \2465 );
and \U$1620 ( \2467 , \2437 , \2465 );
or \U$1621 ( \2468 , \2463 , \2466 , \2467 );
and \U$1622 ( \2469 , \1471 , \1550 );
and \U$1623 ( \2470 , \1354 , \1697 );
and \U$1624 ( \2471 , \2469 , \2470 );
and \U$1625 ( \2472 , \1377 , \1824 );
and \U$1626 ( \2473 , \2470 , \2472 );
and \U$1627 ( \2474 , \2469 , \2472 );
or \U$1628 ( \2475 , \2471 , \2473 , \2474 );
and \U$1629 ( \2476 , \1769 , \1261 );
and \U$1630 ( \2477 , \1633 , \1326 );
and \U$1631 ( \2478 , \2476 , \2477 );
and \U$1632 ( \2479 , \1656 , \1446 );
and \U$1633 ( \2480 , \2477 , \2479 );
and \U$1634 ( \2481 , \2476 , \2479 );
or \U$1635 ( \2482 , \2478 , \2480 , \2481 );
and \U$1636 ( \2483 , \2475 , \2482 );
xor \U$1637 ( \2484 , \2345 , \2346 );
xor \U$1638 ( \2485 , \2484 , \2348 );
and \U$1639 ( \2486 , \2482 , \2485 );
and \U$1640 ( \2487 , \2475 , \2485 );
or \U$1641 ( \2488 , \2483 , \2486 , \2487 );
and \U$1642 ( \2489 , \2468 , \2488 );
xor \U$1643 ( \2490 , \2313 , \2338 );
xor \U$1644 ( \2491 , \2490 , \2341 );
and \U$1645 ( \2492 , \2488 , \2491 );
and \U$1646 ( \2493 , \2468 , \2491 );
or \U$1647 ( \2494 , \2489 , \2492 , \2493 );
and \U$1648 ( \2495 , \2430 , \2494 );
and \U$1649 ( \2496 , \977 , \2336 );
not \U$1650 ( \2497 , \2336 );
nor \U$1651 ( \2498 , \2496 , \2497 );
and \U$1652 ( \2499 , \2494 , \2498 );
and \U$1653 ( \2500 , \2430 , \2498 );
or \U$1654 ( \2501 , \2495 , \2499 , \2500 );
and \U$1655 ( \2502 , \2128 , \1113 );
and \U$1656 ( \2503 , \1966 , \1197 );
and \U$1657 ( \2504 , \2502 , \2503 );
and \U$1658 ( \2505 , \1989 , \1261 );
and \U$1659 ( \2506 , \2503 , \2505 );
and \U$1660 ( \2507 , \2502 , \2505 );
or \U$1661 ( \2508 , \2504 , \2506 , \2507 );
xor \U$1662 ( \2509 , \2476 , \2477 );
xor \U$1663 ( \2510 , \2509 , \2479 );
and \U$1664 ( \2511 , \2508 , \2510 );
xor \U$1665 ( \2512 , \2378 , \2379 );
xor \U$1666 ( \2513 , \2512 , \2381 );
and \U$1667 ( \2514 , \2510 , \2513 );
and \U$1668 ( \2515 , \2508 , \2513 );
or \U$1669 ( \2516 , \2511 , \2514 , \2515 );
xor \U$1670 ( \2517 , \2475 , \2482 );
xor \U$1671 ( \2518 , \2517 , \2485 );
and \U$1672 ( \2519 , \2516 , \2518 );
xor \U$1673 ( \2520 , \2384 , \2386 );
xor \U$1674 ( \2521 , \2520 , \2389 );
and \U$1675 ( \2522 , \2518 , \2521 );
and \U$1676 ( \2523 , \2516 , \2521 );
or \U$1677 ( \2524 , \2519 , \2522 , \2523 );
xor \U$1678 ( \2525 , \2468 , \2488 );
xor \U$1679 ( \2526 , \2525 , \2491 );
and \U$1680 ( \2527 , \2524 , \2526 );
xor \U$1681 ( \2528 , \2392 , \2394 );
xor \U$1682 ( \2529 , \2528 , \2397 );
and \U$1683 ( \2530 , \2526 , \2529 );
and \U$1684 ( \2531 , \2524 , \2529 );
or \U$1685 ( \2532 , \2527 , \2530 , \2531 );
xor \U$1686 ( \2533 , \2430 , \2494 );
xor \U$1687 ( \2534 , \2533 , \2498 );
and \U$1688 ( \2535 , \2532 , \2534 );
xor \U$1689 ( \2536 , \2400 , \2402 );
xor \U$1690 ( \2537 , \2536 , \2405 );
and \U$1691 ( \2538 , \2534 , \2537 );
and \U$1692 ( \2539 , \2532 , \2537 );
or \U$1693 ( \2540 , \2535 , \2538 , \2539 );
and \U$1694 ( \2541 , \2501 , \2540 );
xor \U$1695 ( \2542 , \2408 , \2410 );
xor \U$1696 ( \2543 , \2542 , \2413 );
and \U$1697 ( \2544 , \2540 , \2543 );
and \U$1698 ( \2545 , \2501 , \2543 );
or \U$1699 ( \2546 , \2541 , \2544 , \2545 );
and \U$1700 ( \2547 , \2426 , \2546 );
xor \U$1701 ( \2548 , \2426 , \2546 );
xor \U$1702 ( \2549 , \2501 , \2540 );
xor \U$1703 ( \2550 , \2549 , \2543 );
and \U$1704 ( \2551 , \2438 , \2439 );
and \U$1705 ( \2552 , \2439 , \2461 );
and \U$1706 ( \2553 , \2438 , \2461 );
or \U$1707 ( \2554 , \2551 , \2552 , \2553 );
and \U$1708 ( \2555 , \1471 , \1697 );
and \U$1709 ( \2556 , \1354 , \1824 );
and \U$1710 ( \2557 , \2555 , \2556 );
and \U$1711 ( \2558 , \1377 , \1908 );
and \U$1712 ( \2559 , \2556 , \2558 );
and \U$1713 ( \2560 , \2555 , \2558 );
or \U$1714 ( \2561 , \2557 , \2559 , \2560 );
and \U$1715 ( \2562 , \1769 , \1326 );
and \U$1716 ( \2563 , \1633 , \1446 );
and \U$1717 ( \2564 , \2562 , \2563 );
and \U$1718 ( \2565 , \1656 , \1550 );
and \U$1719 ( \2566 , \2563 , \2565 );
and \U$1720 ( \2567 , \2562 , \2565 );
or \U$1721 ( \2568 , \2564 , \2566 , \2567 );
and \U$1722 ( \2569 , \2561 , \2568 );
xor \U$1723 ( \2570 , \2469 , \2470 );
xor \U$1724 ( \2571 , \2570 , \2472 );
and \U$1725 ( \2572 , \2568 , \2571 );
and \U$1726 ( \2573 , \2561 , \2571 );
or \U$1727 ( \2574 , \2569 , \2572 , \2573 );
and \U$1728 ( \2575 , \1165 , \2067 );
and \U$1729 ( \2576 , \1061 , \2212 );
and \U$1730 ( \2577 , \2575 , \2576 );
and \U$1731 ( \2578 , \1084 , \2336 );
and \U$1732 ( \2579 , \2576 , \2578 );
and \U$1733 ( \2580 , \2575 , \2578 );
or \U$1734 ( \2581 , \2577 , \2579 , \2580 );
xor \U$1735 ( \2582 , \2431 , \2432 );
xor \U$1736 ( \2583 , \2582 , \2434 );
and \U$1737 ( \2584 , \2581 , \2583 );
and \U$1738 ( \2585 , \1012 , \2336 );
and \U$1739 ( \2586 , \863 , \2460 );
xor \U$1740 ( \2587 , \2585 , \2586 );
and \U$1741 ( \2588 , \2583 , \2587 );
and \U$1742 ( \2589 , \2581 , \2587 );
or \U$1743 ( \2590 , \2584 , \2588 , \2589 );
and \U$1744 ( \2591 , \2574 , \2590 );
xor \U$1745 ( \2592 , \2437 , \2462 );
xor \U$1746 ( \2593 , \2592 , \2465 );
and \U$1747 ( \2594 , \2590 , \2593 );
and \U$1748 ( \2595 , \2574 , \2593 );
or \U$1749 ( \2596 , \2591 , \2594 , \2595 );
and \U$1750 ( \2597 , \2554 , \2596 );
and \U$1751 ( \2598 , \977 , \2460 );
not \U$1752 ( \2599 , \2460 );
nor \U$1753 ( \2600 , \2598 , \2599 );
and \U$1754 ( \2601 , \2596 , \2600 );
and \U$1755 ( \2602 , \2554 , \2600 );
or \U$1756 ( \2603 , \2597 , \2601 , \2602 );
and \U$1757 ( \2604 , \2128 , \1197 );
and \U$1758 ( \2605 , \1966 , \1261 );
and \U$1759 ( \2606 , \2604 , \2605 );
and \U$1760 ( \2607 , \1989 , \1326 );
and \U$1761 ( \2608 , \2605 , \2607 );
and \U$1762 ( \2609 , \2604 , \2607 );
or \U$1763 ( \2610 , \2606 , \2608 , \2609 );
xor \U$1764 ( \2611 , \2562 , \2563 );
xor \U$1765 ( \2612 , \2611 , \2565 );
and \U$1766 ( \2613 , \2610 , \2612 );
xor \U$1767 ( \2614 , \2502 , \2503 );
xor \U$1768 ( \2615 , \2614 , \2505 );
and \U$1769 ( \2616 , \2612 , \2615 );
and \U$1770 ( \2617 , \2610 , \2615 );
or \U$1771 ( \2618 , \2613 , \2616 , \2617 );
xor \U$1772 ( \2619 , \2561 , \2568 );
xor \U$1773 ( \2620 , \2619 , \2571 );
and \U$1774 ( \2621 , \2618 , \2620 );
xor \U$1775 ( \2622 , \2508 , \2510 );
xor \U$1776 ( \2623 , \2622 , \2513 );
and \U$1777 ( \2624 , \2620 , \2623 );
and \U$1778 ( \2625 , \2618 , \2623 );
or \U$1779 ( \2626 , \2621 , \2624 , \2625 );
xor \U$1780 ( \2627 , \2574 , \2590 );
xor \U$1781 ( \2628 , \2627 , \2593 );
and \U$1782 ( \2629 , \2626 , \2628 );
xor \U$1783 ( \2630 , \2516 , \2518 );
xor \U$1784 ( \2631 , \2630 , \2521 );
and \U$1785 ( \2632 , \2628 , \2631 );
and \U$1786 ( \2633 , \2626 , \2631 );
or \U$1787 ( \2634 , \2629 , \2632 , \2633 );
xor \U$1788 ( \2635 , \2554 , \2596 );
xor \U$1789 ( \2636 , \2635 , \2600 );
and \U$1790 ( \2637 , \2634 , \2636 );
xor \U$1791 ( \2638 , \2524 , \2526 );
xor \U$1792 ( \2639 , \2638 , \2529 );
and \U$1793 ( \2640 , \2636 , \2639 );
and \U$1794 ( \2641 , \2634 , \2639 );
or \U$1795 ( \2642 , \2637 , \2640 , \2641 );
and \U$1796 ( \2643 , \2603 , \2642 );
xor \U$1797 ( \2644 , \2532 , \2534 );
xor \U$1798 ( \2645 , \2644 , \2537 );
and \U$1799 ( \2646 , \2642 , \2645 );
and \U$1800 ( \2647 , \2603 , \2645 );
or \U$1801 ( \2648 , \2643 , \2646 , \2647 );
and \U$1802 ( \2649 , \2550 , \2648 );
xor \U$1803 ( \2650 , \2550 , \2648 );
xor \U$1804 ( \2651 , \2603 , \2642 );
xor \U$1805 ( \2652 , \2651 , \2645 );
and \U$1806 ( \2653 , \2585 , \2586 );
and \U$1807 ( \2654 , \1165 , \2212 );
and \U$1808 ( \2655 , \1061 , \2336 );
and \U$1809 ( \2656 , \2654 , \2655 );
and \U$1810 ( \2657 , \1084 , \2460 );
and \U$1811 ( \2658 , \2655 , \2657 );
and \U$1812 ( \2659 , \2654 , \2657 );
or \U$1813 ( \2660 , \2656 , \2658 , \2659 );
and \U$1814 ( \2661 , \1012 , \2460 );
and \U$1815 ( \2662 , \2660 , \2661 );
xor \U$1816 ( \2663 , \2575 , \2576 );
xor \U$1817 ( \2664 , \2663 , \2578 );
and \U$1818 ( \2665 , \2661 , \2664 );
and \U$1819 ( \2666 , \2660 , \2664 );
or \U$1820 ( \2667 , \2662 , \2665 , \2666 );
and \U$1821 ( \2668 , \1471 , \1824 );
and \U$1822 ( \2669 , \1354 , \1908 );
and \U$1823 ( \2670 , \2668 , \2669 );
and \U$1824 ( \2671 , \1377 , \2067 );
and \U$1825 ( \2672 , \2669 , \2671 );
and \U$1826 ( \2673 , \2668 , \2671 );
or \U$1827 ( \2674 , \2670 , \2672 , \2673 );
and \U$1828 ( \2675 , \1769 , \1446 );
and \U$1829 ( \2676 , \1633 , \1550 );
and \U$1830 ( \2677 , \2675 , \2676 );
and \U$1831 ( \2678 , \1656 , \1697 );
and \U$1832 ( \2679 , \2676 , \2678 );
and \U$1833 ( \2680 , \2675 , \2678 );
or \U$1834 ( \2681 , \2677 , \2679 , \2680 );
and \U$1835 ( \2682 , \2674 , \2681 );
xor \U$1836 ( \2683 , \2555 , \2556 );
xor \U$1837 ( \2684 , \2683 , \2558 );
and \U$1838 ( \2685 , \2681 , \2684 );
and \U$1839 ( \2686 , \2674 , \2684 );
or \U$1840 ( \2687 , \2682 , \2685 , \2686 );
and \U$1841 ( \2688 , \2667 , \2687 );
xor \U$1842 ( \2689 , \2581 , \2583 );
xor \U$1843 ( \2690 , \2689 , \2587 );
and \U$1844 ( \2691 , \2687 , \2690 );
and \U$1845 ( \2692 , \2667 , \2690 );
or \U$1846 ( \2693 , \2688 , \2691 , \2692 );
and \U$1847 ( \2694 , \2653 , \2693 );
and \U$1848 ( \2695 , \2128 , \1261 );
and \U$1849 ( \2696 , \1966 , \1326 );
and \U$1850 ( \2697 , \2695 , \2696 );
and \U$1851 ( \2698 , \1989 , \1446 );
and \U$1852 ( \2699 , \2696 , \2698 );
and \U$1853 ( \2700 , \2695 , \2698 );
or \U$1854 ( \2701 , \2697 , \2699 , \2700 );
xor \U$1855 ( \2702 , \2675 , \2676 );
xor \U$1856 ( \2703 , \2702 , \2678 );
and \U$1857 ( \2704 , \2701 , \2703 );
xor \U$1858 ( \2705 , \2604 , \2605 );
xor \U$1859 ( \2706 , \2705 , \2607 );
and \U$1860 ( \2707 , \2703 , \2706 );
and \U$1861 ( \2708 , \2701 , \2706 );
or \U$1862 ( \2709 , \2704 , \2707 , \2708 );
xor \U$1863 ( \2710 , \2674 , \2681 );
xor \U$1864 ( \2711 , \2710 , \2684 );
and \U$1865 ( \2712 , \2709 , \2711 );
xor \U$1866 ( \2713 , \2610 , \2612 );
xor \U$1867 ( \2714 , \2713 , \2615 );
and \U$1868 ( \2715 , \2711 , \2714 );
and \U$1869 ( \2716 , \2709 , \2714 );
or \U$1870 ( \2717 , \2712 , \2715 , \2716 );
xor \U$1871 ( \2718 , \2618 , \2620 );
xor \U$1872 ( \2719 , \2718 , \2623 );
and \U$1873 ( \2720 , \2717 , \2719 );
xor \U$1874 ( \2721 , \2667 , \2687 );
xor \U$1875 ( \2722 , \2721 , \2690 );
and \U$1876 ( \2723 , \2719 , \2722 );
and \U$1877 ( \2724 , \2717 , \2722 );
or \U$1878 ( \2725 , \2720 , \2723 , \2724 );
xor \U$1879 ( \2726 , \2626 , \2628 );
xor \U$1880 ( \2727 , \2726 , \2631 );
and \U$1881 ( \2728 , \2725 , \2727 );
xor \U$1882 ( \2729 , \2653 , \2693 );
and \U$1883 ( \2730 , \2727 , \2729 );
and \U$1884 ( \2731 , \2725 , \2729 );
or \U$1885 ( \2732 , \2728 , \2730 , \2731 );
and \U$1886 ( \2733 , \2694 , \2732 );
xor \U$1887 ( \2734 , \2634 , \2636 );
xor \U$1888 ( \2735 , \2734 , \2639 );
and \U$1889 ( \2736 , \2732 , \2735 );
and \U$1890 ( \2737 , \2694 , \2735 );
or \U$1891 ( \2738 , \2733 , \2736 , \2737 );
and \U$1892 ( \2739 , \2652 , \2738 );
xor \U$1893 ( \2740 , \2652 , \2738 );
xor \U$1894 ( \2741 , \2694 , \2732 );
xor \U$1895 ( \2742 , \2741 , \2735 );
xor \U$1896 ( \2743 , \2725 , \2727 );
xor \U$1897 ( \2744 , \2743 , \2729 );
and \U$1898 ( \2745 , \1769 , \1550 );
and \U$1899 ( \2746 , \1633 , \1697 );
and \U$1900 ( \2747 , \2745 , \2746 );
and \U$1901 ( \2748 , \1656 , \1824 );
and \U$1902 ( \2749 , \2746 , \2748 );
and \U$1903 ( \2750 , \2745 , \2748 );
or \U$1904 ( \2751 , \2747 , \2749 , \2750 );
and \U$1905 ( \2752 , \1471 , \1908 );
and \U$1906 ( \2753 , \1354 , \2067 );
and \U$1907 ( \2754 , \2752 , \2753 );
and \U$1908 ( \2755 , \1377 , \2212 );
and \U$1909 ( \2756 , \2753 , \2755 );
and \U$1910 ( \2757 , \2752 , \2755 );
or \U$1911 ( \2758 , \2754 , \2756 , \2757 );
and \U$1912 ( \2759 , \2751 , \2758 );
xor \U$1913 ( \2760 , \2668 , \2669 );
xor \U$1914 ( \2761 , \2760 , \2671 );
and \U$1915 ( \2762 , \2758 , \2761 );
and \U$1916 ( \2763 , \2751 , \2761 );
or \U$1917 ( \2764 , \2759 , \2762 , \2763 );
and \U$1918 ( \2765 , \1165 , \2336 );
and \U$1919 ( \2766 , \1061 , \2460 );
and \U$1920 ( \2767 , \2765 , \2766 );
xor \U$1921 ( \2768 , \2654 , \2655 );
xor \U$1922 ( \2769 , \2768 , \2657 );
and \U$1923 ( \2770 , \2767 , \2769 );
and \U$1924 ( \2771 , \2764 , \2770 );
xor \U$1925 ( \2772 , \2660 , \2661 );
xor \U$1926 ( \2773 , \2772 , \2664 );
and \U$1927 ( \2774 , \2770 , \2773 );
and \U$1928 ( \2775 , \2764 , \2773 );
or \U$1929 ( \2776 , \2771 , \2774 , \2775 );
and \U$1930 ( \2777 , \2128 , \1326 );
and \U$1931 ( \2778 , \1966 , \1446 );
and \U$1932 ( \2779 , \2777 , \2778 );
and \U$1933 ( \2780 , \1989 , \1550 );
and \U$1934 ( \2781 , \2778 , \2780 );
and \U$1935 ( \2782 , \2777 , \2780 );
or \U$1936 ( \2783 , \2779 , \2781 , \2782 );
xor \U$1937 ( \2784 , \2745 , \2746 );
xor \U$1938 ( \2785 , \2784 , \2748 );
and \U$1939 ( \2786 , \2783 , \2785 );
xor \U$1940 ( \2787 , \2695 , \2696 );
xor \U$1941 ( \2788 , \2787 , \2698 );
and \U$1942 ( \2789 , \2785 , \2788 );
and \U$1943 ( \2790 , \2783 , \2788 );
or \U$1944 ( \2791 , \2786 , \2789 , \2790 );
xor \U$1945 ( \2792 , \2751 , \2758 );
xor \U$1946 ( \2793 , \2792 , \2761 );
and \U$1947 ( \2794 , \2791 , \2793 );
xor \U$1948 ( \2795 , \2701 , \2703 );
xor \U$1949 ( \2796 , \2795 , \2706 );
and \U$1950 ( \2797 , \2793 , \2796 );
and \U$1951 ( \2798 , \2791 , \2796 );
or \U$1952 ( \2799 , \2794 , \2797 , \2798 );
xor \U$1953 ( \2800 , \2764 , \2770 );
xor \U$1954 ( \2801 , \2800 , \2773 );
and \U$1955 ( \2802 , \2799 , \2801 );
xor \U$1956 ( \2803 , \2709 , \2711 );
xor \U$1957 ( \2804 , \2803 , \2714 );
and \U$1958 ( \2805 , \2801 , \2804 );
and \U$1959 ( \2806 , \2799 , \2804 );
or \U$1960 ( \2807 , \2802 , \2805 , \2806 );
and \U$1961 ( \2808 , \2776 , \2807 );
xor \U$1962 ( \2809 , \2717 , \2719 );
xor \U$1963 ( \2810 , \2809 , \2722 );
and \U$1964 ( \2811 , \2807 , \2810 );
and \U$1965 ( \2812 , \2776 , \2810 );
or \U$1966 ( \2813 , \2808 , \2811 , \2812 );
and \U$1967 ( \2814 , \2744 , \2813 );
xor \U$1968 ( \2815 , \2744 , \2813 );
xor \U$1969 ( \2816 , \2776 , \2807 );
xor \U$1970 ( \2817 , \2816 , \2810 );
and \U$1971 ( \2818 , \1471 , \2067 );
and \U$1972 ( \2819 , \1354 , \2212 );
and \U$1973 ( \2820 , \2818 , \2819 );
and \U$1974 ( \2821 , \1377 , \2336 );
and \U$1975 ( \2822 , \2819 , \2821 );
and \U$1976 ( \2823 , \2818 , \2821 );
or \U$1977 ( \2824 , \2820 , \2822 , \2823 );
and \U$1978 ( \2825 , \1769 , \1697 );
and \U$1979 ( \2826 , \1633 , \1824 );
and \U$1980 ( \2827 , \2825 , \2826 );
and \U$1981 ( \2828 , \1656 , \1908 );
and \U$1982 ( \2829 , \2826 , \2828 );
and \U$1983 ( \2830 , \2825 , \2828 );
or \U$1984 ( \2831 , \2827 , \2829 , \2830 );
and \U$1985 ( \2832 , \2824 , \2831 );
xor \U$1986 ( \2833 , \2752 , \2753 );
xor \U$1987 ( \2834 , \2833 , \2755 );
and \U$1988 ( \2835 , \2831 , \2834 );
and \U$1989 ( \2836 , \2824 , \2834 );
or \U$1990 ( \2837 , \2832 , \2835 , \2836 );
xor \U$1991 ( \2838 , \2767 , \2769 );
and \U$1992 ( \2839 , \2837 , \2838 );
and \U$1993 ( \2840 , \2128 , \1446 );
and \U$1994 ( \2841 , \1966 , \1550 );
and \U$1995 ( \2842 , \2840 , \2841 );
and \U$1996 ( \2843 , \1989 , \1697 );
and \U$1997 ( \2844 , \2841 , \2843 );
and \U$1998 ( \2845 , \2840 , \2843 );
or \U$1999 ( \2846 , \2842 , \2844 , \2845 );
xor \U$2000 ( \2847 , \2825 , \2826 );
xor \U$2001 ( \2848 , \2847 , \2828 );
and \U$2002 ( \2849 , \2846 , \2848 );
xor \U$2003 ( \2850 , \2777 , \2778 );
xor \U$2004 ( \2851 , \2850 , \2780 );
and \U$2005 ( \2852 , \2848 , \2851 );
and \U$2006 ( \2853 , \2846 , \2851 );
or \U$2007 ( \2854 , \2849 , \2852 , \2853 );
xor \U$2008 ( \2855 , \2783 , \2785 );
xor \U$2009 ( \2856 , \2855 , \2788 );
and \U$2010 ( \2857 , \2854 , \2856 );
xor \U$2011 ( \2858 , \2824 , \2831 );
xor \U$2012 ( \2859 , \2858 , \2834 );
and \U$2013 ( \2860 , \2856 , \2859 );
and \U$2014 ( \2861 , \2854 , \2859 );
or \U$2015 ( \2862 , \2857 , \2860 , \2861 );
xor \U$2016 ( \2863 , \2791 , \2793 );
xor \U$2017 ( \2864 , \2863 , \2796 );
and \U$2018 ( \2865 , \2862 , \2864 );
xor \U$2019 ( \2866 , \2837 , \2838 );
and \U$2020 ( \2867 , \2864 , \2866 );
and \U$2021 ( \2868 , \2862 , \2866 );
or \U$2022 ( \2869 , \2865 , \2867 , \2868 );
and \U$2023 ( \2870 , \2839 , \2869 );
xor \U$2024 ( \2871 , \2799 , \2801 );
xor \U$2025 ( \2872 , \2871 , \2804 );
and \U$2026 ( \2873 , \2869 , \2872 );
and \U$2027 ( \2874 , \2839 , \2872 );
or \U$2028 ( \2875 , \2870 , \2873 , \2874 );
and \U$2029 ( \2876 , \2817 , \2875 );
xor \U$2030 ( \2877 , \2817 , \2875 );
xor \U$2031 ( \2878 , \2839 , \2869 );
xor \U$2032 ( \2879 , \2878 , \2872 );
and \U$2033 ( \2880 , \1471 , \2212 );
and \U$2034 ( \2881 , \1354 , \2336 );
and \U$2035 ( \2882 , \2880 , \2881 );
and \U$2036 ( \2883 , \1377 , \2460 );
and \U$2037 ( \2884 , \2881 , \2883 );
and \U$2038 ( \2885 , \2880 , \2883 );
or \U$2039 ( \2886 , \2882 , \2884 , \2885 );
and \U$2040 ( \2887 , \1769 , \1824 );
and \U$2041 ( \2888 , \1633 , \1908 );
and \U$2042 ( \2889 , \2887 , \2888 );
and \U$2043 ( \2890 , \1656 , \2067 );
and \U$2044 ( \2891 , \2888 , \2890 );
and \U$2045 ( \2892 , \2887 , \2890 );
or \U$2046 ( \2893 , \2889 , \2891 , \2892 );
and \U$2047 ( \2894 , \2886 , \2893 );
xor \U$2048 ( \2895 , \2818 , \2819 );
xor \U$2049 ( \2896 , \2895 , \2821 );
and \U$2050 ( \2897 , \2893 , \2896 );
and \U$2051 ( \2898 , \2886 , \2896 );
or \U$2052 ( \2899 , \2894 , \2897 , \2898 );
xor \U$2053 ( \2900 , \2765 , \2766 );
and \U$2054 ( \2901 , \2899 , \2900 );
and \U$2055 ( \2902 , \2128 , \1550 );
and \U$2056 ( \2903 , \1966 , \1697 );
and \U$2057 ( \2904 , \2902 , \2903 );
and \U$2058 ( \2905 , \1989 , \1824 );
and \U$2059 ( \2906 , \2903 , \2905 );
and \U$2060 ( \2907 , \2902 , \2905 );
or \U$2061 ( \2908 , \2904 , \2906 , \2907 );
xor \U$2062 ( \2909 , \2887 , \2888 );
xor \U$2063 ( \2910 , \2909 , \2890 );
and \U$2064 ( \2911 , \2908 , \2910 );
xor \U$2065 ( \2912 , \2840 , \2841 );
xor \U$2066 ( \2913 , \2912 , \2843 );
and \U$2067 ( \2914 , \2910 , \2913 );
and \U$2068 ( \2915 , \2908 , \2913 );
or \U$2069 ( \2916 , \2911 , \2914 , \2915 );
xor \U$2070 ( \2917 , \2886 , \2893 );
xor \U$2071 ( \2918 , \2917 , \2896 );
and \U$2072 ( \2919 , \2916 , \2918 );
xor \U$2073 ( \2920 , \2846 , \2848 );
xor \U$2074 ( \2921 , \2920 , \2851 );
and \U$2075 ( \2922 , \2918 , \2921 );
and \U$2076 ( \2923 , \2916 , \2921 );
or \U$2077 ( \2924 , \2919 , \2922 , \2923 );
xor \U$2078 ( \2925 , \2854 , \2856 );
xor \U$2079 ( \2926 , \2925 , \2859 );
and \U$2080 ( \2927 , \2924 , \2926 );
xor \U$2081 ( \2928 , \2899 , \2900 );
and \U$2082 ( \2929 , \2926 , \2928 );
and \U$2083 ( \2930 , \2924 , \2928 );
or \U$2084 ( \2931 , \2927 , \2929 , \2930 );
and \U$2085 ( \2932 , \2901 , \2931 );
xor \U$2086 ( \2933 , \2862 , \2864 );
xor \U$2087 ( \2934 , \2933 , \2866 );
and \U$2088 ( \2935 , \2931 , \2934 );
and \U$2089 ( \2936 , \2901 , \2934 );
or \U$2090 ( \2937 , \2932 , \2935 , \2936 );
and \U$2091 ( \2938 , \2879 , \2937 );
xor \U$2092 ( \2939 , \2879 , \2937 );
xor \U$2093 ( \2940 , \2901 , \2931 );
xor \U$2094 ( \2941 , \2940 , \2934 );
and \U$2095 ( \2942 , \1769 , \1908 );
and \U$2096 ( \2943 , \1633 , \2067 );
and \U$2097 ( \2944 , \2942 , \2943 );
and \U$2098 ( \2945 , \1656 , \2212 );
and \U$2099 ( \2946 , \2943 , \2945 );
and \U$2100 ( \2947 , \2942 , \2945 );
or \U$2101 ( \2948 , \2944 , \2946 , \2947 );
and \U$2102 ( \2949 , \1471 , \2336 );
and \U$2103 ( \2950 , \1354 , \2460 );
and \U$2104 ( \2951 , \2949 , \2950 );
and \U$2105 ( \2952 , \2948 , \2951 );
xor \U$2106 ( \2953 , \2880 , \2881 );
xor \U$2107 ( \2954 , \2953 , \2883 );
and \U$2108 ( \2955 , \2951 , \2954 );
and \U$2109 ( \2956 , \2948 , \2954 );
or \U$2110 ( \2957 , \2952 , \2955 , \2956 );
and \U$2111 ( \2958 , \1165 , \2460 );
and \U$2112 ( \2959 , \2957 , \2958 );
and \U$2113 ( \2960 , \2128 , \1697 );
and \U$2114 ( \2961 , \1966 , \1824 );
and \U$2115 ( \2962 , \2960 , \2961 );
and \U$2116 ( \2963 , \1989 , \1908 );
and \U$2117 ( \2964 , \2961 , \2963 );
and \U$2118 ( \2965 , \2960 , \2963 );
or \U$2119 ( \2966 , \2962 , \2964 , \2965 );
xor \U$2120 ( \2967 , \2902 , \2903 );
xor \U$2121 ( \2968 , \2967 , \2905 );
and \U$2122 ( \2969 , \2966 , \2968 );
xor \U$2123 ( \2970 , \2942 , \2943 );
xor \U$2124 ( \2971 , \2970 , \2945 );
and \U$2125 ( \2972 , \2968 , \2971 );
and \U$2126 ( \2973 , \2966 , \2971 );
or \U$2127 ( \2974 , \2969 , \2972 , \2973 );
xor \U$2128 ( \2975 , \2948 , \2951 );
xor \U$2129 ( \2976 , \2975 , \2954 );
and \U$2130 ( \2977 , \2974 , \2976 );
xor \U$2131 ( \2978 , \2908 , \2910 );
xor \U$2132 ( \2979 , \2978 , \2913 );
and \U$2133 ( \2980 , \2976 , \2979 );
and \U$2134 ( \2981 , \2974 , \2979 );
or \U$2135 ( \2982 , \2977 , \2980 , \2981 );
xor \U$2136 ( \2983 , \2916 , \2918 );
xor \U$2137 ( \2984 , \2983 , \2921 );
and \U$2138 ( \2985 , \2982 , \2984 );
xor \U$2139 ( \2986 , \2957 , \2958 );
and \U$2140 ( \2987 , \2984 , \2986 );
and \U$2141 ( \2988 , \2982 , \2986 );
or \U$2142 ( \2989 , \2985 , \2987 , \2988 );
and \U$2143 ( \2990 , \2959 , \2989 );
xor \U$2144 ( \2991 , \2924 , \2926 );
xor \U$2145 ( \2992 , \2991 , \2928 );
and \U$2146 ( \2993 , \2989 , \2992 );
and \U$2147 ( \2994 , \2959 , \2992 );
or \U$2148 ( \2995 , \2990 , \2993 , \2994 );
and \U$2149 ( \2996 , \2941 , \2995 );
xor \U$2150 ( \2997 , \2941 , \2995 );
xor \U$2151 ( \2998 , \2959 , \2989 );
xor \U$2152 ( \2999 , \2998 , \2992 );
xor \U$2153 ( \3000 , \2982 , \2984 );
xor \U$2154 ( \3001 , \3000 , \2986 );
and \U$2155 ( \3002 , \1769 , \2067 );
and \U$2156 ( \3003 , \1633 , \2212 );
and \U$2157 ( \3004 , \3002 , \3003 );
and \U$2158 ( \3005 , \1656 , \2336 );
and \U$2159 ( \3006 , \3003 , \3005 );
and \U$2160 ( \3007 , \3002 , \3005 );
or \U$2161 ( \3008 , \3004 , \3006 , \3007 );
xor \U$2162 ( \3009 , \2949 , \2950 );
and \U$2163 ( \3010 , \3008 , \3009 );
and \U$2164 ( \3011 , \2128 , \1824 );
and \U$2165 ( \3012 , \1966 , \1908 );
and \U$2166 ( \3013 , \3011 , \3012 );
and \U$2167 ( \3014 , \1989 , \2067 );
and \U$2168 ( \3015 , \3012 , \3014 );
and \U$2169 ( \3016 , \3011 , \3014 );
or \U$2170 ( \3017 , \3013 , \3015 , \3016 );
xor \U$2171 ( \3018 , \3002 , \3003 );
xor \U$2172 ( \3019 , \3018 , \3005 );
and \U$2173 ( \3020 , \3017 , \3019 );
xor \U$2174 ( \3021 , \2960 , \2961 );
xor \U$2175 ( \3022 , \3021 , \2963 );
and \U$2176 ( \3023 , \3019 , \3022 );
and \U$2177 ( \3024 , \3017 , \3022 );
or \U$2178 ( \3025 , \3020 , \3023 , \3024 );
xor \U$2179 ( \3026 , \2966 , \2968 );
xor \U$2180 ( \3027 , \3026 , \2971 );
and \U$2181 ( \3028 , \3025 , \3027 );
xor \U$2182 ( \3029 , \3008 , \3009 );
and \U$2183 ( \3030 , \3027 , \3029 );
and \U$2184 ( \3031 , \3025 , \3029 );
or \U$2185 ( \3032 , \3028 , \3030 , \3031 );
and \U$2186 ( \3033 , \3010 , \3032 );
xor \U$2187 ( \3034 , \2974 , \2976 );
xor \U$2188 ( \3035 , \3034 , \2979 );
and \U$2189 ( \3036 , \3032 , \3035 );
and \U$2190 ( \3037 , \3010 , \3035 );
or \U$2191 ( \3038 , \3033 , \3036 , \3037 );
and \U$2192 ( \3039 , \3001 , \3038 );
xor \U$2193 ( \3040 , \3001 , \3038 );
xor \U$2194 ( \3041 , \3010 , \3032 );
xor \U$2195 ( \3042 , \3041 , \3035 );
and \U$2196 ( \3043 , \1769 , \2212 );
and \U$2197 ( \3044 , \1633 , \2336 );
and \U$2198 ( \3045 , \3043 , \3044 );
and \U$2199 ( \3046 , \1656 , \2460 );
and \U$2200 ( \3047 , \3044 , \3046 );
and \U$2201 ( \3048 , \3043 , \3046 );
or \U$2202 ( \3049 , \3045 , \3047 , \3048 );
and \U$2203 ( \3050 , \1471 , \2460 );
and \U$2204 ( \3051 , \3049 , \3050 );
and \U$2205 ( \3052 , \2128 , \1908 );
and \U$2206 ( \3053 , \1966 , \2067 );
and \U$2207 ( \3054 , \3052 , \3053 );
and \U$2208 ( \3055 , \1989 , \2212 );
and \U$2209 ( \3056 , \3053 , \3055 );
and \U$2210 ( \3057 , \3052 , \3055 );
or \U$2211 ( \3058 , \3054 , \3056 , \3057 );
xor \U$2212 ( \3059 , \3043 , \3044 );
xor \U$2213 ( \3060 , \3059 , \3046 );
and \U$2214 ( \3061 , \3058 , \3060 );
xor \U$2215 ( \3062 , \3011 , \3012 );
xor \U$2216 ( \3063 , \3062 , \3014 );
and \U$2217 ( \3064 , \3060 , \3063 );
and \U$2218 ( \3065 , \3058 , \3063 );
or \U$2219 ( \3066 , \3061 , \3064 , \3065 );
xor \U$2220 ( \3067 , \3017 , \3019 );
xor \U$2221 ( \3068 , \3067 , \3022 );
and \U$2222 ( \3069 , \3066 , \3068 );
xor \U$2223 ( \3070 , \3049 , \3050 );
and \U$2224 ( \3071 , \3068 , \3070 );
and \U$2225 ( \3072 , \3066 , \3070 );
or \U$2226 ( \3073 , \3069 , \3071 , \3072 );
and \U$2227 ( \3074 , \3051 , \3073 );
xor \U$2228 ( \3075 , \3025 , \3027 );
xor \U$2229 ( \3076 , \3075 , \3029 );
and \U$2230 ( \3077 , \3073 , \3076 );
and \U$2231 ( \3078 , \3051 , \3076 );
or \U$2232 ( \3079 , \3074 , \3077 , \3078 );
and \U$2233 ( \3080 , \3042 , \3079 );
xor \U$2234 ( \3081 , \3042 , \3079 );
xor \U$2235 ( \3082 , \3051 , \3073 );
xor \U$2236 ( \3083 , \3082 , \3076 );
xor \U$2237 ( \3084 , \3066 , \3068 );
xor \U$2238 ( \3085 , \3084 , \3070 );
and \U$2239 ( \3086 , \1769 , \2336 );
and \U$2240 ( \3087 , \1633 , \2460 );
and \U$2241 ( \3088 , \3086 , \3087 );
and \U$2242 ( \3089 , \2128 , \2067 );
and \U$2243 ( \3090 , \1966 , \2212 );
and \U$2244 ( \3091 , \3089 , \3090 );
and \U$2245 ( \3092 , \1989 , \2336 );
and \U$2246 ( \3093 , \3090 , \3092 );
and \U$2247 ( \3094 , \3089 , \3092 );
or \U$2248 ( \3095 , \3091 , \3093 , \3094 );
xor \U$2249 ( \3096 , \3052 , \3053 );
xor \U$2250 ( \3097 , \3096 , \3055 );
and \U$2251 ( \3098 , \3095 , \3097 );
xor \U$2252 ( \3099 , \3086 , \3087 );
and \U$2253 ( \3100 , \3097 , \3099 );
and \U$2254 ( \3101 , \3095 , \3099 );
or \U$2255 ( \3102 , \3098 , \3100 , \3101 );
and \U$2256 ( \3103 , \3088 , \3102 );
xor \U$2257 ( \3104 , \3058 , \3060 );
xor \U$2258 ( \3105 , \3104 , \3063 );
and \U$2259 ( \3106 , \3102 , \3105 );
and \U$2260 ( \3107 , \3088 , \3105 );
or \U$2261 ( \3108 , \3103 , \3106 , \3107 );
and \U$2262 ( \3109 , \3085 , \3108 );
xor \U$2263 ( \3110 , \3085 , \3108 );
xor \U$2264 ( \3111 , \3088 , \3102 );
xor \U$2265 ( \3112 , \3111 , \3105 );
xor \U$2266 ( \3113 , \3095 , \3097 );
xor \U$2267 ( \3114 , \3113 , \3099 );
and \U$2268 ( \3115 , \2128 , \2212 );
and \U$2269 ( \3116 , \1966 , \2336 );
and \U$2270 ( \3117 , \3115 , \3116 );
and \U$2271 ( \3118 , \1989 , \2460 );
and \U$2272 ( \3119 , \3116 , \3118 );
and \U$2273 ( \3120 , \3115 , \3118 );
or \U$2274 ( \3121 , \3117 , \3119 , \3120 );
and \U$2275 ( \3122 , \1769 , \2460 );
and \U$2276 ( \3123 , \3121 , \3122 );
xor \U$2277 ( \3124 , \3089 , \3090 );
xor \U$2278 ( \3125 , \3124 , \3092 );
and \U$2279 ( \3126 , \3122 , \3125 );
and \U$2280 ( \3127 , \3121 , \3125 );
or \U$2281 ( \3128 , \3123 , \3126 , \3127 );
and \U$2282 ( \3129 , \3114 , \3128 );
xor \U$2283 ( \3130 , \3114 , \3128 );
xor \U$2284 ( \3131 , \3121 , \3122 );
xor \U$2285 ( \3132 , \3131 , \3125 );
xor \U$2286 ( \3133 , \3115 , \3116 );
xor \U$2287 ( \3134 , \3133 , \3118 );
and \U$2288 ( \3135 , \2128 , \2336 );
and \U$2289 ( \3136 , \1966 , \2460 );
and \U$2290 ( \3137 , \3135 , \3136 );
and \U$2291 ( \3138 , \3134 , \3137 );
and \U$2292 ( \3139 , \3132 , \3138 );
and \U$2293 ( \3140 , \3130 , \3139 );
or \U$2294 ( \3141 , \3129 , \3140 );
and \U$2295 ( \3142 , \3112 , \3141 );
and \U$2296 ( \3143 , \3110 , \3142 );
or \U$2297 ( \3144 , \3109 , \3143 );
and \U$2298 ( \3145 , \3083 , \3144 );
and \U$2299 ( \3146 , \3081 , \3145 );
or \U$2300 ( \3147 , \3080 , \3146 );
and \U$2301 ( \3148 , \3040 , \3147 );
or \U$2302 ( \3149 , \3039 , \3148 );
and \U$2303 ( \3150 , \2999 , \3149 );
and \U$2304 ( \3151 , \2997 , \3150 );
or \U$2305 ( \3152 , \2996 , \3151 );
and \U$2306 ( \3153 , \2939 , \3152 );
or \U$2307 ( \3154 , \2938 , \3153 );
and \U$2308 ( \3155 , \2877 , \3154 );
or \U$2309 ( \3156 , \2876 , \3155 );
and \U$2310 ( \3157 , \2815 , \3156 );
or \U$2311 ( \3158 , \2814 , \3157 );
and \U$2312 ( \3159 , \2742 , \3158 );
and \U$2313 ( \3160 , \2740 , \3159 );
or \U$2314 ( \3161 , \2739 , \3160 );
and \U$2315 ( \3162 , \2650 , \3161 );
or \U$2316 ( \3163 , \2649 , \3162 );
and \U$2317 ( \3164 , \2548 , \3163 );
or \U$2318 ( \3165 , \2547 , \3164 );
and \U$2319 ( \3166 , \2424 , \3165 );
or \U$2320 ( \3167 , \2423 , \3166 );
and \U$2321 ( \3168 , \2300 , \3167 );
or \U$2322 ( \3169 , \2299 , \3168 );
and \U$2323 ( \3170 , \2176 , \3169 );
or \U$2324 ( \3171 , \2175 , \3170 );
and \U$2325 ( \3172 , \2031 , \3171 );
or \U$2326 ( \3173 , \2030 , \3172 );
and \U$2327 ( \3174 , \1869 , \3173 );
or \U$2328 ( \3175 , \1868 , \3174 );
and \U$2329 ( \3176 , \1743 , \3175 );
or \U$2330 ( \3177 , \1742 , \3176 );
and \U$2331 ( \3178 , \1600 , \3177 );
or \U$2332 ( \3179 , \1599 , \3178 );
and \U$2333 ( \3180 , \1514 , \3179 );
or \U$2334 ( \3181 , \1513 , \3180 );
and \U$2335 ( \3182 , \1407 , \3181 );
or \U$2336 ( \3183 , \1406 , \3182 );
and \U$2337 ( \3184 , \1290 , \3183 );
or \U$2338 ( \3185 , \1289 , \3184 );
and \U$2339 ( \3186 , \1225 , \3185 );
or \U$2340 ( \3187 , \1224 , \3186 );
and \U$2341 ( \3188 , \1139 , \3187 );
or \U$2342 ( \3189 , \1138 , \3188 );
xor \U$2343 ( \3190 , \990 , \3189 );
buf gcb0_GF_PartitionCandidate( \3191_nGcb0 , \3190 );
buf \U$2344 ( \3192 , \3191_nGcb0 );
xor \U$2345 ( \3193 , \1139 , \3187 );
buf gcb3_GF_PartitionCandidate( \3194_nGcb3 , \3193 );
buf \U$2346 ( \3195 , \3194_nGcb3 );
xor \U$2347 ( \3196 , \1225 , \3185 );
buf gcb6_GF_PartitionCandidate( \3197_nGcb6 , \3196 );
buf \U$2348 ( \3198 , \3197_nGcb6 );
xor \U$2349 ( \3199 , \1290 , \3183 );
buf gcb9_GF_PartitionCandidate( \3200_nGcb9 , \3199 );
buf \U$2350 ( \3201 , \3200_nGcb9 );
xor \U$2351 ( \3202 , \1407 , \3181 );
buf gcbc_GF_PartitionCandidate( \3203_nGcbc , \3202 );
buf \U$2352 ( \3204 , \3203_nGcbc );
xor \U$2353 ( \3205 , \1514 , \3179 );
buf gcbf_GF_PartitionCandidate( \3206_nGcbf , \3205 );
buf \U$2354 ( \3207 , \3206_nGcbf );
xor \U$2355 ( \3208 , \1600 , \3177 );
buf gcc2_GF_PartitionCandidate( \3209_nGcc2 , \3208 );
buf \U$2356 ( \3210 , \3209_nGcc2 );
xor \U$2357 ( \3211 , \1743 , \3175 );
buf gcc5_GF_PartitionCandidate( \3212_nGcc5 , \3211 );
buf \U$2358 ( \3213 , \3212_nGcc5 );
xor \U$2359 ( \3214 , \1869 , \3173 );
buf gcc8_GF_PartitionCandidate( \3215_nGcc8 , \3214 );
buf \U$2360 ( \3216 , \3215_nGcc8 );
xor \U$2361 ( \3217 , \2031 , \3171 );
buf gccb_GF_PartitionCandidate( \3218_nGccb , \3217 );
buf \U$2362 ( \3219 , \3218_nGccb );
xor \U$2363 ( \3220 , \2176 , \3169 );
buf gcce_GF_PartitionCandidate( \3221_nGcce , \3220 );
buf \U$2364 ( \3222 , \3221_nGcce );
xor \U$2365 ( \3223 , \2300 , \3167 );
buf gcd1_GF_PartitionCandidate( \3224_nGcd1 , \3223 );
buf \U$2366 ( \3225 , \3224_nGcd1 );
xor \U$2367 ( \3226 , \2424 , \3165 );
buf gcd4_GF_PartitionCandidate( \3227_nGcd4 , \3226 );
buf \U$2368 ( \3228 , \3227_nGcd4 );
xor \U$2369 ( \3229 , \2548 , \3163 );
buf gcd7_GF_PartitionCandidate( \3230_nGcd7 , \3229 );
buf \U$2370 ( \3231 , \3230_nGcd7 );
xor \U$2371 ( \3232 , \2650 , \3161 );
buf gcda_GF_PartitionCandidate( \3233_nGcda , \3232 );
buf \U$2372 ( \3234 , \3233_nGcda );
xor \U$2373 ( \3235 , \2740 , \3159 );
buf gcdd_GF_PartitionCandidate( \3236_nGcdd , \3235 );
buf \U$2374 ( \3237 , \3236_nGcdd );
xor \U$2375 ( \3238 , \2742 , \3158 );
buf gce0_GF_PartitionCandidate( \3239_nGce0 , \3238 );
buf \U$2376 ( \3240 , \3239_nGce0 );
nor \U$2377 ( \3241 , \817 , \818 , \819 , \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2378 ( \3242 , RI9157ea0_753, \3241 );
nor \U$2379 ( \3243 , RI91589e0_777, \818 , \819 , \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2380 ( \3244 , RI9157720_737, \3243 );
nor \U$2381 ( \3245 , \817 , RI9158968_776, \819 , \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2382 ( \3246 , RI9156fa0_721, \3245 );
nor \U$2383 ( \3247 , RI91589e0_777, RI9158968_776, \819 , \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2384 ( \3248 , RI9156820_705, \3247 );
nor \U$2385 ( \3249 , \817 , \818 , RI91588f0_775, \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2386 ( \3250 , RI91560a0_689, \3249 );
nor \U$2387 ( \3251 , RI91589e0_777, \818 , RI91588f0_775, \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2388 ( \3252 , RI9155920_673, \3251 );
nor \U$2389 ( \3253 , \817 , RI9158968_776, RI91588f0_775, \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2390 ( \3254 , RI91551a0_657, \3253 );
nor \U$2391 ( \3255 , RI91589e0_777, RI9158968_776, RI91588f0_775, \820 , RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2392 ( \3256 , RI9154a20_641, \3255 );
nor \U$2393 ( \3257 , \817 , \818 , \819 , RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2394 ( \3258 , RI91542a0_625, \3257 );
nor \U$2395 ( \3259 , RI91589e0_777, \818 , \819 , RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2396 ( \3260 , RI9153b20_609, \3259 );
nor \U$2397 ( \3261 , \817 , RI9158968_776, \819 , RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2398 ( \3262 , RI91533a0_593, \3261 );
nor \U$2399 ( \3263 , RI91589e0_777, RI9158968_776, \819 , RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2400 ( \3264 , RI9152c20_577, \3263 );
nor \U$2401 ( \3265 , \817 , \818 , RI91588f0_775, RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2402 ( \3266 , RI91524a0_561, \3265 );
nor \U$2403 ( \3267 , RI91589e0_777, \818 , RI91588f0_775, RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2404 ( \3268 , RI9151d20_545, \3267 );
nor \U$2405 ( \3269 , \817 , RI9158968_776, RI91588f0_775, RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2406 ( \3270 , RI91515a0_529, \3269 );
nor \U$2407 ( \3271 , RI91589e0_777, RI9158968_776, RI91588f0_775, RI9158878_774, RI9158800_773, RI9158788_772, RI9158710_771, RI9158698_770, RI9158620_769);
and \U$2408 ( \3272 , RI9150e20_513, \3271 );
or \U$2409 ( \3273 , \3242 , \3244 , \3246 , \3248 , \3250 , \3252 , \3254 , \3256 , \3258 , \3260 , \3262 , \3264 , \3266 , \3268 , \3270 , \3272 );
buf \U$2410 ( \3274 , RI9158800_773);
buf \U$2411 ( \3275 , RI9158788_772);
buf \U$2412 ( \3276 , RI9158710_771);
buf \U$2413 ( \3277 , RI9158698_770);
buf \U$2414 ( \3278 , RI9158620_769);
or \U$2415 ( \3279 , \3274 , \3275 , \3276 , \3277 , \3278 );
buf \U$2416 ( \3280 , \3279 );
_DC gd37 ( \3281_nGd37 , \3273 , \3280 );
buf \U$2417 ( \3282 , \3281_nGd37 );
and \U$2418 ( \3283 , \3240 , \3282 );
xor \U$2419 ( \3284 , \2815 , \3156 );
buf gce3_GF_PartitionCandidate( \3285_nGce3 , \3284 );
buf \U$2420 ( \3286 , \3285_nGce3 );
and \U$2421 ( \3287 , RI9157f18_754, \3241 );
and \U$2422 ( \3288 , RI9157798_738, \3243 );
and \U$2423 ( \3289 , RI9157018_722, \3245 );
and \U$2424 ( \3290 , RI9156898_706, \3247 );
and \U$2425 ( \3291 , RI9156118_690, \3249 );
and \U$2426 ( \3292 , RI9155998_674, \3251 );
and \U$2427 ( \3293 , RI9155218_658, \3253 );
and \U$2428 ( \3294 , RI9154a98_642, \3255 );
and \U$2429 ( \3295 , RI9154318_626, \3257 );
and \U$2430 ( \3296 , RI9153b98_610, \3259 );
and \U$2431 ( \3297 , RI9153418_594, \3261 );
and \U$2432 ( \3298 , RI9152c98_578, \3263 );
and \U$2433 ( \3299 , RI9152518_562, \3265 );
and \U$2434 ( \3300 , RI9151d98_546, \3267 );
and \U$2435 ( \3301 , RI9151618_530, \3269 );
and \U$2436 ( \3302 , RI9150e98_514, \3271 );
or \U$2437 ( \3303 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 );
_DC gd4a ( \3304_nGd4a , \3303 , \3280 );
buf \U$2438 ( \3305 , \3304_nGd4a );
and \U$2439 ( \3306 , \3286 , \3305 );
xor \U$2440 ( \3307 , \2877 , \3154 );
buf gce6_GF_PartitionCandidate( \3308_nGce6 , \3307 );
buf \U$2441 ( \3309 , \3308_nGce6 );
and \U$2442 ( \3310 , RI9157f90_755, \3241 );
and \U$2443 ( \3311 , RI9157810_739, \3243 );
and \U$2444 ( \3312 , RI9157090_723, \3245 );
and \U$2445 ( \3313 , RI9156910_707, \3247 );
and \U$2446 ( \3314 , RI9156190_691, \3249 );
and \U$2447 ( \3315 , RI9155a10_675, \3251 );
and \U$2448 ( \3316 , RI9155290_659, \3253 );
and \U$2449 ( \3317 , RI9154b10_643, \3255 );
and \U$2450 ( \3318 , RI9154390_627, \3257 );
and \U$2451 ( \3319 , RI9153c10_611, \3259 );
and \U$2452 ( \3320 , RI9153490_595, \3261 );
and \U$2453 ( \3321 , RI9152d10_579, \3263 );
and \U$2454 ( \3322 , RI9152590_563, \3265 );
and \U$2455 ( \3323 , RI9151e10_547, \3267 );
and \U$2456 ( \3324 , RI9151690_531, \3269 );
and \U$2457 ( \3325 , RI9150f10_515, \3271 );
or \U$2458 ( \3326 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 );
_DC gd5d ( \3327_nGd5d , \3326 , \3280 );
buf \U$2459 ( \3328 , \3327_nGd5d );
and \U$2460 ( \3329 , \3309 , \3328 );
xor \U$2461 ( \3330 , \2939 , \3152 );
buf gce9_GF_PartitionCandidate( \3331_nGce9 , \3330 );
buf \U$2462 ( \3332 , \3331_nGce9 );
and \U$2463 ( \3333 , RI9158008_756, \3241 );
and \U$2464 ( \3334 , RI9157888_740, \3243 );
and \U$2465 ( \3335 , RI9157108_724, \3245 );
and \U$2466 ( \3336 , RI9156988_708, \3247 );
and \U$2467 ( \3337 , RI9156208_692, \3249 );
and \U$2468 ( \3338 , RI9155a88_676, \3251 );
and \U$2469 ( \3339 , RI9155308_660, \3253 );
and \U$2470 ( \3340 , RI9154b88_644, \3255 );
and \U$2471 ( \3341 , RI9154408_628, \3257 );
and \U$2472 ( \3342 , RI9153c88_612, \3259 );
and \U$2473 ( \3343 , RI9153508_596, \3261 );
and \U$2474 ( \3344 , RI9152d88_580, \3263 );
and \U$2475 ( \3345 , RI9152608_564, \3265 );
and \U$2476 ( \3346 , RI9151e88_548, \3267 );
and \U$2477 ( \3347 , RI9151708_532, \3269 );
and \U$2478 ( \3348 , RI9150f88_516, \3271 );
or \U$2479 ( \3349 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 );
_DC gd70 ( \3350_nGd70 , \3349 , \3280 );
buf \U$2480 ( \3351 , \3350_nGd70 );
and \U$2481 ( \3352 , \3332 , \3351 );
xor \U$2482 ( \3353 , \2997 , \3150 );
buf gcec_GF_PartitionCandidate( \3354_nGcec , \3353 );
buf \U$2483 ( \3355 , \3354_nGcec );
and \U$2484 ( \3356 , RI9158080_757, \3241 );
and \U$2485 ( \3357 , RI9157900_741, \3243 );
and \U$2486 ( \3358 , RI9157180_725, \3245 );
and \U$2487 ( \3359 , RI9156a00_709, \3247 );
and \U$2488 ( \3360 , RI9156280_693, \3249 );
and \U$2489 ( \3361 , RI9155b00_677, \3251 );
and \U$2490 ( \3362 , RI9155380_661, \3253 );
and \U$2491 ( \3363 , RI9154c00_645, \3255 );
and \U$2492 ( \3364 , RI9154480_629, \3257 );
and \U$2493 ( \3365 , RI9153d00_613, \3259 );
and \U$2494 ( \3366 , RI9153580_597, \3261 );
and \U$2495 ( \3367 , RI9152e00_581, \3263 );
and \U$2496 ( \3368 , RI9152680_565, \3265 );
and \U$2497 ( \3369 , RI9151f00_549, \3267 );
and \U$2498 ( \3370 , RI9151780_533, \3269 );
and \U$2499 ( \3371 , RI9151000_517, \3271 );
or \U$2500 ( \3372 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 );
_DC gd83 ( \3373_nGd83 , \3372 , \3280 );
buf \U$2501 ( \3374 , \3373_nGd83 );
and \U$2502 ( \3375 , \3355 , \3374 );
xor \U$2503 ( \3376 , \2999 , \3149 );
buf gcef_GF_PartitionCandidate( \3377_nGcef , \3376 );
buf \U$2504 ( \3378 , \3377_nGcef );
and \U$2505 ( \3379 , RI91580f8_758, \3241 );
and \U$2506 ( \3380 , RI9157978_742, \3243 );
and \U$2507 ( \3381 , RI91571f8_726, \3245 );
and \U$2508 ( \3382 , RI9156a78_710, \3247 );
and \U$2509 ( \3383 , RI91562f8_694, \3249 );
and \U$2510 ( \3384 , RI9155b78_678, \3251 );
and \U$2511 ( \3385 , RI91553f8_662, \3253 );
and \U$2512 ( \3386 , RI9154c78_646, \3255 );
and \U$2513 ( \3387 , RI91544f8_630, \3257 );
and \U$2514 ( \3388 , RI9153d78_614, \3259 );
and \U$2515 ( \3389 , RI91535f8_598, \3261 );
and \U$2516 ( \3390 , RI9152e78_582, \3263 );
and \U$2517 ( \3391 , RI91526f8_566, \3265 );
and \U$2518 ( \3392 , RI9151f78_550, \3267 );
and \U$2519 ( \3393 , RI91517f8_534, \3269 );
and \U$2520 ( \3394 , RI9151078_518, \3271 );
or \U$2521 ( \3395 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 );
_DC gd96 ( \3396_nGd96 , \3395 , \3280 );
buf \U$2522 ( \3397 , \3396_nGd96 );
and \U$2523 ( \3398 , \3378 , \3397 );
xor \U$2524 ( \3399 , \3040 , \3147 );
buf gcf2_GF_PartitionCandidate( \3400_nGcf2 , \3399 );
buf \U$2525 ( \3401 , \3400_nGcf2 );
and \U$2526 ( \3402 , RI9158170_759, \3241 );
and \U$2527 ( \3403 , RI91579f0_743, \3243 );
and \U$2528 ( \3404 , RI9157270_727, \3245 );
and \U$2529 ( \3405 , RI9156af0_711, \3247 );
and \U$2530 ( \3406 , RI9156370_695, \3249 );
and \U$2531 ( \3407 , RI9155bf0_679, \3251 );
and \U$2532 ( \3408 , RI9155470_663, \3253 );
and \U$2533 ( \3409 , RI9154cf0_647, \3255 );
and \U$2534 ( \3410 , RI9154570_631, \3257 );
and \U$2535 ( \3411 , RI9153df0_615, \3259 );
and \U$2536 ( \3412 , RI9153670_599, \3261 );
and \U$2537 ( \3413 , RI9152ef0_583, \3263 );
and \U$2538 ( \3414 , RI9152770_567, \3265 );
and \U$2539 ( \3415 , RI9151ff0_551, \3267 );
and \U$2540 ( \3416 , RI9151870_535, \3269 );
and \U$2541 ( \3417 , RI91510f0_519, \3271 );
or \U$2542 ( \3418 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 );
_DC gda9 ( \3419_nGda9 , \3418 , \3280 );
buf \U$2543 ( \3420 , \3419_nGda9 );
and \U$2544 ( \3421 , \3401 , \3420 );
xor \U$2545 ( \3422 , \3081 , \3145 );
buf gcf5_GF_PartitionCandidate( \3423_nGcf5 , \3422 );
buf \U$2546 ( \3424 , \3423_nGcf5 );
and \U$2547 ( \3425 , RI91581e8_760, \3241 );
and \U$2548 ( \3426 , RI9157a68_744, \3243 );
and \U$2549 ( \3427 , RI91572e8_728, \3245 );
and \U$2550 ( \3428 , RI9156b68_712, \3247 );
and \U$2551 ( \3429 , RI91563e8_696, \3249 );
and \U$2552 ( \3430 , RI9155c68_680, \3251 );
and \U$2553 ( \3431 , RI91554e8_664, \3253 );
and \U$2554 ( \3432 , RI9154d68_648, \3255 );
and \U$2555 ( \3433 , RI91545e8_632, \3257 );
and \U$2556 ( \3434 , RI9153e68_616, \3259 );
and \U$2557 ( \3435 , RI91536e8_600, \3261 );
and \U$2558 ( \3436 , RI9152f68_584, \3263 );
and \U$2559 ( \3437 , RI91527e8_568, \3265 );
and \U$2560 ( \3438 , RI9152068_552, \3267 );
and \U$2561 ( \3439 , RI91518e8_536, \3269 );
and \U$2562 ( \3440 , RI9151168_520, \3271 );
or \U$2563 ( \3441 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 );
_DC gdbc ( \3442_nGdbc , \3441 , \3280 );
buf \U$2564 ( \3443 , \3442_nGdbc );
and \U$2565 ( \3444 , \3424 , \3443 );
xor \U$2566 ( \3445 , \3083 , \3144 );
buf gcf8_GF_PartitionCandidate( \3446_nGcf8 , \3445 );
buf \U$2567 ( \3447 , \3446_nGcf8 );
and \U$2568 ( \3448 , RI9158260_761, \3241 );
and \U$2569 ( \3449 , RI9157ae0_745, \3243 );
and \U$2570 ( \3450 , RI9157360_729, \3245 );
and \U$2571 ( \3451 , RI9156be0_713, \3247 );
and \U$2572 ( \3452 , RI9156460_697, \3249 );
and \U$2573 ( \3453 , RI9155ce0_681, \3251 );
and \U$2574 ( \3454 , RI9155560_665, \3253 );
and \U$2575 ( \3455 , RI9154de0_649, \3255 );
and \U$2576 ( \3456 , RI9154660_633, \3257 );
and \U$2577 ( \3457 , RI9153ee0_617, \3259 );
and \U$2578 ( \3458 , RI9153760_601, \3261 );
and \U$2579 ( \3459 , RI9152fe0_585, \3263 );
and \U$2580 ( \3460 , RI9152860_569, \3265 );
and \U$2581 ( \3461 , RI91520e0_553, \3267 );
and \U$2582 ( \3462 , RI9151960_537, \3269 );
and \U$2583 ( \3463 , RI91511e0_521, \3271 );
or \U$2584 ( \3464 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 );
_DC gdcf ( \3465_nGdcf , \3464 , \3280 );
buf \U$2585 ( \3466 , \3465_nGdcf );
and \U$2586 ( \3467 , \3447 , \3466 );
xor \U$2587 ( \3468 , \3110 , \3142 );
buf gcfb_GF_PartitionCandidate( \3469_nGcfb , \3468 );
buf \U$2588 ( \3470 , \3469_nGcfb );
and \U$2589 ( \3471 , RI91582d8_762, \3241 );
and \U$2590 ( \3472 , RI9157b58_746, \3243 );
and \U$2591 ( \3473 , RI91573d8_730, \3245 );
and \U$2592 ( \3474 , RI9156c58_714, \3247 );
and \U$2593 ( \3475 , RI91564d8_698, \3249 );
and \U$2594 ( \3476 , RI9155d58_682, \3251 );
and \U$2595 ( \3477 , RI91555d8_666, \3253 );
and \U$2596 ( \3478 , RI9154e58_650, \3255 );
and \U$2597 ( \3479 , RI91546d8_634, \3257 );
and \U$2598 ( \3480 , RI9153f58_618, \3259 );
and \U$2599 ( \3481 , RI91537d8_602, \3261 );
and \U$2600 ( \3482 , RI9153058_586, \3263 );
and \U$2601 ( \3483 , RI91528d8_570, \3265 );
and \U$2602 ( \3484 , RI9152158_554, \3267 );
and \U$2603 ( \3485 , RI91519d8_538, \3269 );
and \U$2604 ( \3486 , RI9151258_522, \3271 );
or \U$2605 ( \3487 , \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 , \3486 );
_DC gde2 ( \3488_nGde2 , \3487 , \3280 );
buf \U$2606 ( \3489 , \3488_nGde2 );
and \U$2607 ( \3490 , \3470 , \3489 );
xor \U$2608 ( \3491 , \3112 , \3141 );
buf gcfe_GF_PartitionCandidate( \3492_nGcfe , \3491 );
buf \U$2609 ( \3493 , \3492_nGcfe );
and \U$2610 ( \3494 , RI9158350_763, \3241 );
and \U$2611 ( \3495 , RI9157bd0_747, \3243 );
and \U$2612 ( \3496 , RI9157450_731, \3245 );
and \U$2613 ( \3497 , RI9156cd0_715, \3247 );
and \U$2614 ( \3498 , RI9156550_699, \3249 );
and \U$2615 ( \3499 , RI9155dd0_683, \3251 );
and \U$2616 ( \3500 , RI9155650_667, \3253 );
and \U$2617 ( \3501 , RI9154ed0_651, \3255 );
and \U$2618 ( \3502 , RI9154750_635, \3257 );
and \U$2619 ( \3503 , RI9153fd0_619, \3259 );
and \U$2620 ( \3504 , RI9153850_603, \3261 );
and \U$2621 ( \3505 , RI91530d0_587, \3263 );
and \U$2622 ( \3506 , RI9152950_571, \3265 );
and \U$2623 ( \3507 , RI91521d0_555, \3267 );
and \U$2624 ( \3508 , RI9151a50_539, \3269 );
and \U$2625 ( \3509 , RI91512d0_523, \3271 );
or \U$2626 ( \3510 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 );
_DC gdf5 ( \3511_nGdf5 , \3510 , \3280 );
buf \U$2627 ( \3512 , \3511_nGdf5 );
and \U$2628 ( \3513 , \3493 , \3512 );
xor \U$2629 ( \3514 , \3130 , \3139 );
buf gd01_GF_PartitionCandidate( \3515_nGd01 , \3514 );
buf \U$2630 ( \3516 , \3515_nGd01 );
and \U$2631 ( \3517 , RI91583c8_764, \3241 );
and \U$2632 ( \3518 , RI9157c48_748, \3243 );
and \U$2633 ( \3519 , RI91574c8_732, \3245 );
and \U$2634 ( \3520 , RI9156d48_716, \3247 );
and \U$2635 ( \3521 , RI91565c8_700, \3249 );
and \U$2636 ( \3522 , RI9155e48_684, \3251 );
and \U$2637 ( \3523 , RI91556c8_668, \3253 );
and \U$2638 ( \3524 , RI9154f48_652, \3255 );
and \U$2639 ( \3525 , RI91547c8_636, \3257 );
and \U$2640 ( \3526 , RI9154048_620, \3259 );
and \U$2641 ( \3527 , RI91538c8_604, \3261 );
and \U$2642 ( \3528 , RI9153148_588, \3263 );
and \U$2643 ( \3529 , RI91529c8_572, \3265 );
and \U$2644 ( \3530 , RI9152248_556, \3267 );
and \U$2645 ( \3531 , RI9151ac8_540, \3269 );
and \U$2646 ( \3532 , RI9151348_524, \3271 );
or \U$2647 ( \3533 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 );
_DC ge08 ( \3534_nGe08 , \3533 , \3280 );
buf \U$2648 ( \3535 , \3534_nGe08 );
and \U$2649 ( \3536 , \3516 , \3535 );
xor \U$2650 ( \3537 , \3132 , \3138 );
buf gd04_GF_PartitionCandidate( \3538_nGd04 , \3537 );
buf \U$2651 ( \3539 , \3538_nGd04 );
and \U$2652 ( \3540 , RI9158440_765, \3241 );
and \U$2653 ( \3541 , RI9157cc0_749, \3243 );
and \U$2654 ( \3542 , RI9157540_733, \3245 );
and \U$2655 ( \3543 , RI9156dc0_717, \3247 );
and \U$2656 ( \3544 , RI9156640_701, \3249 );
and \U$2657 ( \3545 , RI9155ec0_685, \3251 );
and \U$2658 ( \3546 , RI9155740_669, \3253 );
and \U$2659 ( \3547 , RI9154fc0_653, \3255 );
and \U$2660 ( \3548 , RI9154840_637, \3257 );
and \U$2661 ( \3549 , RI91540c0_621, \3259 );
and \U$2662 ( \3550 , RI9153940_605, \3261 );
and \U$2663 ( \3551 , RI91531c0_589, \3263 );
and \U$2664 ( \3552 , RI9152a40_573, \3265 );
and \U$2665 ( \3553 , RI91522c0_557, \3267 );
and \U$2666 ( \3554 , RI9151b40_541, \3269 );
and \U$2667 ( \3555 , RI91513c0_525, \3271 );
or \U$2668 ( \3556 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 );
_DC ge1b ( \3557_nGe1b , \3556 , \3280 );
buf \U$2669 ( \3558 , \3557_nGe1b );
and \U$2670 ( \3559 , \3539 , \3558 );
xor \U$2671 ( \3560 , \3134 , \3137 );
buf gd07_GF_PartitionCandidate( \3561_nGd07 , \3560 );
buf \U$2672 ( \3562 , \3561_nGd07 );
and \U$2673 ( \3563 , RI91584b8_766, \3241 );
and \U$2674 ( \3564 , RI9157d38_750, \3243 );
and \U$2675 ( \3565 , RI91575b8_734, \3245 );
and \U$2676 ( \3566 , RI9156e38_718, \3247 );
and \U$2677 ( \3567 , RI91566b8_702, \3249 );
and \U$2678 ( \3568 , RI9155f38_686, \3251 );
and \U$2679 ( \3569 , RI91557b8_670, \3253 );
and \U$2680 ( \3570 , RI9155038_654, \3255 );
and \U$2681 ( \3571 , RI91548b8_638, \3257 );
and \U$2682 ( \3572 , RI9154138_622, \3259 );
and \U$2683 ( \3573 , RI91539b8_606, \3261 );
and \U$2684 ( \3574 , RI9153238_590, \3263 );
and \U$2685 ( \3575 , RI9152ab8_574, \3265 );
and \U$2686 ( \3576 , RI9152338_558, \3267 );
and \U$2687 ( \3577 , RI9151bb8_542, \3269 );
and \U$2688 ( \3578 , RI9151438_526, \3271 );
or \U$2689 ( \3579 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 );
_DC ge2e ( \3580_nGe2e , \3579 , \3280 );
buf \U$2690 ( \3581 , \3580_nGe2e );
and \U$2691 ( \3582 , \3562 , \3581 );
xor \U$2692 ( \3583 , \3135 , \3136 );
buf gd0a_GF_PartitionCandidate( \3584_nGd0a , \3583 );
buf \U$2693 ( \3585 , \3584_nGd0a );
and \U$2694 ( \3586 , RI9158530_767, \3241 );
and \U$2695 ( \3587 , RI9157db0_751, \3243 );
and \U$2696 ( \3588 , RI9157630_735, \3245 );
and \U$2697 ( \3589 , RI9156eb0_719, \3247 );
and \U$2698 ( \3590 , RI9156730_703, \3249 );
and \U$2699 ( \3591 , RI9155fb0_687, \3251 );
and \U$2700 ( \3592 , RI9155830_671, \3253 );
and \U$2701 ( \3593 , RI91550b0_655, \3255 );
and \U$2702 ( \3594 , RI9154930_639, \3257 );
and \U$2703 ( \3595 , RI91541b0_623, \3259 );
and \U$2704 ( \3596 , RI9153a30_607, \3261 );
and \U$2705 ( \3597 , RI91532b0_591, \3263 );
and \U$2706 ( \3598 , RI9152b30_575, \3265 );
and \U$2707 ( \3599 , RI91523b0_559, \3267 );
and \U$2708 ( \3600 , RI9151c30_543, \3269 );
and \U$2709 ( \3601 , RI91514b0_527, \3271 );
or \U$2710 ( \3602 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 );
_DC ge41 ( \3603_nGe41 , \3602 , \3280 );
buf \U$2711 ( \3604 , \3603_nGe41 );
and \U$2712 ( \3605 , \3585 , \3604 );
and \U$2713 ( \3606 , \2128 , \2460 );
buf gd0d_GF_PartitionCandidate( \3607_nGd0d , \3606 );
buf \U$2714 ( \3608 , \3607_nGd0d );
and \U$2715 ( \3609 , RI91585a8_768, \3241 );
and \U$2716 ( \3610 , RI9157e28_752, \3243 );
and \U$2717 ( \3611 , RI91576a8_736, \3245 );
and \U$2718 ( \3612 , RI9156f28_720, \3247 );
and \U$2719 ( \3613 , RI91567a8_704, \3249 );
and \U$2720 ( \3614 , RI9156028_688, \3251 );
and \U$2721 ( \3615 , RI91558a8_672, \3253 );
and \U$2722 ( \3616 , RI9155128_656, \3255 );
and \U$2723 ( \3617 , RI91549a8_640, \3257 );
and \U$2724 ( \3618 , RI9154228_624, \3259 );
and \U$2725 ( \3619 , RI9153aa8_608, \3261 );
and \U$2726 ( \3620 , RI9153328_592, \3263 );
and \U$2727 ( \3621 , RI9152ba8_576, \3265 );
and \U$2728 ( \3622 , RI9152428_560, \3267 );
and \U$2729 ( \3623 , RI9151ca8_544, \3269 );
and \U$2730 ( \3624 , RI9151528_528, \3271 );
or \U$2731 ( \3625 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 );
_DC ge54 ( \3626_nGe54 , \3625 , \3280 );
buf \U$2732 ( \3627 , \3626_nGe54 );
and \U$2733 ( \3628 , \3608 , \3627 );
and \U$2734 ( \3629 , \3604 , \3628 );
and \U$2735 ( \3630 , \3585 , \3628 );
or \U$2736 ( \3631 , \3605 , \3629 , \3630 );
and \U$2737 ( \3632 , \3581 , \3631 );
and \U$2738 ( \3633 , \3562 , \3631 );
or \U$2739 ( \3634 , \3582 , \3632 , \3633 );
and \U$2740 ( \3635 , \3558 , \3634 );
and \U$2741 ( \3636 , \3539 , \3634 );
or \U$2742 ( \3637 , \3559 , \3635 , \3636 );
and \U$2743 ( \3638 , \3535 , \3637 );
and \U$2744 ( \3639 , \3516 , \3637 );
or \U$2745 ( \3640 , \3536 , \3638 , \3639 );
and \U$2746 ( \3641 , \3512 , \3640 );
and \U$2747 ( \3642 , \3493 , \3640 );
or \U$2748 ( \3643 , \3513 , \3641 , \3642 );
and \U$2749 ( \3644 , \3489 , \3643 );
and \U$2750 ( \3645 , \3470 , \3643 );
or \U$2751 ( \3646 , \3490 , \3644 , \3645 );
and \U$2752 ( \3647 , \3466 , \3646 );
and \U$2753 ( \3648 , \3447 , \3646 );
or \U$2754 ( \3649 , \3467 , \3647 , \3648 );
and \U$2755 ( \3650 , \3443 , \3649 );
and \U$2756 ( \3651 , \3424 , \3649 );
or \U$2757 ( \3652 , \3444 , \3650 , \3651 );
and \U$2758 ( \3653 , \3420 , \3652 );
and \U$2759 ( \3654 , \3401 , \3652 );
or \U$2760 ( \3655 , \3421 , \3653 , \3654 );
and \U$2761 ( \3656 , \3397 , \3655 );
and \U$2762 ( \3657 , \3378 , \3655 );
or \U$2763 ( \3658 , \3398 , \3656 , \3657 );
and \U$2764 ( \3659 , \3374 , \3658 );
and \U$2765 ( \3660 , \3355 , \3658 );
or \U$2766 ( \3661 , \3375 , \3659 , \3660 );
and \U$2767 ( \3662 , \3351 , \3661 );
and \U$2768 ( \3663 , \3332 , \3661 );
or \U$2769 ( \3664 , \3352 , \3662 , \3663 );
and \U$2770 ( \3665 , \3328 , \3664 );
and \U$2771 ( \3666 , \3309 , \3664 );
or \U$2772 ( \3667 , \3329 , \3665 , \3666 );
and \U$2773 ( \3668 , \3305 , \3667 );
and \U$2774 ( \3669 , \3286 , \3667 );
or \U$2775 ( \3670 , \3306 , \3668 , \3669 );
and \U$2776 ( \3671 , \3282 , \3670 );
and \U$2777 ( \3672 , \3240 , \3670 );
or \U$2778 ( \3673 , \3283 , \3671 , \3672 );
and \U$2779 ( \3674 , \3237 , \3673 );
and \U$2780 ( \3675 , \3234 , \3674 );
and \U$2781 ( \3676 , \3231 , \3675 );
and \U$2782 ( \3677 , \3228 , \3676 );
and \U$2783 ( \3678 , \3225 , \3677 );
and \U$2784 ( \3679 , \3222 , \3678 );
and \U$2785 ( \3680 , \3219 , \3679 );
and \U$2786 ( \3681 , \3216 , \3680 );
and \U$2787 ( \3682 , \3213 , \3681 );
and \U$2788 ( \3683 , \3210 , \3682 );
and \U$2789 ( \3684 , \3207 , \3683 );
and \U$2790 ( \3685 , \3204 , \3684 );
and \U$2791 ( \3686 , \3201 , \3685 );
and \U$2792 ( \3687 , \3198 , \3686 );
and \U$2793 ( \3688 , \3195 , \3687 );
xor \U$2794 ( \3689 , \3192 , \3688 );
buf \U$2795 ( \3690 , \3689 );
buf \U$2796 ( \3691 , \3690 );
xor \U$2797 ( \3692 , \3195 , \3687 );
buf \U$2798 ( \3693 , \3692 );
buf \U$2799 ( \3694 , \3693 );
xor \U$2800 ( \3695 , \3198 , \3686 );
buf \U$2801 ( \3696 , \3695 );
buf \U$2802 ( \3697 , \3696 );
xor \U$2803 ( \3698 , \3201 , \3685 );
buf \U$2804 ( \3699 , \3698 );
buf \U$2805 ( \3700 , \3699 );
xor \U$2806 ( \3701 , \3204 , \3684 );
buf \U$2807 ( \3702 , \3701 );
buf \U$2808 ( \3703 , \3702 );
xor \U$2809 ( \3704 , \3207 , \3683 );
buf \U$2810 ( \3705 , \3704 );
buf \U$2811 ( \3706 , \3705 );
xor \U$2812 ( \3707 , \3210 , \3682 );
buf \U$2813 ( \3708 , \3707 );
buf \U$2814 ( \3709 , \3708 );
xor \U$2815 ( \3710 , \3213 , \3681 );
buf \U$2816 ( \3711 , \3710 );
buf \U$2817 ( \3712 , \3711 );
xor \U$2818 ( \3713 , \3216 , \3680 );
buf \U$2819 ( \3714 , \3713 );
buf \U$2820 ( \3715 , \3714 );
xor \U$2821 ( \3716 , \3219 , \3679 );
buf \U$2822 ( \3717 , \3716 );
buf \U$2823 ( \3718 , \3717 );
xor \U$2824 ( \3719 , \3222 , \3678 );
buf \U$2825 ( \3720 , \3719 );
buf \U$2826 ( \3721 , \3720 );
xor \U$2827 ( \3722 , \3225 , \3677 );
buf \U$2828 ( \3723 , \3722 );
buf \U$2829 ( \3724 , \3723 );
xor \U$2830 ( \3725 , \3228 , \3676 );
buf \U$2831 ( \3726 , \3725 );
buf \U$2832 ( \3727 , \3726 );
xor \U$2833 ( \3728 , \3231 , \3675 );
buf \U$2834 ( \3729 , \3728 );
buf \U$2835 ( \3730 , \3729 );
xor \U$2836 ( \3731 , \3234 , \3674 );
buf \U$2837 ( \3732 , \3731 );
buf \U$2838 ( \3733 , \3732 );
xor \U$2839 ( \3734 , \3237 , \3673 );
buf \U$2840 ( \3735 , \3734 );
buf \U$2841 ( \3736 , \3735 );
xor \U$2842 ( \3737 , \3240 , \3282 );
xor \U$2843 ( \3738 , \3737 , \3670 );
buf \U$2844 ( \3739 , \3738 );
buf \U$2845 ( \3740 , \3739 );
xor \U$2846 ( \3741 , \3286 , \3305 );
xor \U$2847 ( \3742 , \3741 , \3667 );
buf \U$2848 ( \3743 , \3742 );
buf \U$2849 ( \3744 , \3743 );
xor \U$2850 ( \3745 , \3309 , \3328 );
xor \U$2851 ( \3746 , \3745 , \3664 );
buf \U$2852 ( \3747 , \3746 );
buf \U$2853 ( \3748 , \3747 );
xor \U$2854 ( \3749 , \3332 , \3351 );
xor \U$2855 ( \3750 , \3749 , \3661 );
buf \U$2856 ( \3751 , \3750 );
buf \U$2857 ( \3752 , \3751 );
xor \U$2858 ( \3753 , \3355 , \3374 );
xor \U$2859 ( \3754 , \3753 , \3658 );
buf \U$2860 ( \3755 , \3754 );
buf \U$2861 ( \3756 , \3755 );
xor \U$2862 ( \3757 , \3378 , \3397 );
xor \U$2863 ( \3758 , \3757 , \3655 );
buf \U$2864 ( \3759 , \3758 );
buf \U$2865 ( \3760 , \3759 );
xor \U$2866 ( \3761 , \3401 , \3420 );
xor \U$2867 ( \3762 , \3761 , \3652 );
buf \U$2868 ( \3763 , \3762 );
buf \U$2869 ( \3764 , \3763 );
xor \U$2870 ( \3765 , \3424 , \3443 );
xor \U$2871 ( \3766 , \3765 , \3649 );
buf \U$2872 ( \3767 , \3766 );
buf \U$2873 ( \3768 , \3767 );
xor \U$2874 ( \3769 , \3447 , \3466 );
xor \U$2875 ( \3770 , \3769 , \3646 );
buf \U$2876 ( \3771 , \3770 );
buf \U$2877 ( \3772 , \3771 );
xor \U$2878 ( \3773 , \3470 , \3489 );
xor \U$2879 ( \3774 , \3773 , \3643 );
buf \U$2880 ( \3775 , \3774 );
buf \U$2881 ( \3776 , \3775 );
xor \U$2882 ( \3777 , \3493 , \3512 );
xor \U$2883 ( \3778 , \3777 , \3640 );
buf \U$2884 ( \3779 , \3778 );
buf \U$2885 ( \3780 , \3779 );
endmodule

